module fake_netlist_5_109_n_828 (n_137, n_168, n_164, n_91, n_82, n_122, n_142, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_165, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_60, n_155, n_152, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_125, n_35, n_167, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_157, n_29, n_79, n_131, n_151, n_47, n_25, n_53, n_160, n_8, n_158, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_159, n_163, n_95, n_119, n_169, n_59, n_26, n_133, n_55, n_99, n_2, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_162, n_27, n_170, n_64, n_77, n_102, n_106, n_161, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_134, n_32, n_41, n_104, n_103, n_56, n_51, n_63, n_97, n_141, n_166, n_11, n_171, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_828);

input n_137;
input n_168;
input n_164;
input n_91;
input n_82;
input n_122;
input n_142;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_165;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_60;
input n_155;
input n_152;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_125;
input n_35;
input n_167;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_157;
input n_29;
input n_79;
input n_131;
input n_151;
input n_47;
input n_25;
input n_53;
input n_160;
input n_8;
input n_158;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_159;
input n_163;
input n_95;
input n_119;
input n_169;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_162;
input n_27;
input n_170;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_134;
input n_32;
input n_41;
input n_104;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_166;
input n_11;
input n_171;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_828;

wire n_676;
wire n_294;
wire n_431;
wire n_318;
wire n_419;
wire n_380;
wire n_653;
wire n_611;
wire n_444;
wire n_642;
wire n_469;
wire n_615;
wire n_194;
wire n_316;
wire n_785;
wire n_389;
wire n_549;
wire n_684;
wire n_418;
wire n_248;
wire n_315;
wire n_268;
wire n_523;
wire n_451;
wire n_532;
wire n_705;
wire n_619;
wire n_408;
wire n_678;
wire n_664;
wire n_376;
wire n_697;
wire n_503;
wire n_235;
wire n_226;
wire n_605;
wire n_776;
wire n_667;
wire n_515;
wire n_790;
wire n_353;
wire n_351;
wire n_367;
wire n_643;
wire n_620;
wire n_452;
wire n_397;
wire n_493;
wire n_525;
wire n_703;
wire n_698;
wire n_483;
wire n_544;
wire n_683;
wire n_780;
wire n_649;
wire n_552;
wire n_547;
wire n_721;
wire n_564;
wire n_467;
wire n_802;
wire n_423;
wire n_284;
wire n_245;
wire n_501;
wire n_823;
wire n_725;
wire n_280;
wire n_744;
wire n_590;
wire n_629;
wire n_672;
wire n_378;
wire n_551;
wire n_762;
wire n_581;
wire n_688;
wire n_382;
wire n_554;
wire n_800;
wire n_254;
wire n_690;
wire n_583;
wire n_671;
wire n_718;
wire n_819;
wire n_302;
wire n_265;
wire n_526;
wire n_719;
wire n_293;
wire n_372;
wire n_443;
wire n_244;
wire n_677;
wire n_173;
wire n_821;
wire n_198;
wire n_714;
wire n_447;
wire n_247;
wire n_314;
wire n_368;
wire n_433;
wire n_604;
wire n_321;
wire n_292;
wire n_625;
wire n_621;
wire n_753;
wire n_455;
wire n_674;
wire n_417;
wire n_612;
wire n_212;
wire n_385;
wire n_516;
wire n_498;
wire n_788;
wire n_507;
wire n_497;
wire n_689;
wire n_738;
wire n_606;
wire n_559;
wire n_275;
wire n_640;
wire n_252;
wire n_624;
wire n_825;
wire n_295;
wire n_330;
wire n_508;
wire n_739;
wire n_506;
wire n_737;
wire n_610;
wire n_692;
wire n_755;
wire n_509;
wire n_568;
wire n_373;
wire n_820;
wire n_757;
wire n_307;
wire n_633;
wire n_439;
wire n_530;
wire n_556;
wire n_209;
wire n_259;
wire n_448;
wire n_758;
wire n_668;
wire n_733;
wire n_375;
wire n_301;
wire n_779;
wire n_576;
wire n_804;
wire n_186;
wire n_537;
wire n_191;
wire n_587;
wire n_659;
wire n_492;
wire n_792;
wire n_563;
wire n_756;
wire n_524;
wire n_399;
wire n_341;
wire n_204;
wire n_394;
wire n_250;
wire n_579;
wire n_741;
wire n_548;
wire n_543;
wire n_260;
wire n_812;
wire n_298;
wire n_650;
wire n_320;
wire n_694;
wire n_518;
wire n_505;
wire n_286;
wire n_282;
wire n_752;
wire n_331;
wire n_406;
wire n_519;
wire n_470;
wire n_782;
wire n_325;
wire n_449;
wire n_724;
wire n_546;
wire n_760;
wire n_658;
wire n_281;
wire n_240;
wire n_381;
wire n_189;
wire n_220;
wire n_291;
wire n_231;
wire n_257;
wire n_390;
wire n_731;
wire n_456;
wire n_371;
wire n_481;
wire n_535;
wire n_709;
wire n_540;
wire n_317;
wire n_618;
wire n_323;
wire n_569;
wire n_769;
wire n_195;
wire n_356;
wire n_227;
wire n_592;
wire n_271;
wire n_826;
wire n_335;
wire n_654;
wire n_370;
wire n_234;
wire n_343;
wire n_308;
wire n_379;
wire n_428;
wire n_267;
wire n_514;
wire n_457;
wire n_570;
wire n_297;
wire n_603;
wire n_225;
wire n_377;
wire n_751;
wire n_484;
wire n_775;
wire n_219;
wire n_442;
wire n_814;
wire n_192;
wire n_636;
wire n_786;
wire n_600;
wire n_660;
wire n_223;
wire n_392;
wire n_655;
wire n_704;
wire n_787;
wire n_264;
wire n_669;
wire n_472;
wire n_742;
wire n_750;
wire n_454;
wire n_387;
wire n_771;
wire n_374;
wire n_276;
wire n_339;
wire n_183;
wire n_185;
wire n_243;
wire n_398;
wire n_396;
wire n_635;
wire n_347;
wire n_763;
wire n_550;
wire n_522;
wire n_255;
wire n_696;
wire n_215;
wire n_350;
wire n_196;
wire n_798;
wire n_662;
wire n_459;
wire n_646;
wire n_211;
wire n_218;
wire n_400;
wire n_181;
wire n_436;
wire n_290;
wire n_580;
wire n_221;
wire n_178;
wire n_622;
wire n_723;
wire n_386;
wire n_578;
wire n_287;
wire n_344;
wire n_555;
wire n_783;
wire n_473;
wire n_422;
wire n_475;
wire n_777;
wire n_661;
wire n_682;
wire n_415;
wire n_485;
wire n_496;
wire n_355;
wire n_486;
wire n_670;
wire n_816;
wire n_336;
wire n_584;
wire n_681;
wire n_591;
wire n_521;
wire n_614;
wire n_663;
wire n_430;
wire n_337;
wire n_313;
wire n_631;
wire n_673;
wire n_479;
wire n_528;
wire n_510;
wire n_216;
wire n_680;
wire n_395;
wire n_432;
wire n_553;
wire n_727;
wire n_311;
wire n_813;
wire n_773;
wire n_208;
wire n_743;
wire n_214;
wire n_328;
wire n_801;
wire n_299;
wire n_303;
wire n_369;
wire n_675;
wire n_296;
wire n_613;
wire n_241;
wire n_637;
wire n_357;
wire n_598;
wire n_685;
wire n_608;
wire n_184;
wire n_446;
wire n_445;
wire n_749;
wire n_772;
wire n_691;
wire n_717;
wire n_468;
wire n_499;
wire n_213;
wire n_517;
wire n_342;
wire n_482;
wire n_588;
wire n_361;
wire n_464;
wire n_789;
wire n_363;
wire n_413;
wire n_402;
wire n_734;
wire n_638;
wire n_700;
wire n_197;
wire n_796;
wire n_573;
wire n_236;
wire n_388;
wire n_761;
wire n_249;
wire n_740;
wire n_304;
wire n_329;
wire n_203;
wire n_274;
wire n_577;
wire n_384;
wire n_582;
wire n_460;
wire n_277;
wire n_477;
wire n_338;
wire n_461;
wire n_333;
wire n_571;
wire n_693;
wire n_309;
wire n_512;
wire n_462;
wire n_322;
wire n_567;
wire n_258;
wire n_652;
wire n_778;
wire n_306;
wire n_722;
wire n_458;
wire n_288;
wire n_770;
wire n_188;
wire n_190;
wire n_201;
wire n_263;
wire n_471;
wire n_609;
wire n_224;
wire n_228;
wire n_283;
wire n_383;
wire n_781;
wire n_711;
wire n_474;
wire n_765;
wire n_542;
wire n_463;
wire n_488;
wire n_595;
wire n_736;
wire n_502;
wire n_239;
wire n_466;
wire n_420;
wire n_630;
wire n_489;
wire n_632;
wire n_699;
wire n_617;
wire n_310;
wire n_593;
wire n_504;
wire n_511;
wire n_748;
wire n_586;
wire n_465;
wire n_358;
wire n_362;
wire n_332;
wire n_273;
wire n_349;
wire n_585;
wire n_270;
wire n_616;
wire n_230;
wire n_601;
wire n_279;
wire n_253;
wire n_261;
wire n_174;
wire n_289;
wire n_745;
wire n_627;
wire n_767;
wire n_172;
wire n_206;
wire n_217;
wire n_440;
wire n_726;
wire n_478;
wire n_793;
wire n_545;
wire n_441;
wire n_450;
wire n_648;
wire n_312;
wire n_476;
wire n_818;
wire n_429;
wire n_534;
wire n_345;
wire n_210;
wire n_494;
wire n_641;
wire n_628;
wire n_365;
wire n_774;
wire n_730;
wire n_729;
wire n_176;
wire n_557;
wire n_182;
wire n_354;
wire n_607;
wire n_575;
wire n_480;
wire n_647;
wire n_237;
wire n_425;
wire n_513;
wire n_407;
wire n_527;
wire n_679;
wire n_795;
wire n_707;
wire n_710;
wire n_695;
wire n_180;
wire n_560;
wire n_656;
wire n_340;
wire n_207;
wire n_561;
wire n_346;
wire n_393;
wire n_229;
wire n_487;
wire n_495;
wire n_602;
wire n_665;
wire n_574;
wire n_437;
wire n_177;
wire n_403;
wire n_453;
wire n_421;
wire n_720;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_490;
wire n_805;
wire n_326;
wire n_794;
wire n_768;
wire n_233;
wire n_404;
wire n_686;
wire n_205;
wire n_366;
wire n_572;
wire n_712;
wire n_754;
wire n_815;
wire n_246;
wire n_596;
wire n_179;
wire n_410;
wire n_558;
wire n_708;
wire n_269;
wire n_529;
wire n_735;
wire n_702;
wire n_285;
wire n_822;
wire n_412;
wire n_232;
wire n_327;
wire n_657;
wire n_644;
wire n_728;
wire n_202;
wire n_266;
wire n_272;
wire n_491;
wire n_427;
wire n_791;
wire n_732;
wire n_193;
wire n_251;
wire n_352;
wire n_566;
wire n_426;
wire n_520;
wire n_565;
wire n_808;
wire n_409;
wire n_797;
wire n_589;
wire n_716;
wire n_597;
wire n_500;
wire n_562;
wire n_300;
wire n_651;
wire n_435;
wire n_809;
wire n_334;
wire n_599;
wire n_766;
wire n_811;
wire n_541;
wire n_807;
wire n_391;
wire n_701;
wire n_434;
wire n_645;
wire n_539;
wire n_175;
wire n_538;
wire n_666;
wire n_262;
wire n_803;
wire n_238;
wire n_639;
wire n_799;
wire n_687;
wire n_715;
wire n_411;
wire n_414;
wire n_319;
wire n_364;
wire n_536;
wire n_531;
wire n_242;
wire n_817;
wire n_360;
wire n_594;
wire n_764;
wire n_200;
wire n_759;
wire n_222;
wire n_438;
wire n_806;
wire n_713;
wire n_324;
wire n_810;
wire n_634;
wire n_416;
wire n_199;
wire n_827;
wire n_187;
wire n_401;
wire n_348;
wire n_626;
wire n_424;
wire n_706;
wire n_746;
wire n_256;
wire n_305;
wire n_533;
wire n_747;
wire n_278;
wire n_784;

BUFx2_ASAP7_75t_L g172 ( 
.A(n_24),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_77),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_11),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_154),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_55),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_135),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_159),
.Y(n_178)
);

INVx1_ASAP7_75t_SL g179 ( 
.A(n_101),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_113),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_28),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_74),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_168),
.Y(n_183)
);

BUFx3_ASAP7_75t_L g184 ( 
.A(n_134),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_35),
.Y(n_185)
);

CKINVDCx16_ASAP7_75t_R g186 ( 
.A(n_164),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_60),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_3),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_105),
.Y(n_189)
);

INVx1_ASAP7_75t_SL g190 ( 
.A(n_30),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_152),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_9),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_145),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_17),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g195 ( 
.A(n_8),
.Y(n_195)
);

BUFx5_ASAP7_75t_L g196 ( 
.A(n_76),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g197 ( 
.A(n_108),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_8),
.Y(n_198)
);

INVx1_ASAP7_75t_SL g199 ( 
.A(n_25),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_160),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_53),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_156),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g203 ( 
.A(n_102),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_18),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_31),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_124),
.Y(n_206)
);

CKINVDCx14_ASAP7_75t_R g207 ( 
.A(n_11),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_147),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_116),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_20),
.Y(n_210)
);

BUFx5_ASAP7_75t_L g211 ( 
.A(n_67),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_66),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_25),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_40),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_20),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_36),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_167),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_87),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_89),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_118),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_94),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_39),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_99),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_78),
.Y(n_224)
);

INVx2_ASAP7_75t_SL g225 ( 
.A(n_126),
.Y(n_225)
);

BUFx2_ASAP7_75t_L g226 ( 
.A(n_41),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_43),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_150),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_119),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_103),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_26),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_88),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_195),
.Y(n_233)
);

INVxp67_ASAP7_75t_L g234 ( 
.A(n_172),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_173),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_207),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_174),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_195),
.Y(n_238)
);

INVxp67_ASAP7_75t_L g239 ( 
.A(n_194),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_195),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_226),
.B(n_0),
.Y(n_241)
);

INVxp67_ASAP7_75t_SL g242 ( 
.A(n_184),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_204),
.Y(n_243)
);

INVx1_ASAP7_75t_SL g244 ( 
.A(n_231),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_175),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_177),
.Y(n_246)
);

HB1xp67_ASAP7_75t_L g247 ( 
.A(n_188),
.Y(n_247)
);

BUFx6f_ASAP7_75t_SL g248 ( 
.A(n_197),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_192),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_198),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_178),
.Y(n_251)
);

HB1xp67_ASAP7_75t_L g252 ( 
.A(n_210),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_182),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_183),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_180),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_185),
.Y(n_256)
);

INVxp67_ASAP7_75t_L g257 ( 
.A(n_199),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_187),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_213),
.Y(n_259)
);

CKINVDCx16_ASAP7_75t_R g260 ( 
.A(n_186),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_193),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_209),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_225),
.B(n_0),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_181),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_214),
.Y(n_265)
);

NOR2xp67_ASAP7_75t_L g266 ( 
.A(n_215),
.B(n_1),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_223),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_176),
.Y(n_268)
);

BUFx3_ASAP7_75t_L g269 ( 
.A(n_227),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_197),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_197),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_203),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_202),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_196),
.B(n_1),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_208),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_220),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_203),
.Y(n_277)
);

INVxp67_ASAP7_75t_SL g278 ( 
.A(n_203),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_189),
.Y(n_279)
);

INVx3_ASAP7_75t_L g280 ( 
.A(n_270),
.Y(n_280)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_271),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_272),
.Y(n_282)
);

HB1xp67_ASAP7_75t_L g283 ( 
.A(n_257),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_277),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_235),
.Y(n_285)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_233),
.Y(n_286)
);

INVx3_ASAP7_75t_L g287 ( 
.A(n_238),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_268),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_SL g289 ( 
.A(n_236),
.B(n_179),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_245),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_240),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_246),
.B(n_232),
.Y(n_292)
);

INVx4_ASAP7_75t_L g293 ( 
.A(n_248),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_268),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_278),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_R g296 ( 
.A(n_279),
.B(n_191),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_251),
.B(n_230),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_255),
.B(n_200),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_243),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_274),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_273),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_253),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_254),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_273),
.Y(n_304)
);

INVx3_ASAP7_75t_L g305 ( 
.A(n_269),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_264),
.B(n_229),
.Y(n_306)
);

BUFx2_ASAP7_75t_L g307 ( 
.A(n_236),
.Y(n_307)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_256),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_275),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_241),
.B(n_263),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_258),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_279),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_261),
.Y(n_313)
);

INVx3_ASAP7_75t_L g314 ( 
.A(n_269),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_237),
.Y(n_315)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_262),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_265),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_267),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_242),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_239),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_237),
.Y(n_321)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_248),
.Y(n_322)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_248),
.Y(n_323)
);

BUFx6f_ASAP7_75t_L g324 ( 
.A(n_259),
.Y(n_324)
);

AND2x2_ASAP7_75t_L g325 ( 
.A(n_247),
.B(n_190),
.Y(n_325)
);

INVx3_ASAP7_75t_L g326 ( 
.A(n_259),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_266),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_275),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_252),
.Y(n_329)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_234),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_302),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_310),
.B(n_260),
.Y(n_332)
);

AND2x2_ASAP7_75t_L g333 ( 
.A(n_283),
.B(n_244),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_302),
.Y(n_334)
);

AOI22xp5_ASAP7_75t_L g335 ( 
.A1(n_325),
.A2(n_249),
.B1(n_250),
.B2(n_218),
.Y(n_335)
);

INVx3_ASAP7_75t_L g336 ( 
.A(n_308),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_303),
.Y(n_337)
);

BUFx6f_ASAP7_75t_L g338 ( 
.A(n_308),
.Y(n_338)
);

AND2x4_ASAP7_75t_L g339 ( 
.A(n_305),
.B(n_201),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_303),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_311),
.Y(n_341)
);

INVx2_ASAP7_75t_L g342 ( 
.A(n_280),
.Y(n_342)
);

AOI22xp5_ASAP7_75t_L g343 ( 
.A1(n_325),
.A2(n_249),
.B1(n_250),
.B2(n_219),
.Y(n_343)
);

BUFx3_ASAP7_75t_L g344 ( 
.A(n_305),
.Y(n_344)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_280),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_311),
.Y(n_346)
);

AND2x2_ASAP7_75t_L g347 ( 
.A(n_330),
.B(n_276),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g348 ( 
.A(n_319),
.B(n_205),
.Y(n_348)
);

INVx6_ASAP7_75t_L g349 ( 
.A(n_293),
.Y(n_349)
);

BUFx6f_ASAP7_75t_L g350 ( 
.A(n_316),
.Y(n_350)
);

AND2x2_ASAP7_75t_L g351 ( 
.A(n_330),
.B(n_319),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_300),
.B(n_305),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_313),
.Y(n_353)
);

AND2x2_ASAP7_75t_SL g354 ( 
.A(n_324),
.B(n_196),
.Y(n_354)
);

INVx2_ASAP7_75t_L g355 ( 
.A(n_280),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_300),
.B(n_206),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_296),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_313),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_305),
.B(n_212),
.Y(n_359)
);

AND2x6_ASAP7_75t_L g360 ( 
.A(n_322),
.B(n_196),
.Y(n_360)
);

NAND2x1p5_ASAP7_75t_L g361 ( 
.A(n_324),
.B(n_326),
.Y(n_361)
);

BUFx6f_ASAP7_75t_L g362 ( 
.A(n_316),
.Y(n_362)
);

OAI21xp33_ASAP7_75t_SL g363 ( 
.A1(n_289),
.A2(n_211),
.B(n_196),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_317),
.Y(n_364)
);

HB1xp67_ASAP7_75t_L g365 ( 
.A(n_314),
.Y(n_365)
);

INVx2_ASAP7_75t_L g366 ( 
.A(n_280),
.Y(n_366)
);

INVx4_ASAP7_75t_L g367 ( 
.A(n_314),
.Y(n_367)
);

AND2x6_ASAP7_75t_L g368 ( 
.A(n_322),
.B(n_196),
.Y(n_368)
);

INVx2_ASAP7_75t_L g369 ( 
.A(n_281),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_317),
.Y(n_370)
);

NAND2x1p5_ASAP7_75t_L g371 ( 
.A(n_324),
.B(n_216),
.Y(n_371)
);

AND2x6_ASAP7_75t_L g372 ( 
.A(n_323),
.B(n_196),
.Y(n_372)
);

INVx2_ASAP7_75t_L g373 ( 
.A(n_281),
.Y(n_373)
);

CKINVDCx20_ASAP7_75t_R g374 ( 
.A(n_288),
.Y(n_374)
);

BUFx3_ASAP7_75t_L g375 ( 
.A(n_314),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_314),
.B(n_217),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_295),
.B(n_221),
.Y(n_377)
);

INVx1_ASAP7_75t_SL g378 ( 
.A(n_294),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_295),
.B(n_222),
.Y(n_379)
);

INVx2_ASAP7_75t_L g380 ( 
.A(n_286),
.Y(n_380)
);

INVx1_ASAP7_75t_SL g381 ( 
.A(n_301),
.Y(n_381)
);

BUFx3_ASAP7_75t_L g382 ( 
.A(n_323),
.Y(n_382)
);

BUFx3_ASAP7_75t_L g383 ( 
.A(n_318),
.Y(n_383)
);

INVx4_ASAP7_75t_L g384 ( 
.A(n_324),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_L g385 ( 
.A(n_329),
.B(n_292),
.Y(n_385)
);

INVx2_ASAP7_75t_L g386 ( 
.A(n_286),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_297),
.B(n_224),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_298),
.B(n_306),
.Y(n_388)
);

CKINVDCx20_ASAP7_75t_R g389 ( 
.A(n_304),
.Y(n_389)
);

INVx2_ASAP7_75t_SL g390 ( 
.A(n_326),
.Y(n_390)
);

INVx3_ASAP7_75t_L g391 ( 
.A(n_287),
.Y(n_391)
);

INVx4_ASAP7_75t_L g392 ( 
.A(n_324),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_327),
.B(n_228),
.Y(n_393)
);

OR2x6_ASAP7_75t_L g394 ( 
.A(n_307),
.B(n_276),
.Y(n_394)
);

AND2x2_ASAP7_75t_L g395 ( 
.A(n_327),
.B(n_211),
.Y(n_395)
);

AND2x4_ASAP7_75t_L g396 ( 
.A(n_318),
.B(n_29),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_SL g397 ( 
.A(n_326),
.B(n_211),
.Y(n_397)
);

AND2x4_ASAP7_75t_L g398 ( 
.A(n_383),
.B(n_299),
.Y(n_398)
);

AOI22xp33_ASAP7_75t_L g399 ( 
.A1(n_354),
.A2(n_329),
.B1(n_211),
.B2(n_320),
.Y(n_399)
);

NOR2xp33_ASAP7_75t_L g400 ( 
.A(n_332),
.B(n_315),
.Y(n_400)
);

OR2x6_ASAP7_75t_L g401 ( 
.A(n_394),
.B(n_307),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_L g402 ( 
.A(n_332),
.B(n_321),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_365),
.Y(n_403)
);

OR2x6_ASAP7_75t_L g404 ( 
.A(n_394),
.B(n_320),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_388),
.B(n_285),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_L g406 ( 
.A(n_385),
.B(n_290),
.Y(n_406)
);

NOR2xp33_ASAP7_75t_L g407 ( 
.A(n_385),
.B(n_312),
.Y(n_407)
);

AOI22xp33_ASAP7_75t_L g408 ( 
.A1(n_354),
.A2(n_211),
.B1(n_299),
.B2(n_282),
.Y(n_408)
);

NOR3xp33_ASAP7_75t_L g409 ( 
.A(n_356),
.B(n_284),
.C(n_282),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_365),
.B(n_293),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_352),
.B(n_293),
.Y(n_411)
);

BUFx6f_ASAP7_75t_L g412 ( 
.A(n_344),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_L g413 ( 
.A(n_390),
.B(n_309),
.Y(n_413)
);

AOI21xp5_ASAP7_75t_L g414 ( 
.A1(n_359),
.A2(n_284),
.B(n_293),
.Y(n_414)
);

BUFx3_ASAP7_75t_L g415 ( 
.A(n_374),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_SL g416 ( 
.A(n_384),
.B(n_211),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_383),
.Y(n_417)
);

INVxp67_ASAP7_75t_L g418 ( 
.A(n_333),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_331),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_334),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_367),
.B(n_287),
.Y(n_421)
);

AND2x2_ASAP7_75t_L g422 ( 
.A(n_351),
.B(n_291),
.Y(n_422)
);

INVxp67_ASAP7_75t_L g423 ( 
.A(n_348),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_367),
.B(n_287),
.Y(n_424)
);

INVx2_ASAP7_75t_SL g425 ( 
.A(n_347),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_348),
.B(n_291),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_357),
.Y(n_427)
);

INVx2_ASAP7_75t_L g428 ( 
.A(n_336),
.Y(n_428)
);

AND2x6_ASAP7_75t_SL g429 ( 
.A(n_394),
.B(n_328),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_387),
.B(n_32),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_SL g431 ( 
.A(n_384),
.B(n_2),
.Y(n_431)
);

AOI22xp5_ASAP7_75t_L g432 ( 
.A1(n_339),
.A2(n_84),
.B1(n_170),
.B2(n_169),
.Y(n_432)
);

NOR2xp33_ASAP7_75t_L g433 ( 
.A(n_393),
.B(n_2),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_344),
.B(n_33),
.Y(n_434)
);

OR2x2_ASAP7_75t_L g435 ( 
.A(n_378),
.B(n_3),
.Y(n_435)
);

NOR2xp33_ASAP7_75t_L g436 ( 
.A(n_377),
.B(n_4),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_375),
.B(n_34),
.Y(n_437)
);

NAND2xp33_ASAP7_75t_L g438 ( 
.A(n_361),
.B(n_37),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_337),
.Y(n_439)
);

AOI22xp5_ASAP7_75t_L g440 ( 
.A1(n_339),
.A2(n_86),
.B1(n_166),
.B2(n_165),
.Y(n_440)
);

NAND2xp33_ASAP7_75t_L g441 ( 
.A(n_361),
.B(n_38),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_340),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_341),
.Y(n_443)
);

BUFx12f_ASAP7_75t_L g444 ( 
.A(n_357),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_SL g445 ( 
.A(n_392),
.B(n_4),
.Y(n_445)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_336),
.Y(n_446)
);

NOR2xp33_ASAP7_75t_L g447 ( 
.A(n_379),
.B(n_5),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_SL g448 ( 
.A(n_392),
.B(n_5),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_375),
.B(n_42),
.Y(n_449)
);

BUFx6f_ASAP7_75t_L g450 ( 
.A(n_382),
.Y(n_450)
);

AOI22xp33_ASAP7_75t_L g451 ( 
.A1(n_396),
.A2(n_6),
.B1(n_7),
.B2(n_9),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_346),
.B(n_353),
.Y(n_452)
);

NOR2xp33_ASAP7_75t_L g453 ( 
.A(n_335),
.B(n_6),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_358),
.B(n_44),
.Y(n_454)
);

OR2x2_ASAP7_75t_L g455 ( 
.A(n_381),
.B(n_7),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_SL g456 ( 
.A(n_371),
.B(n_10),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_364),
.B(n_370),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_338),
.B(n_45),
.Y(n_458)
);

AND2x2_ASAP7_75t_L g459 ( 
.A(n_343),
.B(n_10),
.Y(n_459)
);

INVxp67_ASAP7_75t_SL g460 ( 
.A(n_338),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_338),
.B(n_46),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_SL g462 ( 
.A(n_371),
.B(n_12),
.Y(n_462)
);

NOR2xp33_ASAP7_75t_L g463 ( 
.A(n_382),
.B(n_12),
.Y(n_463)
);

AOI22xp33_ASAP7_75t_L g464 ( 
.A1(n_396),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_464)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_369),
.Y(n_465)
);

INVx2_ASAP7_75t_SL g466 ( 
.A(n_339),
.Y(n_466)
);

AOI22xp33_ASAP7_75t_L g467 ( 
.A1(n_396),
.A2(n_397),
.B1(n_395),
.B2(n_368),
.Y(n_467)
);

INVx4_ASAP7_75t_L g468 ( 
.A(n_412),
.Y(n_468)
);

AND2x2_ASAP7_75t_L g469 ( 
.A(n_423),
.B(n_422),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_423),
.B(n_397),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_403),
.Y(n_471)
);

AND3x1_ASAP7_75t_L g472 ( 
.A(n_453),
.B(n_459),
.C(n_407),
.Y(n_472)
);

INVx3_ASAP7_75t_L g473 ( 
.A(n_412),
.Y(n_473)
);

INVx4_ASAP7_75t_L g474 ( 
.A(n_412),
.Y(n_474)
);

AOI221xp5_ASAP7_75t_SL g475 ( 
.A1(n_451),
.A2(n_363),
.B1(n_376),
.B2(n_338),
.C(n_362),
.Y(n_475)
);

AND2x2_ASAP7_75t_L g476 ( 
.A(n_418),
.B(n_391),
.Y(n_476)
);

INVx2_ASAP7_75t_L g477 ( 
.A(n_465),
.Y(n_477)
);

CKINVDCx8_ASAP7_75t_R g478 ( 
.A(n_429),
.Y(n_478)
);

AND2x2_ASAP7_75t_L g479 ( 
.A(n_418),
.B(n_391),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_SL g480 ( 
.A(n_405),
.B(n_350),
.Y(n_480)
);

INVx2_ASAP7_75t_SL g481 ( 
.A(n_398),
.Y(n_481)
);

AND2x2_ASAP7_75t_L g482 ( 
.A(n_466),
.B(n_369),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_406),
.B(n_350),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_419),
.Y(n_484)
);

INVxp67_ASAP7_75t_SL g485 ( 
.A(n_460),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_420),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_426),
.B(n_350),
.Y(n_487)
);

AOI22xp33_ASAP7_75t_L g488 ( 
.A1(n_436),
.A2(n_368),
.B1(n_372),
.B2(n_360),
.Y(n_488)
);

NOR2xp33_ASAP7_75t_L g489 ( 
.A(n_400),
.B(n_374),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_428),
.Y(n_490)
);

NOR3xp33_ASAP7_75t_SL g491 ( 
.A(n_413),
.B(n_389),
.C(n_14),
.Y(n_491)
);

BUFx4f_ASAP7_75t_L g492 ( 
.A(n_450),
.Y(n_492)
);

CKINVDCx5p33_ASAP7_75t_R g493 ( 
.A(n_427),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_SL g494 ( 
.A(n_398),
.B(n_350),
.Y(n_494)
);

INVx3_ASAP7_75t_L g495 ( 
.A(n_412),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_446),
.Y(n_496)
);

NOR2xp33_ASAP7_75t_L g497 ( 
.A(n_402),
.B(n_389),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_SL g498 ( 
.A(n_450),
.B(n_362),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_SL g499 ( 
.A(n_450),
.B(n_362),
.Y(n_499)
);

INVx2_ASAP7_75t_L g500 ( 
.A(n_439),
.Y(n_500)
);

INVx5_ASAP7_75t_L g501 ( 
.A(n_450),
.Y(n_501)
);

NOR2xp33_ASAP7_75t_L g502 ( 
.A(n_425),
.B(n_362),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_467),
.B(n_373),
.Y(n_503)
);

CKINVDCx8_ASAP7_75t_R g504 ( 
.A(n_401),
.Y(n_504)
);

HB1xp67_ASAP7_75t_L g505 ( 
.A(n_435),
.Y(n_505)
);

INVx2_ASAP7_75t_L g506 ( 
.A(n_442),
.Y(n_506)
);

NAND3xp33_ASAP7_75t_SL g507 ( 
.A(n_451),
.B(n_386),
.C(n_380),
.Y(n_507)
);

HB1xp67_ASAP7_75t_L g508 ( 
.A(n_455),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_SL g509 ( 
.A(n_417),
.B(n_373),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_443),
.Y(n_510)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_452),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_467),
.B(n_380),
.Y(n_512)
);

BUFx3_ASAP7_75t_L g513 ( 
.A(n_415),
.Y(n_513)
);

OR2x2_ASAP7_75t_L g514 ( 
.A(n_401),
.B(n_386),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_460),
.B(n_360),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_457),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_421),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_424),
.Y(n_518)
);

AOI22xp5_ASAP7_75t_L g519 ( 
.A1(n_447),
.A2(n_372),
.B1(n_368),
.B2(n_360),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_399),
.B(n_409),
.Y(n_520)
);

INVx2_ASAP7_75t_L g521 ( 
.A(n_458),
.Y(n_521)
);

NAND3xp33_ASAP7_75t_L g522 ( 
.A(n_433),
.B(n_366),
.C(n_355),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_L g523 ( 
.A(n_516),
.B(n_409),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_516),
.B(n_464),
.Y(n_524)
);

BUFx6f_ASAP7_75t_L g525 ( 
.A(n_492),
.Y(n_525)
);

AOI221x1_ASAP7_75t_L g526 ( 
.A1(n_483),
.A2(n_463),
.B1(n_430),
.B2(n_414),
.C(n_454),
.Y(n_526)
);

OAI21x1_ASAP7_75t_L g527 ( 
.A1(n_515),
.A2(n_434),
.B(n_437),
.Y(n_527)
);

AO31x2_ASAP7_75t_L g528 ( 
.A1(n_521),
.A2(n_461),
.A3(n_449),
.B(n_411),
.Y(n_528)
);

OAI21x1_ASAP7_75t_L g529 ( 
.A1(n_521),
.A2(n_416),
.B(n_410),
.Y(n_529)
);

INVx5_ASAP7_75t_L g530 ( 
.A(n_501),
.Y(n_530)
);

OAI21x1_ASAP7_75t_L g531 ( 
.A1(n_503),
.A2(n_408),
.B(n_345),
.Y(n_531)
);

OAI21xp5_ASAP7_75t_L g532 ( 
.A1(n_512),
.A2(n_441),
.B(n_438),
.Y(n_532)
);

AO31x2_ASAP7_75t_L g533 ( 
.A1(n_517),
.A2(n_518),
.A3(n_487),
.B(n_520),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_L g534 ( 
.A(n_511),
.B(n_464),
.Y(n_534)
);

A2O1A1Ixp33_ASAP7_75t_L g535 ( 
.A1(n_511),
.A2(n_462),
.B(n_456),
.C(n_440),
.Y(n_535)
);

INVx5_ASAP7_75t_L g536 ( 
.A(n_501),
.Y(n_536)
);

AO31x2_ASAP7_75t_L g537 ( 
.A1(n_517),
.A2(n_342),
.A3(n_345),
.B(n_355),
.Y(n_537)
);

OAI21xp5_ASAP7_75t_L g538 ( 
.A1(n_470),
.A2(n_448),
.B(n_445),
.Y(n_538)
);

AND2x2_ASAP7_75t_L g539 ( 
.A(n_469),
.B(n_404),
.Y(n_539)
);

AOI21xp5_ASAP7_75t_SL g540 ( 
.A1(n_485),
.A2(n_432),
.B(n_431),
.Y(n_540)
);

INVx3_ASAP7_75t_L g541 ( 
.A(n_468),
.Y(n_541)
);

AOI21xp33_ASAP7_75t_L g542 ( 
.A1(n_489),
.A2(n_497),
.B(n_469),
.Y(n_542)
);

AOI21xp5_ASAP7_75t_L g543 ( 
.A1(n_492),
.A2(n_349),
.B(n_342),
.Y(n_543)
);

INVx2_ASAP7_75t_L g544 ( 
.A(n_477),
.Y(n_544)
);

NOR2xp33_ASAP7_75t_L g545 ( 
.A(n_505),
.B(n_444),
.Y(n_545)
);

OAI21xp5_ASAP7_75t_L g546 ( 
.A1(n_475),
.A2(n_366),
.B(n_372),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_L g547 ( 
.A(n_476),
.B(n_360),
.Y(n_547)
);

OAI21x1_ASAP7_75t_L g548 ( 
.A1(n_498),
.A2(n_372),
.B(n_368),
.Y(n_548)
);

AO31x2_ASAP7_75t_L g549 ( 
.A1(n_518),
.A2(n_502),
.A3(n_500),
.B(n_506),
.Y(n_549)
);

AOI221x1_ASAP7_75t_L g550 ( 
.A1(n_522),
.A2(n_372),
.B1(n_368),
.B2(n_360),
.C(n_404),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_510),
.Y(n_551)
);

INVx5_ASAP7_75t_L g552 ( 
.A(n_501),
.Y(n_552)
);

NAND3xp33_ASAP7_75t_SL g553 ( 
.A(n_493),
.B(n_401),
.C(n_404),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_476),
.B(n_349),
.Y(n_554)
);

INVx1_ASAP7_75t_SL g555 ( 
.A(n_479),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_L g556 ( 
.A(n_479),
.B(n_349),
.Y(n_556)
);

OAI21x1_ASAP7_75t_L g557 ( 
.A1(n_499),
.A2(n_96),
.B(n_163),
.Y(n_557)
);

AOI21xp5_ASAP7_75t_SL g558 ( 
.A1(n_468),
.A2(n_95),
.B(n_162),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_L g559 ( 
.A(n_510),
.B(n_13),
.Y(n_559)
);

AOI21xp5_ASAP7_75t_L g560 ( 
.A1(n_492),
.A2(n_501),
.B(n_480),
.Y(n_560)
);

AOI21xp5_ASAP7_75t_L g561 ( 
.A1(n_501),
.A2(n_97),
.B(n_161),
.Y(n_561)
);

OAI21xp5_ASAP7_75t_L g562 ( 
.A1(n_507),
.A2(n_93),
.B(n_158),
.Y(n_562)
);

AOI21xp5_ASAP7_75t_L g563 ( 
.A1(n_494),
.A2(n_488),
.B(n_519),
.Y(n_563)
);

OAI21x1_ASAP7_75t_L g564 ( 
.A1(n_473),
.A2(n_92),
.B(n_157),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_L g565 ( 
.A(n_500),
.B(n_15),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_506),
.Y(n_566)
);

OAI21xp5_ASAP7_75t_L g567 ( 
.A1(n_477),
.A2(n_486),
.B(n_484),
.Y(n_567)
);

BUFx3_ASAP7_75t_L g568 ( 
.A(n_525),
.Y(n_568)
);

AND2x2_ASAP7_75t_L g569 ( 
.A(n_555),
.B(n_472),
.Y(n_569)
);

A2O1A1Ixp33_ASAP7_75t_L g570 ( 
.A1(n_535),
.A2(n_481),
.B(n_491),
.C(n_514),
.Y(n_570)
);

AND2x2_ASAP7_75t_L g571 ( 
.A(n_555),
.B(n_482),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_551),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_566),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_544),
.Y(n_574)
);

OAI22xp33_ASAP7_75t_L g575 ( 
.A1(n_542),
.A2(n_508),
.B1(n_493),
.B2(n_504),
.Y(n_575)
);

OAI21x1_ASAP7_75t_L g576 ( 
.A1(n_531),
.A2(n_509),
.B(n_473),
.Y(n_576)
);

OR2x6_ASAP7_75t_L g577 ( 
.A(n_540),
.B(n_514),
.Y(n_577)
);

O2A1O1Ixp33_ASAP7_75t_L g578 ( 
.A1(n_523),
.A2(n_481),
.B(n_471),
.C(n_496),
.Y(n_578)
);

BUFx2_ASAP7_75t_L g579 ( 
.A(n_539),
.Y(n_579)
);

AND2x4_ASAP7_75t_L g580 ( 
.A(n_525),
.B(n_482),
.Y(n_580)
);

OA21x2_ASAP7_75t_L g581 ( 
.A1(n_526),
.A2(n_562),
.B(n_532),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_549),
.Y(n_582)
);

OAI21x1_ASAP7_75t_L g583 ( 
.A1(n_546),
.A2(n_495),
.B(n_473),
.Y(n_583)
);

OAI21xp5_ASAP7_75t_L g584 ( 
.A1(n_563),
.A2(n_490),
.B(n_496),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_565),
.Y(n_585)
);

AND2x4_ASAP7_75t_L g586 ( 
.A(n_525),
.B(n_468),
.Y(n_586)
);

OAI22xp33_ASAP7_75t_L g587 ( 
.A1(n_524),
.A2(n_504),
.B1(n_513),
.B2(n_478),
.Y(n_587)
);

INVx2_ASAP7_75t_L g588 ( 
.A(n_537),
.Y(n_588)
);

INVx2_ASAP7_75t_L g589 ( 
.A(n_537),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_L g590 ( 
.A(n_534),
.B(n_490),
.Y(n_590)
);

OAI21x1_ASAP7_75t_L g591 ( 
.A1(n_546),
.A2(n_495),
.B(n_474),
.Y(n_591)
);

BUFx12f_ASAP7_75t_L g592 ( 
.A(n_530),
.Y(n_592)
);

INVx2_ASAP7_75t_L g593 ( 
.A(n_537),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_559),
.Y(n_594)
);

OAI21x1_ASAP7_75t_L g595 ( 
.A1(n_527),
.A2(n_495),
.B(n_474),
.Y(n_595)
);

AOI21xp5_ASAP7_75t_L g596 ( 
.A1(n_530),
.A2(n_474),
.B(n_513),
.Y(n_596)
);

OAI21x1_ASAP7_75t_L g597 ( 
.A1(n_564),
.A2(n_98),
.B(n_171),
.Y(n_597)
);

AO31x2_ASAP7_75t_L g598 ( 
.A1(n_550),
.A2(n_16),
.A3(n_17),
.B(n_18),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_567),
.Y(n_599)
);

HB1xp67_ASAP7_75t_L g600 ( 
.A(n_567),
.Y(n_600)
);

AOI221xp5_ASAP7_75t_L g601 ( 
.A1(n_553),
.A2(n_478),
.B1(n_19),
.B2(n_21),
.C(n_22),
.Y(n_601)
);

INVx3_ASAP7_75t_L g602 ( 
.A(n_530),
.Y(n_602)
);

CKINVDCx5p33_ASAP7_75t_R g603 ( 
.A(n_545),
.Y(n_603)
);

AOI22xp33_ASAP7_75t_L g604 ( 
.A1(n_562),
.A2(n_16),
.B1(n_19),
.B2(n_21),
.Y(n_604)
);

O2A1O1Ixp33_ASAP7_75t_SL g605 ( 
.A1(n_547),
.A2(n_104),
.B(n_153),
.C(n_151),
.Y(n_605)
);

INVx2_ASAP7_75t_SL g606 ( 
.A(n_536),
.Y(n_606)
);

NOR2xp33_ASAP7_75t_L g607 ( 
.A(n_538),
.B(n_22),
.Y(n_607)
);

OAI21x1_ASAP7_75t_L g608 ( 
.A1(n_529),
.A2(n_100),
.B(n_149),
.Y(n_608)
);

OAI21x1_ASAP7_75t_L g609 ( 
.A1(n_557),
.A2(n_91),
.B(n_148),
.Y(n_609)
);

INVx6_ASAP7_75t_L g610 ( 
.A(n_536),
.Y(n_610)
);

INVx2_ASAP7_75t_L g611 ( 
.A(n_572),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_572),
.Y(n_612)
);

INVx2_ASAP7_75t_L g613 ( 
.A(n_588),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_573),
.Y(n_614)
);

AOI221xp5_ASAP7_75t_L g615 ( 
.A1(n_607),
.A2(n_558),
.B1(n_561),
.B2(n_554),
.C(n_556),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_574),
.Y(n_616)
);

INVx2_ASAP7_75t_L g617 ( 
.A(n_588),
.Y(n_617)
);

AND2x4_ASAP7_75t_L g618 ( 
.A(n_580),
.B(n_541),
.Y(n_618)
);

BUFx8_ASAP7_75t_L g619 ( 
.A(n_592),
.Y(n_619)
);

AND2x4_ASAP7_75t_L g620 ( 
.A(n_580),
.B(n_541),
.Y(n_620)
);

OAI22xp5_ASAP7_75t_L g621 ( 
.A1(n_575),
.A2(n_552),
.B1(n_536),
.B2(n_560),
.Y(n_621)
);

OR2x2_ASAP7_75t_L g622 ( 
.A(n_579),
.B(n_533),
.Y(n_622)
);

INVx2_ASAP7_75t_L g623 ( 
.A(n_589),
.Y(n_623)
);

BUFx2_ASAP7_75t_L g624 ( 
.A(n_579),
.Y(n_624)
);

A2O1A1Ixp33_ASAP7_75t_L g625 ( 
.A1(n_604),
.A2(n_543),
.B(n_552),
.C(n_548),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_L g626 ( 
.A(n_594),
.B(n_533),
.Y(n_626)
);

A2O1A1Ixp33_ASAP7_75t_L g627 ( 
.A1(n_601),
.A2(n_552),
.B(n_533),
.C(n_549),
.Y(n_627)
);

BUFx3_ASAP7_75t_L g628 ( 
.A(n_568),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_571),
.B(n_549),
.Y(n_629)
);

AOI22xp33_ASAP7_75t_L g630 ( 
.A1(n_585),
.A2(n_569),
.B1(n_581),
.B2(n_600),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_L g631 ( 
.A(n_571),
.B(n_528),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_582),
.Y(n_632)
);

AND2x2_ASAP7_75t_L g633 ( 
.A(n_569),
.B(n_528),
.Y(n_633)
);

INVx2_ASAP7_75t_L g634 ( 
.A(n_589),
.Y(n_634)
);

NAND2xp33_ASAP7_75t_R g635 ( 
.A(n_581),
.B(n_528),
.Y(n_635)
);

AND2x4_ASAP7_75t_L g636 ( 
.A(n_580),
.B(n_47),
.Y(n_636)
);

AND2x4_ASAP7_75t_L g637 ( 
.A(n_586),
.B(n_48),
.Y(n_637)
);

AND2x2_ASAP7_75t_L g638 ( 
.A(n_568),
.B(n_570),
.Y(n_638)
);

OAI21xp33_ASAP7_75t_L g639 ( 
.A1(n_590),
.A2(n_23),
.B(n_24),
.Y(n_639)
);

AND2x2_ASAP7_75t_L g640 ( 
.A(n_603),
.B(n_23),
.Y(n_640)
);

AOI22xp33_ASAP7_75t_L g641 ( 
.A1(n_581),
.A2(n_26),
.B1(n_27),
.B2(n_49),
.Y(n_641)
);

NAND2x1_ASAP7_75t_L g642 ( 
.A(n_610),
.B(n_602),
.Y(n_642)
);

AND2x4_ASAP7_75t_L g643 ( 
.A(n_586),
.B(n_109),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_582),
.Y(n_644)
);

AOI21xp33_ASAP7_75t_L g645 ( 
.A1(n_578),
.A2(n_577),
.B(n_587),
.Y(n_645)
);

OAI21x1_ASAP7_75t_L g646 ( 
.A1(n_595),
.A2(n_608),
.B(n_576),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_L g647 ( 
.A(n_599),
.B(n_27),
.Y(n_647)
);

INVx4_ASAP7_75t_L g648 ( 
.A(n_592),
.Y(n_648)
);

AND2x2_ASAP7_75t_L g649 ( 
.A(n_603),
.B(n_50),
.Y(n_649)
);

AND2x4_ASAP7_75t_L g650 ( 
.A(n_586),
.B(n_51),
.Y(n_650)
);

CKINVDCx5p33_ASAP7_75t_R g651 ( 
.A(n_577),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_584),
.Y(n_652)
);

CKINVDCx5p33_ASAP7_75t_R g653 ( 
.A(n_577),
.Y(n_653)
);

INVx4_ASAP7_75t_L g654 ( 
.A(n_610),
.Y(n_654)
);

AND2x2_ASAP7_75t_L g655 ( 
.A(n_577),
.B(n_598),
.Y(n_655)
);

INVx2_ASAP7_75t_L g656 ( 
.A(n_593),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_L g657 ( 
.A(n_596),
.B(n_52),
.Y(n_657)
);

AOI22xp33_ASAP7_75t_L g658 ( 
.A1(n_593),
.A2(n_155),
.B1(n_56),
.B2(n_57),
.Y(n_658)
);

AOI22xp33_ASAP7_75t_L g659 ( 
.A1(n_610),
.A2(n_54),
.B1(n_58),
.B2(n_59),
.Y(n_659)
);

OAI221xp5_ASAP7_75t_L g660 ( 
.A1(n_605),
.A2(n_61),
.B1(n_62),
.B2(n_63),
.C(n_64),
.Y(n_660)
);

AOI221x1_ASAP7_75t_L g661 ( 
.A1(n_602),
.A2(n_65),
.B1(n_68),
.B2(n_69),
.C(n_70),
.Y(n_661)
);

OAI221xp5_ASAP7_75t_L g662 ( 
.A1(n_606),
.A2(n_71),
.B1(n_72),
.B2(n_73),
.C(n_75),
.Y(n_662)
);

AND2x2_ASAP7_75t_L g663 ( 
.A(n_598),
.B(n_79),
.Y(n_663)
);

CKINVDCx5p33_ASAP7_75t_R g664 ( 
.A(n_619),
.Y(n_664)
);

AOI222xp33_ASAP7_75t_L g665 ( 
.A1(n_639),
.A2(n_606),
.B1(n_610),
.B2(n_602),
.C1(n_583),
.C2(n_597),
.Y(n_665)
);

AOI22xp33_ASAP7_75t_L g666 ( 
.A1(n_641),
.A2(n_597),
.B1(n_609),
.B2(n_576),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_L g667 ( 
.A(n_624),
.B(n_647),
.Y(n_667)
);

AOI222xp33_ASAP7_75t_L g668 ( 
.A1(n_641),
.A2(n_583),
.B1(n_591),
.B2(n_609),
.C1(n_608),
.C2(n_598),
.Y(n_668)
);

HB1xp67_ASAP7_75t_L g669 ( 
.A(n_613),
.Y(n_669)
);

AOI22xp33_ASAP7_75t_L g670 ( 
.A1(n_645),
.A2(n_591),
.B1(n_595),
.B2(n_598),
.Y(n_670)
);

AO21x2_ASAP7_75t_L g671 ( 
.A1(n_646),
.A2(n_625),
.B(n_627),
.Y(n_671)
);

NAND4xp25_ASAP7_75t_L g672 ( 
.A(n_640),
.B(n_598),
.C(n_81),
.D(n_82),
.Y(n_672)
);

OAI21x1_ASAP7_75t_L g673 ( 
.A1(n_613),
.A2(n_80),
.B(n_83),
.Y(n_673)
);

AOI22xp33_ASAP7_75t_L g674 ( 
.A1(n_638),
.A2(n_85),
.B1(n_90),
.B2(n_106),
.Y(n_674)
);

BUFx4f_ASAP7_75t_SL g675 ( 
.A(n_619),
.Y(n_675)
);

INVx2_ASAP7_75t_L g676 ( 
.A(n_611),
.Y(n_676)
);

NAND3xp33_ASAP7_75t_L g677 ( 
.A(n_658),
.B(n_107),
.C(n_110),
.Y(n_677)
);

INVx2_ASAP7_75t_L g678 ( 
.A(n_611),
.Y(n_678)
);

AOI221xp5_ASAP7_75t_L g679 ( 
.A1(n_660),
.A2(n_111),
.B1(n_112),
.B2(n_114),
.C(n_115),
.Y(n_679)
);

OAI22xp5_ASAP7_75t_L g680 ( 
.A1(n_651),
.A2(n_117),
.B1(n_120),
.B2(n_121),
.Y(n_680)
);

INVx1_ASAP7_75t_SL g681 ( 
.A(n_628),
.Y(n_681)
);

AOI21xp5_ASAP7_75t_L g682 ( 
.A1(n_625),
.A2(n_122),
.B(n_123),
.Y(n_682)
);

AO21x2_ASAP7_75t_L g683 ( 
.A1(n_627),
.A2(n_125),
.B(n_127),
.Y(n_683)
);

AOI22xp33_ASAP7_75t_L g684 ( 
.A1(n_658),
.A2(n_128),
.B1(n_129),
.B2(n_130),
.Y(n_684)
);

AOI21xp5_ASAP7_75t_L g685 ( 
.A1(n_652),
.A2(n_131),
.B(n_132),
.Y(n_685)
);

AOI221xp5_ASAP7_75t_L g686 ( 
.A1(n_630),
.A2(n_133),
.B1(n_136),
.B2(n_137),
.C(n_138),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_612),
.Y(n_687)
);

OAI22xp5_ASAP7_75t_L g688 ( 
.A1(n_653),
.A2(n_139),
.B1(n_140),
.B2(n_141),
.Y(n_688)
);

INVx2_ASAP7_75t_L g689 ( 
.A(n_616),
.Y(n_689)
);

AOI22xp33_ASAP7_75t_L g690 ( 
.A1(n_663),
.A2(n_142),
.B1(n_143),
.B2(n_144),
.Y(n_690)
);

OAI221xp5_ASAP7_75t_L g691 ( 
.A1(n_659),
.A2(n_146),
.B1(n_615),
.B2(n_662),
.C(n_630),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_632),
.Y(n_692)
);

AOI22xp5_ASAP7_75t_L g693 ( 
.A1(n_636),
.A2(n_637),
.B1(n_643),
.B2(n_650),
.Y(n_693)
);

INVx2_ASAP7_75t_L g694 ( 
.A(n_614),
.Y(n_694)
);

OAI22xp5_ASAP7_75t_L g695 ( 
.A1(n_659),
.A2(n_622),
.B1(n_636),
.B2(n_629),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_L g696 ( 
.A(n_633),
.B(n_626),
.Y(n_696)
);

AOI21xp5_ASAP7_75t_SL g697 ( 
.A1(n_637),
.A2(n_643),
.B(n_650),
.Y(n_697)
);

OAI22xp33_ASAP7_75t_L g698 ( 
.A1(n_661),
.A2(n_631),
.B1(n_648),
.B2(n_654),
.Y(n_698)
);

AOI222xp33_ASAP7_75t_L g699 ( 
.A1(n_649),
.A2(n_636),
.B1(n_619),
.B2(n_637),
.C1(n_650),
.C2(n_643),
.Y(n_699)
);

AOI22xp33_ASAP7_75t_L g700 ( 
.A1(n_648),
.A2(n_618),
.B1(n_620),
.B2(n_655),
.Y(n_700)
);

INVx2_ASAP7_75t_SL g701 ( 
.A(n_628),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_644),
.Y(n_702)
);

AOI221xp5_ASAP7_75t_L g703 ( 
.A1(n_621),
.A2(n_648),
.B1(n_657),
.B2(n_620),
.C(n_618),
.Y(n_703)
);

AND2x4_ASAP7_75t_L g704 ( 
.A(n_654),
.B(n_618),
.Y(n_704)
);

HB1xp67_ASAP7_75t_L g705 ( 
.A(n_669),
.Y(n_705)
);

INVx2_ASAP7_75t_L g706 ( 
.A(n_692),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_702),
.Y(n_707)
);

INVx2_ASAP7_75t_L g708 ( 
.A(n_687),
.Y(n_708)
);

INVx2_ASAP7_75t_L g709 ( 
.A(n_676),
.Y(n_709)
);

INVx2_ASAP7_75t_L g710 ( 
.A(n_678),
.Y(n_710)
);

BUFx3_ASAP7_75t_L g711 ( 
.A(n_704),
.Y(n_711)
);

NOR2x1p5_ASAP7_75t_L g712 ( 
.A(n_672),
.B(n_642),
.Y(n_712)
);

AND2x2_ASAP7_75t_L g713 ( 
.A(n_696),
.B(n_617),
.Y(n_713)
);

OR2x2_ASAP7_75t_L g714 ( 
.A(n_667),
.B(n_617),
.Y(n_714)
);

AOI322xp5_ASAP7_75t_L g715 ( 
.A1(n_690),
.A2(n_620),
.A3(n_623),
.B1(n_634),
.B2(n_656),
.C1(n_635),
.C2(n_654),
.Y(n_715)
);

AND2x2_ASAP7_75t_L g716 ( 
.A(n_694),
.B(n_634),
.Y(n_716)
);

AND2x2_ASAP7_75t_L g717 ( 
.A(n_700),
.B(n_656),
.Y(n_717)
);

OAI22xp33_ASAP7_75t_L g718 ( 
.A1(n_691),
.A2(n_635),
.B1(n_677),
.B2(n_693),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_689),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_671),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_671),
.Y(n_721)
);

INVxp67_ASAP7_75t_L g722 ( 
.A(n_683),
.Y(n_722)
);

AND2x4_ASAP7_75t_L g723 ( 
.A(n_683),
.B(n_700),
.Y(n_723)
);

AND2x2_ASAP7_75t_L g724 ( 
.A(n_670),
.B(n_695),
.Y(n_724)
);

INVx3_ASAP7_75t_L g725 ( 
.A(n_673),
.Y(n_725)
);

INVx2_ASAP7_75t_L g726 ( 
.A(n_704),
.Y(n_726)
);

INVx2_ASAP7_75t_L g727 ( 
.A(n_701),
.Y(n_727)
);

AND2x2_ASAP7_75t_L g728 ( 
.A(n_670),
.B(n_668),
.Y(n_728)
);

AND2x2_ASAP7_75t_L g729 ( 
.A(n_690),
.B(n_681),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_698),
.Y(n_730)
);

AND2x2_ASAP7_75t_L g731 ( 
.A(n_665),
.B(n_666),
.Y(n_731)
);

AOI22xp33_ASAP7_75t_L g732 ( 
.A1(n_684),
.A2(n_679),
.B1(n_703),
.B2(n_686),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_L g733 ( 
.A(n_698),
.B(n_682),
.Y(n_733)
);

BUFx6f_ASAP7_75t_L g734 ( 
.A(n_697),
.Y(n_734)
);

OR2x2_ASAP7_75t_L g735 ( 
.A(n_705),
.B(n_666),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_706),
.Y(n_736)
);

CKINVDCx5p33_ASAP7_75t_R g737 ( 
.A(n_727),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_SL g738 ( 
.A(n_734),
.B(n_699),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_714),
.B(n_684),
.Y(n_739)
);

OAI22xp5_ASAP7_75t_L g740 ( 
.A1(n_732),
.A2(n_674),
.B1(n_675),
.B2(n_685),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_706),
.Y(n_741)
);

BUFx12f_ASAP7_75t_L g742 ( 
.A(n_712),
.Y(n_742)
);

NAND3xp33_ASAP7_75t_L g743 ( 
.A(n_733),
.B(n_680),
.C(n_688),
.Y(n_743)
);

OAI21xp5_ASAP7_75t_L g744 ( 
.A1(n_733),
.A2(n_664),
.B(n_675),
.Y(n_744)
);

INVx2_ASAP7_75t_L g745 ( 
.A(n_706),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_L g746 ( 
.A(n_714),
.B(n_713),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_708),
.Y(n_747)
);

OR2x2_ASAP7_75t_L g748 ( 
.A(n_705),
.B(n_708),
.Y(n_748)
);

AND2x2_ASAP7_75t_L g749 ( 
.A(n_724),
.B(n_723),
.Y(n_749)
);

INVx2_ASAP7_75t_L g750 ( 
.A(n_708),
.Y(n_750)
);

AO21x2_ASAP7_75t_L g751 ( 
.A1(n_720),
.A2(n_721),
.B(n_722),
.Y(n_751)
);

BUFx3_ASAP7_75t_L g752 ( 
.A(n_734),
.Y(n_752)
);

AO21x2_ASAP7_75t_L g753 ( 
.A1(n_720),
.A2(n_721),
.B(n_722),
.Y(n_753)
);

INVx2_ASAP7_75t_SL g754 ( 
.A(n_748),
.Y(n_754)
);

AND2x2_ASAP7_75t_L g755 ( 
.A(n_749),
.B(n_723),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_745),
.Y(n_756)
);

AND2x2_ASAP7_75t_L g757 ( 
.A(n_749),
.B(n_723),
.Y(n_757)
);

AND2x2_ASAP7_75t_L g758 ( 
.A(n_746),
.B(n_723),
.Y(n_758)
);

OR2x2_ASAP7_75t_L g759 ( 
.A(n_748),
.B(n_730),
.Y(n_759)
);

INVx2_ASAP7_75t_L g760 ( 
.A(n_745),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_737),
.B(n_730),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_736),
.Y(n_762)
);

INVx5_ASAP7_75t_L g763 ( 
.A(n_742),
.Y(n_763)
);

AND2x4_ASAP7_75t_L g764 ( 
.A(n_752),
.B(n_726),
.Y(n_764)
);

AOI221x1_ASAP7_75t_L g765 ( 
.A1(n_743),
.A2(n_728),
.B1(n_727),
.B2(n_731),
.C(n_724),
.Y(n_765)
);

AND2x2_ASAP7_75t_L g766 ( 
.A(n_745),
.B(n_728),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_L g767 ( 
.A(n_739),
.B(n_713),
.Y(n_767)
);

AND2x2_ASAP7_75t_L g768 ( 
.A(n_755),
.B(n_726),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_L g769 ( 
.A(n_766),
.B(n_747),
.Y(n_769)
);

AND2x2_ASAP7_75t_L g770 ( 
.A(n_755),
.B(n_726),
.Y(n_770)
);

OR2x2_ASAP7_75t_L g771 ( 
.A(n_766),
.B(n_735),
.Y(n_771)
);

INVx2_ASAP7_75t_L g772 ( 
.A(n_764),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_767),
.B(n_758),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_769),
.Y(n_774)
);

AND2x4_ASAP7_75t_L g775 ( 
.A(n_772),
.B(n_763),
.Y(n_775)
);

INVx1_ASAP7_75t_SL g776 ( 
.A(n_771),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_769),
.Y(n_777)
);

AND2x4_ASAP7_75t_L g778 ( 
.A(n_768),
.B(n_763),
.Y(n_778)
);

OAI21xp5_ASAP7_75t_L g779 ( 
.A1(n_775),
.A2(n_765),
.B(n_738),
.Y(n_779)
);

AND2x4_ASAP7_75t_L g780 ( 
.A(n_775),
.B(n_763),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_776),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_L g782 ( 
.A(n_774),
.B(n_773),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_L g783 ( 
.A(n_781),
.B(n_777),
.Y(n_783)
);

O2A1O1Ixp33_ASAP7_75t_L g784 ( 
.A1(n_779),
.A2(n_740),
.B(n_744),
.C(n_718),
.Y(n_784)
);

OR2x2_ASAP7_75t_L g785 ( 
.A(n_783),
.B(n_782),
.Y(n_785)
);

AOI222xp33_ASAP7_75t_L g786 ( 
.A1(n_784),
.A2(n_780),
.B1(n_731),
.B2(n_743),
.C1(n_729),
.C2(n_778),
.Y(n_786)
);

OAI31xp33_ASAP7_75t_L g787 ( 
.A1(n_784),
.A2(n_780),
.A3(n_778),
.B(n_712),
.Y(n_787)
);

NOR3xp33_ASAP7_75t_L g788 ( 
.A(n_785),
.B(n_761),
.C(n_729),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_786),
.B(n_787),
.Y(n_789)
);

OAI21xp5_ASAP7_75t_SL g790 ( 
.A1(n_786),
.A2(n_765),
.B(n_734),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_785),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_785),
.Y(n_792)
);

INVx2_ASAP7_75t_L g793 ( 
.A(n_792),
.Y(n_793)
);

NAND3xp33_ASAP7_75t_L g794 ( 
.A(n_789),
.B(n_763),
.C(n_727),
.Y(n_794)
);

AOI22xp5_ASAP7_75t_L g795 ( 
.A1(n_790),
.A2(n_742),
.B1(n_763),
.B2(n_734),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_SL g796 ( 
.A(n_791),
.B(n_734),
.Y(n_796)
);

AND2x2_ASAP7_75t_L g797 ( 
.A(n_788),
.B(n_770),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_SL g798 ( 
.A(n_791),
.B(n_734),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_793),
.Y(n_799)
);

OAI22xp5_ASAP7_75t_L g800 ( 
.A1(n_795),
.A2(n_742),
.B1(n_759),
.B2(n_752),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_794),
.Y(n_801)
);

NAND5xp2_ASAP7_75t_L g802 ( 
.A(n_797),
.B(n_715),
.C(n_757),
.D(n_758),
.E(n_717),
.Y(n_802)
);

O2A1O1Ixp33_ASAP7_75t_L g803 ( 
.A1(n_796),
.A2(n_752),
.B(n_754),
.C(n_735),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_L g804 ( 
.A(n_801),
.B(n_798),
.Y(n_804)
);

NAND4xp75_ASAP7_75t_L g805 ( 
.A(n_799),
.B(n_757),
.C(n_754),
.D(n_762),
.Y(n_805)
);

NAND4xp75_ASAP7_75t_L g806 ( 
.A(n_803),
.B(n_756),
.C(n_719),
.D(n_707),
.Y(n_806)
);

NOR4xp25_ASAP7_75t_L g807 ( 
.A(n_800),
.B(n_759),
.C(n_756),
.D(n_760),
.Y(n_807)
);

O2A1O1Ixp33_ASAP7_75t_L g808 ( 
.A1(n_802),
.A2(n_725),
.B(n_764),
.C(n_760),
.Y(n_808)
);

NAND2xp33_ASAP7_75t_L g809 ( 
.A(n_801),
.B(n_719),
.Y(n_809)
);

OAI21xp33_ASAP7_75t_L g810 ( 
.A1(n_804),
.A2(n_764),
.B(n_711),
.Y(n_810)
);

HB1xp67_ASAP7_75t_L g811 ( 
.A(n_805),
.Y(n_811)
);

OR3x1_ASAP7_75t_L g812 ( 
.A(n_809),
.B(n_707),
.C(n_747),
.Y(n_812)
);

AOI221xp5_ASAP7_75t_L g813 ( 
.A1(n_807),
.A2(n_808),
.B1(n_806),
.B2(n_725),
.C(n_741),
.Y(n_813)
);

HB1xp67_ASAP7_75t_L g814 ( 
.A(n_804),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_814),
.Y(n_815)
);

CKINVDCx5p33_ASAP7_75t_R g816 ( 
.A(n_811),
.Y(n_816)
);

CKINVDCx5p33_ASAP7_75t_R g817 ( 
.A(n_810),
.Y(n_817)
);

AOI211xp5_ASAP7_75t_L g818 ( 
.A1(n_813),
.A2(n_741),
.B(n_736),
.C(n_725),
.Y(n_818)
);

CKINVDCx5p33_ASAP7_75t_R g819 ( 
.A(n_812),
.Y(n_819)
);

AND2x4_ASAP7_75t_L g820 ( 
.A(n_814),
.B(n_711),
.Y(n_820)
);

INVx2_ASAP7_75t_L g821 ( 
.A(n_815),
.Y(n_821)
);

NAND3xp33_ASAP7_75t_L g822 ( 
.A(n_821),
.B(n_816),
.C(n_817),
.Y(n_822)
);

AOI22xp33_ASAP7_75t_SL g823 ( 
.A1(n_822),
.A2(n_819),
.B1(n_820),
.B2(n_818),
.Y(n_823)
);

OAI22xp5_ASAP7_75t_L g824 ( 
.A1(n_823),
.A2(n_725),
.B1(n_711),
.B2(n_750),
.Y(n_824)
);

AOI21x1_ASAP7_75t_L g825 ( 
.A1(n_824),
.A2(n_750),
.B(n_717),
.Y(n_825)
);

AOI22xp33_ASAP7_75t_SL g826 ( 
.A1(n_825),
.A2(n_753),
.B1(n_751),
.B2(n_750),
.Y(n_826)
);

AOI22xp33_ASAP7_75t_L g827 ( 
.A1(n_826),
.A2(n_751),
.B1(n_753),
.B2(n_709),
.Y(n_827)
);

AOI211xp5_ASAP7_75t_L g828 ( 
.A1(n_827),
.A2(n_709),
.B(n_710),
.C(n_716),
.Y(n_828)
);


endmodule