module fake_netlist_5_2329_n_971 (n_137, n_210, n_168, n_164, n_191, n_91, n_208, n_82, n_122, n_194, n_142, n_176, n_10, n_214, n_140, n_24, n_124, n_86, n_136, n_146, n_182, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_180, n_184, n_226, n_65, n_78, n_74, n_144, n_207, n_114, n_57, n_96, n_37, n_189, n_220, n_165, n_111, n_108, n_213, n_129, n_31, n_13, n_66, n_98, n_177, n_60, n_155, n_152, n_197, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_195, n_42, n_22, n_227, n_1, n_45, n_117, n_46, n_21, n_94, n_203, n_205, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_179, n_125, n_35, n_167, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_225, n_84, n_23, n_202, n_130, n_219, n_157, n_29, n_79, n_193, n_131, n_151, n_47, n_173, n_192, n_25, n_53, n_160, n_198, n_223, n_188, n_190, n_8, n_201, n_158, n_44, n_224, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_228, n_109, n_112, n_212, n_85, n_159, n_163, n_95, n_119, n_183, n_185, n_175, n_169, n_59, n_26, n_133, n_215, n_55, n_196, n_99, n_2, n_211, n_218, n_181, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_178, n_221, n_12, n_67, n_121, n_36, n_76, n_200, n_87, n_150, n_162, n_27, n_170, n_64, n_77, n_102, n_106, n_161, n_209, n_222, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_174, n_186, n_199, n_134, n_187, n_32, n_41, n_104, n_172, n_103, n_56, n_51, n_63, n_97, n_141, n_166, n_11, n_206, n_217, n_171, n_153, n_7, n_15, n_145, n_48, n_204, n_50, n_52, n_88, n_110, n_216, n_971);

input n_137;
input n_210;
input n_168;
input n_164;
input n_191;
input n_91;
input n_208;
input n_82;
input n_122;
input n_194;
input n_142;
input n_176;
input n_10;
input n_214;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_182;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_180;
input n_184;
input n_226;
input n_65;
input n_78;
input n_74;
input n_144;
input n_207;
input n_114;
input n_57;
input n_96;
input n_37;
input n_189;
input n_220;
input n_165;
input n_111;
input n_108;
input n_213;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_177;
input n_60;
input n_155;
input n_152;
input n_197;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_195;
input n_42;
input n_22;
input n_227;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_203;
input n_205;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_179;
input n_125;
input n_35;
input n_167;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_225;
input n_84;
input n_23;
input n_202;
input n_130;
input n_219;
input n_157;
input n_29;
input n_79;
input n_193;
input n_131;
input n_151;
input n_47;
input n_173;
input n_192;
input n_25;
input n_53;
input n_160;
input n_198;
input n_223;
input n_188;
input n_190;
input n_8;
input n_201;
input n_158;
input n_44;
input n_224;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_228;
input n_109;
input n_112;
input n_212;
input n_85;
input n_159;
input n_163;
input n_95;
input n_119;
input n_183;
input n_185;
input n_175;
input n_169;
input n_59;
input n_26;
input n_133;
input n_215;
input n_55;
input n_196;
input n_99;
input n_2;
input n_211;
input n_218;
input n_181;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_178;
input n_221;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_200;
input n_87;
input n_150;
input n_162;
input n_27;
input n_170;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_209;
input n_222;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_174;
input n_186;
input n_199;
input n_134;
input n_187;
input n_32;
input n_41;
input n_104;
input n_172;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_166;
input n_11;
input n_206;
input n_217;
input n_171;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_204;
input n_50;
input n_52;
input n_88;
input n_110;
input n_216;

output n_971;

wire n_924;
wire n_676;
wire n_294;
wire n_431;
wire n_380;
wire n_318;
wire n_419;
wire n_653;
wire n_611;
wire n_444;
wire n_642;
wire n_615;
wire n_469;
wire n_851;
wire n_316;
wire n_785;
wire n_389;
wire n_843;
wire n_855;
wire n_549;
wire n_684;
wire n_850;
wire n_418;
wire n_248;
wire n_315;
wire n_268;
wire n_523;
wire n_451;
wire n_532;
wire n_705;
wire n_619;
wire n_408;
wire n_865;
wire n_913;
wire n_678;
wire n_664;
wire n_376;
wire n_697;
wire n_503;
wire n_967;
wire n_235;
wire n_605;
wire n_776;
wire n_928;
wire n_667;
wire n_515;
wire n_790;
wire n_353;
wire n_351;
wire n_367;
wire n_643;
wire n_620;
wire n_916;
wire n_452;
wire n_885;
wire n_525;
wire n_493;
wire n_397;
wire n_880;
wire n_703;
wire n_698;
wire n_483;
wire n_544;
wire n_683;
wire n_780;
wire n_649;
wire n_552;
wire n_547;
wire n_721;
wire n_841;
wire n_956;
wire n_467;
wire n_564;
wire n_802;
wire n_423;
wire n_840;
wire n_284;
wire n_245;
wire n_501;
wire n_823;
wire n_725;
wire n_280;
wire n_744;
wire n_590;
wire n_629;
wire n_672;
wire n_873;
wire n_378;
wire n_551;
wire n_762;
wire n_581;
wire n_688;
wire n_382;
wire n_554;
wire n_800;
wire n_898;
wire n_254;
wire n_690;
wire n_583;
wire n_718;
wire n_671;
wire n_819;
wire n_302;
wire n_265;
wire n_526;
wire n_915;
wire n_719;
wire n_293;
wire n_372;
wire n_443;
wire n_244;
wire n_677;
wire n_864;
wire n_859;
wire n_951;
wire n_821;
wire n_714;
wire n_447;
wire n_247;
wire n_314;
wire n_368;
wire n_433;
wire n_604;
wire n_321;
wire n_292;
wire n_909;
wire n_625;
wire n_854;
wire n_949;
wire n_621;
wire n_753;
wire n_455;
wire n_674;
wire n_932;
wire n_417;
wire n_946;
wire n_612;
wire n_385;
wire n_516;
wire n_498;
wire n_933;
wire n_788;
wire n_507;
wire n_497;
wire n_689;
wire n_738;
wire n_912;
wire n_606;
wire n_559;
wire n_275;
wire n_640;
wire n_968;
wire n_252;
wire n_624;
wire n_825;
wire n_295;
wire n_330;
wire n_877;
wire n_508;
wire n_739;
wire n_506;
wire n_737;
wire n_610;
wire n_692;
wire n_755;
wire n_509;
wire n_568;
wire n_936;
wire n_373;
wire n_820;
wire n_757;
wire n_947;
wire n_307;
wire n_633;
wire n_530;
wire n_439;
wire n_556;
wire n_259;
wire n_448;
wire n_758;
wire n_668;
wire n_733;
wire n_375;
wire n_301;
wire n_828;
wire n_779;
wire n_576;
wire n_941;
wire n_929;
wire n_804;
wire n_867;
wire n_537;
wire n_902;
wire n_587;
wire n_945;
wire n_659;
wire n_492;
wire n_792;
wire n_563;
wire n_756;
wire n_878;
wire n_524;
wire n_943;
wire n_399;
wire n_579;
wire n_394;
wire n_250;
wire n_341;
wire n_938;
wire n_741;
wire n_548;
wire n_543;
wire n_260;
wire n_812;
wire n_842;
wire n_298;
wire n_650;
wire n_320;
wire n_694;
wire n_518;
wire n_505;
wire n_286;
wire n_883;
wire n_282;
wire n_752;
wire n_331;
wire n_906;
wire n_905;
wire n_406;
wire n_519;
wire n_470;
wire n_919;
wire n_782;
wire n_908;
wire n_325;
wire n_449;
wire n_862;
wire n_900;
wire n_724;
wire n_856;
wire n_546;
wire n_760;
wire n_658;
wire n_281;
wire n_918;
wire n_240;
wire n_942;
wire n_381;
wire n_291;
wire n_231;
wire n_257;
wire n_390;
wire n_731;
wire n_456;
wire n_371;
wire n_959;
wire n_481;
wire n_535;
wire n_709;
wire n_540;
wire n_317;
wire n_618;
wire n_940;
wire n_896;
wire n_323;
wire n_569;
wire n_769;
wire n_356;
wire n_592;
wire n_920;
wire n_894;
wire n_271;
wire n_934;
wire n_831;
wire n_826;
wire n_335;
wire n_886;
wire n_964;
wire n_654;
wire n_370;
wire n_234;
wire n_343;
wire n_308;
wire n_379;
wire n_428;
wire n_267;
wire n_514;
wire n_570;
wire n_833;
wire n_457;
wire n_297;
wire n_853;
wire n_603;
wire n_377;
wire n_751;
wire n_484;
wire n_775;
wire n_442;
wire n_814;
wire n_636;
wire n_786;
wire n_600;
wire n_660;
wire n_392;
wire n_655;
wire n_704;
wire n_787;
wire n_264;
wire n_669;
wire n_472;
wire n_750;
wire n_742;
wire n_454;
wire n_961;
wire n_955;
wire n_387;
wire n_771;
wire n_374;
wire n_276;
wire n_339;
wire n_882;
wire n_243;
wire n_398;
wire n_396;
wire n_635;
wire n_347;
wire n_763;
wire n_550;
wire n_522;
wire n_255;
wire n_696;
wire n_897;
wire n_350;
wire n_798;
wire n_662;
wire n_459;
wire n_646;
wire n_962;
wire n_400;
wire n_930;
wire n_436;
wire n_290;
wire n_580;
wire n_622;
wire n_723;
wire n_386;
wire n_578;
wire n_926;
wire n_287;
wire n_344;
wire n_848;
wire n_555;
wire n_783;
wire n_473;
wire n_422;
wire n_475;
wire n_777;
wire n_661;
wire n_682;
wire n_415;
wire n_485;
wire n_496;
wire n_355;
wire n_958;
wire n_849;
wire n_670;
wire n_486;
wire n_816;
wire n_336;
wire n_584;
wire n_681;
wire n_591;
wire n_922;
wire n_521;
wire n_614;
wire n_663;
wire n_845;
wire n_430;
wire n_337;
wire n_313;
wire n_631;
wire n_673;
wire n_837;
wire n_479;
wire n_528;
wire n_510;
wire n_680;
wire n_395;
wire n_553;
wire n_727;
wire n_839;
wire n_432;
wire n_901;
wire n_311;
wire n_813;
wire n_957;
wire n_830;
wire n_773;
wire n_743;
wire n_328;
wire n_801;
wire n_299;
wire n_303;
wire n_369;
wire n_675;
wire n_888;
wire n_296;
wire n_613;
wire n_871;
wire n_241;
wire n_637;
wire n_357;
wire n_875;
wire n_598;
wire n_685;
wire n_608;
wire n_446;
wire n_445;
wire n_749;
wire n_829;
wire n_858;
wire n_923;
wire n_772;
wire n_691;
wire n_881;
wire n_717;
wire n_468;
wire n_499;
wire n_939;
wire n_342;
wire n_482;
wire n_517;
wire n_588;
wire n_361;
wire n_464;
wire n_789;
wire n_363;
wire n_413;
wire n_402;
wire n_734;
wire n_638;
wire n_700;
wire n_796;
wire n_573;
wire n_866;
wire n_969;
wire n_236;
wire n_388;
wire n_761;
wire n_249;
wire n_903;
wire n_740;
wire n_304;
wire n_329;
wire n_274;
wire n_577;
wire n_384;
wire n_582;
wire n_460;
wire n_889;
wire n_277;
wire n_477;
wire n_571;
wire n_461;
wire n_333;
wire n_693;
wire n_338;
wire n_309;
wire n_512;
wire n_836;
wire n_462;
wire n_322;
wire n_567;
wire n_258;
wire n_652;
wire n_778;
wire n_306;
wire n_907;
wire n_722;
wire n_458;
wire n_288;
wire n_770;
wire n_844;
wire n_263;
wire n_471;
wire n_609;
wire n_852;
wire n_283;
wire n_383;
wire n_711;
wire n_781;
wire n_834;
wire n_474;
wire n_765;
wire n_542;
wire n_463;
wire n_488;
wire n_595;
wire n_736;
wire n_502;
wire n_893;
wire n_892;
wire n_891;
wire n_239;
wire n_466;
wire n_420;
wire n_630;
wire n_632;
wire n_489;
wire n_699;
wire n_617;
wire n_310;
wire n_593;
wire n_504;
wire n_511;
wire n_748;
wire n_586;
wire n_846;
wire n_874;
wire n_465;
wire n_838;
wire n_358;
wire n_362;
wire n_876;
wire n_332;
wire n_273;
wire n_585;
wire n_349;
wire n_270;
wire n_616;
wire n_230;
wire n_953;
wire n_601;
wire n_279;
wire n_917;
wire n_966;
wire n_253;
wire n_261;
wire n_289;
wire n_745;
wire n_963;
wire n_954;
wire n_627;
wire n_767;
wire n_440;
wire n_726;
wire n_478;
wire n_793;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_648;
wire n_312;
wire n_476;
wire n_818;
wire n_429;
wire n_861;
wire n_534;
wire n_948;
wire n_884;
wire n_899;
wire n_345;
wire n_944;
wire n_494;
wire n_641;
wire n_628;
wire n_365;
wire n_774;
wire n_730;
wire n_729;
wire n_970;
wire n_911;
wire n_557;
wire n_354;
wire n_575;
wire n_607;
wire n_647;
wire n_480;
wire n_237;
wire n_425;
wire n_513;
wire n_407;
wire n_527;
wire n_795;
wire n_710;
wire n_707;
wire n_832;
wire n_695;
wire n_857;
wire n_560;
wire n_656;
wire n_340;
wire n_561;
wire n_346;
wire n_937;
wire n_393;
wire n_229;
wire n_487;
wire n_495;
wire n_602;
wire n_665;
wire n_574;
wire n_437;
wire n_403;
wire n_453;
wire n_421;
wire n_879;
wire n_720;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_863;
wire n_910;
wire n_490;
wire n_805;
wire n_326;
wire n_794;
wire n_768;
wire n_921;
wire n_233;
wire n_404;
wire n_686;
wire n_366;
wire n_572;
wire n_712;
wire n_754;
wire n_847;
wire n_815;
wire n_246;
wire n_596;
wire n_410;
wire n_558;
wire n_708;
wire n_269;
wire n_529;
wire n_735;
wire n_702;
wire n_285;
wire n_822;
wire n_412;
wire n_232;
wire n_679;
wire n_327;
wire n_657;
wire n_644;
wire n_728;
wire n_895;
wire n_266;
wire n_272;
wire n_491;
wire n_427;
wire n_791;
wire n_732;
wire n_251;
wire n_352;
wire n_566;
wire n_426;
wire n_520;
wire n_565;
wire n_808;
wire n_409;
wire n_797;
wire n_887;
wire n_589;
wire n_716;
wire n_597;
wire n_500;
wire n_562;
wire n_300;
wire n_651;
wire n_435;
wire n_809;
wire n_870;
wire n_931;
wire n_334;
wire n_599;
wire n_766;
wire n_811;
wire n_952;
wire n_541;
wire n_807;
wire n_391;
wire n_701;
wire n_434;
wire n_645;
wire n_539;
wire n_835;
wire n_538;
wire n_666;
wire n_262;
wire n_803;
wire n_868;
wire n_238;
wire n_639;
wire n_799;
wire n_914;
wire n_687;
wire n_715;
wire n_411;
wire n_414;
wire n_319;
wire n_364;
wire n_965;
wire n_927;
wire n_536;
wire n_531;
wire n_935;
wire n_242;
wire n_817;
wire n_872;
wire n_360;
wire n_594;
wire n_764;
wire n_890;
wire n_960;
wire n_759;
wire n_438;
wire n_806;
wire n_713;
wire n_904;
wire n_869;
wire n_324;
wire n_810;
wire n_634;
wire n_416;
wire n_827;
wire n_401;
wire n_348;
wire n_626;
wire n_925;
wire n_424;
wire n_706;
wire n_746;
wire n_256;
wire n_305;
wire n_533;
wire n_950;
wire n_747;
wire n_278;
wire n_784;

INVx2_ASAP7_75t_L g229 ( 
.A(n_111),
.Y(n_229)
);

INVx2_ASAP7_75t_SL g230 ( 
.A(n_100),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_216),
.Y(n_231)
);

BUFx10_ASAP7_75t_L g232 ( 
.A(n_11),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_124),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_172),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_37),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_25),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_17),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_115),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_101),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_197),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_57),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_102),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_138),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_149),
.Y(n_244)
);

CKINVDCx16_ASAP7_75t_R g245 ( 
.A(n_129),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_13),
.Y(n_246)
);

BUFx8_ASAP7_75t_SL g247 ( 
.A(n_184),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_117),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_167),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_170),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_116),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_113),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_207),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_150),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_225),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_153),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_183),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_7),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_43),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_155),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_147),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_125),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_179),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_3),
.Y(n_264)
);

BUFx10_ASAP7_75t_L g265 ( 
.A(n_65),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_140),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_202),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_94),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_39),
.Y(n_269)
);

BUFx10_ASAP7_75t_L g270 ( 
.A(n_17),
.Y(n_270)
);

BUFx10_ASAP7_75t_L g271 ( 
.A(n_227),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_217),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_157),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_119),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_139),
.Y(n_275)
);

BUFx3_ASAP7_75t_L g276 ( 
.A(n_90),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_143),
.Y(n_277)
);

INVx2_ASAP7_75t_SL g278 ( 
.A(n_112),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_62),
.Y(n_279)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_18),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_224),
.Y(n_281)
);

INVx1_ASAP7_75t_SL g282 ( 
.A(n_173),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_85),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_110),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_26),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_71),
.Y(n_286)
);

BUFx6f_ASAP7_75t_L g287 ( 
.A(n_79),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_151),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_95),
.Y(n_289)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_31),
.Y(n_290)
);

BUFx2_ASAP7_75t_L g291 ( 
.A(n_182),
.Y(n_291)
);

BUFx10_ASAP7_75t_L g292 ( 
.A(n_77),
.Y(n_292)
);

BUFx6f_ASAP7_75t_L g293 ( 
.A(n_44),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_189),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_145),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_208),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_87),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_203),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_160),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_81),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_114),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_222),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_122),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_11),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_162),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_93),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_154),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_130),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_194),
.Y(n_309)
);

INVx2_ASAP7_75t_SL g310 ( 
.A(n_142),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_171),
.Y(n_311)
);

INVx4_ASAP7_75t_R g312 ( 
.A(n_82),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_8),
.Y(n_313)
);

BUFx10_ASAP7_75t_L g314 ( 
.A(n_0),
.Y(n_314)
);

HB1xp67_ASAP7_75t_L g315 ( 
.A(n_92),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_52),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_204),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_164),
.Y(n_318)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_168),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_34),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_188),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_190),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_22),
.Y(n_323)
);

INVx2_ASAP7_75t_SL g324 ( 
.A(n_226),
.Y(n_324)
);

INVx2_ASAP7_75t_SL g325 ( 
.A(n_126),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_177),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_118),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_169),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_20),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_146),
.Y(n_330)
);

INVx2_ASAP7_75t_SL g331 ( 
.A(n_132),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_104),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_16),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_199),
.Y(n_334)
);

BUFx5_ASAP7_75t_L g335 ( 
.A(n_35),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_88),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_103),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_127),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_159),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_37),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_163),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_120),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_61),
.Y(n_343)
);

BUFx10_ASAP7_75t_L g344 ( 
.A(n_166),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_56),
.Y(n_345)
);

BUFx2_ASAP7_75t_L g346 ( 
.A(n_96),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_48),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_152),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_97),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_215),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_22),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_51),
.Y(n_352)
);

BUFx10_ASAP7_75t_L g353 ( 
.A(n_71),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_19),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_133),
.Y(n_355)
);

BUFx10_ASAP7_75t_L g356 ( 
.A(n_54),
.Y(n_356)
);

CKINVDCx20_ASAP7_75t_R g357 ( 
.A(n_91),
.Y(n_357)
);

BUFx10_ASAP7_75t_L g358 ( 
.A(n_49),
.Y(n_358)
);

BUFx10_ASAP7_75t_L g359 ( 
.A(n_128),
.Y(n_359)
);

BUFx3_ASAP7_75t_L g360 ( 
.A(n_9),
.Y(n_360)
);

INVx2_ASAP7_75t_L g361 ( 
.A(n_158),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_76),
.Y(n_362)
);

CKINVDCx20_ASAP7_75t_R g363 ( 
.A(n_201),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_66),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_99),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_83),
.Y(n_366)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_136),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_84),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_66),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_175),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_23),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_137),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_185),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_174),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_0),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_178),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_148),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_141),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_43),
.Y(n_379)
);

BUFx5_ASAP7_75t_L g380 ( 
.A(n_121),
.Y(n_380)
);

CKINVDCx16_ASAP7_75t_R g381 ( 
.A(n_200),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_156),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_191),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_180),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_78),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_74),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_176),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_205),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_86),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_34),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_55),
.Y(n_391)
);

BUFx10_ASAP7_75t_L g392 ( 
.A(n_89),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_123),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_4),
.Y(n_394)
);

BUFx6f_ASAP7_75t_L g395 ( 
.A(n_287),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_231),
.Y(n_396)
);

INVx4_ASAP7_75t_L g397 ( 
.A(n_287),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_335),
.B(n_1),
.Y(n_398)
);

BUFx12f_ASAP7_75t_L g399 ( 
.A(n_232),
.Y(n_399)
);

INVx2_ASAP7_75t_L g400 ( 
.A(n_335),
.Y(n_400)
);

XOR2xp5_ASAP7_75t_L g401 ( 
.A(n_315),
.B(n_2),
.Y(n_401)
);

HB1xp67_ASAP7_75t_L g402 ( 
.A(n_235),
.Y(n_402)
);

AND2x2_ASAP7_75t_L g403 ( 
.A(n_291),
.B(n_2),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_335),
.B(n_4),
.Y(n_404)
);

BUFx2_ASAP7_75t_L g405 ( 
.A(n_360),
.Y(n_405)
);

AND2x4_ASAP7_75t_L g406 ( 
.A(n_276),
.B(n_5),
.Y(n_406)
);

HB1xp67_ASAP7_75t_L g407 ( 
.A(n_236),
.Y(n_407)
);

INVx5_ASAP7_75t_L g408 ( 
.A(n_287),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_335),
.Y(n_409)
);

INVx5_ASAP7_75t_L g410 ( 
.A(n_287),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_335),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_335),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_L g413 ( 
.A(n_346),
.B(n_5),
.Y(n_413)
);

BUFx6f_ASAP7_75t_L g414 ( 
.A(n_276),
.Y(n_414)
);

AND2x6_ASAP7_75t_L g415 ( 
.A(n_229),
.B(n_75),
.Y(n_415)
);

INVx4_ASAP7_75t_L g416 ( 
.A(n_233),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_230),
.B(n_6),
.Y(n_417)
);

BUFx12f_ASAP7_75t_L g418 ( 
.A(n_232),
.Y(n_418)
);

HB1xp67_ASAP7_75t_L g419 ( 
.A(n_246),
.Y(n_419)
);

NOR2xp33_ASAP7_75t_SL g420 ( 
.A(n_245),
.B(n_7),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_278),
.B(n_8),
.Y(n_421)
);

HB1xp67_ASAP7_75t_L g422 ( 
.A(n_258),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_293),
.Y(n_423)
);

AND2x4_ASAP7_75t_L g424 ( 
.A(n_319),
.B(n_9),
.Y(n_424)
);

BUFx3_ASAP7_75t_L g425 ( 
.A(n_271),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_310),
.B(n_10),
.Y(n_426)
);

INVx5_ASAP7_75t_L g427 ( 
.A(n_293),
.Y(n_427)
);

HB1xp67_ASAP7_75t_L g428 ( 
.A(n_259),
.Y(n_428)
);

AND2x4_ASAP7_75t_L g429 ( 
.A(n_319),
.B(n_10),
.Y(n_429)
);

BUFx2_ASAP7_75t_L g430 ( 
.A(n_360),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_293),
.Y(n_431)
);

INVx5_ASAP7_75t_L g432 ( 
.A(n_293),
.Y(n_432)
);

NOR2x1_ASAP7_75t_L g433 ( 
.A(n_361),
.B(n_12),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_280),
.Y(n_434)
);

AND2x4_ASAP7_75t_L g435 ( 
.A(n_361),
.B(n_12),
.Y(n_435)
);

BUFx6f_ASAP7_75t_L g436 ( 
.A(n_367),
.Y(n_436)
);

AND2x4_ASAP7_75t_L g437 ( 
.A(n_367),
.B(n_13),
.Y(n_437)
);

AND2x4_ASAP7_75t_L g438 ( 
.A(n_324),
.B(n_14),
.Y(n_438)
);

BUFx6f_ASAP7_75t_L g439 ( 
.A(n_238),
.Y(n_439)
);

BUFx3_ASAP7_75t_L g440 ( 
.A(n_271),
.Y(n_440)
);

AND2x4_ASAP7_75t_L g441 ( 
.A(n_325),
.B(n_14),
.Y(n_441)
);

AND2x4_ASAP7_75t_L g442 ( 
.A(n_331),
.B(n_15),
.Y(n_442)
);

NOR2xp33_ASAP7_75t_L g443 ( 
.A(n_282),
.B(n_15),
.Y(n_443)
);

BUFx6f_ASAP7_75t_L g444 ( 
.A(n_242),
.Y(n_444)
);

INVx5_ASAP7_75t_L g445 ( 
.A(n_292),
.Y(n_445)
);

AND2x4_ASAP7_75t_L g446 ( 
.A(n_243),
.B(n_18),
.Y(n_446)
);

AND2x4_ASAP7_75t_L g447 ( 
.A(n_244),
.B(n_21),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_234),
.Y(n_448)
);

INVx3_ASAP7_75t_L g449 ( 
.A(n_280),
.Y(n_449)
);

INVx3_ASAP7_75t_L g450 ( 
.A(n_290),
.Y(n_450)
);

BUFx6f_ASAP7_75t_L g451 ( 
.A(n_251),
.Y(n_451)
);

BUFx6f_ASAP7_75t_L g452 ( 
.A(n_252),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_290),
.Y(n_453)
);

INVxp67_ASAP7_75t_L g454 ( 
.A(n_265),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_237),
.Y(n_455)
);

BUFx8_ASAP7_75t_SL g456 ( 
.A(n_247),
.Y(n_456)
);

INVx2_ASAP7_75t_L g457 ( 
.A(n_380),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_241),
.B(n_24),
.Y(n_458)
);

AND2x2_ASAP7_75t_L g459 ( 
.A(n_381),
.B(n_344),
.Y(n_459)
);

AND2x4_ASAP7_75t_L g460 ( 
.A(n_257),
.B(n_24),
.Y(n_460)
);

INVx5_ASAP7_75t_L g461 ( 
.A(n_344),
.Y(n_461)
);

NOR2xp33_ASAP7_75t_L g462 ( 
.A(n_263),
.B(n_27),
.Y(n_462)
);

CKINVDCx11_ASAP7_75t_R g463 ( 
.A(n_265),
.Y(n_463)
);

INVx3_ASAP7_75t_L g464 ( 
.A(n_270),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_264),
.Y(n_465)
);

AND2x4_ASAP7_75t_L g466 ( 
.A(n_267),
.B(n_268),
.Y(n_466)
);

BUFx12f_ASAP7_75t_L g467 ( 
.A(n_314),
.Y(n_467)
);

BUFx2_ASAP7_75t_L g468 ( 
.A(n_285),
.Y(n_468)
);

AND2x4_ASAP7_75t_L g469 ( 
.A(n_273),
.B(n_28),
.Y(n_469)
);

AND2x4_ASAP7_75t_L g470 ( 
.A(n_275),
.B(n_28),
.Y(n_470)
);

BUFx6f_ASAP7_75t_L g471 ( 
.A(n_281),
.Y(n_471)
);

INVx3_ASAP7_75t_L g472 ( 
.A(n_353),
.Y(n_472)
);

NOR2xp33_ASAP7_75t_L g473 ( 
.A(n_283),
.B(n_284),
.Y(n_473)
);

HB1xp67_ASAP7_75t_L g474 ( 
.A(n_286),
.Y(n_474)
);

CKINVDCx20_ASAP7_75t_R g475 ( 
.A(n_262),
.Y(n_475)
);

INVx5_ASAP7_75t_L g476 ( 
.A(n_359),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_269),
.B(n_29),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_394),
.Y(n_478)
);

INVx5_ASAP7_75t_L g479 ( 
.A(n_392),
.Y(n_479)
);

AND2x4_ASAP7_75t_L g480 ( 
.A(n_288),
.B(n_30),
.Y(n_480)
);

AND2x4_ASAP7_75t_L g481 ( 
.A(n_289),
.B(n_31),
.Y(n_481)
);

CKINVDCx5p33_ASAP7_75t_R g482 ( 
.A(n_239),
.Y(n_482)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_279),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_304),
.B(n_313),
.Y(n_484)
);

INVx5_ASAP7_75t_L g485 ( 
.A(n_392),
.Y(n_485)
);

INVx2_ASAP7_75t_L g486 ( 
.A(n_333),
.Y(n_486)
);

INVx3_ASAP7_75t_L g487 ( 
.A(n_356),
.Y(n_487)
);

BUFx6f_ASAP7_75t_L g488 ( 
.A(n_299),
.Y(n_488)
);

AND2x4_ASAP7_75t_L g489 ( 
.A(n_301),
.B(n_32),
.Y(n_489)
);

BUFx6f_ASAP7_75t_L g490 ( 
.A(n_303),
.Y(n_490)
);

INVx2_ASAP7_75t_L g491 ( 
.A(n_340),
.Y(n_491)
);

AND2x4_ASAP7_75t_L g492 ( 
.A(n_305),
.B(n_33),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_343),
.B(n_36),
.Y(n_493)
);

BUFx6f_ASAP7_75t_L g494 ( 
.A(n_318),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_351),
.B(n_38),
.Y(n_495)
);

INVx5_ASAP7_75t_L g496 ( 
.A(n_358),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_352),
.Y(n_497)
);

AND2x4_ASAP7_75t_L g498 ( 
.A(n_326),
.B(n_39),
.Y(n_498)
);

AND2x4_ASAP7_75t_L g499 ( 
.A(n_336),
.B(n_40),
.Y(n_499)
);

NOR2xp33_ASAP7_75t_L g500 ( 
.A(n_339),
.B(n_40),
.Y(n_500)
);

NOR2xp33_ASAP7_75t_L g501 ( 
.A(n_342),
.B(n_41),
.Y(n_501)
);

BUFx6f_ASAP7_75t_L g502 ( 
.A(n_348),
.Y(n_502)
);

BUFx2_ASAP7_75t_L g503 ( 
.A(n_316),
.Y(n_503)
);

INVx2_ASAP7_75t_SL g504 ( 
.A(n_320),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_349),
.B(n_42),
.Y(n_505)
);

AND2x6_ASAP7_75t_L g506 ( 
.A(n_355),
.B(n_80),
.Y(n_506)
);

INVx5_ASAP7_75t_L g507 ( 
.A(n_312),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_364),
.Y(n_508)
);

NOR2xp33_ASAP7_75t_SL g509 ( 
.A(n_323),
.B(n_45),
.Y(n_509)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_395),
.Y(n_510)
);

AND2x2_ASAP7_75t_L g511 ( 
.A(n_507),
.B(n_240),
.Y(n_511)
);

AND2x2_ASAP7_75t_L g512 ( 
.A(n_507),
.B(n_459),
.Y(n_512)
);

AOI22xp5_ASAP7_75t_L g513 ( 
.A1(n_413),
.A2(n_302),
.B1(n_327),
.B2(n_308),
.Y(n_513)
);

INVx2_ASAP7_75t_L g514 ( 
.A(n_395),
.Y(n_514)
);

AO22x2_ASAP7_75t_L g515 ( 
.A1(n_401),
.A2(n_386),
.B1(n_391),
.B2(n_375),
.Y(n_515)
);

OAI22xp33_ASAP7_75t_L g516 ( 
.A1(n_420),
.A2(n_329),
.B1(n_347),
.B2(n_345),
.Y(n_516)
);

AND2x2_ASAP7_75t_L g517 ( 
.A(n_507),
.B(n_248),
.Y(n_517)
);

AOI22xp5_ASAP7_75t_L g518 ( 
.A1(n_509),
.A2(n_363),
.B1(n_357),
.B2(n_266),
.Y(n_518)
);

INVx2_ASAP7_75t_L g519 ( 
.A(n_395),
.Y(n_519)
);

AO22x2_ASAP7_75t_L g520 ( 
.A1(n_406),
.A2(n_365),
.B1(n_372),
.B2(n_362),
.Y(n_520)
);

AND2x2_ASAP7_75t_L g521 ( 
.A(n_402),
.B(n_249),
.Y(n_521)
);

AND2x2_ASAP7_75t_L g522 ( 
.A(n_407),
.B(n_250),
.Y(n_522)
);

NOR2xp33_ASAP7_75t_L g523 ( 
.A(n_416),
.B(n_374),
.Y(n_523)
);

OAI22xp33_ASAP7_75t_L g524 ( 
.A1(n_454),
.A2(n_369),
.B1(n_371),
.B2(n_354),
.Y(n_524)
);

INVx2_ASAP7_75t_SL g525 ( 
.A(n_496),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_423),
.Y(n_526)
);

AOI22xp5_ASAP7_75t_L g527 ( 
.A1(n_443),
.A2(n_390),
.B1(n_379),
.B2(n_254),
.Y(n_527)
);

AND2x2_ASAP7_75t_L g528 ( 
.A(n_419),
.B(n_253),
.Y(n_528)
);

AND2x2_ASAP7_75t_L g529 ( 
.A(n_422),
.B(n_255),
.Y(n_529)
);

OR2x2_ASAP7_75t_L g530 ( 
.A(n_464),
.B(n_46),
.Y(n_530)
);

BUFx10_ASAP7_75t_L g531 ( 
.A(n_396),
.Y(n_531)
);

AND2x2_ASAP7_75t_L g532 ( 
.A(n_428),
.B(n_256),
.Y(n_532)
);

AND2x2_ASAP7_75t_L g533 ( 
.A(n_474),
.B(n_260),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_L g534 ( 
.A(n_448),
.B(n_376),
.Y(n_534)
);

AND2x2_ASAP7_75t_L g535 ( 
.A(n_468),
.B(n_261),
.Y(n_535)
);

OAI22xp33_ASAP7_75t_L g536 ( 
.A1(n_464),
.A2(n_384),
.B1(n_385),
.B2(n_377),
.Y(n_536)
);

AO22x2_ASAP7_75t_L g537 ( 
.A1(n_403),
.A2(n_387),
.B1(n_48),
.B2(n_46),
.Y(n_537)
);

AO22x2_ASAP7_75t_L g538 ( 
.A1(n_438),
.A2(n_50),
.B1(n_47),
.B2(n_49),
.Y(n_538)
);

HB1xp67_ASAP7_75t_L g539 ( 
.A(n_496),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_431),
.Y(n_540)
);

AOI22xp5_ASAP7_75t_L g541 ( 
.A1(n_462),
.A2(n_274),
.B1(n_277),
.B2(n_272),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_431),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_409),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_L g544 ( 
.A(n_482),
.B(n_393),
.Y(n_544)
);

INVx2_ASAP7_75t_L g545 ( 
.A(n_400),
.Y(n_545)
);

CKINVDCx16_ASAP7_75t_R g546 ( 
.A(n_475),
.Y(n_546)
);

INVx3_ASAP7_75t_L g547 ( 
.A(n_414),
.Y(n_547)
);

INVx2_ASAP7_75t_SL g548 ( 
.A(n_496),
.Y(n_548)
);

AO22x2_ASAP7_75t_L g549 ( 
.A1(n_438),
.A2(n_51),
.B1(n_47),
.B2(n_50),
.Y(n_549)
);

BUFx10_ASAP7_75t_L g550 ( 
.A(n_473),
.Y(n_550)
);

CKINVDCx5p33_ASAP7_75t_R g551 ( 
.A(n_456),
.Y(n_551)
);

OAI22xp5_ASAP7_75t_L g552 ( 
.A1(n_503),
.A2(n_295),
.B1(n_296),
.B2(n_294),
.Y(n_552)
);

AND2x2_ASAP7_75t_L g553 ( 
.A(n_504),
.B(n_297),
.Y(n_553)
);

AND2x2_ASAP7_75t_L g554 ( 
.A(n_445),
.B(n_298),
.Y(n_554)
);

OR2x6_ASAP7_75t_L g555 ( 
.A(n_399),
.B(n_418),
.Y(n_555)
);

NOR2xp33_ASAP7_75t_L g556 ( 
.A(n_416),
.B(n_300),
.Y(n_556)
);

AOI22xp5_ASAP7_75t_L g557 ( 
.A1(n_500),
.A2(n_350),
.B1(n_388),
.B2(n_383),
.Y(n_557)
);

OAI22xp33_ASAP7_75t_L g558 ( 
.A1(n_472),
.A2(n_389),
.B1(n_382),
.B2(n_378),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_411),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_L g560 ( 
.A(n_445),
.B(n_306),
.Y(n_560)
);

INVx2_ASAP7_75t_L g561 ( 
.A(n_414),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_L g562 ( 
.A(n_461),
.B(n_373),
.Y(n_562)
);

AND2x2_ASAP7_75t_L g563 ( 
.A(n_461),
.B(n_307),
.Y(n_563)
);

AO22x2_ASAP7_75t_L g564 ( 
.A1(n_441),
.A2(n_53),
.B1(n_54),
.B2(n_56),
.Y(n_564)
);

NOR2xp33_ASAP7_75t_L g565 ( 
.A(n_417),
.B(n_309),
.Y(n_565)
);

INVx3_ASAP7_75t_L g566 ( 
.A(n_414),
.Y(n_566)
);

AND2x2_ASAP7_75t_L g567 ( 
.A(n_476),
.B(n_311),
.Y(n_567)
);

OA22x2_ASAP7_75t_L g568 ( 
.A1(n_405),
.A2(n_430),
.B1(n_487),
.B2(n_472),
.Y(n_568)
);

BUFx4f_ASAP7_75t_L g569 ( 
.A(n_415),
.Y(n_569)
);

XOR2xp5_ASAP7_75t_L g570 ( 
.A(n_425),
.B(n_317),
.Y(n_570)
);

AND2x2_ASAP7_75t_L g571 ( 
.A(n_476),
.B(n_321),
.Y(n_571)
);

NOR2xp33_ASAP7_75t_L g572 ( 
.A(n_421),
.B(n_322),
.Y(n_572)
);

OAI22xp33_ASAP7_75t_L g573 ( 
.A1(n_487),
.A2(n_370),
.B1(n_368),
.B2(n_366),
.Y(n_573)
);

AO22x2_ASAP7_75t_L g574 ( 
.A1(n_441),
.A2(n_53),
.B1(n_58),
.B2(n_59),
.Y(n_574)
);

OAI22xp5_ASAP7_75t_SL g575 ( 
.A1(n_458),
.A2(n_493),
.B1(n_495),
.B2(n_477),
.Y(n_575)
);

INVx2_ASAP7_75t_L g576 ( 
.A(n_436),
.Y(n_576)
);

OR2x2_ASAP7_75t_L g577 ( 
.A(n_440),
.B(n_58),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_L g578 ( 
.A(n_479),
.B(n_328),
.Y(n_578)
);

AO22x2_ASAP7_75t_L g579 ( 
.A1(n_442),
.A2(n_59),
.B1(n_60),
.B2(n_61),
.Y(n_579)
);

AND2x2_ASAP7_75t_L g580 ( 
.A(n_479),
.B(n_330),
.Y(n_580)
);

AO22x2_ASAP7_75t_L g581 ( 
.A1(n_442),
.A2(n_60),
.B1(n_63),
.B2(n_64),
.Y(n_581)
);

AND2x2_ASAP7_75t_L g582 ( 
.A(n_485),
.B(n_332),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_411),
.Y(n_583)
);

AND2x2_ASAP7_75t_SL g584 ( 
.A(n_424),
.B(n_63),
.Y(n_584)
);

AND2x2_ASAP7_75t_L g585 ( 
.A(n_485),
.B(n_334),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_543),
.Y(n_586)
);

XNOR2x2_ASAP7_75t_L g587 ( 
.A(n_518),
.B(n_433),
.Y(n_587)
);

INVx2_ASAP7_75t_L g588 ( 
.A(n_576),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_559),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_559),
.Y(n_590)
);

BUFx3_ASAP7_75t_L g591 ( 
.A(n_547),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_L g592 ( 
.A(n_583),
.B(n_466),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_583),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_566),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_566),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_510),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_514),
.Y(n_597)
);

NAND2x1p5_ASAP7_75t_L g598 ( 
.A(n_569),
.B(n_433),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_519),
.Y(n_599)
);

INVx8_ASAP7_75t_L g600 ( 
.A(n_512),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_561),
.Y(n_601)
);

NAND2xp33_ASAP7_75t_SL g602 ( 
.A(n_575),
.B(n_426),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_545),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_526),
.Y(n_604)
);

OAI21xp5_ASAP7_75t_L g605 ( 
.A1(n_534),
.A2(n_404),
.B(n_398),
.Y(n_605)
);

XOR2xp5_ASAP7_75t_L g606 ( 
.A(n_546),
.B(n_337),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_540),
.Y(n_607)
);

NOR2xp33_ASAP7_75t_L g608 ( 
.A(n_550),
.B(n_516),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_540),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_L g610 ( 
.A(n_542),
.B(n_466),
.Y(n_610)
);

AND2x6_ASAP7_75t_L g611 ( 
.A(n_553),
.B(n_424),
.Y(n_611)
);

INVxp67_ASAP7_75t_SL g612 ( 
.A(n_530),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_568),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_577),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_521),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_522),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_528),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_529),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_532),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_533),
.Y(n_620)
);

CKINVDCx5p33_ASAP7_75t_R g621 ( 
.A(n_531),
.Y(n_621)
);

AND2x2_ASAP7_75t_SL g622 ( 
.A(n_584),
.B(n_429),
.Y(n_622)
);

AND2x2_ASAP7_75t_L g623 ( 
.A(n_535),
.B(n_463),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_520),
.Y(n_624)
);

NAND2xp33_ASAP7_75t_R g625 ( 
.A(n_551),
.B(n_446),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_554),
.Y(n_626)
);

CKINVDCx16_ASAP7_75t_R g627 ( 
.A(n_513),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_563),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_567),
.Y(n_629)
);

XNOR2x2_ASAP7_75t_L g630 ( 
.A(n_538),
.B(n_477),
.Y(n_630)
);

OR2x6_ASAP7_75t_L g631 ( 
.A(n_538),
.B(n_467),
.Y(n_631)
);

NOR2xp33_ASAP7_75t_L g632 ( 
.A(n_565),
.B(n_439),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_571),
.Y(n_633)
);

INVxp33_ASAP7_75t_SL g634 ( 
.A(n_570),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_580),
.Y(n_635)
);

INVx2_ASAP7_75t_L g636 ( 
.A(n_511),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_582),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_585),
.Y(n_638)
);

OR2x2_ASAP7_75t_L g639 ( 
.A(n_527),
.B(n_505),
.Y(n_639)
);

AND2x2_ASAP7_75t_L g640 ( 
.A(n_525),
.B(n_449),
.Y(n_640)
);

NOR2xp33_ASAP7_75t_L g641 ( 
.A(n_572),
.B(n_439),
.Y(n_641)
);

INVx2_ASAP7_75t_L g642 ( 
.A(n_517),
.Y(n_642)
);

NOR2xp33_ASAP7_75t_L g643 ( 
.A(n_544),
.B(n_439),
.Y(n_643)
);

INVx2_ASAP7_75t_L g644 ( 
.A(n_548),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_L g645 ( 
.A(n_523),
.B(n_412),
.Y(n_645)
);

INVxp67_ASAP7_75t_L g646 ( 
.A(n_539),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_560),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_562),
.Y(n_648)
);

NOR2xp33_ASAP7_75t_L g649 ( 
.A(n_527),
.B(n_444),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_578),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_549),
.Y(n_651)
);

INVx2_ASAP7_75t_SL g652 ( 
.A(n_552),
.Y(n_652)
);

INVx2_ASAP7_75t_L g653 ( 
.A(n_549),
.Y(n_653)
);

AND2x2_ASAP7_75t_L g654 ( 
.A(n_605),
.B(n_537),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_632),
.B(n_556),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_632),
.B(n_541),
.Y(n_656)
);

INVx4_ASAP7_75t_L g657 ( 
.A(n_611),
.Y(n_657)
);

HB1xp67_ASAP7_75t_L g658 ( 
.A(n_613),
.Y(n_658)
);

AND2x2_ASAP7_75t_L g659 ( 
.A(n_612),
.B(n_622),
.Y(n_659)
);

INVx2_ASAP7_75t_L g660 ( 
.A(n_586),
.Y(n_660)
);

BUFx3_ASAP7_75t_L g661 ( 
.A(n_600),
.Y(n_661)
);

INVx2_ASAP7_75t_L g662 ( 
.A(n_589),
.Y(n_662)
);

INVx2_ASAP7_75t_L g663 ( 
.A(n_590),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_593),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_L g665 ( 
.A(n_641),
.B(n_541),
.Y(n_665)
);

INVx2_ASAP7_75t_L g666 ( 
.A(n_604),
.Y(n_666)
);

INVx2_ASAP7_75t_L g667 ( 
.A(n_607),
.Y(n_667)
);

INVx3_ASAP7_75t_L g668 ( 
.A(n_588),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_609),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_592),
.Y(n_670)
);

INVx2_ASAP7_75t_SL g671 ( 
.A(n_640),
.Y(n_671)
);

BUFx3_ASAP7_75t_L g672 ( 
.A(n_600),
.Y(n_672)
);

AND2x2_ASAP7_75t_L g673 ( 
.A(n_649),
.B(n_564),
.Y(n_673)
);

INVx4_ASAP7_75t_SL g674 ( 
.A(n_611),
.Y(n_674)
);

AND2x2_ASAP7_75t_L g675 ( 
.A(n_649),
.B(n_574),
.Y(n_675)
);

AND2x2_ASAP7_75t_L g676 ( 
.A(n_636),
.B(n_642),
.Y(n_676)
);

AND2x2_ASAP7_75t_L g677 ( 
.A(n_645),
.B(n_615),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_592),
.Y(n_678)
);

AND2x4_ASAP7_75t_L g679 ( 
.A(n_626),
.B(n_506),
.Y(n_679)
);

BUFx3_ASAP7_75t_L g680 ( 
.A(n_600),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_L g681 ( 
.A(n_643),
.B(n_557),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_603),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_610),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_647),
.B(n_506),
.Y(n_684)
);

BUFx6f_ASAP7_75t_L g685 ( 
.A(n_598),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_610),
.Y(n_686)
);

AND2x4_ASAP7_75t_L g687 ( 
.A(n_628),
.B(n_506),
.Y(n_687)
);

INVx2_ASAP7_75t_L g688 ( 
.A(n_596),
.Y(n_688)
);

INVxp67_ASAP7_75t_L g689 ( 
.A(n_608),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_648),
.B(n_506),
.Y(n_690)
);

AND2x6_ASAP7_75t_L g691 ( 
.A(n_651),
.B(n_435),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_L g692 ( 
.A(n_650),
.B(n_558),
.Y(n_692)
);

AND2x2_ASAP7_75t_L g693 ( 
.A(n_616),
.B(n_579),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_597),
.Y(n_694)
);

AND2x2_ASAP7_75t_L g695 ( 
.A(n_617),
.B(n_579),
.Y(n_695)
);

BUFx3_ASAP7_75t_L g696 ( 
.A(n_611),
.Y(n_696)
);

INVx2_ASAP7_75t_L g697 ( 
.A(n_599),
.Y(n_697)
);

INVx2_ASAP7_75t_L g698 ( 
.A(n_601),
.Y(n_698)
);

INVx3_ASAP7_75t_L g699 ( 
.A(n_611),
.Y(n_699)
);

AND2x2_ASAP7_75t_L g700 ( 
.A(n_618),
.B(n_581),
.Y(n_700)
);

INVx4_ASAP7_75t_L g701 ( 
.A(n_611),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_L g702 ( 
.A(n_629),
.B(n_573),
.Y(n_702)
);

INVx2_ASAP7_75t_L g703 ( 
.A(n_594),
.Y(n_703)
);

AND2x4_ASAP7_75t_L g704 ( 
.A(n_633),
.B(n_447),
.Y(n_704)
);

INVx3_ASAP7_75t_SL g705 ( 
.A(n_621),
.Y(n_705)
);

INVx2_ASAP7_75t_L g706 ( 
.A(n_595),
.Y(n_706)
);

INVx2_ASAP7_75t_SL g707 ( 
.A(n_635),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_637),
.Y(n_708)
);

AND2x2_ASAP7_75t_L g709 ( 
.A(n_619),
.B(n_581),
.Y(n_709)
);

AND2x2_ASAP7_75t_L g710 ( 
.A(n_620),
.B(n_638),
.Y(n_710)
);

AND2x2_ASAP7_75t_L g711 ( 
.A(n_639),
.B(n_460),
.Y(n_711)
);

INVx2_ASAP7_75t_L g712 ( 
.A(n_591),
.Y(n_712)
);

INVx2_ASAP7_75t_L g713 ( 
.A(n_624),
.Y(n_713)
);

AND2x2_ASAP7_75t_L g714 ( 
.A(n_652),
.B(n_460),
.Y(n_714)
);

AOI22xp5_ASAP7_75t_L g715 ( 
.A1(n_602),
.A2(n_501),
.B1(n_469),
.B2(n_470),
.Y(n_715)
);

NOR2xp33_ASAP7_75t_L g716 ( 
.A(n_608),
.B(n_524),
.Y(n_716)
);

INVx2_ASAP7_75t_L g717 ( 
.A(n_644),
.Y(n_717)
);

BUFx3_ASAP7_75t_L g718 ( 
.A(n_653),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_587),
.Y(n_719)
);

BUFx3_ASAP7_75t_L g720 ( 
.A(n_630),
.Y(n_720)
);

AND2x2_ASAP7_75t_SL g721 ( 
.A(n_627),
.B(n_437),
.Y(n_721)
);

AND2x2_ASAP7_75t_L g722 ( 
.A(n_614),
.B(n_470),
.Y(n_722)
);

BUFx3_ASAP7_75t_L g723 ( 
.A(n_631),
.Y(n_723)
);

INVx2_ASAP7_75t_L g724 ( 
.A(n_660),
.Y(n_724)
);

BUFx3_ASAP7_75t_L g725 ( 
.A(n_705),
.Y(n_725)
);

NOR2x1_ASAP7_75t_L g726 ( 
.A(n_661),
.B(n_623),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_660),
.Y(n_727)
);

AND2x4_ASAP7_75t_L g728 ( 
.A(n_661),
.B(n_646),
.Y(n_728)
);

OR2x2_ASAP7_75t_L g729 ( 
.A(n_689),
.B(n_606),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_655),
.B(n_646),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_L g731 ( 
.A(n_670),
.B(n_678),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_658),
.Y(n_732)
);

BUFx6f_ASAP7_75t_L g733 ( 
.A(n_661),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_L g734 ( 
.A(n_683),
.B(n_480),
.Y(n_734)
);

AND2x4_ASAP7_75t_L g735 ( 
.A(n_672),
.B(n_483),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_664),
.Y(n_736)
);

BUFx6f_ASAP7_75t_L g737 ( 
.A(n_672),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_L g738 ( 
.A(n_683),
.B(n_480),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_669),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_669),
.Y(n_740)
);

AND2x4_ASAP7_75t_L g741 ( 
.A(n_672),
.B(n_486),
.Y(n_741)
);

OR2x6_ASAP7_75t_L g742 ( 
.A(n_723),
.B(n_555),
.Y(n_742)
);

NOR2xp33_ASAP7_75t_L g743 ( 
.A(n_656),
.B(n_634),
.Y(n_743)
);

BUFx6f_ASAP7_75t_L g744 ( 
.A(n_680),
.Y(n_744)
);

AND2x4_ASAP7_75t_L g745 ( 
.A(n_680),
.B(n_491),
.Y(n_745)
);

BUFx4f_ASAP7_75t_L g746 ( 
.A(n_705),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_686),
.B(n_481),
.Y(n_747)
);

INVx5_ASAP7_75t_L g748 ( 
.A(n_685),
.Y(n_748)
);

BUFx6f_ASAP7_75t_L g749 ( 
.A(n_680),
.Y(n_749)
);

BUFx6f_ASAP7_75t_L g750 ( 
.A(n_718),
.Y(n_750)
);

AND2x2_ASAP7_75t_L g751 ( 
.A(n_677),
.B(n_515),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_662),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_L g753 ( 
.A(n_665),
.B(n_489),
.Y(n_753)
);

CKINVDCx11_ASAP7_75t_R g754 ( 
.A(n_723),
.Y(n_754)
);

INVx4_ASAP7_75t_L g755 ( 
.A(n_685),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_L g756 ( 
.A(n_714),
.B(n_492),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_663),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_666),
.Y(n_758)
);

INVx3_ASAP7_75t_L g759 ( 
.A(n_666),
.Y(n_759)
);

INVx4_ASAP7_75t_L g760 ( 
.A(n_685),
.Y(n_760)
);

BUFx6f_ASAP7_75t_L g761 ( 
.A(n_718),
.Y(n_761)
);

BUFx6f_ASAP7_75t_L g762 ( 
.A(n_718),
.Y(n_762)
);

AND2x6_ASAP7_75t_L g763 ( 
.A(n_699),
.B(n_498),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_667),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_667),
.Y(n_765)
);

NAND2x1p5_ASAP7_75t_L g766 ( 
.A(n_685),
.B(n_455),
.Y(n_766)
);

AND2x2_ASAP7_75t_L g767 ( 
.A(n_711),
.B(n_508),
.Y(n_767)
);

AND2x4_ASAP7_75t_L g768 ( 
.A(n_676),
.B(n_712),
.Y(n_768)
);

BUFx6f_ASAP7_75t_L g769 ( 
.A(n_685),
.Y(n_769)
);

NOR2xp33_ASAP7_75t_L g770 ( 
.A(n_716),
.B(n_536),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_681),
.B(n_498),
.Y(n_771)
);

AND2x4_ASAP7_75t_L g772 ( 
.A(n_768),
.B(n_713),
.Y(n_772)
);

INVx5_ASAP7_75t_L g773 ( 
.A(n_769),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_727),
.Y(n_774)
);

INVx2_ASAP7_75t_SL g775 ( 
.A(n_750),
.Y(n_775)
);

INVx4_ASAP7_75t_L g776 ( 
.A(n_748),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_L g777 ( 
.A(n_730),
.B(n_659),
.Y(n_777)
);

BUFx3_ASAP7_75t_L g778 ( 
.A(n_725),
.Y(n_778)
);

INVx5_ASAP7_75t_L g779 ( 
.A(n_769),
.Y(n_779)
);

BUFx6f_ASAP7_75t_L g780 ( 
.A(n_733),
.Y(n_780)
);

BUFx3_ASAP7_75t_L g781 ( 
.A(n_746),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_727),
.Y(n_782)
);

BUFx3_ASAP7_75t_L g783 ( 
.A(n_746),
.Y(n_783)
);

BUFx6f_ASAP7_75t_L g784 ( 
.A(n_733),
.Y(n_784)
);

AND2x4_ASAP7_75t_L g785 ( 
.A(n_768),
.B(n_713),
.Y(n_785)
);

INVx4_ASAP7_75t_L g786 ( 
.A(n_755),
.Y(n_786)
);

INVx3_ASAP7_75t_L g787 ( 
.A(n_755),
.Y(n_787)
);

INVx4_ASAP7_75t_L g788 ( 
.A(n_760),
.Y(n_788)
);

BUFx3_ASAP7_75t_L g789 ( 
.A(n_733),
.Y(n_789)
);

INVx2_ASAP7_75t_L g790 ( 
.A(n_752),
.Y(n_790)
);

INVx4_ASAP7_75t_L g791 ( 
.A(n_760),
.Y(n_791)
);

CKINVDCx14_ASAP7_75t_R g792 ( 
.A(n_754),
.Y(n_792)
);

INVx3_ASAP7_75t_L g793 ( 
.A(n_750),
.Y(n_793)
);

INVx3_ASAP7_75t_L g794 ( 
.A(n_761),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_736),
.Y(n_795)
);

INVx2_ASAP7_75t_SL g796 ( 
.A(n_761),
.Y(n_796)
);

BUFx2_ASAP7_75t_SL g797 ( 
.A(n_737),
.Y(n_797)
);

INVx4_ASAP7_75t_L g798 ( 
.A(n_744),
.Y(n_798)
);

AOI22xp33_ASAP7_75t_L g799 ( 
.A1(n_770),
.A2(n_720),
.B1(n_719),
.B2(n_654),
.Y(n_799)
);

BUFx2_ASAP7_75t_R g800 ( 
.A(n_729),
.Y(n_800)
);

AND2x4_ASAP7_75t_L g801 ( 
.A(n_744),
.B(n_659),
.Y(n_801)
);

INVx4_ASAP7_75t_L g802 ( 
.A(n_749),
.Y(n_802)
);

BUFx6f_ASAP7_75t_L g803 ( 
.A(n_749),
.Y(n_803)
);

INVxp67_ASAP7_75t_SL g804 ( 
.A(n_762),
.Y(n_804)
);

INVx2_ASAP7_75t_SL g805 ( 
.A(n_762),
.Y(n_805)
);

INVx1_ASAP7_75t_SL g806 ( 
.A(n_732),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_739),
.Y(n_807)
);

BUFx4f_ASAP7_75t_L g808 ( 
.A(n_749),
.Y(n_808)
);

INVxp67_ASAP7_75t_SL g809 ( 
.A(n_762),
.Y(n_809)
);

BUFx6f_ASAP7_75t_L g810 ( 
.A(n_766),
.Y(n_810)
);

BUFx2_ASAP7_75t_L g811 ( 
.A(n_728),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_740),
.Y(n_812)
);

BUFx5_ASAP7_75t_L g813 ( 
.A(n_763),
.Y(n_813)
);

INVx1_ASAP7_75t_SL g814 ( 
.A(n_751),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_795),
.Y(n_815)
);

AOI22xp33_ASAP7_75t_L g816 ( 
.A1(n_799),
.A2(n_720),
.B1(n_719),
.B2(n_743),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_807),
.Y(n_817)
);

INVx3_ASAP7_75t_L g818 ( 
.A(n_776),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_812),
.Y(n_819)
);

OAI21xp5_ASAP7_75t_SL g820 ( 
.A1(n_814),
.A2(n_715),
.B(n_675),
.Y(n_820)
);

AOI22xp33_ASAP7_75t_SL g821 ( 
.A1(n_777),
.A2(n_721),
.B1(n_675),
.B2(n_673),
.Y(n_821)
);

AND2x4_ASAP7_75t_L g822 ( 
.A(n_801),
.B(n_735),
.Y(n_822)
);

INVxp67_ASAP7_75t_L g823 ( 
.A(n_806),
.Y(n_823)
);

INVx2_ASAP7_75t_SL g824 ( 
.A(n_778),
.Y(n_824)
);

BUFx6f_ASAP7_75t_L g825 ( 
.A(n_808),
.Y(n_825)
);

BUFx6f_ASAP7_75t_L g826 ( 
.A(n_808),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_774),
.Y(n_827)
);

INVx4_ASAP7_75t_L g828 ( 
.A(n_779),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_782),
.Y(n_829)
);

OAI22xp5_ASAP7_75t_L g830 ( 
.A1(n_790),
.A2(n_731),
.B1(n_753),
.B2(n_771),
.Y(n_830)
);

OAI22xp5_ASAP7_75t_L g831 ( 
.A1(n_790),
.A2(n_738),
.B1(n_747),
.B2(n_734),
.Y(n_831)
);

OAI22xp5_ASAP7_75t_SL g832 ( 
.A1(n_792),
.A2(n_692),
.B1(n_742),
.B2(n_708),
.Y(n_832)
);

AND2x2_ASAP7_75t_L g833 ( 
.A(n_811),
.B(n_767),
.Y(n_833)
);

BUFx6f_ASAP7_75t_L g834 ( 
.A(n_808),
.Y(n_834)
);

OAI21xp33_ASAP7_75t_L g835 ( 
.A1(n_800),
.A2(n_702),
.B(n_710),
.Y(n_835)
);

OAI22xp33_ASAP7_75t_L g836 ( 
.A1(n_781),
.A2(n_707),
.B1(n_625),
.B2(n_756),
.Y(n_836)
);

BUFx3_ASAP7_75t_L g837 ( 
.A(n_783),
.Y(n_837)
);

BUFx4f_ASAP7_75t_SL g838 ( 
.A(n_789),
.Y(n_838)
);

AOI22xp5_ASAP7_75t_L g839 ( 
.A1(n_801),
.A2(n_726),
.B1(n_741),
.B2(n_735),
.Y(n_839)
);

BUFx8_ASAP7_75t_L g840 ( 
.A(n_780),
.Y(n_840)
);

CKINVDCx11_ASAP7_75t_R g841 ( 
.A(n_784),
.Y(n_841)
);

INVx2_ASAP7_75t_L g842 ( 
.A(n_772),
.Y(n_842)
);

AOI22xp33_ASAP7_75t_SL g843 ( 
.A1(n_797),
.A2(n_695),
.B1(n_700),
.B2(n_693),
.Y(n_843)
);

AOI22xp33_ASAP7_75t_L g844 ( 
.A1(n_816),
.A2(n_499),
.B1(n_758),
.B2(n_757),
.Y(n_844)
);

AOI22xp33_ASAP7_75t_SL g845 ( 
.A1(n_832),
.A2(n_810),
.B1(n_745),
.B2(n_700),
.Y(n_845)
);

OAI22xp33_ASAP7_75t_L g846 ( 
.A1(n_820),
.A2(n_765),
.B1(n_764),
.B2(n_724),
.Y(n_846)
);

AND2x2_ASAP7_75t_L g847 ( 
.A(n_833),
.B(n_709),
.Y(n_847)
);

AOI211xp5_ASAP7_75t_L g848 ( 
.A1(n_835),
.A2(n_484),
.B(n_722),
.C(n_478),
.Y(n_848)
);

NOR2xp33_ASAP7_75t_L g849 ( 
.A(n_820),
.B(n_772),
.Y(n_849)
);

AOI22xp33_ASAP7_75t_L g850 ( 
.A1(n_821),
.A2(n_785),
.B1(n_682),
.B2(n_694),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_815),
.Y(n_851)
);

INVx3_ASAP7_75t_L g852 ( 
.A(n_825),
.Y(n_852)
);

NAND2x1_ASAP7_75t_L g853 ( 
.A(n_828),
.B(n_776),
.Y(n_853)
);

AOI22xp33_ASAP7_75t_L g854 ( 
.A1(n_830),
.A2(n_704),
.B1(n_759),
.B2(n_697),
.Y(n_854)
);

INVx3_ASAP7_75t_L g855 ( 
.A(n_826),
.Y(n_855)
);

AOI22xp33_ASAP7_75t_L g856 ( 
.A1(n_830),
.A2(n_759),
.B1(n_697),
.B2(n_698),
.Y(n_856)
);

OAI22xp5_ASAP7_75t_L g857 ( 
.A1(n_839),
.A2(n_696),
.B1(n_809),
.B2(n_804),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_L g858 ( 
.A(n_823),
.B(n_671),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_L g859 ( 
.A(n_822),
.B(n_775),
.Y(n_859)
);

AOI22xp33_ASAP7_75t_L g860 ( 
.A1(n_831),
.A2(n_698),
.B1(n_688),
.B2(n_478),
.Y(n_860)
);

OAI222xp33_ASAP7_75t_L g861 ( 
.A1(n_843),
.A2(n_338),
.B1(n_341),
.B2(n_775),
.C1(n_796),
.C2(n_805),
.Y(n_861)
);

AND2x2_ASAP7_75t_L g862 ( 
.A(n_842),
.B(n_796),
.Y(n_862)
);

OAI22xp33_ASAP7_75t_L g863 ( 
.A1(n_817),
.A2(n_787),
.B1(n_788),
.B2(n_786),
.Y(n_863)
);

AOI22xp33_ASAP7_75t_L g864 ( 
.A1(n_831),
.A2(n_688),
.B1(n_497),
.B2(n_465),
.Y(n_864)
);

OAI221xp5_ASAP7_75t_SL g865 ( 
.A1(n_848),
.A2(n_836),
.B1(n_837),
.B2(n_824),
.C(n_819),
.Y(n_865)
);

AOI22xp33_ASAP7_75t_L g866 ( 
.A1(n_849),
.A2(n_415),
.B1(n_706),
.B2(n_703),
.Y(n_866)
);

AOI22xp33_ASAP7_75t_L g867 ( 
.A1(n_845),
.A2(n_841),
.B1(n_684),
.B2(n_690),
.Y(n_867)
);

AOI22xp33_ASAP7_75t_L g868 ( 
.A1(n_850),
.A2(n_793),
.B1(n_794),
.B2(n_827),
.Y(n_868)
);

AOI22xp33_ASAP7_75t_L g869 ( 
.A1(n_850),
.A2(n_793),
.B1(n_794),
.B2(n_829),
.Y(n_869)
);

AOI22xp33_ASAP7_75t_L g870 ( 
.A1(n_846),
.A2(n_794),
.B1(n_834),
.B2(n_826),
.Y(n_870)
);

AOI22xp33_ASAP7_75t_SL g871 ( 
.A1(n_861),
.A2(n_834),
.B1(n_840),
.B2(n_838),
.Y(n_871)
);

AOI22xp33_ASAP7_75t_L g872 ( 
.A1(n_844),
.A2(n_763),
.B1(n_691),
.B2(n_687),
.Y(n_872)
);

OAI221xp5_ASAP7_75t_L g873 ( 
.A1(n_844),
.A2(n_717),
.B1(n_453),
.B2(n_434),
.C(n_449),
.Y(n_873)
);

NAND3xp33_ASAP7_75t_L g874 ( 
.A(n_864),
.B(n_451),
.C(n_444),
.Y(n_874)
);

AOI22xp33_ASAP7_75t_L g875 ( 
.A1(n_847),
.A2(n_763),
.B1(n_691),
.B2(n_687),
.Y(n_875)
);

AND2x2_ASAP7_75t_L g876 ( 
.A(n_851),
.B(n_784),
.Y(n_876)
);

AOI22xp33_ASAP7_75t_SL g877 ( 
.A1(n_857),
.A2(n_813),
.B1(n_691),
.B2(n_818),
.Y(n_877)
);

NOR2xp33_ASAP7_75t_L g878 ( 
.A(n_858),
.B(n_717),
.Y(n_878)
);

AOI22xp33_ASAP7_75t_L g879 ( 
.A1(n_854),
.A2(n_679),
.B1(n_798),
.B2(n_802),
.Y(n_879)
);

AOI22xp33_ASAP7_75t_L g880 ( 
.A1(n_860),
.A2(n_699),
.B1(n_803),
.B2(n_784),
.Y(n_880)
);

AOI22xp33_ASAP7_75t_L g881 ( 
.A1(n_859),
.A2(n_699),
.B1(n_803),
.B2(n_668),
.Y(n_881)
);

AOI21xp33_ASAP7_75t_L g882 ( 
.A1(n_856),
.A2(n_803),
.B(n_668),
.Y(n_882)
);

OAI221xp5_ASAP7_75t_L g883 ( 
.A1(n_856),
.A2(n_434),
.B1(n_453),
.B2(n_450),
.C(n_791),
.Y(n_883)
);

AOI22xp33_ASAP7_75t_L g884 ( 
.A1(n_862),
.A2(n_668),
.B1(n_813),
.B2(n_657),
.Y(n_884)
);

AOI22xp33_ASAP7_75t_L g885 ( 
.A1(n_852),
.A2(n_701),
.B1(n_452),
.B2(n_502),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_863),
.Y(n_886)
);

AOI22xp33_ASAP7_75t_L g887 ( 
.A1(n_852),
.A2(n_471),
.B1(n_490),
.B2(n_494),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_853),
.Y(n_888)
);

AOI22xp33_ASAP7_75t_L g889 ( 
.A1(n_855),
.A2(n_471),
.B1(n_490),
.B2(n_494),
.Y(n_889)
);

NAND3xp33_ASAP7_75t_L g890 ( 
.A(n_865),
.B(n_488),
.C(n_436),
.Y(n_890)
);

OAI21xp5_ASAP7_75t_SL g891 ( 
.A1(n_871),
.A2(n_450),
.B(n_457),
.Y(n_891)
);

AOI221xp5_ASAP7_75t_L g892 ( 
.A1(n_878),
.A2(n_397),
.B1(n_67),
.B2(n_68),
.C(n_69),
.Y(n_892)
);

OAI221xp5_ASAP7_75t_SL g893 ( 
.A1(n_867),
.A2(n_65),
.B1(n_67),
.B2(n_70),
.C(n_72),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_L g894 ( 
.A(n_876),
.B(n_70),
.Y(n_894)
);

AND2x2_ASAP7_75t_L g895 ( 
.A(n_886),
.B(n_73),
.Y(n_895)
);

OAI22xp33_ASAP7_75t_L g896 ( 
.A1(n_874),
.A2(n_773),
.B1(n_397),
.B2(n_410),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_SL g897 ( 
.A(n_870),
.B(n_773),
.Y(n_897)
);

AOI221xp5_ASAP7_75t_L g898 ( 
.A1(n_868),
.A2(n_432),
.B1(n_427),
.B2(n_410),
.C(n_408),
.Y(n_898)
);

OAI21xp5_ASAP7_75t_L g899 ( 
.A1(n_866),
.A2(n_432),
.B(n_427),
.Y(n_899)
);

AOI22xp5_ASAP7_75t_L g900 ( 
.A1(n_877),
.A2(n_674),
.B1(n_427),
.B2(n_410),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_869),
.B(n_98),
.Y(n_901)
);

AND2x2_ASAP7_75t_L g902 ( 
.A(n_888),
.B(n_105),
.Y(n_902)
);

OAI221xp5_ASAP7_75t_SL g903 ( 
.A1(n_872),
.A2(n_106),
.B1(n_107),
.B2(n_108),
.C(n_109),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_879),
.B(n_131),
.Y(n_904)
);

AOI221xp5_ASAP7_75t_L g905 ( 
.A1(n_893),
.A2(n_873),
.B1(n_883),
.B2(n_880),
.C(n_882),
.Y(n_905)
);

NAND3xp33_ASAP7_75t_L g906 ( 
.A(n_892),
.B(n_889),
.C(n_887),
.Y(n_906)
);

NAND3xp33_ASAP7_75t_L g907 ( 
.A(n_890),
.B(n_875),
.C(n_881),
.Y(n_907)
);

NOR3xp33_ASAP7_75t_L g908 ( 
.A(n_903),
.B(n_884),
.C(n_885),
.Y(n_908)
);

NOR3xp33_ASAP7_75t_L g909 ( 
.A(n_891),
.B(n_134),
.C(n_135),
.Y(n_909)
);

INVxp67_ASAP7_75t_L g910 ( 
.A(n_894),
.Y(n_910)
);

INVx2_ASAP7_75t_L g911 ( 
.A(n_902),
.Y(n_911)
);

OR2x6_ASAP7_75t_L g912 ( 
.A(n_897),
.B(n_144),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_895),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_913),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_L g915 ( 
.A(n_910),
.B(n_897),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_911),
.Y(n_916)
);

INVx2_ASAP7_75t_L g917 ( 
.A(n_912),
.Y(n_917)
);

INVx2_ASAP7_75t_L g918 ( 
.A(n_912),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_912),
.Y(n_919)
);

INVx2_ASAP7_75t_L g920 ( 
.A(n_914),
.Y(n_920)
);

INVx2_ASAP7_75t_L g921 ( 
.A(n_916),
.Y(n_921)
);

INVx2_ASAP7_75t_L g922 ( 
.A(n_915),
.Y(n_922)
);

OA22x2_ASAP7_75t_L g923 ( 
.A1(n_919),
.A2(n_900),
.B1(n_901),
.B2(n_904),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_917),
.Y(n_924)
);

AO22x2_ASAP7_75t_L g925 ( 
.A1(n_918),
.A2(n_909),
.B1(n_906),
.B2(n_907),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_920),
.Y(n_926)
);

INVx2_ASAP7_75t_SL g927 ( 
.A(n_924),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_921),
.Y(n_928)
);

AOI22x1_ASAP7_75t_L g929 ( 
.A1(n_925),
.A2(n_899),
.B1(n_908),
.B2(n_905),
.Y(n_929)
);

AOI22x1_ASAP7_75t_L g930 ( 
.A1(n_925),
.A2(n_905),
.B1(n_898),
.B2(n_896),
.Y(n_930)
);

INVx2_ASAP7_75t_L g931 ( 
.A(n_926),
.Y(n_931)
);

INVxp33_ASAP7_75t_L g932 ( 
.A(n_929),
.Y(n_932)
);

INVx1_ASAP7_75t_L g933 ( 
.A(n_928),
.Y(n_933)
);

AOI22x1_ASAP7_75t_L g934 ( 
.A1(n_932),
.A2(n_927),
.B1(n_922),
.B2(n_930),
.Y(n_934)
);

AOI31xp33_ASAP7_75t_L g935 ( 
.A1(n_932),
.A2(n_923),
.A3(n_161),
.B(n_165),
.Y(n_935)
);

INVx2_ASAP7_75t_L g936 ( 
.A(n_931),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_936),
.Y(n_937)
);

OAI22xp5_ASAP7_75t_L g938 ( 
.A1(n_935),
.A2(n_933),
.B1(n_931),
.B2(n_181),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_934),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_937),
.Y(n_940)
);

INVxp67_ASAP7_75t_SL g941 ( 
.A(n_939),
.Y(n_941)
);

INVx1_ASAP7_75t_L g942 ( 
.A(n_938),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_937),
.Y(n_943)
);

NOR2xp33_ASAP7_75t_L g944 ( 
.A(n_942),
.B(n_186),
.Y(n_944)
);

INVx1_ASAP7_75t_L g945 ( 
.A(n_941),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_940),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_943),
.Y(n_947)
);

NOR3xp33_ASAP7_75t_SL g948 ( 
.A(n_945),
.B(n_228),
.C(n_187),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_946),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_947),
.Y(n_950)
);

INVx2_ASAP7_75t_L g951 ( 
.A(n_944),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_949),
.Y(n_952)
);

INVx3_ASAP7_75t_L g953 ( 
.A(n_950),
.Y(n_953)
);

AND2x4_ASAP7_75t_L g954 ( 
.A(n_951),
.B(n_192),
.Y(n_954)
);

INVxp33_ASAP7_75t_SL g955 ( 
.A(n_952),
.Y(n_955)
);

INVx2_ASAP7_75t_SL g956 ( 
.A(n_953),
.Y(n_956)
);

AOI22xp33_ASAP7_75t_L g957 ( 
.A1(n_953),
.A2(n_948),
.B1(n_195),
.B2(n_196),
.Y(n_957)
);

INVx1_ASAP7_75t_L g958 ( 
.A(n_956),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_955),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_957),
.Y(n_960)
);

AOI22xp5_ASAP7_75t_L g961 ( 
.A1(n_958),
.A2(n_959),
.B1(n_960),
.B2(n_954),
.Y(n_961)
);

AOI22xp5_ASAP7_75t_L g962 ( 
.A1(n_958),
.A2(n_193),
.B1(n_198),
.B2(n_206),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_961),
.Y(n_963)
);

INVx1_ASAP7_75t_L g964 ( 
.A(n_962),
.Y(n_964)
);

INVx1_ASAP7_75t_L g965 ( 
.A(n_961),
.Y(n_965)
);

AOI22xp33_ASAP7_75t_SL g966 ( 
.A1(n_963),
.A2(n_209),
.B1(n_210),
.B2(n_211),
.Y(n_966)
);

OAI22xp5_ASAP7_75t_L g967 ( 
.A1(n_965),
.A2(n_212),
.B1(n_213),
.B2(n_214),
.Y(n_967)
);

INVxp67_ASAP7_75t_SL g968 ( 
.A(n_967),
.Y(n_968)
);

INVxp67_ASAP7_75t_R g969 ( 
.A(n_966),
.Y(n_969)
);

AOI221xp5_ASAP7_75t_L g970 ( 
.A1(n_968),
.A2(n_964),
.B1(n_218),
.B2(n_219),
.C(n_220),
.Y(n_970)
);

AOI211xp5_ASAP7_75t_L g971 ( 
.A1(n_970),
.A2(n_969),
.B(n_221),
.C(n_223),
.Y(n_971)
);


endmodule