module fake_netlist_6_1580_n_1887 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_166, n_28, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_127, n_125, n_153, n_168, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_165, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_171, n_31, n_57, n_169, n_53, n_51, n_44, n_56, n_1887);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_127;
input n_125;
input n_153;
input n_168;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_165;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_171;
input n_31;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1887;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_1853;
wire n_783;
wire n_1738;
wire n_798;
wire n_188;
wire n_1575;
wire n_1854;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1688;
wire n_1691;
wire n_1009;
wire n_1743;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_1844;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1803;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1867;
wire n_1704;
wire n_1078;
wire n_544;
wire n_250;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_616;
wire n_658;
wire n_1874;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1842;
wire n_1620;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_1815;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1644;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_1843;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1876;
wire n_1697;
wire n_243;
wire n_979;
wire n_1873;
wire n_905;
wire n_1866;
wire n_1680;
wire n_175;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1865;
wire n_1875;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_210;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_178;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1747;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1802;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_928;
wire n_835;
wire n_1214;
wire n_690;
wire n_850;
wire n_1801;
wire n_1886;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_1709;
wire n_1825;
wire n_1757;
wire n_1796;
wire n_1792;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_595;
wire n_297;
wire n_627;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1858;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_1839;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_1863;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_173;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_1788;
wire n_622;
wire n_1469;
wire n_1838;
wire n_1835;
wire n_1766;
wire n_1776;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_1878;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_1181;
wire n_1822;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_1817;
wire n_927;
wire n_1849;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_216;
wire n_912;
wire n_1857;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_527;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_1837;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_211;
wire n_1483;
wire n_1834;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_1877;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1769;
wire n_1220;
wire n_556;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1775;
wire n_1773;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_1745;
wire n_914;
wire n_759;
wire n_1831;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1881;
wire n_1267;
wire n_1281;
wire n_1806;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_177;
wire n_1855;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_1832;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_1869;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_1871;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_1859;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_198;
wire n_1847;
wire n_179;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1841;
wire n_1639;
wire n_1623;
wire n_183;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1818;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_1870;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_1828;
wire n_1695;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1883;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_1823;
wire n_227;
wire n_1720;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_1846;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_1676;
wire n_833;
wire n_1830;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_1758;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1559;
wire n_1725;
wire n_1872;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1741;
wire n_1325;
wire n_1002;
wire n_1746;
wire n_545;
wire n_489;
wire n_1804;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1860;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1800;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1882;
wire n_1118;
wire n_1076;
wire n_194;
wire n_1007;
wire n_1807;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_1879;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_181;
wire n_1810;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_1729;
wire n_669;
wire n_176;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1785;
wire n_763;
wire n_1147;
wire n_1848;
wire n_360;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_174;
wire n_1173;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_719;
wire n_228;
wire n_1525;
wire n_455;
wire n_1585;
wire n_1851;
wire n_363;
wire n_1799;
wire n_1090;
wire n_592;
wire n_1816;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_1829;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_404;
wire n_271;
wire n_1884;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1819;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_373;
wire n_1632;
wire n_1805;
wire n_257;
wire n_1557;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_1850;
wire n_1868;
wire n_207;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_1836;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1856;
wire n_1862;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1885;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

INVx1_ASAP7_75t_SL g173 ( 
.A(n_29),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_161),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_162),
.Y(n_175)
);

INVx1_ASAP7_75t_SL g176 ( 
.A(n_33),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_55),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_68),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_37),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_50),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_39),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_78),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_19),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_61),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_28),
.Y(n_185)
);

BUFx10_ASAP7_75t_L g186 ( 
.A(n_10),
.Y(n_186)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_15),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_137),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_72),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_95),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_134),
.Y(n_191)
);

INVxp67_ASAP7_75t_L g192 ( 
.A(n_22),
.Y(n_192)
);

BUFx3_ASAP7_75t_L g193 ( 
.A(n_0),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_125),
.Y(n_194)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_153),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_24),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_160),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_2),
.Y(n_198)
);

CKINVDCx16_ASAP7_75t_R g199 ( 
.A(n_126),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_140),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_105),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_86),
.Y(n_202)
);

INVxp67_ASAP7_75t_L g203 ( 
.A(n_0),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_138),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_152),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_13),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_71),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_46),
.Y(n_208)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_18),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_74),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_85),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_23),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_158),
.Y(n_213)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_164),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_120),
.Y(n_215)
);

BUFx6f_ASAP7_75t_L g216 ( 
.A(n_166),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_7),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_133),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_141),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_63),
.Y(n_220)
);

BUFx5_ASAP7_75t_L g221 ( 
.A(n_118),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_73),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_50),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_114),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_21),
.Y(n_225)
);

INVx1_ASAP7_75t_SL g226 ( 
.A(n_53),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_154),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_109),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_139),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_52),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_103),
.Y(n_231)
);

HB1xp67_ASAP7_75t_L g232 ( 
.A(n_112),
.Y(n_232)
);

BUFx5_ASAP7_75t_L g233 ( 
.A(n_35),
.Y(n_233)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_163),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_24),
.Y(n_235)
);

BUFx3_ASAP7_75t_L g236 ( 
.A(n_127),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_39),
.Y(n_237)
);

CKINVDCx16_ASAP7_75t_R g238 ( 
.A(n_30),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_148),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_36),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_145),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_165),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_89),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_9),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_16),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_108),
.Y(n_246)
);

INVx2_ASAP7_75t_SL g247 ( 
.A(n_128),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_37),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_30),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_83),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_171),
.Y(n_251)
);

BUFx6f_ASAP7_75t_L g252 ( 
.A(n_143),
.Y(n_252)
);

CKINVDCx16_ASAP7_75t_R g253 ( 
.A(n_9),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_75),
.Y(n_254)
);

CKINVDCx14_ASAP7_75t_R g255 ( 
.A(n_12),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_81),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_40),
.Y(n_257)
);

BUFx6f_ASAP7_75t_L g258 ( 
.A(n_80),
.Y(n_258)
);

BUFx2_ASAP7_75t_L g259 ( 
.A(n_41),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_14),
.Y(n_260)
);

INVx2_ASAP7_75t_SL g261 ( 
.A(n_111),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_60),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_64),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_48),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_28),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_167),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_117),
.Y(n_267)
);

INVx2_ASAP7_75t_SL g268 ( 
.A(n_6),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_54),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_146),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_48),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_168),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_98),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_2),
.Y(n_274)
);

CKINVDCx14_ASAP7_75t_R g275 ( 
.A(n_10),
.Y(n_275)
);

HB1xp67_ASAP7_75t_L g276 ( 
.A(n_1),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_151),
.Y(n_277)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_84),
.Y(n_278)
);

BUFx3_ASAP7_75t_L g279 ( 
.A(n_51),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_70),
.Y(n_280)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_102),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_129),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_123),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_21),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_79),
.Y(n_285)
);

BUFx2_ASAP7_75t_L g286 ( 
.A(n_35),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_5),
.Y(n_287)
);

INVxp67_ASAP7_75t_L g288 ( 
.A(n_155),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_27),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_76),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_1),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_62),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_23),
.Y(n_293)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_16),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_22),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_87),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_169),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_67),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_101),
.Y(n_299)
);

INVx2_ASAP7_75t_SL g300 ( 
.A(n_57),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_65),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_15),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_121),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_32),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_144),
.Y(n_305)
);

INVx1_ASAP7_75t_SL g306 ( 
.A(n_12),
.Y(n_306)
);

BUFx10_ASAP7_75t_L g307 ( 
.A(n_149),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_170),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_99),
.Y(n_309)
);

BUFx5_ASAP7_75t_L g310 ( 
.A(n_147),
.Y(n_310)
);

BUFx2_ASAP7_75t_SL g311 ( 
.A(n_31),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_4),
.Y(n_312)
);

BUFx3_ASAP7_75t_L g313 ( 
.A(n_49),
.Y(n_313)
);

INVx1_ASAP7_75t_SL g314 ( 
.A(n_93),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_36),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_90),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_25),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_34),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_172),
.Y(n_319)
);

INVx2_ASAP7_75t_L g320 ( 
.A(n_13),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_6),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_4),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_20),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_46),
.Y(n_324)
);

INVx3_ASAP7_75t_L g325 ( 
.A(n_96),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_19),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_130),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_26),
.Y(n_328)
);

BUFx2_ASAP7_75t_L g329 ( 
.A(n_7),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g330 ( 
.A(n_107),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_59),
.Y(n_331)
);

CKINVDCx14_ASAP7_75t_R g332 ( 
.A(n_88),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_32),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_8),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_5),
.Y(n_335)
);

INVx2_ASAP7_75t_SL g336 ( 
.A(n_113),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_31),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_56),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_100),
.Y(n_339)
);

BUFx3_ASAP7_75t_L g340 ( 
.A(n_18),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_26),
.Y(n_341)
);

BUFx10_ASAP7_75t_L g342 ( 
.A(n_20),
.Y(n_342)
);

INVx1_ASAP7_75t_SL g343 ( 
.A(n_157),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_94),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_233),
.Y(n_345)
);

INVxp67_ASAP7_75t_SL g346 ( 
.A(n_232),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g347 ( 
.A(n_174),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_255),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_233),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_233),
.Y(n_350)
);

INVxp67_ASAP7_75t_SL g351 ( 
.A(n_236),
.Y(n_351)
);

CKINVDCx14_ASAP7_75t_R g352 ( 
.A(n_275),
.Y(n_352)
);

INVxp67_ASAP7_75t_SL g353 ( 
.A(n_236),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_233),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_233),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_233),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_233),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_193),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_193),
.Y(n_359)
);

INVxp67_ASAP7_75t_L g360 ( 
.A(n_259),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_313),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_238),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_187),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_253),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_187),
.Y(n_365)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_174),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_179),
.Y(n_367)
);

BUFx6f_ASAP7_75t_L g368 ( 
.A(n_216),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_180),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_181),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_313),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_340),
.Y(n_372)
);

CKINVDCx20_ASAP7_75t_R g373 ( 
.A(n_184),
.Y(n_373)
);

INVxp67_ASAP7_75t_SL g374 ( 
.A(n_279),
.Y(n_374)
);

CKINVDCx20_ASAP7_75t_R g375 ( 
.A(n_184),
.Y(n_375)
);

INVx3_ASAP7_75t_L g376 ( 
.A(n_279),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_340),
.Y(n_377)
);

INVxp33_ASAP7_75t_SL g378 ( 
.A(n_276),
.Y(n_378)
);

INVxp67_ASAP7_75t_SL g379 ( 
.A(n_325),
.Y(n_379)
);

INVxp33_ASAP7_75t_SL g380 ( 
.A(n_196),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_183),
.Y(n_381)
);

HB1xp67_ASAP7_75t_L g382 ( 
.A(n_286),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_185),
.Y(n_383)
);

CKINVDCx20_ASAP7_75t_R g384 ( 
.A(n_219),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_237),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_206),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_260),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_208),
.Y(n_388)
);

INVxp67_ASAP7_75t_SL g389 ( 
.A(n_325),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_264),
.Y(n_390)
);

BUFx6f_ASAP7_75t_L g391 ( 
.A(n_216),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_287),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_289),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_295),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_304),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_312),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_315),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_323),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_212),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_223),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_225),
.Y(n_401)
);

CKINVDCx16_ASAP7_75t_R g402 ( 
.A(n_199),
.Y(n_402)
);

CKINVDCx16_ASAP7_75t_R g403 ( 
.A(n_332),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_333),
.Y(n_404)
);

INVxp33_ASAP7_75t_L g405 ( 
.A(n_329),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_235),
.Y(n_406)
);

CKINVDCx20_ASAP7_75t_R g407 ( 
.A(n_219),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_240),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_335),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_341),
.Y(n_410)
);

INVxp33_ASAP7_75t_SL g411 ( 
.A(n_196),
.Y(n_411)
);

BUFx2_ASAP7_75t_L g412 ( 
.A(n_198),
.Y(n_412)
);

HB1xp67_ASAP7_75t_L g413 ( 
.A(n_198),
.Y(n_413)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_221),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_175),
.Y(n_415)
);

CKINVDCx20_ASAP7_75t_R g416 ( 
.A(n_243),
.Y(n_416)
);

INVxp67_ASAP7_75t_SL g417 ( 
.A(n_325),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_245),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_249),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_178),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_257),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_182),
.Y(n_422)
);

CKINVDCx20_ASAP7_75t_R g423 ( 
.A(n_243),
.Y(n_423)
);

CKINVDCx20_ASAP7_75t_R g424 ( 
.A(n_254),
.Y(n_424)
);

CKINVDCx16_ASAP7_75t_R g425 ( 
.A(n_254),
.Y(n_425)
);

CKINVDCx20_ASAP7_75t_R g426 ( 
.A(n_263),
.Y(n_426)
);

CKINVDCx20_ASAP7_75t_R g427 ( 
.A(n_263),
.Y(n_427)
);

BUFx2_ASAP7_75t_SL g428 ( 
.A(n_299),
.Y(n_428)
);

CKINVDCx20_ASAP7_75t_R g429 ( 
.A(n_299),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_189),
.Y(n_430)
);

INVxp67_ASAP7_75t_L g431 ( 
.A(n_186),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_209),
.Y(n_432)
);

INVx2_ASAP7_75t_L g433 ( 
.A(n_355),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_355),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_376),
.B(n_379),
.Y(n_435)
);

OA21x2_ASAP7_75t_L g436 ( 
.A1(n_414),
.A2(n_294),
.B(n_209),
.Y(n_436)
);

INVx2_ASAP7_75t_L g437 ( 
.A(n_345),
.Y(n_437)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_349),
.Y(n_438)
);

AND2x4_ASAP7_75t_L g439 ( 
.A(n_389),
.B(n_247),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_350),
.Y(n_440)
);

OA21x2_ASAP7_75t_L g441 ( 
.A1(n_414),
.A2(n_320),
.B(n_294),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_354),
.Y(n_442)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_356),
.Y(n_443)
);

BUFx8_ASAP7_75t_L g444 ( 
.A(n_412),
.Y(n_444)
);

INVx4_ASAP7_75t_L g445 ( 
.A(n_368),
.Y(n_445)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_357),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_368),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_368),
.Y(n_448)
);

XNOR2xp5_ASAP7_75t_L g449 ( 
.A(n_347),
.B(n_217),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_368),
.Y(n_450)
);

INVx2_ASAP7_75t_L g451 ( 
.A(n_368),
.Y(n_451)
);

AND3x2_ASAP7_75t_L g452 ( 
.A(n_382),
.B(n_203),
.C(n_192),
.Y(n_452)
);

INVx2_ASAP7_75t_L g453 ( 
.A(n_391),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_391),
.Y(n_454)
);

BUFx6f_ASAP7_75t_L g455 ( 
.A(n_391),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_391),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_376),
.B(n_247),
.Y(n_457)
);

AND2x2_ASAP7_75t_L g458 ( 
.A(n_417),
.B(n_261),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_376),
.B(n_261),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_391),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_363),
.Y(n_461)
);

AND2x2_ASAP7_75t_L g462 ( 
.A(n_351),
.B(n_300),
.Y(n_462)
);

INVx2_ASAP7_75t_L g463 ( 
.A(n_363),
.Y(n_463)
);

INVx3_ASAP7_75t_L g464 ( 
.A(n_365),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_365),
.Y(n_465)
);

AND2x2_ASAP7_75t_L g466 ( 
.A(n_353),
.B(n_374),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_432),
.Y(n_467)
);

BUFx6f_ASAP7_75t_L g468 ( 
.A(n_432),
.Y(n_468)
);

INVx2_ASAP7_75t_L g469 ( 
.A(n_415),
.Y(n_469)
);

HB1xp67_ASAP7_75t_L g470 ( 
.A(n_413),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_381),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_420),
.B(n_300),
.Y(n_472)
);

BUFx6f_ASAP7_75t_L g473 ( 
.A(n_422),
.Y(n_473)
);

AND2x2_ASAP7_75t_L g474 ( 
.A(n_430),
.B(n_336),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_385),
.Y(n_475)
);

INVx2_ASAP7_75t_L g476 ( 
.A(n_387),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_390),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_392),
.Y(n_478)
);

XNOR2xp5_ASAP7_75t_L g479 ( 
.A(n_366),
.B(n_217),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_393),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_358),
.B(n_336),
.Y(n_481)
);

AND2x4_ASAP7_75t_L g482 ( 
.A(n_359),
.B(n_195),
.Y(n_482)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_394),
.Y(n_483)
);

CKINVDCx20_ASAP7_75t_R g484 ( 
.A(n_373),
.Y(n_484)
);

INVx2_ASAP7_75t_L g485 ( 
.A(n_395),
.Y(n_485)
);

BUFx6f_ASAP7_75t_L g486 ( 
.A(n_396),
.Y(n_486)
);

AND2x2_ASAP7_75t_L g487 ( 
.A(n_361),
.B(n_371),
.Y(n_487)
);

INVx2_ASAP7_75t_L g488 ( 
.A(n_397),
.Y(n_488)
);

INVx2_ASAP7_75t_L g489 ( 
.A(n_398),
.Y(n_489)
);

INVx4_ASAP7_75t_L g490 ( 
.A(n_367),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_404),
.Y(n_491)
);

BUFx6f_ASAP7_75t_L g492 ( 
.A(n_409),
.Y(n_492)
);

INVxp67_ASAP7_75t_L g493 ( 
.A(n_412),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_372),
.B(n_191),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_377),
.B(n_191),
.Y(n_495)
);

BUFx6f_ASAP7_75t_L g496 ( 
.A(n_410),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_346),
.B(n_197),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_367),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_369),
.Y(n_499)
);

INVx2_ASAP7_75t_L g500 ( 
.A(n_369),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_403),
.B(n_197),
.Y(n_501)
);

NOR2xp33_ASAP7_75t_L g502 ( 
.A(n_378),
.B(n_288),
.Y(n_502)
);

INVx2_ASAP7_75t_L g503 ( 
.A(n_360),
.Y(n_503)
);

CKINVDCx5p33_ASAP7_75t_R g504 ( 
.A(n_428),
.Y(n_504)
);

AOI22xp5_ASAP7_75t_L g505 ( 
.A1(n_378),
.A2(n_244),
.B1(n_293),
.B2(n_324),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_370),
.Y(n_506)
);

INVx2_ASAP7_75t_L g507 ( 
.A(n_370),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_383),
.Y(n_508)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_383),
.Y(n_509)
);

BUFx6f_ASAP7_75t_L g510 ( 
.A(n_386),
.Y(n_510)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_433),
.Y(n_511)
);

NOR2xp33_ASAP7_75t_L g512 ( 
.A(n_498),
.B(n_402),
.Y(n_512)
);

OAI21xp33_ASAP7_75t_SL g513 ( 
.A1(n_458),
.A2(n_268),
.B(n_320),
.Y(n_513)
);

INVx2_ASAP7_75t_L g514 ( 
.A(n_433),
.Y(n_514)
);

INVx3_ASAP7_75t_L g515 ( 
.A(n_455),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_436),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_436),
.Y(n_517)
);

INVxp67_ASAP7_75t_SL g518 ( 
.A(n_435),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_436),
.Y(n_519)
);

INVx2_ASAP7_75t_L g520 ( 
.A(n_433),
.Y(n_520)
);

NOR2xp33_ASAP7_75t_L g521 ( 
.A(n_498),
.B(n_348),
.Y(n_521)
);

INVx2_ASAP7_75t_SL g522 ( 
.A(n_466),
.Y(n_522)
);

INVx2_ASAP7_75t_L g523 ( 
.A(n_433),
.Y(n_523)
);

INVx3_ASAP7_75t_L g524 ( 
.A(n_455),
.Y(n_524)
);

INVx2_ASAP7_75t_L g525 ( 
.A(n_437),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_436),
.Y(n_526)
);

INVx2_ASAP7_75t_L g527 ( 
.A(n_437),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_435),
.B(n_352),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_439),
.B(n_348),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_436),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_L g531 ( 
.A(n_439),
.B(n_466),
.Y(n_531)
);

INVx2_ASAP7_75t_L g532 ( 
.A(n_437),
.Y(n_532)
);

BUFx3_ASAP7_75t_L g533 ( 
.A(n_487),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_441),
.Y(n_534)
);

INVxp33_ASAP7_75t_SL g535 ( 
.A(n_504),
.Y(n_535)
);

AOI22xp33_ASAP7_75t_L g536 ( 
.A1(n_439),
.A2(n_268),
.B1(n_405),
.B2(n_380),
.Y(n_536)
);

INVx2_ASAP7_75t_L g537 ( 
.A(n_438),
.Y(n_537)
);

INVx2_ASAP7_75t_L g538 ( 
.A(n_438),
.Y(n_538)
);

INVx2_ASAP7_75t_L g539 ( 
.A(n_438),
.Y(n_539)
);

BUFx10_ASAP7_75t_L g540 ( 
.A(n_502),
.Y(n_540)
);

BUFx3_ASAP7_75t_L g541 ( 
.A(n_487),
.Y(n_541)
);

INVx2_ASAP7_75t_L g542 ( 
.A(n_443),
.Y(n_542)
);

INVx2_ASAP7_75t_L g543 ( 
.A(n_443),
.Y(n_543)
);

INVx2_ASAP7_75t_L g544 ( 
.A(n_443),
.Y(n_544)
);

NAND3xp33_ASAP7_75t_L g545 ( 
.A(n_502),
.B(n_388),
.C(n_386),
.Y(n_545)
);

INVx3_ASAP7_75t_L g546 ( 
.A(n_455),
.Y(n_546)
);

AOI22xp33_ASAP7_75t_L g547 ( 
.A1(n_439),
.A2(n_411),
.B1(n_380),
.B2(n_311),
.Y(n_547)
);

INVxp67_ASAP7_75t_SL g548 ( 
.A(n_441),
.Y(n_548)
);

INVx2_ASAP7_75t_L g549 ( 
.A(n_446),
.Y(n_549)
);

INVx2_ASAP7_75t_L g550 ( 
.A(n_446),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_441),
.Y(n_551)
);

XNOR2xp5_ASAP7_75t_L g552 ( 
.A(n_505),
.B(n_375),
.Y(n_552)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_446),
.Y(n_553)
);

NAND3xp33_ASAP7_75t_L g554 ( 
.A(n_493),
.B(n_399),
.C(n_388),
.Y(n_554)
);

INVx2_ASAP7_75t_L g555 ( 
.A(n_468),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_441),
.Y(n_556)
);

INVx2_ASAP7_75t_SL g557 ( 
.A(n_466),
.Y(n_557)
);

CKINVDCx5p33_ASAP7_75t_R g558 ( 
.A(n_504),
.Y(n_558)
);

INVx2_ASAP7_75t_L g559 ( 
.A(n_468),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_441),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_434),
.Y(n_561)
);

NOR2xp33_ASAP7_75t_L g562 ( 
.A(n_499),
.B(n_411),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_468),
.Y(n_563)
);

BUFx6f_ASAP7_75t_L g564 ( 
.A(n_455),
.Y(n_564)
);

AOI22xp5_ASAP7_75t_L g565 ( 
.A1(n_493),
.A2(n_305),
.B1(n_330),
.B2(n_293),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_434),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_468),
.Y(n_567)
);

HB1xp67_ASAP7_75t_L g568 ( 
.A(n_470),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_440),
.Y(n_569)
);

INVx3_ASAP7_75t_L g570 ( 
.A(n_455),
.Y(n_570)
);

INVx2_ASAP7_75t_L g571 ( 
.A(n_468),
.Y(n_571)
);

BUFx10_ASAP7_75t_L g572 ( 
.A(n_510),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_442),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_L g574 ( 
.A(n_439),
.B(n_400),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_458),
.B(n_400),
.Y(n_575)
);

INVx4_ASAP7_75t_L g576 ( 
.A(n_473),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_SL g577 ( 
.A(n_510),
.B(n_401),
.Y(n_577)
);

BUFx6f_ASAP7_75t_L g578 ( 
.A(n_455),
.Y(n_578)
);

BUFx6f_ASAP7_75t_L g579 ( 
.A(n_455),
.Y(n_579)
);

OAI22xp33_ASAP7_75t_SL g580 ( 
.A1(n_497),
.A2(n_431),
.B1(n_195),
.B2(n_278),
.Y(n_580)
);

CKINVDCx6p67_ASAP7_75t_R g581 ( 
.A(n_490),
.Y(n_581)
);

BUFx6f_ASAP7_75t_L g582 ( 
.A(n_473),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_442),
.Y(n_583)
);

INVx3_ASAP7_75t_L g584 ( 
.A(n_445),
.Y(n_584)
);

INVx4_ASAP7_75t_L g585 ( 
.A(n_473),
.Y(n_585)
);

BUFx2_ASAP7_75t_L g586 ( 
.A(n_444),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_469),
.Y(n_587)
);

NOR3xp33_ASAP7_75t_L g588 ( 
.A(n_499),
.B(n_425),
.C(n_364),
.Y(n_588)
);

NOR2xp33_ASAP7_75t_L g589 ( 
.A(n_506),
.B(n_507),
.Y(n_589)
);

INVx3_ASAP7_75t_L g590 ( 
.A(n_445),
.Y(n_590)
);

BUFx6f_ASAP7_75t_L g591 ( 
.A(n_473),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_469),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_469),
.Y(n_593)
);

AO21x2_ASAP7_75t_L g594 ( 
.A1(n_457),
.A2(n_194),
.B(n_190),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_SL g595 ( 
.A(n_510),
.B(n_500),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_486),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_486),
.Y(n_597)
);

NOR2x1p5_ASAP7_75t_L g598 ( 
.A(n_490),
.B(n_362),
.Y(n_598)
);

BUFx2_ASAP7_75t_L g599 ( 
.A(n_444),
.Y(n_599)
);

INVx2_ASAP7_75t_L g600 ( 
.A(n_468),
.Y(n_600)
);

INVx2_ASAP7_75t_L g601 ( 
.A(n_468),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_464),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_486),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_486),
.Y(n_604)
);

NAND3xp33_ASAP7_75t_L g605 ( 
.A(n_503),
.B(n_406),
.C(n_401),
.Y(n_605)
);

NAND2xp33_ASAP7_75t_L g606 ( 
.A(n_500),
.B(n_406),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_486),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_486),
.Y(n_608)
);

NOR2xp33_ASAP7_75t_L g609 ( 
.A(n_506),
.B(n_408),
.Y(n_609)
);

INVx2_ASAP7_75t_L g610 ( 
.A(n_464),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_SL g611 ( 
.A(n_510),
.B(n_408),
.Y(n_611)
);

INVx2_ASAP7_75t_L g612 ( 
.A(n_464),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_486),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_492),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_492),
.Y(n_615)
);

BUFx3_ASAP7_75t_L g616 ( 
.A(n_487),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_L g617 ( 
.A(n_458),
.B(n_418),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_492),
.Y(n_618)
);

BUFx6f_ASAP7_75t_SL g619 ( 
.A(n_510),
.Y(n_619)
);

AND3x1_ASAP7_75t_L g620 ( 
.A(n_505),
.B(n_234),
.C(n_214),
.Y(n_620)
);

BUFx6f_ASAP7_75t_SL g621 ( 
.A(n_510),
.Y(n_621)
);

OAI22xp5_ASAP7_75t_L g622 ( 
.A1(n_500),
.A2(n_418),
.B1(n_419),
.B2(n_421),
.Y(n_622)
);

INVx3_ASAP7_75t_L g623 ( 
.A(n_445),
.Y(n_623)
);

INVx2_ASAP7_75t_L g624 ( 
.A(n_464),
.Y(n_624)
);

INVx2_ASAP7_75t_L g625 ( 
.A(n_464),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_492),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_492),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_492),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_492),
.Y(n_629)
);

AND2x4_ASAP7_75t_L g630 ( 
.A(n_482),
.B(n_214),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_496),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_496),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_L g633 ( 
.A(n_462),
.B(n_419),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_SL g634 ( 
.A(n_500),
.B(n_421),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_L g635 ( 
.A(n_462),
.B(n_226),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_L g636 ( 
.A(n_462),
.B(n_474),
.Y(n_636)
);

INVx2_ASAP7_75t_L g637 ( 
.A(n_463),
.Y(n_637)
);

BUFx6f_ASAP7_75t_L g638 ( 
.A(n_473),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_SL g639 ( 
.A(n_503),
.B(n_507),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_496),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_L g641 ( 
.A(n_474),
.B(n_314),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_496),
.Y(n_642)
);

INVx3_ASAP7_75t_L g643 ( 
.A(n_445),
.Y(n_643)
);

AND2x2_ASAP7_75t_L g644 ( 
.A(n_474),
.B(n_362),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_L g645 ( 
.A(n_497),
.B(n_343),
.Y(n_645)
);

BUFx10_ASAP7_75t_L g646 ( 
.A(n_470),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_496),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_496),
.Y(n_648)
);

INVx3_ASAP7_75t_L g649 ( 
.A(n_445),
.Y(n_649)
);

INVx2_ASAP7_75t_L g650 ( 
.A(n_463),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_496),
.Y(n_651)
);

BUFx10_ASAP7_75t_L g652 ( 
.A(n_452),
.Y(n_652)
);

INVx2_ASAP7_75t_L g653 ( 
.A(n_463),
.Y(n_653)
);

INVx6_ASAP7_75t_L g654 ( 
.A(n_473),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_476),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_476),
.Y(n_656)
);

BUFx3_ASAP7_75t_L g657 ( 
.A(n_471),
.Y(n_657)
);

INVx2_ASAP7_75t_L g658 ( 
.A(n_451),
.Y(n_658)
);

INVx2_ASAP7_75t_L g659 ( 
.A(n_451),
.Y(n_659)
);

INVx4_ASAP7_75t_L g660 ( 
.A(n_482),
.Y(n_660)
);

NOR2xp33_ASAP7_75t_L g661 ( 
.A(n_589),
.B(n_507),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_L g662 ( 
.A(n_518),
.B(n_508),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_SL g663 ( 
.A(n_522),
.B(n_508),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_548),
.B(n_508),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_657),
.Y(n_665)
);

AND2x2_ASAP7_75t_L g666 ( 
.A(n_522),
.B(n_503),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_L g667 ( 
.A(n_516),
.B(n_509),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_516),
.B(n_509),
.Y(n_668)
);

INVxp67_ASAP7_75t_L g669 ( 
.A(n_562),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_SL g670 ( 
.A(n_557),
.B(n_509),
.Y(n_670)
);

AND2x4_ASAP7_75t_L g671 ( 
.A(n_533),
.B(n_471),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_SL g672 ( 
.A(n_557),
.B(n_490),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_SL g673 ( 
.A(n_633),
.B(n_490),
.Y(n_673)
);

INVx2_ASAP7_75t_L g674 ( 
.A(n_511),
.Y(n_674)
);

AND2x4_ASAP7_75t_L g675 ( 
.A(n_533),
.B(n_541),
.Y(n_675)
);

INVx2_ASAP7_75t_L g676 ( 
.A(n_511),
.Y(n_676)
);

AND2x2_ASAP7_75t_L g677 ( 
.A(n_644),
.B(n_490),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_L g678 ( 
.A(n_517),
.B(n_519),
.Y(n_678)
);

AOI22xp5_ASAP7_75t_SL g679 ( 
.A1(n_552),
.A2(n_384),
.B1(n_407),
.B2(n_416),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_657),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_569),
.Y(n_681)
);

INVx3_ASAP7_75t_L g682 ( 
.A(n_660),
.Y(n_682)
);

NOR2xp67_ASAP7_75t_L g683 ( 
.A(n_545),
.B(n_501),
.Y(n_683)
);

AOI22xp5_ASAP7_75t_L g684 ( 
.A1(n_574),
.A2(n_501),
.B1(n_305),
.B2(n_330),
.Y(n_684)
);

NOR2xp67_ASAP7_75t_L g685 ( 
.A(n_554),
.B(n_494),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_SL g686 ( 
.A(n_575),
.B(n_444),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_531),
.B(n_457),
.Y(n_687)
);

NOR2xp33_ASAP7_75t_L g688 ( 
.A(n_609),
.B(n_364),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_L g689 ( 
.A(n_645),
.B(n_459),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_636),
.B(n_459),
.Y(n_690)
);

HB1xp67_ASAP7_75t_L g691 ( 
.A(n_568),
.Y(n_691)
);

INVx2_ASAP7_75t_L g692 ( 
.A(n_514),
.Y(n_692)
);

NOR2xp33_ASAP7_75t_SL g693 ( 
.A(n_586),
.B(n_428),
.Y(n_693)
);

INVx2_ASAP7_75t_L g694 ( 
.A(n_514),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_517),
.B(n_494),
.Y(n_695)
);

INVx2_ASAP7_75t_L g696 ( 
.A(n_520),
.Y(n_696)
);

A2O1A1Ixp33_ASAP7_75t_L g697 ( 
.A1(n_635),
.A2(n_495),
.B(n_234),
.C(n_278),
.Y(n_697)
);

INVx1_ASAP7_75t_SL g698 ( 
.A(n_646),
.Y(n_698)
);

INVx2_ASAP7_75t_L g699 ( 
.A(n_520),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_L g700 ( 
.A(n_561),
.B(n_495),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_519),
.B(n_482),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_L g702 ( 
.A(n_526),
.B(n_482),
.Y(n_702)
);

NOR2xp33_ASAP7_75t_L g703 ( 
.A(n_622),
.B(n_423),
.Y(n_703)
);

NAND2xp33_ASAP7_75t_SL g704 ( 
.A(n_598),
.B(n_244),
.Y(n_704)
);

NAND2x1_ASAP7_75t_L g705 ( 
.A(n_526),
.B(n_451),
.Y(n_705)
);

NAND2x1_ASAP7_75t_L g706 ( 
.A(n_530),
.B(n_453),
.Y(n_706)
);

NOR3xp33_ASAP7_75t_L g707 ( 
.A(n_605),
.B(n_481),
.C(n_472),
.Y(n_707)
);

INVx2_ASAP7_75t_L g708 ( 
.A(n_523),
.Y(n_708)
);

HB1xp67_ASAP7_75t_L g709 ( 
.A(n_644),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_L g710 ( 
.A(n_530),
.B(n_482),
.Y(n_710)
);

NOR3xp33_ASAP7_75t_L g711 ( 
.A(n_634),
.B(n_481),
.C(n_472),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_L g712 ( 
.A(n_561),
.B(n_447),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_L g713 ( 
.A(n_566),
.B(n_447),
.Y(n_713)
);

AOI22xp33_ASAP7_75t_L g714 ( 
.A1(n_630),
.A2(n_281),
.B1(n_273),
.B2(n_277),
.Y(n_714)
);

AND2x2_ASAP7_75t_L g715 ( 
.A(n_536),
.B(n_424),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_SL g716 ( 
.A(n_617),
.B(n_444),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_L g717 ( 
.A(n_566),
.B(n_448),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_L g718 ( 
.A(n_573),
.B(n_583),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_SL g719 ( 
.A(n_529),
.B(n_528),
.Y(n_719)
);

NOR2xp33_ASAP7_75t_L g720 ( 
.A(n_521),
.B(n_426),
.Y(n_720)
);

NAND2xp33_ASAP7_75t_L g721 ( 
.A(n_595),
.B(n_221),
.Y(n_721)
);

AOI21xp5_ASAP7_75t_L g722 ( 
.A1(n_639),
.A2(n_450),
.B(n_448),
.Y(n_722)
);

NOR2xp33_ASAP7_75t_L g723 ( 
.A(n_540),
.B(n_427),
.Y(n_723)
);

BUFx6f_ASAP7_75t_L g724 ( 
.A(n_541),
.Y(n_724)
);

AND2x6_ASAP7_75t_SL g725 ( 
.A(n_512),
.B(n_248),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_L g726 ( 
.A(n_573),
.B(n_450),
.Y(n_726)
);

INVx2_ASAP7_75t_L g727 ( 
.A(n_523),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_583),
.Y(n_728)
);

INVxp67_ASAP7_75t_L g729 ( 
.A(n_646),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_616),
.Y(n_730)
);

INVx2_ASAP7_75t_L g731 ( 
.A(n_525),
.Y(n_731)
);

INVxp67_ASAP7_75t_SL g732 ( 
.A(n_584),
.Y(n_732)
);

INVx1_ASAP7_75t_SL g733 ( 
.A(n_646),
.Y(n_733)
);

AND2x6_ASAP7_75t_L g734 ( 
.A(n_534),
.B(n_281),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_616),
.Y(n_735)
);

INVx2_ASAP7_75t_SL g736 ( 
.A(n_540),
.Y(n_736)
);

A2O1A1Ixp33_ASAP7_75t_L g737 ( 
.A1(n_513),
.A2(n_241),
.B(n_319),
.C(n_297),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_SL g738 ( 
.A(n_547),
.B(n_444),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_587),
.Y(n_739)
);

CKINVDCx5p33_ASAP7_75t_R g740 ( 
.A(n_558),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_SL g741 ( 
.A(n_540),
.B(n_177),
.Y(n_741)
);

INVx2_ASAP7_75t_L g742 ( 
.A(n_525),
.Y(n_742)
);

AOI22xp33_ASAP7_75t_L g743 ( 
.A1(n_630),
.A2(n_269),
.B1(n_227),
.B2(n_316),
.Y(n_743)
);

INVx2_ASAP7_75t_L g744 ( 
.A(n_527),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_L g745 ( 
.A(n_534),
.B(n_454),
.Y(n_745)
);

NOR2xp67_ASAP7_75t_L g746 ( 
.A(n_558),
.B(n_475),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_587),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_592),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_551),
.B(n_454),
.Y(n_749)
);

AND2x2_ASAP7_75t_L g750 ( 
.A(n_641),
.B(n_429),
.Y(n_750)
);

NOR2xp67_ASAP7_75t_SL g751 ( 
.A(n_551),
.B(n_216),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_L g752 ( 
.A(n_556),
.B(n_456),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_592),
.Y(n_753)
);

INVx2_ASAP7_75t_SL g754 ( 
.A(n_652),
.Y(n_754)
);

BUFx5_ASAP7_75t_L g755 ( 
.A(n_556),
.Y(n_755)
);

OAI22xp5_ASAP7_75t_L g756 ( 
.A1(n_620),
.A2(n_324),
.B1(n_248),
.B2(n_302),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_593),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_L g758 ( 
.A(n_560),
.B(n_456),
.Y(n_758)
);

INVx4_ASAP7_75t_L g759 ( 
.A(n_660),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_660),
.B(n_630),
.Y(n_760)
);

AOI22xp5_ASAP7_75t_L g761 ( 
.A1(n_606),
.A2(n_239),
.B1(n_200),
.B2(n_188),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_593),
.Y(n_762)
);

INVxp67_ASAP7_75t_L g763 ( 
.A(n_552),
.Y(n_763)
);

INVx2_ASAP7_75t_L g764 ( 
.A(n_527),
.Y(n_764)
);

NAND2xp33_ASAP7_75t_L g765 ( 
.A(n_598),
.B(n_221),
.Y(n_765)
);

AOI22xp5_ASAP7_75t_L g766 ( 
.A1(n_577),
.A2(n_611),
.B1(n_581),
.B2(n_588),
.Y(n_766)
);

BUFx6f_ASAP7_75t_L g767 ( 
.A(n_630),
.Y(n_767)
);

AO22x2_ASAP7_75t_L g768 ( 
.A1(n_565),
.A2(n_173),
.B1(n_176),
.B2(n_306),
.Y(n_768)
);

INVx2_ASAP7_75t_SL g769 ( 
.A(n_652),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_SL g770 ( 
.A(n_580),
.B(n_201),
.Y(n_770)
);

NOR2x1p5_ASAP7_75t_L g771 ( 
.A(n_581),
.B(n_318),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_655),
.Y(n_772)
);

INVx2_ASAP7_75t_L g773 ( 
.A(n_532),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_656),
.Y(n_774)
);

NOR2xp33_ASAP7_75t_L g775 ( 
.A(n_535),
.B(n_580),
.Y(n_775)
);

INVx2_ASAP7_75t_SL g776 ( 
.A(n_652),
.Y(n_776)
);

AOI22xp33_ASAP7_75t_L g777 ( 
.A1(n_594),
.A2(n_210),
.B1(n_338),
.B2(n_344),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_SL g778 ( 
.A(n_572),
.B(n_202),
.Y(n_778)
);

BUFx6f_ASAP7_75t_L g779 ( 
.A(n_602),
.Y(n_779)
);

OAI22xp33_ASAP7_75t_L g780 ( 
.A1(n_565),
.A2(n_242),
.B1(n_283),
.B2(n_290),
.Y(n_780)
);

INVx2_ASAP7_75t_L g781 ( 
.A(n_532),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_SL g782 ( 
.A(n_572),
.B(n_204),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_L g783 ( 
.A(n_610),
.B(n_460),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_610),
.B(n_460),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_612),
.B(n_624),
.Y(n_785)
);

INVx2_ASAP7_75t_L g786 ( 
.A(n_537),
.Y(n_786)
);

NOR2xp33_ASAP7_75t_L g787 ( 
.A(n_535),
.B(n_449),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_L g788 ( 
.A(n_584),
.B(n_453),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_SL g789 ( 
.A(n_572),
.B(n_205),
.Y(n_789)
);

INVx2_ASAP7_75t_SL g790 ( 
.A(n_594),
.Y(n_790)
);

INVx5_ASAP7_75t_L g791 ( 
.A(n_564),
.Y(n_791)
);

O2A1O1Ixp33_ASAP7_75t_L g792 ( 
.A1(n_513),
.A2(n_491),
.B(n_475),
.C(n_477),
.Y(n_792)
);

NOR2xp33_ASAP7_75t_L g793 ( 
.A(n_584),
.B(n_449),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_SL g794 ( 
.A(n_586),
.B(n_207),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_L g795 ( 
.A(n_590),
.B(n_453),
.Y(n_795)
);

NOR2xp33_ASAP7_75t_L g796 ( 
.A(n_590),
.B(n_449),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_656),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_SL g798 ( 
.A(n_599),
.B(n_211),
.Y(n_798)
);

AOI21xp5_ASAP7_75t_L g799 ( 
.A1(n_590),
.A2(n_476),
.B(n_489),
.Y(n_799)
);

NOR2xp33_ASAP7_75t_L g800 ( 
.A(n_623),
.B(n_479),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_612),
.Y(n_801)
);

NAND3xp33_ASAP7_75t_L g802 ( 
.A(n_599),
.B(n_452),
.C(n_480),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_SL g803 ( 
.A(n_623),
.B(n_213),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_SL g804 ( 
.A(n_623),
.B(n_215),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_L g805 ( 
.A(n_625),
.B(n_483),
.Y(n_805)
);

OR2x2_ASAP7_75t_L g806 ( 
.A(n_594),
.B(n_479),
.Y(n_806)
);

BUFx6f_ASAP7_75t_L g807 ( 
.A(n_625),
.Y(n_807)
);

BUFx5_ASAP7_75t_L g808 ( 
.A(n_596),
.Y(n_808)
);

OR2x2_ASAP7_75t_L g809 ( 
.A(n_658),
.B(n_479),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_SL g810 ( 
.A(n_643),
.B(n_649),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_L g811 ( 
.A(n_537),
.B(n_483),
.Y(n_811)
);

NAND2xp33_ASAP7_75t_L g812 ( 
.A(n_582),
.B(n_221),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_SL g813 ( 
.A(n_643),
.B(n_218),
.Y(n_813)
);

NOR2xp33_ASAP7_75t_L g814 ( 
.A(n_643),
.B(n_484),
.Y(n_814)
);

NOR3xp33_ASAP7_75t_L g815 ( 
.A(n_649),
.B(n_477),
.C(n_478),
.Y(n_815)
);

INVx2_ASAP7_75t_L g816 ( 
.A(n_538),
.Y(n_816)
);

NOR2xp33_ASAP7_75t_L g817 ( 
.A(n_649),
.B(n_484),
.Y(n_817)
);

OR2x6_ASAP7_75t_L g818 ( 
.A(n_637),
.B(n_478),
.Y(n_818)
);

NOR2xp67_ASAP7_75t_SL g819 ( 
.A(n_619),
.B(n_216),
.Y(n_819)
);

BUFx6f_ASAP7_75t_L g820 ( 
.A(n_564),
.Y(n_820)
);

AND2x6_ASAP7_75t_SL g821 ( 
.A(n_596),
.B(n_302),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_SL g822 ( 
.A(n_582),
.B(n_220),
.Y(n_822)
);

INVx2_ASAP7_75t_L g823 ( 
.A(n_538),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_L g824 ( 
.A(n_539),
.B(n_483),
.Y(n_824)
);

A2O1A1Ixp33_ASAP7_75t_L g825 ( 
.A1(n_539),
.A2(n_296),
.B(n_339),
.C(n_491),
.Y(n_825)
);

BUFx6f_ASAP7_75t_L g826 ( 
.A(n_767),
.Y(n_826)
);

BUFx6f_ASAP7_75t_L g827 ( 
.A(n_767),
.Y(n_827)
);

INVx5_ASAP7_75t_L g828 ( 
.A(n_734),
.Y(n_828)
);

INVx2_ASAP7_75t_L g829 ( 
.A(n_675),
.Y(n_829)
);

CKINVDCx5p33_ASAP7_75t_R g830 ( 
.A(n_740),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_675),
.Y(n_831)
);

INVx2_ASAP7_75t_SL g832 ( 
.A(n_691),
.Y(n_832)
);

CKINVDCx5p33_ASAP7_75t_R g833 ( 
.A(n_679),
.Y(n_833)
);

AOI22xp33_ASAP7_75t_L g834 ( 
.A1(n_690),
.A2(n_687),
.B1(n_689),
.B2(n_707),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_SL g835 ( 
.A(n_724),
.B(n_582),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_SL g836 ( 
.A(n_724),
.B(n_582),
.Y(n_836)
);

INVx2_ASAP7_75t_L g837 ( 
.A(n_801),
.Y(n_837)
);

AOI22xp5_ASAP7_75t_L g838 ( 
.A1(n_677),
.A2(n_619),
.B1(n_621),
.B2(n_628),
.Y(n_838)
);

NOR2xp33_ASAP7_75t_L g839 ( 
.A(n_669),
.B(n_688),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_L g840 ( 
.A(n_661),
.B(n_542),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_SL g841 ( 
.A(n_724),
.B(n_582),
.Y(n_841)
);

OAI22xp5_ASAP7_75t_L g842 ( 
.A1(n_678),
.A2(n_321),
.B1(n_621),
.B2(n_619),
.Y(n_842)
);

BUFx3_ASAP7_75t_L g843 ( 
.A(n_754),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_L g844 ( 
.A(n_755),
.B(n_542),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_L g845 ( 
.A(n_755),
.B(n_543),
.Y(n_845)
);

INVx2_ASAP7_75t_SL g846 ( 
.A(n_809),
.Y(n_846)
);

NOR3xp33_ASAP7_75t_SL g847 ( 
.A(n_780),
.B(n_322),
.C(n_318),
.Y(n_847)
);

HB1xp67_ASAP7_75t_L g848 ( 
.A(n_709),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_730),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_755),
.B(n_543),
.Y(n_850)
);

INVx2_ASAP7_75t_SL g851 ( 
.A(n_666),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_L g852 ( 
.A(n_755),
.B(n_544),
.Y(n_852)
);

OR2x4_ASAP7_75t_L g853 ( 
.A(n_775),
.B(n_480),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_755),
.B(n_544),
.Y(n_854)
);

BUFx3_ASAP7_75t_L g855 ( 
.A(n_769),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_SL g856 ( 
.A(n_746),
.B(n_591),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_735),
.Y(n_857)
);

NOR2xp33_ASAP7_75t_L g858 ( 
.A(n_793),
.B(n_621),
.Y(n_858)
);

AOI22xp5_ASAP7_75t_L g859 ( 
.A1(n_719),
.A2(n_608),
.B1(n_607),
.B2(n_597),
.Y(n_859)
);

OAI22xp33_ASAP7_75t_L g860 ( 
.A1(n_684),
.A2(n_321),
.B1(n_489),
.B2(n_488),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_739),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_747),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_748),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_753),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_757),
.Y(n_865)
);

NAND2x1p5_ASAP7_75t_L g866 ( 
.A(n_759),
.B(n_576),
.Y(n_866)
);

AOI22xp33_ASAP7_75t_L g867 ( 
.A1(n_664),
.A2(n_550),
.B1(n_553),
.B2(n_549),
.Y(n_867)
);

AOI22xp5_ASAP7_75t_L g868 ( 
.A1(n_685),
.A2(n_614),
.B1(n_613),
.B2(n_597),
.Y(n_868)
);

NAND2x1p5_ASAP7_75t_L g869 ( 
.A(n_759),
.B(n_576),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_762),
.Y(n_870)
);

INVx2_ASAP7_75t_L g871 ( 
.A(n_731),
.Y(n_871)
);

AND2x6_ASAP7_75t_L g872 ( 
.A(n_678),
.B(n_555),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_755),
.B(n_549),
.Y(n_873)
);

OAI22xp5_ASAP7_75t_SL g874 ( 
.A1(n_763),
.A2(n_322),
.B1(n_274),
.B2(n_271),
.Y(n_874)
);

OAI22xp5_ASAP7_75t_SL g875 ( 
.A1(n_787),
.A2(n_291),
.B1(n_265),
.B2(n_284),
.Y(n_875)
);

INVx2_ASAP7_75t_L g876 ( 
.A(n_742),
.Y(n_876)
);

OR2x6_ASAP7_75t_L g877 ( 
.A(n_776),
.B(n_485),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_772),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_662),
.B(n_550),
.Y(n_879)
);

OAI22xp5_ASAP7_75t_L g880 ( 
.A1(n_667),
.A2(n_317),
.B1(n_337),
.B2(n_326),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_L g881 ( 
.A(n_662),
.B(n_695),
.Y(n_881)
);

NAND3xp33_ASAP7_75t_SL g882 ( 
.A(n_720),
.B(n_334),
.C(n_328),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_774),
.Y(n_883)
);

BUFx4f_ASAP7_75t_L g884 ( 
.A(n_736),
.Y(n_884)
);

INVx2_ASAP7_75t_L g885 ( 
.A(n_744),
.Y(n_885)
);

INVx2_ASAP7_75t_L g886 ( 
.A(n_764),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_L g887 ( 
.A(n_695),
.B(n_553),
.Y(n_887)
);

INVx3_ASAP7_75t_L g888 ( 
.A(n_767),
.Y(n_888)
);

OAI22xp5_ASAP7_75t_L g889 ( 
.A1(n_667),
.A2(n_461),
.B1(n_467),
.B2(n_465),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_797),
.Y(n_890)
);

NAND3xp33_ASAP7_75t_SL g891 ( 
.A(n_703),
.B(n_280),
.C(n_285),
.Y(n_891)
);

INVx6_ASAP7_75t_L g892 ( 
.A(n_671),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_671),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_SL g894 ( 
.A(n_683),
.B(n_591),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_L g895 ( 
.A(n_668),
.B(n_637),
.Y(n_895)
);

AND2x2_ASAP7_75t_L g896 ( 
.A(n_750),
.B(n_485),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_L g897 ( 
.A(n_668),
.B(n_650),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_681),
.Y(n_898)
);

AO22x1_ASAP7_75t_L g899 ( 
.A1(n_796),
.A2(n_270),
.B1(n_251),
.B2(n_250),
.Y(n_899)
);

AOI22xp33_ASAP7_75t_L g900 ( 
.A1(n_664),
.A2(n_650),
.B1(n_653),
.B2(n_603),
.Y(n_900)
);

CKINVDCx5p33_ASAP7_75t_R g901 ( 
.A(n_723),
.Y(n_901)
);

NOR2xp33_ASAP7_75t_L g902 ( 
.A(n_800),
.B(n_603),
.Y(n_902)
);

INVx2_ASAP7_75t_SL g903 ( 
.A(n_698),
.Y(n_903)
);

INVx3_ASAP7_75t_L g904 ( 
.A(n_779),
.Y(n_904)
);

INVx2_ASAP7_75t_L g905 ( 
.A(n_773),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_L g906 ( 
.A(n_700),
.B(n_653),
.Y(n_906)
);

INVx2_ASAP7_75t_SL g907 ( 
.A(n_733),
.Y(n_907)
);

INVx2_ASAP7_75t_L g908 ( 
.A(n_781),
.Y(n_908)
);

INVx5_ASAP7_75t_L g909 ( 
.A(n_734),
.Y(n_909)
);

BUFx3_ASAP7_75t_L g910 ( 
.A(n_665),
.Y(n_910)
);

INVxp67_ASAP7_75t_L g911 ( 
.A(n_715),
.Y(n_911)
);

INVx5_ASAP7_75t_L g912 ( 
.A(n_734),
.Y(n_912)
);

INVx4_ASAP7_75t_L g913 ( 
.A(n_820),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_L g914 ( 
.A(n_732),
.B(n_604),
.Y(n_914)
);

BUFx4f_ASAP7_75t_L g915 ( 
.A(n_806),
.Y(n_915)
);

AND2x6_ASAP7_75t_SL g916 ( 
.A(n_814),
.B(n_461),
.Y(n_916)
);

INVxp67_ASAP7_75t_L g917 ( 
.A(n_817),
.Y(n_917)
);

BUFx4f_ASAP7_75t_L g918 ( 
.A(n_680),
.Y(n_918)
);

BUFx6f_ASAP7_75t_L g919 ( 
.A(n_820),
.Y(n_919)
);

AOI22xp33_ASAP7_75t_L g920 ( 
.A1(n_790),
.A2(n_627),
.B1(n_608),
.B2(n_651),
.Y(n_920)
);

INVx2_ASAP7_75t_SL g921 ( 
.A(n_771),
.Y(n_921)
);

O2A1O1Ixp33_ASAP7_75t_L g922 ( 
.A1(n_663),
.A2(n_489),
.B(n_488),
.C(n_485),
.Y(n_922)
);

INVx2_ASAP7_75t_SL g923 ( 
.A(n_670),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_728),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_805),
.Y(n_925)
);

INVx1_ASAP7_75t_SL g926 ( 
.A(n_756),
.Y(n_926)
);

BUFx2_ASAP7_75t_L g927 ( 
.A(n_704),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_L g928 ( 
.A(n_718),
.B(n_701),
.Y(n_928)
);

AND2x2_ASAP7_75t_L g929 ( 
.A(n_729),
.B(n_488),
.Y(n_929)
);

NOR2xp33_ASAP7_75t_L g930 ( 
.A(n_741),
.B(n_613),
.Y(n_930)
);

BUFx12f_ASAP7_75t_L g931 ( 
.A(n_821),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_805),
.Y(n_932)
);

INVx1_ASAP7_75t_L g933 ( 
.A(n_818),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_L g934 ( 
.A(n_701),
.B(n_614),
.Y(n_934)
);

INVx2_ASAP7_75t_L g935 ( 
.A(n_786),
.Y(n_935)
);

AOI22xp5_ASAP7_75t_L g936 ( 
.A1(n_711),
.A2(n_618),
.B1(n_615),
.B2(n_651),
.Y(n_936)
);

OR2x6_ASAP7_75t_L g937 ( 
.A(n_738),
.B(n_252),
.Y(n_937)
);

AOI22xp33_ASAP7_75t_L g938 ( 
.A1(n_777),
.A2(n_815),
.B1(n_770),
.B2(n_710),
.Y(n_938)
);

BUFx3_ASAP7_75t_L g939 ( 
.A(n_818),
.Y(n_939)
);

OR2x6_ASAP7_75t_L g940 ( 
.A(n_686),
.B(n_716),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_L g941 ( 
.A(n_702),
.B(n_615),
.Y(n_941)
);

INVx2_ASAP7_75t_L g942 ( 
.A(n_816),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_818),
.Y(n_943)
);

CKINVDCx20_ASAP7_75t_R g944 ( 
.A(n_756),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_L g945 ( 
.A(n_682),
.B(n_515),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_785),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_785),
.Y(n_947)
);

HB1xp67_ASAP7_75t_L g948 ( 
.A(n_802),
.Y(n_948)
);

CKINVDCx11_ASAP7_75t_R g949 ( 
.A(n_725),
.Y(n_949)
);

AOI22xp5_ASAP7_75t_L g950 ( 
.A1(n_673),
.A2(n_618),
.B1(n_626),
.B2(n_648),
.Y(n_950)
);

NOR2xp33_ASAP7_75t_L g951 ( 
.A(n_693),
.B(n_626),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_L g952 ( 
.A(n_702),
.B(n_627),
.Y(n_952)
);

INVx1_ASAP7_75t_L g953 ( 
.A(n_811),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_L g954 ( 
.A(n_710),
.B(n_628),
.Y(n_954)
);

BUFx3_ASAP7_75t_L g955 ( 
.A(n_766),
.Y(n_955)
);

BUFx6f_ASAP7_75t_L g956 ( 
.A(n_820),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_811),
.Y(n_957)
);

HB1xp67_ASAP7_75t_L g958 ( 
.A(n_737),
.Y(n_958)
);

INVx5_ASAP7_75t_L g959 ( 
.A(n_734),
.Y(n_959)
);

BUFx2_ASAP7_75t_L g960 ( 
.A(n_768),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_SL g961 ( 
.A(n_682),
.B(n_591),
.Y(n_961)
);

CKINVDCx5p33_ASAP7_75t_R g962 ( 
.A(n_761),
.Y(n_962)
);

NOR2xp33_ASAP7_75t_L g963 ( 
.A(n_672),
.B(n_629),
.Y(n_963)
);

INVx1_ASAP7_75t_L g964 ( 
.A(n_824),
.Y(n_964)
);

AOI22xp33_ASAP7_75t_L g965 ( 
.A1(n_765),
.A2(n_631),
.B1(n_629),
.B2(n_648),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_824),
.Y(n_966)
);

INVx3_ASAP7_75t_L g967 ( 
.A(n_779),
.Y(n_967)
);

NOR2xp67_ASAP7_75t_L g968 ( 
.A(n_794),
.B(n_631),
.Y(n_968)
);

INVx2_ASAP7_75t_L g969 ( 
.A(n_823),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_L g970 ( 
.A(n_745),
.B(n_632),
.Y(n_970)
);

INVx2_ASAP7_75t_L g971 ( 
.A(n_674),
.Y(n_971)
);

AND2x2_ASAP7_75t_L g972 ( 
.A(n_768),
.B(n_186),
.Y(n_972)
);

INVx1_ASAP7_75t_L g973 ( 
.A(n_726),
.Y(n_973)
);

AOI22xp33_ASAP7_75t_L g974 ( 
.A1(n_714),
.A2(n_640),
.B1(n_632),
.B2(n_647),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_L g975 ( 
.A(n_745),
.B(n_640),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_L g976 ( 
.A(n_749),
.B(n_642),
.Y(n_976)
);

CKINVDCx20_ASAP7_75t_R g977 ( 
.A(n_798),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_L g978 ( 
.A(n_749),
.B(n_642),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_712),
.Y(n_979)
);

INVx2_ASAP7_75t_L g980 ( 
.A(n_676),
.Y(n_980)
);

INVx2_ASAP7_75t_L g981 ( 
.A(n_692),
.Y(n_981)
);

INVx2_ASAP7_75t_SL g982 ( 
.A(n_768),
.Y(n_982)
);

INVx2_ASAP7_75t_L g983 ( 
.A(n_694),
.Y(n_983)
);

INVxp67_ASAP7_75t_L g984 ( 
.A(n_721),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_L g985 ( 
.A(n_752),
.B(n_647),
.Y(n_985)
);

AND2x6_ASAP7_75t_SL g986 ( 
.A(n_713),
.B(n_465),
.Y(n_986)
);

NOR2xp33_ASAP7_75t_L g987 ( 
.A(n_810),
.B(n_515),
.Y(n_987)
);

NAND2x1p5_ASAP7_75t_L g988 ( 
.A(n_791),
.B(n_576),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_L g989 ( 
.A(n_752),
.B(n_515),
.Y(n_989)
);

AND2x4_ASAP7_75t_L g990 ( 
.A(n_760),
.B(n_467),
.Y(n_990)
);

BUFx2_ASAP7_75t_L g991 ( 
.A(n_697),
.Y(n_991)
);

INVx1_ASAP7_75t_L g992 ( 
.A(n_717),
.Y(n_992)
);

BUFx3_ASAP7_75t_L g993 ( 
.A(n_807),
.Y(n_993)
);

NOR2xp33_ASAP7_75t_L g994 ( 
.A(n_803),
.B(n_524),
.Y(n_994)
);

INVxp33_ASAP7_75t_L g995 ( 
.A(n_792),
.Y(n_995)
);

OR2x2_ASAP7_75t_SL g996 ( 
.A(n_807),
.B(n_186),
.Y(n_996)
);

BUFx6f_ASAP7_75t_L g997 ( 
.A(n_807),
.Y(n_997)
);

A2O1A1Ixp33_ASAP7_75t_L g998 ( 
.A1(n_799),
.A2(n_659),
.B(n_601),
.C(n_600),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_L g999 ( 
.A(n_758),
.B(n_524),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_L g1000 ( 
.A(n_758),
.B(n_524),
.Y(n_1000)
);

NOR2xp67_ASAP7_75t_L g1001 ( 
.A(n_722),
.B(n_659),
.Y(n_1001)
);

INVxp67_ASAP7_75t_L g1002 ( 
.A(n_783),
.Y(n_1002)
);

NAND2xp33_ASAP7_75t_L g1003 ( 
.A(n_808),
.B(n_221),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_L g1004 ( 
.A(n_808),
.B(n_696),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_SL g1005 ( 
.A(n_791),
.B(n_591),
.Y(n_1005)
);

INVx3_ASAP7_75t_L g1006 ( 
.A(n_705),
.Y(n_1006)
);

NOR2xp33_ASAP7_75t_L g1007 ( 
.A(n_804),
.B(n_546),
.Y(n_1007)
);

HB1xp67_ASAP7_75t_L g1008 ( 
.A(n_783),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_784),
.Y(n_1009)
);

INVx4_ASAP7_75t_L g1010 ( 
.A(n_826),
.Y(n_1010)
);

BUFx6f_ASAP7_75t_L g1011 ( 
.A(n_919),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_L g1012 ( 
.A(n_881),
.B(n_808),
.Y(n_1012)
);

AOI22xp33_ASAP7_75t_L g1013 ( 
.A1(n_955),
.A2(n_743),
.B1(n_813),
.B2(n_822),
.Y(n_1013)
);

AOI21xp5_ASAP7_75t_L g1014 ( 
.A1(n_928),
.A2(n_791),
.B(n_788),
.Y(n_1014)
);

INVx3_ASAP7_75t_L g1015 ( 
.A(n_997),
.Y(n_1015)
);

AOI21xp5_ASAP7_75t_L g1016 ( 
.A1(n_928),
.A2(n_791),
.B(n_795),
.Y(n_1016)
);

NOR2xp33_ASAP7_75t_L g1017 ( 
.A(n_839),
.B(n_778),
.Y(n_1017)
);

OAI21xp33_ASAP7_75t_L g1018 ( 
.A1(n_926),
.A2(n_784),
.B(n_825),
.Y(n_1018)
);

INVx2_ASAP7_75t_L g1019 ( 
.A(n_837),
.Y(n_1019)
);

NOR2xp33_ASAP7_75t_L g1020 ( 
.A(n_917),
.B(n_911),
.Y(n_1020)
);

AOI21xp33_ASAP7_75t_L g1021 ( 
.A1(n_995),
.A2(n_789),
.B(n_782),
.Y(n_1021)
);

NAND2xp5_ASAP7_75t_L g1022 ( 
.A(n_834),
.B(n_808),
.Y(n_1022)
);

OAI22xp5_ASAP7_75t_L g1023 ( 
.A1(n_881),
.A2(n_706),
.B1(n_699),
.B2(n_727),
.Y(n_1023)
);

AND2x2_ASAP7_75t_L g1024 ( 
.A(n_915),
.B(n_342),
.Y(n_1024)
);

INVx1_ASAP7_75t_L g1025 ( 
.A(n_898),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_L g1026 ( 
.A(n_946),
.B(n_808),
.Y(n_1026)
);

BUFx2_ASAP7_75t_L g1027 ( 
.A(n_832),
.Y(n_1027)
);

A2O1A1Ixp33_ASAP7_75t_L g1028 ( 
.A1(n_902),
.A2(n_708),
.B(n_751),
.C(n_812),
.Y(n_1028)
);

NAND2xp5_ASAP7_75t_L g1029 ( 
.A(n_947),
.B(n_808),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_L g1030 ( 
.A(n_1002),
.B(n_546),
.Y(n_1030)
);

AND2x2_ASAP7_75t_L g1031 ( 
.A(n_915),
.B(n_342),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_L g1032 ( 
.A(n_1008),
.B(n_546),
.Y(n_1032)
);

BUFx3_ASAP7_75t_L g1033 ( 
.A(n_830),
.Y(n_1033)
);

O2A1O1Ixp5_ASAP7_75t_L g1034 ( 
.A1(n_858),
.A2(n_819),
.B(n_585),
.C(n_571),
.Y(n_1034)
);

BUFx2_ASAP7_75t_L g1035 ( 
.A(n_853),
.Y(n_1035)
);

NAND2xp5_ASAP7_75t_L g1036 ( 
.A(n_973),
.B(n_570),
.Y(n_1036)
);

OAI22xp5_ASAP7_75t_L g1037 ( 
.A1(n_1009),
.A2(n_853),
.B1(n_906),
.B2(n_887),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_L g1038 ( 
.A(n_979),
.B(n_992),
.Y(n_1038)
);

O2A1O1Ixp33_ASAP7_75t_L g1039 ( 
.A1(n_860),
.A2(n_882),
.B(n_948),
.C(n_842),
.Y(n_1039)
);

NAND2xp5_ASAP7_75t_L g1040 ( 
.A(n_851),
.B(n_570),
.Y(n_1040)
);

INVx3_ASAP7_75t_L g1041 ( 
.A(n_997),
.Y(n_1041)
);

NOR2xp33_ASAP7_75t_L g1042 ( 
.A(n_901),
.B(n_570),
.Y(n_1042)
);

HB1xp67_ASAP7_75t_L g1043 ( 
.A(n_848),
.Y(n_1043)
);

A2O1A1Ixp33_ASAP7_75t_L g1044 ( 
.A1(n_930),
.A2(n_938),
.B(n_958),
.C(n_923),
.Y(n_1044)
);

AND2x2_ASAP7_75t_L g1045 ( 
.A(n_896),
.B(n_342),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_L g1046 ( 
.A(n_925),
.B(n_555),
.Y(n_1046)
);

AOI21x1_ASAP7_75t_L g1047 ( 
.A1(n_879),
.A2(n_559),
.B(n_563),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_L g1048 ( 
.A(n_932),
.B(n_559),
.Y(n_1048)
);

NAND2xp5_ASAP7_75t_L g1049 ( 
.A(n_953),
.B(n_957),
.Y(n_1049)
);

NAND2xp5_ASAP7_75t_L g1050 ( 
.A(n_964),
.B(n_563),
.Y(n_1050)
);

HB1xp67_ASAP7_75t_L g1051 ( 
.A(n_846),
.Y(n_1051)
);

NAND2xp5_ASAP7_75t_SL g1052 ( 
.A(n_918),
.B(n_222),
.Y(n_1052)
);

AND2x4_ASAP7_75t_L g1053 ( 
.A(n_829),
.B(n_567),
.Y(n_1053)
);

INVx2_ASAP7_75t_L g1054 ( 
.A(n_971),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_L g1055 ( 
.A(n_966),
.B(n_567),
.Y(n_1055)
);

A2O1A1Ixp33_ASAP7_75t_L g1056 ( 
.A1(n_991),
.A2(n_571),
.B(n_600),
.C(n_601),
.Y(n_1056)
);

OAI22xp5_ASAP7_75t_SL g1057 ( 
.A1(n_944),
.A2(n_833),
.B1(n_977),
.B2(n_996),
.Y(n_1057)
);

A2O1A1Ixp33_ASAP7_75t_SL g1058 ( 
.A1(n_951),
.A2(n_654),
.B(n_282),
.C(n_272),
.Y(n_1058)
);

OAI22xp5_ASAP7_75t_L g1059 ( 
.A1(n_906),
.A2(n_252),
.B1(n_258),
.B2(n_654),
.Y(n_1059)
);

NOR2xp33_ASAP7_75t_R g1060 ( 
.A(n_891),
.B(n_962),
.Y(n_1060)
);

NAND3xp33_ASAP7_75t_L g1061 ( 
.A(n_847),
.B(n_331),
.C(n_228),
.Y(n_1061)
);

AOI21xp5_ASAP7_75t_L g1062 ( 
.A1(n_970),
.A2(n_638),
.B(n_579),
.Y(n_1062)
);

BUFx6f_ASAP7_75t_L g1063 ( 
.A(n_919),
.Y(n_1063)
);

INVx1_ASAP7_75t_L g1064 ( 
.A(n_924),
.Y(n_1064)
);

BUFx6f_ASAP7_75t_L g1065 ( 
.A(n_919),
.Y(n_1065)
);

NAND2xp33_ASAP7_75t_L g1066 ( 
.A(n_826),
.B(n_221),
.Y(n_1066)
);

AOI21xp5_ASAP7_75t_L g1067 ( 
.A1(n_970),
.A2(n_638),
.B(n_579),
.Y(n_1067)
);

OAI22xp5_ASAP7_75t_L g1068 ( 
.A1(n_840),
.A2(n_252),
.B1(n_258),
.B2(n_654),
.Y(n_1068)
);

A2O1A1Ixp33_ASAP7_75t_L g1069 ( 
.A1(n_918),
.A2(n_224),
.B(n_229),
.C(n_230),
.Y(n_1069)
);

NAND2xp5_ASAP7_75t_L g1070 ( 
.A(n_840),
.B(n_564),
.Y(n_1070)
);

AND2x2_ASAP7_75t_L g1071 ( 
.A(n_893),
.B(n_307),
.Y(n_1071)
);

INVx2_ASAP7_75t_L g1072 ( 
.A(n_980),
.Y(n_1072)
);

OAI22xp5_ASAP7_75t_SL g1073 ( 
.A1(n_875),
.A2(n_231),
.B1(n_246),
.B2(n_327),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_L g1074 ( 
.A(n_879),
.B(n_564),
.Y(n_1074)
);

O2A1O1Ixp33_ASAP7_75t_L g1075 ( 
.A1(n_842),
.A2(n_307),
.B(n_8),
.C(n_11),
.Y(n_1075)
);

AOI22xp33_ASAP7_75t_L g1076 ( 
.A1(n_990),
.A2(n_221),
.B1(n_310),
.B2(n_307),
.Y(n_1076)
);

NAND2xp5_ASAP7_75t_L g1077 ( 
.A(n_975),
.B(n_579),
.Y(n_1077)
);

NAND2xp5_ASAP7_75t_SL g1078 ( 
.A(n_826),
.B(n_301),
.Y(n_1078)
);

INVx1_ASAP7_75t_L g1079 ( 
.A(n_861),
.Y(n_1079)
);

INVx2_ASAP7_75t_L g1080 ( 
.A(n_981),
.Y(n_1080)
);

O2A1O1Ixp33_ASAP7_75t_L g1081 ( 
.A1(n_982),
.A2(n_3),
.B(n_11),
.C(n_14),
.Y(n_1081)
);

AOI22xp33_ASAP7_75t_L g1082 ( 
.A1(n_990),
.A2(n_310),
.B1(n_252),
.B2(n_258),
.Y(n_1082)
);

BUFx2_ASAP7_75t_L g1083 ( 
.A(n_939),
.Y(n_1083)
);

NOR2xp33_ASAP7_75t_R g1084 ( 
.A(n_916),
.B(n_256),
.Y(n_1084)
);

NAND2xp5_ASAP7_75t_L g1085 ( 
.A(n_862),
.B(n_308),
.Y(n_1085)
);

NOR2xp33_ASAP7_75t_L g1086 ( 
.A(n_927),
.B(n_298),
.Y(n_1086)
);

AOI22xp33_ASAP7_75t_L g1087 ( 
.A1(n_937),
.A2(n_310),
.B1(n_258),
.B2(n_303),
.Y(n_1087)
);

BUFx12f_ASAP7_75t_L g1088 ( 
.A(n_949),
.Y(n_1088)
);

INVx1_ASAP7_75t_L g1089 ( 
.A(n_863),
.Y(n_1089)
);

NAND2xp5_ASAP7_75t_L g1090 ( 
.A(n_864),
.B(n_309),
.Y(n_1090)
);

NOR2xp67_ASAP7_75t_L g1091 ( 
.A(n_903),
.B(n_262),
.Y(n_1091)
);

INVx2_ASAP7_75t_L g1092 ( 
.A(n_983),
.Y(n_1092)
);

OAI22xp5_ASAP7_75t_L g1093 ( 
.A1(n_976),
.A2(n_985),
.B1(n_978),
.B2(n_920),
.Y(n_1093)
);

AOI22xp5_ASAP7_75t_L g1094 ( 
.A1(n_892),
.A2(n_940),
.B1(n_831),
.B2(n_929),
.Y(n_1094)
);

BUFx6f_ASAP7_75t_L g1095 ( 
.A(n_956),
.Y(n_1095)
);

INVx1_ASAP7_75t_L g1096 ( 
.A(n_865),
.Y(n_1096)
);

BUFx6f_ASAP7_75t_L g1097 ( 
.A(n_956),
.Y(n_1097)
);

OAI21x1_ASAP7_75t_L g1098 ( 
.A1(n_844),
.A2(n_654),
.B(n_578),
.Y(n_1098)
);

INVx2_ASAP7_75t_L g1099 ( 
.A(n_871),
.Y(n_1099)
);

NAND2xp5_ASAP7_75t_L g1100 ( 
.A(n_978),
.B(n_578),
.Y(n_1100)
);

NOR2xp33_ASAP7_75t_R g1101 ( 
.A(n_907),
.B(n_266),
.Y(n_1101)
);

AOI21x1_ASAP7_75t_L g1102 ( 
.A1(n_985),
.A2(n_578),
.B(n_564),
.Y(n_1102)
);

A2O1A1Ixp33_ASAP7_75t_L g1103 ( 
.A1(n_870),
.A2(n_292),
.B(n_267),
.C(n_578),
.Y(n_1103)
);

O2A1O1Ixp33_ASAP7_75t_L g1104 ( 
.A1(n_880),
.A2(n_3),
.B(n_17),
.C(n_25),
.Y(n_1104)
);

NAND2xp5_ASAP7_75t_SL g1105 ( 
.A(n_827),
.B(n_310),
.Y(n_1105)
);

O2A1O1Ixp33_ASAP7_75t_L g1106 ( 
.A1(n_880),
.A2(n_17),
.B(n_27),
.C(n_29),
.Y(n_1106)
);

O2A1O1Ixp5_ASAP7_75t_L g1107 ( 
.A1(n_894),
.A2(n_310),
.B(n_97),
.C(n_104),
.Y(n_1107)
);

INVx3_ASAP7_75t_L g1108 ( 
.A(n_997),
.Y(n_1108)
);

AND2x4_ASAP7_75t_L g1109 ( 
.A(n_910),
.B(n_92),
.Y(n_1109)
);

OAI21xp5_ASAP7_75t_L g1110 ( 
.A1(n_934),
.A2(n_310),
.B(n_91),
.Y(n_1110)
);

INVx2_ASAP7_75t_L g1111 ( 
.A(n_876),
.Y(n_1111)
);

NAND2xp5_ASAP7_75t_L g1112 ( 
.A(n_934),
.B(n_310),
.Y(n_1112)
);

INVx2_ASAP7_75t_L g1113 ( 
.A(n_885),
.Y(n_1113)
);

XNOR2x2_ASAP7_75t_SL g1114 ( 
.A(n_972),
.B(n_33),
.Y(n_1114)
);

O2A1O1Ixp33_ASAP7_75t_SL g1115 ( 
.A1(n_984),
.A2(n_106),
.B(n_156),
.C(n_150),
.Y(n_1115)
);

INVx1_ASAP7_75t_L g1116 ( 
.A(n_878),
.Y(n_1116)
);

OAI22xp5_ASAP7_75t_L g1117 ( 
.A1(n_838),
.A2(n_34),
.B1(n_38),
.B2(n_40),
.Y(n_1117)
);

A2O1A1Ixp33_ASAP7_75t_L g1118 ( 
.A1(n_883),
.A2(n_38),
.B(n_41),
.C(n_42),
.Y(n_1118)
);

AOI22xp33_ASAP7_75t_L g1119 ( 
.A1(n_937),
.A2(n_940),
.B1(n_849),
.B2(n_857),
.Y(n_1119)
);

O2A1O1Ixp33_ASAP7_75t_L g1120 ( 
.A1(n_940),
.A2(n_42),
.B(n_43),
.C(n_44),
.Y(n_1120)
);

INVx2_ASAP7_75t_L g1121 ( 
.A(n_886),
.Y(n_1121)
);

O2A1O1Ixp33_ASAP7_75t_L g1122 ( 
.A1(n_889),
.A2(n_43),
.B(n_44),
.C(n_45),
.Y(n_1122)
);

INVx6_ASAP7_75t_L g1123 ( 
.A(n_827),
.Y(n_1123)
);

OR2x6_ASAP7_75t_SL g1124 ( 
.A(n_933),
.B(n_45),
.Y(n_1124)
);

INVx1_ASAP7_75t_L g1125 ( 
.A(n_890),
.Y(n_1125)
);

AOI21xp5_ASAP7_75t_L g1126 ( 
.A1(n_989),
.A2(n_116),
.B(n_142),
.Y(n_1126)
);

NOR2xp33_ASAP7_75t_SL g1127 ( 
.A(n_884),
.B(n_115),
.Y(n_1127)
);

INVx1_ASAP7_75t_L g1128 ( 
.A(n_905),
.Y(n_1128)
);

CKINVDCx6p67_ASAP7_75t_R g1129 ( 
.A(n_931),
.Y(n_1129)
);

NOR2xp33_ASAP7_75t_L g1130 ( 
.A(n_892),
.B(n_47),
.Y(n_1130)
);

BUFx12f_ASAP7_75t_L g1131 ( 
.A(n_921),
.Y(n_1131)
);

HB1xp67_ASAP7_75t_L g1132 ( 
.A(n_943),
.Y(n_1132)
);

INVx1_ASAP7_75t_L g1133 ( 
.A(n_908),
.Y(n_1133)
);

BUFx2_ASAP7_75t_L g1134 ( 
.A(n_877),
.Y(n_1134)
);

INVx1_ASAP7_75t_L g1135 ( 
.A(n_935),
.Y(n_1135)
);

OAI22xp5_ASAP7_75t_L g1136 ( 
.A1(n_895),
.A2(n_47),
.B1(n_49),
.B2(n_58),
.Y(n_1136)
);

BUFx2_ASAP7_75t_L g1137 ( 
.A(n_877),
.Y(n_1137)
);

CKINVDCx5p33_ASAP7_75t_R g1138 ( 
.A(n_986),
.Y(n_1138)
);

A2O1A1Ixp33_ASAP7_75t_SL g1139 ( 
.A1(n_994),
.A2(n_66),
.B(n_69),
.C(n_77),
.Y(n_1139)
);

AND2x6_ASAP7_75t_L g1140 ( 
.A(n_827),
.B(n_888),
.Y(n_1140)
);

OAI22xp5_ASAP7_75t_SL g1141 ( 
.A1(n_874),
.A2(n_82),
.B1(n_110),
.B2(n_119),
.Y(n_1141)
);

NAND2xp5_ASAP7_75t_SL g1142 ( 
.A(n_884),
.B(n_122),
.Y(n_1142)
);

NOR2xp33_ASAP7_75t_L g1143 ( 
.A(n_892),
.B(n_124),
.Y(n_1143)
);

A2O1A1Ixp33_ASAP7_75t_SL g1144 ( 
.A1(n_1007),
.A2(n_963),
.B(n_987),
.C(n_888),
.Y(n_1144)
);

O2A1O1Ixp33_ASAP7_75t_L g1145 ( 
.A1(n_889),
.A2(n_131),
.B(n_132),
.C(n_135),
.Y(n_1145)
);

A2O1A1Ixp33_ASAP7_75t_L g1146 ( 
.A1(n_968),
.A2(n_136),
.B(n_159),
.C(n_868),
.Y(n_1146)
);

BUFx2_ASAP7_75t_L g1147 ( 
.A(n_877),
.Y(n_1147)
);

AOI21xp5_ASAP7_75t_L g1148 ( 
.A1(n_989),
.A2(n_999),
.B(n_1000),
.Y(n_1148)
);

OAI22xp5_ASAP7_75t_L g1149 ( 
.A1(n_895),
.A2(n_897),
.B1(n_999),
.B2(n_1000),
.Y(n_1149)
);

NAND2xp5_ASAP7_75t_L g1150 ( 
.A(n_941),
.B(n_952),
.Y(n_1150)
);

A2O1A1Ixp33_ASAP7_75t_L g1151 ( 
.A1(n_922),
.A2(n_936),
.B(n_954),
.C(n_941),
.Y(n_1151)
);

INVx1_ASAP7_75t_L g1152 ( 
.A(n_942),
.Y(n_1152)
);

A2O1A1Ixp33_ASAP7_75t_L g1153 ( 
.A1(n_952),
.A2(n_859),
.B(n_969),
.C(n_897),
.Y(n_1153)
);

INVx1_ASAP7_75t_L g1154 ( 
.A(n_904),
.Y(n_1154)
);

INVx1_ASAP7_75t_L g1155 ( 
.A(n_904),
.Y(n_1155)
);

AND2x2_ASAP7_75t_L g1156 ( 
.A(n_843),
.B(n_855),
.Y(n_1156)
);

BUFx6f_ASAP7_75t_L g1157 ( 
.A(n_956),
.Y(n_1157)
);

NAND2xp5_ASAP7_75t_SL g1158 ( 
.A(n_828),
.B(n_959),
.Y(n_1158)
);

NAND2xp5_ASAP7_75t_SL g1159 ( 
.A(n_828),
.B(n_959),
.Y(n_1159)
);

AND2x6_ASAP7_75t_SL g1160 ( 
.A(n_937),
.B(n_960),
.Y(n_1160)
);

AOI21xp5_ASAP7_75t_L g1161 ( 
.A1(n_1150),
.A2(n_828),
.B(n_959),
.Y(n_1161)
);

NAND2xp5_ASAP7_75t_L g1162 ( 
.A(n_1038),
.B(n_899),
.Y(n_1162)
);

AO31x2_ASAP7_75t_L g1163 ( 
.A1(n_1068),
.A2(n_998),
.A3(n_873),
.B(n_854),
.Y(n_1163)
);

AOI21xp5_ASAP7_75t_L g1164 ( 
.A1(n_1012),
.A2(n_828),
.B(n_959),
.Y(n_1164)
);

INVx1_ASAP7_75t_L g1165 ( 
.A(n_1025),
.Y(n_1165)
);

AOI22xp5_ASAP7_75t_L g1166 ( 
.A1(n_1017),
.A2(n_872),
.B1(n_856),
.B2(n_974),
.Y(n_1166)
);

AOI221xp5_ASAP7_75t_L g1167 ( 
.A1(n_1039),
.A2(n_1003),
.B1(n_867),
.B2(n_900),
.C(n_914),
.Y(n_1167)
);

AOI21xp5_ASAP7_75t_L g1168 ( 
.A1(n_1148),
.A2(n_1149),
.B(n_1093),
.Y(n_1168)
);

NAND2xp5_ASAP7_75t_L g1169 ( 
.A(n_1049),
.B(n_1020),
.Y(n_1169)
);

BUFx3_ASAP7_75t_L g1170 ( 
.A(n_1027),
.Y(n_1170)
);

OAI21xp5_ASAP7_75t_L g1171 ( 
.A1(n_1044),
.A2(n_852),
.B(n_854),
.Y(n_1171)
);

A2O1A1Ixp33_ASAP7_75t_L g1172 ( 
.A1(n_1110),
.A2(n_950),
.B(n_965),
.C(n_912),
.Y(n_1172)
);

BUFx6f_ASAP7_75t_L g1173 ( 
.A(n_1011),
.Y(n_1173)
);

NOR2xp33_ASAP7_75t_L g1174 ( 
.A(n_1043),
.B(n_993),
.Y(n_1174)
);

AOI21xp5_ASAP7_75t_L g1175 ( 
.A1(n_1149),
.A2(n_909),
.B(n_912),
.Y(n_1175)
);

NAND2xp5_ASAP7_75t_L g1176 ( 
.A(n_1045),
.B(n_914),
.Y(n_1176)
);

AND2x6_ASAP7_75t_L g1177 ( 
.A(n_1109),
.B(n_967),
.Y(n_1177)
);

OAI21xp5_ASAP7_75t_L g1178 ( 
.A1(n_1151),
.A2(n_852),
.B(n_873),
.Y(n_1178)
);

BUFx4f_ASAP7_75t_L g1179 ( 
.A(n_1131),
.Y(n_1179)
);

O2A1O1Ixp5_ASAP7_75t_L g1180 ( 
.A1(n_1110),
.A2(n_835),
.B(n_836),
.C(n_841),
.Y(n_1180)
);

O2A1O1Ixp5_ASAP7_75t_L g1181 ( 
.A1(n_1021),
.A2(n_961),
.B(n_1005),
.C(n_850),
.Y(n_1181)
);

AOI21xp5_ASAP7_75t_L g1182 ( 
.A1(n_1093),
.A2(n_912),
.B(n_909),
.Y(n_1182)
);

AOI21x1_ASAP7_75t_L g1183 ( 
.A1(n_1102),
.A2(n_844),
.B(n_845),
.Y(n_1183)
);

INVx5_ASAP7_75t_L g1184 ( 
.A(n_1140),
.Y(n_1184)
);

AND2x2_ASAP7_75t_L g1185 ( 
.A(n_1024),
.B(n_967),
.Y(n_1185)
);

AOI21xp5_ASAP7_75t_L g1186 ( 
.A1(n_1028),
.A2(n_912),
.B(n_909),
.Y(n_1186)
);

INVx1_ASAP7_75t_L g1187 ( 
.A(n_1064),
.Y(n_1187)
);

INVx1_ASAP7_75t_L g1188 ( 
.A(n_1079),
.Y(n_1188)
);

AO31x2_ASAP7_75t_L g1189 ( 
.A1(n_1068),
.A2(n_845),
.A3(n_850),
.B(n_1004),
.Y(n_1189)
);

NAND2xp5_ASAP7_75t_L g1190 ( 
.A(n_1037),
.B(n_872),
.Y(n_1190)
);

AND2x2_ASAP7_75t_L g1191 ( 
.A(n_1031),
.B(n_1004),
.Y(n_1191)
);

CKINVDCx11_ASAP7_75t_R g1192 ( 
.A(n_1088),
.Y(n_1192)
);

INVx3_ASAP7_75t_L g1193 ( 
.A(n_1010),
.Y(n_1193)
);

INVx2_ASAP7_75t_L g1194 ( 
.A(n_1089),
.Y(n_1194)
);

OAI21x1_ASAP7_75t_L g1195 ( 
.A1(n_1098),
.A2(n_945),
.B(n_1006),
.Y(n_1195)
);

AOI21xp5_ASAP7_75t_SL g1196 ( 
.A1(n_1153),
.A2(n_866),
.B(n_869),
.Y(n_1196)
);

A2O1A1Ixp33_ASAP7_75t_L g1197 ( 
.A1(n_1021),
.A2(n_909),
.B(n_1001),
.C(n_872),
.Y(n_1197)
);

BUFx3_ASAP7_75t_L g1198 ( 
.A(n_1033),
.Y(n_1198)
);

INVxp67_ASAP7_75t_L g1199 ( 
.A(n_1051),
.Y(n_1199)
);

BUFx4_ASAP7_75t_SL g1200 ( 
.A(n_1160),
.Y(n_1200)
);

INVx1_ASAP7_75t_L g1201 ( 
.A(n_1096),
.Y(n_1201)
);

AOI21xp5_ASAP7_75t_L g1202 ( 
.A1(n_1014),
.A2(n_988),
.B(n_866),
.Y(n_1202)
);

OAI21x1_ASAP7_75t_SL g1203 ( 
.A1(n_1120),
.A2(n_1145),
.B(n_1081),
.Y(n_1203)
);

INVx3_ASAP7_75t_L g1204 ( 
.A(n_1010),
.Y(n_1204)
);

NOR2xp67_ASAP7_75t_L g1205 ( 
.A(n_1037),
.B(n_913),
.Y(n_1205)
);

AO31x2_ASAP7_75t_L g1206 ( 
.A1(n_1056),
.A2(n_913),
.A3(n_872),
.B(n_988),
.Y(n_1206)
);

AND2x4_ASAP7_75t_L g1207 ( 
.A(n_1035),
.B(n_1134),
.Y(n_1207)
);

AND2x4_ASAP7_75t_L g1208 ( 
.A(n_1137),
.B(n_1147),
.Y(n_1208)
);

AOI21xp5_ASAP7_75t_L g1209 ( 
.A1(n_1016),
.A2(n_1026),
.B(n_1029),
.Y(n_1209)
);

AOI21xp5_ASAP7_75t_L g1210 ( 
.A1(n_1026),
.A2(n_1029),
.B(n_1022),
.Y(n_1210)
);

INVx5_ASAP7_75t_L g1211 ( 
.A(n_1140),
.Y(n_1211)
);

AOI21x1_ASAP7_75t_L g1212 ( 
.A1(n_1112),
.A2(n_1022),
.B(n_1070),
.Y(n_1212)
);

AOI21xp5_ASAP7_75t_SL g1213 ( 
.A1(n_1158),
.A2(n_1159),
.B(n_1146),
.Y(n_1213)
);

AOI21x1_ASAP7_75t_L g1214 ( 
.A1(n_1112),
.A2(n_1070),
.B(n_1074),
.Y(n_1214)
);

INVx2_ASAP7_75t_SL g1215 ( 
.A(n_1156),
.Y(n_1215)
);

AOI21xp33_ASAP7_75t_L g1216 ( 
.A1(n_1086),
.A2(n_1090),
.B(n_1085),
.Y(n_1216)
);

OAI21xp5_ASAP7_75t_L g1217 ( 
.A1(n_1062),
.A2(n_1067),
.B(n_1023),
.Y(n_1217)
);

AOI211x1_ASAP7_75t_L g1218 ( 
.A1(n_1117),
.A2(n_1136),
.B(n_1116),
.C(n_1125),
.Y(n_1218)
);

NAND2xp5_ASAP7_75t_L g1219 ( 
.A(n_1042),
.B(n_1019),
.Y(n_1219)
);

NOR2xp33_ASAP7_75t_L g1220 ( 
.A(n_1057),
.B(n_1138),
.Y(n_1220)
);

OAI21xp5_ASAP7_75t_L g1221 ( 
.A1(n_1023),
.A2(n_1077),
.B(n_1100),
.Y(n_1221)
);

CKINVDCx20_ASAP7_75t_R g1222 ( 
.A(n_1129),
.Y(n_1222)
);

AOI21xp5_ASAP7_75t_L g1223 ( 
.A1(n_1144),
.A2(n_1100),
.B(n_1077),
.Y(n_1223)
);

OAI21x1_ASAP7_75t_L g1224 ( 
.A1(n_1055),
.A2(n_1034),
.B(n_1048),
.Y(n_1224)
);

AOI21xp5_ASAP7_75t_SL g1225 ( 
.A1(n_1143),
.A2(n_1109),
.B(n_1103),
.Y(n_1225)
);

AOI21xp5_ASAP7_75t_L g1226 ( 
.A1(n_1018),
.A2(n_1013),
.B(n_1055),
.Y(n_1226)
);

AOI21xp5_ASAP7_75t_L g1227 ( 
.A1(n_1046),
.A2(n_1050),
.B(n_1036),
.Y(n_1227)
);

INVx1_ASAP7_75t_L g1228 ( 
.A(n_1128),
.Y(n_1228)
);

INVx3_ASAP7_75t_L g1229 ( 
.A(n_1140),
.Y(n_1229)
);

INVx3_ASAP7_75t_L g1230 ( 
.A(n_1140),
.Y(n_1230)
);

NAND2xp5_ASAP7_75t_L g1231 ( 
.A(n_1094),
.B(n_1119),
.Y(n_1231)
);

HB1xp67_ASAP7_75t_L g1232 ( 
.A(n_1083),
.Y(n_1232)
);

O2A1O1Ixp33_ASAP7_75t_SL g1233 ( 
.A1(n_1139),
.A2(n_1069),
.B(n_1142),
.C(n_1118),
.Y(n_1233)
);

HB1xp67_ASAP7_75t_L g1234 ( 
.A(n_1132),
.Y(n_1234)
);

OAI21xp5_ASAP7_75t_L g1235 ( 
.A1(n_1059),
.A2(n_1107),
.B(n_1126),
.Y(n_1235)
);

NAND2xp5_ASAP7_75t_SL g1236 ( 
.A(n_1060),
.B(n_1101),
.Y(n_1236)
);

NAND2xp5_ASAP7_75t_L g1237 ( 
.A(n_1133),
.B(n_1135),
.Y(n_1237)
);

OAI21x1_ASAP7_75t_L g1238 ( 
.A1(n_1105),
.A2(n_1040),
.B(n_1032),
.Y(n_1238)
);

NAND2xp5_ASAP7_75t_L g1239 ( 
.A(n_1152),
.B(n_1092),
.Y(n_1239)
);

NAND3xp33_ASAP7_75t_L g1240 ( 
.A(n_1075),
.B(n_1106),
.C(n_1104),
.Y(n_1240)
);

OAI21x1_ASAP7_75t_L g1241 ( 
.A1(n_1030),
.A2(n_1059),
.B(n_1154),
.Y(n_1241)
);

OAI21xp5_ASAP7_75t_L g1242 ( 
.A1(n_1082),
.A2(n_1076),
.B(n_1117),
.Y(n_1242)
);

AOI21xp5_ASAP7_75t_L g1243 ( 
.A1(n_1058),
.A2(n_1127),
.B(n_1052),
.Y(n_1243)
);

AOI21xp5_ASAP7_75t_SL g1244 ( 
.A1(n_1136),
.A2(n_1122),
.B(n_1157),
.Y(n_1244)
);

OAI21x1_ASAP7_75t_L g1245 ( 
.A1(n_1155),
.A2(n_1108),
.B(n_1015),
.Y(n_1245)
);

O2A1O1Ixp33_ASAP7_75t_L g1246 ( 
.A1(n_1130),
.A2(n_1078),
.B(n_1115),
.C(n_1071),
.Y(n_1246)
);

AO21x2_ASAP7_75t_L g1247 ( 
.A1(n_1066),
.A2(n_1072),
.B(n_1111),
.Y(n_1247)
);

OAI21x1_ASAP7_75t_L g1248 ( 
.A1(n_1015),
.A2(n_1108),
.B(n_1041),
.Y(n_1248)
);

AOI21xp5_ASAP7_75t_L g1249 ( 
.A1(n_1053),
.A2(n_1121),
.B(n_1054),
.Y(n_1249)
);

NAND2xp5_ASAP7_75t_SL g1250 ( 
.A(n_1084),
.B(n_1091),
.Y(n_1250)
);

AO22x2_ASAP7_75t_L g1251 ( 
.A1(n_1114),
.A2(n_1061),
.B1(n_1113),
.B2(n_1080),
.Y(n_1251)
);

AOI21xp5_ASAP7_75t_L g1252 ( 
.A1(n_1053),
.A2(n_1099),
.B(n_1041),
.Y(n_1252)
);

NAND2x1_ASAP7_75t_L g1253 ( 
.A(n_1123),
.B(n_1011),
.Y(n_1253)
);

NOR4xp25_ASAP7_75t_L g1254 ( 
.A(n_1087),
.B(n_1141),
.C(n_1124),
.D(n_1073),
.Y(n_1254)
);

OAI21x1_ASAP7_75t_L g1255 ( 
.A1(n_1123),
.A2(n_1011),
.B(n_1063),
.Y(n_1255)
);

NAND2xp5_ASAP7_75t_L g1256 ( 
.A(n_1123),
.B(n_1157),
.Y(n_1256)
);

OAI21x1_ASAP7_75t_L g1257 ( 
.A1(n_1063),
.A2(n_1065),
.B(n_1095),
.Y(n_1257)
);

OAI22xp5_ASAP7_75t_L g1258 ( 
.A1(n_1063),
.A2(n_1065),
.B1(n_1095),
.B2(n_1097),
.Y(n_1258)
);

OAI22xp5_ASAP7_75t_L g1259 ( 
.A1(n_1095),
.A2(n_1150),
.B1(n_1038),
.B2(n_881),
.Y(n_1259)
);

NAND3xp33_ASAP7_75t_L g1260 ( 
.A(n_1097),
.B(n_839),
.C(n_688),
.Y(n_1260)
);

O2A1O1Ixp5_ASAP7_75t_SL g1261 ( 
.A1(n_1097),
.A2(n_1136),
.B(n_1110),
.C(n_1068),
.Y(n_1261)
);

NAND2xp5_ASAP7_75t_L g1262 ( 
.A(n_1038),
.B(n_839),
.Y(n_1262)
);

AO31x2_ASAP7_75t_L g1263 ( 
.A1(n_1068),
.A2(n_1056),
.A3(n_1059),
.B(n_1149),
.Y(n_1263)
);

OR2x2_ASAP7_75t_L g1264 ( 
.A(n_1038),
.B(n_846),
.Y(n_1264)
);

NAND2xp5_ASAP7_75t_L g1265 ( 
.A(n_1038),
.B(n_839),
.Y(n_1265)
);

INVx3_ASAP7_75t_L g1266 ( 
.A(n_1010),
.Y(n_1266)
);

OAI22xp5_ASAP7_75t_L g1267 ( 
.A1(n_1150),
.A2(n_661),
.B1(n_1038),
.B2(n_834),
.Y(n_1267)
);

OR2x2_ASAP7_75t_L g1268 ( 
.A(n_1038),
.B(n_846),
.Y(n_1268)
);

AO31x2_ASAP7_75t_L g1269 ( 
.A1(n_1068),
.A2(n_1056),
.A3(n_1059),
.B(n_1149),
.Y(n_1269)
);

INVx1_ASAP7_75t_SL g1270 ( 
.A(n_1043),
.Y(n_1270)
);

NOR2xp67_ASAP7_75t_L g1271 ( 
.A(n_1038),
.B(n_522),
.Y(n_1271)
);

AOI21xp5_ASAP7_75t_L g1272 ( 
.A1(n_1150),
.A2(n_682),
.B(n_881),
.Y(n_1272)
);

OAI21x1_ASAP7_75t_L g1273 ( 
.A1(n_1098),
.A2(n_1047),
.B(n_1102),
.Y(n_1273)
);

NAND2xp5_ASAP7_75t_SL g1274 ( 
.A(n_1017),
.B(n_915),
.Y(n_1274)
);

INVx2_ASAP7_75t_L g1275 ( 
.A(n_1025),
.Y(n_1275)
);

AOI21xp5_ASAP7_75t_L g1276 ( 
.A1(n_1150),
.A2(n_682),
.B(n_881),
.Y(n_1276)
);

OAI21x1_ASAP7_75t_L g1277 ( 
.A1(n_1098),
.A2(n_1047),
.B(n_1102),
.Y(n_1277)
);

OAI21xp5_ASAP7_75t_L g1278 ( 
.A1(n_1148),
.A2(n_1044),
.B(n_1149),
.Y(n_1278)
);

OAI21x1_ASAP7_75t_L g1279 ( 
.A1(n_1098),
.A2(n_1047),
.B(n_1102),
.Y(n_1279)
);

OAI22x1_ASAP7_75t_L g1280 ( 
.A1(n_1094),
.A2(n_565),
.B1(n_960),
.B2(n_982),
.Y(n_1280)
);

INVx1_ASAP7_75t_L g1281 ( 
.A(n_1025),
.Y(n_1281)
);

INVx1_ASAP7_75t_L g1282 ( 
.A(n_1025),
.Y(n_1282)
);

INVx2_ASAP7_75t_L g1283 ( 
.A(n_1025),
.Y(n_1283)
);

AND2x4_ASAP7_75t_L g1284 ( 
.A(n_1035),
.B(n_939),
.Y(n_1284)
);

INVxp67_ASAP7_75t_L g1285 ( 
.A(n_1043),
.Y(n_1285)
);

OAI21xp33_ASAP7_75t_SL g1286 ( 
.A1(n_1150),
.A2(n_1012),
.B(n_881),
.Y(n_1286)
);

AOI21xp5_ASAP7_75t_L g1287 ( 
.A1(n_1150),
.A2(n_682),
.B(n_881),
.Y(n_1287)
);

BUFx8_ASAP7_75t_SL g1288 ( 
.A(n_1088),
.Y(n_1288)
);

INVx2_ASAP7_75t_L g1289 ( 
.A(n_1025),
.Y(n_1289)
);

INVx2_ASAP7_75t_L g1290 ( 
.A(n_1025),
.Y(n_1290)
);

OAI22xp5_ASAP7_75t_L g1291 ( 
.A1(n_1150),
.A2(n_661),
.B1(n_1038),
.B2(n_834),
.Y(n_1291)
);

AND2x2_ASAP7_75t_L g1292 ( 
.A(n_1045),
.B(n_915),
.Y(n_1292)
);

OAI21xp5_ASAP7_75t_L g1293 ( 
.A1(n_1148),
.A2(n_1044),
.B(n_1149),
.Y(n_1293)
);

AO21x2_ASAP7_75t_L g1294 ( 
.A1(n_1110),
.A2(n_1148),
.B(n_1047),
.Y(n_1294)
);

AO31x2_ASAP7_75t_L g1295 ( 
.A1(n_1068),
.A2(n_1056),
.A3(n_1059),
.B(n_1149),
.Y(n_1295)
);

NAND2xp5_ASAP7_75t_L g1296 ( 
.A(n_1038),
.B(n_839),
.Y(n_1296)
);

NAND2xp5_ASAP7_75t_L g1297 ( 
.A(n_1038),
.B(n_839),
.Y(n_1297)
);

O2A1O1Ixp5_ASAP7_75t_L g1298 ( 
.A1(n_1110),
.A2(n_858),
.B(n_716),
.C(n_686),
.Y(n_1298)
);

AOI21xp5_ASAP7_75t_L g1299 ( 
.A1(n_1150),
.A2(n_682),
.B(n_881),
.Y(n_1299)
);

A2O1A1Ixp33_ASAP7_75t_L g1300 ( 
.A1(n_1017),
.A2(n_1039),
.B(n_839),
.C(n_661),
.Y(n_1300)
);

AO31x2_ASAP7_75t_L g1301 ( 
.A1(n_1068),
.A2(n_1056),
.A3(n_1059),
.B(n_1149),
.Y(n_1301)
);

NOR2xp33_ASAP7_75t_L g1302 ( 
.A(n_1017),
.B(n_839),
.Y(n_1302)
);

AOI21x1_ASAP7_75t_L g1303 ( 
.A1(n_1102),
.A2(n_1047),
.B(n_1112),
.Y(n_1303)
);

BUFx6f_ASAP7_75t_L g1304 ( 
.A(n_1011),
.Y(n_1304)
);

AOI21xp5_ASAP7_75t_L g1305 ( 
.A1(n_1150),
.A2(n_682),
.B(n_881),
.Y(n_1305)
);

AOI21xp33_ASAP7_75t_L g1306 ( 
.A1(n_1039),
.A2(n_720),
.B(n_839),
.Y(n_1306)
);

AO31x2_ASAP7_75t_L g1307 ( 
.A1(n_1068),
.A2(n_1056),
.A3(n_1059),
.B(n_1149),
.Y(n_1307)
);

A2O1A1Ixp33_ASAP7_75t_L g1308 ( 
.A1(n_1017),
.A2(n_1039),
.B(n_839),
.C(n_661),
.Y(n_1308)
);

INVx2_ASAP7_75t_L g1309 ( 
.A(n_1025),
.Y(n_1309)
);

OA21x2_ASAP7_75t_L g1310 ( 
.A1(n_1110),
.A2(n_1148),
.B(n_1056),
.Y(n_1310)
);

NAND3x1_ASAP7_75t_L g1311 ( 
.A(n_1114),
.B(n_505),
.C(n_565),
.Y(n_1311)
);

AOI22xp5_ASAP7_75t_L g1312 ( 
.A1(n_1302),
.A2(n_1292),
.B1(n_1274),
.B2(n_1311),
.Y(n_1312)
);

BUFx3_ASAP7_75t_L g1313 ( 
.A(n_1170),
.Y(n_1313)
);

BUFx3_ASAP7_75t_L g1314 ( 
.A(n_1198),
.Y(n_1314)
);

BUFx2_ASAP7_75t_L g1315 ( 
.A(n_1208),
.Y(n_1315)
);

INVx1_ASAP7_75t_SL g1316 ( 
.A(n_1270),
.Y(n_1316)
);

AND2x2_ASAP7_75t_L g1317 ( 
.A(n_1191),
.B(n_1262),
.Y(n_1317)
);

INVx2_ASAP7_75t_L g1318 ( 
.A(n_1275),
.Y(n_1318)
);

INVx2_ASAP7_75t_L g1319 ( 
.A(n_1283),
.Y(n_1319)
);

INVx2_ASAP7_75t_L g1320 ( 
.A(n_1289),
.Y(n_1320)
);

INVx2_ASAP7_75t_L g1321 ( 
.A(n_1290),
.Y(n_1321)
);

OR2x2_ASAP7_75t_L g1322 ( 
.A(n_1169),
.B(n_1296),
.Y(n_1322)
);

O2A1O1Ixp33_ASAP7_75t_SL g1323 ( 
.A1(n_1172),
.A2(n_1300),
.B(n_1308),
.C(n_1306),
.Y(n_1323)
);

INVx1_ASAP7_75t_L g1324 ( 
.A(n_1309),
.Y(n_1324)
);

AO31x2_ASAP7_75t_L g1325 ( 
.A1(n_1168),
.A2(n_1223),
.A3(n_1197),
.B(n_1209),
.Y(n_1325)
);

AOI21xp5_ASAP7_75t_L g1326 ( 
.A1(n_1196),
.A2(n_1276),
.B(n_1272),
.Y(n_1326)
);

INVx1_ASAP7_75t_L g1327 ( 
.A(n_1165),
.Y(n_1327)
);

AOI21xp5_ASAP7_75t_L g1328 ( 
.A1(n_1287),
.A2(n_1305),
.B(n_1299),
.Y(n_1328)
);

OAI22xp5_ASAP7_75t_L g1329 ( 
.A1(n_1297),
.A2(n_1260),
.B1(n_1231),
.B2(n_1162),
.Y(n_1329)
);

OAI21x1_ASAP7_75t_L g1330 ( 
.A1(n_1303),
.A2(n_1202),
.B(n_1195),
.Y(n_1330)
);

AOI21xp5_ASAP7_75t_L g1331 ( 
.A1(n_1278),
.A2(n_1293),
.B(n_1267),
.Y(n_1331)
);

OAI22xp5_ASAP7_75t_L g1332 ( 
.A1(n_1260),
.A2(n_1176),
.B1(n_1268),
.B2(n_1264),
.Y(n_1332)
);

NAND2xp5_ASAP7_75t_L g1333 ( 
.A(n_1259),
.B(n_1216),
.Y(n_1333)
);

AND2x4_ASAP7_75t_L g1334 ( 
.A(n_1177),
.B(n_1208),
.Y(n_1334)
);

BUFx4_ASAP7_75t_SL g1335 ( 
.A(n_1222),
.Y(n_1335)
);

OAI21x1_ASAP7_75t_L g1336 ( 
.A1(n_1217),
.A2(n_1224),
.B(n_1214),
.Y(n_1336)
);

OAI21x1_ASAP7_75t_L g1337 ( 
.A1(n_1217),
.A2(n_1212),
.B(n_1186),
.Y(n_1337)
);

OAI21xp5_ASAP7_75t_L g1338 ( 
.A1(n_1298),
.A2(n_1291),
.B(n_1240),
.Y(n_1338)
);

CKINVDCx20_ASAP7_75t_R g1339 ( 
.A(n_1192),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_1187),
.Y(n_1340)
);

INVx1_ASAP7_75t_L g1341 ( 
.A(n_1188),
.Y(n_1341)
);

INVx1_ASAP7_75t_L g1342 ( 
.A(n_1201),
.Y(n_1342)
);

NOR2xp33_ASAP7_75t_L g1343 ( 
.A(n_1270),
.B(n_1285),
.Y(n_1343)
);

AO21x2_ASAP7_75t_L g1344 ( 
.A1(n_1235),
.A2(n_1293),
.B(n_1278),
.Y(n_1344)
);

OAI21x1_ASAP7_75t_L g1345 ( 
.A1(n_1175),
.A2(n_1182),
.B(n_1183),
.Y(n_1345)
);

OAI21x1_ASAP7_75t_L g1346 ( 
.A1(n_1241),
.A2(n_1221),
.B(n_1210),
.Y(n_1346)
);

OAI22xp5_ASAP7_75t_L g1347 ( 
.A1(n_1219),
.A2(n_1166),
.B1(n_1240),
.B2(n_1271),
.Y(n_1347)
);

INVx1_ASAP7_75t_L g1348 ( 
.A(n_1281),
.Y(n_1348)
);

HB1xp67_ASAP7_75t_L g1349 ( 
.A(n_1190),
.Y(n_1349)
);

OAI21x1_ASAP7_75t_L g1350 ( 
.A1(n_1221),
.A2(n_1227),
.B(n_1238),
.Y(n_1350)
);

INVx1_ASAP7_75t_L g1351 ( 
.A(n_1282),
.Y(n_1351)
);

NAND2x1p5_ASAP7_75t_L g1352 ( 
.A(n_1184),
.B(n_1211),
.Y(n_1352)
);

BUFx3_ASAP7_75t_L g1353 ( 
.A(n_1215),
.Y(n_1353)
);

INVx1_ASAP7_75t_L g1354 ( 
.A(n_1237),
.Y(n_1354)
);

INVx1_ASAP7_75t_L g1355 ( 
.A(n_1228),
.Y(n_1355)
);

OAI21xp5_ASAP7_75t_L g1356 ( 
.A1(n_1226),
.A2(n_1246),
.B(n_1261),
.Y(n_1356)
);

OAI21x1_ASAP7_75t_L g1357 ( 
.A1(n_1178),
.A2(n_1235),
.B(n_1171),
.Y(n_1357)
);

OAI21x1_ASAP7_75t_L g1358 ( 
.A1(n_1178),
.A2(n_1171),
.B(n_1164),
.Y(n_1358)
);

INVxp67_ASAP7_75t_L g1359 ( 
.A(n_1232),
.Y(n_1359)
);

OA21x2_ASAP7_75t_L g1360 ( 
.A1(n_1180),
.A2(n_1181),
.B(n_1167),
.Y(n_1360)
);

BUFx3_ASAP7_75t_L g1361 ( 
.A(n_1284),
.Y(n_1361)
);

OAI21x1_ASAP7_75t_L g1362 ( 
.A1(n_1243),
.A2(n_1245),
.B(n_1310),
.Y(n_1362)
);

BUFx3_ASAP7_75t_L g1363 ( 
.A(n_1253),
.Y(n_1363)
);

AND2x2_ASAP7_75t_L g1364 ( 
.A(n_1185),
.B(n_1251),
.Y(n_1364)
);

AO21x2_ASAP7_75t_L g1365 ( 
.A1(n_1294),
.A2(n_1205),
.B(n_1203),
.Y(n_1365)
);

NAND2x1p5_ASAP7_75t_L g1366 ( 
.A(n_1184),
.B(n_1211),
.Y(n_1366)
);

INVx2_ASAP7_75t_L g1367 ( 
.A(n_1247),
.Y(n_1367)
);

AND2x2_ASAP7_75t_L g1368 ( 
.A(n_1251),
.B(n_1207),
.Y(n_1368)
);

INVx1_ASAP7_75t_L g1369 ( 
.A(n_1239),
.Y(n_1369)
);

AND2x6_ASAP7_75t_L g1370 ( 
.A(n_1166),
.B(n_1229),
.Y(n_1370)
);

AND2x2_ASAP7_75t_L g1371 ( 
.A(n_1207),
.B(n_1254),
.Y(n_1371)
);

NOR2xp33_ASAP7_75t_L g1372 ( 
.A(n_1199),
.B(n_1234),
.Y(n_1372)
);

INVx2_ASAP7_75t_L g1373 ( 
.A(n_1247),
.Y(n_1373)
);

O2A1O1Ixp33_ASAP7_75t_L g1374 ( 
.A1(n_1254),
.A2(n_1242),
.B(n_1236),
.C(n_1250),
.Y(n_1374)
);

INVx2_ASAP7_75t_L g1375 ( 
.A(n_1163),
.Y(n_1375)
);

INVx2_ASAP7_75t_L g1376 ( 
.A(n_1163),
.Y(n_1376)
);

OR2x2_ASAP7_75t_L g1377 ( 
.A(n_1174),
.B(n_1280),
.Y(n_1377)
);

OAI21x1_ASAP7_75t_L g1378 ( 
.A1(n_1310),
.A2(n_1161),
.B(n_1249),
.Y(n_1378)
);

AOI22xp33_ASAP7_75t_L g1379 ( 
.A1(n_1242),
.A2(n_1271),
.B1(n_1286),
.B2(n_1177),
.Y(n_1379)
);

OAI21x1_ASAP7_75t_L g1380 ( 
.A1(n_1252),
.A2(n_1248),
.B(n_1213),
.Y(n_1380)
);

OAI221xp5_ASAP7_75t_L g1381 ( 
.A1(n_1225),
.A2(n_1244),
.B1(n_1220),
.B2(n_1286),
.C(n_1233),
.Y(n_1381)
);

AOI21xp33_ASAP7_75t_L g1382 ( 
.A1(n_1294),
.A2(n_1205),
.B(n_1258),
.Y(n_1382)
);

OA21x2_ASAP7_75t_L g1383 ( 
.A1(n_1263),
.A2(n_1307),
.B(n_1301),
.Y(n_1383)
);

OAI21xp5_ASAP7_75t_L g1384 ( 
.A1(n_1177),
.A2(n_1257),
.B(n_1255),
.Y(n_1384)
);

INVx1_ASAP7_75t_L g1385 ( 
.A(n_1218),
.Y(n_1385)
);

NOR2xp33_ASAP7_75t_L g1386 ( 
.A(n_1256),
.B(n_1266),
.Y(n_1386)
);

OA21x2_ASAP7_75t_L g1387 ( 
.A1(n_1263),
.A2(n_1307),
.B(n_1301),
.Y(n_1387)
);

OAI21x1_ASAP7_75t_L g1388 ( 
.A1(n_1229),
.A2(n_1230),
.B(n_1266),
.Y(n_1388)
);

NAND3xp33_ASAP7_75t_L g1389 ( 
.A(n_1218),
.B(n_1211),
.C(n_1184),
.Y(n_1389)
);

NOR2xp67_ASAP7_75t_L g1390 ( 
.A(n_1193),
.B(n_1204),
.Y(n_1390)
);

OAI21x1_ASAP7_75t_L g1391 ( 
.A1(n_1230),
.A2(n_1204),
.B(n_1193),
.Y(n_1391)
);

OR2x6_ASAP7_75t_L g1392 ( 
.A(n_1173),
.B(n_1304),
.Y(n_1392)
);

INVx2_ASAP7_75t_SL g1393 ( 
.A(n_1179),
.Y(n_1393)
);

OAI21x1_ASAP7_75t_L g1394 ( 
.A1(n_1206),
.A2(n_1163),
.B(n_1269),
.Y(n_1394)
);

OAI21x1_ASAP7_75t_L g1395 ( 
.A1(n_1206),
.A2(n_1269),
.B(n_1301),
.Y(n_1395)
);

AND2x4_ASAP7_75t_L g1396 ( 
.A(n_1173),
.B(n_1304),
.Y(n_1396)
);

OAI21x1_ASAP7_75t_L g1397 ( 
.A1(n_1206),
.A2(n_1269),
.B(n_1295),
.Y(n_1397)
);

INVx2_ASAP7_75t_L g1398 ( 
.A(n_1189),
.Y(n_1398)
);

AND2x4_ASAP7_75t_L g1399 ( 
.A(n_1304),
.B(n_1173),
.Y(n_1399)
);

INVx2_ASAP7_75t_L g1400 ( 
.A(n_1189),
.Y(n_1400)
);

INVx1_ASAP7_75t_L g1401 ( 
.A(n_1189),
.Y(n_1401)
);

OAI21x1_ASAP7_75t_L g1402 ( 
.A1(n_1295),
.A2(n_1200),
.B(n_1179),
.Y(n_1402)
);

AOI22xp33_ASAP7_75t_L g1403 ( 
.A1(n_1288),
.A2(n_1302),
.B1(n_1306),
.B2(n_860),
.Y(n_1403)
);

INVx2_ASAP7_75t_SL g1404 ( 
.A(n_1198),
.Y(n_1404)
);

INVx3_ASAP7_75t_L g1405 ( 
.A(n_1184),
.Y(n_1405)
);

AOI21xp5_ASAP7_75t_L g1406 ( 
.A1(n_1196),
.A2(n_1276),
.B(n_1272),
.Y(n_1406)
);

AOI22xp33_ASAP7_75t_L g1407 ( 
.A1(n_1302),
.A2(n_1306),
.B1(n_860),
.B2(n_1240),
.Y(n_1407)
);

OAI21x1_ASAP7_75t_L g1408 ( 
.A1(n_1273),
.A2(n_1279),
.B(n_1277),
.Y(n_1408)
);

INVx1_ASAP7_75t_L g1409 ( 
.A(n_1194),
.Y(n_1409)
);

INVxp67_ASAP7_75t_SL g1410 ( 
.A(n_1259),
.Y(n_1410)
);

INVx1_ASAP7_75t_L g1411 ( 
.A(n_1194),
.Y(n_1411)
);

NOR2xp33_ASAP7_75t_L g1412 ( 
.A(n_1302),
.B(n_1306),
.Y(n_1412)
);

OAI21x1_ASAP7_75t_L g1413 ( 
.A1(n_1273),
.A2(n_1279),
.B(n_1277),
.Y(n_1413)
);

OAI22xp5_ASAP7_75t_L g1414 ( 
.A1(n_1302),
.A2(n_915),
.B1(n_1265),
.B2(n_1262),
.Y(n_1414)
);

INVx1_ASAP7_75t_L g1415 ( 
.A(n_1194),
.Y(n_1415)
);

INVx1_ASAP7_75t_L g1416 ( 
.A(n_1194),
.Y(n_1416)
);

INVx1_ASAP7_75t_L g1417 ( 
.A(n_1194),
.Y(n_1417)
);

OAI21x1_ASAP7_75t_L g1418 ( 
.A1(n_1273),
.A2(n_1279),
.B(n_1277),
.Y(n_1418)
);

OAI22xp5_ASAP7_75t_L g1419 ( 
.A1(n_1302),
.A2(n_915),
.B1(n_1265),
.B2(n_1262),
.Y(n_1419)
);

INVx2_ASAP7_75t_L g1420 ( 
.A(n_1194),
.Y(n_1420)
);

NAND2xp5_ASAP7_75t_SL g1421 ( 
.A(n_1306),
.B(n_1300),
.Y(n_1421)
);

NAND2xp5_ASAP7_75t_SL g1422 ( 
.A(n_1306),
.B(n_1300),
.Y(n_1422)
);

OAI21x1_ASAP7_75t_L g1423 ( 
.A1(n_1273),
.A2(n_1279),
.B(n_1277),
.Y(n_1423)
);

O2A1O1Ixp33_ASAP7_75t_SL g1424 ( 
.A1(n_1172),
.A2(n_1300),
.B(n_1308),
.C(n_1306),
.Y(n_1424)
);

BUFx2_ASAP7_75t_L g1425 ( 
.A(n_1170),
.Y(n_1425)
);

INVx1_ASAP7_75t_L g1426 ( 
.A(n_1194),
.Y(n_1426)
);

AND2x2_ASAP7_75t_L g1427 ( 
.A(n_1292),
.B(n_915),
.Y(n_1427)
);

BUFx12f_ASAP7_75t_L g1428 ( 
.A(n_1192),
.Y(n_1428)
);

HB1xp67_ASAP7_75t_L g1429 ( 
.A(n_1190),
.Y(n_1429)
);

INVx1_ASAP7_75t_L g1430 ( 
.A(n_1194),
.Y(n_1430)
);

AO31x2_ASAP7_75t_L g1431 ( 
.A1(n_1168),
.A2(n_1223),
.A3(n_1197),
.B(n_1209),
.Y(n_1431)
);

BUFx2_ASAP7_75t_L g1432 ( 
.A(n_1170),
.Y(n_1432)
);

OAI21x1_ASAP7_75t_SL g1433 ( 
.A1(n_1246),
.A2(n_1203),
.B(n_1226),
.Y(n_1433)
);

INVx1_ASAP7_75t_L g1434 ( 
.A(n_1194),
.Y(n_1434)
);

CKINVDCx20_ASAP7_75t_R g1435 ( 
.A(n_1192),
.Y(n_1435)
);

OAI21x1_ASAP7_75t_L g1436 ( 
.A1(n_1273),
.A2(n_1279),
.B(n_1277),
.Y(n_1436)
);

AOI22xp33_ASAP7_75t_L g1437 ( 
.A1(n_1302),
.A2(n_1306),
.B1(n_860),
.B2(n_1240),
.Y(n_1437)
);

OAI21x1_ASAP7_75t_L g1438 ( 
.A1(n_1273),
.A2(n_1279),
.B(n_1277),
.Y(n_1438)
);

OAI21x1_ASAP7_75t_L g1439 ( 
.A1(n_1273),
.A2(n_1279),
.B(n_1277),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_1194),
.Y(n_1440)
);

INVx1_ASAP7_75t_L g1441 ( 
.A(n_1194),
.Y(n_1441)
);

INVx1_ASAP7_75t_SL g1442 ( 
.A(n_1270),
.Y(n_1442)
);

OAI21xp5_ASAP7_75t_L g1443 ( 
.A1(n_1300),
.A2(n_1308),
.B(n_1306),
.Y(n_1443)
);

A2O1A1Ixp33_ASAP7_75t_L g1444 ( 
.A1(n_1302),
.A2(n_1308),
.B(n_1300),
.C(n_1110),
.Y(n_1444)
);

O2A1O1Ixp33_ASAP7_75t_L g1445 ( 
.A1(n_1306),
.A2(n_1300),
.B(n_1308),
.C(n_1302),
.Y(n_1445)
);

OAI21xp5_ASAP7_75t_L g1446 ( 
.A1(n_1300),
.A2(n_1308),
.B(n_1306),
.Y(n_1446)
);

AO31x2_ASAP7_75t_L g1447 ( 
.A1(n_1168),
.A2(n_1223),
.A3(n_1197),
.B(n_1209),
.Y(n_1447)
);

OAI21x1_ASAP7_75t_L g1448 ( 
.A1(n_1273),
.A2(n_1279),
.B(n_1277),
.Y(n_1448)
);

OAI21x1_ASAP7_75t_L g1449 ( 
.A1(n_1273),
.A2(n_1279),
.B(n_1277),
.Y(n_1449)
);

INVx1_ASAP7_75t_L g1450 ( 
.A(n_1194),
.Y(n_1450)
);

INVx5_ASAP7_75t_L g1451 ( 
.A(n_1184),
.Y(n_1451)
);

OAI21xp5_ASAP7_75t_L g1452 ( 
.A1(n_1300),
.A2(n_1308),
.B(n_1306),
.Y(n_1452)
);

OR2x6_ASAP7_75t_L g1453 ( 
.A(n_1225),
.B(n_1244),
.Y(n_1453)
);

AND2x2_ASAP7_75t_L g1454 ( 
.A(n_1292),
.B(n_915),
.Y(n_1454)
);

NOR2xp67_ASAP7_75t_R g1455 ( 
.A(n_1451),
.B(n_1428),
.Y(n_1455)
);

OAI22xp5_ASAP7_75t_L g1456 ( 
.A1(n_1407),
.A2(n_1437),
.B1(n_1403),
.B2(n_1412),
.Y(n_1456)
);

OAI22xp5_ASAP7_75t_L g1457 ( 
.A1(n_1407),
.A2(n_1437),
.B1(n_1403),
.B2(n_1412),
.Y(n_1457)
);

OA21x2_ASAP7_75t_L g1458 ( 
.A1(n_1356),
.A2(n_1338),
.B(n_1443),
.Y(n_1458)
);

AOI21xp5_ASAP7_75t_L g1459 ( 
.A1(n_1331),
.A2(n_1453),
.B(n_1406),
.Y(n_1459)
);

BUFx3_ASAP7_75t_L g1460 ( 
.A(n_1314),
.Y(n_1460)
);

NAND2x1p5_ASAP7_75t_L g1461 ( 
.A(n_1451),
.B(n_1380),
.Y(n_1461)
);

NOR2x1_ASAP7_75t_SL g1462 ( 
.A(n_1453),
.B(n_1451),
.Y(n_1462)
);

AND2x2_ASAP7_75t_L g1463 ( 
.A(n_1317),
.B(n_1364),
.Y(n_1463)
);

AND2x2_ASAP7_75t_L g1464 ( 
.A(n_1312),
.B(n_1371),
.Y(n_1464)
);

OA21x2_ASAP7_75t_L g1465 ( 
.A1(n_1446),
.A2(n_1452),
.B(n_1336),
.Y(n_1465)
);

AND2x2_ASAP7_75t_L g1466 ( 
.A(n_1368),
.B(n_1427),
.Y(n_1466)
);

NOR2xp67_ASAP7_75t_L g1467 ( 
.A(n_1393),
.B(n_1359),
.Y(n_1467)
);

NAND2xp5_ASAP7_75t_L g1468 ( 
.A(n_1410),
.B(n_1349),
.Y(n_1468)
);

NAND2xp5_ASAP7_75t_L g1469 ( 
.A(n_1349),
.B(n_1429),
.Y(n_1469)
);

OAI22xp5_ASAP7_75t_L g1470 ( 
.A1(n_1322),
.A2(n_1444),
.B1(n_1453),
.B2(n_1381),
.Y(n_1470)
);

AND2x2_ASAP7_75t_L g1471 ( 
.A(n_1454),
.B(n_1315),
.Y(n_1471)
);

CKINVDCx20_ASAP7_75t_R g1472 ( 
.A(n_1339),
.Y(n_1472)
);

AND2x2_ASAP7_75t_L g1473 ( 
.A(n_1377),
.B(n_1414),
.Y(n_1473)
);

OAI22x1_ASAP7_75t_L g1474 ( 
.A1(n_1421),
.A2(n_1422),
.B1(n_1429),
.B2(n_1389),
.Y(n_1474)
);

INVx1_ASAP7_75t_L g1475 ( 
.A(n_1327),
.Y(n_1475)
);

NAND2xp5_ASAP7_75t_L g1476 ( 
.A(n_1329),
.B(n_1445),
.Y(n_1476)
);

HB1xp67_ASAP7_75t_L g1477 ( 
.A(n_1316),
.Y(n_1477)
);

OA22x2_ASAP7_75t_L g1478 ( 
.A1(n_1419),
.A2(n_1332),
.B1(n_1421),
.B2(n_1422),
.Y(n_1478)
);

CKINVDCx5p33_ASAP7_75t_R g1479 ( 
.A(n_1335),
.Y(n_1479)
);

AOI21xp5_ASAP7_75t_L g1480 ( 
.A1(n_1326),
.A2(n_1344),
.B(n_1444),
.Y(n_1480)
);

AND2x2_ASAP7_75t_L g1481 ( 
.A(n_1361),
.B(n_1386),
.Y(n_1481)
);

AND2x2_ASAP7_75t_L g1482 ( 
.A(n_1386),
.B(n_1318),
.Y(n_1482)
);

AOI21xp5_ASAP7_75t_L g1483 ( 
.A1(n_1344),
.A2(n_1323),
.B(n_1424),
.Y(n_1483)
);

OR2x2_ASAP7_75t_L g1484 ( 
.A(n_1442),
.B(n_1319),
.Y(n_1484)
);

NAND2xp33_ASAP7_75t_SL g1485 ( 
.A(n_1339),
.B(n_1435),
.Y(n_1485)
);

AOI21xp5_ASAP7_75t_L g1486 ( 
.A1(n_1323),
.A2(n_1424),
.B(n_1328),
.Y(n_1486)
);

NAND2xp5_ASAP7_75t_L g1487 ( 
.A(n_1347),
.B(n_1354),
.Y(n_1487)
);

NAND2xp5_ASAP7_75t_L g1488 ( 
.A(n_1385),
.B(n_1369),
.Y(n_1488)
);

OA21x2_ASAP7_75t_L g1489 ( 
.A1(n_1336),
.A2(n_1337),
.B(n_1346),
.Y(n_1489)
);

AOI21xp5_ASAP7_75t_L g1490 ( 
.A1(n_1357),
.A2(n_1382),
.B(n_1433),
.Y(n_1490)
);

OA21x2_ASAP7_75t_L g1491 ( 
.A1(n_1337),
.A2(n_1346),
.B(n_1350),
.Y(n_1491)
);

CKINVDCx5p33_ASAP7_75t_R g1492 ( 
.A(n_1428),
.Y(n_1492)
);

OR2x2_ASAP7_75t_L g1493 ( 
.A(n_1320),
.B(n_1321),
.Y(n_1493)
);

NOR2xp67_ASAP7_75t_L g1494 ( 
.A(n_1404),
.B(n_1343),
.Y(n_1494)
);

AND2x4_ASAP7_75t_L g1495 ( 
.A(n_1405),
.B(n_1396),
.Y(n_1495)
);

AOI21xp5_ASAP7_75t_L g1496 ( 
.A1(n_1360),
.A2(n_1358),
.B(n_1330),
.Y(n_1496)
);

O2A1O1Ixp33_ASAP7_75t_L g1497 ( 
.A1(n_1374),
.A2(n_1343),
.B(n_1372),
.C(n_1353),
.Y(n_1497)
);

O2A1O1Ixp33_ASAP7_75t_L g1498 ( 
.A1(n_1372),
.A2(n_1353),
.B(n_1379),
.C(n_1355),
.Y(n_1498)
);

NAND2xp5_ASAP7_75t_L g1499 ( 
.A(n_1370),
.B(n_1379),
.Y(n_1499)
);

OAI22xp5_ASAP7_75t_L g1500 ( 
.A1(n_1340),
.A2(n_1351),
.B1(n_1348),
.B2(n_1342),
.Y(n_1500)
);

AOI21xp5_ASAP7_75t_SL g1501 ( 
.A1(n_1352),
.A2(n_1366),
.B(n_1363),
.Y(n_1501)
);

O2A1O1Ixp5_ASAP7_75t_L g1502 ( 
.A1(n_1384),
.A2(n_1376),
.B(n_1375),
.C(n_1401),
.Y(n_1502)
);

OAI22xp5_ASAP7_75t_SL g1503 ( 
.A1(n_1435),
.A2(n_1314),
.B1(n_1313),
.B2(n_1425),
.Y(n_1503)
);

CKINVDCx5p33_ASAP7_75t_R g1504 ( 
.A(n_1313),
.Y(n_1504)
);

NAND2xp5_ASAP7_75t_L g1505 ( 
.A(n_1370),
.B(n_1341),
.Y(n_1505)
);

AOI21xp5_ASAP7_75t_L g1506 ( 
.A1(n_1360),
.A2(n_1451),
.B(n_1365),
.Y(n_1506)
);

O2A1O1Ixp5_ASAP7_75t_L g1507 ( 
.A1(n_1375),
.A2(n_1376),
.B(n_1398),
.C(n_1400),
.Y(n_1507)
);

NAND2xp5_ASAP7_75t_L g1508 ( 
.A(n_1370),
.B(n_1420),
.Y(n_1508)
);

O2A1O1Ixp33_ASAP7_75t_L g1509 ( 
.A1(n_1324),
.A2(n_1450),
.B(n_1441),
.C(n_1440),
.Y(n_1509)
);

NAND2xp5_ASAP7_75t_L g1510 ( 
.A(n_1370),
.B(n_1416),
.Y(n_1510)
);

CKINVDCx5p33_ASAP7_75t_R g1511 ( 
.A(n_1432),
.Y(n_1511)
);

OA21x2_ASAP7_75t_L g1512 ( 
.A1(n_1394),
.A2(n_1397),
.B(n_1395),
.Y(n_1512)
);

NAND2xp5_ASAP7_75t_L g1513 ( 
.A(n_1370),
.B(n_1415),
.Y(n_1513)
);

AND2x2_ASAP7_75t_L g1514 ( 
.A(n_1409),
.B(n_1417),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_1411),
.Y(n_1515)
);

NAND2xp5_ASAP7_75t_L g1516 ( 
.A(n_1426),
.B(n_1430),
.Y(n_1516)
);

OAI22xp5_ASAP7_75t_L g1517 ( 
.A1(n_1434),
.A2(n_1366),
.B1(n_1352),
.B2(n_1400),
.Y(n_1517)
);

OAI22xp5_ASAP7_75t_L g1518 ( 
.A1(n_1398),
.A2(n_1405),
.B1(n_1390),
.B2(n_1363),
.Y(n_1518)
);

NOR2xp67_ASAP7_75t_L g1519 ( 
.A(n_1399),
.B(n_1373),
.Y(n_1519)
);

AOI21x1_ASAP7_75t_SL g1520 ( 
.A1(n_1402),
.A2(n_1365),
.B(n_1362),
.Y(n_1520)
);

AND2x2_ASAP7_75t_L g1521 ( 
.A(n_1402),
.B(n_1392),
.Y(n_1521)
);

OAI22xp5_ASAP7_75t_L g1522 ( 
.A1(n_1383),
.A2(n_1387),
.B1(n_1392),
.B2(n_1367),
.Y(n_1522)
);

BUFx2_ASAP7_75t_L g1523 ( 
.A(n_1388),
.Y(n_1523)
);

AND2x2_ASAP7_75t_L g1524 ( 
.A(n_1383),
.B(n_1387),
.Y(n_1524)
);

INVx8_ASAP7_75t_L g1525 ( 
.A(n_1391),
.Y(n_1525)
);

OA21x2_ASAP7_75t_L g1526 ( 
.A1(n_1397),
.A2(n_1362),
.B(n_1345),
.Y(n_1526)
);

CKINVDCx5p33_ASAP7_75t_R g1527 ( 
.A(n_1325),
.Y(n_1527)
);

AND2x2_ASAP7_75t_L g1528 ( 
.A(n_1325),
.B(n_1431),
.Y(n_1528)
);

AND2x2_ASAP7_75t_L g1529 ( 
.A(n_1325),
.B(n_1431),
.Y(n_1529)
);

OA21x2_ASAP7_75t_L g1530 ( 
.A1(n_1345),
.A2(n_1378),
.B(n_1448),
.Y(n_1530)
);

O2A1O1Ixp33_ASAP7_75t_L g1531 ( 
.A1(n_1447),
.A2(n_1436),
.B(n_1438),
.C(n_1423),
.Y(n_1531)
);

HB1xp67_ASAP7_75t_L g1532 ( 
.A(n_1408),
.Y(n_1532)
);

INVx3_ASAP7_75t_L g1533 ( 
.A(n_1408),
.Y(n_1533)
);

AND2x4_ASAP7_75t_SL g1534 ( 
.A(n_1413),
.B(n_1418),
.Y(n_1534)
);

O2A1O1Ixp33_ASAP7_75t_L g1535 ( 
.A1(n_1413),
.A2(n_1418),
.B(n_1439),
.C(n_1448),
.Y(n_1535)
);

OR2x2_ASAP7_75t_L g1536 ( 
.A(n_1439),
.B(n_1449),
.Y(n_1536)
);

AOI21xp5_ASAP7_75t_L g1537 ( 
.A1(n_1449),
.A2(n_1331),
.B(n_1196),
.Y(n_1537)
);

BUFx2_ASAP7_75t_L g1538 ( 
.A(n_1361),
.Y(n_1538)
);

OR2x2_ASAP7_75t_L g1539 ( 
.A(n_1333),
.B(n_1317),
.Y(n_1539)
);

AND2x2_ASAP7_75t_L g1540 ( 
.A(n_1317),
.B(n_1364),
.Y(n_1540)
);

OA21x2_ASAP7_75t_L g1541 ( 
.A1(n_1356),
.A2(n_1338),
.B(n_1443),
.Y(n_1541)
);

AND2x2_ASAP7_75t_L g1542 ( 
.A(n_1317),
.B(n_1364),
.Y(n_1542)
);

AND2x2_ASAP7_75t_L g1543 ( 
.A(n_1317),
.B(n_1364),
.Y(n_1543)
);

OR2x2_ASAP7_75t_L g1544 ( 
.A(n_1333),
.B(n_1317),
.Y(n_1544)
);

OAI22xp5_ASAP7_75t_SL g1545 ( 
.A1(n_1403),
.A2(n_1302),
.B1(n_1412),
.B2(n_1057),
.Y(n_1545)
);

AND2x2_ASAP7_75t_SL g1546 ( 
.A(n_1407),
.B(n_1254),
.Y(n_1546)
);

AND2x4_ASAP7_75t_L g1547 ( 
.A(n_1334),
.B(n_1361),
.Y(n_1547)
);

OAI22xp5_ASAP7_75t_L g1548 ( 
.A1(n_1407),
.A2(n_1302),
.B1(n_1437),
.B2(n_1311),
.Y(n_1548)
);

AOI21xp5_ASAP7_75t_SL g1549 ( 
.A1(n_1453),
.A2(n_621),
.B(n_619),
.Y(n_1549)
);

O2A1O1Ixp33_ASAP7_75t_L g1550 ( 
.A1(n_1412),
.A2(n_1306),
.B(n_1308),
.C(n_1300),
.Y(n_1550)
);

O2A1O1Ixp33_ASAP7_75t_L g1551 ( 
.A1(n_1412),
.A2(n_1306),
.B(n_1308),
.C(n_1300),
.Y(n_1551)
);

BUFx3_ASAP7_75t_L g1552 ( 
.A(n_1314),
.Y(n_1552)
);

AND2x2_ASAP7_75t_L g1553 ( 
.A(n_1317),
.B(n_1364),
.Y(n_1553)
);

OAI22xp5_ASAP7_75t_L g1554 ( 
.A1(n_1407),
.A2(n_1302),
.B1(n_1437),
.B2(n_1311),
.Y(n_1554)
);

BUFx2_ASAP7_75t_L g1555 ( 
.A(n_1512),
.Y(n_1555)
);

AO21x2_ASAP7_75t_L g1556 ( 
.A1(n_1480),
.A2(n_1496),
.B(n_1506),
.Y(n_1556)
);

BUFx3_ASAP7_75t_L g1557 ( 
.A(n_1525),
.Y(n_1557)
);

INVx2_ASAP7_75t_L g1558 ( 
.A(n_1512),
.Y(n_1558)
);

INVx1_ASAP7_75t_L g1559 ( 
.A(n_1507),
.Y(n_1559)
);

HB1xp67_ASAP7_75t_L g1560 ( 
.A(n_1522),
.Y(n_1560)
);

AND2x2_ASAP7_75t_L g1561 ( 
.A(n_1524),
.B(n_1528),
.Y(n_1561)
);

HB1xp67_ASAP7_75t_L g1562 ( 
.A(n_1522),
.Y(n_1562)
);

AO21x2_ASAP7_75t_L g1563 ( 
.A1(n_1537),
.A2(n_1459),
.B(n_1490),
.Y(n_1563)
);

AND2x4_ASAP7_75t_L g1564 ( 
.A(n_1533),
.B(n_1534),
.Y(n_1564)
);

NAND2xp5_ASAP7_75t_L g1565 ( 
.A(n_1469),
.B(n_1468),
.Y(n_1565)
);

INVx2_ASAP7_75t_L g1566 ( 
.A(n_1536),
.Y(n_1566)
);

INVx2_ASAP7_75t_L g1567 ( 
.A(n_1526),
.Y(n_1567)
);

AND2x2_ASAP7_75t_L g1568 ( 
.A(n_1529),
.B(n_1465),
.Y(n_1568)
);

AND2x2_ASAP7_75t_L g1569 ( 
.A(n_1465),
.B(n_1527),
.Y(n_1569)
);

HB1xp67_ASAP7_75t_L g1570 ( 
.A(n_1469),
.Y(n_1570)
);

INVx1_ASAP7_75t_L g1571 ( 
.A(n_1502),
.Y(n_1571)
);

AO21x2_ASAP7_75t_L g1572 ( 
.A1(n_1483),
.A2(n_1476),
.B(n_1486),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_1532),
.Y(n_1573)
);

INVx2_ASAP7_75t_L g1574 ( 
.A(n_1530),
.Y(n_1574)
);

INVx2_ASAP7_75t_L g1575 ( 
.A(n_1530),
.Y(n_1575)
);

OR2x2_ASAP7_75t_L g1576 ( 
.A(n_1458),
.B(n_1541),
.Y(n_1576)
);

AND2x2_ASAP7_75t_L g1577 ( 
.A(n_1458),
.B(n_1541),
.Y(n_1577)
);

AND2x2_ASAP7_75t_L g1578 ( 
.A(n_1473),
.B(n_1491),
.Y(n_1578)
);

OR2x2_ASAP7_75t_L g1579 ( 
.A(n_1468),
.B(n_1491),
.Y(n_1579)
);

AOI22xp33_ASAP7_75t_L g1580 ( 
.A1(n_1546),
.A2(n_1548),
.B1(n_1554),
.B2(n_1457),
.Y(n_1580)
);

AND2x2_ASAP7_75t_L g1581 ( 
.A(n_1489),
.B(n_1505),
.Y(n_1581)
);

OR2x2_ASAP7_75t_L g1582 ( 
.A(n_1489),
.B(n_1505),
.Y(n_1582)
);

NAND2xp5_ASAP7_75t_L g1583 ( 
.A(n_1487),
.B(n_1476),
.Y(n_1583)
);

AND2x2_ASAP7_75t_L g1584 ( 
.A(n_1508),
.B(n_1463),
.Y(n_1584)
);

BUFx3_ASAP7_75t_L g1585 ( 
.A(n_1521),
.Y(n_1585)
);

OA21x2_ASAP7_75t_L g1586 ( 
.A1(n_1486),
.A2(n_1499),
.B(n_1487),
.Y(n_1586)
);

OR2x6_ASAP7_75t_L g1587 ( 
.A(n_1461),
.B(n_1531),
.Y(n_1587)
);

OA21x2_ASAP7_75t_L g1588 ( 
.A1(n_1499),
.A2(n_1513),
.B(n_1510),
.Y(n_1588)
);

AND2x2_ASAP7_75t_L g1589 ( 
.A(n_1508),
.B(n_1523),
.Y(n_1589)
);

OAI21x1_ASAP7_75t_L g1590 ( 
.A1(n_1520),
.A2(n_1535),
.B(n_1461),
.Y(n_1590)
);

AOI21xp5_ASAP7_75t_SL g1591 ( 
.A1(n_1550),
.A2(n_1551),
.B(n_1548),
.Y(n_1591)
);

INVx2_ASAP7_75t_L g1592 ( 
.A(n_1475),
.Y(n_1592)
);

CKINVDCx11_ASAP7_75t_R g1593 ( 
.A(n_1472),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_1500),
.Y(n_1594)
);

NOR2xp33_ASAP7_75t_L g1595 ( 
.A(n_1456),
.B(n_1457),
.Y(n_1595)
);

AOI22xp5_ASAP7_75t_L g1596 ( 
.A1(n_1554),
.A2(n_1456),
.B1(n_1545),
.B2(n_1478),
.Y(n_1596)
);

AND2x2_ASAP7_75t_L g1597 ( 
.A(n_1540),
.B(n_1553),
.Y(n_1597)
);

OA21x2_ASAP7_75t_L g1598 ( 
.A1(n_1488),
.A2(n_1515),
.B(n_1470),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1500),
.Y(n_1599)
);

AO21x2_ASAP7_75t_L g1600 ( 
.A1(n_1517),
.A2(n_1518),
.B(n_1470),
.Y(n_1600)
);

NOR2xp33_ASAP7_75t_L g1601 ( 
.A(n_1478),
.B(n_1544),
.Y(n_1601)
);

AND2x2_ASAP7_75t_L g1602 ( 
.A(n_1542),
.B(n_1543),
.Y(n_1602)
);

OR2x2_ASAP7_75t_L g1603 ( 
.A(n_1539),
.B(n_1474),
.Y(n_1603)
);

AOI22xp33_ASAP7_75t_L g1604 ( 
.A1(n_1464),
.A2(n_1477),
.B1(n_1485),
.B2(n_1471),
.Y(n_1604)
);

HB1xp67_ASAP7_75t_L g1605 ( 
.A(n_1519),
.Y(n_1605)
);

INVx1_ASAP7_75t_L g1606 ( 
.A(n_1592),
.Y(n_1606)
);

AND2x2_ASAP7_75t_L g1607 ( 
.A(n_1561),
.B(n_1578),
.Y(n_1607)
);

AND2x2_ASAP7_75t_L g1608 ( 
.A(n_1561),
.B(n_1482),
.Y(n_1608)
);

INVx2_ASAP7_75t_R g1609 ( 
.A(n_1571),
.Y(n_1609)
);

AND2x4_ASAP7_75t_L g1610 ( 
.A(n_1557),
.B(n_1462),
.Y(n_1610)
);

OR2x2_ASAP7_75t_L g1611 ( 
.A(n_1588),
.B(n_1484),
.Y(n_1611)
);

INVx1_ASAP7_75t_L g1612 ( 
.A(n_1592),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1592),
.Y(n_1613)
);

AOI22xp33_ASAP7_75t_L g1614 ( 
.A1(n_1595),
.A2(n_1466),
.B1(n_1503),
.B2(n_1481),
.Y(n_1614)
);

NAND2xp33_ASAP7_75t_R g1615 ( 
.A(n_1588),
.B(n_1492),
.Y(n_1615)
);

NOR2xp67_ASAP7_75t_L g1616 ( 
.A(n_1566),
.B(n_1516),
.Y(n_1616)
);

OR2x2_ASAP7_75t_L g1617 ( 
.A(n_1588),
.B(n_1493),
.Y(n_1617)
);

INVxp67_ASAP7_75t_L g1618 ( 
.A(n_1570),
.Y(n_1618)
);

CKINVDCx20_ASAP7_75t_R g1619 ( 
.A(n_1593),
.Y(n_1619)
);

BUFx2_ASAP7_75t_L g1620 ( 
.A(n_1564),
.Y(n_1620)
);

AND2x6_ASAP7_75t_SL g1621 ( 
.A(n_1595),
.B(n_1455),
.Y(n_1621)
);

HB1xp67_ASAP7_75t_L g1622 ( 
.A(n_1588),
.Y(n_1622)
);

AOI221xp5_ASAP7_75t_L g1623 ( 
.A1(n_1591),
.A2(n_1497),
.B1(n_1498),
.B2(n_1509),
.C(n_1514),
.Y(n_1623)
);

NAND2xp5_ASAP7_75t_L g1624 ( 
.A(n_1565),
.B(n_1516),
.Y(n_1624)
);

HB1xp67_ASAP7_75t_L g1625 ( 
.A(n_1588),
.Y(n_1625)
);

NAND2x1p5_ASAP7_75t_L g1626 ( 
.A(n_1598),
.B(n_1494),
.Y(n_1626)
);

AO21x2_ASAP7_75t_L g1627 ( 
.A1(n_1556),
.A2(n_1549),
.B(n_1501),
.Y(n_1627)
);

NOR2xp33_ASAP7_75t_L g1628 ( 
.A(n_1593),
.B(n_1511),
.Y(n_1628)
);

AND2x2_ASAP7_75t_L g1629 ( 
.A(n_1561),
.B(n_1547),
.Y(n_1629)
);

HB1xp67_ASAP7_75t_L g1630 ( 
.A(n_1588),
.Y(n_1630)
);

INVx1_ASAP7_75t_SL g1631 ( 
.A(n_1581),
.Y(n_1631)
);

HB1xp67_ASAP7_75t_L g1632 ( 
.A(n_1589),
.Y(n_1632)
);

OA21x2_ASAP7_75t_L g1633 ( 
.A1(n_1574),
.A2(n_1538),
.B(n_1495),
.Y(n_1633)
);

NOR2xp33_ASAP7_75t_L g1634 ( 
.A(n_1583),
.B(n_1504),
.Y(n_1634)
);

OR2x6_ASAP7_75t_L g1635 ( 
.A(n_1587),
.B(n_1547),
.Y(n_1635)
);

INVx2_ASAP7_75t_SL g1636 ( 
.A(n_1605),
.Y(n_1636)
);

INVx3_ASAP7_75t_L g1637 ( 
.A(n_1564),
.Y(n_1637)
);

NAND2xp5_ASAP7_75t_L g1638 ( 
.A(n_1565),
.B(n_1583),
.Y(n_1638)
);

AND2x2_ASAP7_75t_L g1639 ( 
.A(n_1578),
.B(n_1585),
.Y(n_1639)
);

AOI22xp5_ASAP7_75t_SL g1640 ( 
.A1(n_1619),
.A2(n_1601),
.B1(n_1479),
.B2(n_1605),
.Y(n_1640)
);

INVx1_ASAP7_75t_L g1641 ( 
.A(n_1606),
.Y(n_1641)
);

AND2x2_ASAP7_75t_L g1642 ( 
.A(n_1607),
.B(n_1578),
.Y(n_1642)
);

AND2x2_ASAP7_75t_L g1643 ( 
.A(n_1607),
.B(n_1585),
.Y(n_1643)
);

AND2x6_ASAP7_75t_SL g1644 ( 
.A(n_1628),
.B(n_1601),
.Y(n_1644)
);

AND2x4_ASAP7_75t_L g1645 ( 
.A(n_1635),
.B(n_1585),
.Y(n_1645)
);

INVx1_ASAP7_75t_L g1646 ( 
.A(n_1606),
.Y(n_1646)
);

BUFx2_ASAP7_75t_L g1647 ( 
.A(n_1620),
.Y(n_1647)
);

AND2x2_ASAP7_75t_L g1648 ( 
.A(n_1639),
.B(n_1585),
.Y(n_1648)
);

NAND2xp33_ASAP7_75t_R g1649 ( 
.A(n_1610),
.B(n_1603),
.Y(n_1649)
);

AND2x4_ASAP7_75t_L g1650 ( 
.A(n_1635),
.B(n_1637),
.Y(n_1650)
);

AND2x2_ASAP7_75t_L g1651 ( 
.A(n_1639),
.B(n_1569),
.Y(n_1651)
);

HB1xp67_ASAP7_75t_L g1652 ( 
.A(n_1616),
.Y(n_1652)
);

OAI21x1_ASAP7_75t_L g1653 ( 
.A1(n_1626),
.A2(n_1590),
.B(n_1558),
.Y(n_1653)
);

AOI22xp5_ASAP7_75t_L g1654 ( 
.A1(n_1623),
.A2(n_1596),
.B1(n_1580),
.B2(n_1600),
.Y(n_1654)
);

AND2x2_ASAP7_75t_L g1655 ( 
.A(n_1632),
.B(n_1569),
.Y(n_1655)
);

AOI222xp33_ASAP7_75t_L g1656 ( 
.A1(n_1614),
.A2(n_1580),
.B1(n_1596),
.B2(n_1569),
.C1(n_1577),
.C2(n_1604),
.Y(n_1656)
);

INVxp67_ASAP7_75t_SL g1657 ( 
.A(n_1616),
.Y(n_1657)
);

AOI22xp33_ASAP7_75t_L g1658 ( 
.A1(n_1634),
.A2(n_1596),
.B1(n_1603),
.B2(n_1600),
.Y(n_1658)
);

NAND2x1_ASAP7_75t_L g1659 ( 
.A(n_1633),
.B(n_1635),
.Y(n_1659)
);

A2O1A1Ixp33_ASAP7_75t_L g1660 ( 
.A1(n_1622),
.A2(n_1603),
.B(n_1560),
.C(n_1562),
.Y(n_1660)
);

AOI221xp5_ASAP7_75t_L g1661 ( 
.A1(n_1638),
.A2(n_1560),
.B1(n_1562),
.B2(n_1577),
.C(n_1604),
.Y(n_1661)
);

NAND2xp5_ASAP7_75t_L g1662 ( 
.A(n_1638),
.B(n_1584),
.Y(n_1662)
);

AOI221xp5_ASAP7_75t_L g1663 ( 
.A1(n_1625),
.A2(n_1577),
.B1(n_1571),
.B2(n_1584),
.C(n_1597),
.Y(n_1663)
);

AOI22xp5_ASAP7_75t_L g1664 ( 
.A1(n_1615),
.A2(n_1600),
.B1(n_1572),
.B2(n_1563),
.Y(n_1664)
);

INVxp67_ASAP7_75t_SL g1665 ( 
.A(n_1626),
.Y(n_1665)
);

AO21x2_ASAP7_75t_L g1666 ( 
.A1(n_1630),
.A2(n_1571),
.B(n_1558),
.Y(n_1666)
);

AND2x6_ASAP7_75t_SL g1667 ( 
.A(n_1635),
.B(n_1597),
.Y(n_1667)
);

OR2x2_ASAP7_75t_L g1668 ( 
.A(n_1611),
.B(n_1579),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_1612),
.Y(n_1669)
);

NOR4xp25_ASAP7_75t_SL g1670 ( 
.A(n_1620),
.B(n_1555),
.C(n_1559),
.D(n_1573),
.Y(n_1670)
);

BUFx2_ASAP7_75t_L g1671 ( 
.A(n_1637),
.Y(n_1671)
);

AND2x2_ASAP7_75t_L g1672 ( 
.A(n_1631),
.B(n_1568),
.Y(n_1672)
);

AO21x2_ASAP7_75t_L g1673 ( 
.A1(n_1627),
.A2(n_1558),
.B(n_1567),
.Y(n_1673)
);

OAI221xp5_ASAP7_75t_L g1674 ( 
.A1(n_1626),
.A2(n_1576),
.B1(n_1467),
.B2(n_1582),
.C(n_1460),
.Y(n_1674)
);

OAI22xp5_ASAP7_75t_L g1675 ( 
.A1(n_1635),
.A2(n_1594),
.B1(n_1599),
.B2(n_1602),
.Y(n_1675)
);

INVxp67_ASAP7_75t_L g1676 ( 
.A(n_1608),
.Y(n_1676)
);

INVxp67_ASAP7_75t_SL g1677 ( 
.A(n_1611),
.Y(n_1677)
);

INVx1_ASAP7_75t_L g1678 ( 
.A(n_1613),
.Y(n_1678)
);

INVx1_ASAP7_75t_L g1679 ( 
.A(n_1641),
.Y(n_1679)
);

INVx1_ASAP7_75t_SL g1680 ( 
.A(n_1640),
.Y(n_1680)
);

OA21x2_ASAP7_75t_L g1681 ( 
.A1(n_1653),
.A2(n_1574),
.B(n_1575),
.Y(n_1681)
);

INVx1_ASAP7_75t_L g1682 ( 
.A(n_1641),
.Y(n_1682)
);

INVxp67_ASAP7_75t_L g1683 ( 
.A(n_1652),
.Y(n_1683)
);

INVx1_ASAP7_75t_L g1684 ( 
.A(n_1646),
.Y(n_1684)
);

AND2x2_ASAP7_75t_L g1685 ( 
.A(n_1671),
.B(n_1631),
.Y(n_1685)
);

INVx2_ASAP7_75t_L g1686 ( 
.A(n_1666),
.Y(n_1686)
);

NOR2xp33_ASAP7_75t_L g1687 ( 
.A(n_1644),
.B(n_1621),
.Y(n_1687)
);

INVx2_ASAP7_75t_L g1688 ( 
.A(n_1666),
.Y(n_1688)
);

INVx2_ASAP7_75t_L g1689 ( 
.A(n_1666),
.Y(n_1689)
);

AOI21xp5_ASAP7_75t_L g1690 ( 
.A1(n_1664),
.A2(n_1660),
.B(n_1654),
.Y(n_1690)
);

INVx2_ASAP7_75t_L g1691 ( 
.A(n_1673),
.Y(n_1691)
);

INVx1_ASAP7_75t_L g1692 ( 
.A(n_1646),
.Y(n_1692)
);

NAND2xp5_ASAP7_75t_L g1693 ( 
.A(n_1677),
.B(n_1618),
.Y(n_1693)
);

BUFx2_ASAP7_75t_L g1694 ( 
.A(n_1667),
.Y(n_1694)
);

INVx2_ASAP7_75t_L g1695 ( 
.A(n_1673),
.Y(n_1695)
);

INVx2_ASAP7_75t_L g1696 ( 
.A(n_1673),
.Y(n_1696)
);

INVx1_ASAP7_75t_L g1697 ( 
.A(n_1678),
.Y(n_1697)
);

AND2x2_ASAP7_75t_L g1698 ( 
.A(n_1671),
.B(n_1609),
.Y(n_1698)
);

AND2x2_ASAP7_75t_L g1699 ( 
.A(n_1647),
.B(n_1609),
.Y(n_1699)
);

INVx2_ASAP7_75t_SL g1700 ( 
.A(n_1659),
.Y(n_1700)
);

INVx1_ASAP7_75t_L g1701 ( 
.A(n_1678),
.Y(n_1701)
);

OAI21x1_ASAP7_75t_L g1702 ( 
.A1(n_1664),
.A2(n_1590),
.B(n_1575),
.Y(n_1702)
);

INVx1_ASAP7_75t_L g1703 ( 
.A(n_1669),
.Y(n_1703)
);

NAND3xp33_ASAP7_75t_SL g1704 ( 
.A(n_1656),
.B(n_1658),
.C(n_1670),
.Y(n_1704)
);

AND2x2_ASAP7_75t_L g1705 ( 
.A(n_1647),
.B(n_1609),
.Y(n_1705)
);

AND2x2_ASAP7_75t_L g1706 ( 
.A(n_1642),
.B(n_1672),
.Y(n_1706)
);

INVx2_ASAP7_75t_L g1707 ( 
.A(n_1681),
.Y(n_1707)
);

INVx2_ASAP7_75t_L g1708 ( 
.A(n_1681),
.Y(n_1708)
);

OR2x2_ASAP7_75t_L g1709 ( 
.A(n_1693),
.B(n_1668),
.Y(n_1709)
);

INVx1_ASAP7_75t_L g1710 ( 
.A(n_1679),
.Y(n_1710)
);

INVx3_ASAP7_75t_L g1711 ( 
.A(n_1681),
.Y(n_1711)
);

INVx4_ASAP7_75t_L g1712 ( 
.A(n_1694),
.Y(n_1712)
);

INVx1_ASAP7_75t_L g1713 ( 
.A(n_1679),
.Y(n_1713)
);

HB1xp67_ASAP7_75t_L g1714 ( 
.A(n_1683),
.Y(n_1714)
);

NAND2xp5_ASAP7_75t_L g1715 ( 
.A(n_1690),
.B(n_1663),
.Y(n_1715)
);

OR2x6_ASAP7_75t_L g1716 ( 
.A(n_1690),
.B(n_1587),
.Y(n_1716)
);

AND2x2_ASAP7_75t_L g1717 ( 
.A(n_1694),
.B(n_1651),
.Y(n_1717)
);

NOR3xp33_ASAP7_75t_L g1718 ( 
.A(n_1704),
.B(n_1674),
.C(n_1661),
.Y(n_1718)
);

AND2x2_ASAP7_75t_L g1719 ( 
.A(n_1694),
.B(n_1651),
.Y(n_1719)
);

AND2x2_ASAP7_75t_L g1720 ( 
.A(n_1706),
.B(n_1650),
.Y(n_1720)
);

INVxp67_ASAP7_75t_SL g1721 ( 
.A(n_1687),
.Y(n_1721)
);

INVx1_ASAP7_75t_L g1722 ( 
.A(n_1679),
.Y(n_1722)
);

NAND2xp5_ASAP7_75t_L g1723 ( 
.A(n_1683),
.B(n_1676),
.Y(n_1723)
);

AND2x2_ASAP7_75t_L g1724 ( 
.A(n_1706),
.B(n_1650),
.Y(n_1724)
);

OAI211xp5_ASAP7_75t_SL g1725 ( 
.A1(n_1687),
.A2(n_1668),
.B(n_1662),
.C(n_1665),
.Y(n_1725)
);

NAND2xp5_ASAP7_75t_L g1726 ( 
.A(n_1680),
.B(n_1608),
.Y(n_1726)
);

NOR2xp33_ASAP7_75t_L g1727 ( 
.A(n_1680),
.B(n_1552),
.Y(n_1727)
);

AND2x2_ASAP7_75t_L g1728 ( 
.A(n_1706),
.B(n_1650),
.Y(n_1728)
);

NAND2xp5_ASAP7_75t_L g1729 ( 
.A(n_1693),
.B(n_1657),
.Y(n_1729)
);

NAND2xp5_ASAP7_75t_L g1730 ( 
.A(n_1704),
.B(n_1655),
.Y(n_1730)
);

INVx2_ASAP7_75t_L g1731 ( 
.A(n_1681),
.Y(n_1731)
);

AOI221xp5_ASAP7_75t_L g1732 ( 
.A1(n_1682),
.A2(n_1675),
.B1(n_1624),
.B2(n_1577),
.C(n_1655),
.Y(n_1732)
);

INVx1_ASAP7_75t_SL g1733 ( 
.A(n_1699),
.Y(n_1733)
);

NAND4xp25_ASAP7_75t_SL g1734 ( 
.A(n_1699),
.B(n_1648),
.C(n_1643),
.D(n_1672),
.Y(n_1734)
);

INVx1_ASAP7_75t_L g1735 ( 
.A(n_1682),
.Y(n_1735)
);

NOR2xp33_ASAP7_75t_L g1736 ( 
.A(n_1685),
.B(n_1621),
.Y(n_1736)
);

INVx2_ASAP7_75t_L g1737 ( 
.A(n_1681),
.Y(n_1737)
);

NAND2x1_ASAP7_75t_SL g1738 ( 
.A(n_1699),
.B(n_1645),
.Y(n_1738)
);

HB1xp67_ASAP7_75t_L g1739 ( 
.A(n_1697),
.Y(n_1739)
);

INVx1_ASAP7_75t_L g1740 ( 
.A(n_1682),
.Y(n_1740)
);

AND2x2_ASAP7_75t_L g1741 ( 
.A(n_1685),
.B(n_1643),
.Y(n_1741)
);

AND2x2_ASAP7_75t_L g1742 ( 
.A(n_1685),
.B(n_1645),
.Y(n_1742)
);

AND2x2_ASAP7_75t_L g1743 ( 
.A(n_1705),
.B(n_1645),
.Y(n_1743)
);

NAND2xp5_ASAP7_75t_L g1744 ( 
.A(n_1697),
.B(n_1629),
.Y(n_1744)
);

NAND2xp5_ASAP7_75t_L g1745 ( 
.A(n_1701),
.B(n_1642),
.Y(n_1745)
);

INVx1_ASAP7_75t_L g1746 ( 
.A(n_1684),
.Y(n_1746)
);

INVx1_ASAP7_75t_L g1747 ( 
.A(n_1684),
.Y(n_1747)
);

INVx2_ASAP7_75t_L g1748 ( 
.A(n_1712),
.Y(n_1748)
);

INVx1_ASAP7_75t_L g1749 ( 
.A(n_1739),
.Y(n_1749)
);

INVx2_ASAP7_75t_SL g1750 ( 
.A(n_1738),
.Y(n_1750)
);

OR2x2_ASAP7_75t_L g1751 ( 
.A(n_1714),
.B(n_1684),
.Y(n_1751)
);

INVx2_ASAP7_75t_L g1752 ( 
.A(n_1712),
.Y(n_1752)
);

OR2x2_ASAP7_75t_L g1753 ( 
.A(n_1709),
.B(n_1692),
.Y(n_1753)
);

NAND2x1p5_ASAP7_75t_L g1754 ( 
.A(n_1712),
.B(n_1705),
.Y(n_1754)
);

NAND2xp5_ASAP7_75t_L g1755 ( 
.A(n_1721),
.B(n_1636),
.Y(n_1755)
);

OAI22xp33_ASAP7_75t_L g1756 ( 
.A1(n_1715),
.A2(n_1649),
.B1(n_1586),
.B2(n_1576),
.Y(n_1756)
);

NAND2x1p5_ASAP7_75t_L g1757 ( 
.A(n_1712),
.B(n_1717),
.Y(n_1757)
);

BUFx2_ASAP7_75t_L g1758 ( 
.A(n_1738),
.Y(n_1758)
);

INVx1_ASAP7_75t_SL g1759 ( 
.A(n_1717),
.Y(n_1759)
);

AND2x2_ASAP7_75t_L g1760 ( 
.A(n_1719),
.B(n_1705),
.Y(n_1760)
);

NOR2xp67_ASAP7_75t_L g1761 ( 
.A(n_1734),
.B(n_1700),
.Y(n_1761)
);

BUFx2_ASAP7_75t_L g1762 ( 
.A(n_1719),
.Y(n_1762)
);

INVx1_ASAP7_75t_L g1763 ( 
.A(n_1710),
.Y(n_1763)
);

AND2x2_ASAP7_75t_L g1764 ( 
.A(n_1720),
.B(n_1724),
.Y(n_1764)
);

OR2x2_ASAP7_75t_L g1765 ( 
.A(n_1709),
.B(n_1703),
.Y(n_1765)
);

INVx1_ASAP7_75t_L g1766 ( 
.A(n_1710),
.Y(n_1766)
);

INVx1_ASAP7_75t_L g1767 ( 
.A(n_1713),
.Y(n_1767)
);

AND2x2_ASAP7_75t_L g1768 ( 
.A(n_1720),
.B(n_1698),
.Y(n_1768)
);

OR2x2_ASAP7_75t_L g1769 ( 
.A(n_1723),
.B(n_1703),
.Y(n_1769)
);

OR2x2_ASAP7_75t_L g1770 ( 
.A(n_1726),
.B(n_1617),
.Y(n_1770)
);

O2A1O1Ixp33_ASAP7_75t_L g1771 ( 
.A1(n_1718),
.A2(n_1686),
.B(n_1688),
.C(n_1689),
.Y(n_1771)
);

INVx1_ASAP7_75t_L g1772 ( 
.A(n_1713),
.Y(n_1772)
);

INVx1_ASAP7_75t_L g1773 ( 
.A(n_1722),
.Y(n_1773)
);

BUFx2_ASAP7_75t_L g1774 ( 
.A(n_1741),
.Y(n_1774)
);

INVx1_ASAP7_75t_L g1775 ( 
.A(n_1722),
.Y(n_1775)
);

INVx1_ASAP7_75t_L g1776 ( 
.A(n_1735),
.Y(n_1776)
);

INVx1_ASAP7_75t_SL g1777 ( 
.A(n_1727),
.Y(n_1777)
);

AND2x2_ASAP7_75t_L g1778 ( 
.A(n_1724),
.B(n_1698),
.Y(n_1778)
);

OR2x2_ASAP7_75t_L g1779 ( 
.A(n_1723),
.B(n_1692),
.Y(n_1779)
);

OR2x2_ASAP7_75t_L g1780 ( 
.A(n_1745),
.B(n_1692),
.Y(n_1780)
);

INVxp67_ASAP7_75t_SL g1781 ( 
.A(n_1736),
.Y(n_1781)
);

INVxp67_ASAP7_75t_SL g1782 ( 
.A(n_1730),
.Y(n_1782)
);

NAND2xp5_ASAP7_75t_L g1783 ( 
.A(n_1715),
.B(n_1636),
.Y(n_1783)
);

AND2x2_ASAP7_75t_L g1784 ( 
.A(n_1758),
.B(n_1728),
.Y(n_1784)
);

INVxp67_ASAP7_75t_L g1785 ( 
.A(n_1762),
.Y(n_1785)
);

NAND2xp5_ASAP7_75t_L g1786 ( 
.A(n_1777),
.B(n_1741),
.Y(n_1786)
);

INVx3_ASAP7_75t_SL g1787 ( 
.A(n_1748),
.Y(n_1787)
);

AND2x2_ASAP7_75t_L g1788 ( 
.A(n_1764),
.B(n_1728),
.Y(n_1788)
);

NAND2xp5_ASAP7_75t_L g1789 ( 
.A(n_1781),
.B(n_1729),
.Y(n_1789)
);

AND2x2_ASAP7_75t_L g1790 ( 
.A(n_1764),
.B(n_1742),
.Y(n_1790)
);

INVx1_ASAP7_75t_L g1791 ( 
.A(n_1751),
.Y(n_1791)
);

AND2x4_ASAP7_75t_L g1792 ( 
.A(n_1750),
.B(n_1743),
.Y(n_1792)
);

NAND2xp5_ASAP7_75t_L g1793 ( 
.A(n_1782),
.B(n_1732),
.Y(n_1793)
);

NAND2xp5_ASAP7_75t_L g1794 ( 
.A(n_1759),
.B(n_1744),
.Y(n_1794)
);

AND2x2_ASAP7_75t_L g1795 ( 
.A(n_1750),
.B(n_1742),
.Y(n_1795)
);

INVx2_ASAP7_75t_L g1796 ( 
.A(n_1754),
.Y(n_1796)
);

HB1xp67_ASAP7_75t_L g1797 ( 
.A(n_1774),
.Y(n_1797)
);

INVx2_ASAP7_75t_L g1798 ( 
.A(n_1754),
.Y(n_1798)
);

HB1xp67_ASAP7_75t_L g1799 ( 
.A(n_1757),
.Y(n_1799)
);

INVx1_ASAP7_75t_L g1800 ( 
.A(n_1751),
.Y(n_1800)
);

INVx1_ASAP7_75t_L g1801 ( 
.A(n_1763),
.Y(n_1801)
);

OAI22xp5_ASAP7_75t_L g1802 ( 
.A1(n_1756),
.A2(n_1716),
.B1(n_1733),
.B2(n_1586),
.Y(n_1802)
);

AND2x2_ASAP7_75t_L g1803 ( 
.A(n_1761),
.B(n_1743),
.Y(n_1803)
);

OAI22xp5_ASAP7_75t_L g1804 ( 
.A1(n_1757),
.A2(n_1716),
.B1(n_1733),
.B2(n_1745),
.Y(n_1804)
);

AOI22xp33_ASAP7_75t_L g1805 ( 
.A1(n_1756),
.A2(n_1716),
.B1(n_1725),
.B2(n_1563),
.Y(n_1805)
);

NAND2xp5_ASAP7_75t_L g1806 ( 
.A(n_1748),
.B(n_1716),
.Y(n_1806)
);

INVx2_ASAP7_75t_SL g1807 ( 
.A(n_1752),
.Y(n_1807)
);

INVx2_ASAP7_75t_L g1808 ( 
.A(n_1760),
.Y(n_1808)
);

OAI22xp5_ASAP7_75t_L g1809 ( 
.A1(n_1783),
.A2(n_1716),
.B1(n_1700),
.B2(n_1576),
.Y(n_1809)
);

NAND2xp5_ASAP7_75t_L g1810 ( 
.A(n_1797),
.B(n_1752),
.Y(n_1810)
);

NOR2xp33_ASAP7_75t_SL g1811 ( 
.A(n_1799),
.B(n_1755),
.Y(n_1811)
);

INVx1_ASAP7_75t_L g1812 ( 
.A(n_1791),
.Y(n_1812)
);

NAND2xp5_ASAP7_75t_L g1813 ( 
.A(n_1785),
.B(n_1749),
.Y(n_1813)
);

AOI22xp5_ASAP7_75t_L g1814 ( 
.A1(n_1803),
.A2(n_1760),
.B1(n_1768),
.B2(n_1778),
.Y(n_1814)
);

O2A1O1Ixp5_ASAP7_75t_L g1815 ( 
.A1(n_1793),
.A2(n_1779),
.B(n_1769),
.C(n_1753),
.Y(n_1815)
);

AND2x4_ASAP7_75t_L g1816 ( 
.A(n_1792),
.B(n_1768),
.Y(n_1816)
);

AND2x2_ASAP7_75t_L g1817 ( 
.A(n_1784),
.B(n_1778),
.Y(n_1817)
);

NOR2xp33_ASAP7_75t_L g1818 ( 
.A(n_1786),
.B(n_1789),
.Y(n_1818)
);

NOR2xp33_ASAP7_75t_L g1819 ( 
.A(n_1794),
.B(n_1769),
.Y(n_1819)
);

INVx1_ASAP7_75t_SL g1820 ( 
.A(n_1795),
.Y(n_1820)
);

AOI22x1_ASAP7_75t_L g1821 ( 
.A1(n_1796),
.A2(n_1779),
.B1(n_1765),
.B2(n_1753),
.Y(n_1821)
);

AND2x2_ASAP7_75t_SL g1822 ( 
.A(n_1803),
.B(n_1765),
.Y(n_1822)
);

INVx1_ASAP7_75t_L g1823 ( 
.A(n_1791),
.Y(n_1823)
);

O2A1O1Ixp33_ASAP7_75t_SL g1824 ( 
.A1(n_1796),
.A2(n_1771),
.B(n_1700),
.C(n_1775),
.Y(n_1824)
);

OR2x2_ASAP7_75t_L g1825 ( 
.A(n_1808),
.B(n_1770),
.Y(n_1825)
);

AOI21xp5_ASAP7_75t_L g1826 ( 
.A1(n_1802),
.A2(n_1766),
.B(n_1767),
.Y(n_1826)
);

INVx1_ASAP7_75t_L g1827 ( 
.A(n_1800),
.Y(n_1827)
);

NAND2xp5_ASAP7_75t_L g1828 ( 
.A(n_1787),
.B(n_1772),
.Y(n_1828)
);

A2O1A1Ixp33_ASAP7_75t_L g1829 ( 
.A1(n_1805),
.A2(n_1702),
.B(n_1698),
.C(n_1773),
.Y(n_1829)
);

NOR2xp33_ASAP7_75t_SL g1830 ( 
.A(n_1787),
.B(n_1776),
.Y(n_1830)
);

NAND2xp5_ASAP7_75t_L g1831 ( 
.A(n_1820),
.B(n_1787),
.Y(n_1831)
);

NAND2xp5_ASAP7_75t_L g1832 ( 
.A(n_1822),
.B(n_1784),
.Y(n_1832)
);

NOR2xp33_ASAP7_75t_L g1833 ( 
.A(n_1818),
.B(n_1795),
.Y(n_1833)
);

INVxp33_ASAP7_75t_L g1834 ( 
.A(n_1819),
.Y(n_1834)
);

NAND2xp5_ASAP7_75t_L g1835 ( 
.A(n_1817),
.B(n_1790),
.Y(n_1835)
);

NAND2xp5_ASAP7_75t_L g1836 ( 
.A(n_1816),
.B(n_1790),
.Y(n_1836)
);

OR2x2_ASAP7_75t_L g1837 ( 
.A(n_1813),
.B(n_1808),
.Y(n_1837)
);

INVx1_ASAP7_75t_L g1838 ( 
.A(n_1812),
.Y(n_1838)
);

AND2x2_ASAP7_75t_L g1839 ( 
.A(n_1816),
.B(n_1788),
.Y(n_1839)
);

NAND2xp5_ASAP7_75t_L g1840 ( 
.A(n_1810),
.B(n_1800),
.Y(n_1840)
);

INVx1_ASAP7_75t_SL g1841 ( 
.A(n_1811),
.Y(n_1841)
);

NOR2xp33_ASAP7_75t_L g1842 ( 
.A(n_1830),
.B(n_1792),
.Y(n_1842)
);

AOI21xp5_ASAP7_75t_L g1843 ( 
.A1(n_1841),
.A2(n_1834),
.B(n_1830),
.Y(n_1843)
);

OAI211xp5_ASAP7_75t_L g1844 ( 
.A1(n_1842),
.A2(n_1821),
.B(n_1829),
.C(n_1824),
.Y(n_1844)
);

OAI211xp5_ASAP7_75t_SL g1845 ( 
.A1(n_1832),
.A2(n_1815),
.B(n_1828),
.C(n_1827),
.Y(n_1845)
);

AOI222xp33_ASAP7_75t_L g1846 ( 
.A1(n_1842),
.A2(n_1811),
.B1(n_1802),
.B2(n_1823),
.C1(n_1804),
.C2(n_1801),
.Y(n_1846)
);

CKINVDCx5p33_ASAP7_75t_R g1847 ( 
.A(n_1831),
.Y(n_1847)
);

OAI221xp5_ASAP7_75t_SL g1848 ( 
.A1(n_1836),
.A2(n_1826),
.B1(n_1814),
.B2(n_1825),
.C(n_1806),
.Y(n_1848)
);

NOR2xp33_ASAP7_75t_SL g1849 ( 
.A(n_1833),
.B(n_1796),
.Y(n_1849)
);

INVx2_ASAP7_75t_L g1850 ( 
.A(n_1839),
.Y(n_1850)
);

INVx1_ASAP7_75t_L g1851 ( 
.A(n_1837),
.Y(n_1851)
);

AOI221xp5_ASAP7_75t_L g1852 ( 
.A1(n_1840),
.A2(n_1801),
.B1(n_1809),
.B2(n_1807),
.C(n_1808),
.Y(n_1852)
);

INVx1_ASAP7_75t_L g1853 ( 
.A(n_1851),
.Y(n_1853)
);

AOI21xp33_ASAP7_75t_L g1854 ( 
.A1(n_1845),
.A2(n_1835),
.B(n_1798),
.Y(n_1854)
);

OAI211xp5_ASAP7_75t_L g1855 ( 
.A1(n_1844),
.A2(n_1838),
.B(n_1798),
.C(n_1807),
.Y(n_1855)
);

INVx1_ASAP7_75t_L g1856 ( 
.A(n_1850),
.Y(n_1856)
);

AOI22xp33_ASAP7_75t_L g1857 ( 
.A1(n_1846),
.A2(n_1843),
.B1(n_1792),
.B2(n_1847),
.Y(n_1857)
);

NOR2xp33_ASAP7_75t_L g1858 ( 
.A(n_1849),
.B(n_1848),
.Y(n_1858)
);

INVx1_ASAP7_75t_SL g1859 ( 
.A(n_1853),
.Y(n_1859)
);

INVx3_ASAP7_75t_L g1860 ( 
.A(n_1856),
.Y(n_1860)
);

INVxp67_ASAP7_75t_L g1861 ( 
.A(n_1858),
.Y(n_1861)
);

INVxp67_ASAP7_75t_L g1862 ( 
.A(n_1855),
.Y(n_1862)
);

AND2x2_ASAP7_75t_L g1863 ( 
.A(n_1857),
.B(n_1788),
.Y(n_1863)
);

AOI21xp5_ASAP7_75t_L g1864 ( 
.A1(n_1854),
.A2(n_1852),
.B(n_1798),
.Y(n_1864)
);

OR2x2_ASAP7_75t_L g1865 ( 
.A(n_1856),
.B(n_1792),
.Y(n_1865)
);

NOR2x1_ASAP7_75t_L g1866 ( 
.A(n_1860),
.B(n_1735),
.Y(n_1866)
);

INVx1_ASAP7_75t_L g1867 ( 
.A(n_1865),
.Y(n_1867)
);

INVx1_ASAP7_75t_SL g1868 ( 
.A(n_1859),
.Y(n_1868)
);

CKINVDCx20_ASAP7_75t_R g1869 ( 
.A(n_1861),
.Y(n_1869)
);

AND2x4_ASAP7_75t_L g1870 ( 
.A(n_1860),
.B(n_1780),
.Y(n_1870)
);

CKINVDCx12_ASAP7_75t_R g1871 ( 
.A(n_1869),
.Y(n_1871)
);

NOR2x1_ASAP7_75t_L g1872 ( 
.A(n_1867),
.B(n_1863),
.Y(n_1872)
);

NAND2xp5_ASAP7_75t_SL g1873 ( 
.A(n_1870),
.B(n_1864),
.Y(n_1873)
);

NAND4xp75_ASAP7_75t_L g1874 ( 
.A(n_1872),
.B(n_1866),
.C(n_1862),
.D(n_1868),
.Y(n_1874)
);

NOR3xp33_ASAP7_75t_L g1875 ( 
.A(n_1874),
.B(n_1873),
.C(n_1871),
.Y(n_1875)
);

NAND2x1p5_ASAP7_75t_L g1876 ( 
.A(n_1875),
.B(n_1780),
.Y(n_1876)
);

AOI22xp33_ASAP7_75t_L g1877 ( 
.A1(n_1875),
.A2(n_1696),
.B1(n_1691),
.B2(n_1695),
.Y(n_1877)
);

INVx1_ASAP7_75t_L g1878 ( 
.A(n_1876),
.Y(n_1878)
);

NAND2xp5_ASAP7_75t_L g1879 ( 
.A(n_1877),
.B(n_1740),
.Y(n_1879)
);

AOI22xp33_ASAP7_75t_L g1880 ( 
.A1(n_1878),
.A2(n_1711),
.B1(n_1695),
.B2(n_1691),
.Y(n_1880)
);

OAI22xp5_ASAP7_75t_L g1881 ( 
.A1(n_1879),
.A2(n_1747),
.B1(n_1746),
.B2(n_1740),
.Y(n_1881)
);

INVx1_ASAP7_75t_L g1882 ( 
.A(n_1881),
.Y(n_1882)
);

AOI21xp5_ASAP7_75t_L g1883 ( 
.A1(n_1882),
.A2(n_1880),
.B(n_1746),
.Y(n_1883)
);

AOI22xp5_ASAP7_75t_L g1884 ( 
.A1(n_1883),
.A2(n_1747),
.B1(n_1731),
.B2(n_1707),
.Y(n_1884)
);

AOI22xp33_ASAP7_75t_L g1885 ( 
.A1(n_1884),
.A2(n_1691),
.B1(n_1695),
.B2(n_1696),
.Y(n_1885)
);

AOI22xp5_ASAP7_75t_L g1886 ( 
.A1(n_1885),
.A2(n_1711),
.B1(n_1708),
.B2(n_1737),
.Y(n_1886)
);

AOI211xp5_ASAP7_75t_L g1887 ( 
.A1(n_1886),
.A2(n_1696),
.B(n_1695),
.C(n_1691),
.Y(n_1887)
);


endmodule