module fake_jpeg_13799_n_128 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_128);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_128;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_120;
wire n_43;
wire n_118;
wire n_100;
wire n_82;
wire n_96;

INVx2_ASAP7_75t_L g41 ( 
.A(n_23),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_3),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_12),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_25),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

BUFx8_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_28),
.Y(n_47)
);

BUFx4f_ASAP7_75t_SL g48 ( 
.A(n_40),
.Y(n_48)
);

CKINVDCx16_ASAP7_75t_R g49 ( 
.A(n_17),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_19),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_20),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_21),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_0),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_5),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

AND2x2_ASAP7_75t_L g56 ( 
.A(n_29),
.B(n_26),
.Y(n_56)
);

CKINVDCx14_ASAP7_75t_R g57 ( 
.A(n_15),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_42),
.B(n_53),
.Y(n_58)
);

A2O1A1Ixp33_ASAP7_75t_L g79 ( 
.A1(n_58),
.A2(n_62),
.B(n_56),
.C(n_49),
.Y(n_79)
);

INVx13_ASAP7_75t_L g59 ( 
.A(n_57),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g77 ( 
.A(n_59),
.Y(n_77)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_54),
.Y(n_60)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_60),
.Y(n_68)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_46),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_61),
.B(n_64),
.Y(n_71)
);

AOI21xp5_ASAP7_75t_L g62 ( 
.A1(n_56),
.A2(n_14),
.B(n_38),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_48),
.Y(n_63)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_63),
.Y(n_69)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_46),
.Y(n_64)
);

INVx11_ASAP7_75t_L g65 ( 
.A(n_48),
.Y(n_65)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_65),
.Y(n_70)
);

INVx8_ASAP7_75t_L g66 ( 
.A(n_54),
.Y(n_66)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_66),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_L g67 ( 
.A1(n_60),
.A2(n_41),
.B1(n_50),
.B2(n_52),
.Y(n_67)
);

INVx6_ASAP7_75t_L g93 ( 
.A(n_67),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_61),
.A2(n_47),
.B1(n_44),
.B2(n_51),
.Y(n_73)
);

INVxp67_ASAP7_75t_L g80 ( 
.A(n_73),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_59),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_74),
.B(n_76),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_61),
.A2(n_55),
.B1(n_45),
.B2(n_43),
.Y(n_75)
);

CKINVDCx16_ASAP7_75t_R g87 ( 
.A(n_75),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_66),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_64),
.A2(n_57),
.B1(n_1),
.B2(n_2),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_78),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_79),
.B(n_1),
.Y(n_89)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_68),
.Y(n_81)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_81),
.Y(n_104)
);

CKINVDCx14_ASAP7_75t_R g82 ( 
.A(n_71),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_82),
.B(n_85),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_70),
.B(n_0),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_83),
.B(n_88),
.Y(n_103)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_72),
.Y(n_85)
);

INVxp33_ASAP7_75t_L g88 ( 
.A(n_77),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_89),
.B(n_90),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_73),
.B(n_63),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_77),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_91),
.Y(n_100)
);

NOR2x1_ASAP7_75t_L g92 ( 
.A(n_67),
.B(n_2),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_L g98 ( 
.A1(n_92),
.A2(n_86),
.B(n_80),
.Y(n_98)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_69),
.Y(n_94)
);

INVx6_ASAP7_75t_L g107 ( 
.A(n_94),
.Y(n_107)
);

XNOR2xp5_ASAP7_75t_L g95 ( 
.A(n_92),
.B(n_16),
.Y(n_95)
);

XNOR2xp5_ASAP7_75t_SL g113 ( 
.A(n_95),
.B(n_97),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_93),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_96),
.A2(n_102),
.B1(n_13),
.B2(n_18),
.Y(n_110)
);

XNOR2x1_ASAP7_75t_L g97 ( 
.A(n_87),
.B(n_22),
.Y(n_97)
);

AOI21xp5_ASAP7_75t_L g109 ( 
.A1(n_98),
.A2(n_105),
.B(n_11),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_93),
.A2(n_4),
.B1(n_6),
.B2(n_7),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_101),
.B(n_106),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_84),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_L g105 ( 
.A1(n_88),
.A2(n_8),
.B(n_9),
.Y(n_105)
);

XOR2xp5_ASAP7_75t_L g106 ( 
.A(n_92),
.B(n_10),
.Y(n_106)
);

AOI322xp5_ASAP7_75t_SL g117 ( 
.A1(n_109),
.A2(n_114),
.A3(n_99),
.B1(n_97),
.B2(n_106),
.C1(n_95),
.C2(n_37),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_110),
.B(n_116),
.Y(n_118)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_104),
.Y(n_111)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_111),
.Y(n_119)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_107),
.Y(n_112)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_112),
.Y(n_120)
);

FAx1_ASAP7_75t_SL g114 ( 
.A(n_108),
.B(n_24),
.CI(n_27),
.CON(n_114),
.SN(n_114)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_107),
.Y(n_116)
);

AO221x1_ASAP7_75t_L g122 ( 
.A1(n_117),
.A2(n_114),
.B1(n_31),
.B2(n_32),
.C(n_33),
.Y(n_122)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_119),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_121),
.A2(n_122),
.B1(n_118),
.B2(n_100),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_123),
.B(n_118),
.C(n_115),
.Y(n_124)
);

AOI21xp5_ASAP7_75t_SL g125 ( 
.A1(n_124),
.A2(n_115),
.B(n_120),
.Y(n_125)
);

NOR3xp33_ASAP7_75t_L g126 ( 
.A(n_125),
.B(n_103),
.C(n_113),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_126),
.B(n_30),
.Y(n_127)
);

XOR2xp5_ASAP7_75t_L g128 ( 
.A(n_127),
.B(n_39),
.Y(n_128)
);


endmodule