module fake_jpeg_24081_n_308 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_308);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_308;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_208;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_8),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

INVx11_ASAP7_75t_SL g22 ( 
.A(n_17),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_15),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_1),
.B(n_7),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_16),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_0),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_8),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_6),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_17),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_9),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_1),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_14),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_21),
.Y(n_39)
);

INVx5_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_26),
.B(n_0),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_40),
.B(n_42),
.Y(n_63)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_21),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_41),
.B(n_45),
.Y(n_60)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_20),
.Y(n_42)
);

INVx11_ASAP7_75t_L g43 ( 
.A(n_22),
.Y(n_43)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_43),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_21),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_44),
.Y(n_62)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_20),
.Y(n_45)
);

AOI21xp33_ASAP7_75t_L g46 ( 
.A1(n_26),
.A2(n_10),
.B(n_16),
.Y(n_46)
);

A2O1A1Ixp33_ASAP7_75t_L g68 ( 
.A1(n_46),
.A2(n_30),
.B(n_25),
.C(n_18),
.Y(n_68)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_20),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_47),
.B(n_49),
.Y(n_76)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_24),
.Y(n_48)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_48),
.Y(n_77)
);

INVx1_ASAP7_75t_SL g49 ( 
.A(n_32),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_42),
.A2(n_23),
.B1(n_22),
.B2(n_32),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_50),
.A2(n_67),
.B1(n_47),
.B2(n_43),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g52 ( 
.A1(n_42),
.A2(n_23),
.B1(n_24),
.B2(n_35),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_52),
.A2(n_53),
.B1(n_57),
.B2(n_66),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_L g53 ( 
.A1(n_48),
.A2(n_35),
.B1(n_24),
.B2(n_38),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_40),
.B(n_19),
.Y(n_54)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_54),
.B(n_58),
.Y(n_87)
);

HB1xp67_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_55),
.Y(n_83)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

INVx5_ASAP7_75t_L g98 ( 
.A(n_56),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g57 ( 
.A1(n_42),
.A2(n_23),
.B1(n_35),
.B2(n_32),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_40),
.B(n_19),
.Y(n_58)
);

MAJIxp5_ASAP7_75t_L g61 ( 
.A(n_41),
.B(n_37),
.C(n_38),
.Y(n_61)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_61),
.B(n_49),
.C(n_45),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_44),
.B(n_37),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_64),
.B(n_72),
.Y(n_82)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_39),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_65),
.B(n_70),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_L g66 ( 
.A1(n_48),
.A2(n_29),
.B1(n_25),
.B2(n_18),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_42),
.A2(n_36),
.B1(n_28),
.B2(n_29),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_68),
.B(n_14),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_47),
.A2(n_36),
.B1(n_28),
.B2(n_30),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_69),
.A2(n_71),
.B1(n_80),
.B2(n_43),
.Y(n_89)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_39),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_L g71 ( 
.A1(n_48),
.A2(n_33),
.B1(n_27),
.B2(n_31),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_44),
.B(n_33),
.Y(n_72)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_44),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_73),
.B(n_47),
.Y(n_90)
);

CKINVDCx16_ASAP7_75t_R g74 ( 
.A(n_44),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_74),
.B(n_79),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_44),
.B(n_33),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_75),
.B(n_34),
.Y(n_104)
);

HB1xp67_ASAP7_75t_L g78 ( 
.A(n_43),
.Y(n_78)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_78),
.Y(n_88)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_48),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_L g80 ( 
.A1(n_43),
.A2(n_33),
.B1(n_27),
.B2(n_31),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_84),
.A2(n_9),
.B1(n_16),
.B2(n_15),
.Y(n_141)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_78),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_85),
.B(n_92),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_L g128 ( 
.A1(n_89),
.A2(n_74),
.B1(n_77),
.B2(n_79),
.Y(n_128)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_90),
.Y(n_120)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_64),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_91),
.B(n_94),
.Y(n_140)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_55),
.Y(n_92)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_69),
.Y(n_94)
);

INVx8_ASAP7_75t_L g95 ( 
.A(n_62),
.Y(n_95)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_95),
.Y(n_129)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_51),
.Y(n_96)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_96),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_54),
.B(n_1),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_97),
.B(n_99),
.Y(n_124)
);

INVx13_ASAP7_75t_L g100 ( 
.A(n_56),
.Y(n_100)
);

INVx13_ASAP7_75t_L g144 ( 
.A(n_100),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_68),
.A2(n_47),
.B1(n_41),
.B2(n_45),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_101),
.A2(n_112),
.B1(n_2),
.B2(n_3),
.Y(n_139)
);

AND2x2_ASAP7_75t_L g123 ( 
.A(n_102),
.B(n_104),
.Y(n_123)
);

INVx8_ASAP7_75t_L g103 ( 
.A(n_62),
.Y(n_103)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_103),
.Y(n_132)
);

NAND2xp67_ASAP7_75t_SL g105 ( 
.A(n_68),
.B(n_49),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g127 ( 
.A(n_105),
.B(n_107),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_63),
.B(n_41),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_106),
.Y(n_131)
);

OR2x4_ASAP7_75t_L g107 ( 
.A(n_63),
.B(n_49),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_65),
.B(n_49),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_108),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_70),
.B(n_45),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_109),
.Y(n_119)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_56),
.Y(n_110)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_110),
.Y(n_121)
);

AOI32xp33_ASAP7_75t_L g111 ( 
.A1(n_76),
.A2(n_27),
.A3(n_34),
.B1(n_31),
.B2(n_11),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_111),
.B(n_101),
.C(n_115),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_57),
.A2(n_34),
.B1(n_31),
.B2(n_27),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_58),
.B(n_2),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_113),
.B(n_9),
.Y(n_148)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_52),
.Y(n_114)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_114),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_60),
.B(n_10),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_115),
.B(n_12),
.Y(n_134)
);

BUFx2_ASAP7_75t_L g116 ( 
.A(n_62),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_116),
.Y(n_143)
);

BUFx12_ASAP7_75t_L g117 ( 
.A(n_51),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g146 ( 
.A(n_117),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_105),
.A2(n_75),
.B1(n_72),
.B2(n_76),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g162 ( 
.A(n_118),
.Y(n_162)
);

AOI21xp5_ASAP7_75t_L g125 ( 
.A1(n_107),
.A2(n_60),
.B(n_77),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_L g169 ( 
.A1(n_125),
.A2(n_126),
.B(n_134),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_128),
.A2(n_136),
.B1(n_139),
.B2(n_85),
.Y(n_154)
);

AND2x2_ASAP7_75t_L g130 ( 
.A(n_82),
.B(n_61),
.Y(n_130)
);

AND2x2_ASAP7_75t_L g177 ( 
.A(n_130),
.B(n_3),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_SL g181 ( 
.A(n_134),
.B(n_148),
.Y(n_181)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_110),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_135),
.B(n_116),
.Y(n_158)
);

AOI22xp33_ASAP7_75t_L g136 ( 
.A1(n_94),
.A2(n_34),
.B1(n_73),
.B2(n_59),
.Y(n_136)
);

AND2x6_ASAP7_75t_L g137 ( 
.A(n_87),
.B(n_11),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_L g155 ( 
.A(n_137),
.B(n_113),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_82),
.B(n_59),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_138),
.B(n_145),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_141),
.A2(n_142),
.B1(n_147),
.B2(n_97),
.Y(n_156)
);

O2A1O1Ixp33_ASAP7_75t_L g142 ( 
.A1(n_86),
.A2(n_2),
.B(n_3),
.C(n_4),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_91),
.B(n_3),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_114),
.A2(n_104),
.B1(n_99),
.B2(n_102),
.Y(n_147)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_149),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_151),
.B(n_155),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_138),
.B(n_87),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_153),
.B(n_159),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_154),
.A2(n_175),
.B1(n_120),
.B2(n_122),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_156),
.A2(n_157),
.B1(n_137),
.B2(n_124),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_150),
.A2(n_111),
.B1(n_86),
.B2(n_87),
.Y(n_157)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_158),
.Y(n_184)
);

OR2x2_ASAP7_75t_L g159 ( 
.A(n_131),
.B(n_93),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_145),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_160),
.B(n_171),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_140),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_161),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_131),
.B(n_83),
.Y(n_163)
);

CKINVDCx16_ASAP7_75t_R g191 ( 
.A(n_163),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_133),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_164),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_133),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_165),
.Y(n_202)
);

CKINVDCx16_ASAP7_75t_R g166 ( 
.A(n_139),
.Y(n_166)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_166),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_147),
.B(n_89),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_167),
.B(n_126),
.C(n_123),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_119),
.B(n_83),
.Y(n_168)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_168),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_169),
.B(n_177),
.Y(n_205)
);

INVx1_ASAP7_75t_SL g170 ( 
.A(n_125),
.Y(n_170)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_170),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_130),
.B(n_93),
.Y(n_171)
);

AO21x1_ASAP7_75t_L g172 ( 
.A1(n_127),
.A2(n_142),
.B(n_150),
.Y(n_172)
);

AOI21xp5_ASAP7_75t_L g198 ( 
.A1(n_172),
.A2(n_122),
.B(n_146),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_SL g173 ( 
.A1(n_129),
.A2(n_96),
.B1(n_95),
.B2(n_103),
.Y(n_173)
);

OAI22x1_ASAP7_75t_L g190 ( 
.A1(n_173),
.A2(n_179),
.B1(n_116),
.B2(n_132),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_130),
.B(n_88),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_L g199 ( 
.A1(n_174),
.A2(n_176),
.B(n_148),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_118),
.A2(n_112),
.B1(n_88),
.B2(n_92),
.Y(n_175)
);

OR2x2_ASAP7_75t_L g176 ( 
.A(n_127),
.B(n_81),
.Y(n_176)
);

INVx3_ASAP7_75t_L g178 ( 
.A(n_121),
.Y(n_178)
);

HB1xp67_ASAP7_75t_L g189 ( 
.A(n_178),
.Y(n_189)
);

AOI22xp33_ASAP7_75t_SL g179 ( 
.A1(n_129),
.A2(n_95),
.B1(n_103),
.B2(n_98),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_119),
.B(n_117),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_SL g209 ( 
.A(n_180),
.B(n_182),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_120),
.B(n_117),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_183),
.B(n_186),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_L g218 ( 
.A1(n_185),
.A2(n_203),
.B1(n_206),
.B2(n_178),
.Y(n_218)
);

MAJx2_ASAP7_75t_L g186 ( 
.A(n_169),
.B(n_123),
.C(n_127),
.Y(n_186)
);

XOR2x2_ASAP7_75t_L g187 ( 
.A(n_170),
.B(n_123),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_SL g229 ( 
.A1(n_187),
.A2(n_190),
.B(n_198),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_194),
.B(n_155),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_174),
.B(n_124),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_197),
.B(n_171),
.C(n_152),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_L g217 ( 
.A1(n_199),
.A2(n_170),
.B(n_152),
.Y(n_217)
);

OA21x2_ASAP7_75t_L g200 ( 
.A1(n_172),
.A2(n_132),
.B(n_117),
.Y(n_200)
);

AOI21xp5_ASAP7_75t_L g231 ( 
.A1(n_200),
.A2(n_158),
.B(n_182),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_157),
.A2(n_143),
.B1(n_135),
.B2(n_121),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_201),
.A2(n_180),
.B1(n_168),
.B2(n_172),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_166),
.A2(n_143),
.B1(n_98),
.B2(n_146),
.Y(n_203)
);

NAND3xp33_ASAP7_75t_L g204 ( 
.A(n_153),
.B(n_12),
.C(n_17),
.Y(n_204)
);

NAND3xp33_ASAP7_75t_L g215 ( 
.A(n_204),
.B(n_13),
.C(n_7),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_175),
.A2(n_100),
.B1(n_144),
.B2(n_4),
.Y(n_206)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_189),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_211),
.B(n_214),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_212),
.B(n_226),
.C(n_197),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_202),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_213),
.Y(n_250)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_207),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_215),
.B(n_216),
.Y(n_243)
);

NAND3xp33_ASAP7_75t_SL g216 ( 
.A(n_207),
.B(n_161),
.C(n_156),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_217),
.B(n_228),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_218),
.A2(n_219),
.B1(n_222),
.B2(n_193),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_L g219 ( 
.A1(n_208),
.A2(n_162),
.B1(n_164),
.B2(n_165),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_202),
.B(n_163),
.Y(n_220)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_220),
.Y(n_239)
);

AND2x2_ASAP7_75t_L g221 ( 
.A(n_201),
.B(n_176),
.Y(n_221)
);

AOI21xp5_ASAP7_75t_L g236 ( 
.A1(n_221),
.A2(n_231),
.B(n_198),
.Y(n_236)
);

HAxp5_ASAP7_75t_SL g224 ( 
.A(n_208),
.B(n_176),
.CON(n_224),
.SN(n_224)
);

NAND3xp33_ASAP7_75t_L g235 ( 
.A(n_224),
.B(n_195),
.C(n_210),
.Y(n_235)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_203),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_225),
.B(n_233),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_183),
.B(n_167),
.C(n_160),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_210),
.B(n_177),
.Y(n_227)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_227),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_196),
.Y(n_228)
);

HB1xp67_ASAP7_75t_L g230 ( 
.A(n_190),
.Y(n_230)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_230),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_232),
.B(n_205),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_SL g233 ( 
.A(n_192),
.B(n_181),
.Y(n_233)
);

XNOR2x1_ASAP7_75t_L g234 ( 
.A(n_221),
.B(n_187),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_SL g257 ( 
.A(n_234),
.B(n_222),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_235),
.B(n_252),
.Y(n_258)
);

OAI21xp5_ASAP7_75t_SL g263 ( 
.A1(n_236),
.A2(n_244),
.B(n_229),
.Y(n_263)
);

INVxp67_ASAP7_75t_L g240 ( 
.A(n_220),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_240),
.B(n_246),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_242),
.B(n_212),
.C(n_217),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_L g245 ( 
.A1(n_230),
.A2(n_193),
.B1(n_185),
.B2(n_206),
.Y(n_245)
);

CKINVDCx16_ASAP7_75t_R g255 ( 
.A(n_245),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_L g246 ( 
.A1(n_225),
.A2(n_195),
.B1(n_191),
.B2(n_200),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_SL g247 ( 
.A(n_223),
.B(n_186),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_247),
.B(n_248),
.Y(n_259)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_219),
.Y(n_252)
);

OAI22xp33_ASAP7_75t_L g254 ( 
.A1(n_251),
.A2(n_200),
.B1(n_213),
.B2(n_231),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_254),
.A2(n_263),
.B1(n_252),
.B2(n_251),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_242),
.B(n_226),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_256),
.B(n_260),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_257),
.B(n_262),
.C(n_264),
.Y(n_270)
);

INVx13_ASAP7_75t_L g260 ( 
.A(n_250),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_248),
.B(n_223),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_261),
.B(n_265),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_247),
.B(n_232),
.C(n_188),
.Y(n_264)
);

HB1xp67_ASAP7_75t_L g265 ( 
.A(n_234),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_SL g266 ( 
.A(n_244),
.B(n_194),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_266),
.B(n_229),
.C(n_236),
.Y(n_271)
);

AOI322xp5_ASAP7_75t_SL g267 ( 
.A1(n_243),
.A2(n_233),
.A3(n_205),
.B1(n_177),
.B2(n_199),
.C1(n_159),
.C2(n_221),
.Y(n_267)
);

OAI21xp5_ASAP7_75t_L g269 ( 
.A1(n_267),
.A2(n_227),
.B(n_237),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_250),
.B(n_228),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_SL g277 ( 
.A(n_268),
.B(n_239),
.Y(n_277)
);

AOI321xp33_ASAP7_75t_L g284 ( 
.A1(n_269),
.A2(n_275),
.A3(n_279),
.B1(n_209),
.B2(n_181),
.C(n_218),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_271),
.B(n_273),
.C(n_274),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_272),
.B(n_280),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_262),
.B(n_238),
.C(n_241),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_259),
.B(n_238),
.C(n_241),
.Y(n_274)
);

OAI21xp5_ASAP7_75t_L g275 ( 
.A1(n_258),
.A2(n_249),
.B(n_240),
.Y(n_275)
);

AOI21xp5_ASAP7_75t_L g286 ( 
.A1(n_275),
.A2(n_184),
.B(n_151),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_259),
.B(n_264),
.C(n_257),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_276),
.B(n_277),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_255),
.A2(n_249),
.B1(n_239),
.B2(n_214),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_L g283 ( 
.A1(n_271),
.A2(n_253),
.B1(n_263),
.B2(n_260),
.Y(n_283)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_283),
.Y(n_289)
);

OAI321xp33_ASAP7_75t_L g292 ( 
.A1(n_284),
.A2(n_286),
.A3(n_287),
.B1(n_154),
.B2(n_184),
.C(n_282),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_273),
.B(n_254),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_285),
.B(n_274),
.Y(n_290)
);

OAI21x1_ASAP7_75t_L g287 ( 
.A1(n_278),
.A2(n_266),
.B(n_159),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_290),
.B(n_291),
.Y(n_298)
);

AND2x2_ASAP7_75t_L g291 ( 
.A(n_281),
.B(n_270),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_SL g299 ( 
.A(n_292),
.B(n_293),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_285),
.B(n_211),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_288),
.B(n_270),
.C(n_276),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_294),
.B(n_144),
.C(n_100),
.Y(n_300)
);

HB1xp67_ASAP7_75t_L g295 ( 
.A(n_287),
.Y(n_295)
);

CKINVDCx16_ASAP7_75t_R g297 ( 
.A(n_295),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_289),
.A2(n_295),
.B1(n_261),
.B2(n_256),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_296),
.B(n_300),
.C(n_7),
.Y(n_301)
);

INVxp67_ASAP7_75t_L g304 ( 
.A(n_301),
.Y(n_304)
);

INVxp67_ASAP7_75t_L g302 ( 
.A(n_299),
.Y(n_302)
);

AOI322xp5_ASAP7_75t_L g305 ( 
.A1(n_302),
.A2(n_303),
.A3(n_297),
.B1(n_296),
.B2(n_300),
.C1(n_13),
.C2(n_4),
.Y(n_305)
);

AOI322xp5_ASAP7_75t_L g303 ( 
.A1(n_298),
.A2(n_8),
.A3(n_11),
.B1(n_12),
.B2(n_13),
.C1(n_4),
.C2(n_5),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_SL g306 ( 
.A(n_305),
.B(n_5),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_306),
.B(n_304),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_307),
.B(n_5),
.Y(n_308)
);


endmodule