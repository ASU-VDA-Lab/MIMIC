module fake_jpeg_27409_n_72 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_72);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_72;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_23;
wire n_10;
wire n_69;
wire n_27;
wire n_55;
wire n_64;
wire n_47;
wire n_22;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_20;
wire n_18;
wire n_59;
wire n_35;
wire n_48;
wire n_68;
wire n_52;
wire n_71;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_65;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_11;
wire n_62;
wire n_25;
wire n_31;
wire n_17;
wire n_56;
wire n_67;
wire n_37;
wire n_29;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_70;
wire n_15;
wire n_66;

BUFx6f_ASAP7_75t_L g10 ( 
.A(n_9),
.Y(n_10)
);

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_2),
.Y(n_11)
);

BUFx10_ASAP7_75t_L g12 ( 
.A(n_8),
.Y(n_12)
);

INVx6_ASAP7_75t_SL g13 ( 
.A(n_0),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_2),
.Y(n_14)
);

BUFx12f_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_7),
.B(n_1),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_1),
.Y(n_19)
);

CKINVDCx16_ASAP7_75t_R g20 ( 
.A(n_13),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_SL g32 ( 
.A(n_20),
.B(n_25),
.Y(n_32)
);

INVx8_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

CKINVDCx6p67_ASAP7_75t_R g29 ( 
.A(n_21),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_SL g22 ( 
.A1(n_16),
.A2(n_0),
.B1(n_4),
.B2(n_5),
.Y(n_22)
);

AOI22xp33_ASAP7_75t_L g26 ( 
.A1(n_22),
.A2(n_19),
.B1(n_11),
.B2(n_14),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_15),
.B(n_0),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_SL g28 ( 
.A(n_23),
.B(n_16),
.Y(n_28)
);

BUFx12_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_24),
.Y(n_27)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_25),
.B(n_12),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_SL g37 ( 
.A1(n_26),
.A2(n_14),
.B1(n_11),
.B2(n_10),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_SL g41 ( 
.A(n_28),
.B(n_18),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_30),
.B(n_23),
.Y(n_34)
);

OA22x2_ASAP7_75t_L g31 ( 
.A1(n_21),
.A2(n_19),
.B1(n_12),
.B2(n_15),
.Y(n_31)
);

AOI22xp5_ASAP7_75t_L g36 ( 
.A1(n_31),
.A2(n_21),
.B1(n_13),
.B2(n_20),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_32),
.B(n_18),
.Y(n_39)
);

MAJIxp5_ASAP7_75t_SL g33 ( 
.A(n_28),
.B(n_22),
.C(n_17),
.Y(n_33)
);

OR2x2_ASAP7_75t_L g48 ( 
.A(n_33),
.B(n_37),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_34),
.B(n_35),
.Y(n_46)
);

XNOR2xp5_ASAP7_75t_L g35 ( 
.A(n_30),
.B(n_15),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_SL g43 ( 
.A(n_35),
.B(n_38),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_36),
.A2(n_31),
.B1(n_29),
.B2(n_27),
.Y(n_49)
);

XNOR2xp5_ASAP7_75t_L g38 ( 
.A(n_32),
.B(n_24),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_SL g44 ( 
.A(n_39),
.B(n_41),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_27),
.Y(n_40)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_40),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_40),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_42),
.B(n_29),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_46),
.B(n_47),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_38),
.B(n_36),
.Y(n_47)
);

CKINVDCx14_ASAP7_75t_R g50 ( 
.A(n_49),
.Y(n_50)
);

INVx13_ASAP7_75t_L g52 ( 
.A(n_45),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_52),
.B(n_54),
.Y(n_59)
);

XNOR2xp5_ASAP7_75t_SL g53 ( 
.A(n_46),
.B(n_31),
.Y(n_53)
);

MAJIxp5_ASAP7_75t_L g57 ( 
.A(n_53),
.B(n_56),
.C(n_47),
.Y(n_57)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_49),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_45),
.Y(n_55)
);

INVxp67_ASAP7_75t_L g61 ( 
.A(n_55),
.Y(n_61)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_57),
.Y(n_64)
);

MAJIxp5_ASAP7_75t_L g58 ( 
.A(n_53),
.B(n_43),
.C(n_48),
.Y(n_58)
);

AOI21xp5_ASAP7_75t_L g62 ( 
.A1(n_58),
.A2(n_60),
.B(n_51),
.Y(n_62)
);

MAJIxp5_ASAP7_75t_L g60 ( 
.A(n_51),
.B(n_48),
.C(n_44),
.Y(n_60)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_62),
.B(n_64),
.C(n_24),
.Y(n_68)
);

AOI21xp5_ASAP7_75t_L g63 ( 
.A1(n_59),
.A2(n_54),
.B(n_50),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_63),
.B(n_29),
.Y(n_66)
);

OAI321xp33_ASAP7_75t_L g65 ( 
.A1(n_61),
.A2(n_31),
.A3(n_55),
.B1(n_52),
.B2(n_10),
.C(n_8),
.Y(n_65)
);

A2O1A1Ixp33_ASAP7_75t_SL g67 ( 
.A1(n_65),
.A2(n_4),
.B(n_5),
.C(n_6),
.Y(n_67)
);

XOR2xp5_ASAP7_75t_L g69 ( 
.A(n_66),
.B(n_68),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_67),
.A2(n_29),
.B1(n_7),
.B2(n_9),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_70),
.A2(n_6),
.B1(n_24),
.B2(n_69),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_71),
.B(n_24),
.Y(n_72)
);


endmodule