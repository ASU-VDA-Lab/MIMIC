module fake_jpeg_12971_n_172 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_172);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_172;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx3_ASAP7_75t_SL g51 ( 
.A(n_35),
.Y(n_51)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_28),
.Y(n_52)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_12),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_49),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_16),
.Y(n_55)
);

INVx11_ASAP7_75t_L g56 ( 
.A(n_33),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_18),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_38),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_37),
.Y(n_59)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_7),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_4),
.Y(n_61)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_13),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_7),
.Y(n_63)
);

BUFx5_ASAP7_75t_L g64 ( 
.A(n_11),
.Y(n_64)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_23),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_3),
.Y(n_66)
);

BUFx12f_ASAP7_75t_L g67 ( 
.A(n_44),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_41),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_4),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_11),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_22),
.Y(n_71)
);

BUFx12f_ASAP7_75t_L g72 ( 
.A(n_17),
.Y(n_72)
);

NOR3xp33_ASAP7_75t_L g73 ( 
.A(n_51),
.B(n_56),
.C(n_61),
.Y(n_73)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_73),
.Y(n_89)
);

INVx5_ASAP7_75t_L g74 ( 
.A(n_67),
.Y(n_74)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_74),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_66),
.B(n_0),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_75),
.B(n_79),
.Y(n_83)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_67),
.Y(n_76)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_76),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_62),
.A2(n_25),
.B1(n_48),
.B2(n_47),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_77),
.A2(n_53),
.B1(n_69),
.B2(n_63),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_59),
.Y(n_78)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_78),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_70),
.B(n_0),
.Y(n_79)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_52),
.Y(n_80)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_80),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_54),
.B(n_1),
.Y(n_81)
);

OAI21xp5_ASAP7_75t_SL g96 ( 
.A1(n_81),
.A2(n_51),
.B(n_58),
.Y(n_96)
);

BUFx12f_ASAP7_75t_L g82 ( 
.A(n_64),
.Y(n_82)
);

INVx13_ASAP7_75t_L g94 ( 
.A(n_82),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_84),
.A2(n_92),
.B1(n_55),
.B2(n_65),
.Y(n_102)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_80),
.B(n_76),
.Y(n_85)
);

AO21x1_ASAP7_75t_L g107 ( 
.A1(n_85),
.A2(n_91),
.B(n_72),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_77),
.B(n_57),
.C(n_51),
.Y(n_86)
);

AOI21xp5_ASAP7_75t_L g101 ( 
.A1(n_86),
.A2(n_51),
.B(n_68),
.Y(n_101)
);

INVx11_ASAP7_75t_L g90 ( 
.A(n_82),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_90),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_74),
.B(n_72),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_L g92 ( 
.A1(n_78),
.A2(n_53),
.B1(n_60),
.B2(n_59),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_96),
.B(n_55),
.Y(n_110)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_82),
.Y(n_97)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_97),
.Y(n_105)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_93),
.Y(n_98)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_98),
.Y(n_118)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_88),
.Y(n_99)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_99),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_L g136 ( 
.A(n_101),
.B(n_107),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_102),
.A2(n_5),
.B1(n_6),
.B2(n_8),
.Y(n_128)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_95),
.Y(n_103)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_103),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_83),
.B(n_1),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_104),
.B(n_109),
.Y(n_123)
);

INVx2_ASAP7_75t_SL g106 ( 
.A(n_87),
.Y(n_106)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_106),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_89),
.B(n_2),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_108),
.B(n_110),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_85),
.Y(n_109)
);

CKINVDCx16_ASAP7_75t_R g111 ( 
.A(n_90),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_111),
.B(n_113),
.Y(n_129)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_85),
.Y(n_112)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_112),
.Y(n_134)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_87),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_86),
.B(n_2),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_114),
.B(n_115),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_84),
.B(n_3),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_89),
.B(n_5),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_116),
.A2(n_6),
.B1(n_8),
.B2(n_9),
.Y(n_132)
);

AOI32xp33_ASAP7_75t_L g117 ( 
.A1(n_91),
.A2(n_71),
.A3(n_65),
.B1(n_29),
.B2(n_30),
.Y(n_117)
);

A2O1A1O1Ixp25_ASAP7_75t_L g127 ( 
.A1(n_117),
.A2(n_94),
.B(n_26),
.C(n_27),
.D(n_50),
.Y(n_127)
);

INVx13_ASAP7_75t_L g120 ( 
.A(n_106),
.Y(n_120)
);

CKINVDCx5p33_ASAP7_75t_R g144 ( 
.A(n_120),
.Y(n_144)
);

INVx13_ASAP7_75t_L g121 ( 
.A(n_105),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_121),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_107),
.A2(n_71),
.B1(n_91),
.B2(n_94),
.Y(n_122)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_122),
.Y(n_140)
);

NAND3xp33_ASAP7_75t_L g154 ( 
.A(n_127),
.B(n_135),
.C(n_42),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_SL g142 ( 
.A1(n_128),
.A2(n_132),
.B(n_10),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_98),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_130),
.B(n_137),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_101),
.B(n_24),
.C(n_45),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_131),
.B(n_138),
.C(n_19),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_103),
.B(n_9),
.Y(n_135)
);

FAx1_ASAP7_75t_SL g137 ( 
.A(n_100),
.B(n_10),
.CI(n_12),
.CON(n_137),
.SN(n_137)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_113),
.B(n_32),
.C(n_43),
.Y(n_138)
);

AND2x6_ASAP7_75t_L g139 ( 
.A(n_100),
.B(n_31),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_139),
.B(n_20),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_SL g141 ( 
.A(n_134),
.B(n_99),
.Y(n_141)
);

A2O1A1O1Ixp25_ASAP7_75t_L g159 ( 
.A1(n_141),
.A2(n_151),
.B(n_152),
.C(n_137),
.D(n_129),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_142),
.B(n_145),
.Y(n_157)
);

XOR2xp5_ASAP7_75t_L g145 ( 
.A(n_133),
.B(n_34),
.Y(n_145)
);

AOI21xp5_ASAP7_75t_L g146 ( 
.A1(n_124),
.A2(n_13),
.B(n_14),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_L g160 ( 
.A1(n_146),
.A2(n_129),
.B(n_139),
.Y(n_160)
);

XOR2xp5_ASAP7_75t_L g147 ( 
.A(n_136),
.B(n_15),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_147),
.B(n_148),
.Y(n_158)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_149),
.Y(n_161)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_118),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_150),
.A2(n_154),
.B1(n_127),
.B2(n_126),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_123),
.B(n_21),
.C(n_36),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_124),
.B(n_39),
.C(n_40),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_155),
.B(n_159),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_140),
.A2(n_143),
.B1(n_141),
.B2(n_153),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_156),
.A2(n_119),
.B1(n_125),
.B2(n_154),
.Y(n_164)
);

AO221x1_ASAP7_75t_L g163 ( 
.A1(n_160),
.A2(n_158),
.B1(n_157),
.B2(n_161),
.C(n_144),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_SL g162 ( 
.A1(n_159),
.A2(n_144),
.B(n_147),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_162),
.B(n_163),
.C(n_165),
.Y(n_166)
);

INVx1_ASAP7_75t_SL g167 ( 
.A(n_164),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_166),
.B(n_160),
.C(n_164),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_168),
.B(n_167),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_169),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_SL g171 ( 
.A1(n_170),
.A2(n_46),
.B(n_120),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_171),
.B(n_121),
.Y(n_172)
);


endmodule