module real_jpeg_20774_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_336, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_336;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_332;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_83;
wire n_288;
wire n_78;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_286;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_299;
wire n_243;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_0),
.A2(n_26),
.B1(n_33),
.B2(n_134),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_0),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_SL g167 ( 
.A1(n_0),
.A2(n_30),
.B1(n_31),
.B2(n_134),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_0),
.A2(n_46),
.B1(n_47),
.B2(n_134),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_0),
.A2(n_63),
.B1(n_64),
.B2(n_134),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_1),
.Y(n_27)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_2),
.A2(n_30),
.B1(n_31),
.B2(n_129),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_2),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g181 ( 
.A1(n_2),
.A2(n_63),
.B1(n_64),
.B2(n_129),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_SL g227 ( 
.A1(n_2),
.A2(n_46),
.B1(n_47),
.B2(n_129),
.Y(n_227)
);

AOI22xp33_ASAP7_75t_SL g268 ( 
.A1(n_2),
.A2(n_26),
.B1(n_33),
.B2(n_129),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_3),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_3),
.B(n_29),
.Y(n_164)
);

AOI21xp33_ASAP7_75t_L g185 ( 
.A1(n_3),
.A2(n_6),
.B(n_64),
.Y(n_185)
);

AOI22xp33_ASAP7_75t_SL g188 ( 
.A1(n_3),
.A2(n_46),
.B1(n_47),
.B2(n_132),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_3),
.A2(n_106),
.B1(n_111),
.B2(n_194),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_3),
.B(n_88),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_3),
.B(n_31),
.Y(n_220)
);

AOI21xp33_ASAP7_75t_L g224 ( 
.A1(n_3),
.A2(n_31),
.B(n_220),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_4),
.B(n_63),
.Y(n_107)
);

INVx8_ASAP7_75t_L g111 ( 
.A(n_4),
.Y(n_111)
);

INVx6_ASAP7_75t_L g161 ( 
.A(n_4),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_5),
.A2(n_30),
.B1(n_31),
.B2(n_51),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_5),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_5),
.A2(n_46),
.B1(n_47),
.B2(n_51),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_5),
.A2(n_51),
.B1(n_63),
.B2(n_64),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_5),
.A2(n_26),
.B1(n_33),
.B2(n_51),
.Y(n_288)
);

A2O1A1Ixp33_ASAP7_75t_L g60 ( 
.A1(n_6),
.A2(n_46),
.B(n_61),
.C(n_62),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_6),
.B(n_46),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_6),
.A2(n_63),
.B1(n_64),
.B2(n_65),
.Y(n_62)
);

INVx6_ASAP7_75t_SL g65 ( 
.A(n_6),
.Y(n_65)
);

BUFx8_ASAP7_75t_L g64 ( 
.A(n_7),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g35 ( 
.A1(n_8),
.A2(n_26),
.B1(n_33),
.B2(n_36),
.Y(n_35)
);

CKINVDCx14_ASAP7_75t_R g36 ( 
.A(n_8),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_8),
.A2(n_30),
.B1(n_31),
.B2(n_36),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_8),
.A2(n_36),
.B1(n_63),
.B2(n_64),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g260 ( 
.A1(n_8),
.A2(n_36),
.B1(n_46),
.B2(n_47),
.Y(n_260)
);

AOI22xp33_ASAP7_75t_L g126 ( 
.A1(n_9),
.A2(n_30),
.B1(n_31),
.B2(n_127),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_9),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_9),
.A2(n_26),
.B1(n_33),
.B2(n_127),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_SL g178 ( 
.A1(n_9),
.A2(n_63),
.B1(n_64),
.B2(n_127),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_SL g209 ( 
.A1(n_9),
.A2(n_46),
.B1(n_47),
.B2(n_127),
.Y(n_209)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

AOI22xp33_ASAP7_75t_SL g32 ( 
.A1(n_11),
.A2(n_26),
.B1(n_33),
.B2(n_34),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_11),
.Y(n_34)
);

AOI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_11),
.A2(n_34),
.B1(n_46),
.B2(n_47),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_11),
.A2(n_34),
.B1(n_63),
.B2(n_64),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_SL g284 ( 
.A1(n_11),
.A2(n_30),
.B1(n_31),
.B2(n_34),
.Y(n_284)
);

INVx13_ASAP7_75t_L g45 ( 
.A(n_12),
.Y(n_45)
);

INVx13_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_L g29 ( 
.A1(n_13),
.A2(n_25),
.B1(n_30),
.B2(n_31),
.Y(n_29)
);

AOI22xp33_ASAP7_75t_L g57 ( 
.A1(n_14),
.A2(n_30),
.B1(n_31),
.B2(n_58),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_14),
.Y(n_58)
);

OAI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_14),
.A2(n_26),
.B1(n_33),
.B2(n_58),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_L g112 ( 
.A1(n_14),
.A2(n_58),
.B1(n_63),
.B2(n_64),
.Y(n_112)
);

OAI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_14),
.A2(n_46),
.B1(n_47),
.B2(n_58),
.Y(n_116)
);

INVx11_ASAP7_75t_SL g48 ( 
.A(n_15),
.Y(n_48)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_95),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_SL g17 ( 
.A(n_18),
.B(n_93),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_79),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_19),
.B(n_79),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_71),
.C(n_74),
.Y(n_19)
);

AOI22xp5_ASAP7_75t_L g328 ( 
.A1(n_20),
.A2(n_21),
.B1(n_71),
.B2(n_322),
.Y(n_328)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_38),
.B1(n_39),
.B2(n_70),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_22),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g22 ( 
.A1(n_23),
.A2(n_32),
.B1(n_35),
.B2(n_37),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_23),
.A2(n_37),
.B1(n_144),
.B2(n_145),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_23),
.A2(n_37),
.B1(n_145),
.B2(n_268),
.Y(n_267)
);

OAI21xp5_ASAP7_75t_SL g286 ( 
.A1(n_23),
.A2(n_268),
.B(n_287),
.Y(n_286)
);

OAI21xp5_ASAP7_75t_SL g313 ( 
.A1(n_23),
.A2(n_85),
.B(n_314),
.Y(n_313)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_24),
.B(n_73),
.Y(n_72)
);

AOI21xp5_ASAP7_75t_L g82 ( 
.A1(n_24),
.A2(n_83),
.B(n_84),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_24),
.A2(n_29),
.B1(n_131),
.B2(n_133),
.Y(n_130)
);

O2A1O1Ixp33_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_26),
.B(n_28),
.C(n_29),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_25),
.B(n_26),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_25),
.B(n_31),
.Y(n_138)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_26),
.Y(n_33)
);

HAxp5_ASAP7_75t_SL g131 ( 
.A(n_26),
.B(n_132),
.CON(n_131),
.SN(n_131)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_28),
.A2(n_30),
.B1(n_131),
.B2(n_138),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_29),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_29),
.B(n_73),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g287 ( 
.A(n_29),
.B(n_288),
.Y(n_287)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_30),
.Y(n_31)
);

AOI32xp33_ASAP7_75t_L g219 ( 
.A1(n_30),
.A2(n_46),
.A3(n_49),
.B1(n_220),
.B2(n_221),
.Y(n_219)
);

A2O1A1Ixp33_ASAP7_75t_L g54 ( 
.A1(n_31),
.A2(n_43),
.B(n_44),
.C(n_55),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_31),
.B(n_44),
.Y(n_55)
);

OAI21xp5_ASAP7_75t_L g71 ( 
.A1(n_32),
.A2(n_37),
.B(n_72),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_35),
.Y(n_83)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g39 ( 
.A1(n_40),
.A2(n_59),
.B1(n_68),
.B2(n_69),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_40),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_41),
.B(n_52),
.Y(n_40)
);

INVxp67_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

AOI21xp5_ASAP7_75t_L g147 ( 
.A1(n_42),
.A2(n_53),
.B(n_148),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_43),
.B(n_50),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_43),
.B(n_57),
.Y(n_78)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_43),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_43),
.A2(n_54),
.B1(n_126),
.B2(n_128),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_43),
.A2(n_54),
.B1(n_167),
.B2(n_224),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_L g283 ( 
.A1(n_43),
.A2(n_52),
.B(n_284),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_43),
.A2(n_54),
.B1(n_77),
.B2(n_284),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_L g43 ( 
.A1(n_44),
.A2(n_46),
.B1(n_47),
.B2(n_49),
.Y(n_43)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_44),
.Y(n_49)
);

NAND2xp33_ASAP7_75t_SL g221 ( 
.A(n_44),
.B(n_47),
.Y(n_221)
);

INVx11_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

A2O1A1Ixp33_ASAP7_75t_L g184 ( 
.A1(n_47),
.A2(n_65),
.B(n_132),
.C(n_185),
.Y(n_184)
);

INVx11_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_50),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_53),
.B(n_56),
.Y(n_52)
);

AOI21xp5_ASAP7_75t_L g75 ( 
.A1(n_53),
.A2(n_76),
.B(n_78),
.Y(n_75)
);

OAI21xp5_ASAP7_75t_SL g87 ( 
.A1(n_53),
.A2(n_88),
.B(n_89),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_53),
.A2(n_88),
.B1(n_166),
.B2(n_168),
.Y(n_165)
);

AOI21xp5_ASAP7_75t_L g270 ( 
.A1(n_53),
.A2(n_78),
.B(n_89),
.Y(n_270)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_57),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_59),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_59),
.B(n_69),
.C(n_70),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g324 ( 
.A1(n_59),
.A2(n_68),
.B1(n_75),
.B2(n_325),
.Y(n_324)
);

AOI21xp5_ASAP7_75t_SL g59 ( 
.A1(n_60),
.A2(n_62),
.B(n_66),
.Y(n_59)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_60),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_SL g121 ( 
.A1(n_60),
.A2(n_66),
.B(n_122),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_60),
.A2(n_62),
.B1(n_188),
.B2(n_189),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_60),
.A2(n_62),
.B1(n_189),
.B2(n_209),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_60),
.A2(n_62),
.B1(n_209),
.B2(n_227),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_SL g241 ( 
.A1(n_60),
.A2(n_227),
.B(n_242),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_60),
.A2(n_62),
.B1(n_114),
.B2(n_260),
.Y(n_259)
);

OAI21xp5_ASAP7_75t_SL g295 ( 
.A1(n_60),
.A2(n_122),
.B(n_260),
.Y(n_295)
);

OAI21xp5_ASAP7_75t_L g113 ( 
.A1(n_62),
.A2(n_114),
.B(n_115),
.Y(n_113)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_62),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_62),
.B(n_132),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_63),
.B(n_198),
.Y(n_197)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_67),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_67),
.B(n_123),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_68),
.B(n_71),
.C(n_75),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_71),
.A2(n_322),
.B1(n_323),
.B2(n_324),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_71),
.Y(n_322)
);

XNOR2xp5_ASAP7_75t_L g327 ( 
.A(n_74),
.B(n_328),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_75),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_77),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_80),
.A2(n_90),
.B1(n_91),
.B2(n_92),
.Y(n_79)
);

CKINVDCx14_ASAP7_75t_R g92 ( 
.A(n_80),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_81),
.A2(n_82),
.B1(n_86),
.B2(n_87),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_82),
.Y(n_81)
);

CKINVDCx16_ASAP7_75t_R g84 ( 
.A(n_85),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_87),
.Y(n_86)
);

CKINVDCx16_ASAP7_75t_R g90 ( 
.A(n_91),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

OAI321xp33_ASAP7_75t_L g95 ( 
.A1(n_96),
.A2(n_319),
.A3(n_329),
.B1(n_332),
.B2(n_333),
.C(n_336),
.Y(n_95)
);

AOI21xp5_ASAP7_75t_L g96 ( 
.A1(n_97),
.A2(n_299),
.B(n_318),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_SL g97 ( 
.A1(n_98),
.A2(n_275),
.B(n_298),
.Y(n_97)
);

O2A1O1Ixp33_ASAP7_75t_SL g98 ( 
.A1(n_99),
.A2(n_169),
.B(n_251),
.C(n_274),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_150),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_100),
.B(n_150),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_101),
.A2(n_102),
.B1(n_135),
.B2(n_149),
.Y(n_100)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_SL g102 ( 
.A(n_103),
.B(n_119),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_103),
.B(n_119),
.C(n_149),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_104),
.A2(n_105),
.B1(n_113),
.B2(n_118),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g263 ( 
.A(n_104),
.B(n_118),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_105),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_L g105 ( 
.A1(n_106),
.A2(n_108),
.B(n_109),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_106),
.A2(n_108),
.B1(n_111),
.B2(n_140),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_106),
.A2(n_161),
.B1(n_178),
.B2(n_194),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_L g210 ( 
.A1(n_106),
.A2(n_181),
.B(n_211),
.Y(n_210)
);

AOI21xp5_ASAP7_75t_L g293 ( 
.A1(n_106),
.A2(n_111),
.B(n_294),
.Y(n_293)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_107),
.B(n_163),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_107),
.A2(n_177),
.B1(n_179),
.B2(n_180),
.Y(n_176)
);

AOI21xp5_ASAP7_75t_L g218 ( 
.A1(n_107),
.A2(n_110),
.B(n_212),
.Y(n_218)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_111),
.B(n_112),
.Y(n_110)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_111),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_111),
.B(n_132),
.Y(n_198)
);

INVxp67_ASAP7_75t_L g163 ( 
.A(n_112),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_113),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_115),
.B(n_242),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_117),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_116),
.B(n_123),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_120),
.B(n_124),
.C(n_130),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_120),
.A2(n_121),
.B1(n_124),
.B2(n_125),
.Y(n_152)
);

CKINVDCx16_ASAP7_75t_R g120 ( 
.A(n_121),
.Y(n_120)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_126),
.Y(n_168)
);

CKINVDCx16_ASAP7_75t_R g148 ( 
.A(n_128),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_SL g151 ( 
.A(n_130),
.B(n_152),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_133),
.Y(n_144)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_135),
.Y(n_149)
);

XOR2xp5_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_141),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_136),
.B(n_142),
.C(n_147),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_139),
.Y(n_136)
);

XOR2xp5_ASAP7_75t_L g154 ( 
.A(n_137),
.B(n_139),
.Y(n_154)
);

OAI21x1_ASAP7_75t_SL g158 ( 
.A1(n_140),
.A2(n_159),
.B(n_162),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_142),
.A2(n_143),
.B1(n_146),
.B2(n_147),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

CKINVDCx16_ASAP7_75t_R g146 ( 
.A(n_147),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_153),
.C(n_155),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_151),
.B(n_248),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_L g248 ( 
.A1(n_153),
.A2(n_154),
.B1(n_155),
.B2(n_156),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_154),
.Y(n_153)
);

CKINVDCx16_ASAP7_75t_R g155 ( 
.A(n_156),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_164),
.C(n_165),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_157),
.A2(n_158),
.B1(n_164),
.B2(n_238),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_158),
.Y(n_157)
);

INVx4_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_160),
.B(n_212),
.Y(n_211)
);

INVx5_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_162),
.B(n_211),
.Y(n_258)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_164),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_SL g236 ( 
.A(n_165),
.B(n_237),
.Y(n_236)
);

CKINVDCx16_ASAP7_75t_R g166 ( 
.A(n_167),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_SL g169 ( 
.A(n_170),
.B(n_250),
.Y(n_169)
);

AOI21xp5_ASAP7_75t_L g170 ( 
.A1(n_171),
.A2(n_245),
.B(n_249),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_SL g171 ( 
.A1(n_172),
.A2(n_232),
.B(n_244),
.Y(n_171)
);

AOI21xp5_ASAP7_75t_L g172 ( 
.A1(n_173),
.A2(n_214),
.B(n_231),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_SL g173 ( 
.A1(n_174),
.A2(n_201),
.B(n_213),
.Y(n_173)
);

AOI21xp5_ASAP7_75t_L g174 ( 
.A1(n_175),
.A2(n_190),
.B(n_200),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_182),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_176),
.B(n_182),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_178),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_181),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_183),
.A2(n_184),
.B1(n_186),
.B2(n_187),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_184),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_SL g202 ( 
.A(n_184),
.B(n_186),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_187),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_SL g190 ( 
.A1(n_191),
.A2(n_195),
.B(n_199),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_193),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_192),
.B(n_193),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_196),
.B(n_197),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_203),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_202),
.B(n_203),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_210),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_205),
.A2(n_206),
.B1(n_207),
.B2(n_208),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_205),
.B(n_208),
.C(n_210),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_206),
.Y(n_205)
);

CKINVDCx16_ASAP7_75t_R g207 ( 
.A(n_208),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_212),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_216),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_215),
.B(n_216),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_217),
.A2(n_222),
.B1(n_229),
.B2(n_230),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_217),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_219),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_218),
.B(n_219),
.Y(n_243)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_222),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_223),
.A2(n_225),
.B1(n_226),
.B2(n_228),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_223),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_225),
.B(n_228),
.C(n_229),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_226),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_234),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_233),
.B(n_234),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_235),
.A2(n_236),
.B1(n_239),
.B2(n_240),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_235),
.B(n_241),
.C(n_243),
.Y(n_246)
);

CKINVDCx14_ASAP7_75t_R g235 ( 
.A(n_236),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_240),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_243),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_247),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_SL g249 ( 
.A(n_246),
.B(n_247),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_253),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_SL g274 ( 
.A(n_252),
.B(n_253),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_254),
.A2(n_255),
.B1(n_272),
.B2(n_273),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_L g255 ( 
.A1(n_256),
.A2(n_257),
.B1(n_261),
.B2(n_262),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_256),
.B(n_262),
.C(n_273),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_257),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_259),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_258),
.B(n_259),
.Y(n_281)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_263),
.A2(n_264),
.B1(n_265),
.B2(n_271),
.Y(n_262)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_263),
.Y(n_271)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_266),
.A2(n_267),
.B1(n_269),
.B2(n_270),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_266),
.B(n_270),
.C(n_271),
.Y(n_297)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

CKINVDCx14_ASAP7_75t_R g273 ( 
.A(n_272),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_276),
.B(n_277),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_276),
.B(n_277),
.Y(n_298)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_278),
.B(n_297),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_279),
.A2(n_280),
.B1(n_290),
.B2(n_291),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_279),
.B(n_291),
.C(n_297),
.Y(n_300)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_281),
.B(n_282),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_281),
.B(n_285),
.C(n_289),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_283),
.A2(n_285),
.B1(n_286),
.B2(n_289),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_283),
.Y(n_289)
);

CKINVDCx14_ASAP7_75t_R g285 ( 
.A(n_286),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_288),
.Y(n_314)
);

CKINVDCx14_ASAP7_75t_R g290 ( 
.A(n_291),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_L g291 ( 
.A1(n_292),
.A2(n_293),
.B1(n_295),
.B2(n_296),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g312 ( 
.A1(n_292),
.A2(n_293),
.B1(n_313),
.B2(n_315),
.Y(n_312)
);

OAI21xp5_ASAP7_75t_L g326 ( 
.A1(n_292),
.A2(n_309),
.B(n_313),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_293),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_293),
.B(n_295),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_295),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_300),
.B(n_301),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_SL g318 ( 
.A(n_300),
.B(n_301),
.Y(n_318)
);

AOI22xp33_ASAP7_75t_SL g301 ( 
.A1(n_302),
.A2(n_303),
.B1(n_316),
.B2(n_317),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

XOR2xp5_ASAP7_75t_L g303 ( 
.A(n_304),
.B(n_308),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_304),
.B(n_308),
.C(n_317),
.Y(n_330)
);

AOI21xp5_ASAP7_75t_L g304 ( 
.A1(n_305),
.A2(n_306),
.B(n_307),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_305),
.B(n_306),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_307),
.B(n_321),
.C(n_326),
.Y(n_320)
);

FAx1_ASAP7_75t_SL g331 ( 
.A(n_307),
.B(n_321),
.CI(n_326),
.CON(n_331),
.SN(n_331)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_309),
.A2(n_310),
.B1(n_311),
.B2(n_312),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_310),
.Y(n_309)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);

CKINVDCx16_ASAP7_75t_R g315 ( 
.A(n_313),
.Y(n_315)
);

CKINVDCx16_ASAP7_75t_R g317 ( 
.A(n_316),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_320),
.B(n_327),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_320),
.B(n_327),
.Y(n_333)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_330),
.B(n_331),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_SL g332 ( 
.A(n_330),
.B(n_331),
.Y(n_332)
);

BUFx24_ASAP7_75t_SL g335 ( 
.A(n_331),
.Y(n_335)
);


endmodule