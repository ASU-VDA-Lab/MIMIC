module fake_jpeg_6239_n_203 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_203);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_203;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_121;
wire n_130;
wire n_99;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_12),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_1),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_11),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_6),
.Y(n_21)
);

INVx11_ASAP7_75t_SL g22 ( 
.A(n_1),
.Y(n_22)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_13),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_7),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_18),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_31),
.B(n_38),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_18),
.Y(n_32)
);

INVx11_ASAP7_75t_L g51 ( 
.A(n_32),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_18),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_33),
.Y(n_53)
);

INVx11_ASAP7_75t_L g34 ( 
.A(n_26),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_34),
.A2(n_35),
.B1(n_27),
.B2(n_23),
.Y(n_45)
);

INVx11_ASAP7_75t_L g35 ( 
.A(n_26),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_22),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_36),
.Y(n_43)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_22),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_37),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_19),
.B(n_0),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_15),
.Y(n_39)
);

INVx5_ASAP7_75t_L g60 ( 
.A(n_39),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_16),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_40),
.B(n_41),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_16),
.Y(n_41)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_37),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_42),
.B(n_45),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_38),
.B(n_30),
.Y(n_46)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_46),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_34),
.A2(n_27),
.B1(n_20),
.B2(n_23),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_47),
.A2(n_27),
.B1(n_23),
.B2(n_29),
.Y(n_63)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_48),
.Y(n_70)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_39),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_50),
.Y(n_64)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

INVx1_ASAP7_75t_SL g76 ( 
.A(n_52),
.Y(n_76)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_54),
.Y(n_71)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_36),
.Y(n_56)
);

INVx6_ASAP7_75t_SL g75 ( 
.A(n_56),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_40),
.B(n_41),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_57),
.B(n_59),
.Y(n_68)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_36),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_58),
.B(n_36),
.Y(n_65)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_36),
.Y(n_59)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_49),
.B(n_41),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_61),
.B(n_66),
.Y(n_87)
);

OAI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_55),
.A2(n_35),
.B1(n_34),
.B2(n_20),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_L g88 ( 
.A1(n_62),
.A2(n_60),
.B1(n_51),
.B2(n_35),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_63),
.A2(n_77),
.B1(n_66),
.B2(n_61),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_65),
.B(n_74),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_49),
.B(n_40),
.Y(n_66)
);

OR2x2_ASAP7_75t_SL g69 ( 
.A(n_55),
.B(n_24),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_69),
.B(n_77),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_43),
.B(n_31),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_73),
.B(n_48),
.Y(n_90)
);

OR2x2_ASAP7_75t_L g74 ( 
.A(n_43),
.B(n_17),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_60),
.B(n_28),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_69),
.B(n_25),
.Y(n_79)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_79),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_72),
.A2(n_51),
.B1(n_42),
.B2(n_52),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_80),
.A2(n_29),
.B1(n_17),
.B2(n_53),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_63),
.A2(n_34),
.B1(n_35),
.B2(n_50),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_82),
.A2(n_95),
.B1(n_76),
.B2(n_70),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_83),
.A2(n_91),
.B1(n_15),
.B2(n_26),
.Y(n_113)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_73),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_84),
.B(n_85),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_74),
.Y(n_85)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_75),
.Y(n_86)
);

INVx13_ASAP7_75t_L g97 ( 
.A(n_86),
.Y(n_97)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_88),
.Y(n_100)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_75),
.Y(n_89)
);

INVx13_ASAP7_75t_L g110 ( 
.A(n_89),
.Y(n_110)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_90),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_L g91 ( 
.A1(n_61),
.A2(n_54),
.B1(n_24),
.B2(n_30),
.Y(n_91)
);

XNOR2xp5_ASAP7_75t_L g92 ( 
.A(n_66),
.B(n_33),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_92),
.B(n_94),
.C(n_67),
.Y(n_103)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_71),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_93),
.B(n_36),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_65),
.B(n_31),
.C(n_32),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_68),
.A2(n_59),
.B1(n_56),
.B2(n_25),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_L g96 ( 
.A1(n_87),
.A2(n_77),
.B(n_21),
.Y(n_96)
);

AOI21xp5_ASAP7_75t_L g129 ( 
.A1(n_96),
.A2(n_44),
.B(n_15),
.Y(n_129)
);

AOI21xp5_ASAP7_75t_SL g98 ( 
.A1(n_84),
.A2(n_70),
.B(n_19),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_L g117 ( 
.A1(n_98),
.A2(n_87),
.B(n_78),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_101),
.B(n_109),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_82),
.A2(n_71),
.B1(n_76),
.B2(n_67),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_102),
.A2(n_113),
.B1(n_89),
.B2(n_86),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_103),
.B(n_105),
.C(n_83),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_85),
.B(n_28),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_104),
.B(n_107),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_94),
.B(n_58),
.C(n_32),
.Y(n_105)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_106),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_81),
.B(n_21),
.Y(n_107)
);

OA21x2_ASAP7_75t_L g109 ( 
.A1(n_90),
.A2(n_53),
.B(n_33),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_111),
.B(n_15),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_114),
.B(n_125),
.C(n_100),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_108),
.B(n_92),
.Y(n_116)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_116),
.Y(n_142)
);

AOI21xp5_ASAP7_75t_L g146 ( 
.A1(n_117),
.A2(n_131),
.B(n_26),
.Y(n_146)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_98),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_118),
.B(n_119),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g119 ( 
.A(n_112),
.B(n_95),
.Y(n_119)
);

CKINVDCx16_ASAP7_75t_R g120 ( 
.A(n_106),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_120),
.B(n_123),
.Y(n_138)
);

NOR3xp33_ASAP7_75t_L g121 ( 
.A(n_105),
.B(n_78),
.C(n_12),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_121),
.B(n_122),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_98),
.B(n_93),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_108),
.B(n_103),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_124),
.B(n_58),
.Y(n_140)
);

XOR2xp5_ASAP7_75t_L g125 ( 
.A(n_113),
.B(n_33),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_128),
.B(n_64),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_129),
.B(n_130),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_97),
.B(n_64),
.Y(n_130)
);

AOI32xp33_ASAP7_75t_L g131 ( 
.A1(n_101),
.A2(n_96),
.A3(n_109),
.B1(n_102),
.B2(n_111),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_132),
.B(n_139),
.C(n_143),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g135 ( 
.A(n_116),
.B(n_109),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_135),
.B(n_136),
.Y(n_160)
);

AOI322xp5_ASAP7_75t_L g136 ( 
.A1(n_117),
.A2(n_100),
.A3(n_107),
.B1(n_99),
.B2(n_104),
.C1(n_109),
.C2(n_32),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_114),
.B(n_99),
.C(n_110),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_140),
.B(n_115),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_123),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_141),
.B(n_0),
.Y(n_159)
);

XOR2xp5_ASAP7_75t_L g143 ( 
.A(n_124),
.B(n_110),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_144),
.B(n_97),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_120),
.B(n_110),
.C(n_97),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_145),
.B(n_147),
.C(n_129),
.Y(n_156)
);

AOI21xp5_ASAP7_75t_L g152 ( 
.A1(n_146),
.A2(n_126),
.B(n_133),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_115),
.B(n_125),
.C(n_118),
.Y(n_147)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_148),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_149),
.B(n_151),
.Y(n_166)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_138),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_150),
.B(n_153),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_145),
.B(n_122),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_L g173 ( 
.A1(n_152),
.A2(n_156),
.B(n_161),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_134),
.Y(n_153)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_137),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_155),
.B(n_158),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_156),
.B(n_161),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_147),
.A2(n_131),
.B1(n_119),
.B2(n_127),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_157),
.A2(n_139),
.B1(n_44),
.B2(n_2),
.Y(n_170)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_143),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_159),
.B(n_0),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_132),
.B(n_58),
.C(n_44),
.Y(n_161)
);

INVxp67_ASAP7_75t_SL g162 ( 
.A(n_148),
.Y(n_162)
);

AOI21xp5_ASAP7_75t_L g182 ( 
.A1(n_162),
.A2(n_3),
.B(n_4),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_157),
.B(n_135),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_167),
.B(n_168),
.C(n_169),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_SL g168 ( 
.A(n_160),
.B(n_146),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_SL g169 ( 
.A(n_160),
.B(n_142),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_170),
.B(n_154),
.C(n_2),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_SL g180 ( 
.A(n_172),
.B(n_1),
.Y(n_180)
);

AO21x1_ASAP7_75t_L g179 ( 
.A1(n_173),
.A2(n_44),
.B(n_2),
.Y(n_179)
);

OR2x2_ASAP7_75t_L g175 ( 
.A(n_162),
.B(n_152),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_175),
.B(n_5),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_176),
.B(n_177),
.C(n_178),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_L g177 ( 
.A1(n_164),
.A2(n_171),
.B(n_166),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_L g178 ( 
.A1(n_163),
.A2(n_154),
.B(n_165),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_179),
.B(n_181),
.C(n_4),
.Y(n_186)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_180),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_169),
.B(n_3),
.C(n_4),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_182),
.B(n_5),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_174),
.A2(n_173),
.B1(n_168),
.B2(n_6),
.Y(n_183)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_183),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_SL g193 ( 
.A(n_186),
.B(n_7),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_182),
.B(n_5),
.C(n_7),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_187),
.B(n_189),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_188),
.Y(n_192)
);

INVxp67_ASAP7_75t_L g191 ( 
.A(n_188),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_SL g199 ( 
.A1(n_191),
.A2(n_195),
.B(n_10),
.Y(n_199)
);

INVxp67_ASAP7_75t_L g196 ( 
.A(n_193),
.Y(n_196)
);

AOI21xp5_ASAP7_75t_SL g195 ( 
.A1(n_185),
.A2(n_8),
.B(n_9),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_194),
.A2(n_184),
.B1(n_10),
.B2(n_11),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_197),
.B(n_198),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_190),
.B(n_8),
.Y(n_198)
);

O2A1O1Ixp33_ASAP7_75t_L g200 ( 
.A1(n_199),
.A2(n_191),
.B(n_192),
.C(n_10),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_200),
.B(n_196),
.Y(n_202)
);

OR2x2_ASAP7_75t_L g203 ( 
.A(n_202),
.B(n_201),
.Y(n_203)
);


endmodule