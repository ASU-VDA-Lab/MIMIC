module real_jpeg_12611_n_6 (n_5, n_4, n_0, n_1, n_2, n_3, n_6);

input n_5;
input n_4;
input n_0;
input n_1;
input n_2;
input n_3;

output n_6;

wire n_17;
wire n_8;
wire n_21;
wire n_10;
wire n_9;
wire n_12;
wire n_24;
wire n_23;
wire n_11;
wire n_14;
wire n_25;
wire n_7;
wire n_22;
wire n_18;
wire n_27;
wire n_26;
wire n_20;
wire n_19;
wire n_16;
wire n_15;
wire n_13;

OAI331xp33_ASAP7_75t_L g7 ( 
.A1(n_0),
.A2(n_2),
.A3(n_5),
.B1(n_8),
.B2(n_15),
.B3(n_16),
.C1(n_21),
.Y(n_7)
);

AO21x1_ASAP7_75t_L g10 ( 
.A1(n_0),
.A2(n_11),
.B(n_12),
.Y(n_10)
);

NOR2xp33_ASAP7_75t_L g12 ( 
.A(n_0),
.B(n_11),
.Y(n_12)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_0),
.A2(n_12),
.B1(n_22),
.B2(n_27),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_1),
.Y(n_14)
);

AND2x2_ASAP7_75t_L g15 ( 
.A(n_1),
.B(n_3),
.Y(n_15)
);

OAI22xp5_ASAP7_75t_SL g25 ( 
.A1(n_1),
.A2(n_4),
.B1(n_14),
.B2(n_26),
.Y(n_25)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_2),
.B(n_5),
.Y(n_23)
);

AOI21xp5_ASAP7_75t_L g8 ( 
.A1(n_3),
.A2(n_9),
.B(n_13),
.Y(n_8)
);

OAI21xp5_ASAP7_75t_SL g19 ( 
.A1(n_3),
.A2(n_14),
.B(n_20),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_3),
.B(n_14),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_4),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_5),
.Y(n_11)
);

INVx1_ASAP7_75t_L g6 ( 
.A(n_7),
.Y(n_6)
);

CKINVDCx20_ASAP7_75t_R g9 ( 
.A(n_10),
.Y(n_9)
);

NOR2xp33_ASAP7_75t_SL g13 ( 
.A(n_10),
.B(n_14),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_11),
.B(n_25),
.Y(n_24)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_19),
.Y(n_17)
);

OAI21xp33_ASAP7_75t_SL g22 ( 
.A1(n_19),
.A2(n_23),
.B(n_24),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_25),
.Y(n_27)
);


endmodule