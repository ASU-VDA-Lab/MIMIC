module fake_jpeg_13953_n_561 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_561);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_561;

wire n_529;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_511;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx11_ASAP7_75t_L g19 ( 
.A(n_16),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_14),
.Y(n_20)
);

CKINVDCx16_ASAP7_75t_R g21 ( 
.A(n_8),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_14),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_16),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_17),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_1),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_17),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_17),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_12),
.Y(n_35)
);

INVx2_ASAP7_75t_SL g36 ( 
.A(n_13),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_11),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_1),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_0),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_11),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_16),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_0),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_8),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_12),
.Y(n_44)
);

BUFx24_ASAP7_75t_L g45 ( 
.A(n_7),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_4),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_3),
.Y(n_47)
);

BUFx5_ASAP7_75t_L g48 ( 
.A(n_16),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_14),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_10),
.Y(n_50)
);

BUFx5_ASAP7_75t_L g51 ( 
.A(n_13),
.Y(n_51)
);

INVx13_ASAP7_75t_L g52 ( 
.A(n_8),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_31),
.Y(n_53)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_53),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_54),
.Y(n_107)
);

INVx3_ASAP7_75t_SL g55 ( 
.A(n_45),
.Y(n_55)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_55),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g56 ( 
.A(n_20),
.B(n_8),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_56),
.B(n_89),
.Y(n_111)
);

BUFx8_ASAP7_75t_L g57 ( 
.A(n_45),
.Y(n_57)
);

BUFx2_ASAP7_75t_SL g135 ( 
.A(n_57),
.Y(n_135)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_26),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_58),
.Y(n_154)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_33),
.Y(n_59)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_59),
.Y(n_120)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_33),
.Y(n_60)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_60),
.Y(n_123)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_31),
.Y(n_61)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_61),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_38),
.Y(n_62)
);

BUFx2_ASAP7_75t_L g144 ( 
.A(n_62),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_38),
.Y(n_63)
);

INVx5_ASAP7_75t_L g140 ( 
.A(n_63),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_26),
.Y(n_64)
);

INVx5_ASAP7_75t_L g145 ( 
.A(n_64),
.Y(n_145)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_29),
.Y(n_65)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_65),
.Y(n_110)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_48),
.Y(n_66)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_66),
.Y(n_122)
);

BUFx12f_ASAP7_75t_L g67 ( 
.A(n_48),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g147 ( 
.A(n_67),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_26),
.Y(n_68)
);

INVx5_ASAP7_75t_L g164 ( 
.A(n_68),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_27),
.Y(n_69)
);

INVx4_ASAP7_75t_L g117 ( 
.A(n_69),
.Y(n_117)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_48),
.Y(n_70)
);

INVx3_ASAP7_75t_L g168 ( 
.A(n_70),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_27),
.Y(n_71)
);

INVx4_ASAP7_75t_L g126 ( 
.A(n_71),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_27),
.Y(n_72)
);

INVx4_ASAP7_75t_L g128 ( 
.A(n_72),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_20),
.B(n_9),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_73),
.B(n_74),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_22),
.B(n_43),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_51),
.Y(n_75)
);

INVx4_ASAP7_75t_L g151 ( 
.A(n_75),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_22),
.B(n_9),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_76),
.B(n_84),
.Y(n_121)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_37),
.Y(n_77)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_77),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_37),
.Y(n_78)
);

INVx4_ASAP7_75t_L g163 ( 
.A(n_78),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_37),
.Y(n_79)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_79),
.Y(n_143)
);

BUFx5_ASAP7_75t_L g80 ( 
.A(n_51),
.Y(n_80)
);

BUFx8_ASAP7_75t_L g166 ( 
.A(n_80),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_40),
.B(n_9),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_81),
.B(n_21),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_41),
.Y(n_82)
);

INVx3_ASAP7_75t_L g160 ( 
.A(n_82),
.Y(n_160)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_40),
.Y(n_83)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_83),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_43),
.B(n_9),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_41),
.Y(n_85)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_85),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_41),
.Y(n_86)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_86),
.Y(n_139)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_30),
.Y(n_87)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_87),
.Y(n_148)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_34),
.Y(n_88)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_88),
.Y(n_119)
);

CKINVDCx16_ASAP7_75t_R g89 ( 
.A(n_45),
.Y(n_89)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_51),
.Y(n_90)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_90),
.Y(n_149)
);

BUFx3_ASAP7_75t_L g91 ( 
.A(n_25),
.Y(n_91)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_91),
.Y(n_159)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_42),
.Y(n_92)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_92),
.Y(n_130)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_30),
.Y(n_93)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_93),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_32),
.Y(n_94)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_94),
.Y(n_142)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_32),
.Y(n_95)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_95),
.Y(n_155)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_32),
.Y(n_96)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_96),
.Y(n_165)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_30),
.Y(n_97)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_97),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_49),
.B(n_7),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g129 ( 
.A(n_98),
.B(n_17),
.Y(n_129)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_34),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_99),
.B(n_101),
.Y(n_112)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_42),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_100),
.B(n_103),
.Y(n_116)
);

CKINVDCx16_ASAP7_75t_R g101 ( 
.A(n_45),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_35),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_102),
.B(n_105),
.Y(n_125)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_29),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_39),
.Y(n_104)
);

NOR3xp33_ASAP7_75t_L g124 ( 
.A(n_104),
.B(n_19),
.C(n_21),
.Y(n_124)
);

INVx5_ASAP7_75t_L g105 ( 
.A(n_29),
.Y(n_105)
);

AND2x4_ASAP7_75t_SL g108 ( 
.A(n_92),
.B(n_45),
.Y(n_108)
);

AND2x2_ASAP7_75t_L g207 ( 
.A(n_108),
.B(n_113),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_65),
.B(n_103),
.C(n_104),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_115),
.B(n_124),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_100),
.B(n_49),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_SL g177 ( 
.A(n_127),
.B(n_129),
.Y(n_177)
);

NAND2xp67_ASAP7_75t_SL g132 ( 
.A(n_57),
.B(n_19),
.Y(n_132)
);

AND2x2_ASAP7_75t_L g212 ( 
.A(n_132),
.B(n_133),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_94),
.B(n_23),
.C(n_24),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_67),
.B(n_35),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g214 ( 
.A(n_134),
.B(n_137),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_67),
.B(n_44),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_105),
.B(n_44),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_SL g216 ( 
.A(n_141),
.B(n_152),
.Y(n_216)
);

AOI22xp33_ASAP7_75t_L g146 ( 
.A1(n_58),
.A2(n_36),
.B1(n_28),
.B2(n_24),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_146),
.A2(n_156),
.B1(n_79),
.B2(n_78),
.Y(n_189)
);

A2O1A1Ixp33_ASAP7_75t_L g150 ( 
.A1(n_57),
.A2(n_23),
.B(n_19),
.C(n_52),
.Y(n_150)
);

AOI32xp33_ASAP7_75t_L g197 ( 
.A1(n_150),
.A2(n_50),
.A3(n_46),
.B1(n_29),
.B2(n_52),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_77),
.B(n_28),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_L g156 ( 
.A1(n_54),
.A2(n_36),
.B1(n_39),
.B2(n_47),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_62),
.A2(n_36),
.B1(n_39),
.B2(n_52),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_157),
.A2(n_55),
.B1(n_42),
.B2(n_47),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_75),
.B(n_47),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_158),
.B(n_162),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_63),
.B(n_36),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_161),
.B(n_47),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_91),
.B(n_47),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_169),
.A2(n_174),
.B1(n_189),
.B2(n_201),
.Y(n_238)
);

HB1xp67_ASAP7_75t_L g170 ( 
.A(n_155),
.Y(n_170)
);

HB1xp67_ASAP7_75t_L g243 ( 
.A(n_170),
.Y(n_243)
);

AOI22xp33_ASAP7_75t_SL g171 ( 
.A1(n_132),
.A2(n_70),
.B1(n_50),
.B2(n_46),
.Y(n_171)
);

CKINVDCx16_ASAP7_75t_R g268 ( 
.A(n_171),
.Y(n_268)
);

AND2x2_ASAP7_75t_L g264 ( 
.A(n_172),
.B(n_173),
.Y(n_264)
);

AND2x2_ASAP7_75t_SL g173 ( 
.A(n_108),
.B(n_42),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_156),
.A2(n_86),
.B1(n_85),
.B2(n_82),
.Y(n_174)
);

INVx4_ASAP7_75t_L g175 ( 
.A(n_110),
.Y(n_175)
);

INVx3_ASAP7_75t_L g276 ( 
.A(n_175),
.Y(n_276)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_136),
.Y(n_176)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_176),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_125),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_178),
.B(n_196),
.Y(n_259)
);

AOI22xp33_ASAP7_75t_SL g179 ( 
.A1(n_109),
.A2(n_29),
.B1(n_46),
.B2(n_50),
.Y(n_179)
);

OR2x2_ASAP7_75t_L g254 ( 
.A(n_179),
.B(n_209),
.Y(n_254)
);

INVx6_ASAP7_75t_L g180 ( 
.A(n_107),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g232 ( 
.A(n_180),
.Y(n_232)
);

INVx2_ASAP7_75t_SL g181 ( 
.A(n_142),
.Y(n_181)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_181),
.Y(n_231)
);

BUFx3_ASAP7_75t_L g182 ( 
.A(n_147),
.Y(n_182)
);

INVx1_ASAP7_75t_SL g236 ( 
.A(n_182),
.Y(n_236)
);

INVx3_ASAP7_75t_L g183 ( 
.A(n_110),
.Y(n_183)
);

INVx1_ASAP7_75t_SL g256 ( 
.A(n_183),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_133),
.B(n_42),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_184),
.B(n_200),
.Y(n_252)
);

INVx5_ASAP7_75t_L g185 ( 
.A(n_151),
.Y(n_185)
);

HB1xp67_ASAP7_75t_L g257 ( 
.A(n_185),
.Y(n_257)
);

INVx4_ASAP7_75t_L g186 ( 
.A(n_168),
.Y(n_186)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_186),
.Y(n_282)
);

BUFx6f_ASAP7_75t_L g187 ( 
.A(n_107),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g258 ( 
.A(n_187),
.Y(n_258)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_136),
.Y(n_188)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_188),
.Y(n_242)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_153),
.Y(n_190)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_190),
.Y(n_246)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_153),
.Y(n_191)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_191),
.Y(n_249)
);

INVx4_ASAP7_75t_L g193 ( 
.A(n_168),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g267 ( 
.A(n_193),
.Y(n_267)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_114),
.Y(n_194)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_194),
.Y(n_255)
);

INVx3_ASAP7_75t_L g195 ( 
.A(n_151),
.Y(n_195)
);

BUFx6f_ASAP7_75t_L g271 ( 
.A(n_195),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_112),
.Y(n_196)
);

OAI21xp33_ASAP7_75t_SL g239 ( 
.A1(n_197),
.A2(n_206),
.B(n_140),
.Y(n_239)
);

BUFx2_ASAP7_75t_L g198 ( 
.A(n_109),
.Y(n_198)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_198),
.Y(n_281)
);

INVx8_ASAP7_75t_L g199 ( 
.A(n_154),
.Y(n_199)
);

INVx4_ASAP7_75t_SL g235 ( 
.A(n_199),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_118),
.B(n_0),
.Y(n_200)
);

OAI22xp33_ASAP7_75t_SL g201 ( 
.A1(n_157),
.A2(n_72),
.B1(n_71),
.B2(n_69),
.Y(n_201)
);

BUFx2_ASAP7_75t_L g202 ( 
.A(n_145),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_202),
.B(n_204),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_121),
.A2(n_146),
.B1(n_106),
.B2(n_111),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_203),
.A2(n_219),
.B1(n_227),
.B2(n_228),
.Y(n_244)
);

BUFx6f_ASAP7_75t_L g204 ( 
.A(n_154),
.Y(n_204)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_139),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_205),
.B(n_222),
.Y(n_275)
);

AOI22xp33_ASAP7_75t_L g206 ( 
.A1(n_144),
.A2(n_68),
.B1(n_64),
.B2(n_50),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_119),
.B(n_0),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_208),
.B(n_210),
.Y(n_279)
);

AOI22xp33_ASAP7_75t_SL g209 ( 
.A1(n_150),
.A2(n_50),
.B1(n_46),
.B2(n_25),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_120),
.B(n_1),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_165),
.B(n_46),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_SL g234 ( 
.A(n_211),
.B(n_217),
.Y(n_234)
);

INVx5_ASAP7_75t_SL g213 ( 
.A(n_135),
.Y(n_213)
);

OR2x2_ASAP7_75t_L g260 ( 
.A(n_213),
.B(n_221),
.Y(n_260)
);

AO22x1_ASAP7_75t_L g215 ( 
.A1(n_108),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_215)
);

AOI21xp5_ASAP7_75t_SL g278 ( 
.A1(n_215),
.A2(n_2),
.B(n_12),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_167),
.B(n_10),
.Y(n_217)
);

AO22x1_ASAP7_75t_SL g218 ( 
.A1(n_123),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_218),
.A2(n_144),
.B1(n_140),
.B2(n_128),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_L g219 ( 
.A1(n_113),
.A2(n_10),
.B1(n_4),
.B2(n_5),
.Y(n_219)
);

BUFx4f_ASAP7_75t_L g220 ( 
.A(n_145),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_220),
.Y(n_237)
);

AOI22xp33_ASAP7_75t_SL g221 ( 
.A1(n_159),
.A2(n_10),
.B1(n_4),
.B2(n_5),
.Y(n_221)
);

BUFx2_ASAP7_75t_L g222 ( 
.A(n_164),
.Y(n_222)
);

INVx4_ASAP7_75t_L g223 ( 
.A(n_147),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_223),
.B(n_116),
.Y(n_262)
);

INVx3_ASAP7_75t_L g224 ( 
.A(n_164),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_224),
.Y(n_241)
);

AOI22xp33_ASAP7_75t_SL g226 ( 
.A1(n_122),
.A2(n_11),
.B1(n_5),
.B2(n_6),
.Y(n_226)
);

OAI22xp33_ASAP7_75t_SL g248 ( 
.A1(n_226),
.A2(n_215),
.B1(n_198),
.B2(n_222),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_L g227 ( 
.A1(n_138),
.A2(n_11),
.B1(n_5),
.B2(n_6),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_148),
.A2(n_2),
.B1(n_18),
.B2(n_7),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_130),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_229),
.B(n_117),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_230),
.A2(n_233),
.B1(n_253),
.B2(n_274),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_L g233 ( 
.A1(n_184),
.A2(n_160),
.B1(n_143),
.B2(n_126),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g332 ( 
.A1(n_239),
.A2(n_260),
.B1(n_241),
.B2(n_256),
.Y(n_332)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_172),
.B(n_131),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_240),
.B(n_176),
.C(n_205),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_213),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_245),
.B(n_247),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_200),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_248),
.A2(n_261),
.B1(n_202),
.B2(n_195),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_208),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_250),
.B(n_265),
.Y(n_315)
);

AOI22xp33_ASAP7_75t_L g251 ( 
.A1(n_174),
.A2(n_143),
.B1(n_160),
.B2(n_163),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_L g288 ( 
.A1(n_251),
.A2(n_272),
.B1(n_215),
.B2(n_181),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_207),
.A2(n_163),
.B1(n_128),
.B2(n_126),
.Y(n_253)
);

OAI22xp33_ASAP7_75t_SL g261 ( 
.A1(n_212),
.A2(n_122),
.B1(n_117),
.B2(n_149),
.Y(n_261)
);

INVxp67_ASAP7_75t_L g285 ( 
.A(n_262),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_SL g263 ( 
.A(n_177),
.B(n_116),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_SL g287 ( 
.A(n_263),
.B(n_269),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_SL g269 ( 
.A(n_216),
.B(n_13),
.Y(n_269)
);

AOI21xp5_ASAP7_75t_L g270 ( 
.A1(n_207),
.A2(n_166),
.B(n_6),
.Y(n_270)
);

AOI21xp5_ASAP7_75t_L g296 ( 
.A1(n_270),
.A2(n_283),
.B(n_272),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_212),
.A2(n_166),
.B1(n_6),
.B2(n_7),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_207),
.A2(n_166),
.B1(n_2),
.B2(n_15),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_181),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_277),
.B(n_190),
.Y(n_316)
);

OAI21xp5_ASAP7_75t_L g291 ( 
.A1(n_278),
.A2(n_228),
.B(n_218),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_L g280 ( 
.A1(n_210),
.A2(n_15),
.B1(n_18),
.B2(n_192),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g325 ( 
.A1(n_280),
.A2(n_230),
.B1(n_237),
.B2(n_245),
.Y(n_325)
);

A2O1A1Ixp33_ASAP7_75t_L g283 ( 
.A1(n_212),
.A2(n_15),
.B(n_18),
.C(n_173),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_283),
.B(n_218),
.Y(n_304)
);

AND2x2_ASAP7_75t_SL g284 ( 
.A(n_252),
.B(n_173),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g342 ( 
.A(n_284),
.B(n_303),
.Y(n_342)
);

MAJx2_ASAP7_75t_L g286 ( 
.A(n_264),
.B(n_225),
.C(n_194),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_286),
.B(n_321),
.C(n_328),
.Y(n_338)
);

AOI22xp5_ASAP7_75t_L g344 ( 
.A1(n_288),
.A2(n_310),
.B1(n_320),
.B2(n_324),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_SL g289 ( 
.A(n_247),
.B(n_250),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_289),
.B(n_294),
.Y(n_339)
);

AOI22xp33_ASAP7_75t_SL g290 ( 
.A1(n_253),
.A2(n_193),
.B1(n_186),
.B2(n_169),
.Y(n_290)
);

AOI22xp33_ASAP7_75t_SL g345 ( 
.A1(n_290),
.A2(n_256),
.B1(n_237),
.B2(n_236),
.Y(n_345)
);

OAI21xp5_ASAP7_75t_L g337 ( 
.A1(n_291),
.A2(n_296),
.B(n_311),
.Y(n_337)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_242),
.Y(n_292)
);

INVx2_ASAP7_75t_L g346 ( 
.A(n_292),
.Y(n_346)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_255),
.Y(n_293)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_293),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_279),
.B(n_214),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_255),
.Y(n_295)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_295),
.Y(n_352)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_231),
.Y(n_297)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_297),
.Y(n_359)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_231),
.Y(n_298)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_298),
.Y(n_369)
);

INVxp33_ASAP7_75t_L g341 ( 
.A(n_299),
.Y(n_341)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_246),
.Y(n_300)
);

INVx2_ASAP7_75t_L g347 ( 
.A(n_300),
.Y(n_347)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_246),
.Y(n_301)
);

INVx2_ASAP7_75t_L g365 ( 
.A(n_301),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_SL g302 ( 
.A(n_279),
.B(n_229),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_302),
.B(n_312),
.Y(n_340)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_249),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_SL g354 ( 
.A(n_304),
.B(n_308),
.Y(n_354)
);

INVxp67_ASAP7_75t_L g305 ( 
.A(n_270),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g370 ( 
.A(n_305),
.B(n_309),
.Y(n_370)
);

XNOR2xp5_ASAP7_75t_L g306 ( 
.A(n_240),
.B(n_183),
.Y(n_306)
);

XNOR2x1_ASAP7_75t_L g364 ( 
.A(n_306),
.B(n_319),
.Y(n_364)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_249),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_234),
.B(n_175),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_L g310 ( 
.A1(n_238),
.A2(n_199),
.B1(n_180),
.B2(n_204),
.Y(n_310)
);

OAI21xp5_ASAP7_75t_L g311 ( 
.A1(n_278),
.A2(n_182),
.B(n_224),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_252),
.B(n_188),
.Y(n_312)
);

INVxp67_ASAP7_75t_L g313 ( 
.A(n_243),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_313),
.B(n_314),
.Y(n_372)
);

INVxp67_ASAP7_75t_L g314 ( 
.A(n_274),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_SL g362 ( 
.A(n_316),
.B(n_317),
.Y(n_362)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_242),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_SL g320 ( 
.A1(n_238),
.A2(n_191),
.B1(n_187),
.B2(n_185),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_264),
.B(n_223),
.C(n_220),
.Y(n_321)
);

AO22x1_ASAP7_75t_L g322 ( 
.A1(n_233),
.A2(n_220),
.B1(n_15),
.B2(n_18),
.Y(n_322)
);

OA21x2_ASAP7_75t_L g357 ( 
.A1(n_322),
.A2(n_281),
.B(n_282),
.Y(n_357)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_266),
.Y(n_323)
);

INVx3_ASAP7_75t_L g371 ( 
.A(n_323),
.Y(n_371)
);

OAI22xp5_ASAP7_75t_SL g324 ( 
.A1(n_244),
.A2(n_254),
.B1(n_268),
.B2(n_260),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_325),
.B(n_326),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_280),
.B(n_264),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_L g327 ( 
.A1(n_268),
.A2(n_244),
.B1(n_254),
.B2(n_234),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_L g336 ( 
.A1(n_327),
.A2(n_332),
.B1(n_328),
.B2(n_318),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_254),
.B(n_259),
.C(n_265),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_SL g329 ( 
.A(n_277),
.B(n_263),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_329),
.B(n_331),
.Y(n_363)
);

OAI21xp5_ASAP7_75t_L g330 ( 
.A1(n_260),
.A2(n_269),
.B(n_275),
.Y(n_330)
);

OAI21xp5_ASAP7_75t_L g350 ( 
.A1(n_330),
.A2(n_273),
.B(n_236),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_275),
.B(n_241),
.Y(n_331)
);

AND2x2_ASAP7_75t_SL g335 ( 
.A(n_332),
.B(n_276),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_316),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g394 ( 
.A(n_333),
.B(n_349),
.Y(n_394)
);

CKINVDCx14_ASAP7_75t_R g410 ( 
.A(n_335),
.Y(n_410)
);

AOI22xp5_ASAP7_75t_L g376 ( 
.A1(n_336),
.A2(n_348),
.B1(n_357),
.B2(n_361),
.Y(n_376)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_284),
.B(n_257),
.C(n_281),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g377 ( 
.A(n_343),
.B(n_366),
.C(n_367),
.Y(n_377)
);

AOI21xp5_ASAP7_75t_L g391 ( 
.A1(n_345),
.A2(n_351),
.B(n_358),
.Y(n_391)
);

OAI22xp5_ASAP7_75t_SL g348 ( 
.A1(n_327),
.A2(n_273),
.B1(n_232),
.B2(n_258),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g349 ( 
.A(n_331),
.Y(n_349)
);

XOR2xp5_ASAP7_75t_L g396 ( 
.A(n_350),
.B(n_301),
.Y(n_396)
);

AOI21xp5_ASAP7_75t_L g351 ( 
.A1(n_311),
.A2(n_299),
.B(n_307),
.Y(n_351)
);

INVx4_ASAP7_75t_L g355 ( 
.A(n_323),
.Y(n_355)
);

INVx2_ASAP7_75t_L g406 ( 
.A(n_355),
.Y(n_406)
);

CKINVDCx16_ASAP7_75t_R g356 ( 
.A(n_307),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_L g395 ( 
.A(n_356),
.B(n_297),
.Y(n_395)
);

AOI21xp5_ASAP7_75t_L g358 ( 
.A1(n_291),
.A2(n_276),
.B(n_282),
.Y(n_358)
);

AOI22xp33_ASAP7_75t_SL g360 ( 
.A1(n_324),
.A2(n_267),
.B1(n_271),
.B2(n_235),
.Y(n_360)
);

BUFx3_ASAP7_75t_L g380 ( 
.A(n_360),
.Y(n_380)
);

OAI22xp5_ASAP7_75t_SL g361 ( 
.A1(n_318),
.A2(n_232),
.B1(n_258),
.B2(n_267),
.Y(n_361)
);

XOR2xp5_ASAP7_75t_L g366 ( 
.A(n_284),
.B(n_306),
.Y(n_366)
);

MAJIxp5_ASAP7_75t_L g367 ( 
.A(n_284),
.B(n_266),
.C(n_271),
.Y(n_367)
);

OAI22xp5_ASAP7_75t_L g368 ( 
.A1(n_325),
.A2(n_232),
.B1(n_258),
.B2(n_267),
.Y(n_368)
);

AOI22xp5_ASAP7_75t_L g385 ( 
.A1(n_368),
.A2(n_373),
.B1(n_320),
.B2(n_310),
.Y(n_385)
);

OAI22xp5_ASAP7_75t_SL g373 ( 
.A1(n_289),
.A2(n_235),
.B1(n_271),
.B2(n_326),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_302),
.B(n_235),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_374),
.B(n_375),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_312),
.B(n_315),
.Y(n_375)
);

AOI22x1_ASAP7_75t_SL g378 ( 
.A1(n_337),
.A2(n_348),
.B1(n_373),
.B2(n_351),
.Y(n_378)
);

AOI21xp5_ASAP7_75t_L g416 ( 
.A1(n_378),
.A2(n_342),
.B(n_338),
.Y(n_416)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_347),
.Y(n_381)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_381),
.Y(n_425)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_347),
.Y(n_382)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_382),
.Y(n_431)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_365),
.Y(n_383)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_383),
.Y(n_437)
);

CKINVDCx20_ASAP7_75t_R g384 ( 
.A(n_362),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_L g443 ( 
.A(n_384),
.B(n_404),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_385),
.B(n_388),
.Y(n_413)
);

OAI22xp5_ASAP7_75t_SL g386 ( 
.A1(n_353),
.A2(n_304),
.B1(n_315),
.B2(n_296),
.Y(n_386)
);

AOI22xp5_ASAP7_75t_L g423 ( 
.A1(n_386),
.A2(n_390),
.B1(n_398),
.B2(n_409),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_SL g387 ( 
.A(n_356),
.B(n_294),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_SL g434 ( 
.A(n_387),
.B(n_395),
.Y(n_434)
);

AOI22xp5_ASAP7_75t_L g388 ( 
.A1(n_336),
.A2(n_288),
.B1(n_330),
.B2(n_321),
.Y(n_388)
);

AOI22xp5_ASAP7_75t_L g389 ( 
.A1(n_353),
.A2(n_285),
.B1(n_293),
.B2(n_295),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_389),
.B(n_393),
.Y(n_415)
);

OAI22xp5_ASAP7_75t_SL g390 ( 
.A1(n_344),
.A2(n_329),
.B1(n_319),
.B2(n_322),
.Y(n_390)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_365),
.Y(n_392)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_392),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_349),
.B(n_298),
.Y(n_393)
);

XNOR2xp5_ASAP7_75t_SL g444 ( 
.A(n_396),
.B(n_389),
.Y(n_444)
);

NOR2xp33_ASAP7_75t_L g397 ( 
.A(n_354),
.B(n_333),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_SL g442 ( 
.A(n_397),
.B(n_399),
.Y(n_442)
);

OAI22xp5_ASAP7_75t_SL g398 ( 
.A1(n_344),
.A2(n_322),
.B1(n_286),
.B2(n_287),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_L g399 ( 
.A(n_354),
.B(n_287),
.Y(n_399)
);

AOI22xp5_ASAP7_75t_L g400 ( 
.A1(n_335),
.A2(n_300),
.B1(n_303),
.B2(n_308),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_400),
.B(n_401),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_340),
.B(n_317),
.Y(n_401)
);

AOI22xp5_ASAP7_75t_L g402 ( 
.A1(n_335),
.A2(n_286),
.B1(n_292),
.B2(n_337),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_402),
.B(n_403),
.Y(n_435)
);

AOI22xp5_ASAP7_75t_L g403 ( 
.A1(n_335),
.A2(n_361),
.B1(n_357),
.B2(n_368),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_359),
.Y(n_404)
);

CKINVDCx20_ASAP7_75t_R g405 ( 
.A(n_362),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_405),
.B(n_408),
.Y(n_445)
);

XOR2xp5_ASAP7_75t_L g407 ( 
.A(n_364),
.B(n_338),
.Y(n_407)
);

MAJIxp5_ASAP7_75t_L g422 ( 
.A(n_407),
.B(n_369),
.C(n_352),
.Y(n_422)
);

AOI22xp5_ASAP7_75t_L g408 ( 
.A1(n_357),
.A2(n_341),
.B1(n_375),
.B2(n_350),
.Y(n_408)
);

OAI22xp5_ASAP7_75t_SL g409 ( 
.A1(n_339),
.A2(n_358),
.B1(n_363),
.B2(n_340),
.Y(n_409)
);

CKINVDCx14_ASAP7_75t_R g411 ( 
.A(n_372),
.Y(n_411)
);

INVxp67_ASAP7_75t_L g418 ( 
.A(n_411),
.Y(n_418)
);

NOR2xp33_ASAP7_75t_SL g412 ( 
.A(n_339),
.B(n_370),
.Y(n_412)
);

CKINVDCx20_ASAP7_75t_R g420 ( 
.A(n_412),
.Y(n_420)
);

OAI21xp5_ASAP7_75t_L g414 ( 
.A1(n_391),
.A2(n_363),
.B(n_342),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_414),
.B(n_421),
.Y(n_467)
);

OAI22xp5_ASAP7_75t_SL g452 ( 
.A1(n_416),
.A2(n_426),
.B1(n_436),
.B2(n_408),
.Y(n_452)
);

AOI32xp33_ASAP7_75t_L g417 ( 
.A1(n_378),
.A2(n_374),
.A3(n_364),
.B1(n_343),
.B2(n_367),
.Y(n_417)
);

NOR2xp33_ASAP7_75t_L g471 ( 
.A(n_417),
.B(n_429),
.Y(n_471)
);

XNOR2xp5_ASAP7_75t_L g419 ( 
.A(n_407),
.B(n_366),
.Y(n_419)
);

XOR2xp5_ASAP7_75t_L g454 ( 
.A(n_419),
.B(n_430),
.Y(n_454)
);

OAI21xp5_ASAP7_75t_L g421 ( 
.A1(n_391),
.A2(n_369),
.B(n_359),
.Y(n_421)
);

MAJIxp5_ASAP7_75t_L g449 ( 
.A(n_422),
.B(n_428),
.C(n_440),
.Y(n_449)
);

CKINVDCx20_ASAP7_75t_R g424 ( 
.A(n_393),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_424),
.B(n_433),
.Y(n_470)
);

AOI22xp5_ASAP7_75t_L g426 ( 
.A1(n_390),
.A2(n_357),
.B1(n_352),
.B2(n_334),
.Y(n_426)
);

XNOR2x2_ASAP7_75t_SL g427 ( 
.A(n_379),
.B(n_334),
.Y(n_427)
);

XNOR2xp5_ASAP7_75t_L g446 ( 
.A(n_427),
.B(n_401),
.Y(n_446)
);

MAJIxp5_ASAP7_75t_L g428 ( 
.A(n_377),
.B(n_346),
.C(n_371),
.Y(n_428)
);

AOI21xp5_ASAP7_75t_L g429 ( 
.A1(n_378),
.A2(n_346),
.B(n_355),
.Y(n_429)
);

XOR2xp5_ASAP7_75t_L g430 ( 
.A(n_377),
.B(n_371),
.Y(n_430)
);

CKINVDCx20_ASAP7_75t_R g433 ( 
.A(n_394),
.Y(n_433)
);

AOI22xp5_ASAP7_75t_L g436 ( 
.A1(n_398),
.A2(n_410),
.B1(n_386),
.B2(n_409),
.Y(n_436)
);

OAI21xp5_ASAP7_75t_L g439 ( 
.A1(n_410),
.A2(n_397),
.B(n_394),
.Y(n_439)
);

CKINVDCx16_ASAP7_75t_R g463 ( 
.A(n_439),
.Y(n_463)
);

MAJIxp5_ASAP7_75t_L g440 ( 
.A(n_396),
.B(n_388),
.C(n_402),
.Y(n_440)
);

CKINVDCx20_ASAP7_75t_R g441 ( 
.A(n_395),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_441),
.B(n_399),
.Y(n_450)
);

XNOR2xp5_ASAP7_75t_SL g473 ( 
.A(n_444),
.B(n_415),
.Y(n_473)
);

INVx1_ASAP7_75t_SL g494 ( 
.A(n_446),
.Y(n_494)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_443),
.Y(n_447)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_447),
.Y(n_474)
);

AOI22xp5_ASAP7_75t_L g448 ( 
.A1(n_413),
.A2(n_405),
.B1(n_384),
.B2(n_380),
.Y(n_448)
);

OAI22xp5_ASAP7_75t_L g475 ( 
.A1(n_448),
.A2(n_464),
.B1(n_437),
.B2(n_431),
.Y(n_475)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_450),
.Y(n_477)
);

MAJIxp5_ASAP7_75t_L g451 ( 
.A(n_430),
.B(n_387),
.C(n_379),
.Y(n_451)
);

MAJIxp5_ASAP7_75t_L g476 ( 
.A(n_451),
.B(n_453),
.C(n_462),
.Y(n_476)
);

XOR2xp5_ASAP7_75t_L g482 ( 
.A(n_452),
.B(n_473),
.Y(n_482)
);

MAJIxp5_ASAP7_75t_L g453 ( 
.A(n_422),
.B(n_376),
.C(n_400),
.Y(n_453)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_443),
.Y(n_455)
);

NOR2xp33_ASAP7_75t_L g492 ( 
.A(n_455),
.B(n_457),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_SL g456 ( 
.A(n_420),
.B(n_412),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_SL g491 ( 
.A(n_456),
.B(n_459),
.Y(n_491)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_427),
.Y(n_457)
);

OAI22xp5_ASAP7_75t_SL g458 ( 
.A1(n_413),
.A2(n_376),
.B1(n_403),
.B2(n_385),
.Y(n_458)
);

AOI22xp5_ASAP7_75t_L g495 ( 
.A1(n_458),
.A2(n_461),
.B1(n_452),
.B2(n_463),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_SL g459 ( 
.A(n_420),
.B(n_404),
.Y(n_459)
);

XNOR2xp5_ASAP7_75t_L g460 ( 
.A(n_416),
.B(n_381),
.Y(n_460)
);

XNOR2xp5_ASAP7_75t_L g486 ( 
.A(n_460),
.B(n_466),
.Y(n_486)
);

OAI22xp5_ASAP7_75t_SL g461 ( 
.A1(n_426),
.A2(n_380),
.B1(n_382),
.B2(n_383),
.Y(n_461)
);

MAJIxp5_ASAP7_75t_L g462 ( 
.A(n_428),
.B(n_392),
.C(n_406),
.Y(n_462)
);

INVx1_ASAP7_75t_SL g464 ( 
.A(n_425),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_427),
.Y(n_465)
);

NOR2xp33_ASAP7_75t_SL g478 ( 
.A(n_465),
.B(n_442),
.Y(n_478)
);

XNOR2xp5_ASAP7_75t_L g466 ( 
.A(n_419),
.B(n_406),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_433),
.B(n_380),
.Y(n_468)
);

CKINVDCx20_ASAP7_75t_R g480 ( 
.A(n_468),
.Y(n_480)
);

MAJIxp5_ASAP7_75t_L g469 ( 
.A(n_440),
.B(n_444),
.C(n_423),
.Y(n_469)
);

MAJIxp5_ASAP7_75t_L g479 ( 
.A(n_469),
.B(n_435),
.C(n_429),
.Y(n_479)
);

XNOR2xp5_ASAP7_75t_L g472 ( 
.A(n_423),
.B(n_436),
.Y(n_472)
);

XNOR2xp5_ASAP7_75t_L g489 ( 
.A(n_472),
.B(n_432),
.Y(n_489)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_475),
.Y(n_508)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_478),
.Y(n_499)
);

XNOR2xp5_ASAP7_75t_L g497 ( 
.A(n_479),
.B(n_485),
.Y(n_497)
);

MAJIxp5_ASAP7_75t_L g481 ( 
.A(n_449),
.B(n_414),
.C(n_421),
.Y(n_481)
);

MAJIxp5_ASAP7_75t_L g503 ( 
.A(n_481),
.B(n_483),
.C(n_484),
.Y(n_503)
);

MAJIxp5_ASAP7_75t_L g483 ( 
.A(n_449),
.B(n_435),
.C(n_417),
.Y(n_483)
);

MAJIxp5_ASAP7_75t_L g484 ( 
.A(n_454),
.B(n_445),
.C(n_439),
.Y(n_484)
);

XOR2xp5_ASAP7_75t_L g485 ( 
.A(n_454),
.B(n_445),
.Y(n_485)
);

MAJIxp5_ASAP7_75t_L g487 ( 
.A(n_466),
.B(n_441),
.C(n_415),
.Y(n_487)
);

HB1xp67_ASAP7_75t_L g507 ( 
.A(n_487),
.Y(n_507)
);

XNOR2xp5_ASAP7_75t_L g488 ( 
.A(n_451),
.B(n_442),
.Y(n_488)
);

NOR2xp33_ASAP7_75t_L g504 ( 
.A(n_488),
.B(n_493),
.Y(n_504)
);

XNOR2xp5_ASAP7_75t_L g500 ( 
.A(n_489),
.B(n_490),
.Y(n_500)
);

XNOR2xp5_ASAP7_75t_L g490 ( 
.A(n_469),
.B(n_432),
.Y(n_490)
);

CKINVDCx20_ASAP7_75t_R g493 ( 
.A(n_470),
.Y(n_493)
);

OAI22xp5_ASAP7_75t_SL g502 ( 
.A1(n_495),
.A2(n_448),
.B1(n_471),
.B2(n_467),
.Y(n_502)
);

MAJIxp5_ASAP7_75t_L g496 ( 
.A(n_462),
.B(n_424),
.C(n_425),
.Y(n_496)
);

NOR2xp33_ASAP7_75t_L g505 ( 
.A(n_496),
.B(n_476),
.Y(n_505)
);

AND2x2_ASAP7_75t_L g498 ( 
.A(n_480),
.B(n_468),
.Y(n_498)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_498),
.Y(n_515)
);

XNOR2xp5_ASAP7_75t_L g501 ( 
.A(n_490),
.B(n_453),
.Y(n_501)
);

XNOR2xp5_ASAP7_75t_L g516 ( 
.A(n_501),
.B(n_476),
.Y(n_516)
);

AOI22xp5_ASAP7_75t_L g525 ( 
.A1(n_502),
.A2(n_511),
.B1(n_482),
.B2(n_473),
.Y(n_525)
);

NOR2xp33_ASAP7_75t_SL g519 ( 
.A(n_505),
.B(n_513),
.Y(n_519)
);

OAI21xp5_ASAP7_75t_SL g506 ( 
.A1(n_477),
.A2(n_450),
.B(n_460),
.Y(n_506)
);

AOI21xp5_ASAP7_75t_L g517 ( 
.A1(n_506),
.A2(n_514),
.B(n_484),
.Y(n_517)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_474),
.Y(n_509)
);

NOR2xp33_ASAP7_75t_L g521 ( 
.A(n_509),
.B(n_512),
.Y(n_521)
);

OAI22xp5_ASAP7_75t_L g510 ( 
.A1(n_491),
.A2(n_418),
.B1(n_434),
.B2(n_464),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_SL g520 ( 
.A(n_510),
.B(n_494),
.Y(n_520)
);

OAI22xp5_ASAP7_75t_SL g511 ( 
.A1(n_492),
.A2(n_458),
.B1(n_434),
.B2(n_446),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_496),
.Y(n_512)
);

CKINVDCx20_ASAP7_75t_R g513 ( 
.A(n_487),
.Y(n_513)
);

OAI21xp5_ASAP7_75t_SL g514 ( 
.A1(n_479),
.A2(n_461),
.B(n_472),
.Y(n_514)
);

NOR2xp33_ASAP7_75t_L g532 ( 
.A(n_516),
.B(n_525),
.Y(n_532)
);

INVxp67_ASAP7_75t_L g539 ( 
.A(n_517),
.Y(n_539)
);

OAI22xp5_ASAP7_75t_SL g518 ( 
.A1(n_508),
.A2(n_494),
.B1(n_483),
.B2(n_481),
.Y(n_518)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_518),
.Y(n_530)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_520),
.Y(n_534)
);

XOR2xp5_ASAP7_75t_L g522 ( 
.A(n_497),
.B(n_485),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_L g531 ( 
.A(n_522),
.B(n_523),
.Y(n_531)
);

XNOR2xp5_ASAP7_75t_L g523 ( 
.A(n_501),
.B(n_489),
.Y(n_523)
);

INVx6_ASAP7_75t_L g524 ( 
.A(n_504),
.Y(n_524)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_524),
.Y(n_536)
);

BUFx24_ASAP7_75t_SL g526 ( 
.A(n_499),
.Y(n_526)
);

NOR2xp33_ASAP7_75t_SL g533 ( 
.A(n_526),
.B(n_528),
.Y(n_533)
);

OAI21xp5_ASAP7_75t_SL g527 ( 
.A1(n_503),
.A2(n_431),
.B(n_437),
.Y(n_527)
);

HB1xp67_ASAP7_75t_L g535 ( 
.A(n_527),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_SL g528 ( 
.A(n_503),
.B(n_482),
.Y(n_528)
);

MAJIxp5_ASAP7_75t_L g529 ( 
.A(n_512),
.B(n_486),
.C(n_438),
.Y(n_529)
);

NOR2xp33_ASAP7_75t_L g537 ( 
.A(n_529),
.B(n_497),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_SL g543 ( 
.A(n_537),
.B(n_538),
.Y(n_543)
);

OAI22xp5_ASAP7_75t_L g538 ( 
.A1(n_515),
.A2(n_508),
.B1(n_507),
.B2(n_509),
.Y(n_538)
);

BUFx3_ASAP7_75t_L g540 ( 
.A(n_524),
.Y(n_540)
);

XOR2xp5_ASAP7_75t_L g542 ( 
.A(n_540),
.B(n_516),
.Y(n_542)
);

OAI21xp5_ASAP7_75t_SL g541 ( 
.A1(n_517),
.A2(n_498),
.B(n_502),
.Y(n_541)
);

AOI21xp5_ASAP7_75t_L g546 ( 
.A1(n_541),
.A2(n_539),
.B(n_535),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_L g549 ( 
.A(n_542),
.B(n_545),
.Y(n_549)
);

AOI31xp33_ASAP7_75t_L g544 ( 
.A1(n_539),
.A2(n_530),
.A3(n_532),
.B(n_534),
.Y(n_544)
);

MAJIxp5_ASAP7_75t_L g550 ( 
.A(n_544),
.B(n_547),
.C(n_543),
.Y(n_550)
);

XOR2xp5_ASAP7_75t_L g545 ( 
.A(n_531),
.B(n_523),
.Y(n_545)
);

AOI21xp5_ASAP7_75t_L g551 ( 
.A1(n_546),
.A2(n_548),
.B(n_541),
.Y(n_551)
);

XOR2xp5_ASAP7_75t_SL g547 ( 
.A(n_531),
.B(n_518),
.Y(n_547)
);

AOI21xp5_ASAP7_75t_L g548 ( 
.A1(n_536),
.A2(n_519),
.B(n_521),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_L g553 ( 
.A(n_550),
.B(n_551),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g552 ( 
.A(n_544),
.B(n_540),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_L g555 ( 
.A(n_552),
.B(n_529),
.Y(n_555)
);

O2A1O1Ixp33_ASAP7_75t_SL g554 ( 
.A1(n_549),
.A2(n_498),
.B(n_511),
.C(n_506),
.Y(n_554)
);

NOR2xp33_ASAP7_75t_SL g556 ( 
.A(n_554),
.B(n_525),
.Y(n_556)
);

AO21x2_ASAP7_75t_L g557 ( 
.A1(n_555),
.A2(n_533),
.B(n_514),
.Y(n_557)
);

AOI21x1_ASAP7_75t_L g558 ( 
.A1(n_556),
.A2(n_557),
.B(n_553),
.Y(n_558)
);

OAI21xp5_ASAP7_75t_SL g559 ( 
.A1(n_558),
.A2(n_438),
.B(n_522),
.Y(n_559)
);

OAI21xp5_ASAP7_75t_L g560 ( 
.A1(n_559),
.A2(n_500),
.B(n_486),
.Y(n_560)
);

XNOR2xp5_ASAP7_75t_L g561 ( 
.A(n_560),
.B(n_500),
.Y(n_561)
);


endmodule