module real_jpeg_4145_n_15 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_15);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_15;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_286;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_330;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_273;
wire n_253;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_299;
wire n_243;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

INVx8_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g169 ( 
.A(n_1),
.Y(n_169)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_1),
.Y(n_182)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_1),
.Y(n_207)
);

INVx3_ASAP7_75t_L g209 ( 
.A(n_1),
.Y(n_209)
);

BUFx6f_ASAP7_75t_L g214 ( 
.A(n_1),
.Y(n_214)
);

BUFx6f_ASAP7_75t_L g218 ( 
.A(n_1),
.Y(n_218)
);

INVx6_ASAP7_75t_L g221 ( 
.A(n_1),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g47 ( 
.A1(n_2),
.A2(n_38),
.B1(n_48),
.B2(n_50),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_2),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_2),
.A2(n_50),
.B1(n_131),
.B2(n_132),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_L g157 ( 
.A1(n_2),
.A2(n_50),
.B1(n_158),
.B2(n_160),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g217 ( 
.A1(n_2),
.A2(n_50),
.B1(n_218),
.B2(n_219),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_3),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_3),
.B(n_144),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_SL g247 ( 
.A1(n_3),
.A2(n_62),
.B1(n_121),
.B2(n_248),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_3),
.B(n_256),
.C(n_260),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_3),
.B(n_23),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_3),
.B(n_188),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_3),
.B(n_135),
.Y(n_300)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_4),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_4),
.Y(n_88)
);

BUFx3_ASAP7_75t_L g95 ( 
.A(n_4),
.Y(n_95)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

INVx8_ASAP7_75t_L g84 ( 
.A(n_6),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_6),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g188 ( 
.A(n_6),
.Y(n_188)
);

BUFx6f_ASAP7_75t_L g274 ( 
.A(n_6),
.Y(n_274)
);

BUFx5_ASAP7_75t_L g299 ( 
.A(n_6),
.Y(n_299)
);

AOI22xp33_ASAP7_75t_L g190 ( 
.A1(n_7),
.A2(n_158),
.B1(n_191),
.B2(n_192),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_7),
.Y(n_191)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_8),
.Y(n_65)
);

BUFx5_ASAP7_75t_L g67 ( 
.A(n_8),
.Y(n_67)
);

BUFx5_ASAP7_75t_L g174 ( 
.A(n_8),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g204 ( 
.A(n_8),
.Y(n_204)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_9),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_SL g36 ( 
.A1(n_10),
.A2(n_37),
.B1(n_43),
.B2(n_44),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_10),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_L g278 ( 
.A1(n_10),
.A2(n_44),
.B1(n_147),
.B2(n_279),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_L g293 ( 
.A1(n_10),
.A2(n_44),
.B1(n_294),
.B2(n_297),
.Y(n_293)
);

AOI22xp33_ASAP7_75t_L g69 ( 
.A1(n_11),
.A2(n_70),
.B1(n_76),
.B2(n_77),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_11),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g233 ( 
.A1(n_11),
.A2(n_76),
.B1(n_104),
.B2(n_234),
.Y(n_233)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_12),
.A2(n_121),
.B1(n_125),
.B2(n_128),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_12),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_L g225 ( 
.A1(n_12),
.A2(n_128),
.B1(n_226),
.B2(n_228),
.Y(n_225)
);

OAI22xp33_ASAP7_75t_SL g265 ( 
.A1(n_12),
.A2(n_128),
.B1(n_266),
.B2(n_269),
.Y(n_265)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_13),
.Y(n_107)
);

BUFx5_ASAP7_75t_L g109 ( 
.A(n_13),
.Y(n_109)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_13),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_13),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_14),
.A2(n_90),
.B1(n_91),
.B2(n_96),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_14),
.Y(n_96)
);

XOR2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_241),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_239),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_163),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_SL g240 ( 
.A(n_18),
.B(n_163),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_99),
.C(n_136),
.Y(n_18)
);

AOI22xp5_ASAP7_75t_L g328 ( 
.A1(n_19),
.A2(n_20),
.B1(n_329),
.B2(n_330),
.Y(n_328)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

XNOR2xp5_ASAP7_75t_SL g20 ( 
.A(n_21),
.B(n_60),
.Y(n_20)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_21),
.B(n_61),
.C(n_68),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_SL g21 ( 
.A1(n_22),
.A2(n_36),
.B(n_45),
.Y(n_21)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_22),
.A2(n_36),
.B1(n_52),
.B2(n_225),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_22),
.B(n_47),
.Y(n_323)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

OR2x2_ASAP7_75t_L g52 ( 
.A(n_23),
.B(n_53),
.Y(n_52)
);

AO22x2_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_28),
.B1(n_32),
.B2(n_34),
.Y(n_23)
);

INVx6_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_26),
.Y(n_35)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_27),
.Y(n_54)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_27),
.Y(n_57)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_27),
.Y(n_142)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_30),
.Y(n_127)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_31),
.Y(n_33)
);

INVx11_ASAP7_75t_L g105 ( 
.A(n_31),
.Y(n_105)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_31),
.Y(n_111)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_31),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_31),
.Y(n_139)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx5_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx4_ASAP7_75t_SL g38 ( 
.A(n_39),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_39),
.A2(n_49),
.B1(n_64),
.B2(n_66),
.Y(n_63)
);

INVx5_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_41),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g321 ( 
.A(n_41),
.Y(n_321)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_42),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_42),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g177 ( 
.A(n_42),
.Y(n_177)
);

INVx3_ASAP7_75t_L g227 ( 
.A(n_42),
.Y(n_227)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_42),
.Y(n_230)
);

OAI32xp33_ASAP7_75t_L g167 ( 
.A1(n_43),
.A2(n_168),
.A3(n_170),
.B1(n_172),
.B2(n_178),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_46),
.B(n_51),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx4_ASAP7_75t_L g138 ( 
.A(n_48),
.Y(n_138)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

AOI21xp5_ASAP7_75t_L g317 ( 
.A1(n_51),
.A2(n_318),
.B(n_323),
.Y(n_317)
);

INVx2_ASAP7_75t_SL g51 ( 
.A(n_52),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_L g53 ( 
.A1(n_54),
.A2(n_55),
.B1(n_57),
.B2(n_58),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx6_ASAP7_75t_L g150 ( 
.A(n_57),
.Y(n_150)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

XOR2xp5_ASAP7_75t_L g60 ( 
.A(n_61),
.B(n_68),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_62),
.B(n_63),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_62),
.B(n_179),
.Y(n_178)
);

OAI21xp33_ASAP7_75t_SL g211 ( 
.A1(n_62),
.A2(n_178),
.B(n_212),
.Y(n_211)
);

AOI21xp5_ASAP7_75t_L g290 ( 
.A1(n_62),
.A2(n_185),
.B(n_272),
.Y(n_290)
);

OAI21xp33_ASAP7_75t_SL g318 ( 
.A1(n_62),
.A2(n_319),
.B(n_322),
.Y(n_318)
);

AND2x2_ASAP7_75t_L g200 ( 
.A(n_63),
.B(n_201),
.Y(n_200)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_63),
.Y(n_222)
);

INVx6_ASAP7_75t_L g171 ( 
.A(n_64),
.Y(n_171)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_69),
.A2(n_81),
.B1(n_89),
.B2(n_97),
.Y(n_68)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_69),
.Y(n_152)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx4_ASAP7_75t_SL g71 ( 
.A(n_72),
.Y(n_71)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx5_ASAP7_75t_L g80 ( 
.A(n_74),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_74),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g162 ( 
.A(n_75),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g271 ( 
.A(n_75),
.Y(n_271)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

HB1xp67_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g262 ( 
.A(n_80),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_81),
.B(n_157),
.Y(n_156)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_81),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_81),
.A2(n_273),
.B1(n_304),
.B2(n_305),
.Y(n_303)
);

OR2x2_ASAP7_75t_L g81 ( 
.A(n_82),
.B(n_85),
.Y(n_81)
);

INVx8_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_84),
.Y(n_98)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx6_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_88),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_88),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g296 ( 
.A(n_88),
.Y(n_296)
);

INVxp67_ASAP7_75t_L g186 ( 
.A(n_89),
.Y(n_186)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

BUFx8_ASAP7_75t_L g159 ( 
.A(n_95),
.Y(n_159)
);

BUFx5_ASAP7_75t_L g193 ( 
.A(n_95),
.Y(n_193)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

XNOR2xp5_ASAP7_75t_SL g330 ( 
.A(n_99),
.B(n_136),
.Y(n_330)
);

OAI21xp5_ASAP7_75t_SL g99 ( 
.A1(n_100),
.A2(n_120),
.B(n_129),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_SL g246 ( 
.A1(n_100),
.A2(n_129),
.B(n_247),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_100),
.A2(n_120),
.B1(n_232),
.B2(n_278),
.Y(n_315)
);

INVx2_ASAP7_75t_SL g100 ( 
.A(n_101),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_101),
.B(n_130),
.Y(n_237)
);

AND2x2_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_112),
.Y(n_101)
);

OAI22xp33_ASAP7_75t_L g102 ( 
.A1(n_103),
.A2(n_106),
.B1(n_108),
.B2(n_110),
.Y(n_102)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx6_ASAP7_75t_L g134 ( 
.A(n_105),
.Y(n_134)
);

INVx6_ASAP7_75t_L g148 ( 
.A(n_105),
.Y(n_148)
);

INVx5_ASAP7_75t_L g236 ( 
.A(n_105),
.Y(n_236)
);

BUFx6f_ASAP7_75t_L g280 ( 
.A(n_105),
.Y(n_280)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx5_ASAP7_75t_L g259 ( 
.A(n_107),
.Y(n_259)
);

INVx4_ASAP7_75t_SL g108 ( 
.A(n_109),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_112),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_SL g277 ( 
.A1(n_112),
.A2(n_237),
.B(n_278),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_113),
.A2(n_116),
.B1(n_117),
.B2(n_118),
.Y(n_112)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx4_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_121),
.Y(n_131)
);

INVx5_ASAP7_75t_SL g121 ( 
.A(n_122),
.Y(n_121)
);

INVx4_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx4_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_130),
.B(n_135),
.Y(n_129)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx6_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_134),
.Y(n_254)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_135),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_151),
.Y(n_136)
);

XOR2xp5_ASAP7_75t_L g324 ( 
.A(n_137),
.B(n_151),
.Y(n_324)
);

AOI32xp33_ASAP7_75t_L g137 ( 
.A1(n_138),
.A2(n_139),
.A3(n_140),
.B1(n_143),
.B2(n_146),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVx4_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

INVxp33_ASAP7_75t_L g322 ( 
.A(n_143),
.Y(n_322)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

NAND2xp33_ASAP7_75t_SL g146 ( 
.A(n_147),
.B(n_149),
.Y(n_146)
);

INVx8_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVx4_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_L g151 ( 
.A1(n_152),
.A2(n_153),
.B(n_156),
.Y(n_151)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

INVx3_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_L g292 ( 
.A1(n_156),
.A2(n_293),
.B(n_299),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_157),
.B(n_273),
.Y(n_272)
);

INVx8_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

INVx4_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

INVx4_ASAP7_75t_L g268 ( 
.A(n_161),
.Y(n_268)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_197),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_165),
.A2(n_194),
.B1(n_195),
.B2(n_196),
.Y(n_164)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_165),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_166),
.A2(n_167),
.B1(n_183),
.B2(n_184),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

INVx8_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_173),
.B(n_175),
.Y(n_172)
);

INVx6_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

INVx4_ASAP7_75t_L g210 ( 
.A(n_174),
.Y(n_210)
);

INVx1_ASAP7_75t_SL g175 ( 
.A(n_176),
.Y(n_175)
);

INVx6_ASAP7_75t_SL g176 ( 
.A(n_177),
.Y(n_176)
);

INVx3_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

INVx4_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_185),
.A2(n_186),
.B1(n_187),
.B2(n_189),
.Y(n_184)
);

AOI21xp5_ASAP7_75t_L g264 ( 
.A1(n_185),
.A2(n_265),
.B(n_272),
.Y(n_264)
);

BUFx6f_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

INVxp67_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

BUFx2_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

INVx3_ASAP7_75t_L g288 ( 
.A(n_193),
.Y(n_288)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_194),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_198),
.A2(n_199),
.B1(n_223),
.B2(n_238),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

AOI21xp5_ASAP7_75t_L g199 ( 
.A1(n_200),
.A2(n_211),
.B(n_215),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_202),
.A2(n_205),
.B1(n_208),
.B2(n_210),
.Y(n_201)
);

INVx6_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

INVx4_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

INVx5_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

INVx3_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

INVx6_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_222),
.Y(n_216)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_223),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_SL g223 ( 
.A(n_224),
.B(n_231),
.Y(n_223)
);

INVx4_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

INVx6_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

OAI21xp5_ASAP7_75t_SL g231 ( 
.A1(n_232),
.A2(n_233),
.B(n_237),
.Y(n_231)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

INVx5_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

BUFx2_ASAP7_75t_L g249 ( 
.A(n_236),
.Y(n_249)
);

INVxp67_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

AO21x1_ASAP7_75t_SL g241 ( 
.A1(n_242),
.A2(n_326),
.B(n_331),
.Y(n_241)
);

OAI21x1_ASAP7_75t_L g242 ( 
.A1(n_243),
.A2(n_310),
.B(n_325),
.Y(n_242)
);

AOI21xp5_ASAP7_75t_L g243 ( 
.A1(n_244),
.A2(n_283),
.B(n_309),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_263),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_245),
.B(n_263),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_246),
.B(n_250),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_246),
.A2(n_250),
.B1(n_251),
.B2(n_307),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_246),
.Y(n_307)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_255),
.Y(n_251)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

BUFx6f_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

INVx3_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_264),
.B(n_275),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_264),
.B(n_276),
.C(n_282),
.Y(n_311)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_265),
.Y(n_305)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

INVx6_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

INVx4_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

INVx4_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

INVx8_ASAP7_75t_L g298 ( 
.A(n_271),
.Y(n_298)
);

INVx4_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_276),
.A2(n_277),
.B1(n_281),
.B2(n_282),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

INVx11_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

OAI21xp5_ASAP7_75t_L g283 ( 
.A1(n_284),
.A2(n_302),
.B(n_308),
.Y(n_283)
);

AOI21xp5_ASAP7_75t_L g284 ( 
.A1(n_285),
.A2(n_291),
.B(n_301),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_286),
.B(n_290),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_287),
.B(n_289),
.Y(n_286)
);

INVx1_ASAP7_75t_SL g287 ( 
.A(n_288),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g291 ( 
.A(n_292),
.B(n_300),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_292),
.B(n_300),
.Y(n_301)
);

INVxp67_ASAP7_75t_L g304 ( 
.A(n_293),
.Y(n_304)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

INVx3_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

INVx4_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_303),
.B(n_306),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_303),
.B(n_306),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_311),
.B(n_312),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_311),
.B(n_312),
.Y(n_325)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_313),
.B(n_324),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_314),
.A2(n_315),
.B1(n_316),
.B2(n_317),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_315),
.B(n_316),
.C(n_324),
.Y(n_327)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

INVx6_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

INVx6_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_327),
.B(n_328),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_SL g331 ( 
.A(n_327),
.B(n_328),
.Y(n_331)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);


endmodule