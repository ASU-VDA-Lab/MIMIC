module fake_jpeg_1248_n_203 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_203);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_203;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_202;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx8_ASAP7_75t_L g49 ( 
.A(n_24),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_40),
.Y(n_50)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_15),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_47),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_19),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_6),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_3),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_4),
.Y(n_56)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_33),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_16),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_41),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_1),
.Y(n_60)
);

BUFx5_ASAP7_75t_L g61 ( 
.A(n_18),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_16),
.Y(n_62)
);

INVx2_ASAP7_75t_SL g63 ( 
.A(n_48),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_30),
.Y(n_64)
);

BUFx6f_ASAP7_75t_SL g65 ( 
.A(n_2),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_31),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_20),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_36),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_29),
.Y(n_69)
);

INVxp33_ASAP7_75t_L g70 ( 
.A(n_45),
.Y(n_70)
);

BUFx5_ASAP7_75t_L g71 ( 
.A(n_8),
.Y(n_71)
);

BUFx12f_ASAP7_75t_L g72 ( 
.A(n_49),
.Y(n_72)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_72),
.Y(n_93)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_65),
.Y(n_73)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_73),
.Y(n_81)
);

BUFx12f_ASAP7_75t_L g74 ( 
.A(n_49),
.Y(n_74)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_74),
.Y(n_92)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_62),
.Y(n_75)
);

BUFx2_ASAP7_75t_L g86 ( 
.A(n_75),
.Y(n_86)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_51),
.Y(n_76)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_76),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_68),
.Y(n_77)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_77),
.Y(n_90)
);

INVx8_ASAP7_75t_L g78 ( 
.A(n_68),
.Y(n_78)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_78),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_58),
.Y(n_79)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_79),
.Y(n_89)
);

INVx8_ASAP7_75t_L g80 ( 
.A(n_58),
.Y(n_80)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_80),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_76),
.B(n_54),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_84),
.B(n_85),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_72),
.B(n_54),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_79),
.A2(n_51),
.B1(n_62),
.B2(n_57),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_87),
.A2(n_94),
.B1(n_63),
.B2(n_57),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_80),
.A2(n_65),
.B1(n_52),
.B2(n_50),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_88),
.A2(n_78),
.B1(n_70),
.B2(n_60),
.Y(n_105)
);

OR2x2_ASAP7_75t_L g91 ( 
.A(n_73),
.B(n_56),
.Y(n_91)
);

NAND2x1_ASAP7_75t_SL g99 ( 
.A(n_91),
.B(n_67),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_75),
.A2(n_63),
.B1(n_56),
.B2(n_67),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_96),
.A2(n_0),
.B1(n_1),
.B2(n_4),
.Y(n_123)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_81),
.Y(n_97)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_97),
.Y(n_116)
);

OAI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_88),
.A2(n_77),
.B1(n_64),
.B2(n_59),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_98),
.A2(n_105),
.B1(n_112),
.B2(n_93),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_99),
.B(n_101),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_91),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_L g102 ( 
.A1(n_89),
.A2(n_77),
.B1(n_63),
.B2(n_53),
.Y(n_102)
);

OAI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_102),
.A2(n_71),
.B1(n_61),
.B2(n_3),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_86),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g120 ( 
.A(n_103),
.B(n_106),
.Y(n_120)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_90),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_104),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_83),
.B(n_50),
.Y(n_106)
);

XOR2xp5_ASAP7_75t_L g107 ( 
.A(n_83),
.B(n_52),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_107),
.B(n_93),
.C(n_74),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_90),
.B(n_69),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_108),
.B(n_111),
.Y(n_115)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_81),
.Y(n_109)
);

BUFx3_ASAP7_75t_L g118 ( 
.A(n_109),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_86),
.B(n_55),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_110),
.B(n_0),
.Y(n_126)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_95),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_82),
.A2(n_72),
.B1(n_74),
.B2(n_70),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_92),
.A2(n_66),
.B1(n_72),
.B2(n_74),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_113),
.A2(n_71),
.B1(n_61),
.B2(n_2),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_92),
.B(n_35),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_114),
.B(n_6),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_117),
.B(n_134),
.C(n_26),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_119),
.B(n_122),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_121),
.A2(n_7),
.B1(n_10),
.B2(n_11),
.Y(n_143)
);

INVxp67_ASAP7_75t_L g136 ( 
.A(n_123),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_126),
.B(n_130),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_108),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_127),
.B(n_128),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_100),
.B(n_5),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_99),
.B(n_5),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_129),
.B(n_131),
.Y(n_144)
);

AND2x6_ASAP7_75t_L g130 ( 
.A(n_107),
.B(n_22),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_111),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_132),
.B(n_133),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_114),
.B(n_109),
.Y(n_133)
);

XOR2xp5_ASAP7_75t_L g134 ( 
.A(n_97),
.B(n_105),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_104),
.B(n_23),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_135),
.B(n_46),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_119),
.A2(n_113),
.B1(n_112),
.B2(n_9),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_137),
.A2(n_138),
.B1(n_143),
.B2(n_135),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_134),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_138)
);

INVxp67_ASAP7_75t_L g139 ( 
.A(n_120),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_139),
.B(n_157),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_124),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_142),
.B(n_149),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_145),
.B(n_148),
.C(n_151),
.Y(n_176)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_116),
.Y(n_146)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_146),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_117),
.B(n_25),
.C(n_44),
.Y(n_148)
);

AOI21xp5_ASAP7_75t_SL g150 ( 
.A1(n_125),
.A2(n_10),
.B(n_11),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_SL g171 ( 
.A1(n_150),
.A2(n_152),
.B(n_14),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_115),
.B(n_27),
.C(n_42),
.Y(n_151)
);

AOI21xp5_ASAP7_75t_L g152 ( 
.A1(n_116),
.A2(n_12),
.B(n_13),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_124),
.Y(n_153)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_153),
.Y(n_170)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_118),
.Y(n_155)
);

INVx2_ASAP7_75t_SL g175 ( 
.A(n_155),
.Y(n_175)
);

AO22x1_ASAP7_75t_SL g156 ( 
.A1(n_121),
.A2(n_43),
.B1(n_39),
.B2(n_38),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_156),
.B(n_12),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_115),
.B(n_37),
.C(n_34),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_118),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_158),
.B(n_14),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_SL g160 ( 
.A(n_147),
.B(n_132),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_160),
.B(n_162),
.Y(n_183)
);

AOI21xp5_ASAP7_75t_L g163 ( 
.A1(n_140),
.A2(n_130),
.B(n_32),
.Y(n_163)
);

AOI21xp5_ASAP7_75t_L g180 ( 
.A1(n_163),
.A2(n_148),
.B(n_157),
.Y(n_180)
);

CKINVDCx14_ASAP7_75t_R g178 ( 
.A(n_165),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_145),
.B(n_28),
.Y(n_166)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_166),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_138),
.B(n_13),
.Y(n_167)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_167),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_139),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_SL g177 ( 
.A(n_168),
.B(n_169),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_SL g179 ( 
.A1(n_171),
.A2(n_150),
.B(n_167),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_137),
.A2(n_15),
.B1(n_17),
.B2(n_18),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_172),
.A2(n_174),
.B1(n_154),
.B2(n_136),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_144),
.B(n_17),
.Y(n_173)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_173),
.B(n_151),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_143),
.A2(n_19),
.B1(n_20),
.B2(n_21),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_179),
.B(n_171),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_L g191 ( 
.A1(n_180),
.A2(n_159),
.B(n_136),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_181),
.B(n_176),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_184),
.A2(n_162),
.B1(n_172),
.B2(n_163),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_185),
.B(n_176),
.C(n_181),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_186),
.B(n_180),
.C(n_179),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_187),
.B(n_188),
.Y(n_193)
);

OAI322xp33_ASAP7_75t_L g188 ( 
.A1(n_183),
.A2(n_161),
.A3(n_141),
.B1(n_165),
.B2(n_170),
.C1(n_166),
.C2(n_164),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_189),
.B(n_191),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_190),
.A2(n_184),
.B1(n_178),
.B2(n_182),
.Y(n_192)
);

MAJx2_ASAP7_75t_L g196 ( 
.A(n_192),
.B(n_194),
.C(n_188),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_196),
.B(n_197),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_SL g197 ( 
.A(n_193),
.B(n_177),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_L g198 ( 
.A1(n_197),
.A2(n_195),
.B(n_194),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_198),
.B(n_156),
.Y(n_200)
);

O2A1O1Ixp33_ASAP7_75t_L g201 ( 
.A1(n_200),
.A2(n_156),
.B(n_174),
.C(n_199),
.Y(n_201)
);

OAI21x1_ASAP7_75t_L g202 ( 
.A1(n_201),
.A2(n_175),
.B(n_21),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_202),
.B(n_175),
.Y(n_203)
);


endmodule