module fake_jpeg_17928_n_46 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_46);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_46;

wire n_13;
wire n_21;
wire n_33;
wire n_45;
wire n_23;
wire n_10;
wire n_27;
wire n_22;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

INVx8_ASAP7_75t_L g7 ( 
.A(n_2),
.Y(n_7)
);

INVx2_ASAP7_75t_L g8 ( 
.A(n_4),
.Y(n_8)
);

INVx4_ASAP7_75t_L g9 ( 
.A(n_2),
.Y(n_9)
);

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_6),
.Y(n_10)
);

BUFx3_ASAP7_75t_L g11 ( 
.A(n_2),
.Y(n_11)
);

BUFx5_ASAP7_75t_L g12 ( 
.A(n_1),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_6),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_L g14 ( 
.A(n_3),
.B(n_0),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_0),
.B(n_4),
.Y(n_15)
);

AOI22xp5_ASAP7_75t_L g16 ( 
.A1(n_8),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_16)
);

OAI22xp5_ASAP7_75t_SL g27 ( 
.A1(n_16),
.A2(n_23),
.B1(n_7),
.B2(n_13),
.Y(n_27)
);

OR2x2_ASAP7_75t_L g17 ( 
.A(n_10),
.B(n_1),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_17),
.B(n_22),
.Y(n_33)
);

OAI22xp33_ASAP7_75t_SL g18 ( 
.A1(n_9),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_18)
);

AOI22xp5_ASAP7_75t_L g29 ( 
.A1(n_18),
.A2(n_11),
.B1(n_16),
.B2(n_22),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_14),
.B(n_15),
.Y(n_19)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_19),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_20),
.Y(n_28)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_11),
.B(n_5),
.C(n_12),
.Y(n_21)
);

XNOR2xp5_ASAP7_75t_L g30 ( 
.A(n_21),
.B(n_17),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_13),
.Y(n_22)
);

AOI22xp33_ASAP7_75t_SL g23 ( 
.A1(n_8),
.A2(n_5),
.B1(n_9),
.B2(n_7),
.Y(n_23)
);

AOI21xp5_ASAP7_75t_L g24 ( 
.A1(n_14),
.A2(n_15),
.B(n_9),
.Y(n_24)
);

OAI21xp5_ASAP7_75t_L g31 ( 
.A1(n_24),
.A2(n_21),
.B(n_20),
.Y(n_31)
);

AOI32xp33_ASAP7_75t_L g25 ( 
.A1(n_24),
.A2(n_10),
.A3(n_11),
.B1(n_12),
.B2(n_7),
.Y(n_25)
);

XOR2x2_ASAP7_75t_SL g38 ( 
.A(n_25),
.B(n_27),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g36 ( 
.A1(n_27),
.A2(n_29),
.B1(n_33),
.B2(n_26),
.Y(n_36)
);

XOR2xp5_ASAP7_75t_L g34 ( 
.A(n_30),
.B(n_31),
.Y(n_34)
);

XNOR2xp5_ASAP7_75t_L g32 ( 
.A(n_20),
.B(n_24),
.Y(n_32)
);

MAJIxp5_ASAP7_75t_L g39 ( 
.A(n_32),
.B(n_30),
.C(n_29),
.Y(n_39)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_28),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_35),
.B(n_37),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_SL g40 ( 
.A1(n_36),
.A2(n_38),
.B1(n_32),
.B2(n_37),
.Y(n_40)
);

INVxp67_ASAP7_75t_L g37 ( 
.A(n_31),
.Y(n_37)
);

XOR2xp5_ASAP7_75t_L g42 ( 
.A(n_39),
.B(n_34),
.Y(n_42)
);

XNOR2xp5_ASAP7_75t_L g44 ( 
.A(n_40),
.B(n_42),
.Y(n_44)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_41),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_43),
.B(n_40),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_45),
.A2(n_38),
.B1(n_44),
.B2(n_42),
.Y(n_46)
);


endmodule