module real_jpeg_33516_n_8 (n_5, n_4, n_0, n_1, n_2, n_6, n_7, n_3, n_8);

input n_5;
input n_4;
input n_0;
input n_1;
input n_2;
input n_6;
input n_7;
input n_3;

output n_8;

wire n_17;
wire n_43;
wire n_37;
wire n_21;
wire n_38;
wire n_33;
wire n_50;
wire n_35;
wire n_29;
wire n_49;
wire n_10;
wire n_31;
wire n_9;
wire n_52;
wire n_12;
wire n_24;
wire n_34;
wire n_28;
wire n_44;
wire n_46;
wire n_23;
wire n_11;
wire n_14;
wire n_47;
wire n_51;
wire n_45;
wire n_25;
wire n_42;
wire n_22;
wire n_18;
wire n_53;
wire n_39;
wire n_36;
wire n_40;
wire n_41;
wire n_26;
wire n_32;
wire n_27;
wire n_19;
wire n_20;
wire n_48;
wire n_30;
wire n_16;
wire n_15;
wire n_13;

OAI21xp33_ASAP7_75t_L g8 ( 
.A1(n_0),
.A2(n_9),
.B(n_10),
.Y(n_8)
);

NAND2xp5_ASAP7_75t_SL g10 ( 
.A(n_0),
.B(n_11),
.Y(n_10)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

OR2x2_ASAP7_75t_L g31 ( 
.A(n_1),
.B(n_32),
.Y(n_31)
);

OR2x2_ASAP7_75t_L g47 ( 
.A(n_1),
.B(n_45),
.Y(n_47)
);

BUFx2_ASAP7_75t_R g20 ( 
.A(n_2),
.Y(n_20)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_2),
.Y(n_38)
);

NAND2x1p5_ASAP7_75t_L g39 ( 
.A(n_2),
.B(n_18),
.Y(n_39)
);

INVx1_ASAP7_75t_L g9 ( 
.A(n_3),
.Y(n_9)
);

AND2x4_ASAP7_75t_SL g12 ( 
.A(n_4),
.B(n_13),
.Y(n_12)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_4),
.B(n_41),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_4),
.B(n_32),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_4),
.B(n_42),
.Y(n_53)
);

OR2x2_ASAP7_75t_L g25 ( 
.A(n_5),
.B(n_26),
.Y(n_25)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

OA22x2_ASAP7_75t_L g16 ( 
.A1(n_6),
.A2(n_7),
.B1(n_17),
.B2(n_18),
.Y(n_16)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

AO21x1_ASAP7_75t_L g42 ( 
.A1(n_6),
.A2(n_37),
.B(n_39),
.Y(n_42)
);

INVx3_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

AND2x2_ASAP7_75t_L g37 ( 
.A(n_7),
.B(n_38),
.Y(n_37)
);

O2A1O1Ixp33_ASAP7_75t_L g11 ( 
.A1(n_12),
.A2(n_21),
.B(n_24),
.C(n_27),
.Y(n_11)
);

INVx2_ASAP7_75t_L g13 ( 
.A(n_14),
.Y(n_13)
);

AND2x2_ASAP7_75t_L g30 ( 
.A(n_14),
.B(n_23),
.Y(n_30)
);

OA22x2_ASAP7_75t_L g14 ( 
.A1(n_15),
.A2(n_16),
.B1(n_19),
.B2(n_20),
.Y(n_14)
);

INVx2_ASAP7_75t_L g15 ( 
.A(n_16),
.Y(n_15)
);

OA21x2_ASAP7_75t_L g36 ( 
.A1(n_17),
.A2(n_37),
.B(n_39),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_SL g22 ( 
.A(n_19),
.B(n_23),
.Y(n_22)
);

OR2x2_ASAP7_75t_L g28 ( 
.A(n_19),
.B(n_23),
.Y(n_28)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

OR2x2_ASAP7_75t_L g35 ( 
.A(n_23),
.B(n_36),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_25),
.Y(n_24)
);

INVx2_ASAP7_75t_R g44 ( 
.A(n_26),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_26),
.B(n_50),
.Y(n_49)
);

A2O1A1Ixp33_ASAP7_75t_L g27 ( 
.A1(n_28),
.A2(n_29),
.B(n_31),
.C(n_33),
.Y(n_27)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_32),
.Y(n_45)
);

O2A1O1Ixp33_ASAP7_75t_L g33 ( 
.A1(n_34),
.A2(n_40),
.B(n_43),
.C(n_46),
.Y(n_33)
);

CKINVDCx16_ASAP7_75t_R g34 ( 
.A(n_35),
.Y(n_34)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

AND2x2_ASAP7_75t_L g43 ( 
.A(n_44),
.B(n_45),
.Y(n_43)
);

O2A1O1Ixp33_ASAP7_75t_L g46 ( 
.A1(n_47),
.A2(n_48),
.B(n_49),
.C(n_52),
.Y(n_46)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);


endmodule