module real_aes_16597_n_249 (n_17, n_28, n_226, n_76, n_202, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_238, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_230, n_165, n_51, n_195, n_246, n_248, n_176, n_27, n_163, n_222, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_18, n_207, n_104, n_21, n_31, n_8, n_183, n_205, n_220, n_211, n_10, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_234, n_153, n_75, n_178, n_219, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_239, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_95, n_131, n_144, n_164, n_231, n_169, n_242, n_44, n_102, n_188, n_152, n_198, n_201, n_122, n_7, n_228, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_69, n_46, n_109, n_59, n_25, n_203, n_236, n_73, n_77, n_218, n_81, n_133, n_48, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_138, n_50, n_114, n_89, n_170, n_26, n_235, n_86, n_93, n_182, n_154, n_127, n_199, n_245, n_161, n_189, n_13, n_24, n_217, n_2, n_142, n_55, n_168, n_175, n_241, n_145, n_62, n_105, n_223, n_84, n_227, n_67, n_92, n_33, n_206, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_116, n_94, n_229, n_39, n_5, n_45, n_60, n_233, n_240, n_247, n_38, n_155, n_243, n_118, n_143, n_139, n_244, n_192, n_213, n_136, n_87, n_171, n_0, n_157, n_78, n_101, n_63, n_1, n_146, n_237, n_107, n_184, n_53, n_36, n_249);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_238;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_230;
input n_165;
input n_51;
input n_195;
input n_246;
input n_248;
input n_176;
input n_27;
input n_163;
input n_222;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_183;
input n_205;
input n_220;
input n_211;
input n_10;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_234;
input n_153;
input n_75;
input n_178;
input n_219;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_239;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_242;
input n_44;
input n_102;
input n_188;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_69;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_236;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_138;
input n_50;
input n_114;
input n_89;
input n_170;
input n_26;
input n_235;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_245;
input n_161;
input n_189;
input n_13;
input n_24;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_241;
input n_145;
input n_62;
input n_105;
input n_223;
input n_84;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_116;
input n_94;
input n_229;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_240;
input n_247;
input n_38;
input n_155;
input n_243;
input n_118;
input n_143;
input n_139;
input n_244;
input n_192;
input n_213;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_101;
input n_63;
input n_1;
input n_146;
input n_237;
input n_107;
input n_184;
input n_53;
input n_36;
output n_249;
wire n_476;
wire n_887;
wire n_599;
wire n_1279;
wire n_1314;
wire n_830;
wire n_1371;
wire n_624;
wire n_618;
wire n_933;
wire n_485;
wire n_822;
wire n_750;
wire n_503;
wire n_254;
wire n_469;
wire n_1310;
wire n_1376;
wire n_592;
wire n_761;
wire n_421;
wire n_329;
wire n_919;
wire n_1217;
wire n_1423;
wire n_571;
wire n_549;
wire n_1034;
wire n_1328;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_593;
wire n_989;
wire n_431;
wire n_1044;
wire n_963;
wire n_551;
wire n_884;
wire n_260;
wire n_814;
wire n_944;
wire n_1283;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_1313;
wire n_1468;
wire n_870;
wire n_1248;
wire n_271;
wire n_548;
wire n_572;
wire n_815;
wire n_1140;
wire n_1453;
wire n_330;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_292;
wire n_1379;
wire n_400;
wire n_1415;
wire n_1160;
wire n_1287;
wire n_883;
wire n_478;
wire n_553;
wire n_1367;
wire n_744;
wire n_1325;
wire n_1441;
wire n_1382;
wire n_875;
wire n_951;
wire n_1199;
wire n_1225;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_1477;
wire n_595;
wire n_343;
wire n_1282;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_281;
wire n_962;
wire n_755;
wire n_409;
wire n_781;
wire n_576;
wire n_956;
wire n_1242;
wire n_796;
wire n_874;
wire n_1126;
wire n_383;
wire n_455;
wire n_682;
wire n_812;
wire n_817;
wire n_782;
wire n_760;
wire n_608;
wire n_534;
wire n_1454;
wire n_708;
wire n_1020;
wire n_885;
wire n_950;
wire n_381;
wire n_1196;
wire n_1013;
wire n_808;
wire n_1224;
wire n_688;
wire n_1042;
wire n_363;
wire n_1317;
wire n_417;
wire n_323;
wire n_690;
wire n_1419;
wire n_499;
wire n_1142;
wire n_947;
wire n_970;
wire n_1149;
wire n_368;
wire n_527;
wire n_1342;
wire n_1440;
wire n_1346;
wire n_552;
wire n_1383;
wire n_590;
wire n_1293;
wire n_432;
wire n_1131;
wire n_1008;
wire n_805;
wire n_619;
wire n_1095;
wire n_1250;
wire n_1284;
wire n_360;
wire n_1465;
wire n_859;
wire n_1304;
wire n_685;
wire n_1080;
wire n_917;
wire n_1247;
wire n_488;
wire n_501;
wire n_1380;
wire n_954;
wire n_702;
wire n_1007;
wire n_351;
wire n_898;
wire n_562;
wire n_1022;
wire n_404;
wire n_1073;
wire n_728;
wire n_1301;
wire n_1201;
wire n_997;
wire n_1105;
wire n_1243;
wire n_306;
wire n_1003;
wire n_346;
wire n_293;
wire n_749;
wire n_914;
wire n_1286;
wire n_494;
wire n_927;
wire n_723;
wire n_1351;
wire n_972;
wire n_1209;
wire n_411;
wire n_498;
wire n_1397;
wire n_765;
wire n_648;
wire n_939;
wire n_290;
wire n_928;
wire n_1384;
wire n_789;
wire n_738;
wire n_1387;
wire n_922;
wire n_1048;
wire n_1422;
wire n_787;
wire n_1214;
wire n_806;
wire n_715;
wire n_420;
wire n_1258;
wire n_873;
wire n_438;
wire n_446;
wire n_1281;
wire n_712;
wire n_266;
wire n_422;
wire n_861;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_724;
wire n_440;
wire n_1231;
wire n_1305;
wire n_315;
wire n_1161;
wire n_686;
wire n_1299;
wire n_949;
wire n_586;
wire n_1421;
wire n_788;
wire n_441;
wire n_1045;
wire n_1339;
wire n_837;
wire n_1349;
wire n_1445;
wire n_829;
wire n_1030;
wire n_1348;
wire n_1391;
wire n_375;
wire n_597;
wire n_1036;
wire n_687;
wire n_258;
wire n_652;
wire n_500;
wire n_804;
wire n_1173;
wire n_854;
wire n_424;
wire n_877;
wire n_802;
wire n_337;
wire n_264;
wire n_480;
wire n_684;
wire n_1178;
wire n_821;
wire n_1018;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_635;
wire n_792;
wire n_1392;
wire n_665;
wire n_667;
wire n_991;
wire n_1004;
wire n_580;
wire n_1417;
wire n_1370;
wire n_979;
wire n_445;
wire n_596;
wire n_1197;
wire n_657;
wire n_328;
wire n_1260;
wire n_355;
wire n_1129;
wire n_1285;
wire n_742;
wire n_1014;
wire n_1385;
wire n_461;
wire n_1047;
wire n_1016;
wire n_694;
wire n_1350;
wire n_894;
wire n_545;
wire n_1459;
wire n_401;
wire n_538;
wire n_537;
wire n_560;
wire n_1094;
wire n_1220;
wire n_696;
wire n_1147;
wire n_1425;
wire n_704;
wire n_453;
wire n_647;
wire n_948;
wire n_399;
wire n_700;
wire n_677;
wire n_1269;
wire n_378;
wire n_591;
wire n_1366;
wire n_678;
wire n_415;
wire n_1400;
wire n_564;
wire n_638;
wire n_510;
wire n_1361;
wire n_1358;
wire n_1406;
wire n_550;
wire n_966;
wire n_333;
wire n_1368;
wire n_994;
wire n_384;
wire n_1479;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_992;
wire n_813;
wire n_981;
wire n_1338;
wire n_1182;
wire n_872;
wire n_1401;
wire n_1086;
wire n_1070;
wire n_1189;
wire n_535;
wire n_882;
wire n_1210;
wire n_1456;
wire n_746;
wire n_656;
wire n_1148;
wire n_860;
wire n_748;
wire n_1261;
wire n_1062;
wire n_1439;
wire n_651;
wire n_801;
wire n_1271;
wire n_529;
wire n_504;
wire n_973;
wire n_1364;
wire n_659;
wire n_634;
wire n_903;
wire n_565;
wire n_925;
wire n_1389;
wire n_1393;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_311;
wire n_278;
wire n_1362;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_277;
wire n_754;
wire n_508;
wire n_1141;
wire n_1112;
wire n_1408;
wire n_428;
wire n_783;
wire n_1107;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1386;
wire n_406;
wire n_617;
wire n_602;
wire n_402;
wire n_733;
wire n_1404;
wire n_658;
wire n_676;
wire n_531;
wire n_1031;
wire n_1394;
wire n_807;
wire n_255;
wire n_286;
wire n_1011;
wire n_416;
wire n_895;
wire n_799;
wire n_490;
wire n_261;
wire n_391;
wire n_695;
wire n_1181;
wire n_881;
wire n_1145;
wire n_645;
wire n_557;
wire n_985;
wire n_777;
wire n_910;
wire n_642;
wire n_613;
wire n_1125;
wire n_296;
wire n_1347;
wire n_1163;
wire n_1278;
wire n_734;
wire n_735;
wire n_334;
wire n_1179;
wire n_569;
wire n_1171;
wire n_785;
wire n_1203;
wire n_1232;
wire n_471;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1187;
wire n_1000;
wire n_649;
wire n_358;
wire n_1234;
wire n_622;
wire n_1002;
wire n_1353;
wire n_1165;
wire n_1058;
wire n_1216;
wire n_662;
wire n_850;
wire n_265;
wire n_720;
wire n_354;
wire n_1026;
wire n_492;
wire n_407;
wire n_419;
wire n_1023;
wire n_730;
wire n_643;
wire n_1403;
wire n_486;
wire n_291;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_365;
wire n_526;
wire n_268;
wire n_1194;
wire n_282;
wire n_389;
wire n_1462;
wire n_701;
wire n_809;
wire n_679;
wire n_520;
wire n_926;
wire n_942;
wire n_1374;
wire n_1120;
wire n_689;
wire n_946;
wire n_300;
wire n_753;
wire n_1409;
wire n_1188;
wire n_623;
wire n_1032;
wire n_1474;
wire n_1431;
wire n_721;
wire n_1133;
wire n_313;
wire n_739;
wire n_1322;
wire n_1162;
wire n_1463;
wire n_762;
wire n_325;
wire n_1298;
wire n_442;
wire n_740;
wire n_1357;
wire n_639;
wire n_1186;
wire n_1365;
wire n_253;
wire n_459;
wire n_1172;
wire n_998;
wire n_1395;
wire n_1276;
wire n_836;
wire n_1184;
wire n_583;
wire n_347;
wire n_414;
wire n_1336;
wire n_279;
wire n_776;
wire n_1138;
wire n_890;
wire n_1306;
wire n_1413;
wire n_1266;
wire n_497;
wire n_911;
wire n_450;
wire n_473;
wire n_967;
wire n_474;
wire n_1159;
wire n_1315;
wire n_1055;
wire n_611;
wire n_380;
wire n_844;
wire n_968;
wire n_710;
wire n_1040;
wire n_307;
wire n_1102;
wire n_661;
wire n_1185;
wire n_447;
wire n_403;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1069;
wire n_1451;
wire n_842;
wire n_798;
wire n_668;
wire n_862;
wire n_869;
wire n_1066;
wire n_257;
wire n_285;
wire n_1377;
wire n_800;
wire n_1170;
wire n_778;
wire n_1175;
wire n_522;
wire n_1475;
wire n_943;
wire n_977;
wire n_287;
wire n_357;
wire n_905;
wire n_386;
wire n_878;
wire n_1333;
wire n_577;
wire n_759;
wire n_1235;
wire n_299;
wire n_322;
wire n_900;
wire n_841;
wire n_318;
wire n_1218;
wire n_736;
wire n_766;
wire n_1113;
wire n_852;
wire n_1268;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_1302;
wire n_1289;
wire n_937;
wire n_1442;
wire n_773;
wire n_353;
wire n_1446;
wire n_865;
wire n_856;
wire n_594;
wire n_1146;
wire n_1435;
wire n_374;
wire n_932;
wire n_958;
wire n_775;
wire n_763;
wire n_1093;
wire n_427;
wire n_519;
wire n_1116;
wire n_709;
wire n_388;
wire n_332;
wire n_1470;
wire n_816;
wire n_625;
wire n_953;
wire n_289;
wire n_1373;
wire n_716;
wire n_356;
wire n_584;
wire n_896;
wire n_528;
wire n_1078;
wire n_495;
wire n_1072;
wire n_370;
wire n_352;
wire n_935;
wire n_467;
wire n_1213;
wire n_1053;
wire n_263;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_284;
wire n_316;
wire n_1168;
wire n_1309;
wire n_909;
wire n_996;
wire n_523;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1332;
wire n_1411;
wire n_1263;
wire n_1115;
wire n_310;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_454;
wire n_1303;
wire n_1471;
wire n_443;
wire n_1029;
wire n_345;
wire n_1207;
wire n_324;
wire n_664;
wire n_367;
wire n_267;
wire n_1017;
wire n_581;
wire n_936;
wire n_1215;
wire n_582;
wire n_641;
wire n_940;
wire n_745;
wire n_339;
wire n_1167;
wire n_1327;
wire n_609;
wire n_1006;
wire n_1259;
wire n_350;
wire n_561;
wire n_437;
wire n_405;
wire n_1223;
wire n_621;
wire n_1012;
wire n_1241;
wire n_1414;
wire n_502;
wire n_769;
wire n_434;
wire n_250;
wire n_1455;
wire n_1212;
wire n_1054;
wire n_1308;
wire n_1050;
wire n_426;
wire n_1134;
wire n_1319;
wire n_1363;
wire n_616;
wire n_880;
wire n_1103;
wire n_1274;
wire n_832;
wire n_1321;
wire n_1429;
wire n_1060;
wire n_1154;
wire n_361;
wire n_632;
wire n_1344;
wire n_1450;
wire n_714;
wire n_1331;
wire n_1222;
wire n_1041;
wire n_251;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_1335;
wire n_1405;
wire n_912;
wire n_464;
wire n_1227;
wire n_945;
wire n_392;
wire n_288;
wire n_274;
wire n_303;
wire n_563;
wire n_891;
wire n_568;
wire n_413;
wire n_1157;
wire n_902;
wire n_1158;
wire n_1079;
wire n_1330;
wire n_1033;
wire n_1464;
wire n_1028;
wire n_366;
wire n_727;
wire n_1083;
wire n_397;
wire n_1056;
wire n_663;
wire n_588;
wire n_1448;
wire n_707;
wire n_915;
wire n_1001;
wire n_1418;
wire n_711;
wire n_864;
wire n_1169;
wire n_377;
wire n_1139;
wire n_273;
wire n_1038;
wire n_276;
wire n_1085;
wire n_295;
wire n_845;
wire n_1127;
wire n_484;
wire n_326;
wire n_893;
wire n_1068;
wire n_747;
wire n_1244;
wire n_697;
wire n_978;
wire n_847;
wire n_1452;
wire n_826;
wire n_373;
wire n_628;
wire n_487;
wire n_831;
wire n_653;
wire n_692;
wire n_1433;
wire n_1051;
wire n_1355;
wire n_309;
wire n_827;
wire n_472;
wire n_866;
wire n_452;
wire n_262;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_1426;
wire n_858;
wire n_764;
wire n_252;
wire n_741;
wire n_1090;
wire n_456;
wire n_359;
wire n_1469;
wire n_1164;
wire n_433;
wire n_627;
wire n_418;
wire n_771;
wire n_524;
wire n_1378;
wire n_705;
wire n_1191;
wire n_1206;
wire n_1270;
wire n_1399;
wire n_546;
wire n_1010;
wire n_1375;
wire n_1015;
wire n_863;
wire n_525;
wire n_1226;
wire n_644;
wire n_1150;
wire n_1341;
wire n_833;
wire n_1229;
wire n_929;
wire n_1143;
wire n_1190;
wire n_543;
wire n_305;
wire n_585;
wire n_1457;
wire n_465;
wire n_719;
wire n_1343;
wire n_1156;
wire n_988;
wire n_1466;
wire n_1396;
wire n_921;
wire n_640;
wire n_1176;
wire n_1151;
wire n_1254;
wire n_1458;
wire n_646;
wire n_1211;
wire n_650;
wire n_743;
wire n_823;
wire n_393;
wire n_294;
wire n_1480;
wire n_1101;
wire n_1076;
wire n_1251;
wire n_1434;
wire n_1461;
wire n_1449;
wire n_1407;
wire n_1104;
wire n_849;
wire n_1061;
wire n_554;
wire n_1153;
wire n_1337;
wire n_797;
wire n_1177;
wire n_758;
wire n_436;
wire n_390;
wire n_1096;
wire n_1316;
wire n_1420;
wire n_1092;
wire n_846;
wire n_631;
wire n_673;
wire n_1410;
wire n_1067;
wire n_518;
wire n_1192;
wire n_1292;
wire n_1478;
wire n_1240;
wire n_987;
wire n_362;
wire n_1065;
wire n_540;
wire n_1064;
wire n_1075;
wire n_718;
wire n_669;
wire n_1091;
wire n_423;
wire n_1221;
wire n_458;
wire n_1200;
wire n_444;
wire n_319;
wire n_364;
wire n_555;
wire n_1295;
wire n_974;
wire n_1329;
wire n_857;
wire n_1424;
wire n_376;
wire n_308;
wire n_491;
wire n_1294;
wire n_1110;
wire n_1137;
wire n_460;
wire n_317;
wire n_321;
wire n_666;
wire n_320;
wire n_660;
wire n_1359;
wire n_886;
wire n_767;
wire n_889;
wire n_1398;
wire n_379;
wire n_1432;
wire n_1021;
wire n_1297;
wire n_1046;
wire n_1109;
wire n_961;
wire n_1447;
wire n_489;
wire n_1381;
wire n_573;
wire n_1099;
wire n_626;
wire n_539;
wire n_462;
wire n_280;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_1272;
wire n_408;
wire n_372;
wire n_578;
wire n_892;
wire n_938;
wire n_327;
wire n_774;
wire n_466;
wire n_1049;
wire n_559;
wire n_1277;
wire n_984;
wire n_301;
wire n_726;
wire n_369;
wire n_517;
wire n_931;
wire n_780;
wire n_530;
wire n_834;
wire n_693;
wire n_496;
wire n_1360;
wire n_1082;
wire n_1257;
wire n_468;
wire n_1025;
wire n_532;
wire n_298;
wire n_924;
wire n_1264;
wire n_297;
wire n_1245;
wire n_1152;
wire n_1081;
wire n_547;
wire n_1324;
wire n_1198;
wire n_304;
wire n_1307;
wire n_993;
wire n_819;
wire n_737;
wire n_1290;
wire n_1318;
wire n_1135;
wire n_1063;
wire n_828;
wire n_770;
wire n_867;
wire n_398;
wire n_1100;
wire n_425;
wire n_879;
wire n_331;
wire n_449;
wire n_1340;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_1443;
wire n_655;
wire n_654;
wire n_672;
wire n_567;
wire n_916;
wire n_1354;
wire n_1334;
wire n_1291;
wire n_1437;
wire n_1473;
wire n_986;
wire n_451;
wire n_1037;
wire n_1267;
wire n_790;
wire n_1262;
wire n_410;
wire n_1444;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_1356;
wire n_768;
wire n_412;
wire n_542;
wire n_1256;
wire n_1427;
wire n_1077;
wire n_1111;
wire n_1249;
wire n_1416;
wire n_387;
wire n_1239;
wire n_969;
wire n_256;
wire n_1009;
wire n_1202;
wire n_302;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_269;
wire n_430;
wire n_1252;
wire n_1132;
wire n_1275;
wire n_843;
wire n_579;
wire n_533;
wire n_1472;
wire n_385;
wire n_275;
wire n_536;
wire n_470;
wire n_851;
wire n_1155;
wire n_934;
wire n_1027;
wire n_965;
wire n_1296;
wire n_382;
wire n_1043;
wire n_435;
wire n_511;
wire n_1467;
wire n_509;
wire n_1204;
wire n_930;
wire n_1265;
wire n_1057;
wire n_907;
wire n_1430;
wire n_1005;
wire n_1312;
wire n_899;
wire n_637;
wire n_544;
wire n_1476;
wire n_1087;
wire n_344;
wire n_482;
wire n_633;
wire n_971;
wire n_1052;
wire n_1071;
wire n_1311;
wire n_1438;
wire n_1273;
wire n_959;
wire n_349;
wire n_336;
wire n_1130;
wire n_794;
wire n_283;
wire n_314;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1253;
wire n_312;
wire n_1183;
wire n_335;
wire n_516;
wire n_1460;
wire n_521;
wire n_1195;
wire n_575;
wire n_1300;
wire n_338;
wire n_1372;
wire n_698;
wire n_371;
wire n_1345;
wire n_587;
wire n_1428;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_1436;
wire n_793;
wire n_1390;
wire n_272;
wire n_1412;
wire n_757;
wire n_803;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1088;
wire n_1230;
wire n_1326;
wire n_1402;
wire n_1388;
wire n_340;
wire n_483;
wire n_394;
wire n_1352;
wire n_729;
wire n_1280;
wire n_1323;
wire n_703;
wire n_1097;
wire n_1369;
wire n_601;
wire n_463;
wire n_396;
wire n_1236;
wire n_342;
wire n_348;
wire n_603;
wire n_1288;
wire n_868;
wire n_1024;
wire n_259;
wire n_1144;
wire n_475;
wire n_897;
wire n_1320;
wire n_855;
wire n_429;
INVx1_ASAP7_75t_L g697 ( .A(n_0), .Y(n_697) );
INVx1_ASAP7_75t_L g808 ( .A(n_1), .Y(n_808) );
AOI22xp33_ASAP7_75t_L g1209 ( .A1(n_2), .A2(n_6), .B1(n_1167), .B2(n_1170), .Y(n_1209) );
OAI211xp5_ASAP7_75t_L g780 ( .A1(n_3), .A2(n_481), .B(n_665), .C(n_781), .Y(n_780) );
INVx1_ASAP7_75t_L g800 ( .A(n_3), .Y(n_800) );
AOI221x1_ASAP7_75t_SL g820 ( .A1(n_4), .A2(n_241), .B1(n_821), .B2(n_823), .C(n_824), .Y(n_820) );
AOI21xp33_ASAP7_75t_L g886 ( .A1(n_4), .A2(n_346), .B(n_887), .Y(n_886) );
INVx1_ASAP7_75t_L g576 ( .A(n_5), .Y(n_576) );
OAI211xp5_ASAP7_75t_L g619 ( .A1(n_5), .A2(n_620), .B(n_622), .C(n_631), .Y(n_619) );
XNOR2xp5_ASAP7_75t_L g1059 ( .A(n_7), .B(n_1060), .Y(n_1059) );
AOI221xp5_ASAP7_75t_L g1349 ( .A1(n_8), .A2(n_195), .B1(n_333), .B2(n_1350), .C(n_1351), .Y(n_1349) );
INVx1_ASAP7_75t_L g1395 ( .A(n_8), .Y(n_1395) );
INVx1_ASAP7_75t_L g528 ( .A(n_9), .Y(n_528) );
INVx1_ASAP7_75t_L g1352 ( .A(n_10), .Y(n_1352) );
AOI221xp5_ASAP7_75t_L g1396 ( .A1(n_10), .A2(n_136), .B1(n_415), .B2(n_1393), .C(n_1397), .Y(n_1396) );
INVx1_ASAP7_75t_L g907 ( .A(n_11), .Y(n_907) );
OAI211xp5_ASAP7_75t_L g947 ( .A1(n_11), .A2(n_483), .B(n_545), .C(n_948), .Y(n_947) );
INVx1_ASAP7_75t_L g1431 ( .A(n_12), .Y(n_1431) );
OAI22xp33_ASAP7_75t_L g1468 ( .A1(n_12), .A2(n_112), .B1(n_1469), .B2(n_1472), .Y(n_1468) );
INVx1_ASAP7_75t_L g259 ( .A(n_13), .Y(n_259) );
AND2x2_ASAP7_75t_L g390 ( .A(n_13), .B(n_391), .Y(n_390) );
AND2x2_ASAP7_75t_L g413 ( .A(n_13), .B(n_211), .Y(n_413) );
NOR2xp33_ASAP7_75t_L g510 ( .A(n_13), .B(n_269), .Y(n_510) );
OAI211xp5_ASAP7_75t_L g457 ( .A1(n_14), .A2(n_458), .B(n_459), .C(n_468), .Y(n_457) );
INVx1_ASAP7_75t_L g490 ( .A(n_14), .Y(n_490) );
OAI221xp5_ASAP7_75t_L g1434 ( .A1(n_15), .A2(n_242), .B1(n_1435), .B2(n_1438), .C(n_1439), .Y(n_1434) );
INVx1_ASAP7_75t_L g1464 ( .A(n_15), .Y(n_1464) );
OAI22xp33_ASAP7_75t_L g995 ( .A1(n_16), .A2(n_189), .B1(n_497), .B2(n_996), .Y(n_995) );
OAI22xp33_ASAP7_75t_L g1008 ( .A1(n_16), .A2(n_189), .B1(n_444), .B2(n_1009), .Y(n_1008) );
INVx1_ASAP7_75t_L g1068 ( .A(n_17), .Y(n_1068) );
INVx1_ASAP7_75t_L g1093 ( .A(n_18), .Y(n_1093) );
INVx2_ASAP7_75t_L g1163 ( .A(n_19), .Y(n_1163) );
AND2x2_ASAP7_75t_L g1165 ( .A(n_19), .B(n_93), .Y(n_1165) );
AND2x2_ASAP7_75t_L g1171 ( .A(n_19), .B(n_1169), .Y(n_1171) );
OAI22xp5_ASAP7_75t_L g443 ( .A1(n_20), .A2(n_141), .B1(n_444), .B2(n_448), .Y(n_443) );
OAI22xp5_ASAP7_75t_L g494 ( .A1(n_20), .A2(n_141), .B1(n_495), .B2(n_497), .Y(n_494) );
OAI22xp5_ASAP7_75t_L g842 ( .A1(n_21), .A2(n_125), .B1(n_843), .B2(n_846), .Y(n_842) );
OAI221xp5_ASAP7_75t_L g855 ( .A1(n_21), .A2(n_218), .B1(n_856), .B2(n_858), .C(n_860), .Y(n_855) );
OAI22xp33_ASAP7_75t_L g1136 ( .A1(n_22), .A2(n_237), .B1(n_670), .B2(n_1137), .Y(n_1136) );
OAI22xp33_ASAP7_75t_L g1147 ( .A1(n_22), .A2(n_237), .B1(n_802), .B2(n_912), .Y(n_1147) );
INVx1_ASAP7_75t_L g1023 ( .A(n_23), .Y(n_1023) );
AOI22xp5_ASAP7_75t_L g1173 ( .A1(n_24), .A2(n_217), .B1(n_1167), .B2(n_1170), .Y(n_1173) );
XNOR2x2_ASAP7_75t_L g1339 ( .A(n_24), .B(n_1340), .Y(n_1339) );
AOI22xp33_ASAP7_75t_L g1412 ( .A1(n_24), .A2(n_1413), .B1(n_1415), .B2(n_1475), .Y(n_1412) );
OAI22xp33_ASAP7_75t_L g669 ( .A1(n_25), .A2(n_54), .B1(n_670), .B2(n_671), .Y(n_669) );
OAI22xp33_ASAP7_75t_L g682 ( .A1(n_25), .A2(n_54), .B1(n_683), .B2(n_684), .Y(n_682) );
OAI22xp33_ASAP7_75t_L g454 ( .A1(n_26), .A2(n_37), .B1(n_261), .B2(n_455), .Y(n_454) );
OAI22xp33_ASAP7_75t_L g472 ( .A1(n_26), .A2(n_37), .B1(n_473), .B2(n_477), .Y(n_472) );
OAI211xp5_ASAP7_75t_L g1091 ( .A1(n_27), .A2(n_483), .B(n_769), .C(n_1092), .Y(n_1091) );
INVx1_ASAP7_75t_L g1100 ( .A(n_27), .Y(n_1100) );
INVx1_ASAP7_75t_L g1108 ( .A(n_28), .Y(n_1108) );
INVx1_ASAP7_75t_L g961 ( .A(n_29), .Y(n_961) );
OAI22xp5_ASAP7_75t_L g1130 ( .A1(n_30), .A2(n_115), .B1(n_1089), .B2(n_1131), .Y(n_1130) );
OAI22xp5_ASAP7_75t_L g1140 ( .A1(n_30), .A2(n_115), .B1(n_455), .B2(n_1141), .Y(n_1140) );
OAI22xp33_ASAP7_75t_L g779 ( .A1(n_31), .A2(n_162), .B1(n_475), .B2(n_660), .Y(n_779) );
OAI22xp33_ASAP7_75t_L g790 ( .A1(n_31), .A2(n_162), .B1(n_261), .B2(n_687), .Y(n_790) );
INVx1_ASAP7_75t_L g930 ( .A(n_32), .Y(n_930) );
INVx1_ASAP7_75t_L g435 ( .A(n_33), .Y(n_435) );
AOI22xp5_ASAP7_75t_L g1179 ( .A1(n_33), .A2(n_244), .B1(n_1160), .B2(n_1180), .Y(n_1179) );
INVx1_ASAP7_75t_L g525 ( .A(n_34), .Y(n_525) );
AOI22xp33_ASAP7_75t_L g604 ( .A1(n_35), .A2(n_219), .B1(n_605), .B2(n_607), .Y(n_604) );
INVx1_ASAP7_75t_L g623 ( .A(n_35), .Y(n_623) );
INVx1_ASAP7_75t_L g759 ( .A(n_36), .Y(n_759) );
INVx1_ASAP7_75t_L g906 ( .A(n_38), .Y(n_906) );
INVx1_ASAP7_75t_L g1354 ( .A(n_39), .Y(n_1354) );
AOI221xp5_ASAP7_75t_L g1388 ( .A1(n_39), .A2(n_71), .B1(n_1389), .B2(n_1391), .C(n_1394), .Y(n_1388) );
CKINVDCx5p33_ASAP7_75t_R g362 ( .A(n_40), .Y(n_362) );
AOI22xp33_ASAP7_75t_L g316 ( .A1(n_41), .A2(n_75), .B1(n_317), .B2(n_318), .Y(n_316) );
INVx1_ASAP7_75t_L g417 ( .A(n_41), .Y(n_417) );
OAI22xp5_ASAP7_75t_L g908 ( .A1(n_42), .A2(n_143), .B1(n_455), .B2(n_909), .Y(n_908) );
OAI22xp5_ASAP7_75t_L g945 ( .A1(n_42), .A2(n_143), .B1(n_658), .B2(n_946), .Y(n_945) );
AOI22xp5_ASAP7_75t_L g1183 ( .A1(n_43), .A2(n_232), .B1(n_1167), .B2(n_1170), .Y(n_1183) );
AO22x1_ASAP7_75t_L g1159 ( .A1(n_44), .A2(n_58), .B1(n_1160), .B2(n_1164), .Y(n_1159) );
AOI22xp33_ASAP7_75t_SL g594 ( .A1(n_45), .A2(n_102), .B1(n_595), .B2(n_597), .Y(n_594) );
AOI22xp33_ASAP7_75t_L g635 ( .A1(n_45), .A2(n_219), .B1(n_369), .B2(n_630), .Y(n_635) );
OAI221xp5_ASAP7_75t_L g1370 ( .A1(n_46), .A2(n_64), .B1(n_856), .B2(n_858), .C(n_1371), .Y(n_1370) );
INVxp67_ASAP7_75t_SL g1380 ( .A(n_46), .Y(n_1380) );
INVx1_ASAP7_75t_L g667 ( .A(n_47), .Y(n_667) );
AOI221xp5_ASAP7_75t_L g1425 ( .A1(n_48), .A2(n_122), .B1(n_1426), .B2(n_1427), .C(n_1428), .Y(n_1425) );
AOI22xp33_ASAP7_75t_L g1462 ( .A1(n_48), .A2(n_78), .B1(n_335), .B2(n_596), .Y(n_1462) );
AOI22xp33_ASAP7_75t_L g1429 ( .A1(n_49), .A2(n_149), .B1(n_617), .B2(n_836), .Y(n_1429) );
AOI22xp33_ASAP7_75t_L g1461 ( .A1(n_49), .A2(n_94), .B1(n_333), .B2(n_925), .Y(n_1461) );
INVx1_ASAP7_75t_L g521 ( .A(n_50), .Y(n_521) );
INVx1_ASAP7_75t_L g284 ( .A(n_51), .Y(n_284) );
INVx1_ASAP7_75t_L g301 ( .A(n_51), .Y(n_301) );
INVx1_ASAP7_75t_L g603 ( .A(n_52), .Y(n_603) );
AOI22xp33_ASAP7_75t_L g629 ( .A1(n_52), .A2(n_228), .B1(n_369), .B2(n_630), .Y(n_629) );
INVx1_ASAP7_75t_L g749 ( .A(n_53), .Y(n_749) );
INVx1_ASAP7_75t_L g1094 ( .A(n_55), .Y(n_1094) );
OAI211xp5_ASAP7_75t_L g1098 ( .A1(n_55), .A2(n_676), .B(n_1013), .C(n_1099), .Y(n_1098) );
CKINVDCx5p33_ASAP7_75t_R g828 ( .A(n_56), .Y(n_828) );
OAI22xp33_ASAP7_75t_L g1049 ( .A1(n_57), .A2(n_182), .B1(n_477), .B2(n_1050), .Y(n_1049) );
OAI22xp33_ASAP7_75t_L g1052 ( .A1(n_57), .A2(n_182), .B1(n_261), .B2(n_1053), .Y(n_1052) );
OAI22xp5_ASAP7_75t_L g571 ( .A1(n_58), .A2(n_572), .B1(n_573), .B2(n_651), .Y(n_571) );
INVxp67_ASAP7_75t_L g651 ( .A(n_58), .Y(n_651) );
INVx1_ASAP7_75t_L g253 ( .A(n_59), .Y(n_253) );
OAI22xp5_ASAP7_75t_L g1365 ( .A1(n_60), .A2(n_201), .B1(n_1366), .B2(n_1368), .Y(n_1365) );
INVx1_ASAP7_75t_L g1387 ( .A(n_60), .Y(n_1387) );
INVx2_ASAP7_75t_L g292 ( .A(n_61), .Y(n_292) );
INVx1_ASAP7_75t_L g964 ( .A(n_62), .Y(n_964) );
OAI22xp5_ASAP7_75t_L g1343 ( .A1(n_63), .A2(n_174), .B1(n_1344), .B2(n_1347), .Y(n_1343) );
INVx1_ASAP7_75t_L g1382 ( .A(n_63), .Y(n_1382) );
INVx1_ASAP7_75t_L g1405 ( .A(n_64), .Y(n_1405) );
XOR2x2_ASAP7_75t_L g654 ( .A(n_65), .B(n_655), .Y(n_654) );
AOI22xp5_ASAP7_75t_L g1184 ( .A1(n_65), .A2(n_165), .B1(n_1160), .B2(n_1164), .Y(n_1184) );
OAI22xp5_ASAP7_75t_L g1449 ( .A1(n_66), .A2(n_208), .B1(n_431), .B2(n_1450), .Y(n_1449) );
INVx1_ASAP7_75t_L g536 ( .A(n_67), .Y(n_536) );
INVx1_ASAP7_75t_L g1028 ( .A(n_68), .Y(n_1028) );
INVx1_ASAP7_75t_L g1448 ( .A(n_69), .Y(n_1448) );
AO221x2_ASAP7_75t_L g1210 ( .A1(n_70), .A2(n_207), .B1(n_1167), .B2(n_1170), .C(n_1211), .Y(n_1210) );
AOI221xp5_ASAP7_75t_L g1356 ( .A1(n_71), .A2(n_196), .B1(n_333), .B2(n_1357), .C(n_1359), .Y(n_1356) );
OAI211xp5_ASAP7_75t_L g902 ( .A1(n_72), .A2(n_903), .B(n_904), .C(n_905), .Y(n_902) );
INVx1_ASAP7_75t_L g949 ( .A(n_72), .Y(n_949) );
XNOR2xp5_ASAP7_75t_L g1416 ( .A(n_73), .B(n_1417), .Y(n_1416) );
INVxp67_ASAP7_75t_SL g577 ( .A(n_74), .Y(n_577) );
OAI221xp5_ASAP7_75t_L g639 ( .A1(n_74), .A2(n_198), .B1(n_640), .B2(n_641), .C(n_645), .Y(n_639) );
AOI221xp5_ASAP7_75t_L g366 ( .A1(n_75), .A2(n_114), .B1(n_367), .B2(n_373), .C(n_376), .Y(n_366) );
INVx1_ASAP7_75t_L g467 ( .A(n_76), .Y(n_467) );
OAI211xp5_ASAP7_75t_L g480 ( .A1(n_76), .A2(n_481), .B(n_483), .C(n_485), .Y(n_480) );
INVx1_ASAP7_75t_L g713 ( .A(n_77), .Y(n_713) );
INVxp67_ASAP7_75t_SL g1442 ( .A(n_78), .Y(n_1442) );
XOR2x2_ASAP7_75t_L g437 ( .A(n_79), .B(n_438), .Y(n_437) );
INVx1_ASAP7_75t_L g784 ( .A(n_80), .Y(n_784) );
OAI211xp5_ASAP7_75t_L g791 ( .A1(n_80), .A2(n_792), .B(n_793), .C(n_797), .Y(n_791) );
INVx1_ASAP7_75t_L g974 ( .A(n_81), .Y(n_974) );
CKINVDCx5p33_ASAP7_75t_R g357 ( .A(n_82), .Y(n_357) );
INVx1_ASAP7_75t_L g764 ( .A(n_83), .Y(n_764) );
INVx1_ASAP7_75t_L g763 ( .A(n_84), .Y(n_763) );
INVx1_ASAP7_75t_L g1001 ( .A(n_85), .Y(n_1001) );
CKINVDCx5p33_ASAP7_75t_R g583 ( .A(n_86), .Y(n_583) );
OA222x2_ASAP7_75t_L g810 ( .A1(n_87), .A2(n_191), .B1(n_218), .B2(n_811), .C1(n_814), .C2(n_818), .Y(n_810) );
INVx1_ASAP7_75t_L g872 ( .A(n_87), .Y(n_872) );
INVx1_ASAP7_75t_L g1115 ( .A(n_88), .Y(n_1115) );
AOI22xp5_ASAP7_75t_L g898 ( .A1(n_89), .A2(n_899), .B1(n_900), .B2(n_953), .Y(n_898) );
INVxp67_ASAP7_75t_SL g953 ( .A(n_89), .Y(n_953) );
HB1xp67_ASAP7_75t_L g255 ( .A(n_90), .Y(n_255) );
AND2x2_ASAP7_75t_L g1161 ( .A(n_90), .B(n_253), .Y(n_1161) );
INVx1_ASAP7_75t_L g1111 ( .A(n_91), .Y(n_1111) );
CKINVDCx5p33_ASAP7_75t_R g344 ( .A(n_92), .Y(n_344) );
AND2x2_ASAP7_75t_L g1162 ( .A(n_93), .B(n_1163), .Y(n_1162) );
INVx1_ASAP7_75t_L g1169 ( .A(n_93), .Y(n_1169) );
AOI221xp5_ASAP7_75t_L g1443 ( .A1(n_94), .A2(n_140), .B1(n_633), .B2(n_634), .C(n_1389), .Y(n_1443) );
AOI22xp33_ASAP7_75t_L g321 ( .A1(n_95), .A2(n_98), .B1(n_322), .B2(n_326), .Y(n_321) );
INVx1_ASAP7_75t_L g421 ( .A(n_95), .Y(n_421) );
OAI211xp5_ASAP7_75t_SL g997 ( .A1(n_96), .A2(n_483), .B(n_998), .C(n_1000), .Y(n_997) );
INVx1_ASAP7_75t_L g1016 ( .A(n_96), .Y(n_1016) );
INVx1_ASAP7_75t_L g303 ( .A(n_97), .Y(n_303) );
OAI22xp5_ASAP7_75t_L g401 ( .A1(n_97), .A2(n_220), .B1(n_402), .B2(n_403), .Y(n_401) );
INVx1_ASAP7_75t_L g382 ( .A(n_98), .Y(n_382) );
INVx1_ASAP7_75t_L g708 ( .A(n_99), .Y(n_708) );
INVx1_ASAP7_75t_L g1112 ( .A(n_100), .Y(n_1112) );
INVx1_ASAP7_75t_L g1109 ( .A(n_101), .Y(n_1109) );
AOI21xp33_ASAP7_75t_L g625 ( .A1(n_102), .A2(n_626), .B(n_628), .Y(n_625) );
OAI211xp5_ASAP7_75t_L g1132 ( .A1(n_103), .A2(n_663), .B(n_665), .C(n_1133), .Y(n_1132) );
INVx1_ASAP7_75t_L g1146 ( .A(n_103), .Y(n_1146) );
NAND2xp5_ASAP7_75t_L g291 ( .A(n_104), .B(n_292), .Y(n_291) );
INVx2_ASAP7_75t_L g312 ( .A(n_104), .Y(n_312) );
INVx1_ASAP7_75t_L g341 ( .A(n_104), .Y(n_341) );
OAI22xp33_ASAP7_75t_L g785 ( .A1(n_105), .A2(n_225), .B1(n_670), .B2(n_786), .Y(n_785) );
OAI22xp5_ASAP7_75t_L g801 ( .A1(n_105), .A2(n_225), .B1(n_802), .B2(n_803), .Y(n_801) );
INVx1_ASAP7_75t_L g1025 ( .A(n_106), .Y(n_1025) );
OAI22xp33_ASAP7_75t_L g657 ( .A1(n_107), .A2(n_243), .B1(n_658), .B2(n_660), .Y(n_657) );
OAI22xp33_ASAP7_75t_L g686 ( .A1(n_107), .A2(n_243), .B1(n_261), .B2(n_687), .Y(n_686) );
AOI22xp33_ASAP7_75t_L g1208 ( .A1(n_108), .A2(n_202), .B1(n_1160), .B2(n_1164), .Y(n_1208) );
INVx1_ASAP7_75t_L g916 ( .A(n_109), .Y(n_916) );
INVx1_ASAP7_75t_L g1070 ( .A(n_110), .Y(n_1070) );
INVx1_ASAP7_75t_L g1135 ( .A(n_111), .Y(n_1135) );
OAI211xp5_ASAP7_75t_L g1144 ( .A1(n_111), .A2(n_522), .B(n_793), .C(n_1145), .Y(n_1144) );
INVx1_ASAP7_75t_L g1432 ( .A(n_112), .Y(n_1432) );
OAI211xp5_ASAP7_75t_L g1041 ( .A1(n_113), .A2(n_483), .B(n_1042), .C(n_1044), .Y(n_1041) );
INVx1_ASAP7_75t_L g1057 ( .A(n_113), .Y(n_1057) );
AOI22xp33_ASAP7_75t_SL g334 ( .A1(n_114), .A2(n_142), .B1(n_317), .B2(n_335), .Y(n_334) );
AOI22xp33_ASAP7_75t_L g835 ( .A1(n_116), .A2(n_240), .B1(n_617), .B2(n_836), .Y(n_835) );
AOI22xp33_ASAP7_75t_L g888 ( .A1(n_116), .A2(n_222), .B1(n_327), .B2(n_889), .Y(n_888) );
INVx1_ASAP7_75t_L g1064 ( .A(n_117), .Y(n_1064) );
INVx1_ASAP7_75t_L g587 ( .A(n_118), .Y(n_587) );
OAI22xp5_ASAP7_75t_L g611 ( .A1(n_118), .A2(n_150), .B1(n_612), .B2(n_615), .Y(n_611) );
INVx1_ASAP7_75t_L g926 ( .A(n_119), .Y(n_926) );
INVx1_ASAP7_75t_L g968 ( .A(n_120), .Y(n_968) );
INVx1_ASAP7_75t_L g1026 ( .A(n_121), .Y(n_1026) );
AOI22xp33_ASAP7_75t_L g1454 ( .A1(n_122), .A2(n_157), .B1(n_1455), .B2(n_1457), .Y(n_1454) );
INVx1_ASAP7_75t_L g1033 ( .A(n_123), .Y(n_1033) );
INVx1_ASAP7_75t_L g1077 ( .A(n_124), .Y(n_1077) );
INVx1_ASAP7_75t_L g873 ( .A(n_125), .Y(n_873) );
OAI22xp33_ASAP7_75t_L g1095 ( .A1(n_126), .A2(n_144), .B1(n_786), .B2(n_996), .Y(n_1095) );
OAI22xp5_ASAP7_75t_L g1101 ( .A1(n_126), .A2(n_144), .B1(n_684), .B2(n_802), .Y(n_1101) );
INVx1_ASAP7_75t_L g1363 ( .A(n_127), .Y(n_1363) );
CKINVDCx5p33_ASAP7_75t_R g602 ( .A(n_128), .Y(n_602) );
CKINVDCx5p33_ASAP7_75t_R g834 ( .A(n_129), .Y(n_834) );
INVx1_ASAP7_75t_L g535 ( .A(n_130), .Y(n_535) );
INVx1_ASAP7_75t_L g752 ( .A(n_131), .Y(n_752) );
INVx1_ASAP7_75t_L g591 ( .A(n_132), .Y(n_591) );
AOI21xp33_ASAP7_75t_L g632 ( .A1(n_132), .A2(n_633), .B(n_634), .Y(n_632) );
INVx1_ASAP7_75t_L g754 ( .A(n_133), .Y(n_754) );
INVx1_ASAP7_75t_L g1114 ( .A(n_134), .Y(n_1114) );
AO22x1_ASAP7_75t_L g1166 ( .A1(n_135), .A2(n_215), .B1(n_1167), .B2(n_1170), .Y(n_1166) );
INVx1_ASAP7_75t_L g1360 ( .A(n_136), .Y(n_1360) );
BUFx3_ASAP7_75t_L g286 ( .A(n_137), .Y(n_286) );
INVx1_ASAP7_75t_L g929 ( .A(n_138), .Y(n_929) );
INVx1_ASAP7_75t_L g1045 ( .A(n_139), .Y(n_1045) );
AOI22xp33_ASAP7_75t_L g1458 ( .A1(n_140), .A2(n_149), .B1(n_322), .B2(n_1459), .Y(n_1458) );
AOI211xp5_ASAP7_75t_SL g414 ( .A1(n_142), .A2(n_415), .B(n_416), .C(n_420), .Y(n_414) );
AOI22xp33_ASAP7_75t_L g1189 ( .A1(n_145), .A2(n_159), .B1(n_1167), .B2(n_1170), .Y(n_1189) );
BUFx6f_ASAP7_75t_L g266 ( .A(n_146), .Y(n_266) );
AOI22xp33_ASAP7_75t_L g329 ( .A1(n_147), .A2(n_176), .B1(n_330), .B2(n_333), .Y(n_329) );
INVx1_ASAP7_75t_L g381 ( .A(n_147), .Y(n_381) );
INVx1_ASAP7_75t_L g1022 ( .A(n_148), .Y(n_1022) );
INVx1_ASAP7_75t_L g586 ( .A(n_150), .Y(n_586) );
INVx1_ASAP7_75t_L g1078 ( .A(n_151), .Y(n_1078) );
INVx1_ASAP7_75t_L g1046 ( .A(n_152), .Y(n_1046) );
OAI211xp5_ASAP7_75t_L g1055 ( .A1(n_152), .A2(n_904), .B(n_1013), .C(n_1056), .Y(n_1055) );
INVx1_ASAP7_75t_L g1119 ( .A(n_153), .Y(n_1119) );
INVx1_ASAP7_75t_L g1072 ( .A(n_154), .Y(n_1072) );
XNOR2xp5_ASAP7_75t_L g956 ( .A(n_155), .B(n_957), .Y(n_956) );
INVx1_ASAP7_75t_L g668 ( .A(n_156), .Y(n_668) );
OAI211xp5_ASAP7_75t_L g674 ( .A1(n_156), .A2(n_675), .B(n_676), .C(n_677), .Y(n_674) );
INVxp67_ASAP7_75t_SL g1440 ( .A(n_157), .Y(n_1440) );
INVx1_ASAP7_75t_L g512 ( .A(n_158), .Y(n_512) );
OAI22xp33_ASAP7_75t_L g1003 ( .A1(n_160), .A2(n_235), .B1(n_473), .B2(n_1004), .Y(n_1003) );
OAI22xp5_ASAP7_75t_L g1006 ( .A1(n_160), .A2(n_235), .B1(n_455), .B2(n_1007), .Y(n_1006) );
XNOR2xp5_ASAP7_75t_L g1017 ( .A(n_161), .B(n_1018), .Y(n_1017) );
CKINVDCx5p33_ASAP7_75t_R g293 ( .A(n_163), .Y(n_293) );
INVx1_ASAP7_75t_L g1032 ( .A(n_164), .Y(n_1032) );
INVx1_ASAP7_75t_L g462 ( .A(n_166), .Y(n_462) );
AOI22xp5_ASAP7_75t_L g1174 ( .A1(n_167), .A2(n_231), .B1(n_1160), .B2(n_1164), .Y(n_1174) );
INVx1_ASAP7_75t_L g746 ( .A(n_168), .Y(n_746) );
INVx1_ASAP7_75t_L g695 ( .A(n_169), .Y(n_695) );
INVx1_ASAP7_75t_L g703 ( .A(n_170), .Y(n_703) );
INVx1_ASAP7_75t_L g962 ( .A(n_171), .Y(n_962) );
XOR2x2_ASAP7_75t_L g739 ( .A(n_172), .B(n_740), .Y(n_739) );
INVx1_ASAP7_75t_L g970 ( .A(n_173), .Y(n_970) );
INVxp67_ASAP7_75t_SL g1401 ( .A(n_174), .Y(n_1401) );
OAI211xp5_ASAP7_75t_L g661 ( .A1(n_175), .A2(n_662), .B(n_665), .C(n_666), .Y(n_661) );
INVx1_ASAP7_75t_L g681 ( .A(n_175), .Y(n_681) );
INVx1_ASAP7_75t_L g424 ( .A(n_176), .Y(n_424) );
INVx1_ASAP7_75t_L g783 ( .A(n_177), .Y(n_783) );
INVx1_ASAP7_75t_L g1030 ( .A(n_178), .Y(n_1030) );
INVx1_ASAP7_75t_L g1002 ( .A(n_179), .Y(n_1002) );
OAI211xp5_ASAP7_75t_L g1012 ( .A1(n_179), .A2(n_904), .B(n_1013), .C(n_1015), .Y(n_1012) );
INVx1_ASAP7_75t_L g516 ( .A(n_180), .Y(n_516) );
INVx1_ASAP7_75t_L g923 ( .A(n_181), .Y(n_923) );
AOI22xp33_ASAP7_75t_L g1188 ( .A1(n_183), .A2(n_227), .B1(n_1160), .B2(n_1164), .Y(n_1188) );
INVx1_ASAP7_75t_L g1073 ( .A(n_184), .Y(n_1073) );
INVx1_ASAP7_75t_L g700 ( .A(n_185), .Y(n_700) );
BUFx6f_ASAP7_75t_L g265 ( .A(n_186), .Y(n_265) );
INVx1_ASAP7_75t_L g918 ( .A(n_187), .Y(n_918) );
INVx1_ASAP7_75t_L g935 ( .A(n_188), .Y(n_935) );
OAI22xp33_ASAP7_75t_L g1088 ( .A1(n_190), .A2(n_206), .B1(n_660), .B2(n_1089), .Y(n_1088) );
OAI22xp33_ASAP7_75t_L g1097 ( .A1(n_190), .A2(n_206), .B1(n_261), .B2(n_1053), .Y(n_1097) );
INVx1_ASAP7_75t_L g861 ( .A(n_191), .Y(n_861) );
INVx1_ASAP7_75t_L g582 ( .A(n_192), .Y(n_582) );
INVx1_ASAP7_75t_L g973 ( .A(n_193), .Y(n_973) );
CKINVDCx5p33_ASAP7_75t_R g848 ( .A(n_194), .Y(n_848) );
INVx1_ASAP7_75t_L g1398 ( .A(n_195), .Y(n_1398) );
INVx1_ASAP7_75t_L g1399 ( .A(n_196), .Y(n_1399) );
OAI22xp33_ASAP7_75t_L g910 ( .A1(n_197), .A2(n_214), .B1(n_911), .B2(n_912), .Y(n_910) );
OAI22xp33_ASAP7_75t_L g950 ( .A1(n_197), .A2(n_214), .B1(n_497), .B2(n_951), .Y(n_950) );
INVx1_ASAP7_75t_L g580 ( .A(n_198), .Y(n_580) );
AO22x1_ASAP7_75t_L g1204 ( .A1(n_199), .A2(n_216), .B1(n_1160), .B2(n_1205), .Y(n_1204) );
CKINVDCx16_ASAP7_75t_R g1212 ( .A(n_200), .Y(n_1212) );
INVxp67_ASAP7_75t_SL g1374 ( .A(n_201), .Y(n_1374) );
INVx1_ASAP7_75t_L g1066 ( .A(n_203), .Y(n_1066) );
INVx1_ASAP7_75t_L g710 ( .A(n_204), .Y(n_710) );
INVx1_ASAP7_75t_L g758 ( .A(n_205), .Y(n_758) );
OAI211xp5_ASAP7_75t_L g1421 ( .A1(n_208), .A2(n_1422), .B(n_1424), .C(n_1430), .Y(n_1421) );
OAI22xp33_ASAP7_75t_L g1047 ( .A1(n_209), .A2(n_248), .B1(n_497), .B2(n_1048), .Y(n_1047) );
OAI22xp33_ASAP7_75t_L g1054 ( .A1(n_209), .A2(n_248), .B1(n_444), .B2(n_1009), .Y(n_1054) );
AOI22xp5_ASAP7_75t_L g1178 ( .A1(n_210), .A2(n_238), .B1(n_1167), .B2(n_1170), .Y(n_1178) );
BUFx3_ASAP7_75t_L g269 ( .A(n_211), .Y(n_269) );
INVx1_ASAP7_75t_L g391 ( .A(n_211), .Y(n_391) );
XOR2x2_ASAP7_75t_L g1103 ( .A(n_212), .B(n_1104), .Y(n_1103) );
CKINVDCx20_ASAP7_75t_R g1214 ( .A(n_213), .Y(n_1214) );
INVx1_ASAP7_75t_L g429 ( .A(n_220), .Y(n_429) );
INVx1_ASAP7_75t_L g523 ( .A(n_221), .Y(n_523) );
INVx1_ASAP7_75t_L g825 ( .A(n_222), .Y(n_825) );
CKINVDCx5p33_ASAP7_75t_R g833 ( .A(n_223), .Y(n_833) );
INVx1_ASAP7_75t_L g934 ( .A(n_224), .Y(n_934) );
INVx1_ASAP7_75t_L g1134 ( .A(n_226), .Y(n_1134) );
INVx1_ASAP7_75t_L g593 ( .A(n_228), .Y(n_593) );
INVx1_ASAP7_75t_L g290 ( .A(n_229), .Y(n_290) );
INVx2_ASAP7_75t_L g315 ( .A(n_229), .Y(n_315) );
INVx1_ASAP7_75t_L g352 ( .A(n_229), .Y(n_352) );
INVx1_ASAP7_75t_L g716 ( .A(n_230), .Y(n_716) );
INVx1_ASAP7_75t_L g1361 ( .A(n_233), .Y(n_1361) );
INVx1_ASAP7_75t_L g1117 ( .A(n_234), .Y(n_1117) );
CKINVDCx5p33_ASAP7_75t_R g851 ( .A(n_236), .Y(n_851) );
AO22x1_ASAP7_75t_L g1206 ( .A1(n_239), .A2(n_246), .B1(n_1167), .B2(n_1170), .Y(n_1206) );
INVx1_ASAP7_75t_L g884 ( .A(n_240), .Y(n_884) );
INVx1_ASAP7_75t_L g883 ( .A(n_241), .Y(n_883) );
INVx1_ASAP7_75t_L g1466 ( .A(n_242), .Y(n_1466) );
CKINVDCx5p33_ASAP7_75t_R g309 ( .A(n_245), .Y(n_309) );
INVx1_ASAP7_75t_L g965 ( .A(n_247), .Y(n_965) );
AOI21xp5_ASAP7_75t_L g249 ( .A1(n_250), .A2(n_270), .B(n_1151), .Y(n_249) );
AND2x2_ASAP7_75t_L g250 ( .A(n_251), .B(n_256), .Y(n_250) );
INVx1_ASAP7_75t_L g1411 ( .A(n_251), .Y(n_1411) );
NOR2xp33_ASAP7_75t_L g251 ( .A(n_252), .B(n_254), .Y(n_251) );
NOR2xp33_ASAP7_75t_L g1414 ( .A(n_252), .B(n_255), .Y(n_1414) );
INVx1_ASAP7_75t_L g1478 ( .A(n_252), .Y(n_1478) );
HB1xp67_ASAP7_75t_L g252 ( .A(n_253), .Y(n_252) );
INVx1_ASAP7_75t_L g254 ( .A(n_255), .Y(n_254) );
NOR2xp33_ASAP7_75t_L g1480 ( .A(n_255), .B(n_1478), .Y(n_1480) );
NAND2xp5_ASAP7_75t_L g256 ( .A(n_257), .B(n_260), .Y(n_256) );
INVx1_ASAP7_75t_L g257 ( .A(n_258), .Y(n_257) );
AND2x4_ASAP7_75t_L g440 ( .A(n_258), .B(n_441), .Y(n_440) );
NOR2xp33_ASAP7_75t_L g1410 ( .A(n_258), .B(n_1411), .Y(n_1410) );
INVx1_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
AND2x4_ASAP7_75t_L g386 ( .A(n_259), .B(n_268), .Y(n_386) );
AND2x4_ASAP7_75t_L g419 ( .A(n_259), .B(n_269), .Y(n_419) );
INVx1_ASAP7_75t_L g909 ( .A(n_260), .Y(n_909) );
INVxp67_ASAP7_75t_SL g1007 ( .A(n_260), .Y(n_1007) );
AND2x4_ASAP7_75t_SL g1409 ( .A(n_260), .B(n_1410), .Y(n_1409) );
INVx3_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
OR2x6_ASAP7_75t_L g261 ( .A(n_262), .B(n_267), .Y(n_261) );
OR2x6_ASAP7_75t_L g446 ( .A(n_262), .B(n_447), .Y(n_446) );
BUFx4f_ASAP7_75t_L g712 ( .A(n_262), .Y(n_712) );
INVxp67_ASAP7_75t_L g748 ( .A(n_262), .Y(n_748) );
INVx1_ASAP7_75t_L g991 ( .A(n_262), .Y(n_991) );
INVx2_ASAP7_75t_L g262 ( .A(n_263), .Y(n_262) );
INVx3_ASAP7_75t_L g402 ( .A(n_263), .Y(n_402) );
BUFx4f_ASAP7_75t_L g423 ( .A(n_263), .Y(n_423) );
INVx3_ASAP7_75t_L g263 ( .A(n_264), .Y(n_263) );
OR2x2_ASAP7_75t_L g264 ( .A(n_265), .B(n_266), .Y(n_264) );
INVx2_ASAP7_75t_L g371 ( .A(n_265), .Y(n_371) );
INVx2_ASAP7_75t_L g375 ( .A(n_265), .Y(n_375) );
NAND2x1_ASAP7_75t_L g380 ( .A(n_265), .B(n_266), .Y(n_380) );
AND2x2_ASAP7_75t_L g396 ( .A(n_265), .B(n_397), .Y(n_396) );
AND2x2_ASAP7_75t_L g400 ( .A(n_265), .B(n_266), .Y(n_400) );
INVx1_ASAP7_75t_L g466 ( .A(n_265), .Y(n_466) );
INVx1_ASAP7_75t_L g372 ( .A(n_266), .Y(n_372) );
AND2x2_ASAP7_75t_L g374 ( .A(n_266), .B(n_375), .Y(n_374) );
OR2x2_ASAP7_75t_L g385 ( .A(n_266), .B(n_371), .Y(n_385) );
INVx2_ASAP7_75t_L g397 ( .A(n_266), .Y(n_397) );
NAND2xp5_ASAP7_75t_L g404 ( .A(n_266), .B(n_375), .Y(n_404) );
BUFx2_ASAP7_75t_L g409 ( .A(n_266), .Y(n_409) );
OR2x6_ASAP7_75t_L g1143 ( .A(n_267), .B(n_402), .Y(n_1143) );
INVxp67_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
INVx1_ASAP7_75t_L g470 ( .A(n_268), .Y(n_470) );
INVx2_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
BUFx2_ASAP7_75t_L g453 ( .A(n_269), .Y(n_453) );
AND2x4_ASAP7_75t_L g464 ( .A(n_269), .B(n_465), .Y(n_464) );
XNOR2xp5_ASAP7_75t_L g270 ( .A(n_271), .B(n_893), .Y(n_270) );
XNOR2xp5_ASAP7_75t_L g271 ( .A(n_272), .B(n_568), .Y(n_271) );
AOI22xp33_ASAP7_75t_L g272 ( .A1(n_273), .A2(n_274), .B1(n_436), .B2(n_437), .Y(n_272) );
INVx1_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
INVx1_ASAP7_75t_L g274 ( .A(n_275), .Y(n_274) );
XNOR2x1_ASAP7_75t_L g275 ( .A(n_276), .B(n_435), .Y(n_275) );
OR2x2_ASAP7_75t_L g276 ( .A(n_277), .B(n_347), .Y(n_276) );
NAND3xp33_ASAP7_75t_L g277 ( .A(n_278), .B(n_310), .C(n_343), .Y(n_277) );
AOI222xp33_ASAP7_75t_L g278 ( .A1(n_279), .A2(n_293), .B1(n_294), .B2(n_303), .C1(n_304), .C2(n_309), .Y(n_278) );
INVx2_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
AND2x4_ASAP7_75t_L g1450 ( .A(n_280), .B(n_846), .Y(n_1450) );
OR2x2_ASAP7_75t_L g280 ( .A(n_281), .B(n_287), .Y(n_280) );
INVx4_ASAP7_75t_L g482 ( .A(n_281), .Y(n_482) );
INVx3_ASAP7_75t_L g664 ( .A(n_281), .Y(n_664) );
BUFx6f_ASAP7_75t_L g921 ( .A(n_281), .Y(n_921) );
BUFx6f_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
BUFx3_ASAP7_75t_L g547 ( .A(n_282), .Y(n_547) );
BUFx2_ASAP7_75t_L g771 ( .A(n_282), .Y(n_771) );
NAND2x1p5_ASAP7_75t_L g282 ( .A(n_283), .B(n_285), .Y(n_282) );
BUFx2_ASAP7_75t_L g493 ( .A(n_283), .Y(n_493) );
INVx1_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
NAND2xp5_ASAP7_75t_L g308 ( .A(n_284), .B(n_286), .Y(n_308) );
INVx2_ASAP7_75t_L g320 ( .A(n_284), .Y(n_320) );
AND2x4_ASAP7_75t_L g327 ( .A(n_285), .B(n_328), .Y(n_327) );
INVx2_ASAP7_75t_L g356 ( .A(n_285), .Y(n_356) );
BUFx2_ASAP7_75t_L g489 ( .A(n_285), .Y(n_489) );
BUFx6f_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
INVx2_ASAP7_75t_L g298 ( .A(n_286), .Y(n_298) );
AND2x4_ASAP7_75t_L g319 ( .A(n_286), .B(n_320), .Y(n_319) );
OR2x2_ASAP7_75t_L g476 ( .A(n_286), .B(n_300), .Y(n_476) );
INVx1_ASAP7_75t_L g302 ( .A(n_287), .Y(n_302) );
OR2x2_ASAP7_75t_L g305 ( .A(n_287), .B(n_306), .Y(n_305) );
INVx1_ASAP7_75t_L g1471 ( .A(n_287), .Y(n_1471) );
OR2x2_ASAP7_75t_L g287 ( .A(n_288), .B(n_291), .Y(n_287) );
HB1xp67_ASAP7_75t_L g505 ( .A(n_288), .Y(n_505) );
INVx1_ASAP7_75t_L g533 ( .A(n_288), .Y(n_533) );
OR2x2_ASAP7_75t_L g539 ( .A(n_288), .B(n_540), .Y(n_539) );
INVx2_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
BUFx2_ASAP7_75t_L g434 ( .A(n_289), .Y(n_434) );
INVx1_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
INVx1_ASAP7_75t_L g876 ( .A(n_291), .Y(n_876) );
INVx1_ASAP7_75t_L g1346 ( .A(n_291), .Y(n_1346) );
BUFx3_ASAP7_75t_L g313 ( .A(n_292), .Y(n_313) );
INVx3_ASAP7_75t_L g342 ( .A(n_292), .Y(n_342) );
NAND2xp33_ASAP7_75t_SL g540 ( .A(n_292), .B(n_312), .Y(n_540) );
AOI22xp33_ASAP7_75t_L g408 ( .A1(n_293), .A2(n_357), .B1(n_409), .B2(n_410), .Y(n_408) );
AND2x4_ASAP7_75t_L g294 ( .A(n_295), .B(n_302), .Y(n_294) );
INVx2_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
INVx8_ASAP7_75t_L g317 ( .A(n_296), .Y(n_317) );
CKINVDCx5p33_ASAP7_75t_R g862 ( .A(n_296), .Y(n_862) );
INVx3_ASAP7_75t_L g889 ( .A(n_296), .Y(n_889) );
INVx2_ASAP7_75t_L g1350 ( .A(n_296), .Y(n_1350) );
INVx8_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
NAND2x1p5_ASAP7_75t_L g432 ( .A(n_297), .B(n_353), .Y(n_432) );
BUFx3_ASAP7_75t_L g596 ( .A(n_297), .Y(n_596) );
HB1xp67_ASAP7_75t_L g868 ( .A(n_297), .Y(n_868) );
AND2x2_ASAP7_75t_L g1345 ( .A(n_297), .B(n_1346), .Y(n_1345) );
AND2x4_ASAP7_75t_L g297 ( .A(n_298), .B(n_299), .Y(n_297) );
AND2x4_ASAP7_75t_L g324 ( .A(n_298), .B(n_325), .Y(n_324) );
INVx1_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
INVx1_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
INVxp67_ASAP7_75t_L g325 ( .A(n_301), .Y(n_325) );
AND2x4_ASAP7_75t_L g345 ( .A(n_302), .B(n_346), .Y(n_345) );
INVx1_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
AND2x4_ASAP7_75t_L g1447 ( .A(n_305), .B(n_813), .Y(n_1447) );
INVx1_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
BUFx6f_ASAP7_75t_L g553 ( .A(n_307), .Y(n_553) );
INVx1_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
BUFx2_ASAP7_75t_L g499 ( .A(n_308), .Y(n_499) );
A2O1A1Ixp33_ASAP7_75t_L g405 ( .A1(n_309), .A2(n_369), .B(n_406), .C(n_412), .Y(n_405) );
AOI33xp33_ASAP7_75t_L g310 ( .A1(n_311), .A2(n_316), .A3(n_321), .B1(n_329), .B2(n_334), .B3(n_337), .Y(n_310) );
AOI33xp33_ASAP7_75t_L g1453 ( .A1(n_311), .A2(n_337), .A3(n_1454), .B1(n_1458), .B2(n_1461), .B3(n_1462), .Y(n_1453) );
AND3x4_ASAP7_75t_L g311 ( .A(n_312), .B(n_313), .C(n_314), .Y(n_311) );
INVx1_ASAP7_75t_L g354 ( .A(n_312), .Y(n_354) );
HB1xp67_ASAP7_75t_L g503 ( .A(n_312), .Y(n_503) );
AND2x2_ASAP7_75t_L g1355 ( .A(n_312), .B(n_313), .Y(n_1355) );
INVx3_ASAP7_75t_L g488 ( .A(n_313), .Y(n_488) );
INVx1_ASAP7_75t_L g427 ( .A(n_314), .Y(n_427) );
INVx2_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
BUFx2_ASAP7_75t_L g339 ( .A(n_315), .Y(n_339) );
NAND2xp5_ASAP7_75t_L g841 ( .A(n_315), .B(n_413), .Y(n_841) );
AOI22xp33_ASAP7_75t_L g871 ( .A1(n_318), .A2(n_326), .B1(n_872), .B2(n_873), .Y(n_871) );
BUFx2_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
INVx2_ASAP7_75t_L g336 ( .A(n_319), .Y(n_336) );
BUFx2_ASAP7_75t_L g364 ( .A(n_319), .Y(n_364) );
AND2x4_ASAP7_75t_L g484 ( .A(n_319), .B(n_342), .Y(n_484) );
BUFx2_ASAP7_75t_L g584 ( .A(n_319), .Y(n_584) );
BUFx3_ASAP7_75t_L g863 ( .A(n_319), .Y(n_863) );
AND2x2_ASAP7_75t_L g1348 ( .A(n_319), .B(n_1346), .Y(n_1348) );
BUFx2_ASAP7_75t_L g1457 ( .A(n_319), .Y(n_1457) );
INVx1_ASAP7_75t_L g328 ( .A(n_320), .Y(n_328) );
INVx1_ASAP7_75t_L g776 ( .A(n_322), .Y(n_776) );
INVx1_ASAP7_75t_L g1124 ( .A(n_322), .Y(n_1124) );
BUFx6f_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
AND2x4_ASAP7_75t_L g478 ( .A(n_323), .B(n_479), .Y(n_478) );
BUFx6f_ASAP7_75t_L g728 ( .A(n_323), .Y(n_728) );
INVx2_ASAP7_75t_L g1128 ( .A(n_323), .Y(n_1128) );
BUFx6f_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
BUFx6f_ASAP7_75t_L g332 ( .A(n_324), .Y(n_332) );
BUFx8_ASAP7_75t_L g346 ( .A(n_324), .Y(n_346) );
INVx2_ASAP7_75t_L g551 ( .A(n_324), .Y(n_551) );
BUFx3_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
BUFx3_ASAP7_75t_L g333 ( .A(n_327), .Y(n_333) );
AND2x4_ASAP7_75t_L g1369 ( .A(n_327), .B(n_876), .Y(n_1369) );
INVx5_ASAP7_75t_L g1460 ( .A(n_327), .Y(n_1460) );
INVx1_ASAP7_75t_L g361 ( .A(n_328), .Y(n_361) );
INVx2_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
INVx2_ASAP7_75t_SL g331 ( .A(n_332), .Y(n_331) );
HB1xp67_ASAP7_75t_L g556 ( .A(n_332), .Y(n_556) );
INVx5_ASAP7_75t_L g733 ( .A(n_332), .Y(n_733) );
INVx3_ASAP7_75t_L g870 ( .A(n_332), .Y(n_870) );
INVx2_ASAP7_75t_SL g1353 ( .A(n_332), .Y(n_1353) );
INVx1_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
INVx1_ASAP7_75t_L g597 ( .A(n_336), .Y(n_597) );
INVx1_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
OAI33xp33_ASAP7_75t_L g1120 ( .A1(n_338), .A2(n_720), .A3(n_1121), .B1(n_1123), .B2(n_1125), .B3(n_1127), .Y(n_1120) );
OR2x6_ASAP7_75t_L g338 ( .A(n_339), .B(n_340), .Y(n_338) );
AND2x4_ASAP7_75t_L g509 ( .A(n_339), .B(n_510), .Y(n_509) );
INVx1_ASAP7_75t_L g891 ( .A(n_339), .Y(n_891) );
INVx3_ASAP7_75t_L g881 ( .A(n_340), .Y(n_881) );
NAND2x1p5_ASAP7_75t_L g340 ( .A(n_341), .B(n_342), .Y(n_340) );
NAND3x1_ASAP7_75t_L g566 ( .A(n_341), .B(n_342), .C(n_567), .Y(n_566) );
AND2x4_ASAP7_75t_L g353 ( .A(n_342), .B(n_354), .Y(n_353) );
OR2x4_ASAP7_75t_L g475 ( .A(n_342), .B(n_476), .Y(n_475) );
INVx1_ASAP7_75t_L g479 ( .A(n_342), .Y(n_479) );
OR2x6_ASAP7_75t_L g498 ( .A(n_342), .B(n_499), .Y(n_498) );
NAND2xp5_ASAP7_75t_L g343 ( .A(n_344), .B(n_345), .Y(n_343) );
AOI221xp5_ASAP7_75t_L g392 ( .A1(n_344), .A2(n_362), .B1(n_393), .B2(n_398), .C(n_401), .Y(n_392) );
INVx2_ASAP7_75t_L g1472 ( .A(n_345), .Y(n_1472) );
INVx3_ASAP7_75t_L g928 ( .A(n_346), .Y(n_928) );
INVx3_ASAP7_75t_L g1029 ( .A(n_346), .Y(n_1029) );
INVx2_ASAP7_75t_SL g1358 ( .A(n_346), .Y(n_1358) );
NAND3xp33_ASAP7_75t_SL g347 ( .A(n_348), .B(n_365), .C(n_428), .Y(n_347) );
AOI221xp5_ASAP7_75t_L g348 ( .A1(n_349), .A2(n_357), .B1(n_358), .B2(n_362), .C(n_363), .Y(n_348) );
AND2x4_ASAP7_75t_SL g349 ( .A(n_350), .B(n_355), .Y(n_349) );
AND2x4_ASAP7_75t_SL g358 ( .A(n_350), .B(n_359), .Y(n_358) );
AND2x4_ASAP7_75t_L g363 ( .A(n_350), .B(n_364), .Y(n_363) );
AND2x2_ASAP7_75t_L g1465 ( .A(n_350), .B(n_355), .Y(n_1465) );
AND2x4_ASAP7_75t_L g1467 ( .A(n_350), .B(n_359), .Y(n_1467) );
AND2x4_ASAP7_75t_L g350 ( .A(n_351), .B(n_353), .Y(n_350) );
OR2x2_ASAP7_75t_L g813 ( .A(n_351), .B(n_640), .Y(n_813) );
INVx1_ASAP7_75t_L g1385 ( .A(n_351), .Y(n_1385) );
INVx1_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
INVx1_ASAP7_75t_L g567 ( .A(n_352), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g817 ( .A(n_352), .B(n_390), .Y(n_817) );
AND2x6_ASAP7_75t_L g857 ( .A(n_353), .B(n_355), .Y(n_857) );
AND2x2_ASAP7_75t_L g859 ( .A(n_353), .B(n_361), .Y(n_859) );
INVx1_ASAP7_75t_L g865 ( .A(n_353), .Y(n_865) );
INVx3_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
INVx2_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
INVx3_ASAP7_75t_L g1474 ( .A(n_363), .Y(n_1474) );
OAI31xp33_ASAP7_75t_L g365 ( .A1(n_366), .A2(n_387), .A3(n_414), .B(n_427), .Y(n_365) );
INVx1_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
INVx3_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
BUFx6f_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
AND2x2_ASAP7_75t_L g614 ( .A(n_370), .B(n_390), .Y(n_614) );
NAND2xp5_ASAP7_75t_L g640 ( .A(n_370), .B(n_413), .Y(n_640) );
INVx3_ASAP7_75t_L g837 ( .A(n_370), .Y(n_837) );
AND2x2_ASAP7_75t_L g370 ( .A(n_371), .B(n_372), .Y(n_370) );
HB1xp67_ASAP7_75t_L g411 ( .A(n_371), .Y(n_411) );
BUFx3_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
INVx2_ASAP7_75t_L g618 ( .A(n_374), .Y(n_618) );
BUFx6f_ASAP7_75t_L g630 ( .A(n_374), .Y(n_630) );
OAI221xp5_ASAP7_75t_L g376 ( .A1(n_377), .A2(n_381), .B1(n_382), .B2(n_383), .C(n_386), .Y(n_376) );
INVx2_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
INVx1_ASAP7_75t_L g458 ( .A(n_378), .Y(n_458) );
INVx1_ASAP7_75t_L g792 ( .A(n_378), .Y(n_792) );
INVx4_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
BUFx4f_ASAP7_75t_L g522 ( .A(n_379), .Y(n_522) );
BUFx4f_ASAP7_75t_L g675 ( .A(n_379), .Y(n_675) );
BUFx4f_ASAP7_75t_L g709 ( .A(n_379), .Y(n_709) );
OR2x6_ASAP7_75t_L g838 ( .A(n_379), .B(n_839), .Y(n_838) );
BUFx4f_ASAP7_75t_L g903 ( .A(n_379), .Y(n_903) );
BUFx6f_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
BUFx3_ASAP7_75t_L g407 ( .A(n_380), .Y(n_407) );
INVx2_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
INVx2_ASAP7_75t_L g520 ( .A(n_384), .Y(n_520) );
INVx2_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
BUFx3_ASAP7_75t_L g418 ( .A(n_385), .Y(n_418) );
BUFx2_ASAP7_75t_L g707 ( .A(n_385), .Y(n_707) );
INVx1_ASAP7_75t_L g757 ( .A(n_385), .Y(n_757) );
INVx3_ASAP7_75t_L g634 ( .A(n_386), .Y(n_634) );
OAI21xp33_ASAP7_75t_L g387 ( .A1(n_388), .A2(n_392), .B(n_405), .Y(n_387) );
INVxp67_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
BUFx2_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
AND2x2_ASAP7_75t_L g616 ( .A(n_390), .B(n_617), .Y(n_616) );
AND2x4_ASAP7_75t_L g621 ( .A(n_390), .B(n_395), .Y(n_621) );
AND2x4_ASAP7_75t_SL g638 ( .A(n_390), .B(n_399), .Y(n_638) );
AND2x2_ASAP7_75t_L g853 ( .A(n_390), .B(n_395), .Y(n_853) );
AND2x4_ASAP7_75t_L g1423 ( .A(n_390), .B(n_630), .Y(n_1423) );
HB1xp67_ASAP7_75t_L g447 ( .A(n_391), .Y(n_447) );
INVx2_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
INVx2_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
BUFx6f_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
AND2x4_ASAP7_75t_L g456 ( .A(n_396), .B(n_447), .Y(n_456) );
INVx2_ASAP7_75t_L g627 ( .A(n_396), .Y(n_627) );
BUFx3_ASAP7_75t_L g1393 ( .A(n_396), .Y(n_1393) );
BUFx2_ASAP7_75t_L g823 ( .A(n_398), .Y(n_823) );
BUFx6f_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
BUFx3_ASAP7_75t_L g415 ( .A(n_399), .Y(n_415) );
AND2x2_ASAP7_75t_L g469 ( .A(n_399), .B(n_470), .Y(n_469) );
AND2x6_ASAP7_75t_L g648 ( .A(n_399), .B(n_413), .Y(n_648) );
INVx1_ASAP7_75t_L g1390 ( .A(n_399), .Y(n_1390) );
BUFx3_ASAP7_75t_L g1426 ( .A(n_399), .Y(n_1426) );
BUFx6f_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
INVx1_ASAP7_75t_L g796 ( .A(n_400), .Y(n_796) );
BUFx3_ASAP7_75t_L g515 ( .A(n_402), .Y(n_515) );
BUFx3_ASAP7_75t_L g696 ( .A(n_402), .Y(n_696) );
INVx2_ASAP7_75t_SL g762 ( .A(n_402), .Y(n_762) );
INVx8_ASAP7_75t_L g426 ( .A(n_403), .Y(n_426) );
OR2x2_ASAP7_75t_L g452 ( .A(n_403), .B(n_453), .Y(n_452) );
BUFx2_ASAP7_75t_L g1441 ( .A(n_403), .Y(n_1441) );
BUFx6f_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
NAND2xp5_ASAP7_75t_L g406 ( .A(n_407), .B(n_408), .Y(n_406) );
INVx2_ASAP7_75t_SL g527 ( .A(n_407), .Y(n_527) );
BUFx3_ASAP7_75t_L g624 ( .A(n_407), .Y(n_624) );
OR2x2_ASAP7_75t_L g818 ( .A(n_407), .B(n_817), .Y(n_818) );
BUFx2_ASAP7_75t_SL g1085 ( .A(n_407), .Y(n_1085) );
OR2x2_ASAP7_75t_L g1404 ( .A(n_407), .B(n_817), .Y(n_1404) );
AND2x4_ASAP7_75t_L g461 ( .A(n_409), .B(n_453), .Y(n_461) );
INVx1_ASAP7_75t_L g643 ( .A(n_409), .Y(n_643) );
AND2x2_ASAP7_75t_L g678 ( .A(n_409), .B(n_453), .Y(n_678) );
INVx1_ASAP7_75t_L g845 ( .A(n_409), .Y(n_845) );
INVx1_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
HB1xp67_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
INVx1_ASAP7_75t_L g644 ( .A(n_413), .Y(n_644) );
NAND2xp5_ASAP7_75t_L g647 ( .A(n_413), .B(n_465), .Y(n_647) );
OAI21xp33_ASAP7_75t_L g416 ( .A1(n_417), .A2(n_418), .B(n_419), .Y(n_416) );
INVx2_ASAP7_75t_L g702 ( .A(n_418), .Y(n_702) );
HB1xp67_ASAP7_75t_L g985 ( .A(n_418), .Y(n_985) );
OAI22xp5_ASAP7_75t_L g1036 ( .A1(n_418), .A2(n_903), .B1(n_1025), .B2(n_1028), .Y(n_1036) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_419), .B(n_532), .Y(n_531) );
INVx4_ASAP7_75t_L g628 ( .A(n_419), .Y(n_628) );
AND2x4_ASAP7_75t_L g718 ( .A(n_419), .B(n_532), .Y(n_718) );
INVx1_ASAP7_75t_SL g1428 ( .A(n_419), .Y(n_1428) );
OAI22xp5_ASAP7_75t_L g420 ( .A1(n_421), .A2(n_422), .B1(n_424), .B2(n_425), .Y(n_420) );
OAI22xp5_ASAP7_75t_L g1394 ( .A1(n_422), .A2(n_425), .B1(n_1361), .B2(n_1395), .Y(n_1394) );
INVx4_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
INVx3_ASAP7_75t_L g940 ( .A(n_423), .Y(n_940) );
BUFx6f_ASAP7_75t_L g979 ( .A(n_423), .Y(n_979) );
INVx2_ASAP7_75t_L g518 ( .A(n_425), .Y(n_518) );
INVx4_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
INVx2_ASAP7_75t_L g698 ( .A(n_426), .Y(n_698) );
BUFx6f_ASAP7_75t_L g715 ( .A(n_426), .Y(n_715) );
INVx2_ASAP7_75t_SL g750 ( .A(n_426), .Y(n_750) );
INVx2_ASAP7_75t_L g827 ( .A(n_426), .Y(n_827) );
INVx1_ASAP7_75t_L g993 ( .A(n_426), .Y(n_993) );
INVx1_ASAP7_75t_L g1081 ( .A(n_426), .Y(n_1081) );
BUFx2_ASAP7_75t_L g650 ( .A(n_427), .Y(n_650) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_429), .B(n_430), .Y(n_428) );
INVx5_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
OR2x6_ASAP7_75t_L g431 ( .A(n_432), .B(n_433), .Y(n_431) );
INVx2_ASAP7_75t_L g1364 ( .A(n_432), .Y(n_1364) );
INVxp67_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
INVx1_ASAP7_75t_L g441 ( .A(n_434), .Y(n_441) );
OR2x2_ASAP7_75t_L g846 ( .A(n_434), .B(n_647), .Y(n_846) );
INVx1_ASAP7_75t_L g850 ( .A(n_434), .Y(n_850) );
INVx1_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
OAI221xp5_ASAP7_75t_L g438 ( .A1(n_439), .A2(n_442), .B1(n_471), .B2(n_500), .C(n_506), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
BUFx2_ASAP7_75t_SL g688 ( .A(n_440), .Y(n_688) );
BUFx3_ASAP7_75t_L g804 ( .A(n_440), .Y(n_804) );
OAI31xp33_ASAP7_75t_L g901 ( .A1(n_440), .A2(n_902), .A3(n_908), .B(n_910), .Y(n_901) );
BUFx2_ASAP7_75t_L g1148 ( .A(n_440), .Y(n_1148) );
NOR3xp33_ASAP7_75t_L g442 ( .A(n_443), .B(n_454), .C(n_457), .Y(n_442) );
INVx1_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
INVx1_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
BUFx2_ASAP7_75t_L g683 ( .A(n_446), .Y(n_683) );
BUFx6f_ASAP7_75t_L g802 ( .A(n_446), .Y(n_802) );
HB1xp67_ASAP7_75t_L g911 ( .A(n_446), .Y(n_911) );
INVx2_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
INVx2_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
INVx2_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
INVx1_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
INVx2_ASAP7_75t_L g685 ( .A(n_452), .Y(n_685) );
BUFx2_ASAP7_75t_L g1011 ( .A(n_452), .Y(n_1011) );
INVx3_ASAP7_75t_SL g455 ( .A(n_456), .Y(n_455) );
INVx4_ASAP7_75t_L g687 ( .A(n_456), .Y(n_687) );
CKINVDCx16_ASAP7_75t_R g1053 ( .A(n_456), .Y(n_1053) );
AOI22xp33_ASAP7_75t_L g459 ( .A1(n_460), .A2(n_462), .B1(n_463), .B2(n_467), .Y(n_459) );
AOI22xp33_ASAP7_75t_L g905 ( .A1(n_460), .A2(n_463), .B1(n_906), .B2(n_907), .Y(n_905) );
AOI22xp33_ASAP7_75t_L g1015 ( .A1(n_460), .A2(n_679), .B1(n_1001), .B2(n_1016), .Y(n_1015) );
AOI22xp33_ASAP7_75t_L g1056 ( .A1(n_460), .A2(n_679), .B1(n_1045), .B2(n_1057), .Y(n_1056) );
BUFx3_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
AOI22xp33_ASAP7_75t_L g1145 ( .A1(n_461), .A2(n_464), .B1(n_1134), .B2(n_1146), .Y(n_1145) );
AOI22xp33_ASAP7_75t_L g485 ( .A1(n_462), .A2(n_486), .B1(n_490), .B2(n_491), .Y(n_485) );
BUFx3_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
INVx2_ASAP7_75t_L g680 ( .A(n_464), .Y(n_680) );
INVx2_ASAP7_75t_L g799 ( .A(n_464), .Y(n_799) );
INVx1_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
INVx3_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
INVx1_ASAP7_75t_L g676 ( .A(n_469), .Y(n_676) );
INVx1_ASAP7_75t_L g904 ( .A(n_469), .Y(n_904) );
AND2x2_ASAP7_75t_L g794 ( .A(n_470), .B(n_795), .Y(n_794) );
NOR3xp33_ASAP7_75t_L g471 ( .A(n_472), .B(n_480), .C(n_494), .Y(n_471) );
INVx2_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
AOI22xp33_ASAP7_75t_L g585 ( .A1(n_474), .A2(n_586), .B1(n_587), .B2(n_588), .Y(n_585) );
INVx2_ASAP7_75t_SL g474 ( .A(n_475), .Y(n_474) );
INVx2_ASAP7_75t_SL g659 ( .A(n_475), .Y(n_659) );
HB1xp67_ASAP7_75t_L g1050 ( .A(n_475), .Y(n_1050) );
INVx1_ASAP7_75t_L g1090 ( .A(n_475), .Y(n_1090) );
OR2x4_ASAP7_75t_L g496 ( .A(n_476), .B(n_479), .Y(n_496) );
BUFx4f_ASAP7_75t_L g544 ( .A(n_476), .Y(n_544) );
INVx2_ASAP7_75t_L g562 ( .A(n_476), .Y(n_562) );
BUFx3_ASAP7_75t_L g724 ( .A(n_476), .Y(n_724) );
BUFx3_ASAP7_75t_L g880 ( .A(n_476), .Y(n_880) );
INVx1_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
AOI22xp33_ASAP7_75t_L g575 ( .A1(n_478), .A2(n_576), .B1(n_577), .B2(n_578), .Y(n_575) );
INVx2_ASAP7_75t_L g660 ( .A(n_478), .Y(n_660) );
INVx2_ASAP7_75t_L g946 ( .A(n_478), .Y(n_946) );
INVx1_ASAP7_75t_L g1004 ( .A(n_478), .Y(n_1004) );
INVxp67_ASAP7_75t_L g1131 ( .A(n_478), .Y(n_1131) );
OAI22xp33_ASAP7_75t_L g777 ( .A1(n_481), .A2(n_749), .B1(n_759), .B2(n_767), .Y(n_777) );
INVx1_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
INVx1_ASAP7_75t_L g725 ( .A(n_482), .Y(n_725) );
INVx2_ASAP7_75t_L g738 ( .A(n_482), .Y(n_738) );
INVx2_ASAP7_75t_L g879 ( .A(n_482), .Y(n_879) );
INVx1_ASAP7_75t_L g1122 ( .A(n_482), .Y(n_1122) );
NAND4xp25_ASAP7_75t_L g574 ( .A(n_483), .B(n_575), .C(n_579), .D(n_585), .Y(n_574) );
CKINVDCx8_ASAP7_75t_R g483 ( .A(n_484), .Y(n_483) );
CKINVDCx8_ASAP7_75t_R g665 ( .A(n_484), .Y(n_665) );
AOI22xp33_ASAP7_75t_L g948 ( .A1(n_486), .A2(n_491), .B1(n_906), .B2(n_949), .Y(n_948) );
AOI22xp33_ASAP7_75t_L g1000 ( .A1(n_486), .A2(n_491), .B1(n_1001), .B2(n_1002), .Y(n_1000) );
AOI22xp33_ASAP7_75t_L g1044 ( .A1(n_486), .A2(n_491), .B1(n_1045), .B2(n_1046), .Y(n_1044) );
BUFx3_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
BUFx3_ASAP7_75t_L g581 ( .A(n_487), .Y(n_581) );
AND2x2_ASAP7_75t_L g487 ( .A(n_488), .B(n_489), .Y(n_487) );
AND2x4_ASAP7_75t_L g492 ( .A(n_488), .B(n_493), .Y(n_492) );
AND2x4_ASAP7_75t_L g782 ( .A(n_488), .B(n_489), .Y(n_782) );
AOI222xp33_ASAP7_75t_L g579 ( .A1(n_491), .A2(n_580), .B1(n_581), .B2(n_582), .C1(n_583), .C2(n_584), .Y(n_579) );
AOI22xp33_ASAP7_75t_L g1092 ( .A1(n_491), .A2(n_581), .B1(n_1093), .B2(n_1094), .Y(n_1092) );
BUFx6f_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
AOI22xp33_ASAP7_75t_SL g666 ( .A1(n_492), .A2(n_581), .B1(n_667), .B2(n_668), .Y(n_666) );
AOI22xp33_ASAP7_75t_L g781 ( .A1(n_492), .A2(n_782), .B1(n_783), .B2(n_784), .Y(n_781) );
AOI22xp33_ASAP7_75t_L g1133 ( .A1(n_492), .A2(n_782), .B1(n_1134), .B2(n_1135), .Y(n_1133) );
BUFx2_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
INVx2_ASAP7_75t_SL g588 ( .A(n_496), .Y(n_588) );
BUFx3_ASAP7_75t_L g670 ( .A(n_496), .Y(n_670) );
BUFx2_ASAP7_75t_L g996 ( .A(n_496), .Y(n_996) );
BUFx3_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
INVx2_ASAP7_75t_L g578 ( .A(n_498), .Y(n_578) );
INVx1_ASAP7_75t_L g672 ( .A(n_498), .Y(n_672) );
INVx1_ASAP7_75t_L g787 ( .A(n_498), .Y(n_787) );
INVx1_ASAP7_75t_L g731 ( .A(n_499), .Y(n_731) );
BUFx3_ASAP7_75t_L g966 ( .A(n_499), .Y(n_966) );
CKINVDCx14_ASAP7_75t_R g500 ( .A(n_501), .Y(n_500) );
AOI211xp5_ASAP7_75t_L g573 ( .A1(n_501), .A2(n_574), .B(n_589), .C(n_609), .Y(n_573) );
OAI31xp33_ASAP7_75t_L g656 ( .A1(n_501), .A2(n_657), .A3(n_661), .B(n_669), .Y(n_656) );
OAI31xp33_ASAP7_75t_L g1040 ( .A1(n_501), .A2(n_1041), .A3(n_1047), .B(n_1049), .Y(n_1040) );
AND2x4_ASAP7_75t_L g501 ( .A(n_502), .B(n_504), .Y(n_501) );
AND2x2_ASAP7_75t_L g788 ( .A(n_502), .B(n_504), .Y(n_788) );
AND2x2_ASAP7_75t_SL g952 ( .A(n_502), .B(n_504), .Y(n_952) );
AND2x2_ASAP7_75t_L g1138 ( .A(n_502), .B(n_504), .Y(n_1138) );
INVx1_ASAP7_75t_SL g502 ( .A(n_503), .Y(n_502) );
INVx1_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
NOR2xp33_ASAP7_75t_L g506 ( .A(n_507), .B(n_537), .Y(n_506) );
OAI33xp33_ASAP7_75t_L g507 ( .A1(n_508), .A2(n_511), .A3(n_519), .B1(n_524), .B2(n_529), .B3(n_534), .Y(n_507) );
INVx2_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
INVx4_ASAP7_75t_L g693 ( .A(n_509), .Y(n_693) );
INVx2_ASAP7_75t_L g744 ( .A(n_509), .Y(n_744) );
INVx1_ASAP7_75t_L g830 ( .A(n_509), .Y(n_830) );
INVx1_ASAP7_75t_L g976 ( .A(n_509), .Y(n_976) );
AOI222xp33_ASAP7_75t_L g1383 ( .A1(n_509), .A2(n_718), .B1(n_1384), .B2(n_1387), .C1(n_1388), .C2(n_1396), .Y(n_1383) );
OAI22xp5_ASAP7_75t_L g511 ( .A1(n_512), .A2(n_513), .B1(n_516), .B2(n_517), .Y(n_511) );
OAI22xp33_ASAP7_75t_L g541 ( .A1(n_512), .A2(n_525), .B1(n_542), .B2(n_545), .Y(n_541) );
OAI22xp5_ASAP7_75t_L g534 ( .A1(n_513), .A2(n_517), .B1(n_535), .B2(n_536), .Y(n_534) );
INVx2_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
INVx1_ASAP7_75t_L g514 ( .A(n_515), .Y(n_514) );
OAI22xp5_ASAP7_75t_L g824 ( .A1(n_515), .A2(n_825), .B1(n_826), .B2(n_828), .Y(n_824) );
OAI22xp33_ASAP7_75t_L g558 ( .A1(n_516), .A2(n_528), .B1(n_559), .B2(n_563), .Y(n_558) );
OAI22xp5_ASAP7_75t_L g937 ( .A1(n_517), .A2(n_916), .B1(n_934), .B2(n_938), .Y(n_937) );
OAI22xp5_ASAP7_75t_L g943 ( .A1(n_517), .A2(n_926), .B1(n_930), .B2(n_938), .Y(n_943) );
INVx2_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
OAI22xp5_ASAP7_75t_L g519 ( .A1(n_520), .A2(n_521), .B1(n_522), .B2(n_523), .Y(n_519) );
OAI22xp5_ASAP7_75t_L g524 ( .A1(n_520), .A2(n_525), .B1(n_526), .B2(n_528), .Y(n_524) );
OAI22xp5_ASAP7_75t_L g941 ( .A1(n_520), .A2(n_522), .B1(n_923), .B2(n_929), .Y(n_941) );
OAI22xp5_ASAP7_75t_L g942 ( .A1(n_520), .A2(n_522), .B1(n_918), .B2(n_935), .Y(n_942) );
INVx1_ASAP7_75t_L g983 ( .A(n_520), .Y(n_983) );
OAI22xp5_ASAP7_75t_L g548 ( .A1(n_521), .A2(n_535), .B1(n_549), .B2(n_552), .Y(n_548) );
OAI22xp5_ASAP7_75t_L g554 ( .A1(n_523), .A2(n_536), .B1(n_555), .B2(n_557), .Y(n_554) );
OAI22xp5_ASAP7_75t_L g755 ( .A1(n_526), .A2(n_756), .B1(n_758), .B2(n_759), .Y(n_755) );
OAI22xp5_ASAP7_75t_L g981 ( .A1(n_526), .A2(n_964), .B1(n_968), .B2(n_982), .Y(n_981) );
OAI22xp33_ASAP7_75t_L g984 ( .A1(n_526), .A2(n_962), .B1(n_974), .B2(n_985), .Y(n_984) );
OAI22xp5_ASAP7_75t_L g1037 ( .A1(n_526), .A2(n_1023), .B1(n_1033), .B2(n_1038), .Y(n_1037) );
OAI22xp5_ASAP7_75t_L g1082 ( .A1(n_526), .A2(n_705), .B1(n_1064), .B2(n_1077), .Y(n_1082) );
OAI22xp5_ASAP7_75t_L g1110 ( .A1(n_526), .A2(n_705), .B1(n_1111), .B2(n_1112), .Y(n_1110) );
INVx5_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
OAI33xp33_ASAP7_75t_L g936 ( .A1(n_529), .A2(n_830), .A3(n_937), .B1(n_941), .B2(n_942), .B3(n_943), .Y(n_936) );
INVx2_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
INVx1_ASAP7_75t_L g530 ( .A(n_531), .Y(n_530) );
INVx1_ASAP7_75t_L g532 ( .A(n_533), .Y(n_532) );
OAI33xp33_ASAP7_75t_L g537 ( .A1(n_538), .A2(n_541), .A3(n_548), .B1(n_554), .B2(n_558), .B3(n_564), .Y(n_537) );
OAI33xp33_ASAP7_75t_L g959 ( .A1(n_538), .A2(n_564), .A3(n_960), .B1(n_963), .B2(n_967), .B3(n_972), .Y(n_959) );
OAI33xp33_ASAP7_75t_L g1020 ( .A1(n_538), .A2(n_564), .A3(n_1021), .B1(n_1024), .B2(n_1027), .B3(n_1031), .Y(n_1020) );
BUFx4f_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
BUFx4f_ASAP7_75t_L g599 ( .A(n_539), .Y(n_599) );
BUFx8_ASAP7_75t_L g720 ( .A(n_539), .Y(n_720) );
BUFx2_ASAP7_75t_L g887 ( .A(n_540), .Y(n_887) );
INVx2_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
INVx1_ASAP7_75t_L g543 ( .A(n_544), .Y(n_543) );
OAI221xp5_ASAP7_75t_L g1359 ( .A1(n_544), .A2(n_547), .B1(n_881), .B2(n_1360), .C(n_1361), .Y(n_1359) );
OAI22xp5_ASAP7_75t_L g933 ( .A1(n_545), .A2(n_917), .B1(n_934), .B2(n_935), .Y(n_933) );
OAI22xp33_ASAP7_75t_L g1031 ( .A1(n_545), .A2(n_722), .B1(n_1032), .B2(n_1033), .Y(n_1031) );
OAI22xp5_ASAP7_75t_L g1067 ( .A1(n_545), .A2(n_1068), .B1(n_1069), .B2(n_1070), .Y(n_1067) );
OAI22xp33_ASAP7_75t_L g1071 ( .A1(n_545), .A2(n_880), .B1(n_1072), .B2(n_1073), .Y(n_1071) );
INVx2_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
INVx2_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
BUFx6f_ASAP7_75t_L g563 ( .A(n_547), .Y(n_563) );
OAI221xp5_ASAP7_75t_L g1351 ( .A1(n_547), .A2(n_1352), .B1(n_1353), .B2(n_1354), .C(n_1355), .Y(n_1351) );
OAI221xp5_ASAP7_75t_L g590 ( .A1(n_549), .A2(n_591), .B1(n_592), .B2(n_593), .C(n_594), .Y(n_590) );
INVx1_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
INVx1_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
BUFx2_ASAP7_75t_L g601 ( .A(n_551), .Y(n_601) );
INVx3_ASAP7_75t_L g774 ( .A(n_551), .Y(n_774) );
OR2x6_ASAP7_75t_SL g1366 ( .A(n_551), .B(n_1367), .Y(n_1366) );
OAI22xp5_ASAP7_75t_L g922 ( .A1(n_552), .A2(n_923), .B1(n_924), .B2(n_926), .Y(n_922) );
OAI22xp5_ASAP7_75t_L g927 ( .A1(n_552), .A2(n_928), .B1(n_929), .B2(n_930), .Y(n_927) );
INVx3_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
INVx3_ASAP7_75t_L g557 ( .A(n_553), .Y(n_557) );
CKINVDCx8_ASAP7_75t_R g592 ( .A(n_553), .Y(n_592) );
INVx3_ASAP7_75t_L g971 ( .A(n_553), .Y(n_971) );
INVx1_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
OAI221xp5_ASAP7_75t_L g600 ( .A1(n_557), .A2(n_601), .B1(n_602), .B2(n_603), .C(n_604), .Y(n_600) );
OAI22xp5_ASAP7_75t_L g1123 ( .A1(n_557), .A2(n_1111), .B1(n_1117), .B2(n_1124), .Y(n_1123) );
INVx1_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
INVx1_ASAP7_75t_L g917 ( .A(n_560), .Y(n_917) );
INVx2_ASAP7_75t_SL g560 ( .A(n_561), .Y(n_560) );
OR2x2_ASAP7_75t_L g1469 ( .A(n_561), .B(n_1470), .Y(n_1469) );
INVx2_ASAP7_75t_SL g561 ( .A(n_562), .Y(n_561) );
INVx3_ASAP7_75t_L g1069 ( .A(n_562), .Y(n_1069) );
OAI22xp33_ASAP7_75t_L g960 ( .A1(n_563), .A2(n_722), .B1(n_961), .B2(n_962), .Y(n_960) );
OAI22xp33_ASAP7_75t_L g972 ( .A1(n_563), .A2(n_722), .B1(n_973), .B2(n_974), .Y(n_972) );
OAI22xp33_ASAP7_75t_L g1021 ( .A1(n_563), .A2(n_722), .B1(n_1022), .B2(n_1023), .Y(n_1021) );
OAI22xp5_ASAP7_75t_L g589 ( .A1(n_564), .A2(n_590), .B1(n_598), .B2(n_600), .Y(n_589) );
INVx2_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
CKINVDCx5p33_ASAP7_75t_R g1074 ( .A(n_565), .Y(n_1074) );
INVx3_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
INVx3_ASAP7_75t_L g736 ( .A(n_566), .Y(n_736) );
OAI33xp33_ASAP7_75t_L g765 ( .A1(n_566), .A2(n_720), .A3(n_766), .B1(n_772), .B2(n_775), .B3(n_777), .Y(n_765) );
XNOR2xp5_ASAP7_75t_L g568 ( .A(n_569), .B(n_652), .Y(n_568) );
INVx1_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
HB1xp67_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
INVx1_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
INVx2_ASAP7_75t_L g1137 ( .A(n_578), .Y(n_1137) );
AOI211xp5_ASAP7_75t_SL g636 ( .A1(n_582), .A2(n_637), .B(n_639), .C(n_648), .Y(n_636) );
NAND2xp5_ASAP7_75t_L g645 ( .A(n_583), .B(n_646), .Y(n_645) );
INVx1_ASAP7_75t_L g608 ( .A(n_584), .Y(n_608) );
INVx1_ASAP7_75t_L g951 ( .A(n_588), .Y(n_951) );
INVx2_ASAP7_75t_L g1048 ( .A(n_588), .Y(n_1048) );
OAI22xp5_ASAP7_75t_L g772 ( .A1(n_592), .A2(n_752), .B1(n_763), .B2(n_773), .Y(n_772) );
OAI22xp5_ASAP7_75t_L g882 ( .A1(n_592), .A2(n_727), .B1(n_883), .B2(n_884), .Y(n_882) );
OAI22xp5_ASAP7_75t_L g1127 ( .A1(n_592), .A2(n_1112), .B1(n_1119), .B2(n_1128), .Y(n_1127) );
BUFx3_ASAP7_75t_L g595 ( .A(n_596), .Y(n_595) );
INVx1_ASAP7_75t_L g606 ( .A(n_596), .Y(n_606) );
INVx2_ASAP7_75t_SL g1456 ( .A(n_596), .Y(n_1456) );
OAI33xp33_ASAP7_75t_L g914 ( .A1(n_598), .A2(n_915), .A3(n_922), .B1(n_927), .B2(n_931), .B3(n_933), .Y(n_914) );
OAI33xp33_ASAP7_75t_L g1062 ( .A1(n_598), .A2(n_1063), .A3(n_1067), .B1(n_1071), .B2(n_1074), .B3(n_1075), .Y(n_1062) );
BUFx3_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
OAI211xp5_ASAP7_75t_SL g631 ( .A1(n_602), .A2(n_624), .B(n_632), .C(n_635), .Y(n_631) );
INVx1_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
INVx1_ASAP7_75t_L g607 ( .A(n_608), .Y(n_607) );
AOI21xp33_ASAP7_75t_L g609 ( .A1(n_610), .A2(n_636), .B(n_649), .Y(n_609) );
NOR2xp33_ASAP7_75t_L g610 ( .A(n_611), .B(n_619), .Y(n_610) );
INVx1_ASAP7_75t_L g612 ( .A(n_613), .Y(n_612) );
AOI22xp33_ASAP7_75t_L g1430 ( .A1(n_613), .A2(n_1431), .B1(n_1432), .B2(n_1433), .Y(n_1430) );
BUFx6f_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
AND2x4_ASAP7_75t_L g849 ( .A(n_614), .B(n_850), .Y(n_849) );
INVx2_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
AND2x4_ASAP7_75t_L g815 ( .A(n_617), .B(n_816), .Y(n_815) );
INVx3_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
INVx1_ASAP7_75t_L g620 ( .A(n_621), .Y(n_620) );
HB1xp67_ASAP7_75t_L g1433 ( .A(n_621), .Y(n_1433) );
OAI211xp5_ASAP7_75t_L g622 ( .A1(n_623), .A2(n_624), .B(n_625), .C(n_629), .Y(n_622) );
INVx2_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
INVx2_ASAP7_75t_L g633 ( .A(n_627), .Y(n_633) );
INVx2_ASAP7_75t_L g822 ( .A(n_633), .Y(n_822) );
BUFx3_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
INVx2_ASAP7_75t_L g1437 ( .A(n_638), .Y(n_1437) );
INVx1_ASAP7_75t_L g1386 ( .A(n_640), .Y(n_1386) );
BUFx2_ASAP7_75t_L g1438 ( .A(n_641), .Y(n_1438) );
INVx2_ASAP7_75t_L g641 ( .A(n_642), .Y(n_641) );
NOR2x1_ASAP7_75t_L g642 ( .A(n_643), .B(n_644), .Y(n_642) );
INVx1_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
AOI21xp5_ASAP7_75t_SL g1424 ( .A1(n_648), .A2(n_1425), .B(n_1429), .Y(n_1424) );
INVx1_ASAP7_75t_L g1444 ( .A(n_649), .Y(n_1444) );
INVx1_ASAP7_75t_L g649 ( .A(n_650), .Y(n_649) );
OAI22x1_ASAP7_75t_L g652 ( .A1(n_653), .A2(n_805), .B1(n_806), .B2(n_892), .Y(n_652) );
INVx1_ASAP7_75t_L g892 ( .A(n_653), .Y(n_892) );
XNOR2x1_ASAP7_75t_L g653 ( .A(n_654), .B(n_739), .Y(n_653) );
NAND3xp33_ASAP7_75t_L g655 ( .A(n_656), .B(n_673), .C(n_689), .Y(n_655) );
INVx2_ASAP7_75t_SL g658 ( .A(n_659), .Y(n_658) );
HB1xp67_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
OAI211xp5_ASAP7_75t_L g885 ( .A1(n_663), .A2(n_833), .B(n_886), .C(n_888), .Y(n_885) );
INVx2_ASAP7_75t_L g663 ( .A(n_664), .Y(n_663) );
AOI22xp33_ASAP7_75t_L g677 ( .A1(n_667), .A2(n_678), .B1(n_679), .B2(n_681), .Y(n_677) );
INVx1_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
OAI31xp33_ASAP7_75t_L g673 ( .A1(n_674), .A2(n_682), .A3(n_686), .B(n_688), .Y(n_673) );
OAI22xp5_ASAP7_75t_L g699 ( .A1(n_675), .A2(n_700), .B1(n_701), .B2(n_703), .Y(n_699) );
OAI22xp5_ASAP7_75t_L g751 ( .A1(n_675), .A2(n_752), .B1(n_753), .B2(n_754), .Y(n_751) );
INVx1_ASAP7_75t_L g1014 ( .A(n_675), .Y(n_1014) );
OAI22xp5_ASAP7_75t_L g1113 ( .A1(n_675), .A2(n_753), .B1(n_1114), .B2(n_1115), .Y(n_1113) );
AOI22xp33_ASAP7_75t_L g797 ( .A1(n_678), .A2(n_783), .B1(n_798), .B2(n_800), .Y(n_797) );
AOI22xp33_ASAP7_75t_L g1099 ( .A1(n_678), .A2(n_798), .B1(n_1093), .B2(n_1100), .Y(n_1099) );
INVx2_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
INVx1_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
INVx2_ASAP7_75t_L g803 ( .A(n_685), .Y(n_803) );
INVx1_ASAP7_75t_L g912 ( .A(n_685), .Y(n_912) );
OAI31xp33_ASAP7_75t_SL g1005 ( .A1(n_688), .A2(n_1006), .A3(n_1008), .B(n_1012), .Y(n_1005) );
OAI31xp33_ASAP7_75t_L g1051 ( .A1(n_688), .A2(n_1052), .A3(n_1054), .B(n_1055), .Y(n_1051) );
NOR2xp33_ASAP7_75t_L g689 ( .A(n_690), .B(n_719), .Y(n_689) );
OAI33xp33_ASAP7_75t_L g690 ( .A1(n_691), .A2(n_694), .A3(n_699), .B1(n_704), .B2(n_711), .B3(n_717), .Y(n_690) );
OAI33xp33_ASAP7_75t_L g1106 ( .A1(n_691), .A2(n_717), .A3(n_1107), .B1(n_1110), .B2(n_1113), .B3(n_1116), .Y(n_1106) );
INVx1_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
INVx2_ASAP7_75t_SL g692 ( .A(n_693), .Y(n_692) );
OAI22xp33_ASAP7_75t_L g694 ( .A1(n_695), .A2(n_696), .B1(n_697), .B2(n_698), .Y(n_694) );
OAI22xp33_ASAP7_75t_L g721 ( .A1(n_695), .A2(n_708), .B1(n_722), .B2(n_725), .Y(n_721) );
OAI22xp5_ASAP7_75t_L g1086 ( .A1(n_696), .A2(n_980), .B1(n_1066), .B2(n_1078), .Y(n_1086) );
OAI22xp33_ASAP7_75t_L g737 ( .A1(n_697), .A2(n_710), .B1(n_722), .B2(n_738), .Y(n_737) );
OAI22xp5_ASAP7_75t_L g1116 ( .A1(n_698), .A2(n_1117), .B1(n_1118), .B2(n_1119), .Y(n_1116) );
OAI22xp5_ASAP7_75t_L g726 ( .A1(n_700), .A2(n_713), .B1(n_727), .B2(n_729), .Y(n_726) );
INVx3_ASAP7_75t_L g701 ( .A(n_702), .Y(n_701) );
OAI22xp5_ASAP7_75t_L g732 ( .A1(n_703), .A2(n_716), .B1(n_729), .B2(n_733), .Y(n_732) );
OAI22xp5_ASAP7_75t_L g704 ( .A1(n_705), .A2(n_708), .B1(n_709), .B2(n_710), .Y(n_704) );
INVx4_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
INVx2_ASAP7_75t_L g753 ( .A(n_706), .Y(n_753) );
INVx2_ASAP7_75t_L g1038 ( .A(n_706), .Y(n_1038) );
INVx2_ASAP7_75t_L g1084 ( .A(n_706), .Y(n_1084) );
INVx4_ASAP7_75t_L g706 ( .A(n_707), .Y(n_706) );
OAI221xp5_ASAP7_75t_L g832 ( .A1(n_709), .A2(n_756), .B1(n_833), .B2(n_834), .C(n_835), .Y(n_832) );
OAI22xp5_ASAP7_75t_L g711 ( .A1(n_712), .A2(n_713), .B1(n_714), .B2(n_716), .Y(n_711) );
OAI22xp33_ASAP7_75t_L g1080 ( .A1(n_712), .A2(n_1068), .B1(n_1072), .B2(n_1081), .Y(n_1080) );
OAI22xp33_ASAP7_75t_L g1107 ( .A1(n_712), .A2(n_826), .B1(n_1108), .B2(n_1109), .Y(n_1107) );
OAI22xp5_ASAP7_75t_L g760 ( .A1(n_714), .A2(n_761), .B1(n_763), .B2(n_764), .Y(n_760) );
OAI22xp33_ASAP7_75t_L g1039 ( .A1(n_714), .A2(n_988), .B1(n_1026), .B2(n_1030), .Y(n_1039) );
INVx5_ASAP7_75t_L g714 ( .A(n_715), .Y(n_714) );
INVx6_ASAP7_75t_L g980 ( .A(n_715), .Y(n_980) );
OAI33xp33_ASAP7_75t_L g742 ( .A1(n_717), .A2(n_743), .A3(n_745), .B1(n_751), .B2(n_755), .B3(n_760), .Y(n_742) );
OAI21xp5_ASAP7_75t_L g831 ( .A1(n_717), .A2(n_832), .B(n_838), .Y(n_831) );
CKINVDCx5p33_ASAP7_75t_R g717 ( .A(n_718), .Y(n_717) );
INVx2_ASAP7_75t_L g986 ( .A(n_718), .Y(n_986) );
OAI33xp33_ASAP7_75t_L g719 ( .A1(n_720), .A2(n_721), .A3(n_726), .B1(n_732), .B2(n_734), .B3(n_737), .Y(n_719) );
INVx2_ASAP7_75t_L g722 ( .A(n_723), .Y(n_722) );
INVx1_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
INVx1_ASAP7_75t_L g768 ( .A(n_724), .Y(n_768) );
INVx2_ASAP7_75t_L g727 ( .A(n_728), .Y(n_727) );
OAI22xp5_ASAP7_75t_L g775 ( .A1(n_729), .A2(n_754), .B1(n_764), .B2(n_776), .Y(n_775) );
OAI22xp33_ASAP7_75t_SL g1063 ( .A1(n_729), .A2(n_1064), .B1(n_1065), .B2(n_1066), .Y(n_1063) );
INVx3_ASAP7_75t_L g729 ( .A(n_730), .Y(n_729) );
BUFx2_ASAP7_75t_L g730 ( .A(n_731), .Y(n_730) );
INVx8_ASAP7_75t_L g925 ( .A(n_733), .Y(n_925) );
BUFx3_ASAP7_75t_L g1076 ( .A(n_733), .Y(n_1076) );
INVx1_ASAP7_75t_L g734 ( .A(n_735), .Y(n_734) );
BUFx2_ASAP7_75t_L g735 ( .A(n_736), .Y(n_735) );
BUFx2_ASAP7_75t_L g932 ( .A(n_736), .Y(n_932) );
NAND3xp33_ASAP7_75t_L g740 ( .A(n_741), .B(n_778), .C(n_789), .Y(n_740) );
NOR2xp33_ASAP7_75t_L g741 ( .A(n_742), .B(n_765), .Y(n_741) );
BUFx6f_ASAP7_75t_L g743 ( .A(n_744), .Y(n_743) );
OAI22xp33_ASAP7_75t_L g745 ( .A1(n_746), .A2(n_747), .B1(n_749), .B2(n_750), .Y(n_745) );
OAI22xp33_ASAP7_75t_L g766 ( .A1(n_746), .A2(n_758), .B1(n_767), .B2(n_769), .Y(n_766) );
INVx1_ASAP7_75t_L g747 ( .A(n_748), .Y(n_747) );
OAI22xp5_ASAP7_75t_L g1397 ( .A1(n_750), .A2(n_990), .B1(n_1398), .B2(n_1399), .Y(n_1397) );
INVx2_ASAP7_75t_L g756 ( .A(n_757), .Y(n_756) );
OAI221xp5_ASAP7_75t_L g1439 ( .A1(n_761), .A2(n_1440), .B1(n_1441), .B2(n_1442), .C(n_1443), .Y(n_1439) );
INVx2_ASAP7_75t_L g761 ( .A(n_762), .Y(n_761) );
INVx2_ASAP7_75t_L g767 ( .A(n_768), .Y(n_767) );
INVx1_ASAP7_75t_L g769 ( .A(n_770), .Y(n_769) );
INVxp67_ASAP7_75t_SL g1043 ( .A(n_770), .Y(n_1043) );
INVx1_ASAP7_75t_L g770 ( .A(n_771), .Y(n_770) );
INVx1_ASAP7_75t_L g999 ( .A(n_771), .Y(n_999) );
OR2x6_ASAP7_75t_L g1371 ( .A(n_771), .B(n_865), .Y(n_1371) );
INVx2_ASAP7_75t_L g773 ( .A(n_774), .Y(n_773) );
OAI31xp33_ASAP7_75t_L g778 ( .A1(n_779), .A2(n_780), .A3(n_785), .B(n_788), .Y(n_778) );
INVx1_ASAP7_75t_L g786 ( .A(n_787), .Y(n_786) );
OAI31xp33_ASAP7_75t_L g994 ( .A1(n_788), .A2(n_995), .A3(n_997), .B(n_1003), .Y(n_994) );
OAI31xp33_ASAP7_75t_L g1087 ( .A1(n_788), .A2(n_1088), .A3(n_1091), .B(n_1095), .Y(n_1087) );
OAI31xp33_ASAP7_75t_L g789 ( .A1(n_790), .A2(n_791), .A3(n_801), .B(n_804), .Y(n_789) );
INVx2_ASAP7_75t_L g793 ( .A(n_794), .Y(n_793) );
INVx1_ASAP7_75t_L g795 ( .A(n_796), .Y(n_795) );
INVx2_ASAP7_75t_L g798 ( .A(n_799), .Y(n_798) );
OAI31xp33_ASAP7_75t_L g1096 ( .A1(n_804), .A2(n_1097), .A3(n_1098), .B(n_1101), .Y(n_1096) );
INVx1_ASAP7_75t_L g805 ( .A(n_806), .Y(n_805) );
INVx1_ASAP7_75t_L g806 ( .A(n_807), .Y(n_806) );
XNOR2x1_ASAP7_75t_L g807 ( .A(n_808), .B(n_809), .Y(n_807) );
NAND4xp75_ASAP7_75t_L g809 ( .A(n_810), .B(n_819), .C(n_847), .D(n_854), .Y(n_809) );
INVx1_ASAP7_75t_L g811 ( .A(n_812), .Y(n_811) );
INVx1_ASAP7_75t_L g812 ( .A(n_813), .Y(n_812) );
INVx1_ASAP7_75t_L g814 ( .A(n_815), .Y(n_814) );
AOI222xp33_ASAP7_75t_L g1378 ( .A1(n_815), .A2(n_1363), .B1(n_1379), .B2(n_1380), .C1(n_1381), .C2(n_1382), .Y(n_1378) );
INVx1_ASAP7_75t_L g816 ( .A(n_817), .Y(n_816) );
AOI211x1_ASAP7_75t_L g819 ( .A1(n_820), .A2(n_829), .B(n_831), .C(n_842), .Y(n_819) );
INVx2_ASAP7_75t_L g821 ( .A(n_822), .Y(n_821) );
INVx2_ASAP7_75t_L g1427 ( .A(n_822), .Y(n_1427) );
BUFx6f_ASAP7_75t_L g826 ( .A(n_827), .Y(n_826) );
OAI221xp5_ASAP7_75t_L g878 ( .A1(n_828), .A2(n_834), .B1(n_879), .B2(n_880), .C(n_881), .Y(n_878) );
INVx1_ASAP7_75t_L g829 ( .A(n_830), .Y(n_829) );
OAI33xp33_ASAP7_75t_L g1079 ( .A1(n_830), .A2(n_986), .A3(n_1080), .B1(n_1082), .B2(n_1083), .B3(n_1086), .Y(n_1079) );
INVx2_ASAP7_75t_L g836 ( .A(n_837), .Y(n_836) );
CKINVDCx5p33_ASAP7_75t_R g1406 ( .A(n_838), .Y(n_1406) );
INVx1_ASAP7_75t_L g839 ( .A(n_840), .Y(n_839) );
NAND2x2_ASAP7_75t_L g843 ( .A(n_840), .B(n_844), .Y(n_843) );
INVx2_ASAP7_75t_L g840 ( .A(n_841), .Y(n_840) );
INVx1_ASAP7_75t_L g1379 ( .A(n_843), .Y(n_1379) );
INVx2_ASAP7_75t_SL g844 ( .A(n_845), .Y(n_844) );
INVx2_ASAP7_75t_SL g1381 ( .A(n_846), .Y(n_1381) );
AOI22xp5_ASAP7_75t_L g847 ( .A1(n_848), .A2(n_849), .B1(n_851), .B2(n_852), .Y(n_847) );
AOI22xp33_ASAP7_75t_L g867 ( .A1(n_848), .A2(n_851), .B1(n_868), .B2(n_869), .Y(n_867) );
NAND2xp5_ASAP7_75t_L g1400 ( .A(n_849), .B(n_1401), .Y(n_1400) );
AND2x4_ASAP7_75t_L g852 ( .A(n_850), .B(n_853), .Y(n_852) );
INVx1_ASAP7_75t_L g1376 ( .A(n_852), .Y(n_1376) );
OAI31xp67_ASAP7_75t_L g854 ( .A1(n_855), .A2(n_866), .A3(n_877), .B(n_890), .Y(n_854) );
INVx4_ASAP7_75t_L g856 ( .A(n_857), .Y(n_856) );
INVx2_ASAP7_75t_L g858 ( .A(n_859), .Y(n_858) );
A2O1A1Ixp33_ASAP7_75t_L g860 ( .A1(n_861), .A2(n_862), .B(n_863), .C(n_864), .Y(n_860) );
INVx1_ASAP7_75t_L g864 ( .A(n_865), .Y(n_864) );
AOI21xp33_ASAP7_75t_L g866 ( .A1(n_867), .A2(n_871), .B(n_874), .Y(n_866) );
INVx2_ASAP7_75t_L g969 ( .A(n_869), .Y(n_969) );
INVx2_ASAP7_75t_L g869 ( .A(n_870), .Y(n_869) );
INVx1_ASAP7_75t_L g874 ( .A(n_875), .Y(n_874) );
HB1xp67_ASAP7_75t_L g875 ( .A(n_876), .Y(n_875) );
INVx2_ASAP7_75t_L g1367 ( .A(n_876), .Y(n_1367) );
OAI21xp5_ASAP7_75t_SL g877 ( .A1(n_878), .A2(n_882), .B(n_885), .Y(n_877) );
INVx2_ASAP7_75t_L g1372 ( .A(n_890), .Y(n_1372) );
BUFx2_ASAP7_75t_L g890 ( .A(n_891), .Y(n_890) );
HB1xp67_ASAP7_75t_L g893 ( .A(n_894), .Y(n_893) );
AOI22xp5_ASAP7_75t_L g894 ( .A1(n_895), .A2(n_896), .B1(n_954), .B2(n_1150), .Y(n_894) );
INVx1_ASAP7_75t_L g895 ( .A(n_896), .Y(n_895) );
HB1xp67_ASAP7_75t_L g896 ( .A(n_897), .Y(n_896) );
INVx1_ASAP7_75t_L g897 ( .A(n_898), .Y(n_897) );
INVx1_ASAP7_75t_L g899 ( .A(n_900), .Y(n_899) );
NAND3xp33_ASAP7_75t_L g900 ( .A(n_901), .B(n_913), .C(n_944), .Y(n_900) );
NOR2xp33_ASAP7_75t_SL g913 ( .A(n_914), .B(n_936), .Y(n_913) );
OAI22xp5_ASAP7_75t_L g915 ( .A1(n_916), .A2(n_917), .B1(n_918), .B2(n_919), .Y(n_915) );
INVx2_ASAP7_75t_SL g919 ( .A(n_920), .Y(n_919) );
INVx1_ASAP7_75t_L g920 ( .A(n_921), .Y(n_920) );
OAI22xp5_ASAP7_75t_L g963 ( .A1(n_924), .A2(n_964), .B1(n_965), .B2(n_966), .Y(n_963) );
OAI22xp5_ASAP7_75t_L g1024 ( .A1(n_924), .A2(n_966), .B1(n_1025), .B2(n_1026), .Y(n_1024) );
INVx2_ASAP7_75t_L g924 ( .A(n_925), .Y(n_924) );
INVx1_ASAP7_75t_L g1065 ( .A(n_925), .Y(n_1065) );
INVx1_ASAP7_75t_L g931 ( .A(n_932), .Y(n_931) );
INVx2_ASAP7_75t_L g938 ( .A(n_939), .Y(n_938) );
INVx2_ASAP7_75t_SL g939 ( .A(n_940), .Y(n_939) );
OAI31xp33_ASAP7_75t_L g944 ( .A1(n_945), .A2(n_947), .A3(n_950), .B(n_952), .Y(n_944) );
INVx1_ASAP7_75t_L g1150 ( .A(n_954), .Y(n_1150) );
XNOR2xp5_ASAP7_75t_L g954 ( .A(n_955), .B(n_1058), .Y(n_954) );
XOR2xp5_ASAP7_75t_L g955 ( .A(n_956), .B(n_1017), .Y(n_955) );
AND3x1_ASAP7_75t_L g957 ( .A(n_958), .B(n_994), .C(n_1005), .Y(n_957) );
NOR2xp33_ASAP7_75t_L g958 ( .A(n_959), .B(n_975), .Y(n_958) );
OAI22xp33_ASAP7_75t_L g977 ( .A1(n_961), .A2(n_973), .B1(n_978), .B2(n_980), .Y(n_977) );
OAI22xp5_ASAP7_75t_L g987 ( .A1(n_965), .A2(n_970), .B1(n_988), .B2(n_992), .Y(n_987) );
OAI22xp5_ASAP7_75t_L g1075 ( .A1(n_966), .A2(n_1076), .B1(n_1077), .B2(n_1078), .Y(n_1075) );
OAI22xp5_ASAP7_75t_L g967 ( .A1(n_968), .A2(n_969), .B1(n_970), .B2(n_971), .Y(n_967) );
OAI22xp5_ASAP7_75t_L g1027 ( .A1(n_971), .A2(n_1028), .B1(n_1029), .B2(n_1030), .Y(n_1027) );
OAI33xp33_ASAP7_75t_L g975 ( .A1(n_976), .A2(n_977), .A3(n_981), .B1(n_984), .B2(n_986), .B3(n_987), .Y(n_975) );
OAI33xp33_ASAP7_75t_L g1034 ( .A1(n_976), .A2(n_986), .A3(n_1035), .B1(n_1036), .B2(n_1037), .B3(n_1039), .Y(n_1034) );
OAI22xp33_ASAP7_75t_L g1035 ( .A1(n_978), .A2(n_980), .B1(n_1022), .B2(n_1032), .Y(n_1035) );
INVx2_ASAP7_75t_L g978 ( .A(n_979), .Y(n_978) );
INVx3_ASAP7_75t_L g1118 ( .A(n_979), .Y(n_1118) );
INVx1_ASAP7_75t_L g982 ( .A(n_983), .Y(n_982) );
INVx1_ASAP7_75t_L g988 ( .A(n_989), .Y(n_988) );
INVx1_ASAP7_75t_L g989 ( .A(n_990), .Y(n_989) );
INVx1_ASAP7_75t_L g990 ( .A(n_991), .Y(n_990) );
BUFx3_ASAP7_75t_L g992 ( .A(n_993), .Y(n_992) );
INVxp67_ASAP7_75t_L g998 ( .A(n_999), .Y(n_998) );
INVx1_ASAP7_75t_L g1126 ( .A(n_999), .Y(n_1126) );
INVx1_ASAP7_75t_L g1009 ( .A(n_1010), .Y(n_1009) );
INVx2_ASAP7_75t_SL g1010 ( .A(n_1011), .Y(n_1010) );
INVx1_ASAP7_75t_L g1013 ( .A(n_1014), .Y(n_1013) );
AND3x1_ASAP7_75t_L g1018 ( .A(n_1019), .B(n_1040), .C(n_1051), .Y(n_1018) );
NOR2xp33_ASAP7_75t_L g1019 ( .A(n_1020), .B(n_1034), .Y(n_1019) );
HB1xp67_ASAP7_75t_L g1042 ( .A(n_1043), .Y(n_1042) );
OA22x2_ASAP7_75t_L g1058 ( .A1(n_1059), .A2(n_1102), .B1(n_1103), .B2(n_1149), .Y(n_1058) );
INVx1_ASAP7_75t_L g1149 ( .A(n_1059), .Y(n_1149) );
NAND3xp33_ASAP7_75t_L g1060 ( .A(n_1061), .B(n_1087), .C(n_1096), .Y(n_1060) );
NOR2xp33_ASAP7_75t_L g1061 ( .A(n_1062), .B(n_1079), .Y(n_1061) );
OAI22xp33_ASAP7_75t_L g1121 ( .A1(n_1069), .A2(n_1108), .B1(n_1114), .B2(n_1122), .Y(n_1121) );
OAI22xp33_ASAP7_75t_L g1125 ( .A1(n_1069), .A2(n_1109), .B1(n_1115), .B2(n_1126), .Y(n_1125) );
OAI22xp5_ASAP7_75t_L g1083 ( .A1(n_1070), .A2(n_1073), .B1(n_1084), .B2(n_1085), .Y(n_1083) );
INVx1_ASAP7_75t_L g1089 ( .A(n_1090), .Y(n_1089) );
INVx2_ASAP7_75t_SL g1102 ( .A(n_1103), .Y(n_1102) );
NAND3xp33_ASAP7_75t_L g1104 ( .A(n_1105), .B(n_1129), .C(n_1139), .Y(n_1104) );
NOR2xp33_ASAP7_75t_L g1105 ( .A(n_1106), .B(n_1120), .Y(n_1105) );
OAI31xp33_ASAP7_75t_L g1129 ( .A1(n_1130), .A2(n_1132), .A3(n_1136), .B(n_1138), .Y(n_1129) );
OAI31xp33_ASAP7_75t_SL g1139 ( .A1(n_1140), .A2(n_1144), .A3(n_1147), .B(n_1148), .Y(n_1139) );
INVx1_ASAP7_75t_L g1141 ( .A(n_1142), .Y(n_1141) );
INVx1_ASAP7_75t_L g1142 ( .A(n_1143), .Y(n_1142) );
OAI221xp5_ASAP7_75t_L g1151 ( .A1(n_1152), .A2(n_1335), .B1(n_1338), .B2(n_1407), .C(n_1412), .Y(n_1151) );
AOI221xp5_ASAP7_75t_SL g1152 ( .A1(n_1153), .A2(n_1216), .B1(n_1273), .B2(n_1275), .C(n_1302), .Y(n_1152) );
A2O1A1Ixp33_ASAP7_75t_L g1153 ( .A1(n_1154), .A2(n_1190), .B(n_1201), .C(n_1210), .Y(n_1153) );
NAND2xp5_ASAP7_75t_L g1154 ( .A(n_1155), .B(n_1185), .Y(n_1154) );
INVx1_ASAP7_75t_L g1155 ( .A(n_1156), .Y(n_1155) );
NAND2xp5_ASAP7_75t_L g1156 ( .A(n_1157), .B(n_1175), .Y(n_1156) );
NAND2xp5_ASAP7_75t_L g1227 ( .A(n_1157), .B(n_1182), .Y(n_1227) );
INVx1_ASAP7_75t_L g1266 ( .A(n_1157), .Y(n_1266) );
AND2x2_ASAP7_75t_L g1296 ( .A(n_1157), .B(n_1297), .Y(n_1296) );
AND2x2_ASAP7_75t_L g1157 ( .A(n_1158), .B(n_1172), .Y(n_1157) );
INVx2_ASAP7_75t_L g1197 ( .A(n_1158), .Y(n_1197) );
AND2x2_ASAP7_75t_L g1199 ( .A(n_1158), .B(n_1200), .Y(n_1199) );
NAND2xp5_ASAP7_75t_L g1224 ( .A(n_1158), .B(n_1195), .Y(n_1224) );
OR2x2_ASAP7_75t_L g1158 ( .A(n_1159), .B(n_1166), .Y(n_1158) );
INVx2_ASAP7_75t_L g1213 ( .A(n_1160), .Y(n_1213) );
AND2x6_ASAP7_75t_L g1160 ( .A(n_1161), .B(n_1162), .Y(n_1160) );
AND2x2_ASAP7_75t_L g1164 ( .A(n_1161), .B(n_1165), .Y(n_1164) );
AND2x4_ASAP7_75t_L g1167 ( .A(n_1161), .B(n_1168), .Y(n_1167) );
AND2x6_ASAP7_75t_L g1170 ( .A(n_1161), .B(n_1171), .Y(n_1170) );
AND2x2_ASAP7_75t_L g1180 ( .A(n_1161), .B(n_1165), .Y(n_1180) );
AND2x2_ASAP7_75t_L g1205 ( .A(n_1161), .B(n_1165), .Y(n_1205) );
AND2x2_ASAP7_75t_L g1168 ( .A(n_1163), .B(n_1169), .Y(n_1168) );
INVxp67_ASAP7_75t_L g1215 ( .A(n_1164), .Y(n_1215) );
INVx2_ASAP7_75t_L g1337 ( .A(n_1170), .Y(n_1337) );
HB1xp67_ASAP7_75t_L g1477 ( .A(n_1171), .Y(n_1477) );
AND2x2_ASAP7_75t_L g1196 ( .A(n_1172), .B(n_1197), .Y(n_1196) );
INVx1_ASAP7_75t_L g1200 ( .A(n_1172), .Y(n_1200) );
AND3x1_ASAP7_75t_L g1245 ( .A(n_1172), .B(n_1176), .C(n_1197), .Y(n_1245) );
AND2x2_ASAP7_75t_L g1247 ( .A(n_1172), .B(n_1195), .Y(n_1247) );
NAND2xp5_ASAP7_75t_L g1254 ( .A(n_1172), .B(n_1176), .Y(n_1254) );
OAI32xp33_ASAP7_75t_L g1331 ( .A1(n_1172), .A2(n_1246), .A3(n_1256), .B1(n_1332), .B2(n_1334), .Y(n_1331) );
AND2x2_ASAP7_75t_L g1172 ( .A(n_1173), .B(n_1174), .Y(n_1172) );
AND2x2_ASAP7_75t_L g1291 ( .A(n_1175), .B(n_1261), .Y(n_1291) );
AND2x2_ASAP7_75t_L g1300 ( .A(n_1175), .B(n_1196), .Y(n_1300) );
AND2x2_ASAP7_75t_L g1175 ( .A(n_1176), .B(n_1181), .Y(n_1175) );
AND2x2_ASAP7_75t_L g1220 ( .A(n_1176), .B(n_1199), .Y(n_1220) );
OR2x2_ASAP7_75t_L g1314 ( .A(n_1176), .B(n_1268), .Y(n_1314) );
INVx2_ASAP7_75t_L g1176 ( .A(n_1177), .Y(n_1176) );
BUFx2_ASAP7_75t_L g1195 ( .A(n_1177), .Y(n_1195) );
AND2x2_ASAP7_75t_L g1198 ( .A(n_1177), .B(n_1199), .Y(n_1198) );
OR2x2_ASAP7_75t_L g1226 ( .A(n_1177), .B(n_1227), .Y(n_1226) );
OR2x2_ASAP7_75t_L g1265 ( .A(n_1177), .B(n_1266), .Y(n_1265) );
AND2x2_ASAP7_75t_L g1295 ( .A(n_1177), .B(n_1261), .Y(n_1295) );
AND2x2_ASAP7_75t_L g1177 ( .A(n_1178), .B(n_1179), .Y(n_1177) );
NOR2xp33_ASAP7_75t_L g1223 ( .A(n_1181), .B(n_1224), .Y(n_1223) );
INVx1_ASAP7_75t_L g1240 ( .A(n_1181), .Y(n_1240) );
NAND2xp5_ASAP7_75t_L g1246 ( .A(n_1181), .B(n_1247), .Y(n_1246) );
NOR2xp33_ASAP7_75t_L g1249 ( .A(n_1181), .B(n_1250), .Y(n_1249) );
AND2x2_ASAP7_75t_L g1301 ( .A(n_1181), .B(n_1242), .Y(n_1301) );
INVx2_ASAP7_75t_L g1181 ( .A(n_1182), .Y(n_1181) );
INVx1_ASAP7_75t_L g1193 ( .A(n_1182), .Y(n_1193) );
OR2x2_ASAP7_75t_L g1252 ( .A(n_1182), .B(n_1187), .Y(n_1252) );
AND2x2_ASAP7_75t_L g1260 ( .A(n_1182), .B(n_1261), .Y(n_1260) );
NAND2xp5_ASAP7_75t_L g1280 ( .A(n_1182), .B(n_1207), .Y(n_1280) );
AND2x2_ASAP7_75t_L g1282 ( .A(n_1182), .B(n_1187), .Y(n_1282) );
OR2x2_ASAP7_75t_L g1288 ( .A(n_1182), .B(n_1224), .Y(n_1288) );
AND2x2_ASAP7_75t_L g1297 ( .A(n_1182), .B(n_1195), .Y(n_1297) );
AND2x2_ASAP7_75t_L g1326 ( .A(n_1182), .B(n_1253), .Y(n_1326) );
AND2x2_ASAP7_75t_L g1333 ( .A(n_1182), .B(n_1203), .Y(n_1333) );
AND2x2_ASAP7_75t_L g1182 ( .A(n_1183), .B(n_1184), .Y(n_1182) );
INVx2_ASAP7_75t_L g1218 ( .A(n_1185), .Y(n_1218) );
A2O1A1Ixp33_ASAP7_75t_L g1221 ( .A1(n_1185), .A2(n_1222), .B(n_1223), .C(n_1225), .Y(n_1221) );
AND2x2_ASAP7_75t_L g1269 ( .A(n_1185), .B(n_1236), .Y(n_1269) );
OR2x2_ASAP7_75t_L g1318 ( .A(n_1185), .B(n_1319), .Y(n_1318) );
INVx2_ASAP7_75t_L g1185 ( .A(n_1186), .Y(n_1185) );
AND2x2_ASAP7_75t_L g1232 ( .A(n_1186), .B(n_1207), .Y(n_1232) );
AND2x2_ASAP7_75t_L g1309 ( .A(n_1186), .B(n_1236), .Y(n_1309) );
INVx1_ASAP7_75t_L g1186 ( .A(n_1187), .Y(n_1186) );
OR2x2_ASAP7_75t_L g1237 ( .A(n_1187), .B(n_1207), .Y(n_1237) );
AND2x2_ASAP7_75t_L g1242 ( .A(n_1187), .B(n_1243), .Y(n_1242) );
AND2x2_ASAP7_75t_L g1307 ( .A(n_1187), .B(n_1207), .Y(n_1307) );
AND2x2_ASAP7_75t_L g1187 ( .A(n_1188), .B(n_1189), .Y(n_1187) );
OAI22xp5_ASAP7_75t_L g1190 ( .A1(n_1191), .A2(n_1192), .B1(n_1194), .B2(n_1198), .Y(n_1190) );
INVx1_ASAP7_75t_L g1191 ( .A(n_1192), .Y(n_1191) );
AND2x2_ASAP7_75t_L g1219 ( .A(n_1192), .B(n_1220), .Y(n_1219) );
INVx2_ASAP7_75t_L g1192 ( .A(n_1193), .Y(n_1192) );
NAND2xp5_ASAP7_75t_L g1268 ( .A(n_1193), .B(n_1261), .Y(n_1268) );
O2A1O1Ixp33_ASAP7_75t_SL g1270 ( .A1(n_1193), .A2(n_1197), .B(n_1271), .C(n_1272), .Y(n_1270) );
AND2x2_ASAP7_75t_L g1304 ( .A(n_1193), .B(n_1194), .Y(n_1304) );
INVx1_ASAP7_75t_L g1311 ( .A(n_1194), .Y(n_1311) );
AND2x2_ASAP7_75t_L g1194 ( .A(n_1195), .B(n_1196), .Y(n_1194) );
AOI221xp5_ASAP7_75t_L g1228 ( .A1(n_1195), .A2(n_1229), .B1(n_1233), .B2(n_1235), .C(n_1238), .Y(n_1228) );
OR2x2_ASAP7_75t_L g1234 ( .A(n_1195), .B(n_1197), .Y(n_1234) );
INVx1_ASAP7_75t_L g1250 ( .A(n_1196), .Y(n_1250) );
OR2x2_ASAP7_75t_L g1278 ( .A(n_1196), .B(n_1199), .Y(n_1278) );
OAI332xp33_ASAP7_75t_L g1238 ( .A1(n_1197), .A2(n_1203), .A3(n_1207), .B1(n_1239), .B2(n_1241), .B3(n_1242), .C1(n_1244), .C2(n_1246), .Y(n_1238) );
AND2x2_ASAP7_75t_L g1261 ( .A(n_1197), .B(n_1200), .Y(n_1261) );
O2A1O1Ixp33_ASAP7_75t_L g1283 ( .A1(n_1198), .A2(n_1284), .B(n_1286), .C(n_1287), .Y(n_1283) );
AOI22xp5_ASAP7_75t_L g1276 ( .A1(n_1200), .A2(n_1277), .B1(n_1279), .B2(n_1281), .Y(n_1276) );
INVx1_ASAP7_75t_L g1201 ( .A(n_1202), .Y(n_1201) );
AND2x2_ASAP7_75t_L g1202 ( .A(n_1203), .B(n_1207), .Y(n_1202) );
OR2x2_ASAP7_75t_L g1230 ( .A(n_1203), .B(n_1231), .Y(n_1230) );
CKINVDCx6p67_ASAP7_75t_R g1236 ( .A(n_1203), .Y(n_1236) );
CKINVDCx5p33_ASAP7_75t_R g1241 ( .A(n_1203), .Y(n_1241) );
OR2x2_ASAP7_75t_L g1289 ( .A(n_1203), .B(n_1207), .Y(n_1289) );
OR2x6_ASAP7_75t_L g1203 ( .A(n_1204), .B(n_1206), .Y(n_1203) );
OR2x2_ASAP7_75t_L g1222 ( .A(n_1204), .B(n_1206), .Y(n_1222) );
INVx1_ASAP7_75t_L g1243 ( .A(n_1207), .Y(n_1243) );
OR2x2_ASAP7_75t_L g1256 ( .A(n_1207), .B(n_1236), .Y(n_1256) );
AND2x2_ASAP7_75t_L g1281 ( .A(n_1207), .B(n_1282), .Y(n_1281) );
AND2x2_ASAP7_75t_L g1315 ( .A(n_1207), .B(n_1236), .Y(n_1315) );
AND2x4_ASAP7_75t_L g1207 ( .A(n_1208), .B(n_1209), .Y(n_1207) );
INVx2_ASAP7_75t_SL g1262 ( .A(n_1210), .Y(n_1262) );
INVx2_ASAP7_75t_SL g1274 ( .A(n_1210), .Y(n_1274) );
OAI22xp5_ASAP7_75t_SL g1211 ( .A1(n_1212), .A2(n_1213), .B1(n_1214), .B2(n_1215), .Y(n_1211) );
NAND5xp2_ASAP7_75t_SL g1216 ( .A(n_1217), .B(n_1221), .C(n_1228), .D(n_1248), .E(n_1263), .Y(n_1216) );
NAND2xp5_ASAP7_75t_L g1217 ( .A(n_1218), .B(n_1219), .Y(n_1217) );
NAND2xp5_ASAP7_75t_L g1290 ( .A(n_1218), .B(n_1291), .Y(n_1290) );
INVx1_ASAP7_75t_L g1271 ( .A(n_1220), .Y(n_1271) );
OAI211xp5_ASAP7_75t_SL g1275 ( .A1(n_1222), .A2(n_1276), .B(n_1283), .C(n_1292), .Y(n_1275) );
INVx1_ASAP7_75t_L g1334 ( .A(n_1224), .Y(n_1334) );
OAI21xp5_ASAP7_75t_L g1316 ( .A1(n_1225), .A2(n_1241), .B(n_1317), .Y(n_1316) );
INVx1_ASAP7_75t_L g1225 ( .A(n_1226), .Y(n_1225) );
INVx1_ASAP7_75t_L g1229 ( .A(n_1230), .Y(n_1229) );
NOR2xp33_ASAP7_75t_L g1328 ( .A(n_1230), .B(n_1265), .Y(n_1328) );
CKINVDCx6p67_ASAP7_75t_R g1231 ( .A(n_1232), .Y(n_1231) );
NAND2xp5_ASAP7_75t_L g1239 ( .A(n_1232), .B(n_1240), .Y(n_1239) );
AOI221xp5_ASAP7_75t_L g1248 ( .A1(n_1232), .A2(n_1249), .B1(n_1251), .B2(n_1253), .C(n_1255), .Y(n_1248) );
OAI22xp5_ASAP7_75t_L g1292 ( .A1(n_1232), .A2(n_1293), .B1(n_1298), .B2(n_1301), .Y(n_1292) );
O2A1O1Ixp33_ASAP7_75t_L g1329 ( .A1(n_1232), .A2(n_1291), .B(n_1330), .C(n_1331), .Y(n_1329) );
A2O1A1Ixp33_ASAP7_75t_L g1312 ( .A1(n_1233), .A2(n_1240), .B(n_1313), .C(n_1315), .Y(n_1312) );
INVx1_ASAP7_75t_L g1233 ( .A(n_1234), .Y(n_1233) );
AOI221xp5_ASAP7_75t_L g1303 ( .A1(n_1235), .A2(n_1247), .B1(n_1304), .B2(n_1305), .C(n_1310), .Y(n_1303) );
NOR2xp33_ASAP7_75t_L g1235 ( .A(n_1236), .B(n_1237), .Y(n_1235) );
NOR2xp33_ASAP7_75t_L g1251 ( .A(n_1236), .B(n_1252), .Y(n_1251) );
NAND2xp5_ASAP7_75t_L g1285 ( .A(n_1236), .B(n_1259), .Y(n_1285) );
AND2x2_ASAP7_75t_L g1327 ( .A(n_1236), .B(n_1242), .Y(n_1327) );
INVx2_ASAP7_75t_L g1259 ( .A(n_1237), .Y(n_1259) );
AOI21xp33_ASAP7_75t_L g1310 ( .A1(n_1237), .A2(n_1288), .B(n_1311), .Y(n_1310) );
INVx1_ASAP7_75t_L g1272 ( .A(n_1242), .Y(n_1272) );
NAND2xp5_ASAP7_75t_L g1332 ( .A(n_1242), .B(n_1333), .Y(n_1332) );
A2O1A1Ixp33_ASAP7_75t_L g1287 ( .A1(n_1244), .A2(n_1288), .B(n_1289), .C(n_1290), .Y(n_1287) );
INVx2_ASAP7_75t_L g1244 ( .A(n_1245), .Y(n_1244) );
INVx1_ASAP7_75t_L g1257 ( .A(n_1247), .Y(n_1257) );
INVx1_ASAP7_75t_L g1286 ( .A(n_1252), .Y(n_1286) );
INVx1_ASAP7_75t_L g1253 ( .A(n_1254), .Y(n_1253) );
OAI211xp5_ASAP7_75t_SL g1255 ( .A1(n_1256), .A2(n_1257), .B(n_1258), .C(n_1262), .Y(n_1255) );
NAND2xp5_ASAP7_75t_L g1258 ( .A(n_1259), .B(n_1260), .Y(n_1258) );
INVx1_ASAP7_75t_L g1321 ( .A(n_1261), .Y(n_1321) );
O2A1O1Ixp33_ASAP7_75t_L g1263 ( .A1(n_1264), .A2(n_1267), .B(n_1269), .C(n_1270), .Y(n_1263) );
INVx1_ASAP7_75t_L g1264 ( .A(n_1265), .Y(n_1264) );
INVx1_ASAP7_75t_L g1267 ( .A(n_1268), .Y(n_1267) );
NAND3xp33_ASAP7_75t_SL g1323 ( .A(n_1268), .B(n_1324), .C(n_1325), .Y(n_1323) );
NOR2xp33_ASAP7_75t_L g1298 ( .A(n_1272), .B(n_1299), .Y(n_1298) );
INVx3_ASAP7_75t_L g1273 ( .A(n_1274), .Y(n_1273) );
AOI21xp33_ASAP7_75t_L g1305 ( .A1(n_1274), .A2(n_1306), .B(n_1308), .Y(n_1305) );
INVx1_ASAP7_75t_L g1277 ( .A(n_1278), .Y(n_1277) );
INVxp67_ASAP7_75t_L g1279 ( .A(n_1280), .Y(n_1279) );
INVx1_ASAP7_75t_L g1284 ( .A(n_1285), .Y(n_1284) );
INVxp67_ASAP7_75t_L g1293 ( .A(n_1294), .Y(n_1293) );
NOR2xp33_ASAP7_75t_L g1294 ( .A(n_1295), .B(n_1296), .Y(n_1294) );
INVx1_ASAP7_75t_L g1320 ( .A(n_1297), .Y(n_1320) );
INVx1_ASAP7_75t_L g1299 ( .A(n_1300), .Y(n_1299) );
NAND5xp2_ASAP7_75t_L g1302 ( .A(n_1303), .B(n_1312), .C(n_1316), .D(n_1322), .E(n_1329), .Y(n_1302) );
INVx2_ASAP7_75t_L g1306 ( .A(n_1307), .Y(n_1306) );
INVx1_ASAP7_75t_L g1308 ( .A(n_1309), .Y(n_1308) );
INVx1_ASAP7_75t_L g1313 ( .A(n_1314), .Y(n_1313) );
INVx1_ASAP7_75t_L g1324 ( .A(n_1315), .Y(n_1324) );
INVx1_ASAP7_75t_L g1317 ( .A(n_1318), .Y(n_1317) );
INVx1_ASAP7_75t_L g1330 ( .A(n_1319), .Y(n_1330) );
OR2x2_ASAP7_75t_L g1319 ( .A(n_1320), .B(n_1321), .Y(n_1319) );
AOI21xp5_ASAP7_75t_L g1322 ( .A1(n_1323), .A2(n_1327), .B(n_1328), .Y(n_1322) );
INVxp67_ASAP7_75t_L g1325 ( .A(n_1326), .Y(n_1325) );
CKINVDCx20_ASAP7_75t_R g1335 ( .A(n_1336), .Y(n_1335) );
CKINVDCx20_ASAP7_75t_R g1336 ( .A(n_1337), .Y(n_1336) );
INVx1_ASAP7_75t_L g1338 ( .A(n_1339), .Y(n_1338) );
OR2x2_ASAP7_75t_L g1340 ( .A(n_1341), .B(n_1377), .Y(n_1340) );
A2O1A1Ixp33_ASAP7_75t_L g1341 ( .A1(n_1342), .A2(n_1362), .B(n_1372), .C(n_1373), .Y(n_1341) );
NOR3xp33_ASAP7_75t_L g1342 ( .A(n_1343), .B(n_1349), .C(n_1356), .Y(n_1342) );
INVx2_ASAP7_75t_L g1344 ( .A(n_1345), .Y(n_1344) );
INVx1_ASAP7_75t_L g1347 ( .A(n_1348), .Y(n_1347) );
INVx1_ASAP7_75t_L g1357 ( .A(n_1358), .Y(n_1357) );
AOI211xp5_ASAP7_75t_SL g1362 ( .A1(n_1363), .A2(n_1364), .B(n_1365), .C(n_1370), .Y(n_1362) );
INVx3_ASAP7_75t_L g1368 ( .A(n_1369), .Y(n_1368) );
NAND2xp5_ASAP7_75t_L g1373 ( .A(n_1374), .B(n_1375), .Y(n_1373) );
INVx1_ASAP7_75t_L g1375 ( .A(n_1376), .Y(n_1375) );
NAND4xp25_ASAP7_75t_L g1377 ( .A(n_1378), .B(n_1383), .C(n_1400), .D(n_1402), .Y(n_1377) );
AND2x4_ASAP7_75t_L g1384 ( .A(n_1385), .B(n_1386), .Y(n_1384) );
INVx1_ASAP7_75t_L g1389 ( .A(n_1390), .Y(n_1389) );
INVx1_ASAP7_75t_L g1391 ( .A(n_1392), .Y(n_1391) );
INVx1_ASAP7_75t_L g1392 ( .A(n_1393), .Y(n_1392) );
AOI21xp5_ASAP7_75t_L g1402 ( .A1(n_1403), .A2(n_1405), .B(n_1406), .Y(n_1402) );
INVx2_ASAP7_75t_L g1403 ( .A(n_1404), .Y(n_1403) );
INVx2_ASAP7_75t_L g1407 ( .A(n_1408), .Y(n_1407) );
BUFx3_ASAP7_75t_L g1408 ( .A(n_1409), .Y(n_1408) );
HB1xp67_ASAP7_75t_L g1413 ( .A(n_1414), .Y(n_1413) );
INVxp33_ASAP7_75t_SL g1415 ( .A(n_1416), .Y(n_1415) );
INVx1_ASAP7_75t_L g1417 ( .A(n_1418), .Y(n_1417) );
HB1xp67_ASAP7_75t_L g1418 ( .A(n_1419), .Y(n_1418) );
NAND3xp33_ASAP7_75t_L g1419 ( .A(n_1420), .B(n_1445), .C(n_1451), .Y(n_1419) );
OAI21xp33_ASAP7_75t_L g1420 ( .A1(n_1421), .A2(n_1434), .B(n_1444), .Y(n_1420) );
INVx2_ASAP7_75t_SL g1422 ( .A(n_1423), .Y(n_1422) );
INVx1_ASAP7_75t_L g1435 ( .A(n_1436), .Y(n_1435) );
INVx4_ASAP7_75t_L g1436 ( .A(n_1437), .Y(n_1436) );
AOI21xp33_ASAP7_75t_SL g1445 ( .A1(n_1446), .A2(n_1448), .B(n_1449), .Y(n_1445) );
INVx8_ASAP7_75t_L g1446 ( .A(n_1447), .Y(n_1446) );
NOR3xp33_ASAP7_75t_L g1451 ( .A(n_1452), .B(n_1468), .C(n_1473), .Y(n_1451) );
NAND2xp5_ASAP7_75t_SL g1452 ( .A(n_1453), .B(n_1463), .Y(n_1452) );
INVx2_ASAP7_75t_L g1455 ( .A(n_1456), .Y(n_1455) );
INVx2_ASAP7_75t_L g1459 ( .A(n_1460), .Y(n_1459) );
AOI22xp33_ASAP7_75t_L g1463 ( .A1(n_1464), .A2(n_1465), .B1(n_1466), .B2(n_1467), .Y(n_1463) );
INVxp67_ASAP7_75t_L g1470 ( .A(n_1471), .Y(n_1470) );
INVx2_ASAP7_75t_SL g1473 ( .A(n_1474), .Y(n_1473) );
HB1xp67_ASAP7_75t_L g1475 ( .A(n_1476), .Y(n_1475) );
OAI21xp5_ASAP7_75t_L g1476 ( .A1(n_1477), .A2(n_1478), .B(n_1479), .Y(n_1476) );
INVx1_ASAP7_75t_L g1479 ( .A(n_1480), .Y(n_1479) );
endmodule