module fake_jpeg_3296_n_227 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_227);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_227;

wire n_159;
wire n_117;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_122;
wire n_75;
wire n_37;
wire n_121;
wire n_102;
wire n_130;
wire n_99;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_192;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g14 ( 
.A(n_0),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_7),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_10),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_9),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_7),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_5),
.Y(n_23)
);

INVxp67_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_7),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_0),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_11),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_5),
.B(n_9),
.Y(n_28)
);

BUFx12_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_3),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_3),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_1),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_32),
.Y(n_37)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_37),
.Y(n_88)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_33),
.Y(n_38)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_38),
.Y(n_99)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_33),
.Y(n_39)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_39),
.Y(n_85)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_32),
.Y(n_40)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_40),
.Y(n_100)
);

INVx11_ASAP7_75t_L g41 ( 
.A(n_18),
.Y(n_41)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_41),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_20),
.B(n_13),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_42),
.B(n_45),
.Y(n_96)
);

BUFx4f_ASAP7_75t_L g43 ( 
.A(n_18),
.Y(n_43)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_43),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_18),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_44),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_28),
.B(n_1),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_31),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g94 ( 
.A(n_46),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_21),
.B(n_12),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_47),
.B(n_53),
.Y(n_106)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_29),
.Y(n_48)
);

INVx5_ASAP7_75t_L g95 ( 
.A(n_48),
.Y(n_95)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_18),
.Y(n_49)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_49),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_30),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_50),
.Y(n_108)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_30),
.Y(n_51)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_51),
.Y(n_78)
);

BUFx10_ASAP7_75t_L g52 ( 
.A(n_30),
.Y(n_52)
);

BUFx8_ASAP7_75t_L g74 ( 
.A(n_52),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_25),
.B(n_2),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_16),
.Y(n_54)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_54),
.Y(n_79)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_30),
.Y(n_55)
);

INVx8_ASAP7_75t_L g102 ( 
.A(n_55),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_35),
.B(n_2),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_56),
.B(n_71),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_17),
.B(n_2),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_57),
.B(n_61),
.Y(n_77)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_24),
.B(n_4),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_58),
.B(n_60),
.Y(n_76)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_24),
.Y(n_59)
);

INVx5_ASAP7_75t_L g75 ( 
.A(n_59),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g60 ( 
.A(n_17),
.B(n_4),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_27),
.B(n_9),
.Y(n_61)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_14),
.Y(n_62)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_62),
.Y(n_93)
);

INVx4_ASAP7_75t_SL g63 ( 
.A(n_29),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g107 ( 
.A(n_63),
.Y(n_107)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_31),
.Y(n_64)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_64),
.Y(n_109)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_14),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_65),
.B(n_68),
.Y(n_105)
);

INVx11_ASAP7_75t_L g66 ( 
.A(n_34),
.Y(n_66)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_66),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g67 ( 
.A(n_27),
.B(n_6),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_67),
.B(n_69),
.Y(n_82)
);

INVx11_ASAP7_75t_L g68 ( 
.A(n_34),
.Y(n_68)
);

INVx5_ASAP7_75t_L g69 ( 
.A(n_29),
.Y(n_69)
);

INVx4_ASAP7_75t_SL g70 ( 
.A(n_23),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_70),
.B(n_8),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_15),
.Y(n_71)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_23),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_72),
.B(n_36),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_15),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_73),
.B(n_6),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_63),
.A2(n_26),
.B1(n_36),
.B2(n_16),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_81),
.A2(n_83),
.B1(n_107),
.B2(n_74),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_66),
.A2(n_39),
.B1(n_38),
.B2(n_43),
.Y(n_83)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_84),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_70),
.B(n_19),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g129 ( 
.A(n_86),
.B(n_90),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_72),
.B(n_19),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_58),
.B(n_22),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_97),
.B(n_98),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_59),
.B(n_22),
.Y(n_98)
);

XOR2xp5_ASAP7_75t_L g101 ( 
.A(n_52),
.B(n_26),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g115 ( 
.A(n_101),
.B(n_76),
.Y(n_115)
);

AO21x1_ASAP7_75t_L g123 ( 
.A1(n_104),
.A2(n_96),
.B(n_106),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_110),
.B(n_107),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_91),
.B(n_73),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_111),
.B(n_112),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_79),
.B(n_71),
.Y(n_112)
);

OAI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_81),
.A2(n_46),
.B1(n_50),
.B2(n_44),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_113),
.A2(n_133),
.B1(n_114),
.B2(n_128),
.Y(n_153)
);

INVx2_ASAP7_75t_SL g114 ( 
.A(n_109),
.Y(n_114)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_114),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_115),
.B(n_117),
.Y(n_148)
);

INVx8_ASAP7_75t_L g116 ( 
.A(n_107),
.Y(n_116)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_116),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_93),
.B(n_55),
.Y(n_117)
);

CKINVDCx16_ASAP7_75t_R g118 ( 
.A(n_74),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_118),
.B(n_120),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_77),
.B(n_8),
.Y(n_120)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_109),
.Y(n_121)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_121),
.Y(n_156)
);

OAI32xp33_ASAP7_75t_L g122 ( 
.A1(n_82),
.A2(n_52),
.A3(n_64),
.B1(n_48),
.B2(n_8),
.Y(n_122)
);

OA22x2_ASAP7_75t_L g143 ( 
.A1(n_122),
.A2(n_131),
.B1(n_137),
.B2(n_80),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_123),
.B(n_125),
.Y(n_155)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_102),
.Y(n_124)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_124),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_88),
.B(n_48),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_100),
.B(n_78),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_127),
.B(n_128),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_75),
.Y(n_128)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_102),
.Y(n_130)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_130),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_105),
.A2(n_94),
.B1(n_103),
.B2(n_99),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_105),
.B(n_89),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_132),
.A2(n_134),
.B1(n_80),
.B2(n_131),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_L g134 ( 
.A1(n_85),
.A2(n_89),
.B1(n_108),
.B2(n_92),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_85),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_135),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_75),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_136),
.Y(n_154)
);

HB1xp67_ASAP7_75t_L g138 ( 
.A(n_94),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_138),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_92),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_139),
.Y(n_152)
);

OAI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_111),
.A2(n_83),
.B1(n_108),
.B2(n_87),
.Y(n_140)
);

AND2x2_ASAP7_75t_L g170 ( 
.A(n_140),
.B(n_153),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_112),
.A2(n_87),
.B1(n_74),
.B2(n_95),
.Y(n_141)
);

AND2x2_ASAP7_75t_L g163 ( 
.A(n_141),
.B(n_143),
.Y(n_163)
);

AND2x2_ASAP7_75t_L g164 ( 
.A(n_144),
.B(n_146),
.Y(n_164)
);

AOI21xp5_ASAP7_75t_L g145 ( 
.A1(n_132),
.A2(n_117),
.B(n_125),
.Y(n_145)
);

AOI21xp5_ASAP7_75t_L g165 ( 
.A1(n_145),
.A2(n_129),
.B(n_114),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_127),
.A2(n_115),
.B1(n_119),
.B2(n_139),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_119),
.A2(n_122),
.B1(n_126),
.B2(n_136),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_147),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_146),
.B(n_123),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_SL g183 ( 
.A(n_162),
.B(n_169),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_165),
.B(n_166),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g166 ( 
.A(n_148),
.B(n_135),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_159),
.B(n_121),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_167),
.B(n_171),
.Y(n_185)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_151),
.Y(n_168)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_168),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_155),
.B(n_124),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_159),
.B(n_130),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_149),
.B(n_116),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_172),
.B(n_174),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_145),
.B(n_158),
.C(n_147),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_154),
.B(n_157),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_175),
.B(n_176),
.Y(n_186)
);

INVxp67_ASAP7_75t_L g176 ( 
.A(n_142),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_151),
.Y(n_177)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_177),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_166),
.B(n_154),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_178),
.B(n_180),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_173),
.B(n_152),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_176),
.Y(n_181)
);

CKINVDCx16_ASAP7_75t_R g198 ( 
.A(n_181),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_164),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_182),
.A2(n_190),
.B1(n_173),
.B2(n_164),
.Y(n_191)
);

BUFx24_ASAP7_75t_L g188 ( 
.A(n_170),
.Y(n_188)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_188),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_174),
.B(n_157),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_191),
.B(n_196),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_182),
.A2(n_163),
.B1(n_164),
.B2(n_170),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_193),
.A2(n_197),
.B1(n_178),
.B2(n_185),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_184),
.B(n_163),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_194),
.B(n_195),
.C(n_187),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_179),
.B(n_163),
.C(n_161),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_180),
.A2(n_143),
.B1(n_153),
.B2(n_150),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_184),
.A2(n_143),
.B1(n_141),
.B2(n_150),
.Y(n_197)
);

AO21x1_ASAP7_75t_L g199 ( 
.A1(n_188),
.A2(n_143),
.B(n_160),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_199),
.B(n_186),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_198),
.B(n_192),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_201),
.B(n_203),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_202),
.A2(n_204),
.B1(n_200),
.B2(n_197),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_195),
.B(n_183),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_192),
.B(n_181),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_205),
.B(n_187),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_206),
.B(n_194),
.Y(n_211)
);

NOR3xp33_ASAP7_75t_SL g208 ( 
.A(n_204),
.B(n_200),
.C(n_188),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_208),
.B(n_209),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_211),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_212),
.Y(n_215)
);

NAND2x1p5_ASAP7_75t_L g216 ( 
.A(n_208),
.B(n_207),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_216),
.B(n_199),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_214),
.B(n_211),
.C(n_210),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_217),
.B(n_218),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_213),
.A2(n_193),
.B1(n_196),
.B2(n_189),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_219),
.A2(n_216),
.B1(n_142),
.B2(n_160),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_215),
.B(n_189),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_SL g222 ( 
.A(n_220),
.B(n_161),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_221),
.B(n_222),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_223),
.B(n_156),
.C(n_221),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_224),
.B(n_156),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_226),
.B(n_225),
.Y(n_227)
);


endmodule