module real_aes_15567_n_102 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_102);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_102;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_838;
wire n_485;
wire n_822;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_364;
wire n_319;
wire n_421;
wire n_555;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_840;
wire n_570;
wire n_675;
wire n_530;
wire n_835;
wire n_104;
wire n_535;
wire n_732;
wire n_834;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_781;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_455;
wire n_310;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_812;
wire n_817;
wire n_565;
wire n_443;
wire n_782;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_754;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_527;
wire n_434;
wire n_502;
wire n_505;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_402;
wire n_552;
wire n_602;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_807;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_832;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_542;
wire n_163;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_288;
wire n_147;
wire n_150;
wire n_404;
wire n_598;
wire n_756;
wire n_713;
wire n_735;
wire n_728;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_810;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_749;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_765;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_831;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_420;
wire n_349;
wire n_336;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_575;
wire n_210;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_103;
wire n_541;
wire n_224;
wire n_839;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_836;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_837;
wire n_474;
wire n_829;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_601;
wire n_500;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_802;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
AND2x4_ASAP7_75t_L g118 ( .A(n_0), .B(n_119), .Y(n_118) );
AOI22xp5_ASAP7_75t_L g510 ( .A1(n_1), .A2(n_3), .B1(n_186), .B2(n_511), .Y(n_510) );
OAI22x1_ASAP7_75t_R g122 ( .A1(n_2), .A2(n_44), .B1(n_123), .B2(n_124), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_2), .Y(n_123) );
AOI22xp33_ASAP7_75t_L g165 ( .A1(n_4), .A2(n_42), .B1(n_143), .B2(n_166), .Y(n_165) );
AOI22xp33_ASAP7_75t_L g485 ( .A1(n_5), .A2(n_25), .B1(n_166), .B2(n_242), .Y(n_485) );
AOI22xp5_ASAP7_75t_L g220 ( .A1(n_6), .A2(n_16), .B1(n_185), .B2(n_221), .Y(n_220) );
AOI22xp33_ASAP7_75t_L g521 ( .A1(n_7), .A2(n_61), .B1(n_203), .B2(n_244), .Y(n_521) );
AOI22xp5_ASAP7_75t_L g527 ( .A1(n_8), .A2(n_17), .B1(n_142), .B2(n_143), .Y(n_527) );
INVx1_ASAP7_75t_L g119 ( .A(n_9), .Y(n_119) );
CKINVDCx5p33_ASAP7_75t_R g581 ( .A(n_10), .Y(n_581) );
CKINVDCx5p33_ASAP7_75t_R g141 ( .A(n_11), .Y(n_141) );
AOI22xp5_ASAP7_75t_L g201 ( .A1(n_12), .A2(n_18), .B1(n_202), .B2(n_205), .Y(n_201) );
OR2x2_ASAP7_75t_L g109 ( .A(n_13), .B(n_38), .Y(n_109) );
BUFx6f_ASAP7_75t_L g144 ( .A(n_14), .Y(n_144) );
CKINVDCx5p33_ASAP7_75t_R g225 ( .A(n_15), .Y(n_225) );
INVx2_ASAP7_75t_L g823 ( .A(n_19), .Y(n_823) );
AOI22xp5_ASAP7_75t_L g184 ( .A1(n_20), .A2(n_100), .B1(n_185), .B2(n_186), .Y(n_184) );
AOI22xp33_ASAP7_75t_L g217 ( .A1(n_21), .A2(n_39), .B1(n_151), .B2(n_218), .Y(n_217) );
NAND2xp5_ASAP7_75t_SL g145 ( .A(n_22), .B(n_146), .Y(n_145) );
OAI21x1_ASAP7_75t_L g137 ( .A1(n_23), .A2(n_57), .B(n_138), .Y(n_137) );
CKINVDCx5p33_ASAP7_75t_R g490 ( .A(n_24), .Y(n_490) );
CKINVDCx5p33_ASAP7_75t_R g195 ( .A(n_26), .Y(n_195) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_27), .B(n_148), .Y(n_497) );
INVx4_ASAP7_75t_R g539 ( .A(n_28), .Y(n_539) );
AOI22xp33_ASAP7_75t_L g170 ( .A1(n_29), .A2(n_47), .B1(n_171), .B2(n_172), .Y(n_170) );
AOI22xp33_ASAP7_75t_L g280 ( .A1(n_30), .A2(n_54), .B1(n_172), .B2(n_185), .Y(n_280) );
CKINVDCx5p33_ASAP7_75t_R g248 ( .A(n_31), .Y(n_248) );
NAND2xp5_ASAP7_75t_L g150 ( .A(n_32), .B(n_151), .Y(n_150) );
CKINVDCx5p33_ASAP7_75t_R g234 ( .A(n_33), .Y(n_234) );
NAND2xp5_ASAP7_75t_SL g504 ( .A(n_34), .B(n_166), .Y(n_504) );
INVx1_ASAP7_75t_L g513 ( .A(n_35), .Y(n_513) );
A2O1A1Ixp33_ASAP7_75t_SL g579 ( .A1(n_36), .A2(n_143), .B(n_147), .C(n_580), .Y(n_579) );
AOI22xp33_ASAP7_75t_L g486 ( .A1(n_37), .A2(n_55), .B1(n_143), .B2(n_172), .Y(n_486) );
AOI22xp5_ASAP7_75t_L g240 ( .A1(n_40), .A2(n_87), .B1(n_143), .B2(n_241), .Y(n_240) );
AOI22xp33_ASAP7_75t_L g206 ( .A1(n_41), .A2(n_46), .B1(n_142), .B2(n_143), .Y(n_206) );
CKINVDCx5p33_ASAP7_75t_R g577 ( .A(n_43), .Y(n_577) );
CKINVDCx5p33_ASAP7_75t_R g124 ( .A(n_44), .Y(n_124) );
AOI22xp33_ASAP7_75t_L g188 ( .A1(n_45), .A2(n_60), .B1(n_185), .B2(n_189), .Y(n_188) );
INVx1_ASAP7_75t_L g501 ( .A(n_48), .Y(n_501) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_49), .B(n_143), .Y(n_503) );
CKINVDCx5p33_ASAP7_75t_R g560 ( .A(n_50), .Y(n_560) );
INVx2_ASAP7_75t_L g117 ( .A(n_51), .Y(n_117) );
CKINVDCx5p33_ASAP7_75t_R g832 ( .A(n_52), .Y(n_832) );
BUFx3_ASAP7_75t_L g108 ( .A(n_53), .Y(n_108) );
INVx1_ASAP7_75t_L g818 ( .A(n_53), .Y(n_818) );
AOI22xp33_ASAP7_75t_L g528 ( .A1(n_56), .A2(n_88), .B1(n_143), .B2(n_172), .Y(n_528) );
CKINVDCx5p33_ASAP7_75t_R g540 ( .A(n_58), .Y(n_540) );
OAI22xp5_ASAP7_75t_L g120 ( .A1(n_59), .A2(n_121), .B1(n_801), .B2(n_802), .Y(n_120) );
INVx1_ASAP7_75t_L g801 ( .A(n_59), .Y(n_801) );
AOI22xp33_ASAP7_75t_L g279 ( .A1(n_62), .A2(n_75), .B1(n_171), .B2(n_189), .Y(n_279) );
CKINVDCx5p33_ASAP7_75t_R g530 ( .A(n_63), .Y(n_530) );
AOI22xp33_ASAP7_75t_L g232 ( .A1(n_64), .A2(n_78), .B1(n_142), .B2(n_143), .Y(n_232) );
AOI22xp5_ASAP7_75t_L g231 ( .A1(n_65), .A2(n_98), .B1(n_185), .B2(n_205), .Y(n_231) );
INVx1_ASAP7_75t_L g138 ( .A(n_66), .Y(n_138) );
AND2x4_ASAP7_75t_L g157 ( .A(n_67), .B(n_158), .Y(n_157) );
AOI22xp5_ASAP7_75t_L g821 ( .A1(n_68), .A2(n_822), .B1(n_823), .B2(n_824), .Y(n_821) );
CKINVDCx5p33_ASAP7_75t_R g824 ( .A(n_68), .Y(n_824) );
AOI22xp33_ASAP7_75t_L g509 ( .A1(n_69), .A2(n_91), .B1(n_171), .B2(n_172), .Y(n_509) );
AO22x1_ASAP7_75t_L g518 ( .A1(n_70), .A2(n_76), .B1(n_218), .B2(n_519), .Y(n_518) );
INVx1_ASAP7_75t_L g158 ( .A(n_71), .Y(n_158) );
AND2x2_ASAP7_75t_L g582 ( .A(n_72), .B(n_160), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g566 ( .A(n_73), .B(n_244), .Y(n_566) );
CKINVDCx5p33_ASAP7_75t_R g575 ( .A(n_74), .Y(n_575) );
CKINVDCx16_ASAP7_75t_R g825 ( .A(n_77), .Y(n_825) );
AOI22xp33_ASAP7_75t_L g833 ( .A1(n_77), .A2(n_89), .B1(n_834), .B2(n_838), .Y(n_833) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_79), .B(n_166), .Y(n_561) );
INVx2_ASAP7_75t_L g148 ( .A(n_80), .Y(n_148) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_81), .B(n_160), .Y(n_494) );
CKINVDCx5p33_ASAP7_75t_R g536 ( .A(n_82), .Y(n_536) );
AOI22xp33_ASAP7_75t_L g243 ( .A1(n_83), .A2(n_99), .B1(n_172), .B2(n_244), .Y(n_243) );
CKINVDCx5p33_ASAP7_75t_R g282 ( .A(n_84), .Y(n_282) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_85), .B(n_193), .Y(n_522) );
CKINVDCx5p33_ASAP7_75t_R g175 ( .A(n_86), .Y(n_175) );
NAND2xp5_ASAP7_75t_SL g159 ( .A(n_90), .B(n_160), .Y(n_159) );
CKINVDCx5p33_ASAP7_75t_R g212 ( .A(n_92), .Y(n_212) );
NAND2xp5_ASAP7_75t_SL g557 ( .A(n_93), .B(n_160), .Y(n_557) );
INVx1_ASAP7_75t_L g113 ( .A(n_94), .Y(n_113) );
NOR2xp33_ASAP7_75t_L g816 ( .A(n_94), .B(n_817), .Y(n_816) );
NAND2xp33_ASAP7_75t_L g153 ( .A(n_95), .B(n_146), .Y(n_153) );
A2O1A1Ixp33_ASAP7_75t_L g534 ( .A1(n_96), .A2(n_208), .B(n_244), .C(n_535), .Y(n_534) );
AND2x2_ASAP7_75t_L g541 ( .A(n_97), .B(n_542), .Y(n_541) );
NAND2xp33_ASAP7_75t_L g565 ( .A(n_101), .B(n_152), .Y(n_565) );
AOI21xp33_ASAP7_75t_L g102 ( .A1(n_103), .A2(n_120), .B(n_803), .Y(n_102) );
BUFx4f_ASAP7_75t_L g103 ( .A(n_104), .Y(n_103) );
INVx3_ASAP7_75t_SL g104 ( .A(n_105), .Y(n_104) );
OR2x2_ASAP7_75t_L g105 ( .A(n_106), .B(n_110), .Y(n_105) );
BUFx2_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
AND2x2_ASAP7_75t_L g111 ( .A(n_107), .B(n_112), .Y(n_111) );
NOR2x1_ASAP7_75t_L g107 ( .A(n_108), .B(n_109), .Y(n_107) );
INVx1_ASAP7_75t_L g819 ( .A(n_109), .Y(n_819) );
OR2x2_ASAP7_75t_L g110 ( .A(n_111), .B(n_114), .Y(n_110) );
AND2x2_ASAP7_75t_L g834 ( .A(n_111), .B(n_835), .Y(n_834) );
HB1xp67_ASAP7_75t_L g473 ( .A(n_112), .Y(n_473) );
CKINVDCx5p33_ASAP7_75t_R g800 ( .A(n_112), .Y(n_800) );
INVx2_ASAP7_75t_L g112 ( .A(n_113), .Y(n_112) );
NOR2xp33_ASAP7_75t_L g835 ( .A(n_114), .B(n_836), .Y(n_835) );
NAND2xp5_ASAP7_75t_SL g114 ( .A(n_115), .B(n_118), .Y(n_114) );
BUFx2_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
NOR2xp33_ASAP7_75t_L g808 ( .A(n_116), .B(n_809), .Y(n_808) );
INVx3_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
NOR2xp33_ASAP7_75t_L g840 ( .A(n_117), .B(n_828), .Y(n_840) );
INVx2_ASAP7_75t_SL g810 ( .A(n_118), .Y(n_810) );
INVx2_ASAP7_75t_L g802 ( .A(n_121), .Y(n_802) );
XNOR2x1_ASAP7_75t_L g121 ( .A(n_122), .B(n_125), .Y(n_121) );
AOI22x1_ASAP7_75t_L g125 ( .A1(n_126), .A2(n_472), .B1(n_474), .B2(n_798), .Y(n_125) );
XNOR2x1_ASAP7_75t_SL g820 ( .A(n_126), .B(n_821), .Y(n_820) );
NAND2x1p5_ASAP7_75t_L g126 ( .A(n_127), .B(n_416), .Y(n_126) );
NOR3x1_ASAP7_75t_L g127 ( .A(n_128), .B(n_334), .C(n_371), .Y(n_127) );
NAND4xp75_ASAP7_75t_L g128 ( .A(n_129), .B(n_254), .C(n_288), .D(n_318), .Y(n_128) );
INVx1_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
OAI32xp33_ASAP7_75t_L g130 ( .A1(n_131), .A2(n_176), .A3(n_226), .B1(n_235), .B2(n_249), .Y(n_130) );
OR2x2_ASAP7_75t_L g235 ( .A(n_131), .B(n_236), .Y(n_235) );
INVx1_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
OAI21xp5_ASAP7_75t_L g445 ( .A1(n_132), .A2(n_446), .B(n_448), .Y(n_445) );
AND2x2_ASAP7_75t_L g132 ( .A(n_133), .B(n_161), .Y(n_132) );
NAND2xp5_ASAP7_75t_L g286 ( .A(n_133), .B(n_287), .Y(n_286) );
AND2x4_ASAP7_75t_L g317 ( .A(n_133), .B(n_263), .Y(n_317) );
AND2x2_ASAP7_75t_L g412 ( .A(n_133), .B(n_228), .Y(n_412) );
INVx2_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
BUFx2_ASAP7_75t_L g261 ( .A(n_134), .Y(n_261) );
OAI21x1_ASAP7_75t_L g134 ( .A1(n_135), .A2(n_139), .B(n_159), .Y(n_134) );
OAI21x1_ASAP7_75t_L g294 ( .A1(n_135), .A2(n_139), .B(n_159), .Y(n_294) );
INVx2_ASAP7_75t_SL g135 ( .A(n_136), .Y(n_135) );
INVx4_ASAP7_75t_L g160 ( .A(n_136), .Y(n_160) );
NOR2xp33_ASAP7_75t_L g174 ( .A(n_136), .B(n_175), .Y(n_174) );
BUFx3_ASAP7_75t_L g223 ( .A(n_136), .Y(n_223) );
NOR2xp33_ASAP7_75t_L g224 ( .A(n_136), .B(n_225), .Y(n_224) );
NOR2xp33_ASAP7_75t_L g233 ( .A(n_136), .B(n_234), .Y(n_233) );
AND2x2_ASAP7_75t_L g505 ( .A(n_136), .B(n_488), .Y(n_505) );
BUFx6f_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
INVx2_ASAP7_75t_L g193 ( .A(n_137), .Y(n_193) );
OAI21x1_ASAP7_75t_L g139 ( .A1(n_140), .A2(n_149), .B(n_155), .Y(n_139) );
O2A1O1Ixp5_ASAP7_75t_L g140 ( .A1(n_141), .A2(n_142), .B(n_145), .C(n_147), .Y(n_140) );
O2A1O1Ixp33_ASAP7_75t_L g559 ( .A1(n_142), .A2(n_560), .B(n_561), .C(n_562), .Y(n_559) );
INVx4_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
INVx1_ASAP7_75t_L g189 ( .A(n_143), .Y(n_189) );
INVx1_ASAP7_75t_L g205 ( .A(n_143), .Y(n_205) );
INVx3_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
BUFx6f_ASAP7_75t_L g146 ( .A(n_144), .Y(n_146) );
BUFx6f_ASAP7_75t_L g152 ( .A(n_144), .Y(n_152) );
BUFx6f_ASAP7_75t_L g166 ( .A(n_144), .Y(n_166) );
BUFx6f_ASAP7_75t_L g172 ( .A(n_144), .Y(n_172) );
INVx1_ASAP7_75t_L g187 ( .A(n_144), .Y(n_187) );
INVx1_ASAP7_75t_L g204 ( .A(n_144), .Y(n_204) );
INVx1_ASAP7_75t_L g219 ( .A(n_144), .Y(n_219) );
INVx1_ASAP7_75t_L g222 ( .A(n_144), .Y(n_222) );
INVx2_ASAP7_75t_L g242 ( .A(n_144), .Y(n_242) );
INVx1_ASAP7_75t_L g244 ( .A(n_144), .Y(n_244) );
INVx3_ASAP7_75t_L g185 ( .A(n_146), .Y(n_185) );
INVxp67_ASAP7_75t_SL g519 ( .A(n_146), .Y(n_519) );
INVx6_ASAP7_75t_L g154 ( .A(n_147), .Y(n_154) );
A2O1A1Ixp33_ASAP7_75t_L g517 ( .A1(n_147), .A2(n_518), .B(n_520), .C(n_523), .Y(n_517) );
AOI21xp5_ASAP7_75t_L g564 ( .A1(n_147), .A2(n_565), .B(n_566), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g591 ( .A(n_147), .B(n_518), .Y(n_591) );
BUFx8_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
INVx2_ASAP7_75t_L g169 ( .A(n_148), .Y(n_169) );
INVx1_ASAP7_75t_L g208 ( .A(n_148), .Y(n_208) );
INVx1_ASAP7_75t_L g500 ( .A(n_148), .Y(n_500) );
AOI21xp5_ASAP7_75t_L g149 ( .A1(n_150), .A2(n_153), .B(n_154), .Y(n_149) );
INVx1_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
INVx2_ASAP7_75t_L g171 ( .A(n_152), .Y(n_171) );
OAI22xp33_ASAP7_75t_L g538 ( .A1(n_152), .A2(n_222), .B1(n_539), .B2(n_540), .Y(n_538) );
OAI22xp5_ASAP7_75t_L g164 ( .A1(n_154), .A2(n_165), .B1(n_167), .B2(n_170), .Y(n_164) );
OAI22xp5_ASAP7_75t_L g183 ( .A1(n_154), .A2(n_167), .B1(n_184), .B2(n_188), .Y(n_183) );
OAI22xp5_ASAP7_75t_L g200 ( .A1(n_154), .A2(n_201), .B1(n_206), .B2(n_207), .Y(n_200) );
OAI22xp5_ASAP7_75t_L g216 ( .A1(n_154), .A2(n_167), .B1(n_217), .B2(n_220), .Y(n_216) );
OAI22xp5_ASAP7_75t_L g230 ( .A1(n_154), .A2(n_207), .B1(n_231), .B2(n_232), .Y(n_230) );
OAI22xp5_ASAP7_75t_L g239 ( .A1(n_154), .A2(n_240), .B1(n_243), .B2(n_245), .Y(n_239) );
OAI22xp5_ASAP7_75t_L g278 ( .A1(n_154), .A2(n_167), .B1(n_279), .B2(n_280), .Y(n_278) );
OAI22xp5_ASAP7_75t_L g484 ( .A1(n_154), .A2(n_485), .B1(n_486), .B2(n_487), .Y(n_484) );
OAI22xp5_ASAP7_75t_L g508 ( .A1(n_154), .A2(n_245), .B1(n_509), .B2(n_510), .Y(n_508) );
OAI22x1_ASAP7_75t_L g526 ( .A1(n_154), .A2(n_245), .B1(n_527), .B2(n_528), .Y(n_526) );
INVx2_ASAP7_75t_SL g155 ( .A(n_156), .Y(n_155) );
INVx2_ASAP7_75t_SL g246 ( .A(n_156), .Y(n_246) );
INVx1_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
BUFx10_ASAP7_75t_L g163 ( .A(n_157), .Y(n_163) );
BUFx10_ASAP7_75t_L g488 ( .A(n_157), .Y(n_488) );
INVx1_ASAP7_75t_L g524 ( .A(n_157), .Y(n_524) );
INVx2_ASAP7_75t_L g173 ( .A(n_160), .Y(n_173) );
NOR2x1_ASAP7_75t_L g567 ( .A(n_160), .B(n_568), .Y(n_567) );
INVx2_ASAP7_75t_L g285 ( .A(n_161), .Y(n_285) );
NAND2xp5_ASAP7_75t_L g293 ( .A(n_161), .B(n_294), .Y(n_293) );
INVx2_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
HB1xp67_ASAP7_75t_L g272 ( .A(n_162), .Y(n_272) );
INVx1_ASAP7_75t_L g316 ( .A(n_162), .Y(n_316) );
AND2x2_ASAP7_75t_L g360 ( .A(n_162), .B(n_294), .Y(n_360) );
OR2x2_ASAP7_75t_L g414 ( .A(n_162), .B(n_238), .Y(n_414) );
AO31x2_ASAP7_75t_L g162 ( .A1(n_163), .A2(n_164), .A3(n_173), .B(n_174), .Y(n_162) );
INVx2_ASAP7_75t_L g182 ( .A(n_163), .Y(n_182) );
AO31x2_ASAP7_75t_L g199 ( .A1(n_163), .A2(n_200), .A3(n_209), .B(n_211), .Y(n_199) );
AO31x2_ASAP7_75t_L g215 ( .A1(n_163), .A2(n_216), .A3(n_223), .B(n_224), .Y(n_215) );
AO31x2_ASAP7_75t_L g525 ( .A1(n_163), .A2(n_196), .A3(n_526), .B(n_529), .Y(n_525) );
NOR2xp33_ASAP7_75t_L g574 ( .A(n_166), .B(n_575), .Y(n_574) );
INVx2_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
INVx2_ASAP7_75t_L g487 ( .A(n_168), .Y(n_487) );
BUFx3_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
INVx2_ASAP7_75t_L g563 ( .A(n_169), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g498 ( .A(n_172), .B(n_499), .Y(n_498) );
INVx2_ASAP7_75t_L g511 ( .A(n_172), .Y(n_511) );
AO31x2_ASAP7_75t_L g483 ( .A1(n_173), .A2(n_484), .A3(n_488), .B(n_489), .Y(n_483) );
INVx1_ASAP7_75t_L g176 ( .A(n_177), .Y(n_176) );
AOI22xp33_ASAP7_75t_L g431 ( .A1(n_177), .A2(n_340), .B1(n_432), .B2(n_434), .Y(n_431) );
AND2x2_ASAP7_75t_L g177 ( .A(n_178), .B(n_197), .Y(n_177) );
INVx4_ASAP7_75t_L g257 ( .A(n_178), .Y(n_257) );
AOI22xp5_ASAP7_75t_L g268 ( .A1(n_178), .A2(n_237), .B1(n_269), .B2(n_271), .Y(n_268) );
OR2x2_ASAP7_75t_L g274 ( .A(n_178), .B(n_275), .Y(n_274) );
AND2x2_ASAP7_75t_L g393 ( .A(n_178), .B(n_292), .Y(n_393) );
INVx3_ASAP7_75t_L g178 ( .A(n_179), .Y(n_178) );
AND2x2_ASAP7_75t_L g313 ( .A(n_179), .B(n_198), .Y(n_313) );
AND2x2_ASAP7_75t_L g404 ( .A(n_179), .B(n_276), .Y(n_404) );
AND2x2_ASAP7_75t_L g459 ( .A(n_179), .B(n_215), .Y(n_459) );
INVx2_ASAP7_75t_L g179 ( .A(n_180), .Y(n_179) );
INVx2_ASAP7_75t_L g253 ( .A(n_180), .Y(n_253) );
AND2x4_ASAP7_75t_L g380 ( .A(n_180), .B(n_276), .Y(n_380) );
AO31x2_ASAP7_75t_L g180 ( .A1(n_181), .A2(n_183), .A3(n_190), .B(n_194), .Y(n_180) );
AO31x2_ASAP7_75t_L g229 ( .A1(n_181), .A2(n_209), .A3(n_230), .B(n_233), .Y(n_229) );
INVx1_ASAP7_75t_L g181 ( .A(n_182), .Y(n_181) );
AOI21xp5_ASAP7_75t_L g533 ( .A1(n_182), .A2(n_534), .B(n_537), .Y(n_533) );
INVx2_ASAP7_75t_L g186 ( .A(n_187), .Y(n_186) );
NOR2xp33_ASAP7_75t_L g576 ( .A(n_187), .B(n_577), .Y(n_576) );
AO31x2_ASAP7_75t_L g277 ( .A1(n_190), .A2(n_246), .A3(n_278), .B(n_281), .Y(n_277) );
AO21x2_ASAP7_75t_L g532 ( .A1(n_190), .A2(n_533), .B(n_541), .Y(n_532) );
INVx2_ASAP7_75t_L g190 ( .A(n_191), .Y(n_190) );
INVx2_ASAP7_75t_L g191 ( .A(n_192), .Y(n_191) );
NOR2xp33_ASAP7_75t_SL g211 ( .A(n_192), .B(n_212), .Y(n_211) );
NOR2xp33_ASAP7_75t_L g247 ( .A(n_192), .B(n_248), .Y(n_247) );
INVx2_ASAP7_75t_L g192 ( .A(n_193), .Y(n_192) );
INVx2_ASAP7_75t_L g196 ( .A(n_193), .Y(n_196) );
INVx2_ASAP7_75t_L g210 ( .A(n_193), .Y(n_210) );
OAI21xp33_ASAP7_75t_L g523 ( .A1(n_193), .A2(n_522), .B(n_524), .Y(n_523) );
NOR2xp33_ASAP7_75t_L g194 ( .A(n_195), .B(n_196), .Y(n_194) );
NOR2xp33_ASAP7_75t_L g281 ( .A(n_196), .B(n_282), .Y(n_281) );
NAND2x1_ASAP7_75t_L g256 ( .A(n_197), .B(n_257), .Y(n_256) );
NAND2xp5_ASAP7_75t_SL g363 ( .A(n_197), .B(n_364), .Y(n_363) );
AND2x4_ASAP7_75t_L g197 ( .A(n_198), .B(n_213), .Y(n_197) );
INVx2_ASAP7_75t_L g251 ( .A(n_198), .Y(n_251) );
NAND2xp5_ASAP7_75t_L g275 ( .A(n_198), .B(n_276), .Y(n_275) );
INVx1_ASAP7_75t_L g299 ( .A(n_198), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g326 ( .A(n_198), .B(n_301), .Y(n_326) );
AND2x2_ASAP7_75t_L g329 ( .A(n_198), .B(n_330), .Y(n_329) );
INVx1_ASAP7_75t_L g389 ( .A(n_198), .Y(n_389) );
INVx4_ASAP7_75t_SL g198 ( .A(n_199), .Y(n_198) );
NAND2xp5_ASAP7_75t_L g267 ( .A(n_199), .B(n_214), .Y(n_267) );
BUFx2_ASAP7_75t_L g305 ( .A(n_199), .Y(n_305) );
AND2x2_ASAP7_75t_L g354 ( .A(n_199), .B(n_215), .Y(n_354) );
AND2x2_ASAP7_75t_L g396 ( .A(n_199), .B(n_277), .Y(n_396) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_199), .B(n_429), .Y(n_428) );
INVx1_ASAP7_75t_L g202 ( .A(n_203), .Y(n_202) );
INVx2_ASAP7_75t_L g203 ( .A(n_204), .Y(n_203) );
NOR2xp33_ASAP7_75t_L g535 ( .A(n_204), .B(n_536), .Y(n_535) );
INVx1_ASAP7_75t_SL g207 ( .A(n_208), .Y(n_207) );
INVx1_ASAP7_75t_L g245 ( .A(n_208), .Y(n_245) );
AO31x2_ASAP7_75t_L g507 ( .A1(n_209), .A2(n_246), .A3(n_508), .B(n_512), .Y(n_507) );
AOI21x1_ASAP7_75t_L g571 ( .A1(n_209), .A2(n_572), .B(n_582), .Y(n_571) );
BUFx2_ASAP7_75t_L g209 ( .A(n_210), .Y(n_209) );
NOR2xp33_ASAP7_75t_L g489 ( .A(n_210), .B(n_490), .Y(n_489) );
NOR2xp33_ASAP7_75t_L g512 ( .A(n_210), .B(n_513), .Y(n_512) );
NOR2xp33_ASAP7_75t_L g529 ( .A(n_210), .B(n_530), .Y(n_529) );
INVx2_ASAP7_75t_L g542 ( .A(n_210), .Y(n_542) );
INVx1_ASAP7_75t_L g213 ( .A(n_214), .Y(n_213) );
INVx1_ASAP7_75t_L g214 ( .A(n_215), .Y(n_214) );
NAND2xp5_ASAP7_75t_L g300 ( .A(n_215), .B(n_301), .Y(n_300) );
OR2x2_ASAP7_75t_L g307 ( .A(n_215), .B(n_277), .Y(n_307) );
INVx1_ASAP7_75t_L g330 ( .A(n_215), .Y(n_330) );
INVx2_ASAP7_75t_L g350 ( .A(n_215), .Y(n_350) );
HB1xp67_ASAP7_75t_L g395 ( .A(n_215), .Y(n_395) );
OAI21xp33_ASAP7_75t_SL g496 ( .A1(n_218), .A2(n_497), .B(n_498), .Y(n_496) );
INVx1_ASAP7_75t_L g218 ( .A(n_219), .Y(n_218) );
INVx1_ASAP7_75t_L g221 ( .A(n_222), .Y(n_221) );
AO31x2_ASAP7_75t_L g238 ( .A1(n_223), .A2(n_239), .A3(n_246), .B(n_247), .Y(n_238) );
INVx1_ASAP7_75t_L g226 ( .A(n_227), .Y(n_226) );
AND2x2_ASAP7_75t_L g314 ( .A(n_227), .B(n_315), .Y(n_314) );
NOR2x1p5_ASAP7_75t_L g420 ( .A(n_227), .B(n_414), .Y(n_420) );
INVx2_ASAP7_75t_L g227 ( .A(n_228), .Y(n_227) );
AND2x4_ASAP7_75t_L g237 ( .A(n_228), .B(n_238), .Y(n_237) );
INVx3_ASAP7_75t_L g270 ( .A(n_228), .Y(n_270) );
NAND2xp5_ASAP7_75t_L g284 ( .A(n_228), .B(n_285), .Y(n_284) );
NAND2xp5_ASAP7_75t_L g345 ( .A(n_228), .B(n_346), .Y(n_345) );
INVx3_ASAP7_75t_L g228 ( .A(n_229), .Y(n_228) );
AND2x2_ASAP7_75t_L g262 ( .A(n_229), .B(n_263), .Y(n_262) );
AND2x2_ASAP7_75t_L g320 ( .A(n_229), .B(n_238), .Y(n_320) );
BUFx2_ASAP7_75t_L g433 ( .A(n_229), .Y(n_433) );
NAND2xp5_ASAP7_75t_L g258 ( .A(n_235), .B(n_259), .Y(n_258) );
INVx1_ASAP7_75t_L g471 ( .A(n_235), .Y(n_471) );
INVx2_ASAP7_75t_SL g236 ( .A(n_237), .Y(n_236) );
INVx1_ASAP7_75t_L g407 ( .A(n_237), .Y(n_407) );
AND2x4_ASAP7_75t_L g430 ( .A(n_237), .B(n_360), .Y(n_430) );
AND2x2_ASAP7_75t_L g454 ( .A(n_237), .B(n_455), .Y(n_454) );
INVx2_ASAP7_75t_L g263 ( .A(n_238), .Y(n_263) );
BUFx2_ASAP7_75t_L g287 ( .A(n_238), .Y(n_287) );
INVx1_ASAP7_75t_L g343 ( .A(n_238), .Y(n_343) );
OR2x2_ASAP7_75t_L g465 ( .A(n_238), .B(n_322), .Y(n_465) );
INVx2_ASAP7_75t_SL g241 ( .A(n_242), .Y(n_241) );
NOR2xp33_ASAP7_75t_L g580 ( .A(n_242), .B(n_581), .Y(n_580) );
NAND2xp5_ASAP7_75t_SL g537 ( .A(n_245), .B(n_538), .Y(n_537) );
HB1xp67_ASAP7_75t_L g249 ( .A(n_250), .Y(n_249) );
NAND2xp5_ASAP7_75t_L g250 ( .A(n_251), .B(n_252), .Y(n_250) );
INVx2_ASAP7_75t_L g311 ( .A(n_251), .Y(n_311) );
HB1xp67_ASAP7_75t_L g328 ( .A(n_252), .Y(n_328) );
INVx1_ASAP7_75t_L g332 ( .A(n_252), .Y(n_332) );
INVx1_ASAP7_75t_L g252 ( .A(n_253), .Y(n_252) );
INVx2_ASAP7_75t_L g273 ( .A(n_253), .Y(n_273) );
OR2x2_ASAP7_75t_L g310 ( .A(n_253), .B(n_302), .Y(n_310) );
AOI21xp5_ASAP7_75t_L g254 ( .A1(n_255), .A2(n_258), .B(n_264), .Y(n_254) );
INVx2_ASAP7_75t_L g255 ( .A(n_256), .Y(n_255) );
OAI22xp5_ASAP7_75t_L g352 ( .A1(n_259), .A2(n_353), .B1(n_355), .B2(n_358), .Y(n_352) );
INVx1_ASAP7_75t_L g259 ( .A(n_260), .Y(n_259) );
AND2x2_ASAP7_75t_L g260 ( .A(n_261), .B(n_262), .Y(n_260) );
OR2x2_ASAP7_75t_L g398 ( .A(n_261), .B(n_399), .Y(n_398) );
INVx1_ASAP7_75t_L g406 ( .A(n_261), .Y(n_406) );
AND2x2_ASAP7_75t_L g419 ( .A(n_261), .B(n_420), .Y(n_419) );
AND2x2_ASAP7_75t_L g381 ( .A(n_262), .B(n_360), .Y(n_381) );
OAI22xp5_ASAP7_75t_L g264 ( .A1(n_265), .A2(n_268), .B1(n_274), .B2(n_283), .Y(n_264) );
INVx1_ASAP7_75t_L g265 ( .A(n_266), .Y(n_265) );
INVx1_ASAP7_75t_L g266 ( .A(n_267), .Y(n_266) );
INVx1_ASAP7_75t_L g333 ( .A(n_267), .Y(n_333) );
INVx1_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
AND2x4_ASAP7_75t_L g291 ( .A(n_270), .B(n_292), .Y(n_291) );
AND2x2_ASAP7_75t_L g359 ( .A(n_270), .B(n_360), .Y(n_359) );
INVx2_ASAP7_75t_L g368 ( .A(n_270), .Y(n_368) );
NAND2xp5_ASAP7_75t_L g384 ( .A(n_270), .B(n_385), .Y(n_384) );
NAND2xp5_ASAP7_75t_L g439 ( .A(n_271), .B(n_440), .Y(n_439) );
AND2x2_ASAP7_75t_L g271 ( .A(n_272), .B(n_273), .Y(n_271) );
AND2x2_ASAP7_75t_L g356 ( .A(n_273), .B(n_357), .Y(n_356) );
INVx3_ASAP7_75t_L g370 ( .A(n_273), .Y(n_370) );
INVx2_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
INVx2_ASAP7_75t_L g302 ( .A(n_277), .Y(n_302) );
AND2x4_ASAP7_75t_L g349 ( .A(n_277), .B(n_350), .Y(n_349) );
HB1xp67_ASAP7_75t_L g365 ( .A(n_277), .Y(n_365) );
INVx1_ASAP7_75t_L g429 ( .A(n_277), .Y(n_429) );
OR2x2_ASAP7_75t_L g283 ( .A(n_284), .B(n_286), .Y(n_283) );
AND2x4_ASAP7_75t_L g321 ( .A(n_285), .B(n_322), .Y(n_321) );
INVx1_ASAP7_75t_L g338 ( .A(n_285), .Y(n_338) );
INVx1_ASAP7_75t_L g296 ( .A(n_287), .Y(n_296) );
AOI22xp5_ASAP7_75t_L g288 ( .A1(n_289), .A2(n_297), .B1(n_308), .B2(n_314), .Y(n_288) );
INVx1_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
NAND2x1p5_ASAP7_75t_L g290 ( .A(n_291), .B(n_295), .Y(n_290) );
INVx1_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
INVxp67_ASAP7_75t_SL g346 ( .A(n_293), .Y(n_346) );
INVx1_ASAP7_75t_L g322 ( .A(n_294), .Y(n_322) );
INVx1_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
NAND2xp5_ASAP7_75t_SL g297 ( .A(n_298), .B(n_303), .Y(n_297) );
OR2x2_ASAP7_75t_L g298 ( .A(n_299), .B(n_300), .Y(n_298) );
NAND2xp5_ASAP7_75t_L g348 ( .A(n_299), .B(n_349), .Y(n_348) );
INVx1_ASAP7_75t_L g451 ( .A(n_300), .Y(n_451) );
INVx1_ASAP7_75t_L g470 ( .A(n_300), .Y(n_470) );
INVx1_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
INVx1_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
NAND2x1_ASAP7_75t_L g447 ( .A(n_304), .B(n_370), .Y(n_447) );
AND2x4_ASAP7_75t_L g304 ( .A(n_305), .B(n_306), .Y(n_304) );
INVx1_ASAP7_75t_L g463 ( .A(n_305), .Y(n_463) );
INVx2_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
NAND2xp5_ASAP7_75t_L g308 ( .A(n_309), .B(n_312), .Y(n_308) );
INVx2_ASAP7_75t_L g401 ( .A(n_309), .Y(n_401) );
OR2x2_ASAP7_75t_L g309 ( .A(n_310), .B(n_311), .Y(n_309) );
INVx2_ASAP7_75t_L g390 ( .A(n_310), .Y(n_390) );
AND2x4_ASAP7_75t_L g392 ( .A(n_311), .B(n_349), .Y(n_392) );
INVx1_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
AOI22xp5_ASAP7_75t_L g460 ( .A1(n_315), .A2(n_461), .B1(n_464), .B2(n_466), .Y(n_460) );
AND2x4_ASAP7_75t_L g315 ( .A(n_316), .B(n_317), .Y(n_315) );
INVx2_ASAP7_75t_L g385 ( .A(n_316), .Y(n_385) );
INVx1_ASAP7_75t_L g339 ( .A(n_317), .Y(n_339) );
AND2x4_ASAP7_75t_L g432 ( .A(n_317), .B(n_433), .Y(n_432) );
AND2x2_ASAP7_75t_L g440 ( .A(n_317), .B(n_441), .Y(n_440) );
NAND2xp5_ASAP7_75t_L g318 ( .A(n_319), .B(n_323), .Y(n_318) );
AND2x4_ASAP7_75t_SL g319 ( .A(n_320), .B(n_321), .Y(n_319) );
INVx1_ASAP7_75t_SL g383 ( .A(n_320), .Y(n_383) );
INVx2_ASAP7_75t_L g399 ( .A(n_320), .Y(n_399) );
INVx1_ASAP7_75t_L g426 ( .A(n_321), .Y(n_426) );
AND2x2_ASAP7_75t_L g457 ( .A(n_321), .B(n_368), .Y(n_457) );
NAND3xp33_ASAP7_75t_L g323 ( .A(n_324), .B(n_327), .C(n_331), .Y(n_323) );
INVx1_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
INVx1_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
NAND2xp5_ASAP7_75t_L g327 ( .A(n_328), .B(n_329), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g353 ( .A(n_328), .B(n_354), .Y(n_353) );
AND2x2_ASAP7_75t_L g369 ( .A(n_329), .B(n_370), .Y(n_369) );
NAND2xp5_ASAP7_75t_L g437 ( .A(n_329), .B(n_404), .Y(n_437) );
INVx1_ASAP7_75t_L g357 ( .A(n_330), .Y(n_357) );
NAND2xp5_ASAP7_75t_L g331 ( .A(n_332), .B(n_333), .Y(n_331) );
NAND2xp5_ASAP7_75t_L g422 ( .A(n_332), .B(n_396), .Y(n_422) );
INVx1_ASAP7_75t_L g377 ( .A(n_333), .Y(n_377) );
NAND3xp33_ASAP7_75t_L g334 ( .A(n_335), .B(n_351), .C(n_361), .Y(n_334) );
OAI21xp5_ASAP7_75t_L g335 ( .A1(n_336), .A2(n_340), .B(n_347), .Y(n_335) );
INVxp67_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
OR2x2_ASAP7_75t_L g337 ( .A(n_338), .B(n_339), .Y(n_337) );
INVx1_ASAP7_75t_L g455 ( .A(n_338), .Y(n_455) );
AND2x4_ASAP7_75t_L g340 ( .A(n_341), .B(n_344), .Y(n_340) );
INVx1_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
AOI32xp33_ASAP7_75t_L g391 ( .A1(n_342), .A2(n_392), .A3(n_393), .B1(n_394), .B2(n_397), .Y(n_391) );
NOR2xp33_ASAP7_75t_L g425 ( .A(n_342), .B(n_426), .Y(n_425) );
BUFx2_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
INVx1_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
INVx1_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
INVx2_ASAP7_75t_L g375 ( .A(n_349), .Y(n_375) );
NAND2x1p5_ASAP7_75t_L g410 ( .A(n_349), .B(n_370), .Y(n_410) );
INVx1_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_354), .B(n_404), .Y(n_403) );
AND2x2_ASAP7_75t_L g415 ( .A(n_354), .B(n_364), .Y(n_415) );
INVx1_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
INVx1_ASAP7_75t_L g443 ( .A(n_357), .Y(n_443) );
INVx1_ASAP7_75t_SL g358 ( .A(n_359), .Y(n_358) );
AOI22xp33_ASAP7_75t_SL g361 ( .A1(n_359), .A2(n_362), .B1(n_366), .B2(n_369), .Y(n_361) );
NAND2xp5_ASAP7_75t_L g367 ( .A(n_360), .B(n_368), .Y(n_367) );
AOI22xp5_ASAP7_75t_L g456 ( .A1(n_362), .A2(n_420), .B1(n_457), .B2(n_458), .Y(n_456) );
INVx1_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
AND2x2_ASAP7_75t_L g458 ( .A(n_364), .B(n_459), .Y(n_458) );
INVx1_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
AOI22xp33_ASAP7_75t_L g408 ( .A1(n_366), .A2(n_409), .B1(n_411), .B2(n_415), .Y(n_408) );
INVx2_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
INVx2_ASAP7_75t_L g450 ( .A(n_370), .Y(n_450) );
NAND4xp25_ASAP7_75t_L g371 ( .A(n_372), .B(n_391), .C(n_400), .D(n_408), .Y(n_371) );
O2A1O1Ixp5_ASAP7_75t_L g372 ( .A1(n_373), .A2(n_378), .B(n_381), .C(n_382), .Y(n_372) );
NOR2x1_ASAP7_75t_L g373 ( .A(n_374), .B(n_376), .Y(n_373) );
INVx1_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
INVx1_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
INVx2_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
INVx3_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
AND2x4_ASAP7_75t_L g436 ( .A(n_380), .B(n_395), .Y(n_436) );
NAND2xp5_ASAP7_75t_L g462 ( .A(n_380), .B(n_463), .Y(n_462) );
AOI21xp5_ASAP7_75t_L g382 ( .A1(n_383), .A2(n_384), .B(n_386), .Y(n_382) );
INVx1_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
AOI22xp5_ASAP7_75t_L g424 ( .A1(n_387), .A2(n_425), .B1(n_427), .B2(n_430), .Y(n_424) );
AND2x4_ASAP7_75t_L g387 ( .A(n_388), .B(n_390), .Y(n_387) );
INVx1_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
OAI21xp5_ASAP7_75t_L g453 ( .A1(n_392), .A2(n_397), .B(n_454), .Y(n_453) );
AND2x4_ASAP7_75t_L g394 ( .A(n_395), .B(n_396), .Y(n_394) );
INVx1_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
OAI21xp33_ASAP7_75t_L g400 ( .A1(n_401), .A2(n_402), .B(n_405), .Y(n_400) );
INVx2_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
NOR2xp33_ASAP7_75t_R g405 ( .A(n_406), .B(n_407), .Y(n_405) );
INVx2_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
AND2x2_ASAP7_75t_L g411 ( .A(n_412), .B(n_413), .Y(n_411) );
INVx1_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
AOI22xp5_ASAP7_75t_L g468 ( .A1(n_415), .A2(n_432), .B1(n_469), .B2(n_471), .Y(n_468) );
NOR3x1_ASAP7_75t_L g416 ( .A(n_417), .B(n_438), .C(n_452), .Y(n_416) );
NAND2xp5_ASAP7_75t_L g417 ( .A(n_418), .B(n_431), .Y(n_417) );
AOI21xp33_ASAP7_75t_L g418 ( .A1(n_419), .A2(n_421), .B(n_423), .Y(n_418) );
INVx1_ASAP7_75t_L g444 ( .A(n_419), .Y(n_444) );
INVx2_ASAP7_75t_SL g421 ( .A(n_422), .Y(n_421) );
INVxp67_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
INVx1_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
INVx1_ASAP7_75t_L g467 ( .A(n_429), .Y(n_467) );
INVx1_ASAP7_75t_L g441 ( .A(n_433), .Y(n_441) );
NAND2xp5_ASAP7_75t_L g434 ( .A(n_435), .B(n_437), .Y(n_434) );
OAI221xp5_ASAP7_75t_L g438 ( .A1(n_435), .A2(n_439), .B1(n_442), .B2(n_444), .C(n_445), .Y(n_438) );
INVx1_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
INVx1_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
INVx1_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
INVx2_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
NAND2xp5_ASAP7_75t_L g449 ( .A(n_450), .B(n_451), .Y(n_449) );
NAND4xp25_ASAP7_75t_SL g452 ( .A(n_453), .B(n_456), .C(n_460), .D(n_468), .Y(n_452) );
AND2x2_ASAP7_75t_L g466 ( .A(n_459), .B(n_467), .Y(n_466) );
INVxp67_ASAP7_75t_SL g461 ( .A(n_462), .Y(n_461) );
INVxp67_ASAP7_75t_SL g464 ( .A(n_465), .Y(n_464) );
HB1xp67_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
INVx1_ASAP7_75t_SL g472 ( .A(n_473), .Y(n_472) );
INVx2_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
AND2x4_ASAP7_75t_L g475 ( .A(n_476), .B(n_675), .Y(n_475) );
NOR2x1_ASAP7_75t_L g476 ( .A(n_477), .B(n_623), .Y(n_476) );
OAI211xp5_ASAP7_75t_L g477 ( .A1(n_478), .A2(n_514), .B(n_543), .C(n_608), .Y(n_477) );
HB1xp67_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
INVx1_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
OAI21xp5_ASAP7_75t_L g758 ( .A1(n_480), .A2(n_544), .B(n_759), .Y(n_758) );
AND2x4_ASAP7_75t_L g480 ( .A(n_481), .B(n_491), .Y(n_480) );
INVx2_ASAP7_75t_L g604 ( .A(n_481), .Y(n_604) );
NOR2xp33_ASAP7_75t_L g778 ( .A(n_481), .B(n_779), .Y(n_778) );
INVx2_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
AND2x2_ASAP7_75t_L g715 ( .A(n_482), .B(n_493), .Y(n_715) );
BUFx2_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
INVx2_ASAP7_75t_SL g583 ( .A(n_483), .Y(n_583) );
NAND2xp5_ASAP7_75t_L g620 ( .A(n_483), .B(n_507), .Y(n_620) );
AND2x2_ASAP7_75t_L g653 ( .A(n_483), .B(n_570), .Y(n_653) );
OR2x2_ASAP7_75t_L g658 ( .A(n_483), .B(n_507), .Y(n_658) );
AOI21xp5_ASAP7_75t_L g502 ( .A1(n_487), .A2(n_503), .B(n_504), .Y(n_502) );
OAI21x1_ASAP7_75t_L g520 ( .A1(n_487), .A2(n_521), .B(n_522), .Y(n_520) );
INVx1_ASAP7_75t_L g568 ( .A(n_488), .Y(n_568) );
INVx1_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
INVx1_ASAP7_75t_L g797 ( .A(n_492), .Y(n_797) );
OR2x2_ASAP7_75t_L g492 ( .A(n_493), .B(n_506), .Y(n_492) );
AND2x2_ASAP7_75t_L g598 ( .A(n_493), .B(n_507), .Y(n_598) );
INVx3_ASAP7_75t_L g606 ( .A(n_493), .Y(n_606) );
NAND2x1p5_ASAP7_75t_SL g638 ( .A(n_493), .B(n_622), .Y(n_638) );
INVx1_ASAP7_75t_L g656 ( .A(n_493), .Y(n_656) );
NAND2xp5_ASAP7_75t_L g681 ( .A(n_493), .B(n_601), .Y(n_681) );
BUFx2_ASAP7_75t_L g767 ( .A(n_493), .Y(n_767) );
AND2x4_ASAP7_75t_L g493 ( .A(n_494), .B(n_495), .Y(n_493) );
OAI21xp5_ASAP7_75t_L g495 ( .A1(n_496), .A2(n_502), .B(n_505), .Y(n_495) );
NOR2xp33_ASAP7_75t_L g499 ( .A(n_500), .B(n_501), .Y(n_499) );
BUFx4f_ASAP7_75t_L g578 ( .A(n_500), .Y(n_578) );
INVx1_ASAP7_75t_L g506 ( .A(n_507), .Y(n_506) );
INVx1_ASAP7_75t_L g551 ( .A(n_507), .Y(n_551) );
INVx1_ASAP7_75t_L g607 ( .A(n_507), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g680 ( .A(n_507), .B(n_583), .Y(n_680) );
NOR2xp33_ASAP7_75t_L g716 ( .A(n_507), .B(n_570), .Y(n_716) );
OR2x2_ASAP7_75t_L g514 ( .A(n_515), .B(n_531), .Y(n_514) );
INVx1_ASAP7_75t_L g774 ( .A(n_515), .Y(n_774) );
NAND2xp5_ASAP7_75t_L g515 ( .A(n_516), .B(n_525), .Y(n_515) );
OR2x2_ASAP7_75t_L g546 ( .A(n_516), .B(n_547), .Y(n_546) );
INVx2_ASAP7_75t_L g611 ( .A(n_516), .Y(n_611) );
INVx1_ASAP7_75t_L g516 ( .A(n_517), .Y(n_516) );
INVx1_ASAP7_75t_L g590 ( .A(n_520), .Y(n_590) );
INVx1_ASAP7_75t_L g592 ( .A(n_523), .Y(n_592) );
AOI21xp5_ASAP7_75t_L g572 ( .A1(n_524), .A2(n_573), .B(n_579), .Y(n_572) );
INVx2_ASAP7_75t_L g547 ( .A(n_525), .Y(n_547) );
OR2x2_ASAP7_75t_L g612 ( .A(n_525), .B(n_532), .Y(n_612) );
AND2x2_ASAP7_75t_L g617 ( .A(n_525), .B(n_532), .Y(n_617) );
INVx2_ASAP7_75t_L g662 ( .A(n_525), .Y(n_662) );
AND2x2_ASAP7_75t_L g703 ( .A(n_525), .B(n_556), .Y(n_703) );
AND2x2_ASAP7_75t_L g737 ( .A(n_525), .B(n_634), .Y(n_737) );
INVx1_ASAP7_75t_L g548 ( .A(n_531), .Y(n_548) );
INVx1_ASAP7_75t_L g667 ( .A(n_531), .Y(n_667) );
INVx1_ASAP7_75t_L g531 ( .A(n_532), .Y(n_531) );
AND2x2_ASAP7_75t_L g587 ( .A(n_532), .B(n_588), .Y(n_587) );
AND2x4_ASAP7_75t_L g628 ( .A(n_532), .B(n_589), .Y(n_628) );
INVx2_ASAP7_75t_L g634 ( .A(n_532), .Y(n_634) );
AND2x2_ASAP7_75t_L g689 ( .A(n_532), .B(n_556), .Y(n_689) );
AND2x2_ASAP7_75t_L g746 ( .A(n_532), .B(n_555), .Y(n_746) );
AOI22xp5_ASAP7_75t_L g543 ( .A1(n_544), .A2(n_549), .B1(n_584), .B2(n_595), .Y(n_543) );
INVx3_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
OR2x2_ASAP7_75t_L g545 ( .A(n_546), .B(n_548), .Y(n_545) );
NAND3xp33_ASAP7_75t_SL g724 ( .A(n_546), .B(n_725), .C(n_727), .Y(n_724) );
INVx1_ASAP7_75t_L g643 ( .A(n_547), .Y(n_643) );
AND2x2_ASAP7_75t_L g693 ( .A(n_547), .B(n_555), .Y(n_693) );
INVx1_ASAP7_75t_L g793 ( .A(n_548), .Y(n_793) );
AND2x2_ASAP7_75t_L g549 ( .A(n_550), .B(n_552), .Y(n_549) );
NOR2xp33_ASAP7_75t_L g784 ( .A(n_550), .B(n_748), .Y(n_784) );
BUFx3_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
INVx1_ASAP7_75t_L g639 ( .A(n_551), .Y(n_639) );
INVx1_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
OR2x2_ASAP7_75t_L g553 ( .A(n_554), .B(n_569), .Y(n_553) );
INVx1_ASAP7_75t_L g627 ( .A(n_554), .Y(n_627) );
BUFx2_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
AND2x2_ASAP7_75t_L g707 ( .A(n_555), .B(n_588), .Y(n_707) );
AND2x2_ASAP7_75t_L g726 ( .A(n_555), .B(n_633), .Y(n_726) );
INVx2_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
INVx1_ASAP7_75t_L g594 ( .A(n_556), .Y(n_594) );
BUFx3_ASAP7_75t_L g632 ( .A(n_556), .Y(n_632) );
AND2x2_ASAP7_75t_L g661 ( .A(n_556), .B(n_662), .Y(n_661) );
NAND2x1p5_ASAP7_75t_L g556 ( .A(n_557), .B(n_558), .Y(n_556) );
OAI21x1_ASAP7_75t_L g558 ( .A1(n_559), .A2(n_564), .B(n_567), .Y(n_558) );
INVx2_ASAP7_75t_SL g562 ( .A(n_563), .Y(n_562) );
INVx2_ASAP7_75t_L g754 ( .A(n_569), .Y(n_754) );
OR2x2_ASAP7_75t_L g569 ( .A(n_570), .B(n_583), .Y(n_569) );
INVx2_ASAP7_75t_L g622 ( .A(n_570), .Y(n_622) );
INVx2_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
INVx1_ASAP7_75t_L g601 ( .A(n_571), .Y(n_601) );
OAI21xp5_ASAP7_75t_L g573 ( .A1(n_574), .A2(n_576), .B(n_578), .Y(n_573) );
INVx1_ASAP7_75t_L g602 ( .A(n_583), .Y(n_602) );
INVx3_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
OR2x6_ASAP7_75t_L g585 ( .A(n_586), .B(n_593), .Y(n_585) );
INVx2_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
AND2x2_ASAP7_75t_L g641 ( .A(n_587), .B(n_642), .Y(n_641) );
BUFx2_ASAP7_75t_L g771 ( .A(n_587), .Y(n_771) );
INVx1_ASAP7_75t_L g616 ( .A(n_588), .Y(n_616) );
AND2x2_ASAP7_75t_L g696 ( .A(n_588), .B(n_634), .Y(n_696) );
INVx2_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
AND2x2_ASAP7_75t_L g633 ( .A(n_589), .B(n_634), .Y(n_633) );
AOI21x1_ASAP7_75t_L g589 ( .A1(n_590), .A2(n_591), .B(n_592), .Y(n_589) );
INVx1_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
NOR2x1_ASAP7_75t_L g645 ( .A(n_594), .B(n_646), .Y(n_645) );
INVx2_ASAP7_75t_L g729 ( .A(n_594), .Y(n_729) );
NAND2xp5_ASAP7_75t_L g595 ( .A(n_596), .B(n_603), .Y(n_595) );
OAI22xp5_ASAP7_75t_L g636 ( .A1(n_596), .A2(n_637), .B1(n_640), .B2(n_644), .Y(n_636) );
INVx1_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
AOI22xp5_ASAP7_75t_L g654 ( .A1(n_597), .A2(n_617), .B1(n_649), .B2(n_655), .Y(n_654) );
AND2x2_ASAP7_75t_L g597 ( .A(n_598), .B(n_599), .Y(n_597) );
BUFx2_ASAP7_75t_SL g635 ( .A(n_598), .Y(n_635) );
AND2x4_ASAP7_75t_L g753 ( .A(n_598), .B(n_754), .Y(n_753) );
INVx1_ASAP7_75t_L g762 ( .A(n_598), .Y(n_762) );
INVx1_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
INVx1_ASAP7_75t_L g674 ( .A(n_600), .Y(n_674) );
OR2x2_ASAP7_75t_L g600 ( .A(n_601), .B(n_602), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g732 ( .A(n_601), .B(n_606), .Y(n_732) );
INVxp67_ASAP7_75t_L g761 ( .A(n_601), .Y(n_761) );
AND2x2_ASAP7_75t_L g766 ( .A(n_601), .B(n_632), .Y(n_766) );
OR2x2_ASAP7_75t_L g748 ( .A(n_602), .B(n_622), .Y(n_748) );
INVx1_ASAP7_75t_L g629 ( .A(n_603), .Y(n_629) );
NAND2xp5_ASAP7_75t_L g603 ( .A(n_604), .B(n_605), .Y(n_603) );
NAND2xp5_ASAP7_75t_L g686 ( .A(n_604), .B(n_687), .Y(n_686) );
AND2x2_ASAP7_75t_L g668 ( .A(n_605), .B(n_653), .Y(n_668) );
AND2x4_ASAP7_75t_L g605 ( .A(n_606), .B(n_607), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g621 ( .A(n_606), .B(n_622), .Y(n_621) );
INVx2_ASAP7_75t_L g652 ( .A(n_606), .Y(n_652) );
OR2x2_ASAP7_75t_L g747 ( .A(n_606), .B(n_748), .Y(n_747) );
OAI21xp33_ASAP7_75t_L g608 ( .A1(n_609), .A2(n_613), .B(n_618), .Y(n_608) );
INVx1_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
INVx2_ASAP7_75t_L g671 ( .A(n_610), .Y(n_671) );
OR2x2_ASAP7_75t_L g610 ( .A(n_611), .B(n_612), .Y(n_610) );
AND2x2_ASAP7_75t_L g665 ( .A(n_611), .B(n_662), .Y(n_665) );
INVx2_ASAP7_75t_L g789 ( .A(n_611), .Y(n_789) );
INVx2_ASAP7_75t_SL g613 ( .A(n_614), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g614 ( .A(n_615), .B(n_617), .Y(n_614) );
AND2x2_ASAP7_75t_L g718 ( .A(n_615), .B(n_661), .Y(n_718) );
AND2x2_ASAP7_75t_L g743 ( .A(n_615), .B(n_689), .Y(n_743) );
INVx1_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
INVx2_ASAP7_75t_L g646 ( .A(n_616), .Y(n_646) );
AND2x2_ASAP7_75t_L g673 ( .A(n_617), .B(n_627), .Y(n_673) );
NAND2xp5_ASAP7_75t_L g685 ( .A(n_617), .B(n_672), .Y(n_685) );
INVx1_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
OR2x2_ASAP7_75t_L g619 ( .A(n_620), .B(n_621), .Y(n_619) );
INVx1_ASAP7_75t_L g770 ( .A(n_620), .Y(n_770) );
OR2x2_ASAP7_75t_L g786 ( .A(n_620), .B(n_681), .Y(n_786) );
INVx1_ASAP7_75t_L g710 ( .A(n_622), .Y(n_710) );
NAND3xp33_ASAP7_75t_L g623 ( .A(n_624), .B(n_647), .C(n_669), .Y(n_623) );
AOI221xp5_ASAP7_75t_L g624 ( .A1(n_625), .A2(n_629), .B1(n_630), .B2(n_635), .C(n_636), .Y(n_624) );
INVx1_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
NAND2xp5_ASAP7_75t_L g626 ( .A(n_627), .B(n_628), .Y(n_626) );
AND2x2_ASAP7_75t_L g649 ( .A(n_628), .B(n_650), .Y(n_649) );
NAND2xp5_ASAP7_75t_L g777 ( .A(n_628), .B(n_693), .Y(n_777) );
AND2x2_ASAP7_75t_L g630 ( .A(n_631), .B(n_633), .Y(n_630) );
BUFx2_ASAP7_75t_L g631 ( .A(n_632), .Y(n_631) );
INVx3_ASAP7_75t_L g672 ( .A(n_632), .Y(n_672) );
AND3x1_ASAP7_75t_L g768 ( .A(n_632), .B(n_769), .C(n_770), .Y(n_768) );
AND2x2_ASAP7_75t_L g755 ( .A(n_633), .B(n_756), .Y(n_755) );
INVx2_ASAP7_75t_L g765 ( .A(n_633), .Y(n_765) );
INVxp67_ASAP7_75t_L g779 ( .A(n_635), .Y(n_779) );
OR2x2_ASAP7_75t_L g637 ( .A(n_638), .B(n_639), .Y(n_637) );
OR2x2_ASAP7_75t_L g734 ( .A(n_638), .B(n_658), .Y(n_734) );
INVx2_ASAP7_75t_L g769 ( .A(n_638), .Y(n_769) );
INVx1_ASAP7_75t_L g687 ( .A(n_639), .Y(n_687) );
INVx1_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
OAI21xp5_ASAP7_75t_L g688 ( .A1(n_641), .A2(n_689), .B(n_690), .Y(n_688) );
NAND2xp5_ASAP7_75t_L g788 ( .A(n_642), .B(n_789), .Y(n_788) );
INVx1_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
INVx1_ASAP7_75t_L g650 ( .A(n_643), .Y(n_650) );
OR2x2_ASAP7_75t_L g744 ( .A(n_643), .B(n_745), .Y(n_744) );
INVxp67_ASAP7_75t_SL g644 ( .A(n_645), .Y(n_644) );
INVx1_ASAP7_75t_L g704 ( .A(n_646), .Y(n_704) );
NAND2xp5_ASAP7_75t_L g783 ( .A(n_646), .B(n_703), .Y(n_783) );
AND3x1_ASAP7_75t_L g647 ( .A(n_648), .B(n_654), .C(n_659), .Y(n_647) );
NAND2xp5_ASAP7_75t_L g648 ( .A(n_649), .B(n_651), .Y(n_648) );
AND2x2_ASAP7_75t_L g698 ( .A(n_650), .B(n_689), .Y(n_698) );
AOI22xp5_ASAP7_75t_L g717 ( .A1(n_651), .A2(n_718), .B1(n_719), .B2(n_721), .Y(n_717) );
AND2x2_ASAP7_75t_L g651 ( .A(n_652), .B(n_653), .Y(n_651) );
OAI321xp33_ASAP7_75t_L g740 ( .A1(n_652), .A2(n_741), .A3(n_742), .B1(n_744), .B2(n_747), .C(n_749), .Y(n_740) );
AND2x2_ASAP7_75t_L g792 ( .A(n_652), .B(n_657), .Y(n_792) );
AND2x2_ASAP7_75t_L g690 ( .A(n_653), .B(n_656), .Y(n_690) );
INVx2_ASAP7_75t_L g699 ( .A(n_655), .Y(n_699) );
AND2x2_ASAP7_75t_L g708 ( .A(n_655), .B(n_709), .Y(n_708) );
AND2x4_ASAP7_75t_L g655 ( .A(n_656), .B(n_657), .Y(n_655) );
INVx2_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
OR2x2_ASAP7_75t_L g720 ( .A(n_658), .B(n_710), .Y(n_720) );
INVx2_ASAP7_75t_L g752 ( .A(n_658), .Y(n_752) );
OAI21xp33_ASAP7_75t_L g659 ( .A1(n_660), .A2(n_663), .B(n_668), .Y(n_659) );
HB1xp67_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
INVx1_ASAP7_75t_L g756 ( .A(n_662), .Y(n_756) );
NAND2xp5_ASAP7_75t_SL g663 ( .A(n_664), .B(n_666), .Y(n_663) );
INVx1_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
NAND2x1p5_ASAP7_75t_L g682 ( .A(n_665), .B(n_672), .Y(n_682) );
INVxp67_ASAP7_75t_L g666 ( .A(n_667), .Y(n_666) );
OAI21xp5_ASAP7_75t_L g669 ( .A1(n_670), .A2(n_673), .B(n_674), .Y(n_669) );
AND2x2_ASAP7_75t_L g670 ( .A(n_671), .B(n_672), .Y(n_670) );
NAND2xp5_ASAP7_75t_L g722 ( .A(n_672), .B(n_696), .Y(n_722) );
NAND2xp5_ASAP7_75t_L g736 ( .A(n_672), .B(n_737), .Y(n_736) );
AND2x2_ASAP7_75t_L g773 ( .A(n_672), .B(n_774), .Y(n_773) );
INVx1_ASAP7_75t_L g741 ( .A(n_674), .Y(n_741) );
NOR2xp67_ASAP7_75t_L g675 ( .A(n_676), .B(n_738), .Y(n_675) );
NAND3xp33_ASAP7_75t_L g676 ( .A(n_677), .B(n_700), .C(n_723), .Y(n_676) );
NOR2xp33_ASAP7_75t_L g677 ( .A(n_678), .B(n_691), .Y(n_677) );
OAI221xp5_ASAP7_75t_L g678 ( .A1(n_679), .A2(n_682), .B1(n_683), .B2(n_686), .C(n_688), .Y(n_678) );
OR2x2_ASAP7_75t_L g679 ( .A(n_680), .B(n_681), .Y(n_679) );
OR2x2_ASAP7_75t_L g731 ( .A(n_680), .B(n_732), .Y(n_731) );
INVx1_ASAP7_75t_L g683 ( .A(n_684), .Y(n_683) );
INVx1_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
AOI21xp33_ASAP7_75t_SL g691 ( .A1(n_692), .A2(n_697), .B(n_699), .Y(n_691) );
NAND2xp5_ASAP7_75t_L g692 ( .A(n_693), .B(n_694), .Y(n_692) );
INVx1_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
INVx2_ASAP7_75t_L g695 ( .A(n_696), .Y(n_695) );
AND2x2_ASAP7_75t_L g728 ( .A(n_696), .B(n_729), .Y(n_728) );
OAI21xp33_ASAP7_75t_SL g711 ( .A1(n_697), .A2(n_712), .B(n_717), .Y(n_711) );
INVx2_ASAP7_75t_SL g697 ( .A(n_698), .Y(n_697) );
O2A1O1Ixp33_ASAP7_75t_L g700 ( .A1(n_701), .A2(n_705), .B(n_708), .C(n_711), .Y(n_700) );
INVx2_ASAP7_75t_SL g701 ( .A(n_702), .Y(n_701) );
NAND2xp5_ASAP7_75t_L g776 ( .A(n_702), .B(n_777), .Y(n_776) );
NAND2x1_ASAP7_75t_L g702 ( .A(n_703), .B(n_704), .Y(n_702) );
INVx1_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
INVx1_ASAP7_75t_L g706 ( .A(n_707), .Y(n_706) );
INVx1_ASAP7_75t_L g709 ( .A(n_710), .Y(n_709) );
NAND2xp5_ASAP7_75t_L g751 ( .A(n_710), .B(n_752), .Y(n_751) );
INVxp67_ASAP7_75t_L g712 ( .A(n_713), .Y(n_712) );
NAND2xp5_ASAP7_75t_SL g772 ( .A(n_713), .B(n_773), .Y(n_772) );
INVx2_ASAP7_75t_L g713 ( .A(n_714), .Y(n_713) );
NAND2xp5_ASAP7_75t_L g714 ( .A(n_715), .B(n_716), .Y(n_714) );
INVx2_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
INVx1_ASAP7_75t_L g721 ( .A(n_722), .Y(n_721) );
AOI22xp5_ASAP7_75t_L g723 ( .A1(n_724), .A2(n_730), .B1(n_733), .B2(n_735), .Y(n_723) );
INVx1_ASAP7_75t_L g725 ( .A(n_726), .Y(n_725) );
INVx1_ASAP7_75t_L g727 ( .A(n_728), .Y(n_727) );
INVx1_ASAP7_75t_L g730 ( .A(n_731), .Y(n_730) );
HB1xp67_ASAP7_75t_L g795 ( .A(n_732), .Y(n_795) );
INVx1_ASAP7_75t_L g733 ( .A(n_734), .Y(n_733) );
INVx1_ASAP7_75t_L g735 ( .A(n_736), .Y(n_735) );
NAND3xp33_ASAP7_75t_L g738 ( .A(n_739), .B(n_775), .C(n_790), .Y(n_738) );
NOR2xp33_ASAP7_75t_L g739 ( .A(n_740), .B(n_757), .Y(n_739) );
INVx2_ASAP7_75t_L g742 ( .A(n_743), .Y(n_742) );
INVx2_ASAP7_75t_SL g745 ( .A(n_746), .Y(n_745) );
OAI21xp33_ASAP7_75t_L g749 ( .A1(n_750), .A2(n_753), .B(n_755), .Y(n_749) );
INVx1_ASAP7_75t_L g750 ( .A(n_751), .Y(n_750) );
NAND3xp33_ASAP7_75t_L g757 ( .A(n_758), .B(n_763), .C(n_772), .Y(n_757) );
INVx1_ASAP7_75t_L g759 ( .A(n_760), .Y(n_759) );
OR2x2_ASAP7_75t_L g760 ( .A(n_761), .B(n_762), .Y(n_760) );
AOI32xp33_ASAP7_75t_L g763 ( .A1(n_764), .A2(n_766), .A3(n_767), .B1(n_768), .B2(n_771), .Y(n_763) );
INVx3_ASAP7_75t_L g764 ( .A(n_765), .Y(n_764) );
AND2x2_ASAP7_75t_L g791 ( .A(n_766), .B(n_792), .Y(n_791) );
AOI21xp5_ASAP7_75t_L g775 ( .A1(n_776), .A2(n_778), .B(n_780), .Y(n_775) );
INVx1_ASAP7_75t_L g780 ( .A(n_781), .Y(n_780) );
AOI22x1_ASAP7_75t_L g781 ( .A1(n_782), .A2(n_784), .B1(n_785), .B2(n_787), .Y(n_781) );
INVx1_ASAP7_75t_L g782 ( .A(n_783), .Y(n_782) );
AOI21xp33_ASAP7_75t_L g794 ( .A1(n_783), .A2(n_795), .B(n_796), .Y(n_794) );
INVx2_ASAP7_75t_L g785 ( .A(n_786), .Y(n_785) );
INVx1_ASAP7_75t_L g787 ( .A(n_788), .Y(n_787) );
AOI21xp5_ASAP7_75t_L g790 ( .A1(n_791), .A2(n_793), .B(n_794), .Y(n_790) );
INVx1_ASAP7_75t_L g796 ( .A(n_797), .Y(n_796) );
INVx8_ASAP7_75t_L g798 ( .A(n_799), .Y(n_798) );
BUFx12f_ASAP7_75t_L g799 ( .A(n_800), .Y(n_799) );
OAI21xp33_ASAP7_75t_L g803 ( .A1(n_804), .A2(n_811), .B(n_833), .Y(n_803) );
CKINVDCx20_ASAP7_75t_R g804 ( .A(n_805), .Y(n_804) );
CKINVDCx20_ASAP7_75t_R g805 ( .A(n_806), .Y(n_805) );
INVx4_ASAP7_75t_SL g806 ( .A(n_807), .Y(n_806) );
BUFx3_ASAP7_75t_L g807 ( .A(n_808), .Y(n_807) );
OR2x4_ASAP7_75t_L g839 ( .A(n_809), .B(n_840), .Y(n_839) );
BUFx2_ASAP7_75t_L g809 ( .A(n_810), .Y(n_809) );
AOI21xp5_ASAP7_75t_L g811 ( .A1(n_812), .A2(n_825), .B(n_826), .Y(n_811) );
AND2x2_ASAP7_75t_L g812 ( .A(n_813), .B(n_820), .Y(n_812) );
BUFx12f_ASAP7_75t_L g813 ( .A(n_814), .Y(n_813) );
INVx4_ASAP7_75t_L g814 ( .A(n_815), .Y(n_814) );
INVx3_ASAP7_75t_L g828 ( .A(n_815), .Y(n_828) );
CKINVDCx8_ASAP7_75t_R g837 ( .A(n_815), .Y(n_837) );
AND2x6_ASAP7_75t_SL g815 ( .A(n_816), .B(n_819), .Y(n_815) );
INVx1_ASAP7_75t_L g817 ( .A(n_818), .Y(n_817) );
OAI31xp33_ASAP7_75t_SL g826 ( .A1(n_820), .A2(n_825), .A3(n_827), .B(n_829), .Y(n_826) );
CKINVDCx5p33_ASAP7_75t_R g822 ( .A(n_823), .Y(n_822) );
INVx2_ASAP7_75t_L g827 ( .A(n_828), .Y(n_827) );
BUFx2_ASAP7_75t_SL g831 ( .A(n_828), .Y(n_831) );
INVxp67_ASAP7_75t_L g829 ( .A(n_830), .Y(n_829) );
NOR2xp33_ASAP7_75t_L g830 ( .A(n_831), .B(n_832), .Y(n_830) );
INVx3_ASAP7_75t_L g836 ( .A(n_837), .Y(n_836) );
BUFx3_ASAP7_75t_L g838 ( .A(n_839), .Y(n_838) );
endmodule