module fake_jpeg_1395_n_702 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_702);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_702;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_696;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_657;
wire n_27;
wire n_664;
wire n_365;
wire n_179;
wire n_620;
wire n_686;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_678;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_699;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_643;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_647;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_641;
wire n_701;
wire n_48;
wire n_465;
wire n_638;
wire n_200;
wire n_582;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_637;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_672;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_606;
wire n_496;
wire n_166;
wire n_688;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_646;
wire n_319;
wire n_689;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_663;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_658;
wire n_698;
wire n_195;
wire n_450;
wire n_557;
wire n_681;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_666;
wire n_639;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_645;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_694;
wire n_692;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_667;
wire n_92;
wire n_332;
wire n_640;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_653;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_668;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_682;
wire n_305;
wire n_161;
wire n_441;
wire n_697;
wire n_555;
wire n_342;
wire n_642;
wire n_101;
wire n_226;
wire n_509;
wire n_644;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_656;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_649;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_679;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_691;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_615;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_662;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_676;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_648;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_670;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_683;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_690;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_650;
wire n_218;
wire n_63;
wire n_652;
wire n_599;
wire n_239;
wire n_693;
wire n_674;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_378;
wire n_419;
wire n_133;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_655;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_684;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_680;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_695;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_659;
wire n_125;
wire n_661;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_687;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_673;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_665;
wire n_72;
wire n_512;
wire n_654;
wire n_445;
wire n_443;
wire n_677;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_700;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_671;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_669;
wire n_524;
wire n_402;
wire n_563;
wire n_685;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_660;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_651;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_675;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx2_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

INVx6_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

CKINVDCx5p33_ASAP7_75t_R g22 ( 
.A(n_12),
.Y(n_22)
);

INVx2_ASAP7_75t_SL g23 ( 
.A(n_9),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

BUFx8_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

BUFx4f_ASAP7_75t_SL g26 ( 
.A(n_17),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_10),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

BUFx16f_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_9),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_2),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_11),
.B(n_16),
.Y(n_34)
);

BUFx6f_ASAP7_75t_SL g35 ( 
.A(n_4),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_19),
.Y(n_36)
);

INVx6_ASAP7_75t_SL g37 ( 
.A(n_16),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_11),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_18),
.B(n_9),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_18),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_7),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_11),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_12),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_1),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_13),
.Y(n_46)
);

BUFx12_ASAP7_75t_L g47 ( 
.A(n_17),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_13),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_7),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_0),
.Y(n_50)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_13),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_4),
.Y(n_52)
);

CKINVDCx5p33_ASAP7_75t_R g53 ( 
.A(n_19),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_8),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_13),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_19),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_1),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_14),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_3),
.Y(n_59)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_51),
.Y(n_60)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_60),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_34),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_61),
.B(n_68),
.Y(n_140)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_51),
.Y(n_62)
);

INVx3_ASAP7_75t_L g157 ( 
.A(n_62),
.Y(n_157)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_36),
.Y(n_63)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_63),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_44),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_64),
.Y(n_141)
);

BUFx5_ASAP7_75t_L g65 ( 
.A(n_37),
.Y(n_65)
);

INVx4_ASAP7_75t_L g137 ( 
.A(n_65),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_44),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_66),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_34),
.B(n_17),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_67),
.B(n_127),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_39),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_36),
.Y(n_69)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_69),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_44),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_70),
.Y(n_163)
);

BUFx12_ASAP7_75t_L g71 ( 
.A(n_37),
.Y(n_71)
);

BUFx4f_ASAP7_75t_SL g151 ( 
.A(n_71),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_44),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g191 ( 
.A(n_72),
.Y(n_191)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_43),
.Y(n_73)
);

BUFx2_ASAP7_75t_L g205 ( 
.A(n_73),
.Y(n_205)
);

CKINVDCx16_ASAP7_75t_R g74 ( 
.A(n_26),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_74),
.B(n_77),
.Y(n_153)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_55),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g192 ( 
.A(n_75),
.Y(n_192)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_56),
.Y(n_76)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_76),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_39),
.Y(n_77)
);

INVx8_ASAP7_75t_L g78 ( 
.A(n_37),
.Y(n_78)
);

BUFx2_ASAP7_75t_L g218 ( 
.A(n_78),
.Y(n_218)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_20),
.Y(n_79)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_79),
.Y(n_145)
);

BUFx5_ASAP7_75t_L g80 ( 
.A(n_25),
.Y(n_80)
);

INVx4_ASAP7_75t_L g142 ( 
.A(n_80),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_55),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g197 ( 
.A(n_81),
.Y(n_197)
);

BUFx3_ASAP7_75t_L g82 ( 
.A(n_43),
.Y(n_82)
);

BUFx3_ASAP7_75t_L g183 ( 
.A(n_82),
.Y(n_183)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_20),
.Y(n_83)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_83),
.Y(n_147)
);

INVx8_ASAP7_75t_L g84 ( 
.A(n_30),
.Y(n_84)
);

INVx5_ASAP7_75t_L g195 ( 
.A(n_84),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_30),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_85),
.B(n_86),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_41),
.B(n_15),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_56),
.Y(n_87)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_87),
.Y(n_217)
);

BUFx8_ASAP7_75t_L g88 ( 
.A(n_25),
.Y(n_88)
);

INVx13_ASAP7_75t_L g139 ( 
.A(n_88),
.Y(n_139)
);

BUFx12f_ASAP7_75t_L g89 ( 
.A(n_25),
.Y(n_89)
);

INVx5_ASAP7_75t_L g199 ( 
.A(n_89),
.Y(n_199)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_55),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g207 ( 
.A(n_90),
.Y(n_207)
);

INVx8_ASAP7_75t_L g91 ( 
.A(n_30),
.Y(n_91)
);

INVx5_ASAP7_75t_L g219 ( 
.A(n_91),
.Y(n_219)
);

INVx8_ASAP7_75t_L g92 ( 
.A(n_30),
.Y(n_92)
);

INVx6_ASAP7_75t_L g148 ( 
.A(n_92),
.Y(n_148)
);

BUFx16f_ASAP7_75t_L g93 ( 
.A(n_25),
.Y(n_93)
);

BUFx8_ASAP7_75t_L g181 ( 
.A(n_93),
.Y(n_181)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_55),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g215 ( 
.A(n_94),
.Y(n_215)
);

INVx6_ASAP7_75t_SL g95 ( 
.A(n_25),
.Y(n_95)
);

INVx2_ASAP7_75t_R g164 ( 
.A(n_95),
.Y(n_164)
);

BUFx12f_ASAP7_75t_L g96 ( 
.A(n_47),
.Y(n_96)
);

INVx8_ASAP7_75t_L g169 ( 
.A(n_96),
.Y(n_169)
);

OR2x2_ASAP7_75t_L g97 ( 
.A(n_53),
.B(n_29),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_97),
.B(n_99),
.Y(n_190)
);

BUFx5_ASAP7_75t_L g98 ( 
.A(n_26),
.Y(n_98)
);

INVx4_ASAP7_75t_L g161 ( 
.A(n_98),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_40),
.Y(n_99)
);

BUFx3_ASAP7_75t_L g100 ( 
.A(n_43),
.Y(n_100)
);

BUFx3_ASAP7_75t_L g206 ( 
.A(n_100),
.Y(n_206)
);

BUFx3_ASAP7_75t_L g101 ( 
.A(n_50),
.Y(n_101)
);

INVx4_ASAP7_75t_L g162 ( 
.A(n_101),
.Y(n_162)
);

INVx2_ASAP7_75t_SL g102 ( 
.A(n_23),
.Y(n_102)
);

INVx1_ASAP7_75t_SL g135 ( 
.A(n_102),
.Y(n_135)
);

BUFx3_ASAP7_75t_L g103 ( 
.A(n_50),
.Y(n_103)
);

INVx4_ASAP7_75t_L g174 ( 
.A(n_103),
.Y(n_174)
);

BUFx3_ASAP7_75t_L g104 ( 
.A(n_50),
.Y(n_104)
);

INVx4_ASAP7_75t_L g176 ( 
.A(n_104),
.Y(n_176)
);

BUFx3_ASAP7_75t_L g105 ( 
.A(n_51),
.Y(n_105)
);

INVx4_ASAP7_75t_L g177 ( 
.A(n_105),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_40),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_106),
.B(n_110),
.Y(n_209)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_24),
.Y(n_107)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_107),
.Y(n_220)
);

BUFx12f_ASAP7_75t_L g108 ( 
.A(n_47),
.Y(n_108)
);

INVx4_ASAP7_75t_L g204 ( 
.A(n_108),
.Y(n_204)
);

BUFx12f_ASAP7_75t_L g109 ( 
.A(n_47),
.Y(n_109)
);

INVx4_ASAP7_75t_L g211 ( 
.A(n_109),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_40),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_53),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_111),
.B(n_112),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_41),
.B(n_15),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_21),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g227 ( 
.A(n_113),
.Y(n_227)
);

INVx8_ASAP7_75t_L g114 ( 
.A(n_45),
.Y(n_114)
);

INVx6_ASAP7_75t_L g189 ( 
.A(n_114),
.Y(n_189)
);

AND2x2_ASAP7_75t_L g115 ( 
.A(n_53),
.B(n_15),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g149 ( 
.A(n_115),
.B(n_22),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_21),
.Y(n_116)
);

INVx6_ASAP7_75t_L g160 ( 
.A(n_116),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_21),
.Y(n_117)
);

INVx6_ASAP7_75t_L g208 ( 
.A(n_117),
.Y(n_208)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_45),
.Y(n_118)
);

INVx6_ASAP7_75t_L g221 ( 
.A(n_118),
.Y(n_221)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_45),
.Y(n_119)
);

INVx6_ASAP7_75t_L g224 ( 
.A(n_119),
.Y(n_224)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_24),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_120),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_45),
.Y(n_121)
);

BUFx12f_ASAP7_75t_L g133 ( 
.A(n_121),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_45),
.Y(n_122)
);

BUFx12f_ASAP7_75t_L g156 ( 
.A(n_122),
.Y(n_156)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_54),
.Y(n_123)
);

INVx3_ASAP7_75t_L g158 ( 
.A(n_123),
.Y(n_158)
);

INVx8_ASAP7_75t_L g124 ( 
.A(n_54),
.Y(n_124)
);

INVx3_ASAP7_75t_L g188 ( 
.A(n_124),
.Y(n_188)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_54),
.Y(n_125)
);

BUFx12f_ASAP7_75t_L g168 ( 
.A(n_125),
.Y(n_168)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_38),
.Y(n_126)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_126),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_26),
.B(n_16),
.Y(n_127)
);

BUFx4f_ASAP7_75t_L g128 ( 
.A(n_23),
.Y(n_128)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_128),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_54),
.Y(n_129)
);

BUFx12f_ASAP7_75t_L g171 ( 
.A(n_129),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_22),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_130),
.B(n_28),
.Y(n_202)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_27),
.Y(n_131)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_131),
.Y(n_172)
);

BUFx3_ASAP7_75t_L g132 ( 
.A(n_38),
.Y(n_132)
);

INVx4_ASAP7_75t_L g225 ( 
.A(n_132),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_93),
.Y(n_134)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_134),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_115),
.A2(n_54),
.B1(n_57),
.B2(n_46),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_144),
.A2(n_201),
.B1(n_149),
.B2(n_152),
.Y(n_243)
);

INVx11_ASAP7_75t_L g146 ( 
.A(n_88),
.Y(n_146)
);

INVx4_ASAP7_75t_L g232 ( 
.A(n_146),
.Y(n_232)
);

AND2x2_ASAP7_75t_L g267 ( 
.A(n_149),
.B(n_33),
.Y(n_267)
);

AND2x2_ASAP7_75t_L g152 ( 
.A(n_97),
.B(n_22),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g238 ( 
.A(n_152),
.B(n_155),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_113),
.Y(n_155)
);

INVx11_ASAP7_75t_L g165 ( 
.A(n_88),
.Y(n_165)
);

CKINVDCx16_ASAP7_75t_R g248 ( 
.A(n_165),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_116),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_SL g250 ( 
.A(n_167),
.B(n_185),
.Y(n_250)
);

INVx11_ASAP7_75t_L g170 ( 
.A(n_89),
.Y(n_170)
);

INVx1_ASAP7_75t_SL g268 ( 
.A(n_170),
.Y(n_268)
);

CKINVDCx14_ASAP7_75t_R g178 ( 
.A(n_102),
.Y(n_178)
);

NAND2xp33_ASAP7_75t_SL g231 ( 
.A(n_178),
.B(n_35),
.Y(n_231)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_132),
.Y(n_179)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_179),
.Y(n_233)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_128),
.Y(n_180)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_180),
.Y(n_244)
);

AOI22xp33_ASAP7_75t_L g182 ( 
.A1(n_64),
.A2(n_23),
.B1(n_26),
.B2(n_35),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g273 ( 
.A1(n_182),
.A2(n_187),
.B1(n_72),
.B2(n_81),
.Y(n_273)
);

AND2x2_ASAP7_75t_L g185 ( 
.A(n_123),
.B(n_23),
.Y(n_185)
);

INVx11_ASAP7_75t_L g186 ( 
.A(n_89),
.Y(n_186)
);

INVx1_ASAP7_75t_SL g293 ( 
.A(n_186),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_117),
.A2(n_35),
.B1(n_26),
.B2(n_48),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_128),
.B(n_58),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_193),
.B(n_202),
.Y(n_275)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_60),
.Y(n_194)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_194),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_75),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_SL g283 ( 
.A(n_196),
.B(n_228),
.Y(n_283)
);

INVx3_ASAP7_75t_L g198 ( 
.A(n_84),
.Y(n_198)
);

INVx4_ASAP7_75t_SL g271 ( 
.A(n_198),
.Y(n_271)
);

INVx3_ASAP7_75t_L g200 ( 
.A(n_91),
.Y(n_200)
);

INVx4_ASAP7_75t_SL g284 ( 
.A(n_200),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_66),
.A2(n_28),
.B1(n_57),
.B2(n_49),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_62),
.B(n_27),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g287 ( 
.A(n_203),
.B(n_42),
.Y(n_287)
);

INVx3_ASAP7_75t_L g210 ( 
.A(n_92),
.Y(n_210)
);

INVx2_ASAP7_75t_SL g278 ( 
.A(n_210),
.Y(n_278)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_105),
.Y(n_212)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_212),
.Y(n_257)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_129),
.Y(n_213)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_213),
.Y(n_269)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_118),
.Y(n_214)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_214),
.Y(n_290)
);

INVx3_ASAP7_75t_L g216 ( 
.A(n_78),
.Y(n_216)
);

HB1xp67_ASAP7_75t_L g305 ( 
.A(n_216),
.Y(n_305)
);

BUFx12f_ASAP7_75t_L g222 ( 
.A(n_71),
.Y(n_222)
);

INVx5_ASAP7_75t_L g294 ( 
.A(n_222),
.Y(n_294)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_119),
.Y(n_223)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_223),
.Y(n_295)
);

AND2x2_ASAP7_75t_L g228 ( 
.A(n_114),
.B(n_29),
.Y(n_228)
);

INVx3_ASAP7_75t_L g229 ( 
.A(n_124),
.Y(n_229)
);

INVx3_ASAP7_75t_L g236 ( 
.A(n_229),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_138),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g341 ( 
.A(n_230),
.B(n_239),
.Y(n_341)
);

AND2x2_ASAP7_75t_L g319 ( 
.A(n_231),
.B(n_287),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_153),
.B(n_73),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_SL g349 ( 
.A(n_234),
.B(n_247),
.Y(n_349)
);

CKINVDCx12_ASAP7_75t_R g235 ( 
.A(n_181),
.Y(n_235)
);

INVx4_ASAP7_75t_SL g345 ( 
.A(n_235),
.Y(n_345)
);

AOI22x1_ASAP7_75t_SL g237 ( 
.A1(n_184),
.A2(n_125),
.B1(n_122),
.B2(n_121),
.Y(n_237)
);

OAI22xp33_ASAP7_75t_SL g327 ( 
.A1(n_237),
.A2(n_162),
.B1(n_176),
.B2(n_174),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_138),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_166),
.Y(n_240)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_240),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_193),
.B(n_48),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_241),
.B(n_266),
.Y(n_316)
);

OA22x2_ASAP7_75t_L g242 ( 
.A1(n_182),
.A2(n_82),
.B1(n_104),
.B2(n_103),
.Y(n_242)
);

AO22x2_ASAP7_75t_L g329 ( 
.A1(n_242),
.A2(n_261),
.B1(n_288),
.B2(n_249),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_L g352 ( 
.A1(n_243),
.A2(n_276),
.B1(n_300),
.B2(n_304),
.Y(n_352)
);

BUFx6f_ASAP7_75t_L g246 ( 
.A(n_141),
.Y(n_246)
);

BUFx6f_ASAP7_75t_L g320 ( 
.A(n_246),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_178),
.Y(n_247)
);

CKINVDCx9p33_ASAP7_75t_R g249 ( 
.A(n_181),
.Y(n_249)
);

BUFx5_ASAP7_75t_L g318 ( 
.A(n_249),
.Y(n_318)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_173),
.Y(n_251)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_251),
.Y(n_338)
);

INVx3_ASAP7_75t_L g252 ( 
.A(n_148),
.Y(n_252)
);

INVx4_ASAP7_75t_L g321 ( 
.A(n_252),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_209),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_SL g365 ( 
.A(n_253),
.B(n_254),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_153),
.B(n_140),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_220),
.B(n_101),
.C(n_100),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g368 ( 
.A(n_255),
.B(n_211),
.C(n_204),
.Y(n_368)
);

BUFx12f_ASAP7_75t_L g256 ( 
.A(n_169),
.Y(n_256)
);

INVx5_ASAP7_75t_L g325 ( 
.A(n_256),
.Y(n_325)
);

BUFx3_ASAP7_75t_L g258 ( 
.A(n_199),
.Y(n_258)
);

BUFx3_ASAP7_75t_L g375 ( 
.A(n_258),
.Y(n_375)
);

INVx6_ASAP7_75t_L g259 ( 
.A(n_141),
.Y(n_259)
);

BUFx6f_ASAP7_75t_L g357 ( 
.A(n_259),
.Y(n_357)
);

INVx3_ASAP7_75t_L g260 ( 
.A(n_195),
.Y(n_260)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_260),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_208),
.A2(n_70),
.B1(n_94),
.B2(n_90),
.Y(n_261)
);

AOI22xp33_ASAP7_75t_SL g262 ( 
.A1(n_135),
.A2(n_31),
.B1(n_52),
.B2(n_58),
.Y(n_262)
);

AOI22xp33_ASAP7_75t_SL g326 ( 
.A1(n_262),
.A2(n_263),
.B1(n_273),
.B2(n_303),
.Y(n_326)
);

AOI22xp33_ASAP7_75t_SL g263 ( 
.A1(n_185),
.A2(n_31),
.B1(n_52),
.B2(n_59),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_140),
.B(n_108),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_SL g371 ( 
.A(n_264),
.B(n_265),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_154),
.B(n_108),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_154),
.B(n_33),
.Y(n_266)
);

XNOR2x1_ASAP7_75t_L g333 ( 
.A(n_267),
.B(n_311),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_226),
.B(n_96),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_270),
.B(n_272),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_226),
.B(n_175),
.Y(n_272)
);

INVx8_ASAP7_75t_L g274 ( 
.A(n_189),
.Y(n_274)
);

INVx2_ASAP7_75t_L g332 ( 
.A(n_274),
.Y(n_332)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_145),
.A2(n_32),
.B1(n_59),
.B2(n_49),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_217),
.Y(n_277)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_277),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_190),
.B(n_96),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_279),
.B(n_280),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_190),
.B(n_109),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_172),
.B(n_46),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_281),
.B(n_285),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_209),
.B(n_109),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g350 ( 
.A(n_282),
.B(n_297),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_147),
.B(n_42),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_159),
.Y(n_286)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_286),
.Y(n_358)
);

OAI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_150),
.A2(n_32),
.B1(n_47),
.B2(n_98),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_228),
.B(n_0),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_289),
.B(n_161),
.Y(n_322)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_218),
.Y(n_291)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_291),
.Y(n_359)
);

BUFx6f_ASAP7_75t_L g292 ( 
.A(n_143),
.Y(n_292)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_292),
.Y(n_337)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_160),
.Y(n_296)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_296),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_218),
.Y(n_297)
);

INVx6_ASAP7_75t_L g298 ( 
.A(n_143),
.Y(n_298)
);

INVx2_ASAP7_75t_L g356 ( 
.A(n_298),
.Y(n_356)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_158),
.Y(n_299)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_299),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_L g300 ( 
.A1(n_160),
.A2(n_47),
.B1(n_65),
.B2(n_71),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_219),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_301),
.Y(n_336)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_192),
.Y(n_302)
);

INVx2_ASAP7_75t_L g362 ( 
.A(n_302),
.Y(n_362)
);

AOI22xp33_ASAP7_75t_SL g303 ( 
.A1(n_142),
.A2(n_80),
.B1(n_1),
.B2(n_3),
.Y(n_303)
);

AOI22xp33_ASAP7_75t_SL g304 ( 
.A1(n_205),
.A2(n_0),
.B1(n_3),
.B2(n_4),
.Y(n_304)
);

OAI22xp33_ASAP7_75t_SL g307 ( 
.A1(n_227),
.A2(n_0),
.B1(n_3),
.B2(n_4),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_SL g370 ( 
.A1(n_307),
.A2(n_312),
.B1(n_5),
.B2(n_6),
.Y(n_370)
);

BUFx6f_ASAP7_75t_L g308 ( 
.A(n_163),
.Y(n_308)
);

INVx2_ASAP7_75t_L g364 ( 
.A(n_308),
.Y(n_364)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_192),
.Y(n_309)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_309),
.Y(n_363)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_188),
.Y(n_310)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_310),
.Y(n_328)
);

AND2x2_ASAP7_75t_L g311 ( 
.A(n_136),
.B(n_14),
.Y(n_311)
);

AOI22xp33_ASAP7_75t_SL g312 ( 
.A1(n_205),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_275),
.B(n_151),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g396 ( 
.A(n_313),
.B(n_368),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_SL g381 ( 
.A(n_322),
.B(n_351),
.Y(n_381)
);

AND2x2_ASAP7_75t_L g323 ( 
.A(n_231),
.B(n_164),
.Y(n_323)
);

INVx1_ASAP7_75t_SL g414 ( 
.A(n_323),
.Y(n_414)
);

AOI22xp5_ASAP7_75t_SL g402 ( 
.A1(n_327),
.A2(n_355),
.B1(n_366),
.B2(n_248),
.Y(n_402)
);

AND2x2_ASAP7_75t_L g380 ( 
.A(n_329),
.B(n_348),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_241),
.B(n_225),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_330),
.B(n_331),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_285),
.B(n_157),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_281),
.B(n_151),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_334),
.B(n_335),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_289),
.B(n_227),
.Y(n_335)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_244),
.Y(n_339)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_339),
.Y(n_376)
);

AND2x2_ASAP7_75t_SL g342 ( 
.A(n_311),
.B(n_164),
.Y(n_342)
);

CKINVDCx14_ASAP7_75t_R g395 ( 
.A(n_342),
.Y(n_395)
);

AOI22xp33_ASAP7_75t_L g346 ( 
.A1(n_242),
.A2(n_191),
.B1(n_163),
.B2(n_215),
.Y(n_346)
);

OAI22xp33_ASAP7_75t_SL g421 ( 
.A1(n_346),
.A2(n_246),
.B1(n_292),
.B2(n_308),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_311),
.B(n_191),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_347),
.B(n_361),
.Y(n_397)
);

AND2x2_ASAP7_75t_L g348 ( 
.A(n_243),
.B(n_137),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g351 ( 
.A(n_306),
.Y(n_351)
);

CKINVDCx20_ASAP7_75t_R g354 ( 
.A(n_306),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_SL g389 ( 
.A(n_354),
.B(n_373),
.Y(n_389)
);

OAI22xp33_ASAP7_75t_SL g355 ( 
.A1(n_237),
.A2(n_197),
.B1(n_207),
.B2(n_215),
.Y(n_355)
);

AOI21xp5_ASAP7_75t_L g360 ( 
.A1(n_250),
.A2(n_139),
.B(n_177),
.Y(n_360)
);

AOI21xp5_ASAP7_75t_L g406 ( 
.A1(n_360),
.A2(n_372),
.B(n_232),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_283),
.B(n_197),
.Y(n_361)
);

OAI22xp33_ASAP7_75t_SL g366 ( 
.A1(n_276),
.A2(n_207),
.B1(n_183),
.B2(n_206),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_269),
.Y(n_367)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_367),
.Y(n_384)
);

OAI21xp5_ASAP7_75t_L g369 ( 
.A1(n_238),
.A2(n_139),
.B(n_169),
.Y(n_369)
);

AOI21xp5_ASAP7_75t_SL g392 ( 
.A1(n_369),
.A2(n_310),
.B(n_242),
.Y(n_392)
);

INVxp67_ASAP7_75t_L g404 ( 
.A(n_370),
.Y(n_404)
);

AOI21xp5_ASAP7_75t_L g372 ( 
.A1(n_255),
.A2(n_224),
.B(n_221),
.Y(n_372)
);

CKINVDCx20_ASAP7_75t_R g373 ( 
.A(n_305),
.Y(n_373)
);

CKINVDCx20_ASAP7_75t_R g374 ( 
.A(n_294),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_SL g415 ( 
.A(n_374),
.B(n_232),
.Y(n_415)
);

OAI21xp5_ASAP7_75t_L g378 ( 
.A1(n_323),
.A2(n_267),
.B(n_266),
.Y(n_378)
);

OAI21xp5_ASAP7_75t_SL g446 ( 
.A1(n_378),
.A2(n_392),
.B(n_406),
.Y(n_446)
);

CKINVDCx20_ASAP7_75t_R g379 ( 
.A(n_341),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_L g443 ( 
.A(n_379),
.B(n_394),
.Y(n_443)
);

INVx2_ASAP7_75t_L g382 ( 
.A(n_362),
.Y(n_382)
);

INVxp67_ASAP7_75t_L g456 ( 
.A(n_382),
.Y(n_456)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_328),
.Y(n_385)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_385),
.Y(n_434)
);

INVx2_ASAP7_75t_L g386 ( 
.A(n_362),
.Y(n_386)
);

INVxp67_ASAP7_75t_L g466 ( 
.A(n_386),
.Y(n_466)
);

INVx13_ASAP7_75t_L g387 ( 
.A(n_345),
.Y(n_387)
);

INVxp33_ASAP7_75t_L g458 ( 
.A(n_387),
.Y(n_458)
);

AOI22xp5_ASAP7_75t_L g388 ( 
.A1(n_352),
.A2(n_261),
.B1(n_288),
.B2(n_267),
.Y(n_388)
);

OAI22xp5_ASAP7_75t_SL g452 ( 
.A1(n_388),
.A2(n_329),
.B1(n_332),
.B2(n_356),
.Y(n_452)
);

NOR2xp33_ASAP7_75t_L g390 ( 
.A(n_349),
.B(n_299),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_SL g432 ( 
.A(n_390),
.B(n_393),
.Y(n_432)
);

BUFx6f_ASAP7_75t_L g391 ( 
.A(n_320),
.Y(n_391)
);

BUFx2_ASAP7_75t_L g436 ( 
.A(n_391),
.Y(n_436)
);

NOR2xp33_ASAP7_75t_L g393 ( 
.A(n_365),
.B(n_371),
.Y(n_393)
);

CKINVDCx20_ASAP7_75t_R g394 ( 
.A(n_350),
.Y(n_394)
);

CKINVDCx20_ASAP7_75t_R g398 ( 
.A(n_336),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_398),
.B(n_339),
.Y(n_467)
);

AOI22xp33_ASAP7_75t_L g399 ( 
.A1(n_331),
.A2(n_252),
.B1(n_242),
.B2(n_278),
.Y(n_399)
);

AOI22xp33_ASAP7_75t_L g453 ( 
.A1(n_399),
.A2(n_421),
.B1(n_412),
.B2(n_284),
.Y(n_453)
);

OAI22xp5_ASAP7_75t_SL g400 ( 
.A1(n_317),
.A2(n_296),
.B1(n_302),
.B2(n_309),
.Y(n_400)
);

AOI22xp5_ASAP7_75t_L g426 ( 
.A1(n_400),
.A2(n_401),
.B1(n_385),
.B2(n_411),
.Y(n_426)
);

OAI22xp5_ASAP7_75t_SL g401 ( 
.A1(n_317),
.A2(n_259),
.B1(n_298),
.B2(n_274),
.Y(n_401)
);

BUFx2_ASAP7_75t_L g454 ( 
.A(n_402),
.Y(n_454)
);

CKINVDCx20_ASAP7_75t_R g403 ( 
.A(n_325),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_403),
.B(n_405),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_330),
.B(n_269),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_L g407 ( 
.A(n_340),
.B(n_271),
.Y(n_407)
);

NAND3xp33_ASAP7_75t_L g461 ( 
.A(n_407),
.B(n_418),
.C(n_422),
.Y(n_461)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_343),
.Y(n_408)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_408),
.Y(n_459)
);

OR2x2_ASAP7_75t_SL g409 ( 
.A(n_342),
.B(n_236),
.Y(n_409)
);

OAI21xp33_ASAP7_75t_L g464 ( 
.A1(n_409),
.A2(n_329),
.B(n_278),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_316),
.B(n_335),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_410),
.B(n_420),
.Y(n_435)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_328),
.Y(n_411)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_411),
.Y(n_465)
);

OAI21xp5_ASAP7_75t_L g412 ( 
.A1(n_323),
.A2(n_278),
.B(n_236),
.Y(n_412)
);

OAI21xp5_ASAP7_75t_L g433 ( 
.A1(n_412),
.A2(n_423),
.B(n_392),
.Y(n_433)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_343),
.Y(n_413)
);

AOI22xp33_ASAP7_75t_SL g457 ( 
.A1(n_413),
.A2(n_416),
.B1(n_417),
.B2(n_419),
.Y(n_457)
);

CKINVDCx16_ASAP7_75t_R g447 ( 
.A(n_415),
.Y(n_447)
);

INVx8_ASAP7_75t_L g416 ( 
.A(n_320),
.Y(n_416)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_321),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_SL g418 ( 
.A(n_316),
.B(n_233),
.Y(n_418)
);

BUFx24_ASAP7_75t_L g419 ( 
.A(n_345),
.Y(n_419)
);

CKINVDCx20_ASAP7_75t_R g420 ( 
.A(n_325),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_L g422 ( 
.A(n_344),
.B(n_284),
.Y(n_422)
);

AOI21xp5_ASAP7_75t_L g423 ( 
.A1(n_369),
.A2(n_348),
.B(n_360),
.Y(n_423)
);

AOI21xp5_ASAP7_75t_L g450 ( 
.A1(n_423),
.A2(n_314),
.B(n_359),
.Y(n_450)
);

INVxp67_ASAP7_75t_L g424 ( 
.A(n_314),
.Y(n_424)
);

CKINVDCx20_ASAP7_75t_R g428 ( 
.A(n_424),
.Y(n_428)
);

INVx2_ASAP7_75t_L g425 ( 
.A(n_321),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_425),
.B(n_315),
.Y(n_440)
);

AND2x2_ASAP7_75t_L g478 ( 
.A(n_426),
.B(n_464),
.Y(n_478)
);

XNOR2xp5_ASAP7_75t_L g427 ( 
.A(n_396),
.B(n_313),
.Y(n_427)
);

XNOR2xp5_ASAP7_75t_SL g499 ( 
.A(n_427),
.B(n_449),
.Y(n_499)
);

XOR2xp5_ASAP7_75t_L g429 ( 
.A(n_396),
.B(n_410),
.Y(n_429)
);

MAJIxp5_ASAP7_75t_L g488 ( 
.A(n_429),
.B(n_437),
.C(n_444),
.Y(n_488)
);

AOI22xp5_ASAP7_75t_L g430 ( 
.A1(n_380),
.A2(n_348),
.B1(n_372),
.B2(n_319),
.Y(n_430)
);

AOI22xp5_ASAP7_75t_L g470 ( 
.A1(n_430),
.A2(n_438),
.B1(n_448),
.B2(n_452),
.Y(n_470)
);

OAI21xp5_ASAP7_75t_SL g501 ( 
.A1(n_433),
.A2(n_441),
.B(n_442),
.Y(n_501)
);

MAJIxp5_ASAP7_75t_L g437 ( 
.A(n_414),
.B(n_368),
.C(n_333),
.Y(n_437)
);

AOI22xp5_ASAP7_75t_L g438 ( 
.A1(n_380),
.A2(n_319),
.B1(n_334),
.B2(n_361),
.Y(n_438)
);

NOR2x1_ASAP7_75t_L g439 ( 
.A(n_378),
.B(n_319),
.Y(n_439)
);

NOR2xp33_ASAP7_75t_L g469 ( 
.A(n_439),
.B(n_395),
.Y(n_469)
);

INVxp67_ASAP7_75t_L g491 ( 
.A(n_440),
.Y(n_491)
);

OAI21xp5_ASAP7_75t_L g441 ( 
.A1(n_380),
.A2(n_326),
.B(n_322),
.Y(n_441)
);

OAI21xp5_ASAP7_75t_L g442 ( 
.A1(n_414),
.A2(n_370),
.B(n_315),
.Y(n_442)
);

MAJIxp5_ASAP7_75t_L g444 ( 
.A(n_377),
.B(n_333),
.C(n_324),
.Y(n_444)
);

XOR2xp5_ASAP7_75t_L g445 ( 
.A(n_383),
.B(n_342),
.Y(n_445)
);

MAJIxp5_ASAP7_75t_L g504 ( 
.A(n_445),
.B(n_451),
.C(n_455),
.Y(n_504)
);

AOI22xp5_ASAP7_75t_L g448 ( 
.A1(n_388),
.A2(n_329),
.B1(n_347),
.B2(n_332),
.Y(n_448)
);

XNOR2xp5_ASAP7_75t_L g449 ( 
.A(n_377),
.B(n_353),
.Y(n_449)
);

OAI21xp5_ASAP7_75t_L g477 ( 
.A1(n_450),
.A2(n_404),
.B(n_398),
.Y(n_477)
);

XOR2xp5_ASAP7_75t_L g451 ( 
.A(n_383),
.B(n_338),
.Y(n_451)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_453),
.Y(n_468)
);

XOR2xp5_ASAP7_75t_L g455 ( 
.A(n_397),
.B(n_358),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_397),
.B(n_363),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_460),
.B(n_463),
.Y(n_480)
);

AOI21xp5_ASAP7_75t_L g462 ( 
.A1(n_406),
.A2(n_293),
.B(n_268),
.Y(n_462)
);

A2O1A1Ixp33_ASAP7_75t_SL g493 ( 
.A1(n_462),
.A2(n_419),
.B(n_387),
.C(n_400),
.Y(n_493)
);

CKINVDCx20_ASAP7_75t_R g463 ( 
.A(n_389),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_467),
.B(n_449),
.Y(n_483)
);

OAI21xp5_ASAP7_75t_SL g508 ( 
.A1(n_469),
.A2(n_477),
.B(n_500),
.Y(n_508)
);

XNOR2xp5_ASAP7_75t_L g471 ( 
.A(n_429),
.B(n_381),
.Y(n_471)
);

XOR2xp5_ASAP7_75t_L g521 ( 
.A(n_471),
.B(n_459),
.Y(n_521)
);

NOR2xp33_ASAP7_75t_SL g472 ( 
.A(n_443),
.B(n_379),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_SL g523 ( 
.A(n_472),
.B(n_473),
.Y(n_523)
);

CKINVDCx20_ASAP7_75t_R g473 ( 
.A(n_467),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_440),
.Y(n_474)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_474),
.Y(n_510)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_434),
.Y(n_475)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_475),
.Y(n_520)
);

AND2x6_ASAP7_75t_L g476 ( 
.A(n_446),
.B(n_394),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g513 ( 
.A(n_476),
.B(n_484),
.Y(n_513)
);

AND2x2_ASAP7_75t_L g479 ( 
.A(n_433),
.B(n_450),
.Y(n_479)
);

INVxp67_ASAP7_75t_L g517 ( 
.A(n_479),
.Y(n_517)
);

INVx5_ASAP7_75t_L g481 ( 
.A(n_461),
.Y(n_481)
);

BUFx3_ASAP7_75t_L g528 ( 
.A(n_481),
.Y(n_528)
);

MAJIxp5_ASAP7_75t_SL g482 ( 
.A(n_427),
.B(n_409),
.C(n_401),
.Y(n_482)
);

NOR2xp33_ASAP7_75t_SL g509 ( 
.A(n_482),
.B(n_490),
.Y(n_509)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_483),
.Y(n_522)
);

AND2x6_ASAP7_75t_L g484 ( 
.A(n_446),
.B(n_439),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_434),
.Y(n_485)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_485),
.Y(n_529)
);

CKINVDCx16_ASAP7_75t_R g486 ( 
.A(n_431),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_SL g530 ( 
.A(n_486),
.B(n_496),
.Y(n_530)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_465),
.Y(n_487)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_487),
.Y(n_541)
);

INVx13_ASAP7_75t_L g489 ( 
.A(n_458),
.Y(n_489)
);

INVxp33_ASAP7_75t_L g534 ( 
.A(n_489),
.Y(n_534)
);

NOR2xp33_ASAP7_75t_L g490 ( 
.A(n_432),
.B(n_420),
.Y(n_490)
);

AND2x2_ASAP7_75t_L g492 ( 
.A(n_441),
.B(n_405),
.Y(n_492)
);

AND2x2_ASAP7_75t_L g543 ( 
.A(n_492),
.B(n_494),
.Y(n_543)
);

OAI21xp5_ASAP7_75t_L g535 ( 
.A1(n_493),
.A2(n_456),
.B(n_318),
.Y(n_535)
);

AND2x2_ASAP7_75t_L g494 ( 
.A(n_462),
.B(n_403),
.Y(n_494)
);

AND2x6_ASAP7_75t_L g495 ( 
.A(n_430),
.B(n_402),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_495),
.B(n_468),
.Y(n_524)
);

NOR2xp33_ASAP7_75t_SL g496 ( 
.A(n_444),
.B(n_419),
.Y(n_496)
);

CKINVDCx20_ASAP7_75t_R g497 ( 
.A(n_431),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_SL g537 ( 
.A(n_497),
.B(n_413),
.Y(n_537)
);

AND2x2_ASAP7_75t_L g498 ( 
.A(n_442),
.B(n_404),
.Y(n_498)
);

CKINVDCx20_ASAP7_75t_R g515 ( 
.A(n_498),
.Y(n_515)
);

OAI21xp5_ASAP7_75t_L g500 ( 
.A1(n_435),
.A2(n_376),
.B(n_384),
.Y(n_500)
);

INVx2_ASAP7_75t_L g502 ( 
.A(n_465),
.Y(n_502)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_502),
.Y(n_544)
);

AOI22xp5_ASAP7_75t_L g503 ( 
.A1(n_452),
.A2(n_376),
.B1(n_384),
.B2(n_424),
.Y(n_503)
);

OAI22xp5_ASAP7_75t_L g514 ( 
.A1(n_503),
.A2(n_448),
.B1(n_426),
.B2(n_491),
.Y(n_514)
);

XOR2xp5_ASAP7_75t_L g505 ( 
.A(n_437),
.B(n_233),
.Y(n_505)
);

MAJIxp5_ASAP7_75t_L g511 ( 
.A(n_505),
.B(n_445),
.C(n_451),
.Y(n_511)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_435),
.Y(n_506)
);

NOR2xp33_ASAP7_75t_L g526 ( 
.A(n_506),
.B(n_500),
.Y(n_526)
);

AOI22xp5_ASAP7_75t_SL g507 ( 
.A1(n_498),
.A2(n_454),
.B1(n_447),
.B2(n_460),
.Y(n_507)
);

OAI21xp5_ASAP7_75t_SL g570 ( 
.A1(n_507),
.A2(n_524),
.B(n_535),
.Y(n_570)
);

MAJIxp5_ASAP7_75t_L g563 ( 
.A(n_511),
.B(n_536),
.C(n_386),
.Y(n_563)
);

XNOR2xp5_ASAP7_75t_L g512 ( 
.A(n_488),
.B(n_455),
.Y(n_512)
);

XOR2xp5_ASAP7_75t_L g560 ( 
.A(n_512),
.B(n_521),
.Y(n_560)
);

OAI22xp5_ASAP7_75t_L g553 ( 
.A1(n_514),
.A2(n_538),
.B1(n_493),
.B2(n_356),
.Y(n_553)
);

NOR2xp33_ASAP7_75t_SL g516 ( 
.A(n_481),
.B(n_428),
.Y(n_516)
);

NAND3xp33_ASAP7_75t_L g576 ( 
.A(n_516),
.B(n_525),
.C(n_540),
.Y(n_576)
);

OAI22xp5_ASAP7_75t_SL g518 ( 
.A1(n_470),
.A2(n_454),
.B1(n_438),
.B2(n_457),
.Y(n_518)
);

AOI22xp5_ASAP7_75t_L g572 ( 
.A1(n_518),
.A2(n_519),
.B1(n_337),
.B2(n_364),
.Y(n_572)
);

OAI22xp5_ASAP7_75t_SL g519 ( 
.A1(n_470),
.A2(n_459),
.B1(n_466),
.B2(n_456),
.Y(n_519)
);

NOR2xp33_ASAP7_75t_SL g525 ( 
.A(n_480),
.B(n_419),
.Y(n_525)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_526),
.Y(n_567)
);

XOR2xp5_ASAP7_75t_L g527 ( 
.A(n_488),
.B(n_425),
.Y(n_527)
);

XOR2xp5_ASAP7_75t_L g573 ( 
.A(n_527),
.B(n_533),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_L g531 ( 
.A(n_491),
.B(n_466),
.Y(n_531)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_531),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_503),
.B(n_502),
.Y(n_532)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_532),
.Y(n_559)
);

XNOR2xp5_ASAP7_75t_L g533 ( 
.A(n_504),
.B(n_257),
.Y(n_533)
);

MAJIxp5_ASAP7_75t_L g536 ( 
.A(n_505),
.B(n_257),
.C(n_417),
.Y(n_536)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_537),
.Y(n_571)
);

AOI22xp5_ASAP7_75t_L g538 ( 
.A1(n_478),
.A2(n_436),
.B1(n_391),
.B2(n_416),
.Y(n_538)
);

NOR2xp33_ASAP7_75t_L g539 ( 
.A(n_471),
.B(n_375),
.Y(n_539)
);

NOR2xp33_ASAP7_75t_SL g565 ( 
.A(n_539),
.B(n_545),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_SL g540 ( 
.A(n_504),
.B(n_408),
.Y(n_540)
);

CKINVDCx20_ASAP7_75t_R g542 ( 
.A(n_494),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_L g549 ( 
.A(n_542),
.B(n_478),
.Y(n_549)
);

NOR2xp33_ASAP7_75t_SL g545 ( 
.A(n_498),
.B(n_436),
.Y(n_545)
);

OAI22xp5_ASAP7_75t_SL g547 ( 
.A1(n_524),
.A2(n_478),
.B1(n_492),
.B2(n_479),
.Y(n_547)
);

AOI22xp5_ASAP7_75t_L g601 ( 
.A1(n_547),
.A2(n_550),
.B1(n_552),
.B2(n_553),
.Y(n_601)
);

CKINVDCx14_ASAP7_75t_R g548 ( 
.A(n_523),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_L g583 ( 
.A(n_548),
.B(n_555),
.Y(n_583)
);

CKINVDCx20_ASAP7_75t_R g586 ( 
.A(n_549),
.Y(n_586)
);

OAI22xp5_ASAP7_75t_SL g550 ( 
.A1(n_513),
.A2(n_492),
.B1(n_479),
.B2(n_476),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_531),
.B(n_493),
.Y(n_551)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_551),
.Y(n_596)
);

OAI22xp5_ASAP7_75t_SL g552 ( 
.A1(n_513),
.A2(n_477),
.B1(n_495),
.B2(n_494),
.Y(n_552)
);

INVx3_ASAP7_75t_L g554 ( 
.A(n_528),
.Y(n_554)
);

HB1xp67_ASAP7_75t_L g606 ( 
.A(n_554),
.Y(n_606)
);

INVx3_ASAP7_75t_L g555 ( 
.A(n_528),
.Y(n_555)
);

OAI22xp5_ASAP7_75t_SL g556 ( 
.A1(n_515),
.A2(n_501),
.B1(n_484),
.B2(n_493),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_L g594 ( 
.A(n_556),
.B(n_558),
.Y(n_594)
);

OAI22xp5_ASAP7_75t_L g557 ( 
.A1(n_507),
.A2(n_501),
.B1(n_499),
.B2(n_489),
.Y(n_557)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_557),
.Y(n_598)
);

INVxp67_ASAP7_75t_L g558 ( 
.A(n_545),
.Y(n_558)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_544),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_L g597 ( 
.A(n_561),
.B(n_562),
.Y(n_597)
);

OAI22xp5_ASAP7_75t_SL g562 ( 
.A1(n_515),
.A2(n_499),
.B1(n_357),
.B2(n_337),
.Y(n_562)
);

XNOR2xp5_ASAP7_75t_L g587 ( 
.A(n_563),
.B(n_536),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_L g564 ( 
.A(n_532),
.B(n_382),
.Y(n_564)
);

INVxp67_ASAP7_75t_SL g603 ( 
.A(n_564),
.Y(n_603)
);

CKINVDCx20_ASAP7_75t_R g566 ( 
.A(n_543),
.Y(n_566)
);

NOR2xp33_ASAP7_75t_L g595 ( 
.A(n_566),
.B(n_569),
.Y(n_595)
);

OAI22xp5_ASAP7_75t_SL g568 ( 
.A1(n_542),
.A2(n_510),
.B1(n_543),
.B2(n_517),
.Y(n_568)
);

OAI22xp5_ASAP7_75t_SL g581 ( 
.A1(n_568),
.A2(n_572),
.B1(n_574),
.B2(n_578),
.Y(n_581)
);

NOR2xp33_ASAP7_75t_SL g569 ( 
.A(n_530),
.B(n_375),
.Y(n_569)
);

OAI22xp5_ASAP7_75t_SL g574 ( 
.A1(n_510),
.A2(n_357),
.B1(n_364),
.B2(n_260),
.Y(n_574)
);

XOR2xp5_ASAP7_75t_L g575 ( 
.A(n_512),
.B(n_245),
.Y(n_575)
);

XOR2xp5_ASAP7_75t_L g584 ( 
.A(n_575),
.B(n_511),
.Y(n_584)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_520),
.Y(n_577)
);

CKINVDCx16_ASAP7_75t_R g589 ( 
.A(n_577),
.Y(n_589)
);

AOI22xp5_ASAP7_75t_SL g578 ( 
.A1(n_518),
.A2(n_294),
.B1(n_271),
.B2(n_258),
.Y(n_578)
);

CKINVDCx20_ASAP7_75t_R g579 ( 
.A(n_543),
.Y(n_579)
);

AOI21xp5_ASAP7_75t_L g580 ( 
.A1(n_579),
.A2(n_508),
.B(n_517),
.Y(n_580)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_580),
.Y(n_613)
);

MAJIxp5_ASAP7_75t_L g582 ( 
.A(n_563),
.B(n_527),
.C(n_533),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_L g615 ( 
.A(n_582),
.B(n_585),
.Y(n_615)
);

XOR2xp5_ASAP7_75t_L g610 ( 
.A(n_584),
.B(n_607),
.Y(n_610)
);

MAJIxp5_ASAP7_75t_L g585 ( 
.A(n_573),
.B(n_560),
.C(n_575),
.Y(n_585)
);

XNOR2xp5_ASAP7_75t_L g618 ( 
.A(n_587),
.B(n_588),
.Y(n_618)
);

XNOR2xp5_ASAP7_75t_L g588 ( 
.A(n_573),
.B(n_521),
.Y(n_588)
);

MAJIxp5_ASAP7_75t_L g590 ( 
.A(n_560),
.B(n_508),
.C(n_519),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_L g631 ( 
.A(n_590),
.B(n_602),
.Y(n_631)
);

XNOR2xp5_ASAP7_75t_SL g591 ( 
.A(n_550),
.B(n_509),
.Y(n_591)
);

MAJx2_ASAP7_75t_L g612 ( 
.A(n_591),
.B(n_592),
.C(n_604),
.Y(n_612)
);

XOR2xp5_ASAP7_75t_L g592 ( 
.A(n_547),
.B(n_522),
.Y(n_592)
);

OAI21xp5_ASAP7_75t_L g593 ( 
.A1(n_549),
.A2(n_535),
.B(n_538),
.Y(n_593)
);

OAI21xp5_ASAP7_75t_SL g628 ( 
.A1(n_593),
.A2(n_599),
.B(n_570),
.Y(n_628)
);

OAI21xp5_ASAP7_75t_L g599 ( 
.A1(n_551),
.A2(n_544),
.B(n_534),
.Y(n_599)
);

OAI22xp5_ASAP7_75t_SL g600 ( 
.A1(n_559),
.A2(n_522),
.B1(n_529),
.B2(n_541),
.Y(n_600)
);

AOI22xp5_ASAP7_75t_L g619 ( 
.A1(n_600),
.A2(n_546),
.B1(n_561),
.B2(n_564),
.Y(n_619)
);

MAJIxp5_ASAP7_75t_L g602 ( 
.A(n_562),
.B(n_541),
.C(n_529),
.Y(n_602)
);

XOR2xp5_ASAP7_75t_L g604 ( 
.A(n_556),
.B(n_520),
.Y(n_604)
);

NOR3xp33_ASAP7_75t_SL g605 ( 
.A(n_567),
.B(n_318),
.C(n_222),
.Y(n_605)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_605),
.Y(n_617)
);

XOR2xp5_ASAP7_75t_L g607 ( 
.A(n_552),
.B(n_568),
.Y(n_607)
);

MAJIxp5_ASAP7_75t_L g608 ( 
.A(n_582),
.B(n_587),
.C(n_584),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_L g640 ( 
.A(n_608),
.B(n_611),
.Y(n_640)
);

NOR2xp33_ASAP7_75t_L g609 ( 
.A(n_583),
.B(n_555),
.Y(n_609)
);

CKINVDCx14_ASAP7_75t_R g637 ( 
.A(n_609),
.Y(n_637)
);

MAJIxp5_ASAP7_75t_L g611 ( 
.A(n_585),
.B(n_558),
.C(n_559),
.Y(n_611)
);

BUFx24_ASAP7_75t_SL g614 ( 
.A(n_586),
.Y(n_614)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_614),
.Y(n_632)
);

OAI22xp5_ASAP7_75t_SL g616 ( 
.A1(n_601),
.A2(n_572),
.B1(n_546),
.B2(n_578),
.Y(n_616)
);

AOI22xp5_ASAP7_75t_L g645 ( 
.A1(n_616),
.A2(n_295),
.B1(n_290),
.B2(n_293),
.Y(n_645)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_619),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g620 ( 
.A(n_595),
.B(n_571),
.Y(n_620)
);

AOI21xp5_ASAP7_75t_L g638 ( 
.A1(n_620),
.A2(n_627),
.B(n_629),
.Y(n_638)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_600),
.Y(n_621)
);

AOI22xp33_ASAP7_75t_SL g633 ( 
.A1(n_621),
.A2(n_623),
.B1(n_626),
.B2(n_598),
.Y(n_633)
);

XNOR2xp5_ASAP7_75t_L g622 ( 
.A(n_590),
.B(n_570),
.Y(n_622)
);

XNOR2xp5_ASAP7_75t_L g644 ( 
.A(n_622),
.B(n_605),
.Y(n_644)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_603),
.Y(n_623)
);

INVxp67_ASAP7_75t_L g624 ( 
.A(n_599),
.Y(n_624)
);

AND2x2_ASAP7_75t_L g636 ( 
.A(n_624),
.B(n_597),
.Y(n_636)
);

CKINVDCx14_ASAP7_75t_R g625 ( 
.A(n_602),
.Y(n_625)
);

OAI22xp5_ASAP7_75t_L g634 ( 
.A1(n_625),
.A2(n_601),
.B1(n_607),
.B2(n_604),
.Y(n_634)
);

HB1xp67_ASAP7_75t_L g626 ( 
.A(n_606),
.Y(n_626)
);

NOR2xp33_ASAP7_75t_L g627 ( 
.A(n_592),
.B(n_554),
.Y(n_627)
);

AOI21xp5_ASAP7_75t_L g648 ( 
.A1(n_628),
.A2(n_630),
.B(n_245),
.Y(n_648)
);

OAI21xp5_ASAP7_75t_SL g629 ( 
.A1(n_594),
.A2(n_576),
.B(n_565),
.Y(n_629)
);

AOI21xp5_ASAP7_75t_L g630 ( 
.A1(n_593),
.A2(n_574),
.B(n_268),
.Y(n_630)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_633),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_634),
.Y(n_653)
);

XOR2xp5_ASAP7_75t_L g635 ( 
.A(n_610),
.B(n_588),
.Y(n_635)
);

AND2x2_ASAP7_75t_L g661 ( 
.A(n_635),
.B(n_644),
.Y(n_661)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_636),
.Y(n_664)
);

MAJIxp5_ASAP7_75t_L g639 ( 
.A(n_608),
.B(n_591),
.C(n_596),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_L g662 ( 
.A(n_639),
.B(n_641),
.Y(n_662)
);

MAJIxp5_ASAP7_75t_L g641 ( 
.A(n_611),
.B(n_581),
.C(n_589),
.Y(n_641)
);

INVx11_ASAP7_75t_L g642 ( 
.A(n_629),
.Y(n_642)
);

NOR2xp33_ASAP7_75t_L g658 ( 
.A(n_642),
.B(n_612),
.Y(n_658)
);

MAJIxp5_ASAP7_75t_L g643 ( 
.A(n_618),
.B(n_581),
.C(n_290),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_SL g657 ( 
.A(n_643),
.B(n_646),
.Y(n_657)
);

XOR2xp5_ASAP7_75t_L g656 ( 
.A(n_645),
.B(n_647),
.Y(n_656)
);

MAJIxp5_ASAP7_75t_L g646 ( 
.A(n_618),
.B(n_295),
.C(n_244),
.Y(n_646)
);

XNOR2x1_ASAP7_75t_L g647 ( 
.A(n_612),
.B(n_256),
.Y(n_647)
);

XOR2xp5_ASAP7_75t_L g663 ( 
.A(n_648),
.B(n_649),
.Y(n_663)
);

OA21x2_ASAP7_75t_L g649 ( 
.A1(n_616),
.A2(n_256),
.B(n_171),
.Y(n_649)
);

OAI22xp5_ASAP7_75t_SL g650 ( 
.A1(n_613),
.A2(n_171),
.B1(n_168),
.B2(n_156),
.Y(n_650)
);

AOI22xp5_ASAP7_75t_SL g667 ( 
.A1(n_650),
.A2(n_156),
.B1(n_133),
.B2(n_8),
.Y(n_667)
);

AOI21xp5_ASAP7_75t_SL g654 ( 
.A1(n_651),
.A2(n_628),
.B(n_624),
.Y(n_654)
);

AOI21x1_ASAP7_75t_SL g673 ( 
.A1(n_654),
.A2(n_648),
.B(n_642),
.Y(n_673)
);

OAI21x1_ASAP7_75t_L g655 ( 
.A1(n_638),
.A2(n_620),
.B(n_631),
.Y(n_655)
);

OR2x2_ASAP7_75t_L g675 ( 
.A(n_655),
.B(n_658),
.Y(n_675)
);

MAJIxp5_ASAP7_75t_L g659 ( 
.A(n_640),
.B(n_615),
.C(n_610),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_659),
.B(n_660),
.Y(n_669)
);

NOR2xp33_ASAP7_75t_L g660 ( 
.A(n_632),
.B(n_617),
.Y(n_660)
);

MAJIxp5_ASAP7_75t_L g665 ( 
.A(n_641),
.B(n_622),
.C(n_619),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_665),
.B(n_666),
.Y(n_677)
);

MAJIxp5_ASAP7_75t_L g666 ( 
.A(n_639),
.B(n_630),
.C(n_168),
.Y(n_666)
);

OAI21xp5_ASAP7_75t_L g674 ( 
.A1(n_667),
.A2(n_649),
.B(n_644),
.Y(n_674)
);

NOR2xp33_ASAP7_75t_L g668 ( 
.A(n_659),
.B(n_637),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_L g681 ( 
.A(n_668),
.B(n_670),
.Y(n_681)
);

MAJIxp5_ASAP7_75t_L g670 ( 
.A(n_665),
.B(n_635),
.C(n_643),
.Y(n_670)
);

NOR2xp33_ASAP7_75t_L g671 ( 
.A(n_662),
.B(n_636),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_671),
.B(n_672),
.Y(n_687)
);

NOR2xp33_ASAP7_75t_L g672 ( 
.A(n_653),
.B(n_636),
.Y(n_672)
);

OAI21xp5_ASAP7_75t_L g684 ( 
.A1(n_673),
.A2(n_663),
.B(n_649),
.Y(n_684)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_674),
.Y(n_686)
);

NOR2xp33_ASAP7_75t_L g676 ( 
.A(n_652),
.B(n_646),
.Y(n_676)
);

NOR2xp33_ASAP7_75t_SL g685 ( 
.A(n_676),
.B(n_678),
.Y(n_685)
);

CKINVDCx20_ASAP7_75t_R g678 ( 
.A(n_661),
.Y(n_678)
);

NOR2xp33_ASAP7_75t_SL g679 ( 
.A(n_661),
.B(n_650),
.Y(n_679)
);

NOR2xp33_ASAP7_75t_L g688 ( 
.A(n_679),
.B(n_656),
.Y(n_688)
);

AOI22xp5_ASAP7_75t_L g680 ( 
.A1(n_675),
.A2(n_664),
.B1(n_657),
.B2(n_663),
.Y(n_680)
);

INVxp33_ASAP7_75t_L g693 ( 
.A(n_680),
.Y(n_693)
);

XOR2xp5_ASAP7_75t_L g682 ( 
.A(n_670),
.B(n_654),
.Y(n_682)
);

NOR2xp33_ASAP7_75t_L g692 ( 
.A(n_682),
.B(n_684),
.Y(n_692)
);

XNOR2xp5_ASAP7_75t_SL g683 ( 
.A(n_669),
.B(n_647),
.Y(n_683)
);

INVxp67_ASAP7_75t_L g689 ( 
.A(n_683),
.Y(n_689)
);

OAI21xp33_ASAP7_75t_L g691 ( 
.A1(n_688),
.A2(n_673),
.B(n_645),
.Y(n_691)
);

OA21x2_ASAP7_75t_SL g690 ( 
.A1(n_687),
.A2(n_677),
.B(n_675),
.Y(n_690)
);

NOR2xp33_ASAP7_75t_SL g694 ( 
.A(n_690),
.B(n_681),
.Y(n_694)
);

AOI22xp5_ASAP7_75t_L g696 ( 
.A1(n_691),
.A2(n_685),
.B1(n_656),
.B2(n_133),
.Y(n_696)
);

NOR3xp33_ASAP7_75t_L g698 ( 
.A(n_694),
.B(n_692),
.C(n_689),
.Y(n_698)
);

MAJIxp5_ASAP7_75t_L g695 ( 
.A(n_693),
.B(n_686),
.C(n_688),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_695),
.B(n_696),
.Y(n_697)
);

OAI321xp33_ASAP7_75t_L g699 ( 
.A1(n_698),
.A2(n_697),
.A3(n_6),
.B1(n_8),
.B2(n_9),
.C(n_5),
.Y(n_699)
);

OAI21xp5_ASAP7_75t_L g700 ( 
.A1(n_699),
.A2(n_5),
.B(n_6),
.Y(n_700)
);

OAI22xp5_ASAP7_75t_SL g701 ( 
.A1(n_700),
.A2(n_8),
.B1(n_10),
.B2(n_11),
.Y(n_701)
);

O2A1O1Ixp33_ASAP7_75t_SL g702 ( 
.A1(n_701),
.A2(n_10),
.B(n_12),
.C(n_249),
.Y(n_702)
);


endmodule