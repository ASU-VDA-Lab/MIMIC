module fake_jpeg_12606_n_96 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_96);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_96;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_2),
.Y(n_11)
);

BUFx12_ASAP7_75t_L g12 ( 
.A(n_6),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_6),
.Y(n_13)
);

BUFx12f_ASAP7_75t_L g14 ( 
.A(n_4),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_2),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

INVxp67_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

INVx5_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_8),
.B(n_9),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_SL g22 ( 
.A(n_4),
.B(n_0),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_22),
.B(n_0),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_SL g39 ( 
.A(n_24),
.B(n_25),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g25 ( 
.A1(n_18),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_23),
.Y(n_26)
);

OR2x2_ASAP7_75t_L g40 ( 
.A(n_26),
.B(n_13),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_21),
.B(n_3),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_27),
.B(n_29),
.Y(n_38)
);

INVx5_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_28),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_17),
.B(n_3),
.Y(n_29)
);

INVx2_ASAP7_75t_SL g30 ( 
.A(n_14),
.Y(n_30)
);

INVx5_ASAP7_75t_SL g43 ( 
.A(n_30),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_SL g31 ( 
.A(n_23),
.B(n_3),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_31),
.B(n_11),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_L g32 ( 
.A1(n_18),
.A2(n_4),
.B1(n_5),
.B2(n_7),
.Y(n_32)
);

OR2x2_ASAP7_75t_L g44 ( 
.A(n_32),
.B(n_20),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_33),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_35),
.B(n_37),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_31),
.B(n_24),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_40),
.B(n_42),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g41 ( 
.A1(n_30),
.A2(n_20),
.B1(n_17),
.B2(n_14),
.Y(n_41)
);

INVxp67_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_27),
.B(n_13),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_L g51 ( 
.A1(n_44),
.A2(n_30),
.B1(n_28),
.B2(n_33),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_29),
.B(n_11),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_45),
.B(n_15),
.Y(n_52)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_43),
.Y(n_48)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_48),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_40),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_49),
.B(n_52),
.Y(n_64)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_50),
.Y(n_62)
);

CKINVDCx16_ASAP7_75t_R g60 ( 
.A(n_51),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_39),
.A2(n_25),
.B1(n_26),
.B2(n_33),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_53),
.A2(n_44),
.B1(n_38),
.B2(n_36),
.Y(n_63)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_43),
.Y(n_54)
);

OAI21xp33_ASAP7_75t_L g58 ( 
.A1(n_54),
.A2(n_57),
.B(n_48),
.Y(n_58)
);

OAI21xp5_ASAP7_75t_SL g56 ( 
.A1(n_39),
.A2(n_15),
.B(n_12),
.Y(n_56)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_56),
.B(n_16),
.C(n_19),
.Y(n_65)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

XNOR2xp5_ASAP7_75t_L g73 ( 
.A(n_58),
.B(n_65),
.Y(n_73)
);

FAx1_ASAP7_75t_SL g61 ( 
.A(n_47),
.B(n_37),
.CI(n_35),
.CON(n_61),
.SN(n_61)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_61),
.B(n_66),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_63),
.A2(n_67),
.B1(n_54),
.B2(n_55),
.Y(n_75)
);

CKINVDCx16_ASAP7_75t_R g66 ( 
.A(n_51),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_53),
.A2(n_16),
.B1(n_19),
.B2(n_34),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_64),
.B(n_46),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_68),
.B(n_71),
.Y(n_81)
);

XNOR2xp5_ASAP7_75t_L g69 ( 
.A(n_61),
.B(n_47),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_69),
.B(n_70),
.C(n_74),
.Y(n_78)
);

XNOR2xp5_ASAP7_75t_L g70 ( 
.A(n_61),
.B(n_56),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_63),
.B(n_52),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_65),
.B(n_57),
.C(n_55),
.Y(n_74)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_75),
.Y(n_76)
);

XOR2x2_ASAP7_75t_L g77 ( 
.A(n_69),
.B(n_59),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_77),
.A2(n_74),
.B1(n_70),
.B2(n_60),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_SL g79 ( 
.A1(n_72),
.A2(n_60),
.B(n_59),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_79),
.A2(n_67),
.B1(n_62),
.B2(n_34),
.Y(n_84)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_73),
.Y(n_80)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_80),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_82),
.B(n_84),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_76),
.A2(n_62),
.B1(n_50),
.B2(n_34),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_85),
.B(n_86),
.Y(n_89)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_81),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_83),
.B(n_77),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_87),
.B(n_82),
.Y(n_90)
);

AOI21xp5_ASAP7_75t_L g93 ( 
.A1(n_90),
.A2(n_91),
.B(n_92),
.Y(n_93)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_89),
.B(n_85),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_88),
.A2(n_78),
.B1(n_9),
.B2(n_10),
.Y(n_92)
);

AOI21xp5_ASAP7_75t_L g94 ( 
.A1(n_91),
.A2(n_78),
.B(n_8),
.Y(n_94)
);

AOI31xp33_ASAP7_75t_L g95 ( 
.A1(n_94),
.A2(n_12),
.A3(n_42),
.B(n_52),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_95),
.B(n_93),
.Y(n_96)
);


endmodule