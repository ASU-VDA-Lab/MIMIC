module fake_jpeg_14477_n_187 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_187);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_187;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_182;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_93;
wire n_91;
wire n_54;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

INVx3_ASAP7_75t_L g48 ( 
.A(n_29),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_25),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_33),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_7),
.Y(n_51)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_4),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_38),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_42),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_2),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_10),
.Y(n_57)
);

BUFx16f_ASAP7_75t_L g58 ( 
.A(n_36),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_32),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_7),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_17),
.Y(n_61)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_37),
.Y(n_62)
);

CKINVDCx16_ASAP7_75t_R g63 ( 
.A(n_24),
.Y(n_63)
);

BUFx5_ASAP7_75t_L g64 ( 
.A(n_44),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_1),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_13),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_26),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_40),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_45),
.Y(n_69)
);

BUFx5_ASAP7_75t_L g70 ( 
.A(n_21),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_16),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_34),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_46),
.Y(n_73)
);

BUFx5_ASAP7_75t_L g74 ( 
.A(n_5),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_6),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_43),
.Y(n_76)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_47),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_62),
.Y(n_78)
);

INVx8_ASAP7_75t_L g102 ( 
.A(n_78),
.Y(n_102)
);

INVx11_ASAP7_75t_L g79 ( 
.A(n_74),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_79),
.Y(n_91)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_74),
.Y(n_80)
);

BUFx3_ASAP7_75t_L g89 ( 
.A(n_80),
.Y(n_89)
);

BUFx8_ASAP7_75t_L g81 ( 
.A(n_58),
.Y(n_81)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_81),
.Y(n_93)
);

INVx4_ASAP7_75t_SL g82 ( 
.A(n_60),
.Y(n_82)
);

NAND2xp33_ASAP7_75t_SL g100 ( 
.A(n_82),
.B(n_85),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_60),
.Y(n_83)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_83),
.Y(n_96)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_51),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_84),
.B(n_86),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_62),
.Y(n_85)
);

OR2x2_ASAP7_75t_L g86 ( 
.A(n_50),
.B(n_0),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_62),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_87),
.B(n_70),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_53),
.B(n_0),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_88),
.B(n_57),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_L g90 ( 
.A1(n_78),
.A2(n_56),
.B1(n_65),
.B2(n_75),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_90),
.A2(n_98),
.B1(n_103),
.B2(n_64),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_85),
.B(n_52),
.C(n_48),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_94),
.B(n_95),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_97),
.B(n_99),
.Y(n_107)
);

OAI22xp33_ASAP7_75t_L g98 ( 
.A1(n_82),
.A2(n_65),
.B1(n_56),
.B2(n_77),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_88),
.B(n_66),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_81),
.B(n_67),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_101),
.B(n_1),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_83),
.A2(n_77),
.B1(n_48),
.B2(n_73),
.Y(n_103)
);

AOI21xp33_ASAP7_75t_SL g104 ( 
.A1(n_79),
.A2(n_58),
.B(n_63),
.Y(n_104)
);

OAI32xp33_ASAP7_75t_L g108 ( 
.A1(n_104),
.A2(n_59),
.A3(n_61),
.B1(n_68),
.B2(n_70),
.Y(n_108)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_96),
.Y(n_105)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_105),
.Y(n_135)
);

NOR3xp33_ASAP7_75t_L g146 ( 
.A(n_108),
.B(n_12),
.C(n_14),
.Y(n_146)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_96),
.Y(n_109)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_109),
.Y(n_142)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_102),
.Y(n_110)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_110),
.Y(n_145)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_93),
.Y(n_111)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_111),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_92),
.B(n_72),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_112),
.B(n_119),
.Y(n_141)
);

INVx6_ASAP7_75t_L g113 ( 
.A(n_102),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_113),
.B(n_115),
.Y(n_129)
);

INVx8_ASAP7_75t_L g114 ( 
.A(n_93),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_114),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_98),
.Y(n_115)
);

OA22x2_ASAP7_75t_L g116 ( 
.A1(n_100),
.A2(n_76),
.B1(n_71),
.B2(n_69),
.Y(n_116)
);

AND2x2_ASAP7_75t_L g144 ( 
.A(n_116),
.B(n_126),
.Y(n_144)
);

BUFx2_ASAP7_75t_L g117 ( 
.A(n_89),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_117),
.Y(n_133)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_89),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_118),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_94),
.Y(n_119)
);

HB1xp67_ASAP7_75t_L g120 ( 
.A(n_91),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_120),
.Y(n_143)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_91),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_121),
.B(n_122),
.Y(n_130)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_96),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_98),
.A2(n_55),
.B1(n_54),
.B2(n_49),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_123),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_136)
);

INVxp33_ASAP7_75t_L g124 ( 
.A(n_100),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_124),
.B(n_127),
.Y(n_139)
);

INVx8_ASAP7_75t_L g125 ( 
.A(n_102),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_125),
.B(n_15),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_106),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_131),
.B(n_136),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_106),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_L g161 ( 
.A1(n_132),
.A2(n_131),
.B1(n_138),
.B2(n_129),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_107),
.B(n_8),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g152 ( 
.A(n_134),
.B(n_140),
.Y(n_152)
);

CKINVDCx14_ASAP7_75t_R g137 ( 
.A(n_120),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_L g157 ( 
.A1(n_137),
.A2(n_151),
.B(n_143),
.Y(n_157)
);

OR2x2_ASAP7_75t_L g138 ( 
.A(n_116),
.B(n_9),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_138),
.B(n_146),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_107),
.B(n_11),
.Y(n_140)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_147),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_127),
.B(n_18),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g165 ( 
.A(n_148),
.B(n_150),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_106),
.B(n_19),
.Y(n_150)
);

INVxp67_ASAP7_75t_L g153 ( 
.A(n_130),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_153),
.B(n_157),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_SL g155 ( 
.A1(n_139),
.A2(n_20),
.B(n_22),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g168 ( 
.A(n_155),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_141),
.B(n_23),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_SL g170 ( 
.A(n_156),
.B(n_159),
.Y(n_170)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_145),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_158),
.B(n_160),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_144),
.B(n_27),
.C(n_28),
.Y(n_159)
);

NOR2x1_ASAP7_75t_L g160 ( 
.A(n_144),
.B(n_30),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_161),
.A2(n_167),
.B1(n_128),
.B2(n_133),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_149),
.B(n_142),
.Y(n_164)
);

CKINVDCx16_ASAP7_75t_R g173 ( 
.A(n_164),
.Y(n_173)
);

BUFx2_ASAP7_75t_L g166 ( 
.A(n_135),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_166),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_SL g167 ( 
.A(n_151),
.B(n_31),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_L g175 ( 
.A1(n_174),
.A2(n_160),
.B(n_154),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_175),
.A2(n_177),
.B1(n_178),
.B2(n_168),
.Y(n_180)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_172),
.Y(n_176)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_176),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_173),
.B(n_163),
.C(n_162),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_SL g178 ( 
.A(n_169),
.B(n_161),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_180),
.B(n_168),
.Y(n_181)
);

HB1xp67_ASAP7_75t_L g182 ( 
.A(n_181),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_182),
.B(n_179),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_183),
.A2(n_171),
.B1(n_152),
.B2(n_165),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_SL g185 ( 
.A1(n_184),
.A2(n_170),
.B(n_128),
.Y(n_185)
);

MAJx2_ASAP7_75t_L g186 ( 
.A(n_185),
.B(n_170),
.C(n_39),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_186),
.B(n_35),
.Y(n_187)
);


endmodule