module fake_jpeg_2797_n_303 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_303);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_303;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_252;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_21;
wire n_57;
wire n_187;
wire n_234;
wire n_288;
wire n_272;
wire n_284;
wire n_280;
wire n_171;
wire n_263;
wire n_119;
wire n_23;
wire n_301;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_298;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_266;
wire n_218;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_299;
wire n_211;
wire n_300;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_302;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_270;
wire n_112;
wire n_260;
wire n_199;
wire n_222;
wire n_95;
wire n_275;
wire n_256;
wire n_151;
wire n_221;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_140;
wire n_82;
wire n_128;
wire n_100;
wire n_258;
wire n_282;
wire n_96;

BUFx3_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

BUFx24_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_0),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

INVx11_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

INVx1_ASAP7_75t_SL g26 ( 
.A(n_0),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_11),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

BUFx12_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_11),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_1),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_7),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_13),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_15),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_11),
.Y(n_41)
);

OR2x2_ASAP7_75t_L g42 ( 
.A(n_3),
.B(n_7),
.Y(n_42)
);

BUFx16f_ASAP7_75t_L g43 ( 
.A(n_2),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_7),
.B(n_12),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_14),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_15),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_27),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_47),
.Y(n_111)
);

INVx11_ASAP7_75t_L g48 ( 
.A(n_20),
.Y(n_48)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_48),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_26),
.B(n_42),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g96 ( 
.A(n_49),
.B(n_84),
.Y(n_96)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_20),
.Y(n_50)
);

INVx5_ASAP7_75t_L g141 ( 
.A(n_50),
.Y(n_141)
);

BUFx12_ASAP7_75t_L g51 ( 
.A(n_43),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g134 ( 
.A(n_51),
.Y(n_134)
);

BUFx24_ASAP7_75t_L g52 ( 
.A(n_43),
.Y(n_52)
);

BUFx8_ASAP7_75t_L g136 ( 
.A(n_52),
.Y(n_136)
);

INVx11_ASAP7_75t_L g53 ( 
.A(n_20),
.Y(n_53)
);

INVx8_ASAP7_75t_L g112 ( 
.A(n_53),
.Y(n_112)
);

INVx6_ASAP7_75t_SL g54 ( 
.A(n_43),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_54),
.B(n_70),
.Y(n_97)
);

BUFx2_ASAP7_75t_L g55 ( 
.A(n_43),
.Y(n_55)
);

INVx1_ASAP7_75t_SL g113 ( 
.A(n_55),
.Y(n_113)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_21),
.Y(n_56)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_56),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_27),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_57),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_27),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_58),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_30),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_59),
.Y(n_122)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_29),
.Y(n_60)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_60),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_30),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_61),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_44),
.B(n_2),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_62),
.B(n_76),
.Y(n_107)
);

INVx3_ASAP7_75t_SL g63 ( 
.A(n_30),
.Y(n_63)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_63),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_37),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_64),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_37),
.Y(n_65)
);

INVx6_ASAP7_75t_L g143 ( 
.A(n_65),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_37),
.Y(n_66)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_66),
.Y(n_132)
);

INVx11_ASAP7_75t_L g67 ( 
.A(n_20),
.Y(n_67)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_67),
.Y(n_114)
);

INVx5_ASAP7_75t_L g68 ( 
.A(n_16),
.Y(n_68)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_68),
.Y(n_123)
);

INVx3_ASAP7_75t_SL g69 ( 
.A(n_35),
.Y(n_69)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_69),
.Y(n_125)
);

CKINVDCx16_ASAP7_75t_R g70 ( 
.A(n_17),
.Y(n_70)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_21),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_71),
.B(n_72),
.Y(n_98)
);

INVx1_ASAP7_75t_SL g72 ( 
.A(n_19),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_16),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_73),
.Y(n_130)
);

BUFx12f_ASAP7_75t_L g74 ( 
.A(n_34),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_74),
.B(n_75),
.Y(n_100)
);

INVx8_ASAP7_75t_L g75 ( 
.A(n_17),
.Y(n_75)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_29),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_42),
.B(n_2),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_77),
.B(n_79),
.Y(n_104)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_35),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_78),
.B(n_81),
.Y(n_109)
);

INVx13_ASAP7_75t_L g79 ( 
.A(n_17),
.Y(n_79)
);

INVx8_ASAP7_75t_L g80 ( 
.A(n_17),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_80),
.B(n_82),
.Y(n_105)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_38),
.Y(n_81)
);

BUFx8_ASAP7_75t_L g82 ( 
.A(n_34),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_25),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_83),
.B(n_86),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_26),
.B(n_4),
.Y(n_84)
);

INVx5_ASAP7_75t_L g85 ( 
.A(n_25),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_85),
.B(n_87),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_31),
.Y(n_86)
);

BUFx12f_ASAP7_75t_L g87 ( 
.A(n_34),
.Y(n_87)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_46),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_88),
.B(n_92),
.Y(n_118)
);

INVx11_ASAP7_75t_L g89 ( 
.A(n_34),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_89),
.A2(n_32),
.B1(n_33),
.B2(n_24),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_31),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_90),
.B(n_91),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_38),
.Y(n_91)
);

INVx8_ASAP7_75t_L g92 ( 
.A(n_18),
.Y(n_92)
);

BUFx2_ASAP7_75t_L g161 ( 
.A(n_94),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_L g95 ( 
.A1(n_91),
.A2(n_28),
.B1(n_45),
.B2(n_18),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_95),
.A2(n_101),
.B1(n_106),
.B2(n_110),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_75),
.A2(n_28),
.B1(n_45),
.B2(n_39),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_49),
.B(n_40),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g149 ( 
.A(n_102),
.B(n_121),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_80),
.A2(n_39),
.B1(n_41),
.B2(n_36),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_55),
.A2(n_41),
.B1(n_33),
.B2(n_24),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_L g116 ( 
.A1(n_47),
.A2(n_22),
.B1(n_36),
.B2(n_32),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_116),
.A2(n_124),
.B1(n_140),
.B2(n_101),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_77),
.A2(n_42),
.B1(n_44),
.B2(n_19),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_119),
.A2(n_127),
.B1(n_61),
.B2(n_65),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_84),
.B(n_46),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_82),
.A2(n_23),
.B1(n_22),
.B2(n_40),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_57),
.A2(n_23),
.B1(n_6),
.B2(n_9),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_92),
.B(n_4),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g158 ( 
.A(n_128),
.B(n_129),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_74),
.B(n_4),
.Y(n_129)
);

FAx1_ASAP7_75t_L g133 ( 
.A(n_79),
.B(n_6),
.CI(n_9),
.CON(n_133),
.SN(n_133)
);

AOI21xp5_ASAP7_75t_L g155 ( 
.A1(n_133),
.A2(n_104),
.B(n_140),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_69),
.B(n_9),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g168 ( 
.A(n_137),
.B(n_138),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_63),
.B(n_10),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_87),
.A2(n_10),
.B1(n_13),
.B2(n_14),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_73),
.B(n_90),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_142),
.B(n_86),
.Y(n_147)
);

INVx3_ASAP7_75t_L g144 ( 
.A(n_136),
.Y(n_144)
);

BUFx4f_ASAP7_75t_SL g196 ( 
.A(n_144),
.Y(n_196)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_118),
.Y(n_145)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_145),
.Y(n_213)
);

INVx5_ASAP7_75t_L g146 ( 
.A(n_136),
.Y(n_146)
);

INVx3_ASAP7_75t_L g189 ( 
.A(n_146),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_147),
.B(n_166),
.Y(n_195)
);

AND2x2_ASAP7_75t_L g148 ( 
.A(n_109),
.B(n_52),
.Y(n_148)
);

AND2x2_ASAP7_75t_L g208 ( 
.A(n_148),
.B(n_155),
.Y(n_208)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_93),
.Y(n_150)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_150),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_97),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_151),
.B(n_160),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_107),
.B(n_64),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_152),
.B(n_182),
.Y(n_200)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_125),
.Y(n_153)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_153),
.Y(n_188)
);

AOI22xp33_ASAP7_75t_SL g154 ( 
.A1(n_133),
.A2(n_83),
.B1(n_58),
.B2(n_59),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_SL g205 ( 
.A1(n_154),
.A2(n_176),
.B1(n_177),
.B2(n_178),
.Y(n_205)
);

INVx4_ASAP7_75t_L g156 ( 
.A(n_141),
.Y(n_156)
);

INVx3_ASAP7_75t_L g199 ( 
.A(n_156),
.Y(n_199)
);

INVx6_ASAP7_75t_L g157 ( 
.A(n_111),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g197 ( 
.A(n_157),
.Y(n_197)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_113),
.Y(n_162)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_162),
.Y(n_192)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_113),
.Y(n_163)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_163),
.Y(n_194)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_93),
.Y(n_164)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_164),
.Y(n_217)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_132),
.Y(n_165)
);

INVx3_ASAP7_75t_L g210 ( 
.A(n_165),
.Y(n_210)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_132),
.Y(n_166)
);

CKINVDCx14_ASAP7_75t_R g167 ( 
.A(n_136),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_167),
.B(n_170),
.Y(n_198)
);

HB1xp67_ASAP7_75t_L g169 ( 
.A(n_123),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_169),
.Y(n_186)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_143),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_98),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_171),
.B(n_172),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_99),
.B(n_66),
.C(n_51),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_135),
.Y(n_173)
);

NOR2x1_ASAP7_75t_L g202 ( 
.A(n_173),
.B(n_181),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_96),
.B(n_119),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_SL g203 ( 
.A(n_174),
.B(n_184),
.Y(n_203)
);

INVx6_ASAP7_75t_L g175 ( 
.A(n_111),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_175),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_127),
.A2(n_133),
.B1(n_103),
.B2(n_106),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_SL g178 ( 
.A1(n_130),
.A2(n_105),
.B1(n_131),
.B2(n_100),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_115),
.A2(n_122),
.B1(n_139),
.B2(n_126),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_179),
.A2(n_175),
.B1(n_157),
.B2(n_161),
.Y(n_209)
);

INVx4_ASAP7_75t_L g180 ( 
.A(n_141),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_SL g216 ( 
.A1(n_180),
.A2(n_183),
.B1(n_185),
.B2(n_146),
.Y(n_216)
);

CKINVDCx16_ASAP7_75t_R g181 ( 
.A(n_117),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_110),
.B(n_124),
.Y(n_182)
);

HB1xp67_ASAP7_75t_L g183 ( 
.A(n_114),
.Y(n_183)
);

OAI211xp5_ASAP7_75t_L g184 ( 
.A1(n_94),
.A2(n_134),
.B(n_143),
.C(n_131),
.Y(n_184)
);

INVx8_ASAP7_75t_L g185 ( 
.A(n_134),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_155),
.A2(n_122),
.B1(n_126),
.B2(n_115),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_191),
.A2(n_193),
.B1(n_204),
.B2(n_207),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_152),
.A2(n_139),
.B1(n_120),
.B2(n_108),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_177),
.B(n_120),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_201),
.B(n_211),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_182),
.A2(n_108),
.B1(n_112),
.B2(n_134),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_SL g206 ( 
.A(n_149),
.B(n_112),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_206),
.B(n_196),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_161),
.A2(n_160),
.B1(n_148),
.B2(n_159),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_209),
.A2(n_214),
.B1(n_193),
.B2(n_191),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_148),
.B(n_168),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_179),
.A2(n_170),
.B1(n_165),
.B2(n_166),
.Y(n_214)
);

INVxp67_ASAP7_75t_L g218 ( 
.A(n_216),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_217),
.Y(n_219)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_219),
.Y(n_242)
);

INVxp67_ASAP7_75t_L g222 ( 
.A(n_198),
.Y(n_222)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_222),
.Y(n_241)
);

NOR2x1_ASAP7_75t_L g223 ( 
.A(n_208),
.B(n_172),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_223),
.B(n_224),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_200),
.B(n_158),
.Y(n_224)
);

HB1xp67_ASAP7_75t_L g225 ( 
.A(n_210),
.Y(n_225)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_225),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_212),
.B(n_150),
.C(n_156),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_226),
.B(n_227),
.C(n_233),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_200),
.B(n_208),
.C(n_201),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_217),
.Y(n_228)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_228),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_205),
.A2(n_180),
.B1(n_144),
.B2(n_185),
.Y(n_229)
);

AND2x2_ASAP7_75t_L g254 ( 
.A(n_229),
.B(n_235),
.Y(n_254)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_187),
.Y(n_230)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_230),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_213),
.B(n_202),
.Y(n_231)
);

CKINVDCx16_ASAP7_75t_R g250 ( 
.A(n_231),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_195),
.B(n_215),
.Y(n_232)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_232),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_208),
.B(n_211),
.C(n_207),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_202),
.B(n_186),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_234),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_192),
.B(n_194),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_188),
.B(n_210),
.Y(n_236)
);

MAJx2_ASAP7_75t_L g256 ( 
.A(n_236),
.B(n_192),
.C(n_187),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_197),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_L g251 ( 
.A1(n_237),
.A2(n_238),
.B1(n_239),
.B2(n_240),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_L g239 ( 
.A1(n_203),
.A2(n_190),
.B1(n_204),
.B2(n_197),
.Y(n_239)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_219),
.Y(n_249)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_249),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_220),
.A2(n_214),
.B1(n_188),
.B2(n_194),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_252),
.B(n_236),
.Y(n_263)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_228),
.Y(n_255)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_255),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_SL g259 ( 
.A(n_256),
.B(n_227),
.Y(n_259)
);

A2O1A1Ixp33_ASAP7_75t_L g257 ( 
.A1(n_245),
.A2(n_233),
.B(n_224),
.C(n_220),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_257),
.B(n_258),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_252),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_259),
.B(n_243),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_SL g262 ( 
.A(n_245),
.B(n_232),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_262),
.B(n_264),
.C(n_256),
.Y(n_277)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_263),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_243),
.B(n_223),
.C(n_226),
.Y(n_264)
);

A2O1A1Ixp33_ASAP7_75t_L g265 ( 
.A1(n_248),
.A2(n_223),
.B(n_222),
.C(n_229),
.Y(n_265)
);

OAI21xp5_ASAP7_75t_L g279 ( 
.A1(n_265),
.A2(n_255),
.B(n_249),
.Y(n_279)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_246),
.Y(n_266)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_266),
.Y(n_271)
);

OAI322xp33_ASAP7_75t_L g267 ( 
.A1(n_248),
.A2(n_230),
.A3(n_237),
.B1(n_239),
.B2(n_196),
.C1(n_221),
.C2(n_218),
.Y(n_267)
);

NOR3xp33_ASAP7_75t_SL g275 ( 
.A(n_267),
.B(n_241),
.C(n_247),
.Y(n_275)
);

AOI21xp5_ASAP7_75t_L g268 ( 
.A1(n_254),
.A2(n_218),
.B(n_221),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_SL g276 ( 
.A1(n_268),
.A2(n_269),
.B(n_247),
.Y(n_276)
);

AOI21xp5_ASAP7_75t_L g269 ( 
.A1(n_254),
.A2(n_238),
.B(n_189),
.Y(n_269)
);

AOI21xp5_ASAP7_75t_SL g272 ( 
.A1(n_263),
.A2(n_251),
.B(n_254),
.Y(n_272)
);

OAI21xp5_ASAP7_75t_L g280 ( 
.A1(n_272),
.A2(n_275),
.B(n_276),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_273),
.B(n_274),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_L g274 ( 
.A1(n_269),
.A2(n_253),
.B1(n_241),
.B2(n_250),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_277),
.B(n_279),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_277),
.B(n_264),
.C(n_259),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_281),
.B(n_272),
.C(n_270),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_SL g283 ( 
.A(n_278),
.B(n_262),
.Y(n_283)
);

OR2x2_ASAP7_75t_L g291 ( 
.A(n_283),
.B(n_285),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_SL g285 ( 
.A(n_271),
.B(n_257),
.Y(n_285)
);

AOI321xp33_ASAP7_75t_L g286 ( 
.A1(n_279),
.A2(n_261),
.A3(n_260),
.B1(n_265),
.B2(n_246),
.C(n_242),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_286),
.B(n_275),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_287),
.B(n_199),
.C(n_289),
.Y(n_294)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_288),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_284),
.B(n_244),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_289),
.B(n_292),
.Y(n_295)
);

O2A1O1Ixp33_ASAP7_75t_L g290 ( 
.A1(n_280),
.A2(n_276),
.B(n_268),
.C(n_244),
.Y(n_290)
);

AOI22xp33_ASAP7_75t_SL g293 ( 
.A1(n_290),
.A2(n_282),
.B1(n_281),
.B2(n_189),
.Y(n_293)
);

AO21x1_ASAP7_75t_L g292 ( 
.A1(n_282),
.A2(n_196),
.B(n_199),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_293),
.B(n_294),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_293),
.B(n_291),
.C(n_292),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_297),
.B(n_299),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_296),
.B(n_295),
.Y(n_298)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_298),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_300),
.B(n_297),
.Y(n_302)
);

OR2x2_ASAP7_75t_L g303 ( 
.A(n_302),
.B(n_301),
.Y(n_303)
);


endmodule