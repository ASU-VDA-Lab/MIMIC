module real_jpeg_1508_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_176;
wire n_104;
wire n_153;
wire n_161;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_164;
wire n_48;
wire n_140;
wire n_126;
wire n_113;
wire n_120;
wire n_155;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_170;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_172;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_100;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_30;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_185;
wire n_55;
wire n_180;
wire n_58;
wire n_52;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_187;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_179;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_0),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_1),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g44 ( 
.A1(n_2),
.A2(n_36),
.B1(n_42),
.B2(n_45),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_2),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_3),
.A2(n_24),
.B1(n_25),
.B2(n_57),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_3),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_3),
.A2(n_30),
.B1(n_32),
.B2(n_57),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_3),
.A2(n_50),
.B1(n_51),
.B2(n_57),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_3),
.A2(n_36),
.B1(n_42),
.B2(n_57),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_4),
.A2(n_36),
.B1(n_42),
.B2(n_108),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_4),
.Y(n_108)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_5),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_6),
.A2(n_24),
.B1(n_25),
.B2(n_60),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_6),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_6),
.A2(n_30),
.B1(n_32),
.B2(n_60),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_6),
.A2(n_50),
.B1(n_51),
.B2(n_60),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_6),
.A2(n_36),
.B1(n_42),
.B2(n_60),
.Y(n_170)
);

BUFx8_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_8),
.B(n_32),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_8),
.B(n_63),
.Y(n_62)
);

AOI21xp5_ASAP7_75t_L g74 ( 
.A1(n_8),
.A2(n_31),
.B(n_32),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_8),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_8),
.B(n_49),
.Y(n_138)
);

AOI21xp33_ASAP7_75t_L g145 ( 
.A1(n_8),
.A2(n_24),
.B(n_146),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_8),
.B(n_36),
.C(n_85),
.Y(n_154)
);

OAI22xp33_ASAP7_75t_SL g157 ( 
.A1(n_8),
.A2(n_50),
.B1(n_51),
.B2(n_125),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_8),
.B(n_39),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_8),
.B(n_90),
.Y(n_168)
);

BUFx16f_ASAP7_75t_L g85 ( 
.A(n_9),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_11),
.A2(n_50),
.B1(n_51),
.B2(n_82),
.Y(n_81)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_11),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_11),
.A2(n_24),
.B1(n_25),
.B2(n_82),
.Y(n_102)
);

OAI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_11),
.A2(n_36),
.B1(n_42),
.B2(n_82),
.Y(n_129)
);

OAI22xp33_ASAP7_75t_L g67 ( 
.A1(n_12),
.A2(n_36),
.B1(n_42),
.B2(n_68),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_12),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_12),
.A2(n_50),
.B1(n_51),
.B2(n_68),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_L g40 ( 
.A1(n_14),
.A2(n_36),
.B1(n_41),
.B2(n_42),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_14),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_L g111 ( 
.A1(n_14),
.A2(n_41),
.B1(n_50),
.B2(n_51),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_15),
.A2(n_24),
.B1(n_25),
.B2(n_79),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_15),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_15),
.A2(n_50),
.B1(n_51),
.B2(n_79),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_15),
.A2(n_36),
.B1(n_42),
.B2(n_79),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_16),
.Y(n_52)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

OAI22xp5_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_114),
.B1(n_186),
.B2(n_187),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_19),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_113),
.Y(n_19)
);

OR2x2_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_93),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_21),
.B(n_93),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_21),
.B(n_116),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_21),
.B(n_116),
.Y(n_185)
);

FAx1_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_46),
.CI(n_69),
.CON(n_21),
.SN(n_21)
);

XNOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_34),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_23),
.B(n_34),
.Y(n_95)
);

AOI32xp33_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_27),
.A3(n_30),
.B1(n_31),
.B2(n_33),
.Y(n_23)
);

AOI22xp33_ASAP7_75t_L g55 ( 
.A1(n_24),
.A2(n_25),
.B1(n_53),
.B2(n_54),
.Y(n_55)
);

OA22x2_ASAP7_75t_L g64 ( 
.A1(n_24),
.A2(n_25),
.B1(n_27),
.B2(n_28),
.Y(n_64)
);

OAI32xp33_ASAP7_75t_L g123 ( 
.A1(n_24),
.A2(n_51),
.A3(n_53),
.B1(n_124),
.B2(n_126),
.Y(n_123)
);

INVx8_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

NAND2xp33_ASAP7_75t_SL g33 ( 
.A(n_25),
.B(n_28),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_25),
.B(n_125),
.Y(n_124)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_27),
.A2(n_28),
.B1(n_30),
.B2(n_32),
.Y(n_73)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

BUFx4f_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_30),
.Y(n_32)
);

AOI22xp5_ASAP7_75t_L g34 ( 
.A1(n_35),
.A2(n_39),
.B1(n_40),
.B2(n_43),
.Y(n_34)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_35),
.A2(n_39),
.B1(n_40),
.B2(n_67),
.Y(n_66)
);

INVx1_ASAP7_75t_SL g106 ( 
.A(n_35),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_35),
.A2(n_39),
.B1(n_129),
.B2(n_140),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_35),
.A2(n_39),
.B1(n_125),
.B2(n_166),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_35),
.A2(n_39),
.B1(n_166),
.B2(n_170),
.Y(n_169)
);

AND2x2_ASAP7_75t_L g35 ( 
.A(n_36),
.B(n_38),
.Y(n_35)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_36),
.Y(n_42)
);

OA22x2_ASAP7_75t_L g87 ( 
.A1(n_36),
.A2(n_42),
.B1(n_85),
.B2(n_86),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_36),
.B(n_164),
.Y(n_163)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_38),
.A2(n_44),
.B1(n_106),
.B2(n_107),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_38),
.A2(n_106),
.B1(n_128),
.B2(n_130),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_38),
.A2(n_106),
.B1(n_174),
.B2(n_175),
.Y(n_173)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

MAJIxp5_ASAP7_75t_L g46 ( 
.A(n_47),
.B(n_61),
.C(n_65),
.Y(n_46)
);

XOR2xp5_ASAP7_75t_L g117 ( 
.A(n_47),
.B(n_118),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g47 ( 
.A1(n_48),
.A2(n_56),
.B1(n_58),
.B2(n_59),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_48),
.A2(n_58),
.B1(n_59),
.B2(n_78),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_48),
.A2(n_58),
.B1(n_78),
.B2(n_101),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_48),
.A2(n_56),
.B1(n_58),
.B2(n_145),
.Y(n_144)
);

OR2x2_ASAP7_75t_L g48 ( 
.A(n_49),
.B(n_55),
.Y(n_48)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_49),
.Y(n_58)
);

AO22x2_ASAP7_75t_SL g49 ( 
.A1(n_50),
.A2(n_51),
.B1(n_53),
.B2(n_54),
.Y(n_49)
);

OAI22xp33_ASAP7_75t_L g84 ( 
.A1(n_50),
.A2(n_51),
.B1(n_85),
.B2(n_86),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_50),
.B(n_54),
.Y(n_126)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_51),
.B(n_154),
.Y(n_153)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx3_ASAP7_75t_SL g54 ( 
.A(n_53),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_61),
.A2(n_62),
.B1(n_65),
.B2(n_66),
.Y(n_118)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_64),
.A2(n_71),
.B1(n_74),
.B2(n_75),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_64),
.B(n_73),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_64),
.A2(n_71),
.B1(n_75),
.B2(n_98),
.Y(n_97)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_67),
.Y(n_130)
);

XOR2xp5_ASAP7_75t_L g69 ( 
.A(n_70),
.B(n_76),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_70),
.B(n_77),
.C(n_92),
.Y(n_112)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_77),
.A2(n_80),
.B1(n_91),
.B2(n_92),
.Y(n_76)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_77),
.Y(n_91)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_80),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_81),
.A2(n_83),
.B1(n_88),
.B2(n_90),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_81),
.A2(n_83),
.B1(n_90),
.B2(n_120),
.Y(n_119)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_83),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_83),
.A2(n_90),
.B1(n_136),
.B2(n_137),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_83),
.A2(n_90),
.B1(n_136),
.B2(n_157),
.Y(n_156)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_87),
.Y(n_83)
);

INVx11_ASAP7_75t_L g86 ( 
.A(n_85),
.Y(n_86)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_87),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_87),
.A2(n_89),
.B1(n_110),
.B2(n_111),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_87),
.A2(n_110),
.B1(n_121),
.B2(n_148),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

XNOR2xp5_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_103),
.Y(n_93)
);

XNOR2xp5_ASAP7_75t_SL g94 ( 
.A(n_95),
.B(n_96),
.Y(n_94)
);

XOR2xp5_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_100),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

CKINVDCx14_ASAP7_75t_R g101 ( 
.A(n_102),
.Y(n_101)
);

XOR2xp5_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_112),
.Y(n_103)
);

XNOR2xp5_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_109),
.Y(n_104)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_114),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_L g114 ( 
.A1(n_115),
.A2(n_131),
.B(n_185),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_119),
.C(n_122),
.Y(n_116)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_117),
.B(n_182),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_119),
.B(n_122),
.Y(n_182)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_127),
.Y(n_122)
);

XOR2xp5_ASAP7_75t_L g142 ( 
.A(n_123),
.B(n_127),
.Y(n_142)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_124),
.Y(n_146)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

AOI21xp5_ASAP7_75t_SL g131 ( 
.A1(n_132),
.A2(n_180),
.B(n_184),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_L g132 ( 
.A1(n_133),
.A2(n_149),
.B(n_179),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_141),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_134),
.B(n_141),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_138),
.C(n_139),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_135),
.B(n_138),
.Y(n_159)
);

INVxp67_ASAP7_75t_L g148 ( 
.A(n_137),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_139),
.B(n_159),
.Y(n_158)
);

INVxp67_ASAP7_75t_L g175 ( 
.A(n_140),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_143),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_142),
.B(n_144),
.C(n_147),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_147),
.Y(n_143)
);

AOI21xp5_ASAP7_75t_L g149 ( 
.A1(n_150),
.A2(n_160),
.B(n_178),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_158),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_151),
.B(n_158),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_155),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_152),
.A2(n_153),
.B1(n_155),
.B2(n_156),
.Y(n_176)
);

CKINVDCx16_ASAP7_75t_R g152 ( 
.A(n_153),
.Y(n_152)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_L g160 ( 
.A1(n_161),
.A2(n_172),
.B(n_177),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_L g161 ( 
.A1(n_162),
.A2(n_167),
.B(n_171),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_165),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_168),
.B(n_169),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_168),
.B(n_169),
.Y(n_171)
);

INVxp67_ASAP7_75t_L g174 ( 
.A(n_170),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_173),
.B(n_176),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_173),
.B(n_176),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_181),
.B(n_183),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_181),
.B(n_183),
.Y(n_184)
);


endmodule