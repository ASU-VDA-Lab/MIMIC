module fake_jpeg_13052_n_375 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_375);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_375;

wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_10),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_13),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_7),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_4),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_8),
.Y(n_21)
);

CKINVDCx16_ASAP7_75t_R g22 ( 
.A(n_9),
.Y(n_22)
);

BUFx16f_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_1),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_2),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_8),
.Y(n_27)
);

BUFx16f_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_13),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_11),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_5),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_8),
.Y(n_36)
);

BUFx4f_ASAP7_75t_L g37 ( 
.A(n_4),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_9),
.Y(n_38)
);

INVx13_ASAP7_75t_L g39 ( 
.A(n_2),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_6),
.Y(n_40)
);

INVx1_ASAP7_75t_SL g41 ( 
.A(n_0),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_15),
.Y(n_42)
);

INVx6_ASAP7_75t_L g102 ( 
.A(n_42),
.Y(n_102)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_23),
.Y(n_43)
);

INVx2_ASAP7_75t_SL g127 ( 
.A(n_43),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_15),
.Y(n_44)
);

BUFx2_ASAP7_75t_L g128 ( 
.A(n_44),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_15),
.Y(n_45)
);

INVx5_ASAP7_75t_L g103 ( 
.A(n_45),
.Y(n_103)
);

INVx2_ASAP7_75t_SL g46 ( 
.A(n_26),
.Y(n_46)
);

INVx5_ASAP7_75t_SL g112 ( 
.A(n_46),
.Y(n_112)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_26),
.Y(n_47)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_47),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_15),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g104 ( 
.A(n_48),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_17),
.Y(n_49)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_49),
.Y(n_121)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_26),
.Y(n_50)
);

INVx4_ASAP7_75t_L g122 ( 
.A(n_50),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_16),
.B(n_12),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_51),
.B(n_54),
.Y(n_117)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_29),
.Y(n_52)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_52),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_36),
.B(n_0),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_53),
.B(n_77),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_16),
.B(n_12),
.Y(n_54)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_20),
.Y(n_55)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_55),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_17),
.Y(n_56)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_56),
.Y(n_106)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_17),
.Y(n_57)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_57),
.Y(n_118)
);

INVx6_ASAP7_75t_SL g58 ( 
.A(n_23),
.Y(n_58)
);

CKINVDCx16_ASAP7_75t_R g126 ( 
.A(n_58),
.Y(n_126)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_30),
.Y(n_59)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_59),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_32),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_60),
.B(n_62),
.Y(n_82)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_30),
.Y(n_61)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_61),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_32),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_17),
.Y(n_63)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_63),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_23),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_64),
.B(n_66),
.Y(n_83)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_23),
.Y(n_65)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_65),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_23),
.Y(n_66)
);

INVx11_ASAP7_75t_L g67 ( 
.A(n_39),
.Y(n_67)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_67),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_28),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_68),
.B(n_70),
.Y(n_95)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_30),
.Y(n_69)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_69),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_31),
.B(n_12),
.Y(n_70)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_36),
.Y(n_71)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_71),
.B(n_73),
.Y(n_97)
);

INVx6_ASAP7_75t_SL g72 ( 
.A(n_28),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_72),
.B(n_74),
.Y(n_108)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_36),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_28),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_28),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_75),
.B(n_76),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_33),
.Y(n_76)
);

HB1xp67_ASAP7_75t_L g77 ( 
.A(n_20),
.Y(n_77)
);

BUFx12f_ASAP7_75t_L g78 ( 
.A(n_20),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_78),
.A2(n_39),
.B1(n_35),
.B2(n_22),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_28),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_79),
.B(n_80),
.Y(n_86)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_37),
.Y(n_80)
);

BUFx5_ASAP7_75t_L g81 ( 
.A(n_33),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_81),
.B(n_41),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_L g87 ( 
.A1(n_57),
.A2(n_33),
.B1(n_40),
.B2(n_24),
.Y(n_87)
);

OAI22xp33_ASAP7_75t_L g170 ( 
.A1(n_87),
.A2(n_88),
.B1(n_115),
.B2(n_123),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_L g88 ( 
.A1(n_42),
.A2(n_33),
.B1(n_40),
.B2(n_24),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_53),
.A2(n_34),
.B1(n_41),
.B2(n_29),
.Y(n_89)
);

OA22x2_ASAP7_75t_L g148 ( 
.A1(n_89),
.A2(n_69),
.B1(n_72),
.B2(n_81),
.Y(n_148)
);

INVxp67_ASAP7_75t_L g140 ( 
.A(n_90),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_71),
.B(n_38),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_91),
.B(n_101),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_60),
.A2(n_31),
.B1(n_38),
.B2(n_27),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_94),
.A2(n_99),
.B1(n_111),
.B2(n_124),
.Y(n_160)
);

OAI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_73),
.A2(n_41),
.B1(n_34),
.B2(n_35),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_52),
.B(n_18),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_66),
.B(n_34),
.C(n_35),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_105),
.B(n_7),
.C(n_97),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_79),
.B(n_18),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_107),
.B(n_114),
.Y(n_135)
);

AOI21xp5_ASAP7_75t_L g156 ( 
.A1(n_110),
.A2(n_4),
.B(n_5),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_62),
.A2(n_27),
.B1(n_25),
.B2(n_21),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_80),
.B(n_25),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_L g115 ( 
.A1(n_44),
.A2(n_21),
.B1(n_19),
.B2(n_22),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_46),
.A2(n_19),
.B1(n_39),
.B2(n_37),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_119),
.A2(n_129),
.B1(n_67),
.B2(n_59),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_L g123 ( 
.A1(n_45),
.A2(n_37),
.B1(n_39),
.B2(n_2),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_48),
.A2(n_37),
.B1(n_10),
.B2(n_2),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_49),
.A2(n_37),
.B1(n_10),
.B2(n_3),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_125),
.A2(n_61),
.B1(n_47),
.B2(n_55),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_46),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_129)
);

BUFx2_ASAP7_75t_L g130 ( 
.A(n_112),
.Y(n_130)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_130),
.Y(n_183)
);

INVx4_ASAP7_75t_L g132 ( 
.A(n_93),
.Y(n_132)
);

BUFx2_ASAP7_75t_L g189 ( 
.A(n_132),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_82),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_133),
.B(n_150),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_117),
.B(n_43),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g193 ( 
.A(n_134),
.B(n_137),
.Y(n_193)
);

AOI22xp33_ASAP7_75t_L g136 ( 
.A1(n_125),
.A2(n_63),
.B1(n_76),
.B2(n_56),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_136),
.A2(n_145),
.B1(n_122),
.B2(n_127),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_95),
.B(n_78),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_84),
.B(n_65),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_138),
.B(n_141),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g139 ( 
.A(n_84),
.B(n_58),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_139),
.B(n_168),
.C(n_141),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_91),
.B(n_0),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_SL g179 ( 
.A1(n_142),
.A2(n_172),
.B1(n_175),
.B2(n_122),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_83),
.B(n_78),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_143),
.B(n_149),
.Y(n_203)
);

BUFx12f_ASAP7_75t_L g144 ( 
.A(n_112),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g198 ( 
.A(n_144),
.Y(n_198)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_118),
.Y(n_146)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_146),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_114),
.B(n_1),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_147),
.B(n_154),
.Y(n_197)
);

AND2x2_ASAP7_75t_L g196 ( 
.A(n_148),
.B(n_161),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_107),
.B(n_50),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_101),
.B(n_50),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_108),
.B(n_1),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_151),
.B(n_152),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_86),
.Y(n_152)
);

OR2x2_ASAP7_75t_L g153 ( 
.A(n_89),
.B(n_3),
.Y(n_153)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_153),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_86),
.B(n_3),
.Y(n_154)
);

INVx6_ASAP7_75t_L g155 ( 
.A(n_102),
.Y(n_155)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_155),
.Y(n_195)
);

AOI21xp5_ASAP7_75t_L g209 ( 
.A1(n_156),
.A2(n_165),
.B(n_139),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_92),
.B(n_4),
.Y(n_157)
);

CKINVDCx14_ASAP7_75t_R g188 ( 
.A(n_157),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_92),
.B(n_5),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_158),
.B(n_166),
.Y(n_202)
);

INVx3_ASAP7_75t_L g159 ( 
.A(n_93),
.Y(n_159)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_159),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_105),
.B(n_113),
.Y(n_161)
);

INVx3_ASAP7_75t_L g162 ( 
.A(n_104),
.Y(n_162)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_162),
.Y(n_180)
);

BUFx8_ASAP7_75t_L g163 ( 
.A(n_126),
.Y(n_163)
);

INVx13_ASAP7_75t_L g194 ( 
.A(n_163),
.Y(n_194)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_97),
.Y(n_164)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_164),
.Y(n_181)
);

A2O1A1Ixp33_ASAP7_75t_L g165 ( 
.A1(n_90),
.A2(n_5),
.B(n_6),
.C(n_7),
.Y(n_165)
);

A2O1A1Ixp33_ASAP7_75t_L g187 ( 
.A1(n_165),
.A2(n_127),
.B(n_109),
.C(n_85),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_97),
.B(n_6),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_96),
.B(n_6),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_167),
.Y(n_182)
);

INVx1_ASAP7_75t_SL g169 ( 
.A(n_98),
.Y(n_169)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_169),
.Y(n_204)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_127),
.Y(n_171)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_171),
.Y(n_206)
);

AOI22xp33_ASAP7_75t_SL g172 ( 
.A1(n_85),
.A2(n_109),
.B1(n_120),
.B2(n_116),
.Y(n_172)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_118),
.Y(n_173)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_173),
.Y(n_207)
);

OAI22xp33_ASAP7_75t_SL g174 ( 
.A1(n_106),
.A2(n_121),
.B1(n_128),
.B2(n_100),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_174),
.A2(n_104),
.B1(n_130),
.B2(n_170),
.Y(n_192)
);

INVx6_ASAP7_75t_L g175 ( 
.A(n_102),
.Y(n_175)
);

AND2x2_ASAP7_75t_L g248 ( 
.A(n_176),
.B(n_192),
.Y(n_248)
);

INVxp67_ASAP7_75t_L g229 ( 
.A(n_179),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_160),
.A2(n_100),
.B1(n_106),
.B2(n_121),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_186),
.A2(n_190),
.B1(n_191),
.B2(n_208),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_187),
.B(n_211),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_160),
.A2(n_103),
.B1(n_128),
.B2(n_120),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_138),
.A2(n_103),
.B1(n_104),
.B2(n_140),
.Y(n_191)
);

INVx13_ASAP7_75t_L g199 ( 
.A(n_163),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_199),
.Y(n_236)
);

AND2x6_ASAP7_75t_L g200 ( 
.A(n_135),
.B(n_131),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_200),
.B(n_196),
.Y(n_216)
);

INVx13_ASAP7_75t_L g201 ( 
.A(n_163),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_201),
.Y(n_220)
);

AOI22xp33_ASAP7_75t_L g205 ( 
.A1(n_170),
.A2(n_164),
.B1(n_140),
.B2(n_148),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_205),
.A2(n_156),
.B1(n_144),
.B2(n_132),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_131),
.A2(n_135),
.B1(n_153),
.B2(n_145),
.Y(n_208)
);

AOI21xp5_ASAP7_75t_L g237 ( 
.A1(n_209),
.A2(n_187),
.B(n_203),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_210),
.B(n_162),
.C(n_144),
.Y(n_218)
);

AO22x1_ASAP7_75t_SL g211 ( 
.A1(n_148),
.A2(n_154),
.B1(n_169),
.B2(n_168),
.Y(n_211)
);

OAI22xp33_ASAP7_75t_SL g214 ( 
.A1(n_148),
.A2(n_147),
.B1(n_158),
.B2(n_159),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_214),
.A2(n_181),
.B1(n_210),
.B2(n_211),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_146),
.B(n_173),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_215),
.B(n_207),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_216),
.B(n_239),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_217),
.A2(n_233),
.B1(n_248),
.B2(n_219),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_218),
.B(n_241),
.Y(n_257)
);

OAI21xp5_ASAP7_75t_L g219 ( 
.A1(n_209),
.A2(n_155),
.B(n_175),
.Y(n_219)
);

AOI21xp5_ASAP7_75t_SL g264 ( 
.A1(n_219),
.A2(n_221),
.B(n_244),
.Y(n_264)
);

OAI21xp5_ASAP7_75t_L g221 ( 
.A1(n_196),
.A2(n_213),
.B(n_193),
.Y(n_221)
);

AOI22xp33_ASAP7_75t_SL g223 ( 
.A1(n_186),
.A2(n_213),
.B1(n_191),
.B2(n_183),
.Y(n_223)
);

INVxp67_ASAP7_75t_L g275 ( 
.A(n_223),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_196),
.A2(n_211),
.B1(n_178),
.B2(n_181),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_225),
.A2(n_231),
.B1(n_222),
.B2(n_230),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_226),
.B(n_230),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_215),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_227),
.B(n_228),
.Y(n_259)
);

BUFx24_ASAP7_75t_SL g228 ( 
.A(n_177),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_178),
.B(n_197),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_182),
.B(n_188),
.Y(n_232)
);

CKINVDCx14_ASAP7_75t_R g265 ( 
.A(n_232),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_200),
.A2(n_192),
.B1(n_197),
.B2(n_202),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_202),
.B(n_185),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_234),
.B(n_243),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_206),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_235),
.B(n_242),
.Y(n_263)
);

OAI21xp5_ASAP7_75t_SL g273 ( 
.A1(n_237),
.A2(n_246),
.B(n_247),
.Y(n_273)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_206),
.Y(n_238)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_238),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_182),
.B(n_204),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_207),
.Y(n_240)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_240),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_204),
.B(n_180),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_SL g277 ( 
.A(n_241),
.B(n_248),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_184),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_183),
.B(n_184),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_L g244 ( 
.A1(n_198),
.A2(n_180),
.B(n_212),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_212),
.B(n_189),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_245),
.B(n_235),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_195),
.A2(n_189),
.B1(n_198),
.B2(n_194),
.Y(n_246)
);

AO22x1_ASAP7_75t_L g247 ( 
.A1(n_195),
.A2(n_194),
.B1(n_199),
.B2(n_201),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_249),
.A2(n_255),
.B1(n_264),
.B2(n_275),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_236),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_251),
.B(n_256),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_253),
.B(n_254),
.Y(n_282)
);

INVx1_ASAP7_75t_SL g254 ( 
.A(n_236),
.Y(n_254)
);

OR2x2_ASAP7_75t_L g255 ( 
.A(n_224),
.B(n_225),
.Y(n_255)
);

NAND2xp33_ASAP7_75t_SL g293 ( 
.A(n_255),
.B(n_268),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_243),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_257),
.B(n_252),
.C(n_277),
.Y(n_291)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_238),
.Y(n_260)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_260),
.Y(n_300)
);

OAI21xp5_ASAP7_75t_L g261 ( 
.A1(n_237),
.A2(n_224),
.B(n_221),
.Y(n_261)
);

OAI21xp5_ASAP7_75t_L g285 ( 
.A1(n_261),
.A2(n_267),
.B(n_220),
.Y(n_285)
);

OAI21xp5_ASAP7_75t_L g267 ( 
.A1(n_231),
.A2(n_216),
.B(n_233),
.Y(n_267)
);

CKINVDCx16_ASAP7_75t_R g268 ( 
.A(n_239),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_269),
.A2(n_274),
.B1(n_267),
.B2(n_268),
.Y(n_296)
);

OAI21xp33_ASAP7_75t_SL g270 ( 
.A1(n_229),
.A2(n_227),
.B(n_217),
.Y(n_270)
);

BUFx12f_ASAP7_75t_SL g288 ( 
.A(n_270),
.Y(n_288)
);

INVx6_ASAP7_75t_L g271 ( 
.A(n_247),
.Y(n_271)
);

BUFx5_ASAP7_75t_L g278 ( 
.A(n_271),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_234),
.B(n_226),
.Y(n_272)
);

CKINVDCx14_ASAP7_75t_R g279 ( 
.A(n_272),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_222),
.A2(n_248),
.B1(n_218),
.B2(n_232),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_220),
.B(n_240),
.Y(n_276)
);

CKINVDCx16_ASAP7_75t_R g289 ( 
.A(n_276),
.Y(n_289)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_277),
.B(n_244),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_257),
.B(n_247),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_280),
.B(n_283),
.C(n_291),
.Y(n_304)
);

XOR2xp5_ASAP7_75t_L g301 ( 
.A(n_281),
.B(n_285),
.Y(n_301)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_261),
.B(n_245),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_263),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g312 ( 
.A(n_284),
.B(n_299),
.Y(n_312)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_250),
.Y(n_286)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_286),
.Y(n_317)
);

AOI21xp5_ASAP7_75t_L g287 ( 
.A1(n_273),
.A2(n_246),
.B(n_242),
.Y(n_287)
);

HB1xp67_ASAP7_75t_L g315 ( 
.A(n_287),
.Y(n_315)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_250),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_290),
.B(n_292),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_272),
.B(n_262),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_262),
.B(n_266),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_295),
.B(n_298),
.C(n_255),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_L g311 ( 
.A1(n_296),
.A2(n_249),
.B1(n_256),
.B2(n_265),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_297),
.A2(n_274),
.B1(n_275),
.B2(n_264),
.Y(n_305)
);

XOR2xp5_ASAP7_75t_L g298 ( 
.A(n_269),
.B(n_252),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_260),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_SL g303 ( 
.A(n_289),
.B(n_259),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_SL g325 ( 
.A(n_303),
.B(n_306),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_SL g335 ( 
.A1(n_305),
.A2(n_278),
.B1(n_290),
.B2(n_299),
.Y(n_335)
);

CKINVDCx16_ASAP7_75t_R g306 ( 
.A(n_282),
.Y(n_306)
);

BUFx3_ASAP7_75t_L g307 ( 
.A(n_296),
.Y(n_307)
);

HB1xp67_ASAP7_75t_L g331 ( 
.A(n_307),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_SL g329 ( 
.A(n_308),
.B(n_300),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_291),
.B(n_266),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_309),
.B(n_314),
.C(n_298),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_294),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_310),
.B(n_318),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_311),
.Y(n_323)
);

OAI22xp5_ASAP7_75t_L g313 ( 
.A1(n_279),
.A2(n_271),
.B1(n_253),
.B2(n_251),
.Y(n_313)
);

INVxp33_ASAP7_75t_L g324 ( 
.A(n_313),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_280),
.B(n_273),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_L g316 ( 
.A1(n_292),
.A2(n_271),
.B1(n_254),
.B2(n_258),
.Y(n_316)
);

BUFx2_ASAP7_75t_L g328 ( 
.A(n_316),
.Y(n_328)
);

INVx3_ASAP7_75t_SL g318 ( 
.A(n_278),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_L g319 ( 
.A1(n_282),
.A2(n_258),
.B1(n_287),
.B2(n_285),
.Y(n_319)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_319),
.Y(n_333)
);

XOR2xp5_ASAP7_75t_L g342 ( 
.A(n_320),
.B(n_309),
.Y(n_342)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_304),
.B(n_281),
.C(n_283),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_321),
.B(n_304),
.C(n_320),
.Y(n_343)
);

OAI22xp5_ASAP7_75t_L g326 ( 
.A1(n_307),
.A2(n_293),
.B1(n_297),
.B2(n_288),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_L g338 ( 
.A1(n_326),
.A2(n_335),
.B1(n_315),
.B2(n_318),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_310),
.B(n_295),
.Y(n_327)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_327),
.Y(n_336)
);

XNOR2xp5_ASAP7_75t_L g346 ( 
.A(n_329),
.B(n_301),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_303),
.B(n_288),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_330),
.B(n_332),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_312),
.B(n_286),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_302),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_334),
.B(n_302),
.Y(n_345)
);

INVxp67_ASAP7_75t_L g337 ( 
.A(n_322),
.Y(n_337)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_337),
.Y(n_349)
);

XNOR2xp5_ASAP7_75t_L g356 ( 
.A(n_338),
.B(n_342),
.Y(n_356)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_325),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_339),
.B(n_340),
.Y(n_352)
);

HB1xp67_ASAP7_75t_L g340 ( 
.A(n_331),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_324),
.B(n_308),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_341),
.B(n_343),
.Y(n_355)
);

A2O1A1Ixp33_ASAP7_75t_L g348 ( 
.A1(n_345),
.A2(n_327),
.B(n_333),
.C(n_323),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_L g350 ( 
.A(n_346),
.B(n_347),
.Y(n_350)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_322),
.Y(n_347)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_348),
.Y(n_359)
);

AOI21xp5_ASAP7_75t_L g351 ( 
.A1(n_344),
.A2(n_333),
.B(n_323),
.Y(n_351)
);

OAI21xp5_ASAP7_75t_SL g357 ( 
.A1(n_351),
.A2(n_354),
.B(n_337),
.Y(n_357)
);

MAJIxp5_ASAP7_75t_L g353 ( 
.A(n_342),
.B(n_321),
.C(n_335),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_353),
.B(n_343),
.Y(n_358)
);

AOI21xp5_ASAP7_75t_L g354 ( 
.A1(n_346),
.A2(n_305),
.B(n_301),
.Y(n_354)
);

AOI21xp5_ASAP7_75t_L g366 ( 
.A1(n_357),
.A2(n_360),
.B(n_363),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_L g364 ( 
.A(n_358),
.B(n_356),
.Y(n_364)
);

MAJIxp5_ASAP7_75t_L g360 ( 
.A(n_356),
.B(n_338),
.C(n_336),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_L g361 ( 
.A(n_355),
.B(n_328),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_SL g367 ( 
.A(n_361),
.B(n_362),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_L g362 ( 
.A(n_352),
.B(n_328),
.Y(n_362)
);

AOI22xp5_ASAP7_75t_SL g363 ( 
.A1(n_349),
.A2(n_326),
.B1(n_328),
.B2(n_334),
.Y(n_363)
);

INVxp67_ASAP7_75t_L g369 ( 
.A(n_364),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_L g365 ( 
.A(n_360),
.B(n_350),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_L g368 ( 
.A(n_365),
.B(n_359),
.Y(n_368)
);

MAJIxp5_ASAP7_75t_L g372 ( 
.A(n_368),
.B(n_370),
.C(n_314),
.Y(n_372)
);

MAJIxp5_ASAP7_75t_L g370 ( 
.A(n_366),
.B(n_353),
.C(n_363),
.Y(n_370)
);

OA21x2_ASAP7_75t_SL g371 ( 
.A1(n_369),
.A2(n_367),
.B(n_348),
.Y(n_371)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_371),
.Y(n_373)
);

MAJIxp5_ASAP7_75t_L g374 ( 
.A(n_373),
.B(n_372),
.C(n_317),
.Y(n_374)
);

FAx1_ASAP7_75t_SL g375 ( 
.A(n_374),
.B(n_317),
.CI(n_372),
.CON(n_375),
.SN(n_375)
);


endmodule