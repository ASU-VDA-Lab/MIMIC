module fake_netlist_5_1213_n_1719 (n_137, n_91, n_82, n_122, n_142, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_60, n_152, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_125, n_35, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_29, n_79, n_131, n_151, n_47, n_25, n_53, n_8, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_109, n_112, n_85, n_95, n_119, n_59, n_26, n_133, n_55, n_99, n_2, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_27, n_64, n_77, n_102, n_106, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_134, n_32, n_41, n_104, n_103, n_56, n_51, n_63, n_97, n_141, n_11, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_1719);

input n_137;
input n_91;
input n_82;
input n_122;
input n_142;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_60;
input n_152;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_125;
input n_35;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_29;
input n_79;
input n_131;
input n_151;
input n_47;
input n_25;
input n_53;
input n_8;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_109;
input n_112;
input n_85;
input n_95;
input n_119;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_27;
input n_64;
input n_77;
input n_102;
input n_106;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_134;
input n_32;
input n_41;
input n_104;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_11;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_1719;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1166;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1677;
wire n_1150;
wire n_226;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_155;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1021;
wire n_551;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1695;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_1666;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_1545;
wire n_864;
wire n_173;
wire n_859;
wire n_951;
wire n_1264;
wire n_447;
wire n_247;
wire n_1494;
wire n_292;
wire n_625;
wire n_854;
wire n_1462;
wire n_1580;
wire n_674;
wire n_417;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_1607;
wire n_1563;
wire n_606;
wire n_275;
wire n_877;
wire n_1696;
wire n_755;
wire n_1118;
wire n_1686;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1359;
wire n_530;
wire n_1107;
wire n_556;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_929;
wire n_1124;
wire n_902;
wire n_1576;
wire n_191;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1705;
wire n_1257;
wire n_171;
wire n_1182;
wire n_579;
wire n_1698;
wire n_1261;
wire n_938;
wire n_1098;
wire n_320;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_406;
wire n_519;
wire n_1016;
wire n_1243;
wire n_546;
wire n_1280;
wire n_281;
wire n_240;
wire n_291;
wire n_231;
wire n_257;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_317;
wire n_1236;
wire n_1633;
wire n_569;
wire n_227;
wire n_920;
wire n_1289;
wire n_1517;
wire n_335;
wire n_1669;
wire n_370;
wire n_976;
wire n_343;
wire n_1449;
wire n_308;
wire n_1566;
wire n_297;
wire n_156;
wire n_1078;
wire n_1670;
wire n_775;
wire n_219;
wire n_157;
wire n_600;
wire n_1484;
wire n_1374;
wire n_1328;
wire n_223;
wire n_264;
wire n_1598;
wire n_955;
wire n_163;
wire n_339;
wire n_1146;
wire n_882;
wire n_183;
wire n_243;
wire n_1036;
wire n_1097;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_215;
wire n_350;
wire n_196;
wire n_798;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_290;
wire n_580;
wire n_1040;
wire n_578;
wire n_926;
wire n_344;
wire n_1218;
wire n_422;
wire n_475;
wire n_777;
wire n_1070;
wire n_1547;
wire n_1030;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_663;
wire n_845;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_680;
wire n_1473;
wire n_1587;
wire n_395;
wire n_164;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_214;
wire n_1672;
wire n_675;
wire n_888;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1556;
wire n_1384;
wire n_184;
wire n_446;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_1706;
wire n_468;
wire n_213;
wire n_342;
wire n_464;
wire n_363;
wire n_1582;
wire n_197;
wire n_1069;
wire n_1075;
wire n_1450;
wire n_1322;
wire n_1471;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_1700;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1599;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_907;
wire n_1447;
wire n_1377;
wire n_190;
wire n_989;
wire n_1039;
wire n_228;
wire n_283;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_310;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_1667;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1248;
wire n_230;
wire n_1331;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_476;
wire n_1527;
wire n_534;
wire n_884;
wire n_345;
wire n_944;
wire n_1623;
wire n_1565;
wire n_182;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_832;
wire n_857;
wire n_207;
wire n_561;
wire n_1319;
wire n_1712;
wire n_1387;
wire n_1532;
wire n_1027;
wire n_971;
wire n_1156;
wire n_326;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_1709;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1538;
wire n_1199;
wire n_352;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_1660;
wire n_887;
wire n_154;
wire n_300;
wire n_809;
wire n_870;
wire n_931;
wire n_599;
wire n_1711;
wire n_1662;
wire n_1481;
wire n_434;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1629;
wire n_1293;
wire n_965;
wire n_935;
wire n_1175;
wire n_817;
wire n_360;
wire n_1479;
wire n_759;
wire n_806;
wire n_1477;
wire n_324;
wire n_1635;
wire n_1571;
wire n_187;
wire n_1189;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_784;
wire n_1244;
wire n_431;
wire n_1194;
wire n_615;
wire n_851;
wire n_843;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_1679;
wire n_776;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1647;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_1674;
wire n_1710;
wire n_284;
wire n_1128;
wire n_744;
wire n_590;
wire n_629;
wire n_1308;
wire n_254;
wire n_1680;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_526;
wire n_372;
wire n_293;
wire n_677;
wire n_244;
wire n_1333;
wire n_1121;
wire n_368;
wire n_314;
wire n_433;
wire n_604;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_498;
wire n_1468;
wire n_1559;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_252;
wire n_624;
wire n_1380;
wire n_1617;
wire n_295;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_610;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_448;
wire n_259;
wire n_758;
wire n_999;
wire n_1656;
wire n_1158;
wire n_1509;
wire n_563;
wire n_1145;
wire n_878;
wire n_524;
wire n_394;
wire n_204;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_331;
wire n_906;
wire n_1163;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_658;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_592;
wire n_1169;
wire n_1596;
wire n_1692;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_1095;
wire n_1614;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_1431;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1640;
wire n_1009;
wire n_1148;
wire n_742;
wire n_750;
wire n_995;
wire n_454;
wire n_1609;
wire n_374;
wire n_185;
wire n_396;
wire n_1383;
wire n_1073;
wire n_255;
wire n_662;
wire n_459;
wire n_218;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1574;
wire n_473;
wire n_1309;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_1548;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_168;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_208;
wire n_743;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_1240;
wire n_829;
wire n_1612;
wire n_1416;
wire n_361;
wire n_700;
wire n_1237;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1568;
wire n_1006;
wire n_329;
wire n_274;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_309;
wire n_512;
wire n_1591;
wire n_322;
wire n_1682;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1349;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_224;
wire n_1562;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_239;
wire n_630;
wire n_504;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_1304;
wire n_1324;
wire n_987;
wire n_261;
wire n_174;
wire n_1455;
wire n_767;
wire n_993;
wire n_1407;
wire n_1551;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_729;
wire n_1131;
wire n_1084;
wire n_970;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_340;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_1645;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_1684;
wire n_233;
wire n_1717;
wire n_572;
wire n_366;
wire n_815;
wire n_327;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_1708;
wire n_426;
wire n_1438;
wire n_1082;
wire n_589;
wire n_716;
wire n_1630;
wire n_562;
wire n_1436;
wire n_1691;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_531;
wire n_890;
wire n_764;
wire n_1056;
wire n_1424;
wire n_162;
wire n_960;
wire n_222;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_634;
wire n_199;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_1519;
wire n_256;
wire n_950;
wire n_1553;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1060;
wire n_1141;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_912;
wire n_315;
wire n_968;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_1699;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_1608;
wire n_983;
wire n_280;
wire n_1305;
wire n_873;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_1644;
wire n_690;
wire n_583;
wire n_302;
wire n_1343;
wire n_1203;
wire n_1631;
wire n_821;
wire n_321;
wire n_1179;
wire n_753;
wire n_621;
wire n_455;
wire n_1048;
wire n_1288;
wire n_385;
wire n_212;
wire n_507;
wire n_1560;
wire n_1605;
wire n_330;
wire n_1228;
wire n_972;
wire n_692;
wire n_820;
wire n_1200;
wire n_1301;
wire n_1363;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_1688;
wire n_945;
wire n_492;
wire n_1504;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_286;
wire n_1643;
wire n_883;
wire n_470;
wire n_449;
wire n_325;
wire n_1594;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_856;
wire n_918;
wire n_942;
wire n_189;
wire n_1147;
wire n_1557;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_195;
wire n_356;
wire n_894;
wire n_1636;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1470;
wire n_1096;
wire n_234;
wire n_1575;
wire n_1697;
wire n_833;
wire n_1646;
wire n_225;
wire n_1307;
wire n_988;
wire n_814;
wire n_192;
wire n_1549;
wire n_1201;
wire n_1114;
wire n_655;
wire n_1616;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_387;
wire n_1149;
wire n_398;
wire n_1671;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_211;
wire n_1219;
wire n_1204;
wire n_178;
wire n_1035;
wire n_287;
wire n_555;
wire n_783;
wire n_1188;
wire n_661;
wire n_849;
wire n_336;
wire n_584;
wire n_681;
wire n_1638;
wire n_430;
wire n_510;
wire n_216;
wire n_311;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_1655;
wire n_445;
wire n_749;
wire n_1134;
wire n_1358;
wire n_717;
wire n_165;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_249;
wire n_304;
wire n_1338;
wire n_577;
wire n_1522;
wire n_1687;
wire n_1637;
wire n_1419;
wire n_338;
wire n_1653;
wire n_693;
wire n_1506;
wire n_836;
wire n_990;
wire n_1389;
wire n_975;
wire n_1256;
wire n_1702;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_306;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1164;
wire n_1659;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_1572;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1685;
wire n_601;
wire n_917;
wire n_1714;
wire n_966;
wire n_253;
wire n_1116;
wire n_1661;
wire n_1212;
wire n_1541;
wire n_172;
wire n_206;
wire n_217;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_818;
wire n_861;
wire n_1713;
wire n_1183;
wire n_1658;
wire n_899;
wire n_1253;
wire n_210;
wire n_774;
wire n_1628;
wire n_1335;
wire n_1514;
wire n_1059;
wire n_1345;
wire n_176;
wire n_1133;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_1168;
wire n_707;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_1584;
wire n_665;
wire n_1440;
wire n_177;
wire n_421;
wire n_1356;
wire n_910;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_205;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_179;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_735;
wire n_232;
wire n_1109;
wire n_895;
wire n_1310;
wire n_202;
wire n_427;
wire n_1399;
wire n_1543;
wire n_791;
wire n_732;
wire n_1533;
wire n_193;
wire n_808;
wire n_797;
wire n_1025;
wire n_500;
wire n_1067;
wire n_435;
wire n_159;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_594;
wire n_200;
wire n_1291;
wire n_1297;
wire n_1155;
wire n_1418;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_985;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1703;
wire n_1352;
wire n_626;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_305;
wire n_676;
wire n_294;
wire n_318;
wire n_653;
wire n_642;
wire n_1602;
wire n_194;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_268;
wire n_664;
wire n_503;
wire n_235;
wire n_1372;
wire n_605;
wire n_1273;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_581;
wire n_382;
wire n_554;
wire n_1625;
wire n_898;
wire n_1013;
wire n_1452;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_198;
wire n_714;
wire n_1683;
wire n_909;
wire n_1497;
wire n_1530;
wire n_997;
wire n_932;
wire n_612;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_508;
wire n_506;
wire n_1320;
wire n_1663;
wire n_737;
wire n_1718;
wire n_986;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1715;
wire n_1281;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_209;
wire n_1564;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1376;
wire n_941;
wire n_981;
wire n_1569;
wire n_867;
wire n_186;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_518;
wire n_505;
wire n_282;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1620;
wire n_381;
wire n_220;
wire n_390;
wire n_1330;
wire n_481;
wire n_1675;
wire n_1554;
wire n_769;
wire n_1046;
wire n_271;
wire n_934;
wire n_1618;
wire n_826;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_167;
wire n_428;
wire n_379;
wire n_1341;
wire n_570;
wire n_1641;
wire n_1361;
wire n_1707;
wire n_853;
wire n_377;
wire n_751;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_158;
wire n_704;
wire n_787;
wire n_961;
wire n_771;
wire n_276;
wire n_1716;
wire n_1225;
wire n_1520;
wire n_169;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_181;
wire n_1411;
wire n_221;
wire n_622;
wire n_1577;
wire n_1087;
wire n_386;
wire n_994;
wire n_1701;
wire n_848;
wire n_1550;
wire n_1498;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1344;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_432;
wire n_839;
wire n_1210;
wire n_1364;
wire n_328;
wire n_1250;
wire n_369;
wire n_871;
wire n_598;
wire n_685;
wire n_608;
wire n_928;
wire n_1367;
wire n_1460;
wire n_772;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_413;
wire n_402;
wire n_1086;
wire n_796;
wire n_1619;
wire n_236;
wire n_1502;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_903;
wire n_1525;
wire n_740;
wire n_203;
wire n_384;
wire n_1404;
wire n_1315;
wire n_277;
wire n_1061;
wire n_333;
wire n_1298;
wire n_1652;
wire n_462;
wire n_1193;
wire n_1676;
wire n_1255;
wire n_258;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_188;
wire n_844;
wire n_201;
wire n_471;
wire n_852;
wire n_1487;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_1673;
wire n_465;
wire n_362;
wire n_1321;
wire n_170;
wire n_161;
wire n_273;
wire n_585;
wire n_270;
wire n_616;
wire n_745;
wire n_1654;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_641;
wire n_730;
wire n_1325;
wire n_1595;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_180;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_229;
wire n_437;
wire n_1642;
wire n_453;
wire n_403;
wire n_1130;
wire n_720;
wire n_1526;
wire n_863;
wire n_805;
wire n_1604;
wire n_1275;
wire n_712;
wire n_246;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_269;
wire n_285;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_1621;
wire n_251;
wire n_160;
wire n_566;
wire n_565;
wire n_1448;
wire n_1507;
wire n_1398;
wire n_597;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_651;
wire n_1340;
wire n_334;
wire n_811;
wire n_1558;
wire n_807;
wire n_835;
wire n_175;
wire n_666;
wire n_262;
wire n_1433;
wire n_1704;
wire n_1254;
wire n_1026;
wire n_1234;
wire n_319;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_242;
wire n_1681;
wire n_1018;
wire n_1693;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_166;
wire n_1180;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;
wire n_278;

INVxp67_ASAP7_75t_L g154 ( 
.A(n_54),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_26),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_101),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_94),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_63),
.Y(n_158)
);

CKINVDCx5p33_ASAP7_75t_R g159 ( 
.A(n_19),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_97),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_119),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_46),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_126),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_140),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_29),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_48),
.Y(n_166)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_88),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_50),
.Y(n_168)
);

BUFx3_ASAP7_75t_L g169 ( 
.A(n_38),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_91),
.Y(n_170)
);

BUFx3_ASAP7_75t_L g171 ( 
.A(n_83),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_61),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_107),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_92),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_41),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_5),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_105),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_96),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_124),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_120),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_85),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_111),
.Y(n_182)
);

INVx1_ASAP7_75t_SL g183 ( 
.A(n_19),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_69),
.Y(n_184)
);

BUFx5_ASAP7_75t_L g185 ( 
.A(n_13),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_136),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_40),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_55),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_44),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_135),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_108),
.Y(n_191)
);

INVx2_ASAP7_75t_SL g192 ( 
.A(n_51),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_104),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_128),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_43),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_109),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_137),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_36),
.Y(n_198)
);

BUFx6f_ASAP7_75t_L g199 ( 
.A(n_152),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_58),
.Y(n_200)
);

CKINVDCx16_ASAP7_75t_R g201 ( 
.A(n_103),
.Y(n_201)
);

INVxp67_ASAP7_75t_L g202 ( 
.A(n_147),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_13),
.Y(n_203)
);

INVx1_ASAP7_75t_SL g204 ( 
.A(n_144),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_6),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_20),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_134),
.Y(n_207)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_74),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_86),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_55),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_84),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_15),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_125),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_15),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_81),
.Y(n_215)
);

BUFx2_ASAP7_75t_L g216 ( 
.A(n_142),
.Y(n_216)
);

CKINVDCx16_ASAP7_75t_R g217 ( 
.A(n_110),
.Y(n_217)
);

INVx2_ASAP7_75t_SL g218 ( 
.A(n_20),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_146),
.Y(n_219)
);

BUFx8_ASAP7_75t_SL g220 ( 
.A(n_62),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_34),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_37),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_100),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_118),
.Y(n_224)
);

BUFx2_ASAP7_75t_L g225 ( 
.A(n_141),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_9),
.Y(n_226)
);

INVx1_ASAP7_75t_SL g227 ( 
.A(n_59),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_16),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_16),
.Y(n_229)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_30),
.Y(n_230)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_78),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_17),
.Y(n_232)
);

CKINVDCx16_ASAP7_75t_R g233 ( 
.A(n_95),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_145),
.Y(n_234)
);

BUFx10_ASAP7_75t_L g235 ( 
.A(n_149),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_57),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_90),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_153),
.Y(n_238)
);

INVx1_ASAP7_75t_SL g239 ( 
.A(n_130),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_18),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_127),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_50),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_76),
.Y(n_243)
);

BUFx3_ASAP7_75t_L g244 ( 
.A(n_10),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_36),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_51),
.Y(n_246)
);

HB1xp67_ASAP7_75t_L g247 ( 
.A(n_0),
.Y(n_247)
);

BUFx2_ASAP7_75t_L g248 ( 
.A(n_73),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_40),
.Y(n_249)
);

INVx1_ASAP7_75t_SL g250 ( 
.A(n_1),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_53),
.Y(n_251)
);

CKINVDCx16_ASAP7_75t_R g252 ( 
.A(n_114),
.Y(n_252)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_25),
.Y(n_253)
);

INVx1_ASAP7_75t_SL g254 ( 
.A(n_7),
.Y(n_254)
);

INVx2_ASAP7_75t_SL g255 ( 
.A(n_87),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_133),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_106),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_131),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_23),
.Y(n_259)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_1),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_68),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_132),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_47),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_22),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_29),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_22),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_139),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_12),
.Y(n_268)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_42),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_102),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_37),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_79),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_72),
.Y(n_273)
);

INVx1_ASAP7_75t_SL g274 ( 
.A(n_82),
.Y(n_274)
);

INVx2_ASAP7_75t_SL g275 ( 
.A(n_56),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_31),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_53),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_26),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_32),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_31),
.Y(n_280)
);

INVx1_ASAP7_75t_SL g281 ( 
.A(n_21),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_0),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_150),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_71),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_148),
.Y(n_285)
);

INVx2_ASAP7_75t_SL g286 ( 
.A(n_99),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_11),
.Y(n_287)
);

BUFx10_ASAP7_75t_L g288 ( 
.A(n_129),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_6),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_93),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_60),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_32),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_138),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_80),
.Y(n_294)
);

INVx1_ASAP7_75t_SL g295 ( 
.A(n_17),
.Y(n_295)
);

BUFx5_ASAP7_75t_L g296 ( 
.A(n_47),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_44),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_116),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_7),
.Y(n_299)
);

INVx1_ASAP7_75t_SL g300 ( 
.A(n_64),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_46),
.Y(n_301)
);

HB1xp67_ASAP7_75t_L g302 ( 
.A(n_48),
.Y(n_302)
);

BUFx6f_ASAP7_75t_L g303 ( 
.A(n_42),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_43),
.Y(n_304)
);

BUFx3_ASAP7_75t_L g305 ( 
.A(n_65),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_185),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_216),
.B(n_2),
.Y(n_307)
);

BUFx6f_ASAP7_75t_L g308 ( 
.A(n_199),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_185),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_185),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_157),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_220),
.Y(n_312)
);

INVxp33_ASAP7_75t_SL g313 ( 
.A(n_247),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_158),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_161),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_163),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_172),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_164),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_174),
.Y(n_319)
);

INVxp67_ASAP7_75t_SL g320 ( 
.A(n_216),
.Y(n_320)
);

INVxp67_ASAP7_75t_SL g321 ( 
.A(n_225),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_185),
.B(n_2),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_177),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_185),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_223),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_237),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_185),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_185),
.Y(n_328)
);

CKINVDCx14_ASAP7_75t_R g329 ( 
.A(n_225),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_185),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_185),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_296),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_296),
.Y(n_333)
);

INVxp67_ASAP7_75t_L g334 ( 
.A(n_302),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_296),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_296),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_262),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_296),
.Y(n_338)
);

INVxp67_ASAP7_75t_L g339 ( 
.A(n_168),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_296),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_296),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_178),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_182),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_296),
.Y(n_344)
);

CKINVDCx16_ASAP7_75t_R g345 ( 
.A(n_201),
.Y(n_345)
);

CKINVDCx20_ASAP7_75t_R g346 ( 
.A(n_267),
.Y(n_346)
);

HB1xp67_ASAP7_75t_L g347 ( 
.A(n_159),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_184),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_296),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_186),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_303),
.Y(n_351)
);

INVxp33_ASAP7_75t_SL g352 ( 
.A(n_165),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_303),
.Y(n_353)
);

INVxp67_ASAP7_75t_SL g354 ( 
.A(n_248),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_190),
.Y(n_355)
);

INVx1_ASAP7_75t_SL g356 ( 
.A(n_155),
.Y(n_356)
);

AND2x2_ASAP7_75t_L g357 ( 
.A(n_244),
.B(n_3),
.Y(n_357)
);

CKINVDCx20_ASAP7_75t_R g358 ( 
.A(n_291),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_303),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g360 ( 
.A(n_201),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_303),
.Y(n_361)
);

BUFx3_ASAP7_75t_L g362 ( 
.A(n_171),
.Y(n_362)
);

INVxp67_ASAP7_75t_SL g363 ( 
.A(n_248),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g364 ( 
.A(n_217),
.Y(n_364)
);

NOR2xp67_ASAP7_75t_L g365 ( 
.A(n_154),
.B(n_3),
.Y(n_365)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_217),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_303),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_230),
.Y(n_368)
);

CKINVDCx20_ASAP7_75t_R g369 ( 
.A(n_233),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_191),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_193),
.Y(n_371)
);

INVxp67_ASAP7_75t_SL g372 ( 
.A(n_171),
.Y(n_372)
);

BUFx6f_ASAP7_75t_SL g373 ( 
.A(n_235),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_230),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_253),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_253),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_260),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_260),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_269),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_269),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_372),
.B(n_255),
.Y(n_381)
);

BUFx6f_ASAP7_75t_L g382 ( 
.A(n_308),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_351),
.Y(n_383)
);

AND2x2_ASAP7_75t_L g384 ( 
.A(n_357),
.B(n_362),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_351),
.Y(n_385)
);

BUFx6f_ASAP7_75t_L g386 ( 
.A(n_308),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_353),
.Y(n_387)
);

OA21x2_ASAP7_75t_L g388 ( 
.A1(n_322),
.A2(n_187),
.B(n_168),
.Y(n_388)
);

BUFx6f_ASAP7_75t_L g389 ( 
.A(n_308),
.Y(n_389)
);

BUFx6f_ASAP7_75t_L g390 ( 
.A(n_308),
.Y(n_390)
);

INVx3_ASAP7_75t_L g391 ( 
.A(n_308),
.Y(n_391)
);

BUFx3_ASAP7_75t_L g392 ( 
.A(n_353),
.Y(n_392)
);

AND2x2_ASAP7_75t_L g393 ( 
.A(n_357),
.B(n_362),
.Y(n_393)
);

AND2x6_ASAP7_75t_L g394 ( 
.A(n_306),
.B(n_167),
.Y(n_394)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_333),
.Y(n_395)
);

BUFx6f_ASAP7_75t_L g396 ( 
.A(n_306),
.Y(n_396)
);

INVx2_ASAP7_75t_L g397 ( 
.A(n_335),
.Y(n_397)
);

AND2x6_ASAP7_75t_L g398 ( 
.A(n_309),
.B(n_167),
.Y(n_398)
);

INVxp67_ASAP7_75t_L g399 ( 
.A(n_347),
.Y(n_399)
);

NOR2x1_ASAP7_75t_L g400 ( 
.A(n_359),
.B(n_305),
.Y(n_400)
);

AND2x2_ASAP7_75t_L g401 ( 
.A(n_359),
.B(n_361),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_361),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_367),
.B(n_255),
.Y(n_403)
);

INVx2_ASAP7_75t_L g404 ( 
.A(n_309),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_367),
.B(n_286),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_310),
.Y(n_406)
);

AND2x4_ASAP7_75t_L g407 ( 
.A(n_310),
.B(n_305),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_324),
.B(n_286),
.Y(n_408)
);

INVx3_ASAP7_75t_L g409 ( 
.A(n_324),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_327),
.B(n_196),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_327),
.Y(n_411)
);

INVx3_ASAP7_75t_L g412 ( 
.A(n_328),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_328),
.Y(n_413)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_330),
.Y(n_414)
);

CKINVDCx9p33_ASAP7_75t_R g415 ( 
.A(n_307),
.Y(n_415)
);

INVx3_ASAP7_75t_L g416 ( 
.A(n_330),
.Y(n_416)
);

AND2x4_ASAP7_75t_L g417 ( 
.A(n_331),
.B(n_305),
.Y(n_417)
);

AND2x4_ASAP7_75t_L g418 ( 
.A(n_331),
.B(n_208),
.Y(n_418)
);

AND2x4_ASAP7_75t_L g419 ( 
.A(n_332),
.B(n_208),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_332),
.Y(n_420)
);

INVx3_ASAP7_75t_L g421 ( 
.A(n_336),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_336),
.Y(n_422)
);

INVx3_ASAP7_75t_L g423 ( 
.A(n_338),
.Y(n_423)
);

AND2x4_ASAP7_75t_L g424 ( 
.A(n_338),
.B(n_231),
.Y(n_424)
);

AND2x4_ASAP7_75t_L g425 ( 
.A(n_340),
.B(n_231),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_340),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_341),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_341),
.Y(n_428)
);

BUFx2_ASAP7_75t_L g429 ( 
.A(n_360),
.Y(n_429)
);

INVx2_ASAP7_75t_L g430 ( 
.A(n_344),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_344),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_349),
.B(n_197),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_349),
.Y(n_433)
);

OR2x2_ASAP7_75t_L g434 ( 
.A(n_320),
.B(n_192),
.Y(n_434)
);

NOR2xp33_ASAP7_75t_SL g435 ( 
.A(n_345),
.B(n_233),
.Y(n_435)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_368),
.Y(n_436)
);

AND2x4_ASAP7_75t_L g437 ( 
.A(n_368),
.B(n_156),
.Y(n_437)
);

BUFx6f_ASAP7_75t_L g438 ( 
.A(n_374),
.Y(n_438)
);

INVx2_ASAP7_75t_L g439 ( 
.A(n_374),
.Y(n_439)
);

BUFx2_ASAP7_75t_L g440 ( 
.A(n_364),
.Y(n_440)
);

INVx3_ASAP7_75t_L g441 ( 
.A(n_380),
.Y(n_441)
);

OA21x2_ASAP7_75t_L g442 ( 
.A1(n_375),
.A2(n_221),
.B(n_187),
.Y(n_442)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_375),
.Y(n_443)
);

BUFx6f_ASAP7_75t_L g444 ( 
.A(n_376),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_321),
.B(n_200),
.Y(n_445)
);

AND2x2_ASAP7_75t_L g446 ( 
.A(n_354),
.B(n_244),
.Y(n_446)
);

INVx2_ASAP7_75t_L g447 ( 
.A(n_376),
.Y(n_447)
);

AND2x4_ASAP7_75t_L g448 ( 
.A(n_377),
.B(n_156),
.Y(n_448)
);

INVxp67_ASAP7_75t_L g449 ( 
.A(n_363),
.Y(n_449)
);

INVx3_ASAP7_75t_L g450 ( 
.A(n_382),
.Y(n_450)
);

INVxp67_ASAP7_75t_SL g451 ( 
.A(n_409),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_401),
.Y(n_452)
);

NAND3xp33_ASAP7_75t_L g453 ( 
.A(n_449),
.B(n_329),
.C(n_334),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_SL g454 ( 
.A(n_435),
.B(n_314),
.Y(n_454)
);

INVx3_ASAP7_75t_L g455 ( 
.A(n_382),
.Y(n_455)
);

INVx4_ASAP7_75t_L g456 ( 
.A(n_396),
.Y(n_456)
);

INVx2_ASAP7_75t_L g457 ( 
.A(n_404),
.Y(n_457)
);

HB1xp67_ASAP7_75t_L g458 ( 
.A(n_384),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_401),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_401),
.Y(n_460)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_404),
.Y(n_461)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_404),
.Y(n_462)
);

INVx2_ASAP7_75t_L g463 ( 
.A(n_404),
.Y(n_463)
);

INVx2_ASAP7_75t_L g464 ( 
.A(n_414),
.Y(n_464)
);

AND2x2_ASAP7_75t_SL g465 ( 
.A(n_435),
.B(n_252),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_406),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_406),
.Y(n_467)
);

CKINVDCx5p33_ASAP7_75t_R g468 ( 
.A(n_429),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_SL g469 ( 
.A(n_449),
.B(n_315),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_406),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_411),
.Y(n_471)
);

BUFx6f_ASAP7_75t_L g472 ( 
.A(n_382),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_411),
.Y(n_473)
);

BUFx3_ASAP7_75t_L g474 ( 
.A(n_388),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_411),
.Y(n_475)
);

INVx2_ASAP7_75t_L g476 ( 
.A(n_414),
.Y(n_476)
);

AOI22xp33_ASAP7_75t_L g477 ( 
.A1(n_388),
.A2(n_313),
.B1(n_275),
.B2(n_192),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_413),
.Y(n_478)
);

INVx5_ASAP7_75t_L g479 ( 
.A(n_394),
.Y(n_479)
);

INVxp67_ASAP7_75t_L g480 ( 
.A(n_445),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_410),
.B(n_316),
.Y(n_481)
);

INVx2_ASAP7_75t_L g482 ( 
.A(n_414),
.Y(n_482)
);

BUFx3_ASAP7_75t_L g483 ( 
.A(n_388),
.Y(n_483)
);

INVx4_ASAP7_75t_SL g484 ( 
.A(n_394),
.Y(n_484)
);

INVx3_ASAP7_75t_L g485 ( 
.A(n_382),
.Y(n_485)
);

BUFx4f_ASAP7_75t_L g486 ( 
.A(n_388),
.Y(n_486)
);

INVx2_ASAP7_75t_L g487 ( 
.A(n_414),
.Y(n_487)
);

BUFx10_ASAP7_75t_L g488 ( 
.A(n_407),
.Y(n_488)
);

INVxp33_ASAP7_75t_L g489 ( 
.A(n_446),
.Y(n_489)
);

AO22x2_ASAP7_75t_L g490 ( 
.A1(n_434),
.A2(n_218),
.B1(n_275),
.B2(n_246),
.Y(n_490)
);

NOR2xp33_ASAP7_75t_L g491 ( 
.A(n_445),
.B(n_352),
.Y(n_491)
);

AOI22xp33_ASAP7_75t_L g492 ( 
.A1(n_388),
.A2(n_218),
.B1(n_244),
.B2(n_169),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_410),
.B(n_318),
.Y(n_493)
);

NOR2x1p5_ASAP7_75t_L g494 ( 
.A(n_434),
.B(n_312),
.Y(n_494)
);

INVx8_ASAP7_75t_L g495 ( 
.A(n_384),
.Y(n_495)
);

INVx2_ASAP7_75t_L g496 ( 
.A(n_430),
.Y(n_496)
);

AND3x1_ASAP7_75t_L g497 ( 
.A(n_446),
.B(n_246),
.C(n_221),
.Y(n_497)
);

BUFx2_ASAP7_75t_L g498 ( 
.A(n_399),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_413),
.Y(n_499)
);

AOI22xp33_ASAP7_75t_L g500 ( 
.A1(n_388),
.A2(n_169),
.B1(n_287),
.B2(n_266),
.Y(n_500)
);

INVx2_ASAP7_75t_SL g501 ( 
.A(n_384),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_432),
.B(n_319),
.Y(n_502)
);

OR2x2_ASAP7_75t_L g503 ( 
.A(n_434),
.B(n_356),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_413),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_420),
.Y(n_505)
);

NAND2xp33_ASAP7_75t_L g506 ( 
.A(n_394),
.B(n_199),
.Y(n_506)
);

OR2x6_ASAP7_75t_L g507 ( 
.A(n_446),
.B(n_365),
.Y(n_507)
);

INVx2_ASAP7_75t_SL g508 ( 
.A(n_393),
.Y(n_508)
);

AOI22xp33_ASAP7_75t_L g509 ( 
.A1(n_407),
.A2(n_277),
.B1(n_266),
.B2(n_268),
.Y(n_509)
);

AND3x1_ASAP7_75t_L g510 ( 
.A(n_415),
.B(n_271),
.C(n_268),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_SL g511 ( 
.A(n_399),
.B(n_323),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_420),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_420),
.Y(n_513)
);

NOR2xp33_ASAP7_75t_L g514 ( 
.A(n_393),
.B(n_342),
.Y(n_514)
);

INVx3_ASAP7_75t_L g515 ( 
.A(n_382),
.Y(n_515)
);

NOR2xp33_ASAP7_75t_L g516 ( 
.A(n_393),
.B(n_343),
.Y(n_516)
);

NOR2xp33_ASAP7_75t_L g517 ( 
.A(n_381),
.B(n_348),
.Y(n_517)
);

AOI22xp33_ASAP7_75t_L g518 ( 
.A1(n_407),
.A2(n_271),
.B1(n_277),
.B2(n_282),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_422),
.Y(n_519)
);

NAND2xp33_ASAP7_75t_L g520 ( 
.A(n_394),
.B(n_199),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_SL g521 ( 
.A(n_381),
.B(n_350),
.Y(n_521)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_430),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_422),
.Y(n_523)
);

AND2x4_ASAP7_75t_L g524 ( 
.A(n_407),
.B(n_160),
.Y(n_524)
);

NOR2xp33_ASAP7_75t_L g525 ( 
.A(n_432),
.B(n_355),
.Y(n_525)
);

INVx4_ASAP7_75t_L g526 ( 
.A(n_396),
.Y(n_526)
);

NOR2xp33_ASAP7_75t_L g527 ( 
.A(n_422),
.B(n_370),
.Y(n_527)
);

INVxp67_ASAP7_75t_SL g528 ( 
.A(n_409),
.Y(n_528)
);

INVx2_ASAP7_75t_L g529 ( 
.A(n_395),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_426),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_426),
.Y(n_531)
);

NOR2xp33_ASAP7_75t_SL g532 ( 
.A(n_429),
.B(n_252),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_426),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_427),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_407),
.B(n_417),
.Y(n_535)
);

NOR2xp33_ASAP7_75t_L g536 ( 
.A(n_427),
.B(n_371),
.Y(n_536)
);

BUFx6f_ASAP7_75t_L g537 ( 
.A(n_382),
.Y(n_537)
);

INVx2_ASAP7_75t_L g538 ( 
.A(n_395),
.Y(n_538)
);

INVx3_ASAP7_75t_L g539 ( 
.A(n_382),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_407),
.B(n_204),
.Y(n_540)
);

AND2x2_ASAP7_75t_L g541 ( 
.A(n_417),
.B(n_380),
.Y(n_541)
);

AOI22xp33_ASAP7_75t_L g542 ( 
.A1(n_417),
.A2(n_287),
.B1(n_282),
.B2(n_373),
.Y(n_542)
);

BUFx6f_ASAP7_75t_L g543 ( 
.A(n_382),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_427),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_428),
.Y(n_545)
);

INVx5_ASAP7_75t_L g546 ( 
.A(n_394),
.Y(n_546)
);

INVx5_ASAP7_75t_L g547 ( 
.A(n_394),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_428),
.Y(n_548)
);

OR2x2_ASAP7_75t_L g549 ( 
.A(n_417),
.B(n_339),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_SL g550 ( 
.A(n_417),
.B(n_366),
.Y(n_550)
);

NOR3xp33_ASAP7_75t_L g551 ( 
.A(n_429),
.B(n_250),
.C(n_183),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_428),
.Y(n_552)
);

AOI22xp5_ASAP7_75t_L g553 ( 
.A1(n_417),
.A2(n_369),
.B1(n_373),
.B2(n_325),
.Y(n_553)
);

INVx4_ASAP7_75t_L g554 ( 
.A(n_396),
.Y(n_554)
);

INVx2_ASAP7_75t_L g555 ( 
.A(n_395),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_431),
.Y(n_556)
);

INVxp67_ASAP7_75t_L g557 ( 
.A(n_440),
.Y(n_557)
);

INVx4_ASAP7_75t_L g558 ( 
.A(n_396),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_SL g559 ( 
.A(n_437),
.B(n_235),
.Y(n_559)
);

INVxp33_ASAP7_75t_SL g560 ( 
.A(n_440),
.Y(n_560)
);

INVx2_ASAP7_75t_L g561 ( 
.A(n_395),
.Y(n_561)
);

INVxp33_ASAP7_75t_SL g562 ( 
.A(n_440),
.Y(n_562)
);

AND2x2_ASAP7_75t_L g563 ( 
.A(n_437),
.B(n_377),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_431),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_431),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_L g566 ( 
.A(n_433),
.B(n_227),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_SL g567 ( 
.A(n_448),
.B(n_235),
.Y(n_567)
);

BUFx3_ASAP7_75t_L g568 ( 
.A(n_442),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_397),
.Y(n_569)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_397),
.Y(n_570)
);

INVx2_ASAP7_75t_L g571 ( 
.A(n_397),
.Y(n_571)
);

AOI22xp33_ASAP7_75t_L g572 ( 
.A1(n_418),
.A2(n_373),
.B1(n_170),
.B2(n_160),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_397),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_433),
.Y(n_574)
);

AND2x2_ASAP7_75t_L g575 ( 
.A(n_437),
.B(n_378),
.Y(n_575)
);

CKINVDCx14_ASAP7_75t_R g576 ( 
.A(n_437),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_L g577 ( 
.A(n_433),
.B(n_239),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_442),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_442),
.Y(n_579)
);

BUFx6f_ASAP7_75t_L g580 ( 
.A(n_382),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_442),
.Y(n_581)
);

INVx2_ASAP7_75t_L g582 ( 
.A(n_383),
.Y(n_582)
);

AOI22xp33_ASAP7_75t_L g583 ( 
.A1(n_418),
.A2(n_257),
.B1(n_241),
.B2(n_272),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_L g584 ( 
.A(n_409),
.B(n_412),
.Y(n_584)
);

OR2x2_ASAP7_75t_L g585 ( 
.A(n_408),
.B(n_254),
.Y(n_585)
);

INVx2_ASAP7_75t_L g586 ( 
.A(n_383),
.Y(n_586)
);

OR2x6_ASAP7_75t_L g587 ( 
.A(n_442),
.B(n_170),
.Y(n_587)
);

INVx2_ASAP7_75t_L g588 ( 
.A(n_383),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_L g589 ( 
.A(n_409),
.B(n_274),
.Y(n_589)
);

NOR2xp33_ASAP7_75t_L g590 ( 
.A(n_408),
.B(n_311),
.Y(n_590)
);

BUFx4f_ASAP7_75t_L g591 ( 
.A(n_442),
.Y(n_591)
);

BUFx4f_ASAP7_75t_L g592 ( 
.A(n_396),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_409),
.Y(n_593)
);

INVx2_ASAP7_75t_L g594 ( 
.A(n_385),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_412),
.Y(n_595)
);

NOR2xp33_ASAP7_75t_L g596 ( 
.A(n_412),
.B(n_317),
.Y(n_596)
);

AOI22xp33_ASAP7_75t_L g597 ( 
.A1(n_568),
.A2(n_425),
.B1(n_424),
.B2(n_419),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_L g598 ( 
.A(n_525),
.B(n_412),
.Y(n_598)
);

NOR2xp33_ASAP7_75t_L g599 ( 
.A(n_480),
.B(n_281),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_L g600 ( 
.A(n_517),
.B(n_412),
.Y(n_600)
);

NOR2xp33_ASAP7_75t_L g601 ( 
.A(n_489),
.B(n_491),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_541),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_L g603 ( 
.A(n_481),
.B(n_416),
.Y(n_603)
);

AND2x2_ASAP7_75t_L g604 ( 
.A(n_498),
.B(n_503),
.Y(n_604)
);

AOI22xp33_ASAP7_75t_L g605 ( 
.A1(n_568),
.A2(n_425),
.B1(n_424),
.B2(n_418),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g606 ( 
.A(n_493),
.B(n_416),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_541),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_SL g608 ( 
.A(n_590),
.B(n_585),
.Y(n_608)
);

BUFx2_ASAP7_75t_L g609 ( 
.A(n_468),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_SL g610 ( 
.A(n_585),
.B(n_300),
.Y(n_610)
);

INVx2_ASAP7_75t_L g611 ( 
.A(n_582),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_L g612 ( 
.A(n_502),
.B(n_416),
.Y(n_612)
);

INVx2_ASAP7_75t_L g613 ( 
.A(n_582),
.Y(n_613)
);

INVx2_ASAP7_75t_L g614 ( 
.A(n_586),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_SL g615 ( 
.A(n_465),
.B(n_527),
.Y(n_615)
);

INVx2_ASAP7_75t_L g616 ( 
.A(n_586),
.Y(n_616)
);

OA22x2_ASAP7_75t_L g617 ( 
.A1(n_507),
.A2(n_415),
.B1(n_295),
.B2(n_448),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_458),
.Y(n_618)
);

NOR2xp33_ASAP7_75t_L g619 ( 
.A(n_521),
.B(n_416),
.Y(n_619)
);

OAI221xp5_ASAP7_75t_L g620 ( 
.A1(n_477),
.A2(n_518),
.B1(n_509),
.B2(n_583),
.C(n_492),
.Y(n_620)
);

BUFx2_ASAP7_75t_L g621 ( 
.A(n_468),
.Y(n_621)
);

NOR2xp33_ASAP7_75t_L g622 ( 
.A(n_536),
.B(n_416),
.Y(n_622)
);

NOR2x1p5_ASAP7_75t_L g623 ( 
.A(n_503),
.B(n_166),
.Y(n_623)
);

NOR3xp33_ASAP7_75t_L g624 ( 
.A(n_550),
.B(n_202),
.C(n_176),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_501),
.B(n_421),
.Y(n_625)
);

INVx2_ASAP7_75t_L g626 ( 
.A(n_588),
.Y(n_626)
);

INVx3_ASAP7_75t_L g627 ( 
.A(n_495),
.Y(n_627)
);

INVx2_ASAP7_75t_L g628 ( 
.A(n_588),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_501),
.B(n_421),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_L g630 ( 
.A(n_508),
.B(n_421),
.Y(n_630)
);

AND2x2_ASAP7_75t_L g631 ( 
.A(n_508),
.B(n_326),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_SL g632 ( 
.A(n_591),
.B(n_418),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_SL g633 ( 
.A(n_591),
.B(n_486),
.Y(n_633)
);

OAI221xp5_ASAP7_75t_L g634 ( 
.A1(n_500),
.A2(n_257),
.B1(n_181),
.B2(n_180),
.C(n_179),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_L g635 ( 
.A(n_452),
.B(n_421),
.Y(n_635)
);

NOR2xp33_ASAP7_75t_L g636 ( 
.A(n_469),
.B(n_421),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_L g637 ( 
.A(n_452),
.B(n_421),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_459),
.Y(n_638)
);

INVx3_ASAP7_75t_L g639 ( 
.A(n_495),
.Y(n_639)
);

BUFx6f_ASAP7_75t_L g640 ( 
.A(n_488),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_L g641 ( 
.A(n_459),
.B(n_423),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_SL g642 ( 
.A(n_591),
.B(n_418),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_L g643 ( 
.A(n_460),
.B(n_423),
.Y(n_643)
);

INVxp67_ASAP7_75t_L g644 ( 
.A(n_532),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_460),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_L g646 ( 
.A(n_451),
.B(n_423),
.Y(n_646)
);

INVxp67_ASAP7_75t_L g647 ( 
.A(n_453),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_563),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_528),
.B(n_423),
.Y(n_649)
);

OAI22xp5_ASAP7_75t_L g650 ( 
.A1(n_486),
.A2(n_337),
.B1(n_346),
.B2(n_358),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_SL g651 ( 
.A(n_465),
.B(n_207),
.Y(n_651)
);

AOI22xp33_ASAP7_75t_L g652 ( 
.A1(n_474),
.A2(n_419),
.B1(n_424),
.B2(n_425),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_L g653 ( 
.A(n_589),
.B(n_423),
.Y(n_653)
);

INVx2_ASAP7_75t_SL g654 ( 
.A(n_507),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_563),
.Y(n_655)
);

INVx4_ASAP7_75t_L g656 ( 
.A(n_495),
.Y(n_656)
);

INVx2_ASAP7_75t_SL g657 ( 
.A(n_507),
.Y(n_657)
);

NOR2xp33_ASAP7_75t_L g658 ( 
.A(n_514),
.B(n_423),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_575),
.Y(n_659)
);

INVx2_ASAP7_75t_L g660 ( 
.A(n_594),
.Y(n_660)
);

INVxp67_ASAP7_75t_SL g661 ( 
.A(n_578),
.Y(n_661)
);

NOR2xp33_ASAP7_75t_L g662 ( 
.A(n_516),
.B(n_175),
.Y(n_662)
);

OR2x6_ASAP7_75t_L g663 ( 
.A(n_557),
.B(n_437),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_540),
.B(n_418),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_SL g665 ( 
.A(n_486),
.B(n_419),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_575),
.Y(n_666)
);

INVx2_ASAP7_75t_SL g667 ( 
.A(n_507),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_535),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_466),
.Y(n_669)
);

OAI22xp5_ASAP7_75t_L g670 ( 
.A1(n_576),
.A2(n_549),
.B1(n_474),
.B2(n_483),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_466),
.B(n_419),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_467),
.B(n_419),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_SL g673 ( 
.A(n_483),
.B(n_419),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_SL g674 ( 
.A(n_488),
.B(n_424),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_467),
.B(n_424),
.Y(n_675)
);

NOR2xp33_ASAP7_75t_L g676 ( 
.A(n_549),
.B(n_511),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_SL g677 ( 
.A(n_488),
.B(n_424),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_SL g678 ( 
.A(n_578),
.B(n_425),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_SL g679 ( 
.A(n_579),
.B(n_425),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_470),
.B(n_471),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_SL g681 ( 
.A(n_579),
.B(n_425),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_SL g682 ( 
.A(n_581),
.B(n_396),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_SL g683 ( 
.A(n_581),
.B(n_396),
.Y(n_683)
);

BUFx8_ASAP7_75t_SL g684 ( 
.A(n_560),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_L g685 ( 
.A(n_470),
.B(n_396),
.Y(n_685)
);

BUFx6f_ASAP7_75t_L g686 ( 
.A(n_495),
.Y(n_686)
);

OAI22xp5_ASAP7_75t_L g687 ( 
.A1(n_542),
.A2(n_173),
.B1(n_179),
.B2(n_180),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_SL g688 ( 
.A(n_524),
.B(n_396),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_471),
.Y(n_689)
);

OAI22xp5_ASAP7_75t_L g690 ( 
.A1(n_596),
.A2(n_173),
.B1(n_181),
.B2(n_194),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_L g691 ( 
.A(n_473),
.B(n_475),
.Y(n_691)
);

INVx2_ASAP7_75t_L g692 ( 
.A(n_594),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_L g693 ( 
.A(n_473),
.B(n_392),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_L g694 ( 
.A(n_475),
.B(n_392),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_SL g695 ( 
.A(n_566),
.B(n_209),
.Y(n_695)
);

INVx2_ASAP7_75t_L g696 ( 
.A(n_478),
.Y(n_696)
);

INVxp33_ASAP7_75t_L g697 ( 
.A(n_551),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_SL g698 ( 
.A(n_524),
.B(n_199),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_478),
.B(n_392),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_L g700 ( 
.A(n_499),
.B(n_392),
.Y(n_700)
);

O2A1O1Ixp33_ASAP7_75t_L g701 ( 
.A1(n_587),
.A2(n_403),
.B(n_405),
.C(n_448),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_504),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_504),
.Y(n_703)
);

INVx2_ASAP7_75t_L g704 ( 
.A(n_505),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_L g705 ( 
.A(n_505),
.B(n_437),
.Y(n_705)
);

NOR2xp33_ASAP7_75t_L g706 ( 
.A(n_577),
.B(n_188),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_512),
.B(n_448),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_L g708 ( 
.A(n_512),
.B(n_513),
.Y(n_708)
);

A2O1A1Ixp33_ASAP7_75t_L g709 ( 
.A1(n_524),
.A2(n_448),
.B(n_284),
.C(n_194),
.Y(n_709)
);

INVx2_ASAP7_75t_L g710 ( 
.A(n_513),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_519),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_523),
.Y(n_712)
);

NAND2xp33_ASAP7_75t_L g713 ( 
.A(n_593),
.B(n_211),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_L g714 ( 
.A(n_523),
.B(n_448),
.Y(n_714)
);

INVx2_ASAP7_75t_L g715 ( 
.A(n_530),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_SL g716 ( 
.A(n_572),
.B(n_213),
.Y(n_716)
);

NOR2xp33_ASAP7_75t_L g717 ( 
.A(n_454),
.B(n_530),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_L g718 ( 
.A(n_531),
.B(n_441),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_L g719 ( 
.A(n_531),
.B(n_441),
.Y(n_719)
);

AOI22xp5_ASAP7_75t_L g720 ( 
.A1(n_559),
.A2(n_243),
.B1(n_273),
.B2(n_219),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_533),
.B(n_441),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_SL g722 ( 
.A(n_533),
.B(n_199),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_534),
.Y(n_723)
);

AO22x2_ASAP7_75t_L g724 ( 
.A1(n_567),
.A2(n_215),
.B1(n_241),
.B2(n_272),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_L g725 ( 
.A(n_534),
.B(n_441),
.Y(n_725)
);

BUFx8_ASAP7_75t_L g726 ( 
.A(n_560),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_L g727 ( 
.A(n_544),
.B(n_441),
.Y(n_727)
);

NOR2xp33_ASAP7_75t_L g728 ( 
.A(n_544),
.B(n_189),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_545),
.Y(n_729)
);

INVx2_ASAP7_75t_L g730 ( 
.A(n_545),
.Y(n_730)
);

INVx2_ASAP7_75t_L g731 ( 
.A(n_548),
.Y(n_731)
);

HB1xp67_ASAP7_75t_L g732 ( 
.A(n_497),
.Y(n_732)
);

OR2x2_ASAP7_75t_L g733 ( 
.A(n_553),
.B(n_195),
.Y(n_733)
);

BUFx6f_ASAP7_75t_L g734 ( 
.A(n_472),
.Y(n_734)
);

AND2x2_ASAP7_75t_L g735 ( 
.A(n_494),
.B(n_400),
.Y(n_735)
);

NOR2xp33_ASAP7_75t_L g736 ( 
.A(n_548),
.B(n_552),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_SL g737 ( 
.A(n_552),
.B(n_224),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_556),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_556),
.B(n_394),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_564),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_564),
.Y(n_741)
);

AOI22xp5_ASAP7_75t_L g742 ( 
.A1(n_510),
.A2(n_293),
.B1(n_283),
.B2(n_234),
.Y(n_742)
);

OR2x6_ASAP7_75t_L g743 ( 
.A(n_494),
.B(n_215),
.Y(n_743)
);

AOI22xp5_ASAP7_75t_L g744 ( 
.A1(n_587),
.A2(n_294),
.B1(n_236),
.B2(n_238),
.Y(n_744)
);

INVxp67_ASAP7_75t_L g745 ( 
.A(n_490),
.Y(n_745)
);

OAI22xp5_ASAP7_75t_SL g746 ( 
.A1(n_562),
.A2(n_265),
.B1(n_162),
.B2(n_276),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_565),
.B(n_394),
.Y(n_747)
);

NAND2xp33_ASAP7_75t_L g748 ( 
.A(n_593),
.B(n_256),
.Y(n_748)
);

INVx2_ASAP7_75t_L g749 ( 
.A(n_574),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_L g750 ( 
.A(n_574),
.B(n_394),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_L g751 ( 
.A(n_595),
.B(n_398),
.Y(n_751)
);

OR2x6_ASAP7_75t_L g752 ( 
.A(n_490),
.B(n_285),
.Y(n_752)
);

BUFx3_ASAP7_75t_L g753 ( 
.A(n_587),
.Y(n_753)
);

AOI221xp5_ASAP7_75t_L g754 ( 
.A1(n_490),
.A2(n_214),
.B1(n_198),
.B2(n_203),
.C(n_205),
.Y(n_754)
);

AOI22xp5_ASAP7_75t_L g755 ( 
.A1(n_490),
.A2(n_584),
.B1(n_261),
.B2(n_270),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_L g756 ( 
.A(n_450),
.B(n_398),
.Y(n_756)
);

NOR2xp33_ASAP7_75t_L g757 ( 
.A(n_456),
.B(n_206),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_L g758 ( 
.A(n_450),
.B(n_455),
.Y(n_758)
);

BUFx6f_ASAP7_75t_L g759 ( 
.A(n_472),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_SL g760 ( 
.A(n_562),
.B(n_258),
.Y(n_760)
);

AND2x2_ASAP7_75t_L g761 ( 
.A(n_529),
.B(n_400),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_529),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_661),
.B(n_457),
.Y(n_763)
);

A2O1A1Ixp33_ASAP7_75t_L g764 ( 
.A1(n_717),
.A2(n_285),
.B(n_290),
.C(n_298),
.Y(n_764)
);

AND2x2_ASAP7_75t_L g765 ( 
.A(n_604),
.B(n_378),
.Y(n_765)
);

AOI21xp5_ASAP7_75t_L g766 ( 
.A1(n_632),
.A2(n_592),
.B(n_558),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_SL g767 ( 
.A(n_601),
.B(n_676),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_L g768 ( 
.A(n_668),
.B(n_457),
.Y(n_768)
);

NOR2x1_ASAP7_75t_L g769 ( 
.A(n_608),
.B(n_403),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_L g770 ( 
.A(n_622),
.B(n_461),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_622),
.B(n_461),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_SL g772 ( 
.A(n_601),
.B(n_676),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_658),
.B(n_462),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_L g774 ( 
.A(n_658),
.B(n_462),
.Y(n_774)
);

AOI21xp5_ASAP7_75t_L g775 ( 
.A1(n_632),
.A2(n_592),
.B(n_558),
.Y(n_775)
);

OAI22xp5_ASAP7_75t_L g776 ( 
.A1(n_753),
.A2(n_592),
.B1(n_290),
.B2(n_298),
.Y(n_776)
);

AOI21xp5_ASAP7_75t_L g777 ( 
.A1(n_642),
.A2(n_665),
.B(n_674),
.Y(n_777)
);

AOI21xp5_ASAP7_75t_L g778 ( 
.A1(n_642),
.A2(n_554),
.B(n_456),
.Y(n_778)
);

AND2x2_ASAP7_75t_L g779 ( 
.A(n_599),
.B(n_379),
.Y(n_779)
);

AOI21xp5_ASAP7_75t_L g780 ( 
.A1(n_665),
.A2(n_677),
.B(n_674),
.Y(n_780)
);

NOR2xp33_ASAP7_75t_L g781 ( 
.A(n_599),
.B(n_662),
.Y(n_781)
);

BUFx6f_ASAP7_75t_L g782 ( 
.A(n_686),
.Y(n_782)
);

BUFx6f_ASAP7_75t_L g783 ( 
.A(n_686),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_696),
.Y(n_784)
);

AOI21xp33_ASAP7_75t_L g785 ( 
.A1(n_662),
.A2(n_279),
.B(n_210),
.Y(n_785)
);

AOI21xp5_ASAP7_75t_L g786 ( 
.A1(n_677),
.A2(n_554),
.B(n_456),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_L g787 ( 
.A(n_638),
.B(n_463),
.Y(n_787)
);

AOI21xp5_ASAP7_75t_L g788 ( 
.A1(n_673),
.A2(n_526),
.B(n_554),
.Y(n_788)
);

INVx5_ASAP7_75t_L g789 ( 
.A(n_686),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_L g790 ( 
.A(n_645),
.B(n_706),
.Y(n_790)
);

AOI21xp5_ASAP7_75t_L g791 ( 
.A1(n_673),
.A2(n_526),
.B(n_558),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_706),
.B(n_463),
.Y(n_792)
);

OAI22xp5_ASAP7_75t_L g793 ( 
.A1(n_753),
.A2(n_555),
.B1(n_573),
.B2(n_571),
.Y(n_793)
);

O2A1O1Ixp5_ASAP7_75t_L g794 ( 
.A1(n_615),
.A2(n_538),
.B(n_573),
.C(n_571),
.Y(n_794)
);

HB1xp67_ASAP7_75t_L g795 ( 
.A(n_631),
.Y(n_795)
);

NOR2x1p5_ASAP7_75t_L g796 ( 
.A(n_733),
.B(n_212),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_598),
.B(n_600),
.Y(n_797)
);

AOI21xp5_ASAP7_75t_L g798 ( 
.A1(n_597),
.A2(n_526),
.B(n_537),
.Y(n_798)
);

OAI21xp5_ASAP7_75t_L g799 ( 
.A1(n_678),
.A2(n_487),
.B(n_464),
.Y(n_799)
);

AOI21xp5_ASAP7_75t_L g800 ( 
.A1(n_605),
.A2(n_580),
.B(n_543),
.Y(n_800)
);

AOI21x1_ASAP7_75t_L g801 ( 
.A1(n_682),
.A2(n_522),
.B(n_487),
.Y(n_801)
);

AOI21xp5_ASAP7_75t_L g802 ( 
.A1(n_633),
.A2(n_580),
.B(n_543),
.Y(n_802)
);

INVx2_ASAP7_75t_L g803 ( 
.A(n_704),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_L g804 ( 
.A(n_602),
.B(n_464),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_L g805 ( 
.A(n_607),
.B(n_476),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_L g806 ( 
.A(n_648),
.B(n_476),
.Y(n_806)
);

AOI21xp5_ASAP7_75t_L g807 ( 
.A1(n_633),
.A2(n_580),
.B(n_543),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_710),
.Y(n_808)
);

NOR2xp33_ASAP7_75t_L g809 ( 
.A(n_697),
.B(n_222),
.Y(n_809)
);

AOI21xp5_ASAP7_75t_L g810 ( 
.A1(n_678),
.A2(n_681),
.B(n_679),
.Y(n_810)
);

AOI21xp33_ASAP7_75t_L g811 ( 
.A1(n_651),
.A2(n_610),
.B(n_647),
.Y(n_811)
);

AOI21xp5_ASAP7_75t_L g812 ( 
.A1(n_679),
.A2(n_580),
.B(n_543),
.Y(n_812)
);

NOR2xp33_ASAP7_75t_L g813 ( 
.A(n_644),
.B(n_226),
.Y(n_813)
);

AND2x2_ASAP7_75t_L g814 ( 
.A(n_618),
.B(n_379),
.Y(n_814)
);

INVx4_ASAP7_75t_L g815 ( 
.A(n_686),
.Y(n_815)
);

AOI21xp5_ASAP7_75t_L g816 ( 
.A1(n_681),
.A2(n_580),
.B(n_472),
.Y(n_816)
);

AO21x1_ASAP7_75t_L g817 ( 
.A1(n_670),
.A2(n_405),
.B(n_506),
.Y(n_817)
);

INVx2_ASAP7_75t_L g818 ( 
.A(n_710),
.Y(n_818)
);

BUFx6f_ASAP7_75t_L g819 ( 
.A(n_734),
.Y(n_819)
);

INVx2_ASAP7_75t_SL g820 ( 
.A(n_623),
.Y(n_820)
);

BUFx6f_ASAP7_75t_L g821 ( 
.A(n_734),
.Y(n_821)
);

AOI21xp5_ASAP7_75t_L g822 ( 
.A1(n_652),
.A2(n_537),
.B(n_472),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_L g823 ( 
.A(n_655),
.B(n_482),
.Y(n_823)
);

AOI21xp5_ASAP7_75t_L g824 ( 
.A1(n_664),
.A2(n_543),
.B(n_537),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_L g825 ( 
.A(n_659),
.B(n_496),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_L g826 ( 
.A(n_666),
.B(n_522),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_L g827 ( 
.A(n_669),
.B(n_450),
.Y(n_827)
);

OAI22xp5_ASAP7_75t_L g828 ( 
.A1(n_620),
.A2(n_570),
.B1(n_569),
.B2(n_561),
.Y(n_828)
);

O2A1O1Ixp33_ASAP7_75t_L g829 ( 
.A1(n_745),
.A2(n_506),
.B(n_520),
.C(n_561),
.Y(n_829)
);

NOR2xp33_ASAP7_75t_L g830 ( 
.A(n_650),
.B(n_228),
.Y(n_830)
);

AOI21xp5_ASAP7_75t_L g831 ( 
.A1(n_688),
.A2(n_472),
.B(n_537),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_L g832 ( 
.A(n_689),
.B(n_455),
.Y(n_832)
);

O2A1O1Ixp33_ASAP7_75t_L g833 ( 
.A1(n_690),
.A2(n_520),
.B(n_569),
.C(n_555),
.Y(n_833)
);

INVx2_ASAP7_75t_L g834 ( 
.A(n_715),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_L g835 ( 
.A(n_736),
.B(n_538),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_730),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_SL g837 ( 
.A(n_640),
.B(n_537),
.Y(n_837)
);

AOI21xp5_ASAP7_75t_L g838 ( 
.A1(n_688),
.A2(n_515),
.B(n_455),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_L g839 ( 
.A(n_736),
.B(n_570),
.Y(n_839)
);

INVx1_ASAP7_75t_SL g840 ( 
.A(n_609),
.Y(n_840)
);

AOI21xp5_ASAP7_75t_L g841 ( 
.A1(n_682),
.A2(n_683),
.B(n_606),
.Y(n_841)
);

NOR2xp33_ASAP7_75t_L g842 ( 
.A(n_732),
.B(n_229),
.Y(n_842)
);

INVx2_ASAP7_75t_L g843 ( 
.A(n_731),
.Y(n_843)
);

OAI21x1_ASAP7_75t_L g844 ( 
.A1(n_758),
.A2(n_539),
.B(n_515),
.Y(n_844)
);

OAI21xp33_ASAP7_75t_L g845 ( 
.A1(n_728),
.A2(n_245),
.B(n_232),
.Y(n_845)
);

AOI21xp5_ASAP7_75t_L g846 ( 
.A1(n_683),
.A2(n_539),
.B(n_515),
.Y(n_846)
);

INVx4_ASAP7_75t_L g847 ( 
.A(n_640),
.Y(n_847)
);

O2A1O1Ixp5_ASAP7_75t_L g848 ( 
.A1(n_737),
.A2(n_539),
.B(n_485),
.C(n_385),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_731),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_702),
.B(n_485),
.Y(n_850)
);

OAI22xp5_ASAP7_75t_L g851 ( 
.A1(n_603),
.A2(n_485),
.B1(n_240),
.B2(n_278),
.Y(n_851)
);

AOI21xp5_ASAP7_75t_L g852 ( 
.A1(n_612),
.A2(n_479),
.B(n_546),
.Y(n_852)
);

AO21x1_ASAP7_75t_L g853 ( 
.A1(n_701),
.A2(n_402),
.B(n_387),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_749),
.Y(n_854)
);

AOI22xp5_ASAP7_75t_L g855 ( 
.A1(n_636),
.A2(n_398),
.B1(n_385),
.B2(n_387),
.Y(n_855)
);

AOI22xp33_ASAP7_75t_L g856 ( 
.A1(n_617),
.A2(n_398),
.B1(n_288),
.B2(n_235),
.Y(n_856)
);

AOI21xp5_ASAP7_75t_L g857 ( 
.A1(n_653),
.A2(n_479),
.B(n_546),
.Y(n_857)
);

AOI21xp5_ASAP7_75t_L g858 ( 
.A1(n_627),
.A2(n_479),
.B(n_546),
.Y(n_858)
);

BUFx6f_ASAP7_75t_L g859 ( 
.A(n_734),
.Y(n_859)
);

A2O1A1Ixp33_ASAP7_75t_L g860 ( 
.A1(n_619),
.A2(n_387),
.B(n_402),
.C(n_436),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_L g861 ( 
.A(n_703),
.B(n_398),
.Y(n_861)
);

OR2x6_ASAP7_75t_L g862 ( 
.A(n_621),
.B(n_436),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_SL g863 ( 
.A(n_640),
.B(n_288),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_711),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_712),
.B(n_398),
.Y(n_865)
);

BUFx12f_ASAP7_75t_L g866 ( 
.A(n_726),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_723),
.B(n_398),
.Y(n_867)
);

OAI22xp5_ASAP7_75t_L g868 ( 
.A1(n_619),
.A2(n_242),
.B1(n_249),
.B2(n_251),
.Y(n_868)
);

INVx2_ASAP7_75t_L g869 ( 
.A(n_611),
.Y(n_869)
);

AOI21x1_ASAP7_75t_L g870 ( 
.A1(n_680),
.A2(n_708),
.B(n_691),
.Y(n_870)
);

AOI21xp5_ASAP7_75t_L g871 ( 
.A1(n_627),
.A2(n_479),
.B(n_547),
.Y(n_871)
);

OAI21xp5_ASAP7_75t_L g872 ( 
.A1(n_635),
.A2(n_398),
.B(n_479),
.Y(n_872)
);

OAI22xp5_ASAP7_75t_L g873 ( 
.A1(n_625),
.A2(n_259),
.B1(n_263),
.B2(n_264),
.Y(n_873)
);

AOI21xp5_ASAP7_75t_L g874 ( 
.A1(n_639),
.A2(n_547),
.B(n_546),
.Y(n_874)
);

AOI21xp5_ASAP7_75t_L g875 ( 
.A1(n_639),
.A2(n_547),
.B(n_546),
.Y(n_875)
);

OAI21xp5_ASAP7_75t_L g876 ( 
.A1(n_637),
.A2(n_398),
.B(n_546),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_L g877 ( 
.A(n_729),
.B(n_402),
.Y(n_877)
);

NOR2xp33_ASAP7_75t_L g878 ( 
.A(n_760),
.B(n_280),
.Y(n_878)
);

OAI21xp5_ASAP7_75t_L g879 ( 
.A1(n_641),
.A2(n_547),
.B(n_391),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_738),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_SL g881 ( 
.A(n_640),
.B(n_288),
.Y(n_881)
);

AOI21xp5_ASAP7_75t_L g882 ( 
.A1(n_734),
.A2(n_547),
.B(n_390),
.Y(n_882)
);

A2O1A1Ixp33_ASAP7_75t_L g883 ( 
.A1(n_728),
.A2(n_755),
.B(n_757),
.C(n_707),
.Y(n_883)
);

AOI21xp5_ASAP7_75t_L g884 ( 
.A1(n_759),
.A2(n_547),
.B(n_390),
.Y(n_884)
);

AND2x4_ASAP7_75t_L g885 ( 
.A(n_654),
.B(n_484),
.Y(n_885)
);

O2A1O1Ixp33_ASAP7_75t_L g886 ( 
.A1(n_687),
.A2(n_447),
.B(n_443),
.C(n_439),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_SL g887 ( 
.A(n_657),
.B(n_288),
.Y(n_887)
);

NAND2xp33_ASAP7_75t_L g888 ( 
.A(n_759),
.B(n_289),
.Y(n_888)
);

AOI21xp5_ASAP7_75t_L g889 ( 
.A1(n_759),
.A2(n_390),
.B(n_386),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_L g890 ( 
.A(n_740),
.B(n_438),
.Y(n_890)
);

AND2x4_ASAP7_75t_L g891 ( 
.A(n_667),
.B(n_484),
.Y(n_891)
);

BUFx6f_ASAP7_75t_L g892 ( 
.A(n_759),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_L g893 ( 
.A(n_741),
.B(n_438),
.Y(n_893)
);

AOI21xp33_ASAP7_75t_L g894 ( 
.A1(n_617),
.A2(n_292),
.B(n_297),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_L g895 ( 
.A(n_643),
.B(n_444),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_L g896 ( 
.A(n_629),
.B(n_444),
.Y(n_896)
);

OAI22xp33_ASAP7_75t_L g897 ( 
.A1(n_752),
.A2(n_299),
.B1(n_301),
.B2(n_304),
.Y(n_897)
);

NOR2xp67_ASAP7_75t_L g898 ( 
.A(n_742),
.B(n_66),
.Y(n_898)
);

BUFx4f_ASAP7_75t_L g899 ( 
.A(n_743),
.Y(n_899)
);

AOI21xp5_ASAP7_75t_L g900 ( 
.A1(n_630),
.A2(n_386),
.B(n_390),
.Y(n_900)
);

INVx4_ASAP7_75t_L g901 ( 
.A(n_656),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_L g902 ( 
.A(n_705),
.B(n_438),
.Y(n_902)
);

AOI21xp5_ASAP7_75t_L g903 ( 
.A1(n_671),
.A2(n_386),
.B(n_390),
.Y(n_903)
);

AOI21xp5_ASAP7_75t_L g904 ( 
.A1(n_672),
.A2(n_386),
.B(n_390),
.Y(n_904)
);

AOI21xp5_ASAP7_75t_L g905 ( 
.A1(n_675),
.A2(n_386),
.B(n_390),
.Y(n_905)
);

NOR2xp33_ASAP7_75t_L g906 ( 
.A(n_746),
.B(n_4),
.Y(n_906)
);

HB1xp67_ASAP7_75t_L g907 ( 
.A(n_663),
.Y(n_907)
);

OAI21xp33_ASAP7_75t_L g908 ( 
.A1(n_754),
.A2(n_447),
.B(n_443),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_714),
.B(n_438),
.Y(n_909)
);

NOR2xp33_ASAP7_75t_L g910 ( 
.A(n_735),
.B(n_695),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_L g911 ( 
.A(n_611),
.B(n_438),
.Y(n_911)
);

AOI21xp5_ASAP7_75t_L g912 ( 
.A1(n_646),
.A2(n_386),
.B(n_390),
.Y(n_912)
);

INVx2_ASAP7_75t_SL g913 ( 
.A(n_663),
.Y(n_913)
);

INVx2_ASAP7_75t_L g914 ( 
.A(n_613),
.Y(n_914)
);

AOI21x1_ASAP7_75t_L g915 ( 
.A1(n_756),
.A2(n_447),
.B(n_443),
.Y(n_915)
);

AOI21xp5_ASAP7_75t_L g916 ( 
.A1(n_649),
.A2(n_386),
.B(n_390),
.Y(n_916)
);

AOI21xp5_ASAP7_75t_L g917 ( 
.A1(n_693),
.A2(n_694),
.B(n_699),
.Y(n_917)
);

INVx2_ASAP7_75t_L g918 ( 
.A(n_613),
.Y(n_918)
);

OAI21xp5_ASAP7_75t_L g919 ( 
.A1(n_685),
.A2(n_391),
.B(n_447),
.Y(n_919)
);

AOI21xp5_ASAP7_75t_L g920 ( 
.A1(n_700),
.A2(n_386),
.B(n_389),
.Y(n_920)
);

BUFx6f_ASAP7_75t_L g921 ( 
.A(n_663),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_L g922 ( 
.A(n_614),
.B(n_616),
.Y(n_922)
);

AND2x4_ASAP7_75t_SL g923 ( 
.A(n_743),
.B(n_443),
.Y(n_923)
);

NOR3xp33_ASAP7_75t_L g924 ( 
.A(n_624),
.B(n_439),
.C(n_436),
.Y(n_924)
);

AOI22xp33_ASAP7_75t_L g925 ( 
.A1(n_634),
.A2(n_444),
.B1(n_438),
.B2(n_439),
.Y(n_925)
);

BUFx2_ASAP7_75t_L g926 ( 
.A(n_726),
.Y(n_926)
);

AOI21xp5_ASAP7_75t_L g927 ( 
.A1(n_656),
.A2(n_386),
.B(n_389),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_L g928 ( 
.A(n_614),
.B(n_616),
.Y(n_928)
);

AOI22xp5_ASAP7_75t_L g929 ( 
.A1(n_757),
.A2(n_439),
.B1(n_436),
.B2(n_484),
.Y(n_929)
);

OAI21xp5_ASAP7_75t_L g930 ( 
.A1(n_718),
.A2(n_391),
.B(n_484),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_L g931 ( 
.A(n_626),
.B(n_444),
.Y(n_931)
);

OAI21xp5_ASAP7_75t_L g932 ( 
.A1(n_719),
.A2(n_391),
.B(n_389),
.Y(n_932)
);

AOI21x1_ASAP7_75t_L g933 ( 
.A1(n_721),
.A2(n_391),
.B(n_389),
.Y(n_933)
);

INVx2_ASAP7_75t_SL g934 ( 
.A(n_743),
.Y(n_934)
);

OAI21xp5_ASAP7_75t_L g935 ( 
.A1(n_725),
.A2(n_389),
.B(n_438),
.Y(n_935)
);

A2O1A1Ixp33_ASAP7_75t_L g936 ( 
.A1(n_744),
.A2(n_444),
.B(n_438),
.C(n_389),
.Y(n_936)
);

AOI21xp5_ASAP7_75t_L g937 ( 
.A1(n_727),
.A2(n_389),
.B(n_444),
.Y(n_937)
);

OAI21xp33_ASAP7_75t_L g938 ( 
.A1(n_737),
.A2(n_444),
.B(n_438),
.Y(n_938)
);

O2A1O1Ixp33_ASAP7_75t_L g939 ( 
.A1(n_752),
.A2(n_4),
.B(n_5),
.C(n_8),
.Y(n_939)
);

O2A1O1Ixp33_ASAP7_75t_L g940 ( 
.A1(n_752),
.A2(n_8),
.B(n_9),
.C(n_10),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_L g941 ( 
.A(n_626),
.B(n_444),
.Y(n_941)
);

AND2x4_ASAP7_75t_L g942 ( 
.A(n_913),
.B(n_761),
.Y(n_942)
);

O2A1O1Ixp33_ASAP7_75t_SL g943 ( 
.A1(n_883),
.A2(n_709),
.B(n_698),
.C(n_750),
.Y(n_943)
);

AND2x2_ASAP7_75t_L g944 ( 
.A(n_779),
.B(n_724),
.Y(n_944)
);

NOR2xp33_ASAP7_75t_L g945 ( 
.A(n_781),
.B(n_726),
.Y(n_945)
);

AOI22xp5_ASAP7_75t_L g946 ( 
.A1(n_910),
.A2(n_716),
.B1(n_720),
.B2(n_713),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_SL g947 ( 
.A(n_790),
.B(n_660),
.Y(n_947)
);

A2O1A1Ixp33_ASAP7_75t_SL g948 ( 
.A1(n_878),
.A2(n_748),
.B(n_660),
.C(n_692),
.Y(n_948)
);

INVx4_ASAP7_75t_L g949 ( 
.A(n_789),
.Y(n_949)
);

O2A1O1Ixp33_ASAP7_75t_L g950 ( 
.A1(n_785),
.A2(n_722),
.B(n_698),
.C(n_739),
.Y(n_950)
);

INVxp67_ASAP7_75t_L g951 ( 
.A(n_795),
.Y(n_951)
);

BUFx6f_ASAP7_75t_L g952 ( 
.A(n_782),
.Y(n_952)
);

BUFx6f_ASAP7_75t_L g953 ( 
.A(n_782),
.Y(n_953)
);

NAND2xp33_ASAP7_75t_R g954 ( 
.A(n_830),
.B(n_809),
.Y(n_954)
);

CKINVDCx20_ASAP7_75t_R g955 ( 
.A(n_926),
.Y(n_955)
);

AOI21xp5_ASAP7_75t_L g956 ( 
.A1(n_780),
.A2(n_751),
.B(n_747),
.Y(n_956)
);

NOR2x1p5_ASAP7_75t_L g957 ( 
.A(n_866),
.B(n_684),
.Y(n_957)
);

AND2x2_ASAP7_75t_L g958 ( 
.A(n_765),
.B(n_724),
.Y(n_958)
);

BUFx8_ASAP7_75t_SL g959 ( 
.A(n_899),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_SL g960 ( 
.A(n_767),
.B(n_692),
.Y(n_960)
);

AOI21xp5_ASAP7_75t_L g961 ( 
.A1(n_810),
.A2(n_628),
.B(n_762),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_784),
.Y(n_962)
);

OAI21xp5_ASAP7_75t_L g963 ( 
.A1(n_841),
.A2(n_822),
.B(n_800),
.Y(n_963)
);

NAND3xp33_ASAP7_75t_L g964 ( 
.A(n_906),
.B(n_722),
.C(n_628),
.Y(n_964)
);

NOR2xp33_ASAP7_75t_L g965 ( 
.A(n_772),
.B(n_11),
.Y(n_965)
);

AOI21xp5_ASAP7_75t_L g966 ( 
.A1(n_797),
.A2(n_389),
.B(n_724),
.Y(n_966)
);

AND2x2_ASAP7_75t_L g967 ( 
.A(n_842),
.B(n_813),
.Y(n_967)
);

AOI21xp5_ASAP7_75t_L g968 ( 
.A1(n_798),
.A2(n_389),
.B(n_444),
.Y(n_968)
);

BUFx2_ASAP7_75t_L g969 ( 
.A(n_840),
.Y(n_969)
);

OAI22xp5_ASAP7_75t_L g970 ( 
.A1(n_792),
.A2(n_839),
.B1(n_835),
.B2(n_768),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_L g971 ( 
.A(n_864),
.B(n_880),
.Y(n_971)
);

O2A1O1Ixp33_ASAP7_75t_L g972 ( 
.A1(n_811),
.A2(n_12),
.B(n_14),
.C(n_18),
.Y(n_972)
);

AND2x2_ASAP7_75t_SL g973 ( 
.A(n_899),
.B(n_151),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_SL g974 ( 
.A(n_921),
.B(n_143),
.Y(n_974)
);

AOI21xp5_ASAP7_75t_L g975 ( 
.A1(n_789),
.A2(n_123),
.B(n_122),
.Y(n_975)
);

NOR3xp33_ASAP7_75t_SL g976 ( 
.A(n_897),
.B(n_14),
.C(n_21),
.Y(n_976)
);

AOI21xp5_ASAP7_75t_SL g977 ( 
.A1(n_901),
.A2(n_121),
.B(n_117),
.Y(n_977)
);

AOI21xp5_ASAP7_75t_L g978 ( 
.A1(n_789),
.A2(n_115),
.B(n_113),
.Y(n_978)
);

A2O1A1Ixp33_ASAP7_75t_L g979 ( 
.A1(n_845),
.A2(n_23),
.B(n_24),
.C(n_25),
.Y(n_979)
);

OAI21xp5_ASAP7_75t_L g980 ( 
.A1(n_794),
.A2(n_112),
.B(n_98),
.Y(n_980)
);

NOR2xp33_ASAP7_75t_R g981 ( 
.A(n_782),
.B(n_89),
.Y(n_981)
);

CKINVDCx16_ASAP7_75t_R g982 ( 
.A(n_862),
.Y(n_982)
);

AOI21xp5_ASAP7_75t_L g983 ( 
.A1(n_789),
.A2(n_77),
.B(n_75),
.Y(n_983)
);

O2A1O1Ixp33_ASAP7_75t_L g984 ( 
.A1(n_764),
.A2(n_24),
.B(n_27),
.C(n_28),
.Y(n_984)
);

NOR2xp33_ASAP7_75t_L g985 ( 
.A(n_769),
.B(n_27),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_L g986 ( 
.A(n_773),
.B(n_28),
.Y(n_986)
);

AOI21xp5_ASAP7_75t_L g987 ( 
.A1(n_773),
.A2(n_70),
.B(n_67),
.Y(n_987)
);

AOI21xp5_ASAP7_75t_L g988 ( 
.A1(n_774),
.A2(n_30),
.B(n_33),
.Y(n_988)
);

INVx3_ASAP7_75t_L g989 ( 
.A(n_847),
.Y(n_989)
);

AOI22xp33_ASAP7_75t_L g990 ( 
.A1(n_808),
.A2(n_33),
.B1(n_34),
.B2(n_35),
.Y(n_990)
);

O2A1O1Ixp33_ASAP7_75t_L g991 ( 
.A1(n_894),
.A2(n_863),
.B(n_881),
.C(n_939),
.Y(n_991)
);

OR2x2_ASAP7_75t_L g992 ( 
.A(n_862),
.B(n_35),
.Y(n_992)
);

AOI21xp5_ASAP7_75t_L g993 ( 
.A1(n_774),
.A2(n_38),
.B(n_39),
.Y(n_993)
);

O2A1O1Ixp33_ASAP7_75t_L g994 ( 
.A1(n_940),
.A2(n_39),
.B(n_41),
.C(n_45),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_L g995 ( 
.A(n_836),
.B(n_45),
.Y(n_995)
);

NOR2xp33_ASAP7_75t_L g996 ( 
.A(n_907),
.B(n_49),
.Y(n_996)
);

AOI21xp5_ASAP7_75t_L g997 ( 
.A1(n_766),
.A2(n_49),
.B(n_52),
.Y(n_997)
);

A2O1A1Ixp33_ASAP7_75t_L g998 ( 
.A1(n_938),
.A2(n_52),
.B(n_54),
.C(n_56),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_L g999 ( 
.A(n_849),
.B(n_854),
.Y(n_999)
);

INVx1_ASAP7_75t_L g1000 ( 
.A(n_803),
.Y(n_1000)
);

NOR2xp33_ASAP7_75t_L g1001 ( 
.A(n_868),
.B(n_921),
.Y(n_1001)
);

O2A1O1Ixp33_ASAP7_75t_L g1002 ( 
.A1(n_887),
.A2(n_873),
.B(n_851),
.C(n_888),
.Y(n_1002)
);

OAI22xp5_ASAP7_75t_L g1003 ( 
.A1(n_835),
.A2(n_839),
.B1(n_768),
.B2(n_770),
.Y(n_1003)
);

NOR2xp33_ASAP7_75t_L g1004 ( 
.A(n_921),
.B(n_862),
.Y(n_1004)
);

AOI21xp5_ASAP7_75t_L g1005 ( 
.A1(n_775),
.A2(n_770),
.B(n_771),
.Y(n_1005)
);

AOI21xp5_ASAP7_75t_L g1006 ( 
.A1(n_771),
.A2(n_824),
.B(n_778),
.Y(n_1006)
);

AOI21xp5_ASAP7_75t_L g1007 ( 
.A1(n_788),
.A2(n_791),
.B(n_786),
.Y(n_1007)
);

NOR2xp33_ASAP7_75t_L g1008 ( 
.A(n_934),
.B(n_820),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_818),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_SL g1010 ( 
.A(n_847),
.B(n_783),
.Y(n_1010)
);

A2O1A1Ixp33_ASAP7_75t_L g1011 ( 
.A1(n_829),
.A2(n_898),
.B(n_936),
.C(n_917),
.Y(n_1011)
);

AOI22xp5_ASAP7_75t_L g1012 ( 
.A1(n_796),
.A2(n_891),
.B1(n_885),
.B2(n_856),
.Y(n_1012)
);

AOI221x1_ASAP7_75t_L g1013 ( 
.A1(n_776),
.A2(n_924),
.B1(n_908),
.B2(n_860),
.C(n_793),
.Y(n_1013)
);

AO21x2_ASAP7_75t_L g1014 ( 
.A1(n_853),
.A2(n_817),
.B(n_844),
.Y(n_1014)
);

AOI21xp5_ASAP7_75t_L g1015 ( 
.A1(n_763),
.A2(n_902),
.B(n_909),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_L g1016 ( 
.A(n_834),
.B(n_843),
.Y(n_1016)
);

HB1xp67_ASAP7_75t_L g1017 ( 
.A(n_819),
.Y(n_1017)
);

AOI21xp5_ASAP7_75t_L g1018 ( 
.A1(n_763),
.A2(n_909),
.B(n_902),
.Y(n_1018)
);

AOI22xp5_ASAP7_75t_L g1019 ( 
.A1(n_885),
.A2(n_891),
.B1(n_923),
.B2(n_814),
.Y(n_1019)
);

INVx2_ASAP7_75t_SL g1020 ( 
.A(n_783),
.Y(n_1020)
);

OAI22xp5_ASAP7_75t_L g1021 ( 
.A1(n_929),
.A2(n_870),
.B1(n_930),
.B2(n_825),
.Y(n_1021)
);

NAND2xp5_ASAP7_75t_L g1022 ( 
.A(n_922),
.B(n_928),
.Y(n_1022)
);

INVx1_ASAP7_75t_L g1023 ( 
.A(n_869),
.Y(n_1023)
);

INVx1_ASAP7_75t_L g1024 ( 
.A(n_914),
.Y(n_1024)
);

OAI22xp5_ASAP7_75t_L g1025 ( 
.A1(n_804),
.A2(n_806),
.B1(n_826),
.B2(n_823),
.Y(n_1025)
);

AOI21xp5_ASAP7_75t_L g1026 ( 
.A1(n_812),
.A2(n_816),
.B(n_837),
.Y(n_1026)
);

A2O1A1Ixp33_ASAP7_75t_L g1027 ( 
.A1(n_848),
.A2(n_861),
.B(n_865),
.C(n_867),
.Y(n_1027)
);

NOR2xp33_ASAP7_75t_L g1028 ( 
.A(n_805),
.B(n_850),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_918),
.Y(n_1029)
);

OR2x2_ASAP7_75t_L g1030 ( 
.A(n_877),
.B(n_787),
.Y(n_1030)
);

HB1xp67_ASAP7_75t_L g1031 ( 
.A(n_819),
.Y(n_1031)
);

AOI22xp5_ASAP7_75t_L g1032 ( 
.A1(n_861),
.A2(n_865),
.B1(n_867),
.B2(n_877),
.Y(n_1032)
);

INVx1_ASAP7_75t_L g1033 ( 
.A(n_922),
.Y(n_1033)
);

BUFx2_ASAP7_75t_L g1034 ( 
.A(n_819),
.Y(n_1034)
);

OAI22xp5_ASAP7_75t_L g1035 ( 
.A1(n_850),
.A2(n_901),
.B1(n_783),
.B2(n_928),
.Y(n_1035)
);

INVx1_ASAP7_75t_L g1036 ( 
.A(n_890),
.Y(n_1036)
);

OAI22xp5_ASAP7_75t_SL g1037 ( 
.A1(n_815),
.A2(n_859),
.B1(n_892),
.B2(n_821),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_SL g1038 ( 
.A(n_815),
.B(n_821),
.Y(n_1038)
);

NAND2xp5_ASAP7_75t_L g1039 ( 
.A(n_895),
.B(n_832),
.Y(n_1039)
);

NAND2x1p5_ASAP7_75t_L g1040 ( 
.A(n_821),
.B(n_892),
.Y(n_1040)
);

NAND2xp5_ASAP7_75t_SL g1041 ( 
.A(n_859),
.B(n_892),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_L g1042 ( 
.A(n_895),
.B(n_827),
.Y(n_1042)
);

NOR2xp33_ASAP7_75t_L g1043 ( 
.A(n_893),
.B(n_859),
.Y(n_1043)
);

INVx1_ASAP7_75t_L g1044 ( 
.A(n_911),
.Y(n_1044)
);

BUFx2_ASAP7_75t_L g1045 ( 
.A(n_799),
.Y(n_1045)
);

NOR2xp33_ASAP7_75t_L g1046 ( 
.A(n_896),
.B(n_828),
.Y(n_1046)
);

NOR3xp33_ASAP7_75t_SL g1047 ( 
.A(n_872),
.B(n_876),
.C(n_831),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_L g1048 ( 
.A(n_896),
.B(n_941),
.Y(n_1048)
);

NAND2xp5_ASAP7_75t_L g1049 ( 
.A(n_911),
.B(n_941),
.Y(n_1049)
);

OAI21xp33_ASAP7_75t_L g1050 ( 
.A1(n_855),
.A2(n_931),
.B(n_925),
.Y(n_1050)
);

AOI21xp5_ASAP7_75t_L g1051 ( 
.A1(n_802),
.A2(n_807),
.B(n_879),
.Y(n_1051)
);

OAI22xp5_ASAP7_75t_L g1052 ( 
.A1(n_932),
.A2(n_838),
.B1(n_846),
.B2(n_935),
.Y(n_1052)
);

AND2x4_ASAP7_75t_L g1053 ( 
.A(n_915),
.B(n_801),
.Y(n_1053)
);

OAI22xp5_ASAP7_75t_L g1054 ( 
.A1(n_919),
.A2(n_931),
.B1(n_833),
.B2(n_916),
.Y(n_1054)
);

AND2x4_ASAP7_75t_L g1055 ( 
.A(n_933),
.B(n_912),
.Y(n_1055)
);

AND2x4_ASAP7_75t_L g1056 ( 
.A(n_857),
.B(n_905),
.Y(n_1056)
);

INVx2_ASAP7_75t_L g1057 ( 
.A(n_886),
.Y(n_1057)
);

HB1xp67_ASAP7_75t_L g1058 ( 
.A(n_903),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_904),
.Y(n_1059)
);

NOR2xp33_ASAP7_75t_L g1060 ( 
.A(n_900),
.B(n_920),
.Y(n_1060)
);

NAND2xp5_ASAP7_75t_SL g1061 ( 
.A(n_852),
.B(n_937),
.Y(n_1061)
);

AOI21xp5_ASAP7_75t_L g1062 ( 
.A1(n_927),
.A2(n_858),
.B(n_871),
.Y(n_1062)
);

AND3x1_ASAP7_75t_L g1063 ( 
.A(n_889),
.B(n_882),
.C(n_884),
.Y(n_1063)
);

INVx3_ASAP7_75t_L g1064 ( 
.A(n_874),
.Y(n_1064)
);

NOR2xp33_ASAP7_75t_L g1065 ( 
.A(n_875),
.B(n_781),
.Y(n_1065)
);

O2A1O1Ixp33_ASAP7_75t_SL g1066 ( 
.A1(n_883),
.A2(n_764),
.B(n_615),
.C(n_781),
.Y(n_1066)
);

NAND2xp5_ASAP7_75t_L g1067 ( 
.A(n_781),
.B(n_601),
.Y(n_1067)
);

BUFx2_ASAP7_75t_R g1068 ( 
.A(n_926),
.Y(n_1068)
);

AOI21xp5_ASAP7_75t_L g1069 ( 
.A1(n_777),
.A2(n_633),
.B(n_591),
.Y(n_1069)
);

INVx1_ASAP7_75t_L g1070 ( 
.A(n_784),
.Y(n_1070)
);

NOR2xp33_ASAP7_75t_L g1071 ( 
.A(n_781),
.B(n_601),
.Y(n_1071)
);

AND2x4_ASAP7_75t_L g1072 ( 
.A(n_913),
.B(n_907),
.Y(n_1072)
);

O2A1O1Ixp33_ASAP7_75t_L g1073 ( 
.A1(n_781),
.A2(n_785),
.B(n_608),
.C(n_615),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_L g1074 ( 
.A(n_781),
.B(n_601),
.Y(n_1074)
);

BUFx3_ASAP7_75t_L g1075 ( 
.A(n_866),
.Y(n_1075)
);

NAND2xp5_ASAP7_75t_SL g1076 ( 
.A(n_781),
.B(n_601),
.Y(n_1076)
);

NAND2xp5_ASAP7_75t_L g1077 ( 
.A(n_1071),
.B(n_1067),
.Y(n_1077)
);

INVx2_ASAP7_75t_L g1078 ( 
.A(n_962),
.Y(n_1078)
);

CKINVDCx5p33_ASAP7_75t_R g1079 ( 
.A(n_959),
.Y(n_1079)
);

INVx6_ASAP7_75t_L g1080 ( 
.A(n_982),
.Y(n_1080)
);

O2A1O1Ixp33_ASAP7_75t_SL g1081 ( 
.A1(n_979),
.A2(n_998),
.B(n_1011),
.C(n_986),
.Y(n_1081)
);

INVx1_ASAP7_75t_L g1082 ( 
.A(n_971),
.Y(n_1082)
);

BUFx2_ASAP7_75t_L g1083 ( 
.A(n_969),
.Y(n_1083)
);

NAND2xp5_ASAP7_75t_L g1084 ( 
.A(n_1074),
.B(n_1076),
.Y(n_1084)
);

OR2x2_ASAP7_75t_L g1085 ( 
.A(n_951),
.B(n_967),
.Y(n_1085)
);

OAI21xp5_ASAP7_75t_L g1086 ( 
.A1(n_1046),
.A2(n_1018),
.B(n_1015),
.Y(n_1086)
);

AOI21xp5_ASAP7_75t_L g1087 ( 
.A1(n_1005),
.A2(n_1006),
.B(n_1007),
.Y(n_1087)
);

AND2x2_ASAP7_75t_L g1088 ( 
.A(n_945),
.B(n_958),
.Y(n_1088)
);

OAI21x1_ASAP7_75t_L g1089 ( 
.A1(n_1062),
.A2(n_968),
.B(n_961),
.Y(n_1089)
);

BUFx2_ASAP7_75t_SL g1090 ( 
.A(n_955),
.Y(n_1090)
);

OAI21xp5_ASAP7_75t_L g1091 ( 
.A1(n_1046),
.A2(n_1065),
.B(n_966),
.Y(n_1091)
);

AOI22xp33_ASAP7_75t_L g1092 ( 
.A1(n_965),
.A2(n_985),
.B1(n_942),
.B2(n_944),
.Y(n_1092)
);

AOI21xp5_ASAP7_75t_L g1093 ( 
.A1(n_963),
.A2(n_970),
.B(n_1003),
.Y(n_1093)
);

AOI21xp5_ASAP7_75t_L g1094 ( 
.A1(n_1051),
.A2(n_1060),
.B(n_1066),
.Y(n_1094)
);

AND2x2_ASAP7_75t_L g1095 ( 
.A(n_945),
.B(n_951),
.Y(n_1095)
);

NAND2xp5_ASAP7_75t_L g1096 ( 
.A(n_965),
.B(n_1033),
.Y(n_1096)
);

AOI21xp5_ASAP7_75t_L g1097 ( 
.A1(n_1060),
.A2(n_1065),
.B(n_1069),
.Y(n_1097)
);

OR2x2_ASAP7_75t_L g1098 ( 
.A(n_942),
.B(n_1072),
.Y(n_1098)
);

AOI21xp5_ASAP7_75t_L g1099 ( 
.A1(n_1022),
.A2(n_1054),
.B(n_1021),
.Y(n_1099)
);

AOI22xp5_ASAP7_75t_L g1100 ( 
.A1(n_954),
.A2(n_985),
.B1(n_1001),
.B2(n_973),
.Y(n_1100)
);

NAND2xp5_ASAP7_75t_L g1101 ( 
.A(n_1030),
.B(n_1028),
.Y(n_1101)
);

BUFx4_ASAP7_75t_SL g1102 ( 
.A(n_1075),
.Y(n_1102)
);

INVx1_ASAP7_75t_L g1103 ( 
.A(n_1070),
.Y(n_1103)
);

NOR2x1_ASAP7_75t_SL g1104 ( 
.A(n_949),
.B(n_1035),
.Y(n_1104)
);

INVx1_ASAP7_75t_L g1105 ( 
.A(n_1023),
.Y(n_1105)
);

AOI21xp5_ASAP7_75t_L g1106 ( 
.A1(n_1039),
.A2(n_1042),
.B(n_1052),
.Y(n_1106)
);

AND2x4_ASAP7_75t_L g1107 ( 
.A(n_1072),
.B(n_1004),
.Y(n_1107)
);

OAI21x1_ASAP7_75t_L g1108 ( 
.A1(n_1026),
.A2(n_956),
.B(n_1061),
.Y(n_1108)
);

OAI22xp5_ASAP7_75t_L g1109 ( 
.A1(n_990),
.A2(n_973),
.B1(n_946),
.B2(n_1019),
.Y(n_1109)
);

NAND2xp5_ASAP7_75t_SL g1110 ( 
.A(n_1073),
.B(n_1001),
.Y(n_1110)
);

AND2x2_ASAP7_75t_L g1111 ( 
.A(n_996),
.B(n_992),
.Y(n_1111)
);

INVx1_ASAP7_75t_SL g1112 ( 
.A(n_1034),
.Y(n_1112)
);

AOI221x1_ASAP7_75t_L g1113 ( 
.A1(n_997),
.A2(n_988),
.B1(n_993),
.B2(n_980),
.C(n_1056),
.Y(n_1113)
);

AOI22xp5_ASAP7_75t_L g1114 ( 
.A1(n_996),
.A2(n_1012),
.B1(n_976),
.B2(n_990),
.Y(n_1114)
);

AOI21xp5_ASAP7_75t_L g1115 ( 
.A1(n_1025),
.A2(n_1048),
.B(n_1058),
.Y(n_1115)
);

NAND2xp5_ASAP7_75t_L g1116 ( 
.A(n_1036),
.B(n_1044),
.Y(n_1116)
);

AO32x2_ASAP7_75t_L g1117 ( 
.A1(n_1037),
.A2(n_1014),
.A3(n_976),
.B1(n_994),
.B2(n_1020),
.Y(n_1117)
);

OA21x2_ASAP7_75t_L g1118 ( 
.A1(n_1013),
.A2(n_1059),
.B(n_1027),
.Y(n_1118)
);

O2A1O1Ixp33_ASAP7_75t_SL g1119 ( 
.A1(n_974),
.A2(n_948),
.B(n_960),
.C(n_947),
.Y(n_1119)
);

OAI22xp5_ASAP7_75t_L g1120 ( 
.A1(n_1045),
.A2(n_964),
.B1(n_999),
.B2(n_1050),
.Y(n_1120)
);

AOI21xp5_ASAP7_75t_L g1121 ( 
.A1(n_1058),
.A2(n_943),
.B(n_1056),
.Y(n_1121)
);

AOI22xp5_ASAP7_75t_L g1122 ( 
.A1(n_995),
.A2(n_1009),
.B1(n_1000),
.B2(n_1008),
.Y(n_1122)
);

NAND2xp5_ASAP7_75t_L g1123 ( 
.A(n_1043),
.B(n_1049),
.Y(n_1123)
);

AOI21xp5_ASAP7_75t_L g1124 ( 
.A1(n_1055),
.A2(n_950),
.B(n_1002),
.Y(n_1124)
);

AOI21x1_ASAP7_75t_L g1125 ( 
.A1(n_1055),
.A2(n_1053),
.B(n_1057),
.Y(n_1125)
);

O2A1O1Ixp5_ASAP7_75t_SL g1126 ( 
.A1(n_1064),
.A2(n_1041),
.B(n_1024),
.C(n_1029),
.Y(n_1126)
);

OAI22xp5_ASAP7_75t_L g1127 ( 
.A1(n_1043),
.A2(n_1032),
.B1(n_991),
.B2(n_1016),
.Y(n_1127)
);

OAI21x1_ASAP7_75t_L g1128 ( 
.A1(n_1063),
.A2(n_987),
.B(n_983),
.Y(n_1128)
);

A2O1A1Ixp33_ASAP7_75t_L g1129 ( 
.A1(n_972),
.A2(n_984),
.B(n_1047),
.C(n_978),
.Y(n_1129)
);

AOI21xp5_ASAP7_75t_L g1130 ( 
.A1(n_949),
.A2(n_1053),
.B(n_1014),
.Y(n_1130)
);

A2O1A1Ixp33_ASAP7_75t_L g1131 ( 
.A1(n_1047),
.A2(n_975),
.B(n_989),
.C(n_1010),
.Y(n_1131)
);

OAI21xp5_ASAP7_75t_L g1132 ( 
.A1(n_977),
.A2(n_1038),
.B(n_1017),
.Y(n_1132)
);

AOI221x1_ASAP7_75t_L g1133 ( 
.A1(n_989),
.A2(n_952),
.B1(n_953),
.B2(n_981),
.C(n_1068),
.Y(n_1133)
);

OAI21x1_ASAP7_75t_L g1134 ( 
.A1(n_1040),
.A2(n_1017),
.B(n_1031),
.Y(n_1134)
);

AO22x2_ASAP7_75t_L g1135 ( 
.A1(n_1031),
.A2(n_1040),
.B1(n_953),
.B2(n_952),
.Y(n_1135)
);

AOI21x1_ASAP7_75t_L g1136 ( 
.A1(n_952),
.A2(n_953),
.B(n_957),
.Y(n_1136)
);

OAI21xp5_ASAP7_75t_L g1137 ( 
.A1(n_1046),
.A2(n_781),
.B(n_883),
.Y(n_1137)
);

BUFx2_ASAP7_75t_L g1138 ( 
.A(n_969),
.Y(n_1138)
);

AOI21xp5_ASAP7_75t_L g1139 ( 
.A1(n_1005),
.A2(n_1011),
.B(n_1015),
.Y(n_1139)
);

NAND2xp5_ASAP7_75t_L g1140 ( 
.A(n_1071),
.B(n_1067),
.Y(n_1140)
);

OA21x2_ASAP7_75t_L g1141 ( 
.A1(n_963),
.A2(n_1005),
.B(n_1006),
.Y(n_1141)
);

NAND3xp33_ASAP7_75t_SL g1142 ( 
.A(n_1071),
.B(n_781),
.C(n_967),
.Y(n_1142)
);

INVx1_ASAP7_75t_SL g1143 ( 
.A(n_969),
.Y(n_1143)
);

INVx3_ASAP7_75t_L g1144 ( 
.A(n_949),
.Y(n_1144)
);

OAI21x1_ASAP7_75t_L g1145 ( 
.A1(n_1062),
.A2(n_844),
.B(n_968),
.Y(n_1145)
);

AND2x2_ASAP7_75t_L g1146 ( 
.A(n_1071),
.B(n_604),
.Y(n_1146)
);

AND2x2_ASAP7_75t_L g1147 ( 
.A(n_1071),
.B(n_604),
.Y(n_1147)
);

AND2x2_ASAP7_75t_L g1148 ( 
.A(n_1071),
.B(n_604),
.Y(n_1148)
);

AND2x2_ASAP7_75t_L g1149 ( 
.A(n_1071),
.B(n_604),
.Y(n_1149)
);

INVx1_ASAP7_75t_L g1150 ( 
.A(n_971),
.Y(n_1150)
);

NAND2xp5_ASAP7_75t_L g1151 ( 
.A(n_1071),
.B(n_1067),
.Y(n_1151)
);

AOI21xp5_ASAP7_75t_L g1152 ( 
.A1(n_1005),
.A2(n_1011),
.B(n_1015),
.Y(n_1152)
);

AO32x2_ASAP7_75t_L g1153 ( 
.A1(n_1003),
.A2(n_970),
.A3(n_1054),
.B1(n_1021),
.B2(n_690),
.Y(n_1153)
);

AOI221xp5_ASAP7_75t_L g1154 ( 
.A1(n_1071),
.A2(n_781),
.B1(n_599),
.B2(n_1074),
.C(n_1067),
.Y(n_1154)
);

OAI21x1_ASAP7_75t_L g1155 ( 
.A1(n_1062),
.A2(n_844),
.B(n_968),
.Y(n_1155)
);

INVx3_ASAP7_75t_L g1156 ( 
.A(n_949),
.Y(n_1156)
);

AO32x2_ASAP7_75t_L g1157 ( 
.A1(n_1003),
.A2(n_970),
.A3(n_1054),
.B1(n_1021),
.B2(n_690),
.Y(n_1157)
);

NAND3xp33_ASAP7_75t_SL g1158 ( 
.A(n_1071),
.B(n_781),
.C(n_967),
.Y(n_1158)
);

AOI21xp5_ASAP7_75t_L g1159 ( 
.A1(n_1005),
.A2(n_1011),
.B(n_1015),
.Y(n_1159)
);

NAND2xp5_ASAP7_75t_L g1160 ( 
.A(n_1071),
.B(n_1067),
.Y(n_1160)
);

AO32x2_ASAP7_75t_L g1161 ( 
.A1(n_1003),
.A2(n_970),
.A3(n_1054),
.B1(n_1021),
.B2(n_690),
.Y(n_1161)
);

OAI21x1_ASAP7_75t_L g1162 ( 
.A1(n_1062),
.A2(n_844),
.B(n_968),
.Y(n_1162)
);

INVxp67_ASAP7_75t_L g1163 ( 
.A(n_969),
.Y(n_1163)
);

CKINVDCx5p33_ASAP7_75t_R g1164 ( 
.A(n_959),
.Y(n_1164)
);

NOR2xp33_ASAP7_75t_L g1165 ( 
.A(n_1071),
.B(n_781),
.Y(n_1165)
);

AOI21xp5_ASAP7_75t_L g1166 ( 
.A1(n_1005),
.A2(n_1011),
.B(n_1015),
.Y(n_1166)
);

O2A1O1Ixp33_ASAP7_75t_SL g1167 ( 
.A1(n_979),
.A2(n_883),
.B(n_998),
.C(n_781),
.Y(n_1167)
);

NAND2xp5_ASAP7_75t_L g1168 ( 
.A(n_1071),
.B(n_1067),
.Y(n_1168)
);

AOI21xp5_ASAP7_75t_L g1169 ( 
.A1(n_1005),
.A2(n_1011),
.B(n_1015),
.Y(n_1169)
);

NAND2xp5_ASAP7_75t_L g1170 ( 
.A(n_1071),
.B(n_1067),
.Y(n_1170)
);

OAI21xp5_ASAP7_75t_L g1171 ( 
.A1(n_1046),
.A2(n_781),
.B(n_883),
.Y(n_1171)
);

BUFx12f_ASAP7_75t_L g1172 ( 
.A(n_957),
.Y(n_1172)
);

AOI21xp5_ASAP7_75t_L g1173 ( 
.A1(n_1005),
.A2(n_1011),
.B(n_1015),
.Y(n_1173)
);

CKINVDCx8_ASAP7_75t_R g1174 ( 
.A(n_969),
.Y(n_1174)
);

INVx1_ASAP7_75t_L g1175 ( 
.A(n_971),
.Y(n_1175)
);

NAND2xp5_ASAP7_75t_L g1176 ( 
.A(n_1071),
.B(n_1067),
.Y(n_1176)
);

AO32x2_ASAP7_75t_L g1177 ( 
.A1(n_1003),
.A2(n_970),
.A3(n_1054),
.B1(n_1021),
.B2(n_690),
.Y(n_1177)
);

O2A1O1Ixp33_ASAP7_75t_SL g1178 ( 
.A1(n_979),
.A2(n_883),
.B(n_998),
.C(n_781),
.Y(n_1178)
);

OAI21x1_ASAP7_75t_L g1179 ( 
.A1(n_1062),
.A2(n_844),
.B(n_968),
.Y(n_1179)
);

AO31x2_ASAP7_75t_L g1180 ( 
.A1(n_1054),
.A2(n_853),
.A3(n_817),
.B(n_1011),
.Y(n_1180)
);

O2A1O1Ixp33_ASAP7_75t_SL g1181 ( 
.A1(n_979),
.A2(n_883),
.B(n_998),
.C(n_781),
.Y(n_1181)
);

INVx1_ASAP7_75t_L g1182 ( 
.A(n_971),
.Y(n_1182)
);

AOI21xp5_ASAP7_75t_L g1183 ( 
.A1(n_1005),
.A2(n_1011),
.B(n_1015),
.Y(n_1183)
);

NAND2xp5_ASAP7_75t_L g1184 ( 
.A(n_1071),
.B(n_1067),
.Y(n_1184)
);

O2A1O1Ixp33_ASAP7_75t_L g1185 ( 
.A1(n_1071),
.A2(n_781),
.B(n_1074),
.C(n_1067),
.Y(n_1185)
);

INVx1_ASAP7_75t_L g1186 ( 
.A(n_971),
.Y(n_1186)
);

OA21x2_ASAP7_75t_L g1187 ( 
.A1(n_963),
.A2(n_1005),
.B(n_1006),
.Y(n_1187)
);

AOI221xp5_ASAP7_75t_SL g1188 ( 
.A1(n_979),
.A2(n_781),
.B1(n_998),
.B2(n_745),
.C(n_965),
.Y(n_1188)
);

BUFx2_ASAP7_75t_R g1189 ( 
.A(n_959),
.Y(n_1189)
);

A2O1A1Ixp33_ASAP7_75t_L g1190 ( 
.A1(n_1073),
.A2(n_781),
.B(n_1071),
.C(n_830),
.Y(n_1190)
);

NAND2xp5_ASAP7_75t_L g1191 ( 
.A(n_1071),
.B(n_1067),
.Y(n_1191)
);

NOR2xp33_ASAP7_75t_L g1192 ( 
.A(n_1071),
.B(n_781),
.Y(n_1192)
);

NAND3xp33_ASAP7_75t_SL g1193 ( 
.A(n_1071),
.B(n_781),
.C(n_967),
.Y(n_1193)
);

NAND2xp5_ASAP7_75t_L g1194 ( 
.A(n_1071),
.B(n_1067),
.Y(n_1194)
);

INVx1_ASAP7_75t_L g1195 ( 
.A(n_971),
.Y(n_1195)
);

INVx1_ASAP7_75t_L g1196 ( 
.A(n_971),
.Y(n_1196)
);

NOR2xp33_ASAP7_75t_L g1197 ( 
.A(n_1071),
.B(n_781),
.Y(n_1197)
);

OR2x2_ASAP7_75t_L g1198 ( 
.A(n_1067),
.B(n_1074),
.Y(n_1198)
);

AO31x2_ASAP7_75t_L g1199 ( 
.A1(n_1054),
.A2(n_853),
.A3(n_817),
.B(n_1011),
.Y(n_1199)
);

BUFx6f_ASAP7_75t_L g1200 ( 
.A(n_952),
.Y(n_1200)
);

OAI21x1_ASAP7_75t_L g1201 ( 
.A1(n_1062),
.A2(n_844),
.B(n_968),
.Y(n_1201)
);

AND2x4_ASAP7_75t_L g1202 ( 
.A(n_1072),
.B(n_942),
.Y(n_1202)
);

INVx2_ASAP7_75t_SL g1203 ( 
.A(n_969),
.Y(n_1203)
);

NOR2x1_ASAP7_75t_R g1204 ( 
.A(n_1075),
.B(n_866),
.Y(n_1204)
);

INVx3_ASAP7_75t_SL g1205 ( 
.A(n_955),
.Y(n_1205)
);

AND2x4_ASAP7_75t_L g1206 ( 
.A(n_1072),
.B(n_942),
.Y(n_1206)
);

BUFx2_ASAP7_75t_L g1207 ( 
.A(n_969),
.Y(n_1207)
);

CKINVDCx11_ASAP7_75t_R g1208 ( 
.A(n_955),
.Y(n_1208)
);

AO31x2_ASAP7_75t_L g1209 ( 
.A1(n_1054),
.A2(n_853),
.A3(n_817),
.B(n_1011),
.Y(n_1209)
);

NAND2xp5_ASAP7_75t_L g1210 ( 
.A(n_1071),
.B(n_1067),
.Y(n_1210)
);

AND2x6_ASAP7_75t_L g1211 ( 
.A(n_989),
.B(n_1033),
.Y(n_1211)
);

HB1xp67_ASAP7_75t_L g1212 ( 
.A(n_969),
.Y(n_1212)
);

OAI21x1_ASAP7_75t_L g1213 ( 
.A1(n_1062),
.A2(n_844),
.B(n_968),
.Y(n_1213)
);

INVx6_ASAP7_75t_L g1214 ( 
.A(n_1080),
.Y(n_1214)
);

INVx6_ASAP7_75t_L g1215 ( 
.A(n_1080),
.Y(n_1215)
);

CKINVDCx16_ASAP7_75t_R g1216 ( 
.A(n_1172),
.Y(n_1216)
);

AOI22xp33_ASAP7_75t_L g1217 ( 
.A1(n_1165),
.A2(n_1197),
.B1(n_1192),
.B2(n_1154),
.Y(n_1217)
);

CKINVDCx5p33_ASAP7_75t_R g1218 ( 
.A(n_1208),
.Y(n_1218)
);

AOI22xp33_ASAP7_75t_L g1219 ( 
.A1(n_1142),
.A2(n_1193),
.B1(n_1158),
.B2(n_1171),
.Y(n_1219)
);

INVx6_ASAP7_75t_L g1220 ( 
.A(n_1200),
.Y(n_1220)
);

CKINVDCx6p67_ASAP7_75t_R g1221 ( 
.A(n_1205),
.Y(n_1221)
);

NAND2xp5_ASAP7_75t_L g1222 ( 
.A(n_1151),
.B(n_1168),
.Y(n_1222)
);

OAI22xp5_ASAP7_75t_L g1223 ( 
.A1(n_1100),
.A2(n_1190),
.B1(n_1101),
.B2(n_1210),
.Y(n_1223)
);

CKINVDCx11_ASAP7_75t_R g1224 ( 
.A(n_1174),
.Y(n_1224)
);

OAI22xp33_ASAP7_75t_L g1225 ( 
.A1(n_1100),
.A2(n_1114),
.B1(n_1077),
.B2(n_1140),
.Y(n_1225)
);

INVx1_ASAP7_75t_SL g1226 ( 
.A(n_1143),
.Y(n_1226)
);

HB1xp67_ASAP7_75t_L g1227 ( 
.A(n_1125),
.Y(n_1227)
);

OAI22xp5_ASAP7_75t_L g1228 ( 
.A1(n_1170),
.A2(n_1176),
.B1(n_1184),
.B2(n_1191),
.Y(n_1228)
);

AOI22xp33_ASAP7_75t_SL g1229 ( 
.A1(n_1109),
.A2(n_1137),
.B1(n_1171),
.B2(n_1194),
.Y(n_1229)
);

INVxp67_ASAP7_75t_L g1230 ( 
.A(n_1212),
.Y(n_1230)
);

INVx6_ASAP7_75t_L g1231 ( 
.A(n_1200),
.Y(n_1231)
);

AOI22xp33_ASAP7_75t_L g1232 ( 
.A1(n_1137),
.A2(n_1109),
.B1(n_1110),
.B2(n_1114),
.Y(n_1232)
);

AOI22xp33_ASAP7_75t_L g1233 ( 
.A1(n_1077),
.A2(n_1140),
.B1(n_1160),
.B2(n_1091),
.Y(n_1233)
);

AOI22xp33_ASAP7_75t_SL g1234 ( 
.A1(n_1160),
.A2(n_1111),
.B1(n_1086),
.B2(n_1093),
.Y(n_1234)
);

AOI22xp33_ASAP7_75t_L g1235 ( 
.A1(n_1091),
.A2(n_1092),
.B1(n_1147),
.B2(n_1146),
.Y(n_1235)
);

INVx4_ASAP7_75t_L g1236 ( 
.A(n_1138),
.Y(n_1236)
);

AND2x2_ASAP7_75t_L g1237 ( 
.A(n_1148),
.B(n_1149),
.Y(n_1237)
);

INVx1_ASAP7_75t_L g1238 ( 
.A(n_1103),
.Y(n_1238)
);

INVx6_ASAP7_75t_L g1239 ( 
.A(n_1107),
.Y(n_1239)
);

INVx1_ASAP7_75t_L g1240 ( 
.A(n_1105),
.Y(n_1240)
);

CKINVDCx11_ASAP7_75t_R g1241 ( 
.A(n_1143),
.Y(n_1241)
);

CKINVDCx6p67_ASAP7_75t_R g1242 ( 
.A(n_1090),
.Y(n_1242)
);

CKINVDCx6p67_ASAP7_75t_R g1243 ( 
.A(n_1207),
.Y(n_1243)
);

AOI22xp33_ASAP7_75t_SL g1244 ( 
.A1(n_1086),
.A2(n_1088),
.B1(n_1096),
.B2(n_1095),
.Y(n_1244)
);

CKINVDCx11_ASAP7_75t_R g1245 ( 
.A(n_1112),
.Y(n_1245)
);

CKINVDCx11_ASAP7_75t_R g1246 ( 
.A(n_1112),
.Y(n_1246)
);

INVx4_ASAP7_75t_L g1247 ( 
.A(n_1079),
.Y(n_1247)
);

CKINVDCx11_ASAP7_75t_R g1248 ( 
.A(n_1102),
.Y(n_1248)
);

OAI22xp5_ASAP7_75t_L g1249 ( 
.A1(n_1198),
.A2(n_1185),
.B1(n_1085),
.B2(n_1182),
.Y(n_1249)
);

OAI22xp5_ASAP7_75t_L g1250 ( 
.A1(n_1082),
.A2(n_1186),
.B1(n_1196),
.B2(n_1150),
.Y(n_1250)
);

NAND2xp5_ASAP7_75t_L g1251 ( 
.A(n_1084),
.B(n_1175),
.Y(n_1251)
);

BUFx3_ASAP7_75t_L g1252 ( 
.A(n_1203),
.Y(n_1252)
);

AOI22xp33_ASAP7_75t_L g1253 ( 
.A1(n_1195),
.A2(n_1120),
.B1(n_1127),
.B2(n_1099),
.Y(n_1253)
);

BUFx6f_ASAP7_75t_L g1254 ( 
.A(n_1107),
.Y(n_1254)
);

AOI22xp33_ASAP7_75t_L g1255 ( 
.A1(n_1120),
.A2(n_1127),
.B1(n_1097),
.B2(n_1123),
.Y(n_1255)
);

BUFx2_ASAP7_75t_L g1256 ( 
.A(n_1202),
.Y(n_1256)
);

INVx1_ASAP7_75t_SL g1257 ( 
.A(n_1098),
.Y(n_1257)
);

AND2x2_ASAP7_75t_L g1258 ( 
.A(n_1202),
.B(n_1206),
.Y(n_1258)
);

INVx4_ASAP7_75t_L g1259 ( 
.A(n_1164),
.Y(n_1259)
);

BUFx8_ASAP7_75t_L g1260 ( 
.A(n_1189),
.Y(n_1260)
);

OAI22xp5_ASAP7_75t_L g1261 ( 
.A1(n_1122),
.A2(n_1163),
.B1(n_1116),
.B2(n_1123),
.Y(n_1261)
);

AOI22xp33_ASAP7_75t_L g1262 ( 
.A1(n_1094),
.A2(n_1124),
.B1(n_1106),
.B2(n_1115),
.Y(n_1262)
);

INVx1_ASAP7_75t_L g1263 ( 
.A(n_1135),
.Y(n_1263)
);

INVx1_ASAP7_75t_L g1264 ( 
.A(n_1135),
.Y(n_1264)
);

BUFx3_ASAP7_75t_L g1265 ( 
.A(n_1134),
.Y(n_1265)
);

CKINVDCx5p33_ASAP7_75t_R g1266 ( 
.A(n_1211),
.Y(n_1266)
);

INVx2_ASAP7_75t_SL g1267 ( 
.A(n_1144),
.Y(n_1267)
);

INVx4_ASAP7_75t_L g1268 ( 
.A(n_1156),
.Y(n_1268)
);

INVx1_ASAP7_75t_L g1269 ( 
.A(n_1211),
.Y(n_1269)
);

BUFx8_ASAP7_75t_SL g1270 ( 
.A(n_1136),
.Y(n_1270)
);

AOI22xp33_ASAP7_75t_L g1271 ( 
.A1(n_1118),
.A2(n_1166),
.B1(n_1139),
.B2(n_1159),
.Y(n_1271)
);

OAI22xp33_ASAP7_75t_L g1272 ( 
.A1(n_1133),
.A2(n_1121),
.B1(n_1113),
.B2(n_1169),
.Y(n_1272)
);

INVx5_ASAP7_75t_L g1273 ( 
.A(n_1211),
.Y(n_1273)
);

NAND2xp5_ASAP7_75t_L g1274 ( 
.A(n_1188),
.B(n_1178),
.Y(n_1274)
);

INVx4_ASAP7_75t_L g1275 ( 
.A(n_1156),
.Y(n_1275)
);

AOI22xp33_ASAP7_75t_L g1276 ( 
.A1(n_1118),
.A2(n_1152),
.B1(n_1173),
.B2(n_1183),
.Y(n_1276)
);

INVx1_ASAP7_75t_L g1277 ( 
.A(n_1117),
.Y(n_1277)
);

BUFx2_ASAP7_75t_L g1278 ( 
.A(n_1132),
.Y(n_1278)
);

BUFx6f_ASAP7_75t_SL g1279 ( 
.A(n_1204),
.Y(n_1279)
);

AOI22xp5_ASAP7_75t_L g1280 ( 
.A1(n_1167),
.A2(n_1181),
.B1(n_1188),
.B2(n_1081),
.Y(n_1280)
);

BUFx2_ASAP7_75t_L g1281 ( 
.A(n_1132),
.Y(n_1281)
);

INVx1_ASAP7_75t_L g1282 ( 
.A(n_1117),
.Y(n_1282)
);

INVx4_ASAP7_75t_L g1283 ( 
.A(n_1141),
.Y(n_1283)
);

BUFx2_ASAP7_75t_L g1284 ( 
.A(n_1117),
.Y(n_1284)
);

BUFx3_ASAP7_75t_L g1285 ( 
.A(n_1128),
.Y(n_1285)
);

BUFx12f_ASAP7_75t_L g1286 ( 
.A(n_1119),
.Y(n_1286)
);

OAI22xp33_ASAP7_75t_L g1287 ( 
.A1(n_1153),
.A2(n_1157),
.B1(n_1177),
.B2(n_1161),
.Y(n_1287)
);

HB1xp67_ASAP7_75t_L g1288 ( 
.A(n_1180),
.Y(n_1288)
);

OAI21xp5_ASAP7_75t_SL g1289 ( 
.A1(n_1129),
.A2(n_1131),
.B(n_1087),
.Y(n_1289)
);

INVx6_ASAP7_75t_L g1290 ( 
.A(n_1104),
.Y(n_1290)
);

BUFx12f_ASAP7_75t_L g1291 ( 
.A(n_1126),
.Y(n_1291)
);

AOI22xp33_ASAP7_75t_SL g1292 ( 
.A1(n_1187),
.A2(n_1161),
.B1(n_1177),
.B2(n_1157),
.Y(n_1292)
);

OAI22xp33_ASAP7_75t_L g1293 ( 
.A1(n_1153),
.A2(n_1161),
.B1(n_1177),
.B2(n_1157),
.Y(n_1293)
);

NAND2xp5_ASAP7_75t_L g1294 ( 
.A(n_1199),
.B(n_1209),
.Y(n_1294)
);

INVx1_ASAP7_75t_L g1295 ( 
.A(n_1199),
.Y(n_1295)
);

AOI22xp33_ASAP7_75t_L g1296 ( 
.A1(n_1130),
.A2(n_1153),
.B1(n_1108),
.B2(n_1089),
.Y(n_1296)
);

INVx1_ASAP7_75t_L g1297 ( 
.A(n_1209),
.Y(n_1297)
);

AOI22xp33_ASAP7_75t_L g1298 ( 
.A1(n_1145),
.A2(n_1155),
.B1(n_1162),
.B2(n_1179),
.Y(n_1298)
);

AOI22xp33_ASAP7_75t_SL g1299 ( 
.A1(n_1201),
.A2(n_1165),
.B1(n_1197),
.B2(n_1192),
.Y(n_1299)
);

INVx1_ASAP7_75t_L g1300 ( 
.A(n_1213),
.Y(n_1300)
);

NAND2xp5_ASAP7_75t_L g1301 ( 
.A(n_1165),
.B(n_1071),
.Y(n_1301)
);

BUFx8_ASAP7_75t_L g1302 ( 
.A(n_1172),
.Y(n_1302)
);

AOI22xp33_ASAP7_75t_L g1303 ( 
.A1(n_1165),
.A2(n_781),
.B1(n_1197),
.B2(n_1192),
.Y(n_1303)
);

INVx1_ASAP7_75t_L g1304 ( 
.A(n_1078),
.Y(n_1304)
);

INVx1_ASAP7_75t_SL g1305 ( 
.A(n_1143),
.Y(n_1305)
);

OAI22xp5_ASAP7_75t_L g1306 ( 
.A1(n_1165),
.A2(n_781),
.B1(n_1197),
.B2(n_1192),
.Y(n_1306)
);

NAND2xp5_ASAP7_75t_L g1307 ( 
.A(n_1165),
.B(n_1071),
.Y(n_1307)
);

INVx6_ASAP7_75t_L g1308 ( 
.A(n_1080),
.Y(n_1308)
);

CKINVDCx20_ASAP7_75t_R g1309 ( 
.A(n_1208),
.Y(n_1309)
);

OAI22xp33_ASAP7_75t_L g1310 ( 
.A1(n_1100),
.A2(n_954),
.B1(n_1192),
.B2(n_1165),
.Y(n_1310)
);

INVx6_ASAP7_75t_L g1311 ( 
.A(n_1080),
.Y(n_1311)
);

INVx2_ASAP7_75t_SL g1312 ( 
.A(n_1080),
.Y(n_1312)
);

INVx4_ASAP7_75t_L g1313 ( 
.A(n_1200),
.Y(n_1313)
);

AOI22xp33_ASAP7_75t_SL g1314 ( 
.A1(n_1165),
.A2(n_1192),
.B1(n_1197),
.B2(n_781),
.Y(n_1314)
);

CKINVDCx11_ASAP7_75t_R g1315 ( 
.A(n_1208),
.Y(n_1315)
);

INVx4_ASAP7_75t_L g1316 ( 
.A(n_1200),
.Y(n_1316)
);

BUFx2_ASAP7_75t_L g1317 ( 
.A(n_1083),
.Y(n_1317)
);

INVx6_ASAP7_75t_L g1318 ( 
.A(n_1080),
.Y(n_1318)
);

AND2x2_ASAP7_75t_L g1319 ( 
.A(n_1146),
.B(n_1147),
.Y(n_1319)
);

AOI22xp33_ASAP7_75t_L g1320 ( 
.A1(n_1165),
.A2(n_781),
.B1(n_1197),
.B2(n_1192),
.Y(n_1320)
);

AOI22xp33_ASAP7_75t_L g1321 ( 
.A1(n_1165),
.A2(n_781),
.B1(n_1197),
.B2(n_1192),
.Y(n_1321)
);

BUFx8_ASAP7_75t_L g1322 ( 
.A(n_1172),
.Y(n_1322)
);

OAI22xp5_ASAP7_75t_L g1323 ( 
.A1(n_1165),
.A2(n_781),
.B1(n_1197),
.B2(n_1192),
.Y(n_1323)
);

INVx6_ASAP7_75t_L g1324 ( 
.A(n_1080),
.Y(n_1324)
);

NAND2x1p5_ASAP7_75t_L g1325 ( 
.A(n_1144),
.B(n_847),
.Y(n_1325)
);

NAND2xp5_ASAP7_75t_L g1326 ( 
.A(n_1228),
.B(n_1217),
.Y(n_1326)
);

OR2x2_ASAP7_75t_L g1327 ( 
.A(n_1294),
.B(n_1295),
.Y(n_1327)
);

INVx1_ASAP7_75t_L g1328 ( 
.A(n_1297),
.Y(n_1328)
);

INVx1_ASAP7_75t_L g1329 ( 
.A(n_1288),
.Y(n_1329)
);

INVx3_ASAP7_75t_L g1330 ( 
.A(n_1285),
.Y(n_1330)
);

BUFx3_ASAP7_75t_L g1331 ( 
.A(n_1273),
.Y(n_1331)
);

AO21x2_ASAP7_75t_L g1332 ( 
.A1(n_1272),
.A2(n_1293),
.B(n_1287),
.Y(n_1332)
);

HB1xp67_ASAP7_75t_L g1333 ( 
.A(n_1230),
.Y(n_1333)
);

INVx1_ASAP7_75t_SL g1334 ( 
.A(n_1226),
.Y(n_1334)
);

INVx1_ASAP7_75t_L g1335 ( 
.A(n_1288),
.Y(n_1335)
);

AND2x2_ASAP7_75t_L g1336 ( 
.A(n_1229),
.B(n_1234),
.Y(n_1336)
);

INVx1_ASAP7_75t_L g1337 ( 
.A(n_1227),
.Y(n_1337)
);

INVx1_ASAP7_75t_L g1338 ( 
.A(n_1227),
.Y(n_1338)
);

INVx1_ASAP7_75t_L g1339 ( 
.A(n_1277),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_1282),
.Y(n_1340)
);

INVx1_ASAP7_75t_L g1341 ( 
.A(n_1263),
.Y(n_1341)
);

AND2x2_ASAP7_75t_L g1342 ( 
.A(n_1229),
.B(n_1234),
.Y(n_1342)
);

INVx1_ASAP7_75t_L g1343 ( 
.A(n_1264),
.Y(n_1343)
);

AND2x2_ASAP7_75t_L g1344 ( 
.A(n_1232),
.B(n_1244),
.Y(n_1344)
);

HB1xp67_ASAP7_75t_L g1345 ( 
.A(n_1230),
.Y(n_1345)
);

BUFx2_ASAP7_75t_L g1346 ( 
.A(n_1278),
.Y(n_1346)
);

AND2x4_ASAP7_75t_L g1347 ( 
.A(n_1265),
.B(n_1273),
.Y(n_1347)
);

AOI22xp33_ASAP7_75t_L g1348 ( 
.A1(n_1232),
.A2(n_1310),
.B1(n_1314),
.B2(n_1217),
.Y(n_1348)
);

INVx1_ASAP7_75t_L g1349 ( 
.A(n_1284),
.Y(n_1349)
);

INVx2_ASAP7_75t_L g1350 ( 
.A(n_1283),
.Y(n_1350)
);

INVxp33_ASAP7_75t_L g1351 ( 
.A(n_1237),
.Y(n_1351)
);

INVx2_ASAP7_75t_L g1352 ( 
.A(n_1300),
.Y(n_1352)
);

INVxp33_ASAP7_75t_L g1353 ( 
.A(n_1319),
.Y(n_1353)
);

INVx1_ASAP7_75t_L g1354 ( 
.A(n_1238),
.Y(n_1354)
);

INVx4_ASAP7_75t_SL g1355 ( 
.A(n_1290),
.Y(n_1355)
);

CKINVDCx6p67_ASAP7_75t_R g1356 ( 
.A(n_1248),
.Y(n_1356)
);

INVx2_ASAP7_75t_L g1357 ( 
.A(n_1240),
.Y(n_1357)
);

INVx1_ASAP7_75t_L g1358 ( 
.A(n_1274),
.Y(n_1358)
);

BUFx2_ASAP7_75t_L g1359 ( 
.A(n_1281),
.Y(n_1359)
);

NAND2xp5_ASAP7_75t_L g1360 ( 
.A(n_1233),
.B(n_1314),
.Y(n_1360)
);

INVx1_ASAP7_75t_L g1361 ( 
.A(n_1280),
.Y(n_1361)
);

INVx2_ASAP7_75t_SL g1362 ( 
.A(n_1214),
.Y(n_1362)
);

INVx1_ASAP7_75t_L g1363 ( 
.A(n_1292),
.Y(n_1363)
);

INVx1_ASAP7_75t_L g1364 ( 
.A(n_1293),
.Y(n_1364)
);

INVx1_ASAP7_75t_L g1365 ( 
.A(n_1304),
.Y(n_1365)
);

BUFx3_ASAP7_75t_L g1366 ( 
.A(n_1273),
.Y(n_1366)
);

OAI21xp33_ASAP7_75t_SL g1367 ( 
.A1(n_1262),
.A2(n_1253),
.B(n_1255),
.Y(n_1367)
);

AOI21xp5_ASAP7_75t_L g1368 ( 
.A1(n_1272),
.A2(n_1262),
.B(n_1289),
.Y(n_1368)
);

OAI21xp5_ASAP7_75t_L g1369 ( 
.A1(n_1306),
.A2(n_1323),
.B(n_1310),
.Y(n_1369)
);

NAND2x1p5_ASAP7_75t_L g1370 ( 
.A(n_1273),
.B(n_1269),
.Y(n_1370)
);

INVx1_ASAP7_75t_L g1371 ( 
.A(n_1255),
.Y(n_1371)
);

INVx1_ASAP7_75t_L g1372 ( 
.A(n_1253),
.Y(n_1372)
);

INVx2_ASAP7_75t_SL g1373 ( 
.A(n_1214),
.Y(n_1373)
);

AND2x2_ASAP7_75t_L g1374 ( 
.A(n_1244),
.B(n_1299),
.Y(n_1374)
);

AND2x2_ASAP7_75t_L g1375 ( 
.A(n_1299),
.B(n_1233),
.Y(n_1375)
);

HB1xp67_ASAP7_75t_L g1376 ( 
.A(n_1305),
.Y(n_1376)
);

OA21x2_ASAP7_75t_L g1377 ( 
.A1(n_1296),
.A2(n_1271),
.B(n_1276),
.Y(n_1377)
);

BUFx2_ASAP7_75t_L g1378 ( 
.A(n_1291),
.Y(n_1378)
);

BUFx6f_ASAP7_75t_L g1379 ( 
.A(n_1286),
.Y(n_1379)
);

NAND2xp5_ASAP7_75t_L g1380 ( 
.A(n_1303),
.B(n_1320),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_1250),
.Y(n_1381)
);

AND2x2_ASAP7_75t_L g1382 ( 
.A(n_1219),
.B(n_1235),
.Y(n_1382)
);

AOI21xp5_ASAP7_75t_L g1383 ( 
.A1(n_1271),
.A2(n_1276),
.B(n_1223),
.Y(n_1383)
);

INVx2_ASAP7_75t_SL g1384 ( 
.A(n_1214),
.Y(n_1384)
);

OAI21x1_ASAP7_75t_L g1385 ( 
.A1(n_1298),
.A2(n_1296),
.B(n_1219),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_1261),
.Y(n_1386)
);

INVx1_ASAP7_75t_L g1387 ( 
.A(n_1225),
.Y(n_1387)
);

INVx1_ASAP7_75t_L g1388 ( 
.A(n_1225),
.Y(n_1388)
);

INVx1_ASAP7_75t_SL g1389 ( 
.A(n_1317),
.Y(n_1389)
);

INVx1_ASAP7_75t_L g1390 ( 
.A(n_1249),
.Y(n_1390)
);

AOI22xp5_ASAP7_75t_L g1391 ( 
.A1(n_1303),
.A2(n_1320),
.B1(n_1321),
.B2(n_1307),
.Y(n_1391)
);

INVx1_ASAP7_75t_L g1392 ( 
.A(n_1251),
.Y(n_1392)
);

AND2x2_ASAP7_75t_L g1393 ( 
.A(n_1254),
.B(n_1257),
.Y(n_1393)
);

INVx1_ASAP7_75t_L g1394 ( 
.A(n_1267),
.Y(n_1394)
);

NAND2x1_ASAP7_75t_L g1395 ( 
.A(n_1268),
.B(n_1275),
.Y(n_1395)
);

INVxp33_ASAP7_75t_L g1396 ( 
.A(n_1258),
.Y(n_1396)
);

OAI21x1_ASAP7_75t_L g1397 ( 
.A1(n_1325),
.A2(n_1222),
.B(n_1321),
.Y(n_1397)
);

INVxp67_ASAP7_75t_L g1398 ( 
.A(n_1252),
.Y(n_1398)
);

AOI22xp33_ASAP7_75t_L g1399 ( 
.A1(n_1301),
.A2(n_1241),
.B1(n_1256),
.B2(n_1245),
.Y(n_1399)
);

OAI21x1_ASAP7_75t_L g1400 ( 
.A1(n_1270),
.A2(n_1266),
.B(n_1220),
.Y(n_1400)
);

OAI21x1_ASAP7_75t_L g1401 ( 
.A1(n_1220),
.A2(n_1231),
.B(n_1242),
.Y(n_1401)
);

NOR2xp33_ASAP7_75t_L g1402 ( 
.A(n_1351),
.B(n_1353),
.Y(n_1402)
);

A2O1A1Ixp33_ASAP7_75t_L g1403 ( 
.A1(n_1369),
.A2(n_1312),
.B(n_1218),
.C(n_1309),
.Y(n_1403)
);

INVx3_ASAP7_75t_L g1404 ( 
.A(n_1347),
.Y(n_1404)
);

OR2x6_ASAP7_75t_L g1405 ( 
.A(n_1383),
.B(n_1236),
.Y(n_1405)
);

INVx1_ASAP7_75t_L g1406 ( 
.A(n_1328),
.Y(n_1406)
);

OA21x2_ASAP7_75t_L g1407 ( 
.A1(n_1385),
.A2(n_1231),
.B(n_1313),
.Y(n_1407)
);

OAI21xp5_ASAP7_75t_L g1408 ( 
.A1(n_1348),
.A2(n_1236),
.B(n_1316),
.Y(n_1408)
);

OA21x2_ASAP7_75t_L g1409 ( 
.A1(n_1368),
.A2(n_1313),
.B(n_1239),
.Y(n_1409)
);

A2O1A1Ixp33_ASAP7_75t_L g1410 ( 
.A1(n_1367),
.A2(n_1241),
.B(n_1245),
.C(n_1246),
.Y(n_1410)
);

AOI221xp5_ASAP7_75t_L g1411 ( 
.A1(n_1326),
.A2(n_1279),
.B1(n_1259),
.B2(n_1247),
.C(n_1216),
.Y(n_1411)
);

A2O1A1Ixp33_ASAP7_75t_L g1412 ( 
.A1(n_1367),
.A2(n_1224),
.B(n_1243),
.C(n_1279),
.Y(n_1412)
);

INVxp67_ASAP7_75t_L g1413 ( 
.A(n_1376),
.Y(n_1413)
);

BUFx2_ASAP7_75t_SL g1414 ( 
.A(n_1379),
.Y(n_1414)
);

INVxp33_ASAP7_75t_L g1415 ( 
.A(n_1393),
.Y(n_1415)
);

OAI22xp5_ASAP7_75t_SL g1416 ( 
.A1(n_1391),
.A2(n_1215),
.B1(n_1318),
.B2(n_1311),
.Y(n_1416)
);

INVxp67_ASAP7_75t_L g1417 ( 
.A(n_1333),
.Y(n_1417)
);

HB1xp67_ASAP7_75t_L g1418 ( 
.A(n_1346),
.Y(n_1418)
);

AND2x2_ASAP7_75t_L g1419 ( 
.A(n_1363),
.B(n_1221),
.Y(n_1419)
);

OAI21xp5_ASAP7_75t_L g1420 ( 
.A1(n_1391),
.A2(n_1247),
.B(n_1259),
.Y(n_1420)
);

AND2x6_ASAP7_75t_L g1421 ( 
.A(n_1331),
.B(n_1260),
.Y(n_1421)
);

AND2x2_ASAP7_75t_L g1422 ( 
.A(n_1363),
.B(n_1215),
.Y(n_1422)
);

AO22x2_ASAP7_75t_L g1423 ( 
.A1(n_1336),
.A2(n_1224),
.B1(n_1315),
.B2(n_1311),
.Y(n_1423)
);

OAI21xp5_ASAP7_75t_L g1424 ( 
.A1(n_1360),
.A2(n_1315),
.B(n_1311),
.Y(n_1424)
);

O2A1O1Ixp33_ASAP7_75t_L g1425 ( 
.A1(n_1380),
.A2(n_1215),
.B(n_1308),
.C(n_1318),
.Y(n_1425)
);

OA21x2_ASAP7_75t_L g1426 ( 
.A1(n_1329),
.A2(n_1308),
.B(n_1318),
.Y(n_1426)
);

O2A1O1Ixp33_ASAP7_75t_L g1427 ( 
.A1(n_1386),
.A2(n_1324),
.B(n_1260),
.C(n_1322),
.Y(n_1427)
);

BUFx2_ASAP7_75t_L g1428 ( 
.A(n_1359),
.Y(n_1428)
);

AOI22xp5_ASAP7_75t_L g1429 ( 
.A1(n_1382),
.A2(n_1302),
.B1(n_1322),
.B2(n_1336),
.Y(n_1429)
);

OAI21xp5_ASAP7_75t_L g1430 ( 
.A1(n_1382),
.A2(n_1397),
.B(n_1342),
.Y(n_1430)
);

OA21x2_ASAP7_75t_L g1431 ( 
.A1(n_1329),
.A2(n_1335),
.B(n_1375),
.Y(n_1431)
);

AND2x4_ASAP7_75t_L g1432 ( 
.A(n_1330),
.B(n_1355),
.Y(n_1432)
);

AND2x2_ASAP7_75t_L g1433 ( 
.A(n_1364),
.B(n_1341),
.Y(n_1433)
);

AOI221xp5_ASAP7_75t_L g1434 ( 
.A1(n_1342),
.A2(n_1375),
.B1(n_1374),
.B2(n_1344),
.C(n_1390),
.Y(n_1434)
);

AND2x2_ASAP7_75t_L g1435 ( 
.A(n_1341),
.B(n_1343),
.Y(n_1435)
);

BUFx3_ASAP7_75t_L g1436 ( 
.A(n_1401),
.Y(n_1436)
);

NOR2xp33_ASAP7_75t_L g1437 ( 
.A(n_1396),
.B(n_1398),
.Y(n_1437)
);

AND2x2_ASAP7_75t_L g1438 ( 
.A(n_1343),
.B(n_1374),
.Y(n_1438)
);

AND2x2_ASAP7_75t_L g1439 ( 
.A(n_1357),
.B(n_1332),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_1357),
.Y(n_1440)
);

A2O1A1Ixp33_ASAP7_75t_L g1441 ( 
.A1(n_1344),
.A2(n_1387),
.B(n_1388),
.C(n_1371),
.Y(n_1441)
);

INVx1_ASAP7_75t_L g1442 ( 
.A(n_1352),
.Y(n_1442)
);

OAI22xp5_ASAP7_75t_L g1443 ( 
.A1(n_1399),
.A2(n_1372),
.B1(n_1371),
.B2(n_1389),
.Y(n_1443)
);

AOI211xp5_ASAP7_75t_L g1444 ( 
.A1(n_1387),
.A2(n_1388),
.B(n_1378),
.C(n_1372),
.Y(n_1444)
);

OAI21xp5_ASAP7_75t_L g1445 ( 
.A1(n_1397),
.A2(n_1361),
.B(n_1381),
.Y(n_1445)
);

AO32x2_ASAP7_75t_L g1446 ( 
.A1(n_1332),
.A2(n_1349),
.A3(n_1327),
.B1(n_1378),
.B2(n_1340),
.Y(n_1446)
);

HB1xp67_ASAP7_75t_L g1447 ( 
.A(n_1345),
.Y(n_1447)
);

AND2x2_ASAP7_75t_L g1448 ( 
.A(n_1332),
.B(n_1354),
.Y(n_1448)
);

AND2x2_ASAP7_75t_L g1449 ( 
.A(n_1438),
.B(n_1439),
.Y(n_1449)
);

AND2x2_ASAP7_75t_L g1450 ( 
.A(n_1438),
.B(n_1350),
.Y(n_1450)
);

AND2x4_ASAP7_75t_SL g1451 ( 
.A(n_1432),
.B(n_1347),
.Y(n_1451)
);

NAND2xp5_ASAP7_75t_L g1452 ( 
.A(n_1448),
.B(n_1337),
.Y(n_1452)
);

BUFx3_ASAP7_75t_L g1453 ( 
.A(n_1426),
.Y(n_1453)
);

INVx1_ASAP7_75t_L g1454 ( 
.A(n_1406),
.Y(n_1454)
);

NAND2xp5_ASAP7_75t_L g1455 ( 
.A(n_1448),
.B(n_1338),
.Y(n_1455)
);

AOI22xp33_ASAP7_75t_SL g1456 ( 
.A1(n_1416),
.A2(n_1332),
.B1(n_1366),
.B2(n_1400),
.Y(n_1456)
);

OR2x2_ASAP7_75t_L g1457 ( 
.A(n_1439),
.B(n_1338),
.Y(n_1457)
);

AND2x2_ASAP7_75t_L g1458 ( 
.A(n_1430),
.B(n_1350),
.Y(n_1458)
);

CKINVDCx6p67_ASAP7_75t_R g1459 ( 
.A(n_1421),
.Y(n_1459)
);

AND2x2_ASAP7_75t_SL g1460 ( 
.A(n_1409),
.B(n_1377),
.Y(n_1460)
);

INVx1_ASAP7_75t_L g1461 ( 
.A(n_1440),
.Y(n_1461)
);

INVx1_ASAP7_75t_L g1462 ( 
.A(n_1440),
.Y(n_1462)
);

OR2x2_ASAP7_75t_L g1463 ( 
.A(n_1418),
.B(n_1327),
.Y(n_1463)
);

INVx2_ASAP7_75t_L g1464 ( 
.A(n_1442),
.Y(n_1464)
);

BUFx6f_ASAP7_75t_L g1465 ( 
.A(n_1407),
.Y(n_1465)
);

AND2x2_ASAP7_75t_L g1466 ( 
.A(n_1415),
.B(n_1433),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_1442),
.Y(n_1467)
);

HB1xp67_ASAP7_75t_L g1468 ( 
.A(n_1428),
.Y(n_1468)
);

BUFx3_ASAP7_75t_L g1469 ( 
.A(n_1426),
.Y(n_1469)
);

OR2x2_ASAP7_75t_L g1470 ( 
.A(n_1428),
.B(n_1340),
.Y(n_1470)
);

AND2x2_ASAP7_75t_L g1471 ( 
.A(n_1435),
.B(n_1339),
.Y(n_1471)
);

OAI222xp33_ASAP7_75t_L g1472 ( 
.A1(n_1429),
.A2(n_1392),
.B1(n_1389),
.B2(n_1358),
.C1(n_1334),
.C2(n_1370),
.Y(n_1472)
);

NAND2xp5_ASAP7_75t_L g1473 ( 
.A(n_1447),
.B(n_1445),
.Y(n_1473)
);

NOR2xp33_ASAP7_75t_SL g1474 ( 
.A(n_1472),
.B(n_1412),
.Y(n_1474)
);

OR2x2_ASAP7_75t_L g1475 ( 
.A(n_1452),
.B(n_1431),
.Y(n_1475)
);

INVx2_ASAP7_75t_L g1476 ( 
.A(n_1464),
.Y(n_1476)
);

NAND2xp5_ASAP7_75t_L g1477 ( 
.A(n_1452),
.B(n_1431),
.Y(n_1477)
);

INVx3_ASAP7_75t_L g1478 ( 
.A(n_1465),
.Y(n_1478)
);

NAND3xp33_ASAP7_75t_L g1479 ( 
.A(n_1456),
.B(n_1444),
.C(n_1410),
.Y(n_1479)
);

AND2x2_ASAP7_75t_L g1480 ( 
.A(n_1460),
.B(n_1431),
.Y(n_1480)
);

AND2x2_ASAP7_75t_L g1481 ( 
.A(n_1460),
.B(n_1431),
.Y(n_1481)
);

AND2x2_ASAP7_75t_L g1482 ( 
.A(n_1460),
.B(n_1446),
.Y(n_1482)
);

OAI31xp33_ASAP7_75t_L g1483 ( 
.A1(n_1472),
.A2(n_1423),
.A3(n_1403),
.B(n_1441),
.Y(n_1483)
);

AND2x2_ASAP7_75t_L g1484 ( 
.A(n_1449),
.B(n_1446),
.Y(n_1484)
);

INVx1_ASAP7_75t_L g1485 ( 
.A(n_1461),
.Y(n_1485)
);

INVx1_ASAP7_75t_L g1486 ( 
.A(n_1461),
.Y(n_1486)
);

BUFx2_ASAP7_75t_L g1487 ( 
.A(n_1453),
.Y(n_1487)
);

AND2x2_ASAP7_75t_L g1488 ( 
.A(n_1449),
.B(n_1446),
.Y(n_1488)
);

INVx1_ASAP7_75t_SL g1489 ( 
.A(n_1457),
.Y(n_1489)
);

INVx1_ASAP7_75t_L g1490 ( 
.A(n_1462),
.Y(n_1490)
);

INVx1_ASAP7_75t_L g1491 ( 
.A(n_1462),
.Y(n_1491)
);

OAI21xp33_ASAP7_75t_L g1492 ( 
.A1(n_1473),
.A2(n_1434),
.B(n_1423),
.Y(n_1492)
);

INVx1_ASAP7_75t_L g1493 ( 
.A(n_1467),
.Y(n_1493)
);

NOR2xp33_ASAP7_75t_SL g1494 ( 
.A(n_1459),
.B(n_1414),
.Y(n_1494)
);

NOR2xp67_ASAP7_75t_L g1495 ( 
.A(n_1453),
.B(n_1404),
.Y(n_1495)
);

INVxp67_ASAP7_75t_SL g1496 ( 
.A(n_1455),
.Y(n_1496)
);

AND2x2_ASAP7_75t_L g1497 ( 
.A(n_1465),
.B(n_1446),
.Y(n_1497)
);

NOR2xp33_ASAP7_75t_R g1498 ( 
.A(n_1459),
.B(n_1356),
.Y(n_1498)
);

OAI33xp33_ASAP7_75t_L g1499 ( 
.A1(n_1473),
.A2(n_1443),
.A3(n_1417),
.B1(n_1413),
.B2(n_1394),
.B3(n_1365),
.Y(n_1499)
);

AND2x2_ASAP7_75t_SL g1500 ( 
.A(n_1465),
.B(n_1377),
.Y(n_1500)
);

AND2x2_ASAP7_75t_L g1501 ( 
.A(n_1465),
.B(n_1446),
.Y(n_1501)
);

INVxp67_ASAP7_75t_SL g1502 ( 
.A(n_1455),
.Y(n_1502)
);

HB1xp67_ASAP7_75t_L g1503 ( 
.A(n_1457),
.Y(n_1503)
);

INVx2_ASAP7_75t_L g1504 ( 
.A(n_1465),
.Y(n_1504)
);

AND2x2_ASAP7_75t_L g1505 ( 
.A(n_1453),
.B(n_1377),
.Y(n_1505)
);

NOR2xp33_ASAP7_75t_L g1506 ( 
.A(n_1458),
.B(n_1419),
.Y(n_1506)
);

AND2x2_ASAP7_75t_L g1507 ( 
.A(n_1480),
.B(n_1469),
.Y(n_1507)
);

AND2x2_ASAP7_75t_L g1508 ( 
.A(n_1480),
.B(n_1469),
.Y(n_1508)
);

OR2x2_ASAP7_75t_L g1509 ( 
.A(n_1496),
.B(n_1463),
.Y(n_1509)
);

AND2x2_ASAP7_75t_L g1510 ( 
.A(n_1480),
.B(n_1469),
.Y(n_1510)
);

NAND2xp5_ASAP7_75t_L g1511 ( 
.A(n_1496),
.B(n_1502),
.Y(n_1511)
);

OR2x2_ASAP7_75t_L g1512 ( 
.A(n_1502),
.B(n_1463),
.Y(n_1512)
);

AND2x4_ASAP7_75t_L g1513 ( 
.A(n_1495),
.B(n_1451),
.Y(n_1513)
);

INVx1_ASAP7_75t_L g1514 ( 
.A(n_1485),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_1485),
.Y(n_1515)
);

AND2x4_ASAP7_75t_L g1516 ( 
.A(n_1495),
.B(n_1451),
.Y(n_1516)
);

HB1xp67_ASAP7_75t_L g1517 ( 
.A(n_1485),
.Y(n_1517)
);

NAND2xp5_ASAP7_75t_L g1518 ( 
.A(n_1477),
.B(n_1468),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_1486),
.Y(n_1519)
);

INVx1_ASAP7_75t_L g1520 ( 
.A(n_1486),
.Y(n_1520)
);

BUFx3_ASAP7_75t_L g1521 ( 
.A(n_1487),
.Y(n_1521)
);

NOR2x1p5_ASAP7_75t_L g1522 ( 
.A(n_1479),
.B(n_1459),
.Y(n_1522)
);

HB1xp67_ASAP7_75t_L g1523 ( 
.A(n_1486),
.Y(n_1523)
);

OR2x2_ASAP7_75t_L g1524 ( 
.A(n_1489),
.B(n_1470),
.Y(n_1524)
);

INVx2_ASAP7_75t_L g1525 ( 
.A(n_1476),
.Y(n_1525)
);

HB1xp67_ASAP7_75t_L g1526 ( 
.A(n_1490),
.Y(n_1526)
);

INVx1_ASAP7_75t_L g1527 ( 
.A(n_1490),
.Y(n_1527)
);

NAND2xp5_ASAP7_75t_L g1528 ( 
.A(n_1477),
.B(n_1471),
.Y(n_1528)
);

HB1xp67_ASAP7_75t_L g1529 ( 
.A(n_1490),
.Y(n_1529)
);

INVx1_ASAP7_75t_L g1530 ( 
.A(n_1491),
.Y(n_1530)
);

AND3x1_ASAP7_75t_L g1531 ( 
.A(n_1483),
.B(n_1411),
.C(n_1427),
.Y(n_1531)
);

INVx1_ASAP7_75t_L g1532 ( 
.A(n_1491),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_1491),
.Y(n_1533)
);

NOR2x1_ASAP7_75t_L g1534 ( 
.A(n_1479),
.B(n_1436),
.Y(n_1534)
);

AND2x2_ASAP7_75t_L g1535 ( 
.A(n_1484),
.B(n_1458),
.Y(n_1535)
);

OR2x2_ASAP7_75t_L g1536 ( 
.A(n_1489),
.B(n_1503),
.Y(n_1536)
);

INVxp67_ASAP7_75t_SL g1537 ( 
.A(n_1476),
.Y(n_1537)
);

AND2x2_ASAP7_75t_L g1538 ( 
.A(n_1480),
.B(n_1450),
.Y(n_1538)
);

AND2x2_ASAP7_75t_L g1539 ( 
.A(n_1481),
.B(n_1450),
.Y(n_1539)
);

BUFx2_ASAP7_75t_L g1540 ( 
.A(n_1498),
.Y(n_1540)
);

AND2x2_ASAP7_75t_L g1541 ( 
.A(n_1484),
.B(n_1466),
.Y(n_1541)
);

NOR2xp67_ASAP7_75t_L g1542 ( 
.A(n_1481),
.B(n_1454),
.Y(n_1542)
);

INVx1_ASAP7_75t_L g1543 ( 
.A(n_1493),
.Y(n_1543)
);

INVx1_ASAP7_75t_L g1544 ( 
.A(n_1517),
.Y(n_1544)
);

INVx1_ASAP7_75t_L g1545 ( 
.A(n_1517),
.Y(n_1545)
);

INVx1_ASAP7_75t_L g1546 ( 
.A(n_1523),
.Y(n_1546)
);

OR2x2_ASAP7_75t_L g1547 ( 
.A(n_1528),
.B(n_1492),
.Y(n_1547)
);

INVx1_ASAP7_75t_L g1548 ( 
.A(n_1523),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_1526),
.Y(n_1549)
);

NAND2xp5_ASAP7_75t_SL g1550 ( 
.A(n_1534),
.B(n_1483),
.Y(n_1550)
);

NAND2xp5_ASAP7_75t_L g1551 ( 
.A(n_1534),
.B(n_1492),
.Y(n_1551)
);

NAND2xp5_ASAP7_75t_L g1552 ( 
.A(n_1522),
.B(n_1492),
.Y(n_1552)
);

INVx1_ASAP7_75t_L g1553 ( 
.A(n_1526),
.Y(n_1553)
);

INVxp33_ASAP7_75t_L g1554 ( 
.A(n_1540),
.Y(n_1554)
);

NAND2x2_ASAP7_75t_L g1555 ( 
.A(n_1522),
.B(n_1362),
.Y(n_1555)
);

INVx1_ASAP7_75t_L g1556 ( 
.A(n_1529),
.Y(n_1556)
);

AND2x4_ASAP7_75t_L g1557 ( 
.A(n_1513),
.B(n_1495),
.Y(n_1557)
);

NAND4xp25_ASAP7_75t_L g1558 ( 
.A(n_1540),
.B(n_1483),
.C(n_1479),
.D(n_1474),
.Y(n_1558)
);

OR2x2_ASAP7_75t_L g1559 ( 
.A(n_1528),
.B(n_1506),
.Y(n_1559)
);

INVx1_ASAP7_75t_L g1560 ( 
.A(n_1529),
.Y(n_1560)
);

INVx1_ASAP7_75t_L g1561 ( 
.A(n_1514),
.Y(n_1561)
);

AND2x2_ASAP7_75t_L g1562 ( 
.A(n_1513),
.B(n_1484),
.Y(n_1562)
);

AND2x2_ASAP7_75t_L g1563 ( 
.A(n_1513),
.B(n_1484),
.Y(n_1563)
);

INVx1_ASAP7_75t_L g1564 ( 
.A(n_1514),
.Y(n_1564)
);

NAND2xp5_ASAP7_75t_L g1565 ( 
.A(n_1518),
.B(n_1506),
.Y(n_1565)
);

INVx1_ASAP7_75t_L g1566 ( 
.A(n_1515),
.Y(n_1566)
);

INVx2_ASAP7_75t_L g1567 ( 
.A(n_1521),
.Y(n_1567)
);

NAND2xp5_ASAP7_75t_L g1568 ( 
.A(n_1518),
.B(n_1481),
.Y(n_1568)
);

INVxp67_ASAP7_75t_SL g1569 ( 
.A(n_1521),
.Y(n_1569)
);

NOR2x1_ASAP7_75t_L g1570 ( 
.A(n_1521),
.B(n_1487),
.Y(n_1570)
);

INVxp67_ASAP7_75t_L g1571 ( 
.A(n_1531),
.Y(n_1571)
);

OR2x2_ASAP7_75t_L g1572 ( 
.A(n_1509),
.B(n_1503),
.Y(n_1572)
);

NAND2xp5_ASAP7_75t_L g1573 ( 
.A(n_1509),
.B(n_1481),
.Y(n_1573)
);

INVx1_ASAP7_75t_L g1574 ( 
.A(n_1515),
.Y(n_1574)
);

OAI31xp33_ASAP7_75t_L g1575 ( 
.A1(n_1531),
.A2(n_1474),
.A3(n_1423),
.B(n_1482),
.Y(n_1575)
);

INVx2_ASAP7_75t_SL g1576 ( 
.A(n_1513),
.Y(n_1576)
);

NAND2xp5_ASAP7_75t_L g1577 ( 
.A(n_1512),
.B(n_1422),
.Y(n_1577)
);

AND2x2_ASAP7_75t_L g1578 ( 
.A(n_1516),
.B(n_1488),
.Y(n_1578)
);

INVx1_ASAP7_75t_L g1579 ( 
.A(n_1519),
.Y(n_1579)
);

OR2x6_ASAP7_75t_L g1580 ( 
.A(n_1511),
.B(n_1423),
.Y(n_1580)
);

HB1xp67_ASAP7_75t_L g1581 ( 
.A(n_1519),
.Y(n_1581)
);

OR2x2_ASAP7_75t_L g1582 ( 
.A(n_1512),
.B(n_1466),
.Y(n_1582)
);

NAND3xp33_ASAP7_75t_SL g1583 ( 
.A(n_1511),
.B(n_1498),
.C(n_1482),
.Y(n_1583)
);

AND2x2_ASAP7_75t_L g1584 ( 
.A(n_1516),
.B(n_1488),
.Y(n_1584)
);

HB1xp67_ASAP7_75t_L g1585 ( 
.A(n_1520),
.Y(n_1585)
);

INVx2_ASAP7_75t_L g1586 ( 
.A(n_1581),
.Y(n_1586)
);

OR2x2_ASAP7_75t_L g1587 ( 
.A(n_1559),
.B(n_1536),
.Y(n_1587)
);

NAND2xp5_ASAP7_75t_L g1588 ( 
.A(n_1571),
.B(n_1535),
.Y(n_1588)
);

INVx1_ASAP7_75t_L g1589 ( 
.A(n_1581),
.Y(n_1589)
);

NAND4xp25_ASAP7_75t_L g1590 ( 
.A(n_1558),
.B(n_1424),
.C(n_1425),
.D(n_1420),
.Y(n_1590)
);

AND2x2_ASAP7_75t_L g1591 ( 
.A(n_1580),
.B(n_1516),
.Y(n_1591)
);

OR2x2_ASAP7_75t_L g1592 ( 
.A(n_1572),
.B(n_1536),
.Y(n_1592)
);

NAND2xp5_ASAP7_75t_L g1593 ( 
.A(n_1554),
.B(n_1535),
.Y(n_1593)
);

INVx2_ASAP7_75t_L g1594 ( 
.A(n_1585),
.Y(n_1594)
);

OAI22xp5_ASAP7_75t_L g1595 ( 
.A1(n_1550),
.A2(n_1500),
.B1(n_1482),
.B2(n_1405),
.Y(n_1595)
);

HB1xp67_ASAP7_75t_L g1596 ( 
.A(n_1570),
.Y(n_1596)
);

AND2x2_ASAP7_75t_L g1597 ( 
.A(n_1580),
.B(n_1516),
.Y(n_1597)
);

INVx1_ASAP7_75t_L g1598 ( 
.A(n_1585),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1561),
.Y(n_1599)
);

NOR2x2_ASAP7_75t_L g1600 ( 
.A(n_1580),
.B(n_1504),
.Y(n_1600)
);

OR2x2_ASAP7_75t_L g1601 ( 
.A(n_1582),
.B(n_1475),
.Y(n_1601)
);

NAND2xp5_ASAP7_75t_L g1602 ( 
.A(n_1554),
.B(n_1538),
.Y(n_1602)
);

NAND2xp5_ASAP7_75t_L g1603 ( 
.A(n_1552),
.B(n_1575),
.Y(n_1603)
);

NAND2xp5_ASAP7_75t_L g1604 ( 
.A(n_1551),
.B(n_1565),
.Y(n_1604)
);

INVx2_ASAP7_75t_L g1605 ( 
.A(n_1567),
.Y(n_1605)
);

INVx2_ASAP7_75t_L g1606 ( 
.A(n_1567),
.Y(n_1606)
);

AND2x2_ASAP7_75t_L g1607 ( 
.A(n_1580),
.B(n_1538),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_1564),
.Y(n_1608)
);

INVx2_ASAP7_75t_L g1609 ( 
.A(n_1566),
.Y(n_1609)
);

INVx1_ASAP7_75t_L g1610 ( 
.A(n_1574),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_1579),
.Y(n_1611)
);

AND2x2_ASAP7_75t_L g1612 ( 
.A(n_1576),
.B(n_1538),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1544),
.Y(n_1613)
);

NAND2xp5_ASAP7_75t_L g1614 ( 
.A(n_1550),
.B(n_1539),
.Y(n_1614)
);

INVxp67_ASAP7_75t_SL g1615 ( 
.A(n_1569),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_1545),
.Y(n_1616)
);

OR2x2_ASAP7_75t_L g1617 ( 
.A(n_1547),
.B(n_1475),
.Y(n_1617)
);

AND2x2_ASAP7_75t_L g1618 ( 
.A(n_1576),
.B(n_1539),
.Y(n_1618)
);

NAND2xp5_ASAP7_75t_SL g1619 ( 
.A(n_1557),
.B(n_1494),
.Y(n_1619)
);

INVx1_ASAP7_75t_SL g1620 ( 
.A(n_1546),
.Y(n_1620)
);

INVx1_ASAP7_75t_L g1621 ( 
.A(n_1586),
.Y(n_1621)
);

AOI22xp5_ASAP7_75t_L g1622 ( 
.A1(n_1603),
.A2(n_1583),
.B1(n_1555),
.B2(n_1499),
.Y(n_1622)
);

OAI22xp5_ASAP7_75t_L g1623 ( 
.A1(n_1614),
.A2(n_1555),
.B1(n_1482),
.B2(n_1500),
.Y(n_1623)
);

INVx1_ASAP7_75t_L g1624 ( 
.A(n_1586),
.Y(n_1624)
);

NAND2xp5_ASAP7_75t_L g1625 ( 
.A(n_1615),
.B(n_1548),
.Y(n_1625)
);

AOI221xp5_ASAP7_75t_L g1626 ( 
.A1(n_1595),
.A2(n_1499),
.B1(n_1568),
.B2(n_1573),
.C(n_1560),
.Y(n_1626)
);

INVx1_ASAP7_75t_L g1627 ( 
.A(n_1586),
.Y(n_1627)
);

AND2x2_ASAP7_75t_SL g1628 ( 
.A(n_1596),
.B(n_1494),
.Y(n_1628)
);

INVx1_ASAP7_75t_L g1629 ( 
.A(n_1594),
.Y(n_1629)
);

AOI21xp33_ASAP7_75t_L g1630 ( 
.A1(n_1620),
.A2(n_1553),
.B(n_1549),
.Y(n_1630)
);

OAI221xp5_ASAP7_75t_L g1631 ( 
.A1(n_1595),
.A2(n_1556),
.B1(n_1577),
.B2(n_1487),
.C(n_1542),
.Y(n_1631)
);

OR2x2_ASAP7_75t_L g1632 ( 
.A(n_1588),
.B(n_1524),
.Y(n_1632)
);

INVx1_ASAP7_75t_SL g1633 ( 
.A(n_1620),
.Y(n_1633)
);

AND2x2_ASAP7_75t_L g1634 ( 
.A(n_1591),
.B(n_1562),
.Y(n_1634)
);

NOR2x1_ASAP7_75t_L g1635 ( 
.A(n_1589),
.B(n_1598),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_1594),
.Y(n_1636)
);

INVx2_ASAP7_75t_SL g1637 ( 
.A(n_1612),
.Y(n_1637)
);

NOR2xp33_ASAP7_75t_L g1638 ( 
.A(n_1604),
.B(n_1356),
.Y(n_1638)
);

OR2x2_ASAP7_75t_L g1639 ( 
.A(n_1587),
.B(n_1593),
.Y(n_1639)
);

INVx2_ASAP7_75t_L g1640 ( 
.A(n_1612),
.Y(n_1640)
);

NOR2xp33_ASAP7_75t_L g1641 ( 
.A(n_1587),
.B(n_1362),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_1594),
.Y(n_1642)
);

AO21x1_ASAP7_75t_L g1643 ( 
.A1(n_1589),
.A2(n_1557),
.B(n_1508),
.Y(n_1643)
);

AOI322xp5_ASAP7_75t_L g1644 ( 
.A1(n_1607),
.A2(n_1497),
.A3(n_1501),
.B1(n_1510),
.B2(n_1507),
.C1(n_1508),
.C2(n_1584),
.Y(n_1644)
);

AOI221xp5_ASAP7_75t_L g1645 ( 
.A1(n_1613),
.A2(n_1616),
.B1(n_1602),
.B2(n_1590),
.C(n_1607),
.Y(n_1645)
);

NAND2xp5_ASAP7_75t_SL g1646 ( 
.A(n_1628),
.B(n_1592),
.Y(n_1646)
);

INVx2_ASAP7_75t_L g1647 ( 
.A(n_1634),
.Y(n_1647)
);

OAI21xp33_ASAP7_75t_L g1648 ( 
.A1(n_1622),
.A2(n_1619),
.B(n_1590),
.Y(n_1648)
);

AOI22xp5_ASAP7_75t_L g1649 ( 
.A1(n_1643),
.A2(n_1591),
.B1(n_1597),
.B2(n_1618),
.Y(n_1649)
);

AND2x2_ASAP7_75t_L g1650 ( 
.A(n_1637),
.B(n_1597),
.Y(n_1650)
);

OAI22xp5_ASAP7_75t_L g1651 ( 
.A1(n_1633),
.A2(n_1592),
.B1(n_1618),
.B2(n_1617),
.Y(n_1651)
);

OAI222xp33_ASAP7_75t_L g1652 ( 
.A1(n_1631),
.A2(n_1617),
.B1(n_1600),
.B2(n_1613),
.C1(n_1616),
.C2(n_1601),
.Y(n_1652)
);

AOI21xp33_ASAP7_75t_L g1653 ( 
.A1(n_1633),
.A2(n_1606),
.B(n_1605),
.Y(n_1653)
);

NAND2xp5_ASAP7_75t_L g1654 ( 
.A(n_1645),
.B(n_1605),
.Y(n_1654)
);

INVx1_ASAP7_75t_SL g1655 ( 
.A(n_1635),
.Y(n_1655)
);

AOI221xp5_ASAP7_75t_L g1656 ( 
.A1(n_1630),
.A2(n_1598),
.B1(n_1606),
.B2(n_1605),
.C(n_1608),
.Y(n_1656)
);

O2A1O1Ixp33_ASAP7_75t_L g1657 ( 
.A1(n_1630),
.A2(n_1606),
.B(n_1610),
.C(n_1599),
.Y(n_1657)
);

NOR2xp33_ASAP7_75t_L g1658 ( 
.A(n_1638),
.B(n_1599),
.Y(n_1658)
);

AOI22xp5_ASAP7_75t_L g1659 ( 
.A1(n_1640),
.A2(n_1557),
.B1(n_1500),
.B2(n_1608),
.Y(n_1659)
);

INVx1_ASAP7_75t_L g1660 ( 
.A(n_1621),
.Y(n_1660)
);

OR2x2_ASAP7_75t_L g1661 ( 
.A(n_1639),
.B(n_1601),
.Y(n_1661)
);

INVx1_ASAP7_75t_L g1662 ( 
.A(n_1624),
.Y(n_1662)
);

OAI22xp33_ASAP7_75t_L g1663 ( 
.A1(n_1623),
.A2(n_1542),
.B1(n_1475),
.B2(n_1524),
.Y(n_1663)
);

OAI22xp5_ASAP7_75t_L g1664 ( 
.A1(n_1632),
.A2(n_1578),
.B1(n_1562),
.B2(n_1563),
.Y(n_1664)
);

AND2x2_ASAP7_75t_L g1665 ( 
.A(n_1650),
.B(n_1625),
.Y(n_1665)
);

NAND2xp5_ASAP7_75t_L g1666 ( 
.A(n_1647),
.B(n_1641),
.Y(n_1666)
);

INVx2_ASAP7_75t_L g1667 ( 
.A(n_1655),
.Y(n_1667)
);

OAI222xp33_ASAP7_75t_L g1668 ( 
.A1(n_1655),
.A2(n_1623),
.B1(n_1625),
.B2(n_1636),
.C1(n_1627),
.C2(n_1629),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_1657),
.Y(n_1669)
);

INVx1_ASAP7_75t_L g1670 ( 
.A(n_1660),
.Y(n_1670)
);

INVxp67_ASAP7_75t_L g1671 ( 
.A(n_1646),
.Y(n_1671)
);

INVxp33_ASAP7_75t_L g1672 ( 
.A(n_1658),
.Y(n_1672)
);

INVx1_ASAP7_75t_L g1673 ( 
.A(n_1662),
.Y(n_1673)
);

AND2x4_ASAP7_75t_SL g1674 ( 
.A(n_1649),
.B(n_1642),
.Y(n_1674)
);

AND2x2_ASAP7_75t_L g1675 ( 
.A(n_1651),
.B(n_1563),
.Y(n_1675)
);

NOR2x1_ASAP7_75t_SL g1676 ( 
.A(n_1667),
.B(n_1661),
.Y(n_1676)
);

AOI211xp5_ASAP7_75t_L g1677 ( 
.A1(n_1668),
.A2(n_1648),
.B(n_1652),
.C(n_1654),
.Y(n_1677)
);

INVx1_ASAP7_75t_SL g1678 ( 
.A(n_1665),
.Y(n_1678)
);

OAI21xp33_ASAP7_75t_L g1679 ( 
.A1(n_1674),
.A2(n_1659),
.B(n_1644),
.Y(n_1679)
);

OAI21xp33_ASAP7_75t_L g1680 ( 
.A1(n_1674),
.A2(n_1664),
.B(n_1653),
.Y(n_1680)
);

NAND3xp33_ASAP7_75t_L g1681 ( 
.A(n_1669),
.B(n_1656),
.C(n_1626),
.Y(n_1681)
);

NOR2xp33_ASAP7_75t_L g1682 ( 
.A(n_1672),
.B(n_1663),
.Y(n_1682)
);

NOR2xp33_ASAP7_75t_L g1683 ( 
.A(n_1671),
.B(n_1610),
.Y(n_1683)
);

AOI21xp5_ASAP7_75t_L g1684 ( 
.A1(n_1669),
.A2(n_1667),
.B(n_1666),
.Y(n_1684)
);

OAI21xp5_ASAP7_75t_L g1685 ( 
.A1(n_1665),
.A2(n_1611),
.B(n_1609),
.Y(n_1685)
);

O2A1O1Ixp33_ASAP7_75t_L g1686 ( 
.A1(n_1677),
.A2(n_1673),
.B(n_1670),
.C(n_1675),
.Y(n_1686)
);

OAI22xp5_ASAP7_75t_L g1687 ( 
.A1(n_1681),
.A2(n_1675),
.B1(n_1673),
.B2(n_1670),
.Y(n_1687)
);

NAND2xp5_ASAP7_75t_L g1688 ( 
.A(n_1676),
.B(n_1611),
.Y(n_1688)
);

AOI221xp5_ASAP7_75t_L g1689 ( 
.A1(n_1679),
.A2(n_1609),
.B1(n_1507),
.B2(n_1510),
.C(n_1508),
.Y(n_1689)
);

OAI221xp5_ASAP7_75t_L g1690 ( 
.A1(n_1680),
.A2(n_1609),
.B1(n_1334),
.B2(n_1437),
.C(n_1584),
.Y(n_1690)
);

XNOR2x2_ASAP7_75t_L g1691 ( 
.A(n_1684),
.B(n_1497),
.Y(n_1691)
);

AOI21xp5_ASAP7_75t_L g1692 ( 
.A1(n_1682),
.A2(n_1537),
.B(n_1510),
.Y(n_1692)
);

OAI31xp33_ASAP7_75t_L g1693 ( 
.A1(n_1687),
.A2(n_1678),
.A3(n_1683),
.B(n_1685),
.Y(n_1693)
);

OA222x2_ASAP7_75t_L g1694 ( 
.A1(n_1688),
.A2(n_1478),
.B1(n_1504),
.B2(n_1475),
.C1(n_1405),
.C2(n_1436),
.Y(n_1694)
);

AOI22xp5_ASAP7_75t_L g1695 ( 
.A1(n_1689),
.A2(n_1690),
.B1(n_1692),
.B2(n_1578),
.Y(n_1695)
);

NOR3xp33_ASAP7_75t_L g1696 ( 
.A(n_1686),
.B(n_1384),
.C(n_1373),
.Y(n_1696)
);

OAI221xp5_ASAP7_75t_L g1697 ( 
.A1(n_1691),
.A2(n_1384),
.B1(n_1507),
.B2(n_1419),
.C(n_1379),
.Y(n_1697)
);

AOI221xp5_ASAP7_75t_L g1698 ( 
.A1(n_1686),
.A2(n_1497),
.B1(n_1501),
.B2(n_1504),
.C(n_1505),
.Y(n_1698)
);

OR2x2_ASAP7_75t_L g1699 ( 
.A(n_1693),
.B(n_1695),
.Y(n_1699)
);

NAND2x1p5_ASAP7_75t_L g1700 ( 
.A(n_1696),
.B(n_1379),
.Y(n_1700)
);

NOR2x1_ASAP7_75t_L g1701 ( 
.A(n_1697),
.B(n_1379),
.Y(n_1701)
);

AND2x4_ASAP7_75t_L g1702 ( 
.A(n_1694),
.B(n_1539),
.Y(n_1702)
);

AOI22xp5_ASAP7_75t_L g1703 ( 
.A1(n_1698),
.A2(n_1379),
.B1(n_1504),
.B2(n_1421),
.Y(n_1703)
);

INVxp67_ASAP7_75t_L g1704 ( 
.A(n_1702),
.Y(n_1704)
);

NAND2xp5_ASAP7_75t_SL g1705 ( 
.A(n_1701),
.B(n_1379),
.Y(n_1705)
);

AND2x2_ASAP7_75t_L g1706 ( 
.A(n_1700),
.B(n_1541),
.Y(n_1706)
);

NAND2xp5_ASAP7_75t_L g1707 ( 
.A(n_1704),
.B(n_1699),
.Y(n_1707)
);

INVx2_ASAP7_75t_L g1708 ( 
.A(n_1707),
.Y(n_1708)
);

INVx1_ASAP7_75t_L g1709 ( 
.A(n_1708),
.Y(n_1709)
);

OAI22xp33_ASAP7_75t_SL g1710 ( 
.A1(n_1708),
.A2(n_1705),
.B1(n_1703),
.B2(n_1706),
.Y(n_1710)
);

HB1xp67_ASAP7_75t_L g1711 ( 
.A(n_1709),
.Y(n_1711)
);

INVx2_ASAP7_75t_L g1712 ( 
.A(n_1710),
.Y(n_1712)
);

AOI22xp5_ASAP7_75t_SL g1713 ( 
.A1(n_1711),
.A2(n_1414),
.B1(n_1421),
.B2(n_1537),
.Y(n_1713)
);

OAI22xp5_ASAP7_75t_SL g1714 ( 
.A1(n_1712),
.A2(n_1395),
.B1(n_1366),
.B2(n_1525),
.Y(n_1714)
);

XNOR2xp5_ASAP7_75t_L g1715 ( 
.A(n_1714),
.B(n_1422),
.Y(n_1715)
);

OAI21xp5_ASAP7_75t_L g1716 ( 
.A1(n_1715),
.A2(n_1713),
.B(n_1402),
.Y(n_1716)
);

AOI221xp5_ASAP7_75t_L g1717 ( 
.A1(n_1716),
.A2(n_1543),
.B1(n_1520),
.B2(n_1533),
.C(n_1532),
.Y(n_1717)
);

AOI221xp5_ASAP7_75t_L g1718 ( 
.A1(n_1717),
.A2(n_1543),
.B1(n_1533),
.B2(n_1532),
.C(n_1530),
.Y(n_1718)
);

AOI211xp5_ASAP7_75t_L g1719 ( 
.A1(n_1718),
.A2(n_1408),
.B(n_1394),
.C(n_1527),
.Y(n_1719)
);


endmodule