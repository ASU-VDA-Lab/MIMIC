module fake_jpeg_27177_n_309 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_309);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_309;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_13;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_5),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_6),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_4),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

BUFx10_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

CKINVDCx16_ASAP7_75t_R g20 ( 
.A(n_2),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

BUFx12_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_2),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_0),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

OR2x2_ASAP7_75t_L g32 ( 
.A(n_15),
.B(n_12),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_32),
.B(n_37),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_15),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_33),
.B(n_35),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_22),
.Y(n_34)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_34),
.Y(n_60)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_31),
.Y(n_35)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_22),
.Y(n_36)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_31),
.B(n_11),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_31),
.Y(n_38)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_22),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_22),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_31),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_41),
.B(n_42),
.Y(n_56)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

INVx6_ASAP7_75t_SL g43 ( 
.A(n_17),
.Y(n_43)
);

CKINVDCx16_ASAP7_75t_R g59 ( 
.A(n_43),
.Y(n_59)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_13),
.Y(n_44)
);

AND2x2_ASAP7_75t_L g57 ( 
.A(n_44),
.B(n_13),
.Y(n_57)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_13),
.Y(n_45)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_45),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_37),
.B(n_13),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_46),
.B(n_17),
.Y(n_61)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_45),
.Y(n_49)
);

INVx8_ASAP7_75t_L g105 ( 
.A(n_49),
.Y(n_105)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_45),
.Y(n_50)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_50),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_38),
.A2(n_30),
.B1(n_25),
.B2(n_24),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_55),
.A2(n_20),
.B1(n_43),
.B2(n_25),
.Y(n_62)
);

OAI21xp5_ASAP7_75t_SL g83 ( 
.A1(n_57),
.A2(n_20),
.B(n_35),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_61),
.B(n_64),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_62),
.A2(n_29),
.B1(n_18),
.B2(n_26),
.Y(n_121)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_56),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_63),
.B(n_72),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_46),
.B(n_32),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_47),
.B(n_33),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g132 ( 
.A(n_65),
.B(n_66),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_58),
.B(n_32),
.Y(n_66)
);

INVx11_ASAP7_75t_L g68 ( 
.A(n_52),
.Y(n_68)
);

INVx8_ASAP7_75t_L g133 ( 
.A(n_68),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_46),
.B(n_17),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_69),
.B(n_79),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_47),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g134 ( 
.A(n_70),
.B(n_71),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_56),
.B(n_28),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_52),
.Y(n_72)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_51),
.Y(n_73)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_73),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_54),
.Y(n_74)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_74),
.Y(n_114)
);

OR2x4_ASAP7_75t_L g75 ( 
.A(n_58),
.B(n_57),
.Y(n_75)
);

OAI21xp5_ASAP7_75t_L g109 ( 
.A1(n_75),
.A2(n_94),
.B(n_103),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_L g76 ( 
.A1(n_60),
.A2(n_44),
.B1(n_42),
.B2(n_41),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_76),
.A2(n_81),
.B1(n_29),
.B2(n_18),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_58),
.B(n_16),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_77),
.B(n_78),
.Y(n_138)
);

INVx1_ASAP7_75t_SL g78 ( 
.A(n_57),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_57),
.B(n_17),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_51),
.Y(n_80)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_80),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_54),
.A2(n_30),
.B1(n_28),
.B2(n_16),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_59),
.B(n_34),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_82),
.B(n_84),
.Y(n_141)
);

AOI21xp5_ASAP7_75t_L g113 ( 
.A1(n_83),
.A2(n_0),
.B(n_1),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_59),
.B(n_24),
.Y(n_84)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_51),
.Y(n_85)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_85),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_55),
.B(n_17),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_86),
.B(n_97),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_52),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_87),
.Y(n_116)
);

AND2x2_ASAP7_75t_SL g88 ( 
.A(n_52),
.B(n_34),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_88),
.B(n_39),
.C(n_27),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_60),
.A2(n_43),
.B1(n_36),
.B2(n_45),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_89),
.A2(n_99),
.B1(n_26),
.B2(n_19),
.Y(n_127)
);

INVx5_ASAP7_75t_L g90 ( 
.A(n_53),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_90),
.A2(n_100),
.B1(n_91),
.B2(n_102),
.Y(n_124)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_53),
.Y(n_91)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_91),
.Y(n_117)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_48),
.Y(n_92)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_92),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_54),
.B(n_40),
.Y(n_93)
);

CKINVDCx16_ASAP7_75t_R g110 ( 
.A(n_93),
.Y(n_110)
);

A2O1A1Ixp33_ASAP7_75t_L g94 ( 
.A1(n_60),
.A2(n_23),
.B(n_21),
.C(n_35),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_53),
.B(n_21),
.Y(n_95)
);

CKINVDCx16_ASAP7_75t_R g137 ( 
.A(n_95),
.Y(n_137)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_48),
.Y(n_96)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_96),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_53),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_48),
.Y(n_98)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_98),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_60),
.A2(n_36),
.B1(n_45),
.B2(n_23),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_49),
.Y(n_100)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_49),
.Y(n_101)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_101),
.Y(n_140)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_50),
.Y(n_102)
);

CKINVDCx16_ASAP7_75t_R g139 ( 
.A(n_102),
.Y(n_139)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_50),
.B(n_40),
.Y(n_103)
);

HB1xp67_ASAP7_75t_L g104 ( 
.A(n_51),
.Y(n_104)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_104),
.Y(n_130)
);

MAJx2_ASAP7_75t_L g107 ( 
.A(n_75),
.B(n_22),
.C(n_39),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_107),
.B(n_136),
.C(n_14),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_108),
.A2(n_127),
.B1(n_131),
.B2(n_103),
.Y(n_149)
);

AND2x2_ASAP7_75t_L g160 ( 
.A(n_111),
.B(n_74),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_SL g143 ( 
.A1(n_113),
.A2(n_88),
.B(n_120),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_121),
.A2(n_128),
.B1(n_99),
.B2(n_88),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_61),
.B(n_27),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_122),
.B(n_126),
.Y(n_154)
);

INVxp67_ASAP7_75t_L g153 ( 
.A(n_124),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_69),
.B(n_27),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_78),
.A2(n_29),
.B1(n_18),
.B2(n_19),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_86),
.A2(n_79),
.B1(n_63),
.B2(n_64),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g136 ( 
.A(n_83),
.B(n_26),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_L g142 ( 
.A1(n_109),
.A2(n_94),
.B(n_103),
.Y(n_142)
);

A2O1A1Ixp33_ASAP7_75t_SL g200 ( 
.A1(n_142),
.A2(n_166),
.B(n_169),
.C(n_1),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_143),
.B(n_157),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_144),
.A2(n_160),
.B1(n_167),
.B2(n_145),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_106),
.B(n_80),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_145),
.B(n_146),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_134),
.B(n_85),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_132),
.B(n_73),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_147),
.B(n_148),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_141),
.B(n_137),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_149),
.A2(n_121),
.B1(n_130),
.B2(n_119),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_110),
.B(n_98),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_150),
.B(n_156),
.Y(n_193)
);

CKINVDCx16_ASAP7_75t_R g151 ( 
.A(n_125),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_151),
.B(n_161),
.Y(n_174)
);

OR2x2_ASAP7_75t_L g152 ( 
.A(n_120),
.B(n_89),
.Y(n_152)
);

OR2x2_ASAP7_75t_L g195 ( 
.A(n_152),
.B(n_159),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_131),
.A2(n_72),
.B1(n_97),
.B2(n_90),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_155),
.A2(n_158),
.B1(n_115),
.B2(n_135),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_106),
.B(n_92),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_127),
.A2(n_68),
.B1(n_101),
.B2(n_96),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_SL g159 ( 
.A(n_138),
.B(n_9),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_122),
.B(n_67),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_126),
.B(n_118),
.Y(n_162)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_162),
.Y(n_194)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_133),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_163),
.B(n_133),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_118),
.B(n_67),
.Y(n_164)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_164),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_SL g165 ( 
.A1(n_113),
.A2(n_105),
.B(n_19),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_165),
.B(n_128),
.Y(n_171)
);

AOI21xp5_ASAP7_75t_L g166 ( 
.A1(n_109),
.A2(n_0),
.B(n_1),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_136),
.B(n_111),
.Y(n_167)
);

CKINVDCx14_ASAP7_75t_R g176 ( 
.A(n_167),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_116),
.B(n_105),
.Y(n_168)
);

OAI32xp33_ASAP7_75t_L g179 ( 
.A1(n_168),
.A2(n_135),
.A3(n_119),
.B1(n_115),
.B2(n_114),
.Y(n_179)
);

AO21x1_ASAP7_75t_L g169 ( 
.A1(n_107),
.A2(n_14),
.B(n_2),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_116),
.B(n_14),
.Y(n_170)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_170),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_SL g216 ( 
.A1(n_171),
.A2(n_187),
.B(n_200),
.Y(n_216)
);

BUFx24_ASAP7_75t_SL g172 ( 
.A(n_148),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_172),
.B(n_175),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_168),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_150),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_177),
.B(n_178),
.Y(n_223)
);

CKINVDCx16_ASAP7_75t_R g178 ( 
.A(n_170),
.Y(n_178)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_179),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_180),
.A2(n_186),
.B1(n_197),
.B2(n_144),
.Y(n_204)
);

HB1xp67_ASAP7_75t_L g182 ( 
.A(n_161),
.Y(n_182)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_182),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_183),
.A2(n_154),
.B1(n_162),
.B2(n_142),
.Y(n_213)
);

OAI21x1_ASAP7_75t_L g187 ( 
.A1(n_169),
.A2(n_130),
.B(n_12),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_146),
.Y(n_188)
);

AOI22xp33_ASAP7_75t_SL g202 ( 
.A1(n_188),
.A2(n_190),
.B1(n_191),
.B2(n_192),
.Y(n_202)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_189),
.Y(n_220)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_147),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_164),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_155),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_157),
.B(n_140),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_196),
.B(n_199),
.C(n_160),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_149),
.A2(n_114),
.B1(n_117),
.B2(n_129),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_157),
.B(n_140),
.Y(n_199)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_179),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_203),
.B(n_209),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_204),
.A2(n_214),
.B1(n_217),
.B2(n_209),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_205),
.B(n_196),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_193),
.B(n_156),
.Y(n_207)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_207),
.Y(n_234)
);

BUFx6f_ASAP7_75t_L g208 ( 
.A(n_197),
.Y(n_208)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_208),
.Y(n_229)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_180),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_L g210 ( 
.A1(n_195),
.A2(n_142),
.B(n_166),
.Y(n_210)
);

AOI21xp33_ASAP7_75t_L g236 ( 
.A1(n_210),
.A2(n_185),
.B(n_184),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_193),
.B(n_181),
.Y(n_212)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_212),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_213),
.A2(n_219),
.B1(n_199),
.B2(n_112),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_198),
.A2(n_160),
.B1(n_153),
.B2(n_143),
.Y(n_214)
);

AOI21xp5_ASAP7_75t_L g215 ( 
.A1(n_200),
.A2(n_165),
.B(n_169),
.Y(n_215)
);

CKINVDCx14_ASAP7_75t_R g233 ( 
.A(n_215),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_198),
.A2(n_160),
.B1(n_152),
.B2(n_151),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_SL g218 ( 
.A1(n_200),
.A2(n_152),
.B(n_158),
.Y(n_218)
);

CKINVDCx14_ASAP7_75t_R g243 ( 
.A(n_218),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_183),
.A2(n_154),
.B1(n_163),
.B2(n_117),
.Y(n_219)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_174),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_221),
.B(n_224),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_181),
.B(n_159),
.Y(n_222)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_222),
.Y(n_242)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_185),
.Y(n_224)
);

AOI21xp5_ASAP7_75t_L g225 ( 
.A1(n_200),
.A2(n_139),
.B(n_123),
.Y(n_225)
);

CKINVDCx16_ASAP7_75t_R g231 ( 
.A(n_225),
.Y(n_231)
);

O2A1O1Ixp33_ASAP7_75t_L g226 ( 
.A1(n_195),
.A2(n_129),
.B(n_112),
.C(n_123),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_226),
.B(n_194),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_SL g259 ( 
.A1(n_228),
.A2(n_241),
.B(n_218),
.Y(n_259)
);

INVx1_ASAP7_75t_SL g230 ( 
.A(n_212),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_230),
.B(n_244),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_232),
.B(n_246),
.C(n_222),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_SL g249 ( 
.A(n_236),
.B(n_237),
.C(n_210),
.Y(n_249)
);

XNOR2x1_ASAP7_75t_L g237 ( 
.A(n_205),
.B(n_173),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_214),
.B(n_173),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_238),
.B(n_217),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_L g239 ( 
.A1(n_203),
.A2(n_194),
.B1(n_171),
.B2(n_176),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_L g257 ( 
.A1(n_239),
.A2(n_206),
.B1(n_202),
.B2(n_221),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_223),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_245),
.B(n_204),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_219),
.B(n_11),
.C(n_10),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_247),
.B(n_251),
.Y(n_277)
);

HB1xp67_ASAP7_75t_L g248 ( 
.A(n_235),
.Y(n_248)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_248),
.Y(n_272)
);

MAJx2_ASAP7_75t_L g275 ( 
.A(n_249),
.B(n_256),
.C(n_215),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_250),
.A2(n_257),
.B1(n_243),
.B2(n_231),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_238),
.B(n_216),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_232),
.B(n_216),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_252),
.B(n_254),
.C(n_258),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_245),
.B(n_224),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_235),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_255),
.A2(n_261),
.B1(n_264),
.B2(n_234),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_237),
.B(n_201),
.C(n_207),
.Y(n_258)
);

INVxp67_ASAP7_75t_L g274 ( 
.A(n_259),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_244),
.B(n_211),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_L g266 ( 
.A1(n_260),
.A2(n_262),
.B1(n_242),
.B2(n_240),
.Y(n_266)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_241),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_230),
.B(n_220),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_242),
.B(n_201),
.Y(n_263)
);

OAI21xp5_ASAP7_75t_L g268 ( 
.A1(n_263),
.A2(n_226),
.B(n_225),
.Y(n_268)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_227),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_265),
.B(n_2),
.Y(n_285)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_266),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_L g267 ( 
.A1(n_253),
.A2(n_227),
.B1(n_229),
.B2(n_246),
.Y(n_267)
);

INVxp67_ASAP7_75t_L g280 ( 
.A(n_267),
.Y(n_280)
);

AOI21xp5_ASAP7_75t_L g282 ( 
.A1(n_268),
.A2(n_269),
.B(n_252),
.Y(n_282)
);

AND2x2_ASAP7_75t_L g269 ( 
.A(n_251),
.B(n_233),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_258),
.B(n_240),
.C(n_234),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_271),
.B(n_275),
.C(n_270),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_273),
.B(n_1),
.Y(n_284)
);

BUFx6f_ASAP7_75t_L g276 ( 
.A(n_259),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_276),
.B(n_3),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_274),
.A2(n_229),
.B1(n_254),
.B2(n_247),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_279),
.A2(n_283),
.B1(n_269),
.B2(n_275),
.Y(n_292)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_281),
.B(n_282),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_274),
.A2(n_208),
.B1(n_256),
.B2(n_3),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_SL g289 ( 
.A(n_284),
.B(n_4),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_285),
.A2(n_271),
.B1(n_6),
.B2(n_7),
.Y(n_293)
);

CKINVDCx16_ASAP7_75t_R g291 ( 
.A(n_286),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_283),
.B(n_276),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_288),
.B(n_289),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_280),
.B(n_272),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_290),
.B(n_292),
.Y(n_296)
);

INVxp67_ASAP7_75t_L g299 ( 
.A(n_293),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_280),
.A2(n_277),
.B1(n_270),
.B2(n_7),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_294),
.A2(n_278),
.B1(n_279),
.B2(n_7),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_297),
.B(n_298),
.Y(n_300)
);

AOI21xp5_ASAP7_75t_L g298 ( 
.A1(n_292),
.A2(n_281),
.B(n_277),
.Y(n_298)
);

AOI21xp5_ASAP7_75t_L g301 ( 
.A1(n_296),
.A2(n_287),
.B(n_294),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_L g303 ( 
.A1(n_301),
.A2(n_299),
.B1(n_300),
.B2(n_287),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_295),
.B(n_291),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_302),
.B(n_5),
.C(n_6),
.Y(n_304)
);

AOI21xp5_ASAP7_75t_SL g305 ( 
.A1(n_303),
.A2(n_304),
.B(n_5),
.Y(n_305)
);

BUFx24_ASAP7_75t_SL g306 ( 
.A(n_305),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g307 ( 
.A(n_306),
.B(n_8),
.Y(n_307)
);

OAI21xp5_ASAP7_75t_L g308 ( 
.A1(n_307),
.A2(n_6),
.B(n_7),
.Y(n_308)
);

XOR2xp5_ASAP7_75t_L g309 ( 
.A(n_308),
.B(n_8),
.Y(n_309)
);


endmodule