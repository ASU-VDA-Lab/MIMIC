module fake_netlist_1_3644_n_557 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_6, n_4, n_40, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_557);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_6;
input n_4;
input n_40;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_557;
wire n_117;
wire n_361;
wire n_513;
wire n_185;
wire n_407;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_154;
wire n_328;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_353;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_532;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_411;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_366;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_244;
wire n_540;
wire n_119;
wire n_141;
wire n_517;
wire n_479;
wire n_97;
wire n_167;
wire n_554;
wire n_447;
wire n_171;
wire n_196;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_367;
wire n_250;
wire n_85;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_172;
wire n_329;
wire n_251;
wire n_525;
wire n_218;
wire n_507;
wire n_271;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_107;
wire n_403;
wire n_516;
wire n_254;
wire n_549;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_87;
wire n_379;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_370;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_245;
wire n_357;
wire n_90;
wire n_260;
wire n_78;
wire n_539;
wire n_201;
wire n_197;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_126;
wire n_178;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_376;
wire n_552;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_435;
wire n_216;
wire n_147;
wire n_148;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_497;
wire n_339;
wire n_240;
wire n_378;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_335;
wire n_272;
wire n_534;
wire n_531;
wire n_397;
wire n_146;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_198;
wire n_169;
wire n_424;
wire n_156;
wire n_124;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_258;
wire n_253;
wire n_515;
wire n_84;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_521;
wire n_469;
wire n_123;
wire n_457;
wire n_223;
wire n_494;
wire n_480;
wire n_372;
wire n_453;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_425;
wire n_332;
wire n_414;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_132;
wire n_109;
wire n_99;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g78 ( .A(n_47), .Y(n_78) );
CKINVDCx5p33_ASAP7_75t_R g79 ( .A(n_17), .Y(n_79) );
CKINVDCx20_ASAP7_75t_R g80 ( .A(n_21), .Y(n_80) );
BUFx3_ASAP7_75t_L g81 ( .A(n_72), .Y(n_81) );
INVxp33_ASAP7_75t_SL g82 ( .A(n_62), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_26), .Y(n_83) );
INVx1_ASAP7_75t_SL g84 ( .A(n_53), .Y(n_84) );
CKINVDCx5p33_ASAP7_75t_R g85 ( .A(n_73), .Y(n_85) );
CKINVDCx20_ASAP7_75t_R g86 ( .A(n_20), .Y(n_86) );
CKINVDCx16_ASAP7_75t_R g87 ( .A(n_11), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_6), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_18), .Y(n_89) );
CKINVDCx5p33_ASAP7_75t_R g90 ( .A(n_32), .Y(n_90) );
BUFx6f_ASAP7_75t_L g91 ( .A(n_10), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_41), .Y(n_92) );
CKINVDCx5p33_ASAP7_75t_R g93 ( .A(n_75), .Y(n_93) );
INVx2_ASAP7_75t_SL g94 ( .A(n_13), .Y(n_94) );
BUFx10_ASAP7_75t_L g95 ( .A(n_0), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_68), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_77), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_64), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_7), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_34), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_25), .Y(n_101) );
CKINVDCx20_ASAP7_75t_R g102 ( .A(n_65), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_66), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_37), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_18), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_3), .Y(n_106) );
INVxp67_ASAP7_75t_SL g107 ( .A(n_42), .Y(n_107) );
BUFx10_ASAP7_75t_L g108 ( .A(n_8), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_58), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_5), .Y(n_110) );
CKINVDCx5p33_ASAP7_75t_R g111 ( .A(n_3), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_15), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_9), .Y(n_113) );
INVxp33_ASAP7_75t_SL g114 ( .A(n_79), .Y(n_114) );
INVx1_ASAP7_75t_SL g115 ( .A(n_80), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_78), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_83), .Y(n_117) );
OR2x6_ASAP7_75t_L g118 ( .A(n_94), .B(n_35), .Y(n_118) );
BUFx6f_ASAP7_75t_L g119 ( .A(n_81), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_92), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_96), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_97), .Y(n_122) );
HB1xp67_ASAP7_75t_L g123 ( .A(n_79), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_98), .Y(n_124) );
AND2x2_ASAP7_75t_L g125 ( .A(n_87), .B(n_0), .Y(n_125) );
OAI21x1_ASAP7_75t_L g126 ( .A1(n_100), .A2(n_36), .B(n_74), .Y(n_126) );
INVx3_ASAP7_75t_L g127 ( .A(n_91), .Y(n_127) );
BUFx6f_ASAP7_75t_L g128 ( .A(n_81), .Y(n_128) );
CKINVDCx20_ASAP7_75t_R g129 ( .A(n_80), .Y(n_129) );
INVx1_ASAP7_75t_L g130 ( .A(n_101), .Y(n_130) );
BUFx6f_ASAP7_75t_L g131 ( .A(n_91), .Y(n_131) );
INVx1_ASAP7_75t_L g132 ( .A(n_103), .Y(n_132) );
INVx3_ASAP7_75t_L g133 ( .A(n_91), .Y(n_133) );
OAI22xp5_ASAP7_75t_SL g134 ( .A1(n_111), .A2(n_1), .B1(n_2), .B2(n_4), .Y(n_134) );
INVx5_ASAP7_75t_L g135 ( .A(n_91), .Y(n_135) );
BUFx2_ASAP7_75t_L g136 ( .A(n_111), .Y(n_136) );
INVx1_ASAP7_75t_L g137 ( .A(n_104), .Y(n_137) );
CKINVDCx20_ASAP7_75t_R g138 ( .A(n_129), .Y(n_138) );
NAND2xp5_ASAP7_75t_L g139 ( .A(n_136), .B(n_85), .Y(n_139) );
INVx1_ASAP7_75t_L g140 ( .A(n_127), .Y(n_140) );
NAND2xp5_ASAP7_75t_SL g141 ( .A(n_114), .B(n_85), .Y(n_141) );
INVx1_ASAP7_75t_L g142 ( .A(n_127), .Y(n_142) );
BUFx6f_ASAP7_75t_L g143 ( .A(n_131), .Y(n_143) );
NAND2x1p5_ASAP7_75t_L g144 ( .A(n_126), .B(n_109), .Y(n_144) );
INVx2_ASAP7_75t_SL g145 ( .A(n_136), .Y(n_145) );
BUFx6f_ASAP7_75t_L g146 ( .A(n_131), .Y(n_146) );
BUFx6f_ASAP7_75t_L g147 ( .A(n_131), .Y(n_147) );
AND2x4_ASAP7_75t_L g148 ( .A(n_116), .B(n_94), .Y(n_148) );
INVx2_ASAP7_75t_L g149 ( .A(n_119), .Y(n_149) );
INVx2_ASAP7_75t_L g150 ( .A(n_119), .Y(n_150) );
BUFx2_ASAP7_75t_L g151 ( .A(n_123), .Y(n_151) );
CKINVDCx5p33_ASAP7_75t_R g152 ( .A(n_115), .Y(n_152) );
NAND2xp33_ASAP7_75t_L g153 ( .A(n_116), .B(n_90), .Y(n_153) );
NOR2xp33_ASAP7_75t_L g154 ( .A(n_117), .B(n_82), .Y(n_154) );
INVxp67_ASAP7_75t_L g155 ( .A(n_123), .Y(n_155) );
AOI22xp5_ASAP7_75t_L g156 ( .A1(n_125), .A2(n_102), .B1(n_86), .B2(n_82), .Y(n_156) );
BUFx4f_ASAP7_75t_L g157 ( .A(n_118), .Y(n_157) );
INVxp33_ASAP7_75t_L g158 ( .A(n_125), .Y(n_158) );
AND2x4_ASAP7_75t_L g159 ( .A(n_117), .B(n_88), .Y(n_159) );
NOR2xp33_ASAP7_75t_R g160 ( .A(n_120), .B(n_86), .Y(n_160) );
AND2x2_ASAP7_75t_L g161 ( .A(n_120), .B(n_95), .Y(n_161) );
BUFx10_ASAP7_75t_L g162 ( .A(n_118), .Y(n_162) );
OAI22xp5_ASAP7_75t_L g163 ( .A1(n_118), .A2(n_102), .B1(n_112), .B2(n_110), .Y(n_163) );
INVx2_ASAP7_75t_L g164 ( .A(n_119), .Y(n_164) );
NAND2xp5_ASAP7_75t_L g165 ( .A(n_154), .B(n_121), .Y(n_165) );
NAND2xp5_ASAP7_75t_L g166 ( .A(n_161), .B(n_121), .Y(n_166) );
INVx5_ASAP7_75t_L g167 ( .A(n_162), .Y(n_167) );
INVx2_ASAP7_75t_L g168 ( .A(n_149), .Y(n_168) );
NAND2xp5_ASAP7_75t_L g169 ( .A(n_161), .B(n_122), .Y(n_169) );
AOI22xp5_ASAP7_75t_L g170 ( .A1(n_163), .A2(n_118), .B1(n_134), .B2(n_115), .Y(n_170) );
INVx4_ASAP7_75t_L g171 ( .A(n_157), .Y(n_171) );
AND2x2_ASAP7_75t_L g172 ( .A(n_151), .B(n_95), .Y(n_172) );
A2O1A1Ixp33_ASAP7_75t_L g173 ( .A1(n_157), .A2(n_126), .B(n_124), .C(n_130), .Y(n_173) );
HB1xp67_ASAP7_75t_L g174 ( .A(n_151), .Y(n_174) );
INVx1_ASAP7_75t_L g175 ( .A(n_148), .Y(n_175) );
NOR3xp33_ASAP7_75t_L g176 ( .A(n_152), .B(n_134), .C(n_113), .Y(n_176) );
NAND2xp5_ASAP7_75t_SL g177 ( .A(n_157), .B(n_122), .Y(n_177) );
INVx1_ASAP7_75t_L g178 ( .A(n_148), .Y(n_178) );
BUFx4f_ASAP7_75t_L g179 ( .A(n_145), .Y(n_179) );
AOI22xp5_ASAP7_75t_L g180 ( .A1(n_155), .A2(n_118), .B1(n_137), .B2(n_132), .Y(n_180) );
INVx2_ASAP7_75t_SL g181 ( .A(n_145), .Y(n_181) );
OR2x6_ASAP7_75t_L g182 ( .A(n_148), .B(n_118), .Y(n_182) );
INVx1_ASAP7_75t_L g183 ( .A(n_148), .Y(n_183) );
NAND2xp5_ASAP7_75t_L g184 ( .A(n_159), .B(n_124), .Y(n_184) );
AND2x4_ASAP7_75t_L g185 ( .A(n_159), .B(n_130), .Y(n_185) );
NAND2xp5_ASAP7_75t_SL g186 ( .A(n_162), .B(n_132), .Y(n_186) );
NOR2xp33_ASAP7_75t_R g187 ( .A(n_152), .B(n_90), .Y(n_187) );
BUFx3_ASAP7_75t_L g188 ( .A(n_162), .Y(n_188) );
INVx2_ASAP7_75t_SL g189 ( .A(n_160), .Y(n_189) );
AOI22xp33_ASAP7_75t_SL g190 ( .A1(n_139), .A2(n_108), .B1(n_95), .B2(n_93), .Y(n_190) );
INVx1_ASAP7_75t_L g191 ( .A(n_159), .Y(n_191) );
OAI22xp5_ASAP7_75t_L g192 ( .A1(n_158), .A2(n_137), .B1(n_89), .B2(n_99), .Y(n_192) );
INVx1_ASAP7_75t_L g193 ( .A(n_159), .Y(n_193) );
BUFx6f_ASAP7_75t_L g194 ( .A(n_144), .Y(n_194) );
INVx1_ASAP7_75t_L g195 ( .A(n_153), .Y(n_195) );
NAND2xp5_ASAP7_75t_SL g196 ( .A(n_144), .B(n_126), .Y(n_196) );
BUFx6f_ASAP7_75t_L g197 ( .A(n_144), .Y(n_197) );
OR2x6_ASAP7_75t_L g198 ( .A(n_141), .B(n_105), .Y(n_198) );
BUFx3_ASAP7_75t_L g199 ( .A(n_149), .Y(n_199) );
INVx1_ASAP7_75t_L g200 ( .A(n_140), .Y(n_200) );
AOI21xp5_ASAP7_75t_L g201 ( .A1(n_196), .A2(n_164), .B(n_150), .Y(n_201) );
OAI22xp5_ASAP7_75t_L g202 ( .A1(n_180), .A2(n_156), .B1(n_93), .B2(n_106), .Y(n_202) );
CKINVDCx8_ASAP7_75t_R g203 ( .A(n_167), .Y(n_203) );
OAI22xp5_ASAP7_75t_L g204 ( .A1(n_170), .A2(n_156), .B1(n_107), .B2(n_91), .Y(n_204) );
HB1xp67_ASAP7_75t_L g205 ( .A(n_174), .Y(n_205) );
NAND2xp5_ASAP7_75t_SL g206 ( .A(n_167), .B(n_84), .Y(n_206) );
INVx2_ASAP7_75t_L g207 ( .A(n_200), .Y(n_207) );
INVx1_ASAP7_75t_L g208 ( .A(n_191), .Y(n_208) );
NAND2xp5_ASAP7_75t_L g209 ( .A(n_185), .B(n_108), .Y(n_209) );
O2A1O1Ixp33_ASAP7_75t_L g210 ( .A1(n_192), .A2(n_142), .B(n_140), .C(n_127), .Y(n_210) );
AOI22xp5_ASAP7_75t_L g211 ( .A1(n_185), .A2(n_119), .B1(n_128), .B2(n_108), .Y(n_211) );
A2O1A1Ixp33_ASAP7_75t_L g212 ( .A1(n_175), .A2(n_127), .B(n_133), .C(n_142), .Y(n_212) );
INVx3_ASAP7_75t_L g213 ( .A(n_171), .Y(n_213) );
AOI22xp5_ASAP7_75t_L g214 ( .A1(n_185), .A2(n_119), .B1(n_128), .B2(n_133), .Y(n_214) );
NAND2xp5_ASAP7_75t_L g215 ( .A(n_166), .B(n_119), .Y(n_215) );
AND2x4_ASAP7_75t_L g216 ( .A(n_171), .B(n_1), .Y(n_216) );
AND2x2_ASAP7_75t_L g217 ( .A(n_174), .B(n_128), .Y(n_217) );
NOR2xp33_ASAP7_75t_L g218 ( .A(n_181), .B(n_138), .Y(n_218) );
AOI21xp5_ASAP7_75t_L g219 ( .A1(n_196), .A2(n_164), .B(n_150), .Y(n_219) );
AOI22xp33_ASAP7_75t_L g220 ( .A1(n_193), .A2(n_128), .B1(n_133), .B2(n_135), .Y(n_220) );
AOI22xp33_ASAP7_75t_L g221 ( .A1(n_178), .A2(n_128), .B1(n_133), .B2(n_135), .Y(n_221) );
BUFx3_ASAP7_75t_L g222 ( .A(n_167), .Y(n_222) );
NAND2xp5_ASAP7_75t_L g223 ( .A(n_169), .B(n_128), .Y(n_223) );
INVx2_ASAP7_75t_L g224 ( .A(n_168), .Y(n_224) );
NOR2xp33_ASAP7_75t_L g225 ( .A(n_172), .B(n_2), .Y(n_225) );
AND2x4_ASAP7_75t_L g226 ( .A(n_167), .B(n_4), .Y(n_226) );
AND2x4_ASAP7_75t_L g227 ( .A(n_188), .B(n_5), .Y(n_227) );
BUFx2_ASAP7_75t_L g228 ( .A(n_187), .Y(n_228) );
INVx1_ASAP7_75t_L g229 ( .A(n_183), .Y(n_229) );
AOI22xp33_ASAP7_75t_L g230 ( .A1(n_182), .A2(n_135), .B1(n_131), .B2(n_143), .Y(n_230) );
AND2x2_ASAP7_75t_L g231 ( .A(n_184), .B(n_6), .Y(n_231) );
INVx2_ASAP7_75t_L g232 ( .A(n_168), .Y(n_232) );
AOI22xp33_ASAP7_75t_L g233 ( .A1(n_182), .A2(n_135), .B1(n_131), .B2(n_143), .Y(n_233) );
BUFx6f_ASAP7_75t_L g234 ( .A(n_194), .Y(n_234) );
INVx4_ASAP7_75t_L g235 ( .A(n_182), .Y(n_235) );
OAI21x1_ASAP7_75t_L g236 ( .A1(n_201), .A2(n_177), .B(n_186), .Y(n_236) );
INVx1_ASAP7_75t_L g237 ( .A(n_207), .Y(n_237) );
NOR2xp33_ASAP7_75t_L g238 ( .A(n_205), .B(n_198), .Y(n_238) );
INVx1_ASAP7_75t_L g239 ( .A(n_207), .Y(n_239) );
INVx2_ASAP7_75t_L g240 ( .A(n_234), .Y(n_240) );
INVx6_ASAP7_75t_L g241 ( .A(n_235), .Y(n_241) );
NAND3x1_ASAP7_75t_L g242 ( .A(n_225), .B(n_176), .C(n_165), .Y(n_242) );
OAI21xp5_ASAP7_75t_L g243 ( .A1(n_212), .A2(n_173), .B(n_177), .Y(n_243) );
INVx1_ASAP7_75t_L g244 ( .A(n_207), .Y(n_244) );
INVx1_ASAP7_75t_L g245 ( .A(n_229), .Y(n_245) );
AND2x4_ASAP7_75t_L g246 ( .A(n_235), .B(n_188), .Y(n_246) );
INVx1_ASAP7_75t_L g247 ( .A(n_229), .Y(n_247) );
OAI21x1_ASAP7_75t_L g248 ( .A1(n_219), .A2(n_186), .B(n_195), .Y(n_248) );
CKINVDCx16_ASAP7_75t_R g249 ( .A(n_228), .Y(n_249) );
INVx3_ASAP7_75t_L g250 ( .A(n_203), .Y(n_250) );
NAND2xp5_ASAP7_75t_L g251 ( .A(n_204), .B(n_187), .Y(n_251) );
OR2x6_ASAP7_75t_L g252 ( .A(n_235), .B(n_227), .Y(n_252) );
AOI21xp5_ASAP7_75t_L g253 ( .A1(n_224), .A2(n_173), .B(n_197), .Y(n_253) );
OAI21xp33_ASAP7_75t_SL g254 ( .A1(n_235), .A2(n_198), .B(n_189), .Y(n_254) );
HB1xp67_ASAP7_75t_L g255 ( .A(n_227), .Y(n_255) );
HB1xp67_ASAP7_75t_L g256 ( .A(n_227), .Y(n_256) );
INVx1_ASAP7_75t_L g257 ( .A(n_208), .Y(n_257) );
BUFx6f_ASAP7_75t_L g258 ( .A(n_234), .Y(n_258) );
OAI21x1_ASAP7_75t_L g259 ( .A1(n_215), .A2(n_197), .B(n_194), .Y(n_259) );
INVx2_ASAP7_75t_L g260 ( .A(n_234), .Y(n_260) );
INVx1_ASAP7_75t_L g261 ( .A(n_208), .Y(n_261) );
OAI21x1_ASAP7_75t_L g262 ( .A1(n_223), .A2(n_197), .B(n_194), .Y(n_262) );
AOI222xp33_ASAP7_75t_L g263 ( .A1(n_202), .A2(n_179), .B1(n_190), .B2(n_198), .C1(n_194), .C2(n_197), .Y(n_263) );
AOI222xp33_ASAP7_75t_L g264 ( .A1(n_238), .A2(n_179), .B1(n_218), .B2(n_216), .C1(n_228), .C2(n_227), .Y(n_264) );
INVx1_ASAP7_75t_L g265 ( .A(n_237), .Y(n_265) );
NAND3xp33_ASAP7_75t_L g266 ( .A(n_243), .B(n_211), .C(n_226), .Y(n_266) );
AOI22xp33_ASAP7_75t_L g267 ( .A1(n_263), .A2(n_216), .B1(n_231), .B2(n_226), .Y(n_267) );
BUFx2_ASAP7_75t_L g268 ( .A(n_252), .Y(n_268) );
AND2x4_ASAP7_75t_L g269 ( .A(n_252), .B(n_222), .Y(n_269) );
INVx1_ASAP7_75t_L g270 ( .A(n_237), .Y(n_270) );
AOI22xp33_ASAP7_75t_L g271 ( .A1(n_252), .A2(n_216), .B1(n_231), .B2(n_226), .Y(n_271) );
AOI22xp33_ASAP7_75t_L g272 ( .A1(n_252), .A2(n_216), .B1(n_226), .B2(n_217), .Y(n_272) );
OA21x2_ASAP7_75t_L g273 ( .A1(n_259), .A2(n_211), .B(n_214), .Y(n_273) );
INVx2_ASAP7_75t_L g274 ( .A(n_239), .Y(n_274) );
NAND2xp5_ASAP7_75t_L g275 ( .A(n_245), .B(n_213), .Y(n_275) );
O2A1O1Ixp33_ASAP7_75t_L g276 ( .A1(n_254), .A2(n_209), .B(n_206), .C(n_210), .Y(n_276) );
OAI21xp5_ASAP7_75t_L g277 ( .A1(n_253), .A2(n_217), .B(n_214), .Y(n_277) );
AOI221xp5_ASAP7_75t_L g278 ( .A1(n_254), .A2(n_213), .B1(n_221), .B2(n_220), .C(n_230), .Y(n_278) );
INVx1_ASAP7_75t_L g279 ( .A(n_239), .Y(n_279) );
AOI22xp33_ASAP7_75t_L g280 ( .A1(n_252), .A2(n_213), .B1(n_222), .B2(n_233), .Y(n_280) );
BUFx3_ASAP7_75t_L g281 ( .A(n_241), .Y(n_281) );
INVx2_ASAP7_75t_L g282 ( .A(n_244), .Y(n_282) );
AOI221xp5_ASAP7_75t_L g283 ( .A1(n_245), .A2(n_213), .B1(n_222), .B2(n_224), .C(n_232), .Y(n_283) );
CKINVDCx5p33_ASAP7_75t_R g284 ( .A(n_249), .Y(n_284) );
OAI221xp5_ASAP7_75t_L g285 ( .A1(n_251), .A2(n_203), .B1(n_232), .B2(n_135), .C(n_234), .Y(n_285) );
AOI21xp33_ASAP7_75t_L g286 ( .A1(n_242), .A2(n_234), .B(n_131), .Y(n_286) );
INVx1_ASAP7_75t_L g287 ( .A(n_274), .Y(n_287) );
AND2x4_ASAP7_75t_L g288 ( .A(n_274), .B(n_244), .Y(n_288) );
AND2x4_ASAP7_75t_L g289 ( .A(n_274), .B(n_240), .Y(n_289) );
INVx2_ASAP7_75t_L g290 ( .A(n_282), .Y(n_290) );
AND2x2_ASAP7_75t_L g291 ( .A(n_282), .B(n_255), .Y(n_291) );
INVx2_ASAP7_75t_L g292 ( .A(n_282), .Y(n_292) );
INVx2_ASAP7_75t_L g293 ( .A(n_265), .Y(n_293) );
INVx1_ASAP7_75t_L g294 ( .A(n_265), .Y(n_294) );
AND2x4_ASAP7_75t_L g295 ( .A(n_269), .B(n_240), .Y(n_295) );
AND2x2_ASAP7_75t_L g296 ( .A(n_270), .B(n_256), .Y(n_296) );
BUFx3_ASAP7_75t_L g297 ( .A(n_269), .Y(n_297) );
OAI22xp5_ASAP7_75t_L g298 ( .A1(n_267), .A2(n_242), .B1(n_261), .B2(n_257), .Y(n_298) );
AND2x2_ASAP7_75t_L g299 ( .A(n_270), .B(n_247), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g300 ( .A(n_279), .B(n_247), .Y(n_300) );
OAI222xp33_ASAP7_75t_L g301 ( .A1(n_271), .A2(n_249), .B1(n_250), .B2(n_257), .C1(n_261), .C2(n_246), .Y(n_301) );
INVx1_ASAP7_75t_L g302 ( .A(n_279), .Y(n_302) );
NAND2xp5_ASAP7_75t_L g303 ( .A(n_275), .B(n_260), .Y(n_303) );
INVx1_ASAP7_75t_SL g304 ( .A(n_269), .Y(n_304) );
HB1xp67_ASAP7_75t_L g305 ( .A(n_268), .Y(n_305) );
INVx1_ASAP7_75t_L g306 ( .A(n_275), .Y(n_306) );
OR2x2_ASAP7_75t_L g307 ( .A(n_268), .B(n_246), .Y(n_307) );
INVx1_ASAP7_75t_L g308 ( .A(n_277), .Y(n_308) );
INVx2_ASAP7_75t_L g309 ( .A(n_273), .Y(n_309) );
AND2x2_ASAP7_75t_L g310 ( .A(n_308), .B(n_277), .Y(n_310) );
AND2x2_ASAP7_75t_L g311 ( .A(n_308), .B(n_273), .Y(n_311) );
BUFx2_ASAP7_75t_L g312 ( .A(n_305), .Y(n_312) );
INVx1_ASAP7_75t_L g313 ( .A(n_293), .Y(n_313) );
BUFx2_ASAP7_75t_L g314 ( .A(n_305), .Y(n_314) );
AND2x2_ASAP7_75t_L g315 ( .A(n_290), .B(n_273), .Y(n_315) );
INVx1_ASAP7_75t_L g316 ( .A(n_293), .Y(n_316) );
NOR2x1p5_ASAP7_75t_L g317 ( .A(n_297), .B(n_269), .Y(n_317) );
AOI211xp5_ASAP7_75t_L g318 ( .A1(n_298), .A2(n_286), .B(n_284), .C(n_285), .Y(n_318) );
INVx2_ASAP7_75t_L g319 ( .A(n_290), .Y(n_319) );
INVx2_ASAP7_75t_L g320 ( .A(n_309), .Y(n_320) );
HB1xp67_ASAP7_75t_L g321 ( .A(n_290), .Y(n_321) );
INVx4_ASAP7_75t_L g322 ( .A(n_288), .Y(n_322) );
AO21x2_ASAP7_75t_L g323 ( .A1(n_298), .A2(n_286), .B(n_266), .Y(n_323) );
INVx1_ASAP7_75t_L g324 ( .A(n_293), .Y(n_324) );
INVx2_ASAP7_75t_SL g325 ( .A(n_292), .Y(n_325) );
CKINVDCx5p33_ASAP7_75t_R g326 ( .A(n_297), .Y(n_326) );
BUFx2_ASAP7_75t_L g327 ( .A(n_292), .Y(n_327) );
OA211x2_ASAP7_75t_L g328 ( .A1(n_300), .A2(n_272), .B(n_266), .C(n_283), .Y(n_328) );
AOI33xp33_ASAP7_75t_L g329 ( .A1(n_294), .A2(n_276), .A3(n_280), .B1(n_9), .B2(n_10), .B3(n_11), .Y(n_329) );
AND2x2_ASAP7_75t_L g330 ( .A(n_292), .B(n_273), .Y(n_330) );
AND2x2_ASAP7_75t_L g331 ( .A(n_287), .B(n_259), .Y(n_331) );
AND2x2_ASAP7_75t_L g332 ( .A(n_287), .B(n_262), .Y(n_332) );
AND4x1_ASAP7_75t_L g333 ( .A(n_301), .B(n_264), .C(n_278), .D(n_12), .Y(n_333) );
HB1xp67_ASAP7_75t_L g334 ( .A(n_288), .Y(n_334) );
AND2x2_ASAP7_75t_L g335 ( .A(n_309), .B(n_262), .Y(n_335) );
AND2x2_ASAP7_75t_L g336 ( .A(n_309), .B(n_264), .Y(n_336) );
NAND4xp25_ASAP7_75t_L g337 ( .A(n_294), .B(n_285), .C(n_281), .D(n_250), .Y(n_337) );
INVx4_ASAP7_75t_L g338 ( .A(n_288), .Y(n_338) );
BUFx3_ASAP7_75t_L g339 ( .A(n_297), .Y(n_339) );
INVxp67_ASAP7_75t_SL g340 ( .A(n_288), .Y(n_340) );
INVx4_ASAP7_75t_L g341 ( .A(n_289), .Y(n_341) );
AND2x2_ASAP7_75t_L g342 ( .A(n_310), .B(n_302), .Y(n_342) );
INVx1_ASAP7_75t_L g343 ( .A(n_313), .Y(n_343) );
AND2x2_ASAP7_75t_L g344 ( .A(n_310), .B(n_302), .Y(n_344) );
INVx1_ASAP7_75t_L g345 ( .A(n_313), .Y(n_345) );
INVx2_ASAP7_75t_L g346 ( .A(n_325), .Y(n_346) );
INVx1_ASAP7_75t_L g347 ( .A(n_316), .Y(n_347) );
NOR3xp33_ASAP7_75t_L g348 ( .A(n_329), .B(n_301), .C(n_250), .Y(n_348) );
INVx1_ASAP7_75t_L g349 ( .A(n_316), .Y(n_349) );
INVx1_ASAP7_75t_L g350 ( .A(n_324), .Y(n_350) );
NAND2xp5_ASAP7_75t_SL g351 ( .A(n_318), .B(n_299), .Y(n_351) );
AND2x2_ASAP7_75t_L g352 ( .A(n_310), .B(n_304), .Y(n_352) );
NAND2xp5_ASAP7_75t_L g353 ( .A(n_336), .B(n_299), .Y(n_353) );
OR2x2_ASAP7_75t_L g354 ( .A(n_334), .B(n_304), .Y(n_354) );
AND2x2_ASAP7_75t_L g355 ( .A(n_325), .B(n_327), .Y(n_355) );
INVx1_ASAP7_75t_L g356 ( .A(n_324), .Y(n_356) );
AOI22xp5_ASAP7_75t_L g357 ( .A1(n_328), .A2(n_337), .B1(n_336), .B2(n_318), .Y(n_357) );
INVx1_ASAP7_75t_SL g358 ( .A(n_326), .Y(n_358) );
AND2x2_ASAP7_75t_L g359 ( .A(n_325), .B(n_289), .Y(n_359) );
AND2x2_ASAP7_75t_L g360 ( .A(n_327), .B(n_311), .Y(n_360) );
NAND2xp5_ASAP7_75t_L g361 ( .A(n_336), .B(n_306), .Y(n_361) );
INVx1_ASAP7_75t_L g362 ( .A(n_321), .Y(n_362) );
INVx2_ASAP7_75t_L g363 ( .A(n_327), .Y(n_363) );
HB1xp67_ASAP7_75t_L g364 ( .A(n_312), .Y(n_364) );
INVx1_ASAP7_75t_L g365 ( .A(n_321), .Y(n_365) );
INVx1_ASAP7_75t_SL g366 ( .A(n_334), .Y(n_366) );
INVx1_ASAP7_75t_L g367 ( .A(n_312), .Y(n_367) );
AND2x2_ASAP7_75t_L g368 ( .A(n_311), .B(n_289), .Y(n_368) );
NAND2xp5_ASAP7_75t_L g369 ( .A(n_340), .B(n_306), .Y(n_369) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_340), .B(n_296), .Y(n_370) );
INVx1_ASAP7_75t_L g371 ( .A(n_312), .Y(n_371) );
INVx6_ASAP7_75t_L g372 ( .A(n_322), .Y(n_372) );
AND2x4_ASAP7_75t_L g373 ( .A(n_322), .B(n_295), .Y(n_373) );
BUFx3_ASAP7_75t_L g374 ( .A(n_339), .Y(n_374) );
OR2x2_ASAP7_75t_L g375 ( .A(n_314), .B(n_307), .Y(n_375) );
AND2x2_ASAP7_75t_L g376 ( .A(n_311), .B(n_289), .Y(n_376) );
OR2x2_ASAP7_75t_L g377 ( .A(n_314), .B(n_307), .Y(n_377) );
AND2x2_ASAP7_75t_L g378 ( .A(n_331), .B(n_295), .Y(n_378) );
OR2x2_ASAP7_75t_L g379 ( .A(n_314), .B(n_303), .Y(n_379) );
NAND2xp5_ASAP7_75t_SL g380 ( .A(n_329), .B(n_300), .Y(n_380) );
OR2x2_ASAP7_75t_L g381 ( .A(n_322), .B(n_303), .Y(n_381) );
INVx1_ASAP7_75t_L g382 ( .A(n_319), .Y(n_382) );
AND2x4_ASAP7_75t_L g383 ( .A(n_322), .B(n_295), .Y(n_383) );
INVx2_ASAP7_75t_L g384 ( .A(n_320), .Y(n_384) );
AND2x4_ASAP7_75t_L g385 ( .A(n_322), .B(n_295), .Y(n_385) );
AND2x2_ASAP7_75t_L g386 ( .A(n_331), .B(n_291), .Y(n_386) );
AND2x4_ASAP7_75t_L g387 ( .A(n_338), .B(n_296), .Y(n_387) );
AND2x4_ASAP7_75t_SL g388 ( .A(n_338), .B(n_291), .Y(n_388) );
NAND2xp5_ASAP7_75t_L g389 ( .A(n_342), .B(n_331), .Y(n_389) );
NAND2xp5_ASAP7_75t_L g390 ( .A(n_342), .B(n_332), .Y(n_390) );
INVxp67_ASAP7_75t_SL g391 ( .A(n_364), .Y(n_391) );
XNOR2xp5_ASAP7_75t_L g392 ( .A(n_358), .B(n_333), .Y(n_392) );
OAI22xp5_ASAP7_75t_L g393 ( .A1(n_351), .A2(n_317), .B1(n_338), .B2(n_328), .Y(n_393) );
NAND2xp5_ASAP7_75t_L g394 ( .A(n_344), .B(n_353), .Y(n_394) );
NAND2xp5_ASAP7_75t_L g395 ( .A(n_344), .B(n_332), .Y(n_395) );
OR2x2_ASAP7_75t_L g396 ( .A(n_386), .B(n_338), .Y(n_396) );
INVx1_ASAP7_75t_SL g397 ( .A(n_388), .Y(n_397) );
INVx2_ASAP7_75t_L g398 ( .A(n_384), .Y(n_398) );
INVx1_ASAP7_75t_L g399 ( .A(n_345), .Y(n_399) );
OR2x2_ASAP7_75t_L g400 ( .A(n_386), .B(n_338), .Y(n_400) );
AND2x4_ASAP7_75t_L g401 ( .A(n_388), .B(n_317), .Y(n_401) );
NAND3xp33_ASAP7_75t_SL g402 ( .A(n_348), .B(n_333), .C(n_332), .Y(n_402) );
INVxp67_ASAP7_75t_L g403 ( .A(n_379), .Y(n_403) );
NAND2xp5_ASAP7_75t_L g404 ( .A(n_361), .B(n_319), .Y(n_404) );
NOR2xp33_ASAP7_75t_L g405 ( .A(n_357), .B(n_7), .Y(n_405) );
OR2x2_ASAP7_75t_L g406 ( .A(n_370), .B(n_319), .Y(n_406) );
AND2x2_ASAP7_75t_L g407 ( .A(n_378), .B(n_341), .Y(n_407) );
NAND4xp25_ASAP7_75t_L g408 ( .A(n_380), .B(n_337), .C(n_339), .D(n_341), .Y(n_408) );
AND2x2_ASAP7_75t_L g409 ( .A(n_378), .B(n_341), .Y(n_409) );
OR2x2_ASAP7_75t_L g410 ( .A(n_379), .B(n_341), .Y(n_410) );
AND2x2_ASAP7_75t_L g411 ( .A(n_368), .B(n_341), .Y(n_411) );
NAND2x1_ASAP7_75t_L g412 ( .A(n_372), .B(n_320), .Y(n_412) );
INVx1_ASAP7_75t_L g413 ( .A(n_345), .Y(n_413) );
INVx1_ASAP7_75t_L g414 ( .A(n_347), .Y(n_414) );
INVx1_ASAP7_75t_SL g415 ( .A(n_372), .Y(n_415) );
AND2x2_ASAP7_75t_L g416 ( .A(n_368), .B(n_339), .Y(n_416) );
AND2x2_ASAP7_75t_L g417 ( .A(n_376), .B(n_339), .Y(n_417) );
INVx1_ASAP7_75t_SL g418 ( .A(n_372), .Y(n_418) );
AND2x2_ASAP7_75t_L g419 ( .A(n_376), .B(n_330), .Y(n_419) );
OR2x2_ASAP7_75t_L g420 ( .A(n_381), .B(n_320), .Y(n_420) );
AND2x2_ASAP7_75t_L g421 ( .A(n_387), .B(n_330), .Y(n_421) );
AND2x4_ASAP7_75t_L g422 ( .A(n_387), .B(n_330), .Y(n_422) );
INVx1_ASAP7_75t_L g423 ( .A(n_347), .Y(n_423) );
AND2x2_ASAP7_75t_L g424 ( .A(n_387), .B(n_315), .Y(n_424) );
OAI22xp5_ASAP7_75t_L g425 ( .A1(n_381), .A2(n_320), .B1(n_315), .B2(n_335), .Y(n_425) );
AND2x4_ASAP7_75t_L g426 ( .A(n_374), .B(n_315), .Y(n_426) );
AOI21xp5_ASAP7_75t_L g427 ( .A1(n_369), .A2(n_323), .B(n_335), .Y(n_427) );
INVx1_ASAP7_75t_L g428 ( .A(n_356), .Y(n_428) );
NAND2xp5_ASAP7_75t_L g429 ( .A(n_356), .B(n_323), .Y(n_429) );
AND2x2_ASAP7_75t_L g430 ( .A(n_352), .B(n_335), .Y(n_430) );
OR2x2_ASAP7_75t_L g431 ( .A(n_360), .B(n_323), .Y(n_431) );
AND2x2_ASAP7_75t_L g432 ( .A(n_352), .B(n_323), .Y(n_432) );
INVx1_ASAP7_75t_L g433 ( .A(n_343), .Y(n_433) );
AND2x2_ASAP7_75t_L g434 ( .A(n_360), .B(n_323), .Y(n_434) );
INVxp67_ASAP7_75t_L g435 ( .A(n_374), .Y(n_435) );
AND2x2_ASAP7_75t_L g436 ( .A(n_359), .B(n_8), .Y(n_436) );
OR2x2_ASAP7_75t_L g437 ( .A(n_375), .B(n_12), .Y(n_437) );
INVxp67_ASAP7_75t_L g438 ( .A(n_367), .Y(n_438) );
AND2x4_ASAP7_75t_L g439 ( .A(n_373), .B(n_281), .Y(n_439) );
NAND2xp5_ASAP7_75t_L g440 ( .A(n_349), .B(n_13), .Y(n_440) );
INVx1_ASAP7_75t_L g441 ( .A(n_350), .Y(n_441) );
AOI221xp5_ASAP7_75t_L g442 ( .A1(n_402), .A2(n_371), .B1(n_366), .B2(n_365), .C(n_362), .Y(n_442) );
AOI221xp5_ASAP7_75t_L g443 ( .A1(n_405), .A2(n_362), .B1(n_365), .B2(n_355), .C(n_377), .Y(n_443) );
INVx1_ASAP7_75t_L g444 ( .A(n_433), .Y(n_444) );
INVx2_ASAP7_75t_L g445 ( .A(n_420), .Y(n_445) );
INVx2_ASAP7_75t_L g446 ( .A(n_396), .Y(n_446) );
A2O1A1Ixp33_ASAP7_75t_L g447 ( .A1(n_408), .A2(n_385), .B(n_383), .C(n_373), .Y(n_447) );
AOI22xp5_ASAP7_75t_L g448 ( .A1(n_393), .A2(n_372), .B1(n_385), .B2(n_383), .Y(n_448) );
INVx1_ASAP7_75t_SL g449 ( .A(n_397), .Y(n_449) );
AO22x1_ASAP7_75t_L g450 ( .A1(n_401), .A2(n_385), .B1(n_383), .B2(n_373), .Y(n_450) );
AND2x2_ASAP7_75t_L g451 ( .A(n_421), .B(n_359), .Y(n_451) );
NOR3xp33_ASAP7_75t_L g452 ( .A(n_440), .B(n_250), .C(n_281), .Y(n_452) );
OR2x2_ASAP7_75t_L g453 ( .A(n_389), .B(n_377), .Y(n_453) );
OAI322xp33_ASAP7_75t_L g454 ( .A1(n_431), .A2(n_375), .A3(n_354), .B1(n_363), .B2(n_346), .C1(n_355), .C2(n_382), .Y(n_454) );
NAND2xp5_ASAP7_75t_L g455 ( .A(n_403), .B(n_363), .Y(n_455) );
NAND2xp5_ASAP7_75t_L g456 ( .A(n_394), .B(n_346), .Y(n_456) );
OR2x2_ASAP7_75t_L g457 ( .A(n_389), .B(n_354), .Y(n_457) );
AOI22xp33_ASAP7_75t_SL g458 ( .A1(n_401), .A2(n_384), .B1(n_241), .B2(n_246), .Y(n_458) );
INVx1_ASAP7_75t_L g459 ( .A(n_441), .Y(n_459) );
NOR2xp33_ASAP7_75t_L g460 ( .A(n_392), .B(n_14), .Y(n_460) );
AND2x2_ASAP7_75t_L g461 ( .A(n_424), .B(n_422), .Y(n_461) );
AOI221xp5_ASAP7_75t_L g462 ( .A1(n_434), .A2(n_135), .B1(n_246), .B2(n_16), .C(n_17), .Y(n_462) );
NAND2xp5_ASAP7_75t_SL g463 ( .A(n_397), .B(n_258), .Y(n_463) );
OAI32xp33_ASAP7_75t_L g464 ( .A1(n_400), .A2(n_260), .A3(n_15), .B1(n_16), .B2(n_14), .Y(n_464) );
NAND2xp5_ASAP7_75t_L g465 ( .A(n_394), .B(n_135), .Y(n_465) );
OAI21xp5_ASAP7_75t_L g466 ( .A1(n_393), .A2(n_248), .B(n_236), .Y(n_466) );
OAI21xp5_ASAP7_75t_L g467 ( .A1(n_437), .A2(n_248), .B(n_236), .Y(n_467) );
OAI22xp33_ASAP7_75t_SL g468 ( .A1(n_412), .A2(n_241), .B1(n_22), .B2(n_23), .Y(n_468) );
NAND2xp5_ASAP7_75t_SL g469 ( .A(n_415), .B(n_258), .Y(n_469) );
OR2x2_ASAP7_75t_L g470 ( .A(n_390), .B(n_258), .Y(n_470) );
OAI31xp33_ASAP7_75t_L g471 ( .A1(n_415), .A2(n_241), .A3(n_24), .B(n_27), .Y(n_471) );
OAI21xp33_ASAP7_75t_L g472 ( .A1(n_432), .A2(n_147), .B(n_146), .Y(n_472) );
AND2x2_ASAP7_75t_L g473 ( .A(n_422), .B(n_258), .Y(n_473) );
OAI21xp33_ASAP7_75t_SL g474 ( .A1(n_418), .A2(n_19), .B(n_28), .Y(n_474) );
INVxp67_ASAP7_75t_L g475 ( .A(n_391), .Y(n_475) );
NAND2x1_ASAP7_75t_L g476 ( .A(n_426), .B(n_258), .Y(n_476) );
INVx1_ASAP7_75t_L g477 ( .A(n_399), .Y(n_477) );
INVx1_ASAP7_75t_L g478 ( .A(n_413), .Y(n_478) );
OAI221xp5_ASAP7_75t_L g479 ( .A1(n_435), .A2(n_147), .B1(n_146), .B2(n_143), .C(n_199), .Y(n_479) );
HB1xp67_ASAP7_75t_L g480 ( .A(n_426), .Y(n_480) );
OAI21xp5_ASAP7_75t_SL g481 ( .A1(n_418), .A2(n_147), .B(n_146), .Y(n_481) );
NOR2xp33_ASAP7_75t_L g482 ( .A(n_390), .B(n_29), .Y(n_482) );
AND2x2_ASAP7_75t_L g483 ( .A(n_416), .B(n_30), .Y(n_483) );
OAI22xp5_ASAP7_75t_L g484 ( .A1(n_410), .A2(n_425), .B1(n_395), .B2(n_436), .Y(n_484) );
NAND2xp5_ASAP7_75t_L g485 ( .A(n_395), .B(n_31), .Y(n_485) );
NOR4xp25_ASAP7_75t_L g486 ( .A(n_440), .B(n_33), .C(n_38), .D(n_39), .Y(n_486) );
AND2x2_ASAP7_75t_L g487 ( .A(n_480), .B(n_430), .Y(n_487) );
INVx1_ASAP7_75t_L g488 ( .A(n_456), .Y(n_488) );
INVx2_ASAP7_75t_L g489 ( .A(n_477), .Y(n_489) );
OAI21xp33_ASAP7_75t_L g490 ( .A1(n_460), .A2(n_427), .B(n_429), .Y(n_490) );
NAND2xp5_ASAP7_75t_SL g491 ( .A(n_442), .B(n_425), .Y(n_491) );
INVx1_ASAP7_75t_L g492 ( .A(n_444), .Y(n_492) );
NAND2xp33_ASAP7_75t_L g493 ( .A(n_447), .B(n_411), .Y(n_493) );
CKINVDCx14_ASAP7_75t_R g494 ( .A(n_448), .Y(n_494) );
INVx1_ASAP7_75t_L g495 ( .A(n_459), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_484), .B(n_438), .Y(n_496) );
AOI222xp33_ASAP7_75t_L g497 ( .A1(n_443), .A2(n_429), .B1(n_404), .B2(n_428), .C1(n_423), .C2(n_414), .Y(n_497) );
NAND2xp5_ASAP7_75t_L g498 ( .A(n_475), .B(n_419), .Y(n_498) );
INVx1_ASAP7_75t_L g499 ( .A(n_457), .Y(n_499) );
AOI22xp33_ASAP7_75t_L g500 ( .A1(n_452), .A2(n_439), .B1(n_417), .B2(n_409), .Y(n_500) );
INVx1_ASAP7_75t_L g501 ( .A(n_478), .Y(n_501) );
AOI32xp33_ASAP7_75t_L g502 ( .A1(n_449), .A2(n_407), .A3(n_439), .B1(n_404), .B2(n_406), .Y(n_502) );
AOI31xp33_ASAP7_75t_L g503 ( .A1(n_442), .A2(n_398), .A3(n_43), .B(n_44), .Y(n_503) );
OR2x2_ASAP7_75t_L g504 ( .A(n_453), .B(n_40), .Y(n_504) );
OAI211xp5_ASAP7_75t_L g505 ( .A1(n_443), .A2(n_147), .B(n_146), .C(n_143), .Y(n_505) );
OAI21xp5_ASAP7_75t_SL g506 ( .A1(n_458), .A2(n_147), .B(n_146), .Y(n_506) );
INVx1_ASAP7_75t_L g507 ( .A(n_455), .Y(n_507) );
INVx1_ASAP7_75t_L g508 ( .A(n_475), .Y(n_508) );
INVx2_ASAP7_75t_L g509 ( .A(n_470), .Y(n_509) );
AOI22xp5_ASAP7_75t_L g510 ( .A1(n_450), .A2(n_143), .B1(n_199), .B2(n_48), .Y(n_510) );
XNOR2xp5_ASAP7_75t_L g511 ( .A(n_461), .B(n_45), .Y(n_511) );
AOI221xp5_ASAP7_75t_L g512 ( .A1(n_454), .A2(n_46), .B1(n_49), .B2(n_50), .C(n_51), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_446), .B(n_52), .Y(n_513) );
NOR2xp33_ASAP7_75t_L g514 ( .A(n_451), .B(n_465), .Y(n_514) );
INVx1_ASAP7_75t_SL g515 ( .A(n_483), .Y(n_515) );
INVx2_ASAP7_75t_L g516 ( .A(n_445), .Y(n_516) );
OAI21xp33_ASAP7_75t_L g517 ( .A1(n_490), .A2(n_466), .B(n_458), .Y(n_517) );
OAI21xp5_ASAP7_75t_L g518 ( .A1(n_491), .A2(n_474), .B(n_486), .Y(n_518) );
AOI22xp5_ASAP7_75t_L g519 ( .A1(n_494), .A2(n_452), .B1(n_462), .B2(n_482), .Y(n_519) );
AOI211xp5_ASAP7_75t_SL g520 ( .A1(n_503), .A2(n_468), .B(n_462), .C(n_481), .Y(n_520) );
AOI21xp5_ASAP7_75t_L g521 ( .A1(n_491), .A2(n_471), .B(n_476), .Y(n_521) );
OAI221xp5_ASAP7_75t_L g522 ( .A1(n_500), .A2(n_467), .B1(n_485), .B2(n_472), .C(n_463), .Y(n_522) );
INVxp67_ASAP7_75t_L g523 ( .A(n_508), .Y(n_523) );
OAI22xp33_ASAP7_75t_L g524 ( .A1(n_496), .A2(n_469), .B1(n_473), .B2(n_479), .Y(n_524) );
INVxp67_ASAP7_75t_SL g525 ( .A(n_505), .Y(n_525) );
AOI221xp5_ASAP7_75t_L g526 ( .A1(n_494), .A2(n_464), .B1(n_55), .B2(n_56), .C(n_57), .Y(n_526) );
INVx1_ASAP7_75t_L g527 ( .A(n_489), .Y(n_527) );
AND2x4_ASAP7_75t_L g528 ( .A(n_507), .B(n_54), .Y(n_528) );
O2A1O1Ixp33_ASAP7_75t_L g529 ( .A1(n_506), .A2(n_59), .B(n_60), .C(n_61), .Y(n_529) );
AND2x2_ASAP7_75t_L g530 ( .A(n_509), .B(n_63), .Y(n_530) );
OAI21xp5_ASAP7_75t_SL g531 ( .A1(n_511), .A2(n_76), .B(n_69), .Y(n_531) );
INVx1_ASAP7_75t_L g532 ( .A(n_489), .Y(n_532) );
O2A1O1Ixp33_ASAP7_75t_L g533 ( .A1(n_493), .A2(n_67), .B(n_70), .C(n_71), .Y(n_533) );
AOI222xp33_ASAP7_75t_L g534 ( .A1(n_518), .A2(n_500), .B1(n_492), .B2(n_495), .C1(n_488), .C2(n_512), .Y(n_534) );
INVx1_ASAP7_75t_SL g535 ( .A(n_528), .Y(n_535) );
AND2x2_ASAP7_75t_L g536 ( .A(n_523), .B(n_509), .Y(n_536) );
INVx2_ASAP7_75t_L g537 ( .A(n_527), .Y(n_537) );
AOI221xp5_ASAP7_75t_SL g538 ( .A1(n_521), .A2(n_515), .B1(n_514), .B2(n_498), .C(n_499), .Y(n_538) );
INVx1_ASAP7_75t_L g539 ( .A(n_532), .Y(n_539) );
AOI211xp5_ASAP7_75t_L g540 ( .A1(n_517), .A2(n_504), .B(n_510), .C(n_514), .Y(n_540) );
NAND4xp25_ASAP7_75t_SL g541 ( .A(n_519), .B(n_502), .C(n_497), .D(n_487), .Y(n_541) );
OAI221xp5_ASAP7_75t_SL g542 ( .A1(n_525), .A2(n_501), .B1(n_513), .B2(n_516), .C(n_526), .Y(n_542) );
BUFx2_ASAP7_75t_L g543 ( .A(n_535), .Y(n_543) );
NOR2x1_ASAP7_75t_L g544 ( .A(n_541), .B(n_533), .Y(n_544) );
NAND3xp33_ASAP7_75t_SL g545 ( .A(n_534), .B(n_520), .C(n_531), .Y(n_545) );
OR2x2_ASAP7_75t_L g546 ( .A(n_539), .B(n_524), .Y(n_546) );
NOR2xp33_ASAP7_75t_L g547 ( .A(n_542), .B(n_522), .Y(n_547) );
AOI22xp5_ASAP7_75t_L g548 ( .A1(n_545), .A2(n_538), .B1(n_540), .B2(n_536), .Y(n_548) );
AND2x2_ASAP7_75t_L g549 ( .A(n_543), .B(n_536), .Y(n_549) );
BUFx2_ASAP7_75t_L g550 ( .A(n_544), .Y(n_550) );
INVx1_ASAP7_75t_L g551 ( .A(n_549), .Y(n_551) );
INVx1_ASAP7_75t_L g552 ( .A(n_550), .Y(n_552) );
INVx1_ASAP7_75t_L g553 ( .A(n_551), .Y(n_553) );
INVx1_ASAP7_75t_L g554 ( .A(n_553), .Y(n_554) );
AOI222xp33_ASAP7_75t_SL g555 ( .A1(n_554), .A2(n_552), .B1(n_548), .B2(n_547), .C1(n_546), .C2(n_537), .Y(n_555) );
OAI21x1_ASAP7_75t_SL g556 ( .A1(n_555), .A2(n_529), .B(n_537), .Y(n_556) );
AOI21xp5_ASAP7_75t_L g557 ( .A1(n_556), .A2(n_528), .B(n_530), .Y(n_557) );
endmodule