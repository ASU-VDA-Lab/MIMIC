module fake_aes_12221_n_19 (n_1, n_2, n_4, n_3, n_5, n_0, n_19);
input n_1;
input n_2;
input n_4;
input n_3;
input n_5;
input n_0;
output n_19;
wire n_8;
wire n_11;
wire n_16;
wire n_13;
wire n_18;
wire n_12;
wire n_9;
wire n_17;
wire n_14;
wire n_10;
wire n_15;
wire n_6;
wire n_7;
INVx2_ASAP7_75t_L g6 ( .A(n_5), .Y(n_6) );
BUFx3_ASAP7_75t_L g7 ( .A(n_5), .Y(n_7) );
INVx2_ASAP7_75t_L g8 ( .A(n_1), .Y(n_8) );
NAND2xp5_ASAP7_75t_SL g9 ( .A(n_2), .B(n_4), .Y(n_9) );
INVx2_ASAP7_75t_L g10 ( .A(n_0), .Y(n_10) );
OAI21x1_ASAP7_75t_L g11 ( .A1(n_8), .A2(n_0), .B(n_1), .Y(n_11) );
O2A1O1Ixp33_ASAP7_75t_SL g12 ( .A1(n_9), .A2(n_0), .B(n_1), .C(n_2), .Y(n_12) );
OAI21x1_ASAP7_75t_L g13 ( .A1(n_10), .A2(n_2), .B(n_3), .Y(n_13) );
NAND2xp5_ASAP7_75t_L g14 ( .A(n_11), .B(n_7), .Y(n_14) );
NAND2xp5_ASAP7_75t_L g15 ( .A(n_14), .B(n_13), .Y(n_15) );
OAI211xp5_ASAP7_75t_SL g16 ( .A1(n_15), .A2(n_9), .B(n_12), .C(n_6), .Y(n_16) );
AND3x4_ASAP7_75t_L g17 ( .A(n_16), .B(n_3), .C(n_4), .Y(n_17) );
CKINVDCx20_ASAP7_75t_R g18 ( .A(n_17), .Y(n_18) );
INVx3_ASAP7_75t_L g19 ( .A(n_18), .Y(n_19) );
endmodule