module fake_jpeg_28322_n_195 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_195);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_195;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx16f_ASAP7_75t_L g16 ( 
.A(n_14),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_8),
.Y(n_17)
);

INVx11_ASAP7_75t_SL g18 ( 
.A(n_11),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_5),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_13),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_11),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_3),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

INVx11_ASAP7_75t_SL g26 ( 
.A(n_8),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_1),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_4),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_25),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_33),
.Y(n_45)
);

INVx11_ASAP7_75t_L g34 ( 
.A(n_26),
.Y(n_34)
);

INVx5_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_22),
.B(n_0),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_35),
.B(n_25),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_22),
.Y(n_36)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_22),
.Y(n_37)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_38),
.B(n_39),
.Y(n_53)
);

CKINVDCx16_ASAP7_75t_R g39 ( 
.A(n_26),
.Y(n_39)
);

INVx2_ASAP7_75t_SL g40 ( 
.A(n_18),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_40),
.B(n_42),
.Y(n_55)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

INVx5_ASAP7_75t_L g42 ( 
.A(n_16),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_18),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_43),
.B(n_28),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g44 ( 
.A1(n_35),
.A2(n_29),
.B1(n_32),
.B2(n_19),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_44),
.A2(n_17),
.B1(n_24),
.B2(n_30),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g46 ( 
.A(n_35),
.B(n_17),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g69 ( 
.A(n_46),
.B(n_61),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_38),
.A2(n_29),
.B1(n_32),
.B2(n_19),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_49),
.A2(n_40),
.B1(n_31),
.B2(n_23),
.Y(n_83)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_41),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_51),
.B(n_63),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_52),
.B(n_57),
.Y(n_68)
);

INVx11_ASAP7_75t_L g54 ( 
.A(n_33),
.Y(n_54)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_54),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_36),
.B(n_30),
.Y(n_57)
);

BUFx5_ASAP7_75t_L g58 ( 
.A(n_33),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_58),
.B(n_60),
.Y(n_75)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_59),
.Y(n_78)
);

BUFx5_ASAP7_75t_L g60 ( 
.A(n_33),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_36),
.B(n_31),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_36),
.B(n_24),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_SL g79 ( 
.A(n_62),
.B(n_27),
.Y(n_79)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_41),
.Y(n_63)
);

OAI21xp33_ASAP7_75t_L g65 ( 
.A1(n_46),
.A2(n_42),
.B(n_38),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_65),
.A2(n_23),
.B1(n_40),
.B2(n_27),
.Y(n_87)
);

XOR2xp5_ASAP7_75t_L g66 ( 
.A(n_52),
.B(n_37),
.Y(n_66)
);

XOR2xp5_ASAP7_75t_L g95 ( 
.A(n_66),
.B(n_73),
.Y(n_95)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_54),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_67),
.B(n_71),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_L g70 ( 
.A1(n_57),
.A2(n_42),
.B1(n_37),
.B2(n_25),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_70),
.A2(n_74),
.B1(n_83),
.B2(n_34),
.Y(n_97)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_54),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_44),
.B(n_37),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g105 ( 
.A(n_72),
.B(n_79),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_61),
.B(n_33),
.C(n_25),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_50),
.A2(n_40),
.B1(n_34),
.B2(n_39),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_77),
.A2(n_48),
.B1(n_59),
.B2(n_55),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_62),
.B(n_20),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_80),
.B(n_81),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_55),
.Y(n_81)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_50),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_82),
.B(n_45),
.Y(n_94)
);

AND2x2_ASAP7_75t_SL g84 ( 
.A(n_63),
.B(n_43),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_84),
.B(n_45),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_75),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_85),
.B(n_87),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_L g111 ( 
.A1(n_86),
.A2(n_93),
.B(n_99),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_64),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_88),
.B(n_101),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_90),
.A2(n_97),
.B1(n_86),
.B2(n_88),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_66),
.B(n_48),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_92),
.B(n_96),
.Y(n_116)
);

AOI32xp33_ASAP7_75t_L g93 ( 
.A1(n_81),
.A2(n_53),
.A3(n_16),
.B1(n_56),
.B2(n_21),
.Y(n_93)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_94),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_68),
.B(n_51),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_68),
.B(n_53),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_98),
.B(n_100),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_L g99 ( 
.A1(n_72),
.A2(n_78),
.B(n_69),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_69),
.B(n_45),
.Y(n_100)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_64),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_78),
.B(n_45),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_102),
.B(n_104),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_79),
.B(n_21),
.Y(n_103)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_103),
.Y(n_122)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_77),
.Y(n_104)
);

O2A1O1Ixp33_ASAP7_75t_SL g106 ( 
.A1(n_104),
.A2(n_84),
.B(n_74),
.C(n_73),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_L g127 ( 
.A1(n_106),
.A2(n_86),
.B(n_105),
.Y(n_127)
);

XOR2xp5_ASAP7_75t_L g107 ( 
.A(n_95),
.B(n_84),
.Y(n_107)
);

XOR2xp5_ASAP7_75t_L g138 ( 
.A(n_107),
.B(n_109),
.Y(n_138)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_89),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_108),
.B(n_112),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_95),
.B(n_84),
.C(n_82),
.Y(n_109)
);

INVx5_ASAP7_75t_SL g112 ( 
.A(n_85),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_114),
.A2(n_93),
.B1(n_56),
.B2(n_67),
.Y(n_134)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_102),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_115),
.B(n_117),
.Y(n_129)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_96),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_92),
.B(n_76),
.C(n_71),
.Y(n_120)
);

XOR2xp5_ASAP7_75t_L g141 ( 
.A(n_120),
.B(n_121),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_SL g121 ( 
.A(n_98),
.B(n_16),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_99),
.B(n_76),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_124),
.B(n_87),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_114),
.A2(n_101),
.B1(n_100),
.B2(n_90),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_125),
.A2(n_134),
.B1(n_47),
.B2(n_43),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_122),
.B(n_91),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_126),
.B(n_128),
.Y(n_152)
);

XOR2xp5_ASAP7_75t_L g142 ( 
.A(n_127),
.B(n_124),
.Y(n_142)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_123),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_119),
.B(n_105),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_130),
.B(n_133),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_106),
.A2(n_115),
.B1(n_117),
.B2(n_113),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_132),
.A2(n_118),
.B1(n_116),
.B2(n_109),
.Y(n_143)
);

CKINVDCx16_ASAP7_75t_R g135 ( 
.A(n_123),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_135),
.B(n_137),
.Y(n_154)
);

AOI21xp33_ASAP7_75t_L g136 ( 
.A1(n_111),
.A2(n_20),
.B(n_12),
.Y(n_136)
);

AOI221xp5_ASAP7_75t_L g151 ( 
.A1(n_136),
.A2(n_140),
.B1(n_14),
.B2(n_12),
.C(n_2),
.Y(n_151)
);

INVxp67_ASAP7_75t_L g137 ( 
.A(n_120),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g139 ( 
.A(n_118),
.B(n_15),
.Y(n_139)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_139),
.Y(n_145)
);

A2O1A1O1Ixp25_ASAP7_75t_L g140 ( 
.A1(n_111),
.A2(n_28),
.B(n_58),
.C(n_60),
.D(n_15),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_142),
.B(n_146),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_SL g159 ( 
.A1(n_143),
.A2(n_144),
.B(n_133),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_125),
.A2(n_140),
.B1(n_137),
.B2(n_112),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_138),
.B(n_107),
.C(n_116),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_138),
.B(n_121),
.C(n_110),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_147),
.B(n_149),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_132),
.A2(n_108),
.B1(n_106),
.B2(n_47),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_148),
.A2(n_150),
.B1(n_151),
.B2(n_153),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_141),
.B(n_43),
.C(n_28),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_128),
.A2(n_47),
.B1(n_1),
.B2(n_2),
.Y(n_153)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_152),
.Y(n_158)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_158),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_159),
.B(n_0),
.Y(n_171)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_154),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_L g174 ( 
.A1(n_160),
.A2(n_162),
.B(n_165),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_155),
.B(n_129),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_161),
.B(n_164),
.Y(n_170)
);

AOI21xp5_ASAP7_75t_L g162 ( 
.A1(n_142),
.A2(n_127),
.B(n_131),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_144),
.B(n_130),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_153),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_SL g166 ( 
.A(n_145),
.B(n_141),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_166),
.B(n_146),
.C(n_147),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_167),
.B(n_169),
.Y(n_175)
);

BUFx4f_ASAP7_75t_SL g168 ( 
.A(n_157),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_168),
.B(n_173),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_156),
.B(n_149),
.C(n_150),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_171),
.B(n_161),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g173 ( 
.A(n_163),
.B(n_1),
.Y(n_173)
);

AOI21xp5_ASAP7_75t_L g177 ( 
.A1(n_172),
.A2(n_159),
.B(n_164),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_177),
.B(n_181),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_178),
.A2(n_173),
.B1(n_168),
.B2(n_5),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_170),
.B(n_162),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_179),
.B(n_180),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_174),
.B(n_156),
.Y(n_180)
);

AOI21xp5_ASAP7_75t_L g181 ( 
.A1(n_171),
.A2(n_163),
.B(n_3),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_183),
.B(n_7),
.Y(n_188)
);

OAI221xp5_ASAP7_75t_L g185 ( 
.A1(n_175),
.A2(n_168),
.B1(n_3),
.B2(n_5),
.C(n_6),
.Y(n_185)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_185),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_176),
.B(n_2),
.C(n_6),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_186),
.B(n_184),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_182),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_187)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_187),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_188),
.B(n_190),
.Y(n_191)
);

AOI321xp33_ASAP7_75t_L g193 ( 
.A1(n_192),
.A2(n_189),
.A3(n_184),
.B1(n_186),
.B2(n_9),
.C(n_7),
.Y(n_193)
);

XNOR2x2_ASAP7_75t_SL g195 ( 
.A(n_193),
.B(n_194),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_L g194 ( 
.A1(n_191),
.A2(n_189),
.B(n_9),
.Y(n_194)
);


endmodule