module real_aes_5429_n_8 (n_4, n_0, n_3, n_5, n_2, n_7, n_6, n_1, n_8);
input n_4;
input n_0;
input n_3;
input n_5;
input n_2;
input n_7;
input n_6;
input n_1;
output n_8;
wire n_28;
wire n_17;
wire n_22;
wire n_13;
wire n_24;
wire n_12;
wire n_19;
wire n_25;
wire n_14;
wire n_11;
wire n_16;
wire n_15;
wire n_27;
wire n_23;
wire n_9;
wire n_29;
wire n_20;
wire n_18;
wire n_26;
wire n_21;
wire n_10;
NAND3xp33_ASAP7_75t_SL g22 ( .A(n_0), .B(n_23), .C(n_25), .Y(n_22) );
HB1xp67_ASAP7_75t_L g24 ( .A(n_1), .Y(n_24) );
NAND2xp5_ASAP7_75t_L g17 ( .A(n_2), .B(n_6), .Y(n_17) );
BUFx6f_ASAP7_75t_L g27 ( .A(n_3), .Y(n_27) );
INVx2_ASAP7_75t_SL g12 ( .A(n_4), .Y(n_12) );
INVx1_ASAP7_75t_L g19 ( .A(n_5), .Y(n_19) );
HB1xp67_ASAP7_75t_L g14 ( .A(n_7), .Y(n_14) );
AOI32xp33_ASAP7_75t_L g8 ( .A1(n_9), .A2(n_15), .A3(n_18), .B1(n_20), .B2(n_29), .Y(n_8) );
NOR2xp33_ASAP7_75t_L g9 ( .A(n_10), .B(n_13), .Y(n_9) );
OAI21xp33_ASAP7_75t_SL g20 ( .A1(n_10), .A2(n_15), .B(n_21), .Y(n_20) );
AOI21xp5_ASAP7_75t_L g21 ( .A1(n_10), .A2(n_22), .B(n_28), .Y(n_21) );
NOR2xp33_ASAP7_75t_L g28 ( .A(n_10), .B(n_14), .Y(n_28) );
HB1xp67_ASAP7_75t_L g10 ( .A(n_11), .Y(n_10) );
HB1xp67_ASAP7_75t_L g11 ( .A(n_12), .Y(n_11) );
CKINVDCx5p33_ASAP7_75t_R g13 ( .A(n_14), .Y(n_13) );
CKINVDCx5p33_ASAP7_75t_R g15 ( .A(n_16), .Y(n_15) );
HB1xp67_ASAP7_75t_L g16 ( .A(n_17), .Y(n_16) );
CKINVDCx20_ASAP7_75t_R g29 ( .A(n_18), .Y(n_29) );
HB1xp67_ASAP7_75t_L g18 ( .A(n_19), .Y(n_18) );
INVx1_ASAP7_75t_L g23 ( .A(n_24), .Y(n_23) );
BUFx2_ASAP7_75t_L g25 ( .A(n_26), .Y(n_25) );
HB1xp67_ASAP7_75t_L g26 ( .A(n_27), .Y(n_26) );
endmodule