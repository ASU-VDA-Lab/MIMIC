module fake_jpeg_15687_n_136 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_136);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_136;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

INVx11_ASAP7_75t_SL g41 ( 
.A(n_0),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_30),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_29),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_38),
.B(n_3),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_16),
.Y(n_47)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_27),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_1),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_6),
.Y(n_50)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_25),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_11),
.Y(n_52)
);

BUFx12_ASAP7_75t_L g53 ( 
.A(n_8),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_21),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_31),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_24),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_43),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g72 ( 
.A(n_58),
.B(n_60),
.Y(n_72)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_56),
.Y(n_59)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_59),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_50),
.B(n_0),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_42),
.Y(n_61)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_61),
.Y(n_67)
);

BUFx24_ASAP7_75t_L g62 ( 
.A(n_41),
.Y(n_62)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_62),
.Y(n_68)
);

BUFx16f_ASAP7_75t_L g63 ( 
.A(n_41),
.Y(n_63)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_63),
.Y(n_77)
);

BUFx12_ASAP7_75t_L g64 ( 
.A(n_44),
.Y(n_64)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_64),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_42),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_65),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_63),
.B(n_49),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_66),
.B(n_71),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_65),
.A2(n_51),
.B1(n_48),
.B2(n_57),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_69),
.A2(n_74),
.B1(n_2),
.B2(n_3),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_61),
.A2(n_51),
.B1(n_48),
.B2(n_52),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_L g81 ( 
.A1(n_70),
.A2(n_80),
.B1(n_1),
.B2(n_2),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_64),
.A2(n_55),
.B1(n_53),
.B2(n_47),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_64),
.A2(n_44),
.B1(n_47),
.B2(n_46),
.Y(n_74)
);

OA22x2_ASAP7_75t_L g75 ( 
.A1(n_62),
.A2(n_46),
.B1(n_53),
.B2(n_54),
.Y(n_75)
);

OAI32xp33_ASAP7_75t_L g85 ( 
.A1(n_75),
.A2(n_69),
.A3(n_73),
.B1(n_72),
.B2(n_67),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_62),
.Y(n_79)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_79),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_60),
.A2(n_45),
.B1(n_18),
.B2(n_19),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_81),
.B(n_82),
.Y(n_97)
);

INVxp67_ASAP7_75t_L g82 ( 
.A(n_74),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_84),
.A2(n_85),
.B1(n_5),
.B2(n_6),
.Y(n_103)
);

BUFx3_ASAP7_75t_L g86 ( 
.A(n_76),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_86),
.B(n_87),
.Y(n_102)
);

CKINVDCx16_ASAP7_75t_R g87 ( 
.A(n_79),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_76),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_89),
.B(n_91),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_77),
.B(n_4),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_90),
.B(n_92),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_73),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_75),
.Y(n_92)
);

BUFx3_ASAP7_75t_L g93 ( 
.A(n_78),
.Y(n_93)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_93),
.Y(n_99)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_75),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_94),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_68),
.Y(n_95)
);

INVx13_ASAP7_75t_L g106 ( 
.A(n_95),
.Y(n_106)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_68),
.Y(n_96)
);

INVx13_ASAP7_75t_L g107 ( 
.A(n_96),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_83),
.A2(n_20),
.B1(n_40),
.B2(n_36),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_98),
.A2(n_84),
.B1(n_81),
.B2(n_9),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_L g100 ( 
.A1(n_83),
.A2(n_4),
.B(n_5),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_100),
.B(n_86),
.C(n_8),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_103),
.A2(n_7),
.B1(n_9),
.B2(n_10),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_104),
.B(n_88),
.Y(n_108)
);

XNOR2xp5_ASAP7_75t_L g114 ( 
.A(n_108),
.B(n_109),
.Y(n_114)
);

INVxp33_ASAP7_75t_L g110 ( 
.A(n_105),
.Y(n_110)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_110),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_L g117 ( 
.A1(n_111),
.A2(n_100),
.B(n_101),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_112),
.A2(n_113),
.B1(n_98),
.B2(n_99),
.Y(n_118)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_102),
.Y(n_113)
);

XOR2xp5_ASAP7_75t_L g115 ( 
.A(n_111),
.B(n_97),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g119 ( 
.A(n_115),
.B(n_118),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_117),
.B(n_115),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_120),
.A2(n_121),
.B1(n_107),
.B2(n_93),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_116),
.A2(n_110),
.B1(n_106),
.B2(n_99),
.Y(n_121)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_114),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_122),
.A2(n_7),
.B1(n_12),
.B2(n_13),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_114),
.B(n_106),
.Y(n_123)
);

XNOR2xp5_ASAP7_75t_SL g125 ( 
.A(n_123),
.B(n_107),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_L g127 ( 
.A(n_124),
.B(n_125),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_127),
.B(n_126),
.Y(n_128)
);

AOI21xp5_ASAP7_75t_SL g129 ( 
.A1(n_128),
.A2(n_123),
.B(n_119),
.Y(n_129)
);

AOI21xp5_ASAP7_75t_L g130 ( 
.A1(n_129),
.A2(n_14),
.B(n_15),
.Y(n_130)
);

NOR2xp67_ASAP7_75t_L g131 ( 
.A(n_130),
.B(n_17),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_131),
.A2(n_22),
.B1(n_23),
.B2(n_26),
.Y(n_132)
);

NOR3xp33_ASAP7_75t_L g133 ( 
.A(n_132),
.B(n_28),
.C(n_32),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_L g134 ( 
.A(n_133),
.B(n_34),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_134),
.B(n_35),
.Y(n_135)
);

BUFx24_ASAP7_75t_SL g136 ( 
.A(n_135),
.Y(n_136)
);


endmodule