module fake_jpeg_23333_n_219 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_219);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_219;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_182;
wire n_19;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_207;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

INVx4_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

BUFx12_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_3),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

BUFx8_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

INVx1_ASAP7_75t_SL g28 ( 
.A(n_8),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_10),
.Y(n_29)
);

INVx2_ASAP7_75t_SL g30 ( 
.A(n_10),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_6),
.B(n_14),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_25),
.Y(n_34)
);

INVx11_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_19),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_SL g47 ( 
.A(n_35),
.B(n_37),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g36 ( 
.A(n_33),
.B(n_1),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_36),
.B(n_40),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_19),
.Y(n_37)
);

BUFx12_ASAP7_75t_L g38 ( 
.A(n_25),
.Y(n_38)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_38),
.Y(n_65)
);

INVx5_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

BUFx2_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_28),
.B(n_1),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_25),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_41),
.Y(n_64)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_16),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_42),
.B(n_23),
.Y(n_62)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_17),
.Y(n_43)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_43),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_29),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_SL g59 ( 
.A(n_44),
.B(n_18),
.Y(n_59)
);

MAJIxp5_ASAP7_75t_L g45 ( 
.A(n_28),
.B(n_2),
.C(n_3),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g52 ( 
.A(n_45),
.B(n_2),
.Y(n_52)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_34),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_48),
.B(n_54),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_L g50 ( 
.A1(n_35),
.A2(n_16),
.B1(n_28),
.B2(n_29),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_L g79 ( 
.A1(n_50),
.A2(n_21),
.B1(n_24),
.B2(n_20),
.Y(n_79)
);

AOI21xp5_ASAP7_75t_L g98 ( 
.A1(n_52),
.A2(n_69),
.B(n_24),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_37),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_53),
.Y(n_73)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_45),
.A2(n_16),
.B1(n_23),
.B2(n_18),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_56),
.A2(n_66),
.B1(n_68),
.B2(n_30),
.Y(n_89)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_57),
.B(n_58),
.Y(n_84)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_34),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_59),
.B(n_27),
.Y(n_90)
);

CKINVDCx12_ASAP7_75t_R g60 ( 
.A(n_39),
.Y(n_60)
);

CKINVDCx14_ASAP7_75t_R g87 ( 
.A(n_60),
.Y(n_87)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_40),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_61),
.B(n_23),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_62),
.Y(n_71)
);

A2O1A1Ixp33_ASAP7_75t_L g63 ( 
.A1(n_44),
.A2(n_33),
.B(n_32),
.C(n_31),
.Y(n_63)
);

OAI21xp5_ASAP7_75t_SL g92 ( 
.A1(n_63),
.A2(n_21),
.B(n_22),
.Y(n_92)
);

OAI22xp33_ASAP7_75t_L g66 ( 
.A1(n_42),
.A2(n_30),
.B1(n_31),
.B2(n_32),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_34),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_67),
.Y(n_83)
);

OA22x2_ASAP7_75t_L g68 ( 
.A1(n_41),
.A2(n_30),
.B1(n_31),
.B2(n_32),
.Y(n_68)
);

NAND2x1_ASAP7_75t_SL g69 ( 
.A(n_45),
.B(n_26),
.Y(n_69)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_70),
.Y(n_124)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_46),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_72),
.B(n_74),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_47),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_63),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_75),
.B(n_76),
.Y(n_110)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_48),
.Y(n_76)
);

BUFx2_ASAP7_75t_L g77 ( 
.A(n_64),
.Y(n_77)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_77),
.Y(n_119)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_55),
.Y(n_78)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_78),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_79),
.A2(n_86),
.B1(n_89),
.B2(n_90),
.Y(n_105)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_58),
.Y(n_80)
);

HB1xp67_ASAP7_75t_L g111 ( 
.A(n_80),
.Y(n_111)
);

A2O1A1Ixp33_ASAP7_75t_SL g82 ( 
.A1(n_69),
.A2(n_32),
.B(n_31),
.C(n_41),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_SL g115 ( 
.A1(n_82),
.A2(n_92),
.B(n_97),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_53),
.B(n_36),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_85),
.B(n_91),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_61),
.A2(n_30),
.B1(n_20),
.B2(n_27),
.Y(n_86)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_64),
.Y(n_88)
);

BUFx2_ASAP7_75t_L g112 ( 
.A(n_88),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_52),
.B(n_42),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_49),
.B(n_17),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_93),
.B(n_94),
.Y(n_118)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_55),
.Y(n_94)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_67),
.Y(n_95)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_95),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_49),
.B(n_17),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_96),
.B(n_99),
.Y(n_122)
);

OR2x2_ASAP7_75t_SL g97 ( 
.A(n_69),
.B(n_26),
.Y(n_97)
);

XNOR2xp5_ASAP7_75t_L g123 ( 
.A(n_98),
.B(n_7),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_54),
.B(n_17),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_68),
.B(n_4),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_100),
.B(n_26),
.C(n_6),
.Y(n_114)
);

INVx8_ASAP7_75t_L g102 ( 
.A(n_83),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_102),
.B(n_126),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_75),
.A2(n_68),
.B1(n_46),
.B2(n_66),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_103),
.A2(n_104),
.B1(n_107),
.B2(n_108),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_89),
.A2(n_68),
.B1(n_43),
.B2(n_39),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_91),
.A2(n_43),
.B1(n_57),
.B2(n_65),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_98),
.A2(n_65),
.B1(n_41),
.B2(n_22),
.Y(n_108)
);

AOI32xp33_ASAP7_75t_L g109 ( 
.A1(n_97),
.A2(n_38),
.A3(n_51),
.B1(n_26),
.B2(n_12),
.Y(n_109)
);

MAJx2_ASAP7_75t_L g138 ( 
.A(n_109),
.B(n_114),
.C(n_123),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_92),
.A2(n_51),
.B1(n_26),
.B2(n_38),
.Y(n_113)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_113),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g136 ( 
.A(n_114),
.B(n_123),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_82),
.A2(n_5),
.B1(n_7),
.B2(n_8),
.Y(n_117)
);

CKINVDCx14_ASAP7_75t_R g144 ( 
.A(n_117),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_82),
.A2(n_5),
.B1(n_7),
.B2(n_9),
.Y(n_120)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_120),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_73),
.B(n_9),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_125),
.B(n_127),
.Y(n_146)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_72),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_73),
.B(n_9),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_L g128 ( 
.A1(n_110),
.A2(n_82),
.B(n_100),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_L g156 ( 
.A1(n_128),
.A2(n_141),
.B(n_127),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_124),
.B(n_74),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_130),
.B(n_140),
.Y(n_152)
);

AND2x2_ASAP7_75t_L g131 ( 
.A(n_108),
.B(n_82),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_SL g160 ( 
.A1(n_131),
.A2(n_138),
.B(n_121),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_115),
.B(n_81),
.C(n_84),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_132),
.B(n_133),
.C(n_148),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_115),
.B(n_87),
.C(n_94),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_111),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_134),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_112),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_135),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_112),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_137),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_104),
.A2(n_100),
.B1(n_80),
.B2(n_76),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_139),
.A2(n_105),
.B1(n_103),
.B2(n_122),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_116),
.B(n_101),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_L g141 ( 
.A1(n_116),
.A2(n_71),
.B(n_78),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_118),
.B(n_71),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_145),
.B(n_149),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_107),
.B(n_95),
.C(n_88),
.Y(n_148)
);

INVx5_ASAP7_75t_L g149 ( 
.A(n_126),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_142),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_150),
.B(n_154),
.Y(n_172)
);

AOI21xp5_ASAP7_75t_L g151 ( 
.A1(n_133),
.A2(n_122),
.B(n_118),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_SL g167 ( 
.A1(n_151),
.A2(n_160),
.B(n_143),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_156),
.B(n_158),
.Y(n_168)
);

AOI322xp5_ASAP7_75t_SL g158 ( 
.A1(n_138),
.A2(n_125),
.A3(n_121),
.B1(n_13),
.B2(n_14),
.C1(n_15),
.C2(n_11),
.Y(n_158)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_148),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_161),
.B(n_132),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_141),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_162),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_146),
.B(n_119),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_163),
.B(n_147),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_149),
.B(n_119),
.Y(n_165)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_165),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_146),
.B(n_106),
.Y(n_166)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_166),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_167),
.B(n_173),
.C(n_176),
.Y(n_190)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_170),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_162),
.A2(n_143),
.B1(n_144),
.B2(n_129),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_174),
.A2(n_180),
.B1(n_154),
.B2(n_151),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_164),
.B(n_136),
.C(n_129),
.Y(n_176)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_159),
.Y(n_177)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_177),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_164),
.B(n_136),
.C(n_128),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_SL g186 ( 
.A(n_178),
.B(n_156),
.Y(n_186)
);

AOI21xp5_ASAP7_75t_L g179 ( 
.A1(n_160),
.A2(n_131),
.B(n_134),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_SL g181 ( 
.A1(n_179),
.A2(n_163),
.B(n_166),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_161),
.A2(n_139),
.B1(n_131),
.B2(n_102),
.Y(n_180)
);

AOI21xp5_ASAP7_75t_SL g198 ( 
.A1(n_181),
.A2(n_179),
.B(n_169),
.Y(n_198)
);

BUFx24_ASAP7_75t_SL g184 ( 
.A(n_168),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_184),
.B(n_168),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_185),
.A2(n_171),
.B1(n_176),
.B2(n_180),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_186),
.B(n_178),
.C(n_167),
.Y(n_197)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_170),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_187),
.B(n_188),
.Y(n_194)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_175),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_172),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_189),
.B(n_191),
.Y(n_195)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_174),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_181),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_192),
.B(n_196),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_193),
.A2(n_195),
.B1(n_197),
.B2(n_190),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_182),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_197),
.B(n_199),
.Y(n_205)
);

AOI21xp5_ASAP7_75t_L g206 ( 
.A1(n_198),
.A2(n_157),
.B(n_152),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_190),
.B(n_157),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_L g204 ( 
.A1(n_200),
.A2(n_183),
.B(n_188),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_201),
.B(n_204),
.C(n_202),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_194),
.B(n_183),
.Y(n_202)
);

AOI21xp5_ASAP7_75t_L g210 ( 
.A1(n_202),
.A2(n_206),
.B(n_198),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_207),
.B(n_208),
.C(n_209),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_203),
.B(n_200),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_205),
.B(n_150),
.C(n_155),
.Y(n_209)
);

AOI21xp5_ASAP7_75t_L g213 ( 
.A1(n_210),
.A2(n_152),
.B(n_158),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_L g212 ( 
.A1(n_208),
.A2(n_155),
.B(n_153),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_212),
.B(n_213),
.C(n_165),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_211),
.B(n_153),
.Y(n_214)
);

O2A1O1Ixp33_ASAP7_75t_L g217 ( 
.A1(n_214),
.A2(n_11),
.B(n_12),
.C(n_77),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_215),
.A2(n_177),
.B1(n_106),
.B2(n_15),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_216),
.B(n_217),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_218),
.B(n_83),
.Y(n_219)
);


endmodule