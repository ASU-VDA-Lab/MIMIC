module fake_jpeg_9229_n_337 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_337);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_337;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g17 ( 
.A(n_16),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

INVx11_ASAP7_75t_SL g21 ( 
.A(n_0),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_1),
.Y(n_23)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

BUFx10_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_8),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_5),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

BUFx10_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_4),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

BUFx16f_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_5),
.Y(n_35)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_22),
.Y(n_36)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_36),
.Y(n_64)
);

INVx2_ASAP7_75t_SL g37 ( 
.A(n_24),
.Y(n_37)
);

INVx3_ASAP7_75t_SL g49 ( 
.A(n_37),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_21),
.Y(n_38)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_38),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_21),
.Y(n_39)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_22),
.Y(n_40)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_22),
.Y(n_41)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_22),
.Y(n_42)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_42),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_22),
.Y(n_43)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_43),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_22),
.Y(n_44)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_44),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_45),
.Y(n_54)
);

INVx11_ASAP7_75t_L g46 ( 
.A(n_31),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_46),
.Y(n_63)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_47),
.B(n_24),
.Y(n_58)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_46),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_50),
.B(n_51),
.Y(n_79)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_46),
.Y(n_51)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_46),
.Y(n_52)
);

INVx11_ASAP7_75t_L g82 ( 
.A(n_52),
.Y(n_82)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_46),
.Y(n_53)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_53),
.Y(n_74)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_45),
.Y(n_55)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_55),
.Y(n_98)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_37),
.Y(n_57)
);

HB1xp67_ASAP7_75t_L g77 ( 
.A(n_57),
.Y(n_77)
);

CKINVDCx16_ASAP7_75t_R g73 ( 
.A(n_58),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_47),
.B(n_27),
.Y(n_61)
);

CKINVDCx14_ASAP7_75t_R g97 ( 
.A(n_61),
.Y(n_97)
);

OA22x2_ASAP7_75t_L g62 ( 
.A1(n_37),
.A2(n_34),
.B1(n_35),
.B2(n_28),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_L g71 ( 
.A1(n_62),
.A2(n_20),
.B1(n_24),
.B2(n_37),
.Y(n_71)
);

INVx5_ASAP7_75t_L g68 ( 
.A(n_38),
.Y(n_68)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_68),
.Y(n_78)
);

CKINVDCx14_ASAP7_75t_R g69 ( 
.A(n_47),
.Y(n_69)
);

INVx1_ASAP7_75t_SL g94 ( 
.A(n_69),
.Y(n_94)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_37),
.Y(n_70)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_70),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_L g99 ( 
.A1(n_71),
.A2(n_36),
.B1(n_42),
.B2(n_59),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g72 ( 
.A(n_49),
.Y(n_72)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_72),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_L g75 ( 
.A1(n_60),
.A2(n_20),
.B1(n_37),
.B2(n_17),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_75),
.A2(n_67),
.B1(n_26),
.B2(n_33),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_60),
.A2(n_20),
.B1(n_17),
.B2(n_29),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_80),
.A2(n_89),
.B1(n_95),
.B2(n_26),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_L g81 ( 
.A1(n_62),
.A2(n_18),
.B(n_33),
.Y(n_81)
);

XNOR2xp5_ASAP7_75t_L g106 ( 
.A(n_81),
.B(n_87),
.Y(n_106)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_68),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_83),
.B(n_85),
.Y(n_102)
);

CKINVDCx16_ASAP7_75t_R g84 ( 
.A(n_49),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_84),
.B(n_38),
.Y(n_124)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_54),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_54),
.Y(n_86)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_86),
.Y(n_110)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_62),
.B(n_34),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g111 ( 
.A(n_87),
.B(n_88),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_66),
.B(n_34),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_65),
.A2(n_17),
.B1(n_19),
.B2(n_29),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_63),
.Y(n_90)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_90),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_59),
.Y(n_91)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_91),
.Y(n_117)
);

INVx13_ASAP7_75t_L g92 ( 
.A(n_66),
.Y(n_92)
);

INVx5_ASAP7_75t_L g125 ( 
.A(n_92),
.Y(n_125)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_65),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_93),
.B(n_39),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_67),
.A2(n_29),
.B1(n_19),
.B2(n_27),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_63),
.Y(n_96)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_96),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_99),
.A2(n_105),
.B1(n_109),
.B2(n_126),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_87),
.A2(n_42),
.B1(n_36),
.B2(n_64),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_100),
.A2(n_104),
.B1(n_85),
.B2(n_93),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_81),
.B(n_47),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_101),
.B(n_113),
.Y(n_129)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_82),
.Y(n_103)
);

INVx2_ASAP7_75t_SL g145 ( 
.A(n_103),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_73),
.A2(n_42),
.B1(n_36),
.B2(n_64),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g136 ( 
.A(n_106),
.B(n_0),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_97),
.B(n_27),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g153 ( 
.A(n_108),
.B(n_118),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_73),
.A2(n_36),
.B1(n_42),
.B2(n_56),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_88),
.B(n_41),
.Y(n_113)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_82),
.Y(n_114)
);

CKINVDCx16_ASAP7_75t_R g133 ( 
.A(n_114),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_84),
.A2(n_19),
.B1(n_18),
.B2(n_33),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_116),
.A2(n_30),
.B1(n_25),
.B2(n_31),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_94),
.B(n_23),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_79),
.Y(n_119)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_119),
.Y(n_132)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_120),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_121),
.A2(n_86),
.B1(n_23),
.B2(n_32),
.Y(n_130)
);

AND2x2_ASAP7_75t_L g122 ( 
.A(n_88),
.B(n_0),
.Y(n_122)
);

AOI21xp5_ASAP7_75t_L g150 ( 
.A1(n_122),
.A2(n_28),
.B(n_25),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_76),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_123),
.B(n_127),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_124),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_L g126 ( 
.A1(n_94),
.A2(n_18),
.B1(n_26),
.B2(n_35),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_72),
.B(n_40),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_76),
.A2(n_56),
.B1(n_48),
.B2(n_35),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_128),
.A2(n_78),
.B1(n_32),
.B2(n_28),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_130),
.A2(n_141),
.B1(n_146),
.B2(n_116),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_101),
.B(n_98),
.Y(n_134)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_134),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_106),
.B(n_98),
.C(n_74),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_135),
.B(n_119),
.C(n_107),
.Y(n_167)
);

XOR2x1_ASAP7_75t_L g182 ( 
.A(n_136),
.B(n_25),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_111),
.B(n_74),
.Y(n_137)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_137),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_SL g138 ( 
.A1(n_113),
.A2(n_91),
.B(n_45),
.Y(n_138)
);

AO21x1_ASAP7_75t_L g166 ( 
.A1(n_138),
.A2(n_149),
.B(n_110),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_100),
.A2(n_76),
.B1(n_92),
.B2(n_83),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_142),
.A2(n_143),
.B1(n_107),
.B2(n_110),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_111),
.A2(n_92),
.B1(n_78),
.B2(n_48),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_111),
.B(n_122),
.Y(n_147)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_147),
.Y(n_162)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_102),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_148),
.B(n_155),
.Y(n_180)
);

NAND3xp33_ASAP7_75t_L g149 ( 
.A(n_122),
.B(n_16),
.C(n_15),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_L g161 ( 
.A1(n_150),
.A2(n_154),
.B(n_124),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_151),
.A2(n_152),
.B1(n_112),
.B2(n_115),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_123),
.A2(n_77),
.B1(n_44),
.B2(n_43),
.Y(n_152)
);

AOI21xp5_ASAP7_75t_L g154 ( 
.A1(n_105),
.A2(n_45),
.B(n_30),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_127),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_L g193 ( 
.A1(n_157),
.A2(n_161),
.B1(n_179),
.B2(n_140),
.Y(n_193)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_152),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_159),
.B(n_169),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_160),
.A2(n_176),
.B1(n_184),
.B2(n_151),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_135),
.B(n_108),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_163),
.B(n_165),
.C(n_167),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_164),
.A2(n_173),
.B1(n_134),
.B2(n_137),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_135),
.B(n_109),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_SL g205 ( 
.A1(n_166),
.A2(n_170),
.B(n_177),
.Y(n_205)
);

HB1xp67_ASAP7_75t_L g168 ( 
.A(n_145),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_168),
.B(n_175),
.Y(n_204)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_131),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_130),
.A2(n_117),
.B1(n_125),
.B2(n_104),
.Y(n_170)
);

CKINVDCx14_ASAP7_75t_R g171 ( 
.A(n_142),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_171),
.B(n_172),
.Y(n_213)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_131),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_130),
.A2(n_117),
.B1(n_125),
.B2(n_112),
.Y(n_173)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_129),
.B(n_128),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_174),
.B(n_147),
.C(n_150),
.Y(n_192)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_143),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_141),
.A2(n_115),
.B1(n_44),
.B2(n_43),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g177 ( 
.A(n_138),
.Y(n_177)
);

CKINVDCx16_ASAP7_75t_R g178 ( 
.A(n_146),
.Y(n_178)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_178),
.Y(n_187)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_145),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g181 ( 
.A(n_145),
.Y(n_181)
);

CKINVDCx16_ASAP7_75t_R g188 ( 
.A(n_181),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_SL g194 ( 
.A(n_182),
.B(n_149),
.Y(n_194)
);

OA22x2_ASAP7_75t_L g183 ( 
.A1(n_154),
.A2(n_31),
.B1(n_40),
.B2(n_41),
.Y(n_183)
);

A2O1A1Ixp33_ASAP7_75t_SL g202 ( 
.A1(n_183),
.A2(n_90),
.B(n_96),
.C(n_31),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_129),
.A2(n_43),
.B1(n_44),
.B2(n_40),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_185),
.A2(n_193),
.B1(n_145),
.B2(n_103),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_177),
.A2(n_155),
.B1(n_144),
.B2(n_140),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_189),
.A2(n_206),
.B1(n_207),
.B2(n_25),
.Y(n_237)
);

CKINVDCx14_ASAP7_75t_R g216 ( 
.A(n_190),
.Y(n_216)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_180),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_191),
.B(n_197),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_192),
.B(n_211),
.C(n_118),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_SL g228 ( 
.A(n_194),
.B(n_198),
.Y(n_228)
);

AND2x6_ASAP7_75t_L g196 ( 
.A(n_165),
.B(n_136),
.Y(n_196)
);

BUFx2_ASAP7_75t_L g223 ( 
.A(n_196),
.Y(n_223)
);

INVx1_ASAP7_75t_SL g197 ( 
.A(n_181),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_SL g198 ( 
.A(n_163),
.B(n_182),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_184),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_199),
.B(n_203),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_176),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_200),
.B(n_201),
.Y(n_235)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_164),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_202),
.A2(n_209),
.B1(n_133),
.B2(n_114),
.Y(n_220)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_174),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_159),
.A2(n_148),
.B1(n_139),
.B2(n_153),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_160),
.A2(n_139),
.B1(n_153),
.B2(n_132),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_170),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_208),
.B(n_210),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_158),
.A2(n_162),
.B1(n_156),
.B2(n_161),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_183),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_167),
.B(n_136),
.C(n_132),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_166),
.B(n_136),
.Y(n_212)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_212),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_214),
.B(n_215),
.C(n_219),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_198),
.B(n_183),
.Y(n_215)
);

HB1xp67_ASAP7_75t_L g217 ( 
.A(n_197),
.Y(n_217)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_217),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_186),
.B(n_183),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_220),
.A2(n_224),
.B1(n_226),
.B2(n_229),
.Y(n_242)
);

OAI21xp5_ASAP7_75t_L g221 ( 
.A1(n_195),
.A2(n_133),
.B(n_16),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_SL g254 ( 
.A(n_221),
.B(n_237),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_206),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_222),
.B(n_227),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_187),
.A2(n_199),
.B1(n_209),
.B2(n_203),
.Y(n_224)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_204),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_213),
.A2(n_205),
.B1(n_196),
.B2(n_189),
.Y(n_229)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_188),
.Y(n_230)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_230),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_207),
.B(n_14),
.Y(n_231)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_231),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_L g232 ( 
.A1(n_185),
.A2(n_90),
.B1(n_96),
.B2(n_30),
.Y(n_232)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_232),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_186),
.B(n_45),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_234),
.B(n_40),
.Y(n_253)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_205),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_236),
.B(n_192),
.Y(n_246)
);

HB1xp67_ASAP7_75t_L g239 ( 
.A(n_202),
.Y(n_239)
);

CKINVDCx16_ASAP7_75t_R g257 ( 
.A(n_239),
.Y(n_257)
);

OAI21x1_ASAP7_75t_L g240 ( 
.A1(n_229),
.A2(n_194),
.B(n_212),
.Y(n_240)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_240),
.Y(n_271)
);

INVxp67_ASAP7_75t_L g244 ( 
.A(n_233),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_244),
.B(n_235),
.Y(n_263)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_246),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_L g248 ( 
.A1(n_220),
.A2(n_202),
.B1(n_211),
.B2(n_14),
.Y(n_248)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_248),
.Y(n_278)
);

HB1xp67_ASAP7_75t_L g249 ( 
.A(n_230),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_249),
.B(n_39),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_219),
.B(n_202),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_250),
.B(n_255),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_225),
.A2(n_12),
.B1(n_15),
.B2(n_14),
.Y(n_251)
);

OAI21xp5_ASAP7_75t_L g276 ( 
.A1(n_251),
.A2(n_245),
.B(n_254),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_253),
.B(n_258),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_234),
.B(n_45),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_214),
.B(n_41),
.C(n_40),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_256),
.B(n_260),
.C(n_261),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_215),
.B(n_44),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_224),
.B(n_43),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_259),
.B(n_238),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_238),
.B(n_41),
.C(n_39),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_228),
.B(n_41),
.Y(n_261)
);

INVxp67_ASAP7_75t_L g295 ( 
.A(n_263),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_265),
.B(n_258),
.Y(n_285)
);

AND2x2_ASAP7_75t_L g266 ( 
.A(n_260),
.B(n_223),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_266),
.B(n_270),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_L g269 ( 
.A1(n_262),
.A2(n_216),
.B1(n_223),
.B2(n_218),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_269),
.A2(n_274),
.B1(n_10),
.B2(n_11),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_SL g270 ( 
.A(n_247),
.B(n_237),
.Y(n_270)
);

AOI21xp5_ASAP7_75t_L g272 ( 
.A1(n_257),
.A2(n_241),
.B(n_242),
.Y(n_272)
);

OAI21xp5_ASAP7_75t_L g287 ( 
.A1(n_272),
.A2(n_273),
.B(n_276),
.Y(n_287)
);

AOI21xp5_ASAP7_75t_L g273 ( 
.A1(n_244),
.A2(n_243),
.B(n_221),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_254),
.A2(n_228),
.B1(n_2),
.B2(n_3),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_275),
.B(n_279),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_251),
.B(n_9),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_SL g280 ( 
.A(n_256),
.B(n_9),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_280),
.B(n_1),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_267),
.B(n_252),
.C(n_253),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_281),
.B(n_289),
.C(n_292),
.Y(n_297)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_283),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_285),
.B(n_266),
.Y(n_300)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_267),
.B(n_261),
.Y(n_286)
);

XOR2xp5_ASAP7_75t_L g298 ( 
.A(n_286),
.B(n_290),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_265),
.B(n_252),
.Y(n_288)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_288),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_268),
.B(n_39),
.C(n_38),
.Y(n_289)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_264),
.B(n_10),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_291),
.A2(n_293),
.B1(n_271),
.B2(n_263),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_268),
.B(n_39),
.C(n_38),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_278),
.A2(n_25),
.B1(n_30),
.B2(n_10),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_264),
.B(n_25),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_294),
.B(n_276),
.C(n_277),
.Y(n_302)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_299),
.Y(n_314)
);

XOR2xp5_ASAP7_75t_L g311 ( 
.A(n_300),
.B(n_7),
.Y(n_311)
);

XOR2xp5_ASAP7_75t_L g301 ( 
.A(n_286),
.B(n_272),
.Y(n_301)
);

AND2x2_ASAP7_75t_L g313 ( 
.A(n_301),
.B(n_303),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_302),
.B(n_306),
.C(n_308),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_281),
.B(n_273),
.C(n_266),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_282),
.B(n_274),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_SL g317 ( 
.A(n_305),
.B(n_307),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_287),
.B(n_284),
.C(n_290),
.Y(n_306)
);

AND2x2_ASAP7_75t_L g307 ( 
.A(n_295),
.B(n_9),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_289),
.B(n_30),
.C(n_8),
.Y(n_308)
);

AOI21x1_ASAP7_75t_L g309 ( 
.A1(n_301),
.A2(n_295),
.B(n_292),
.Y(n_309)
);

OAI22x1_ASAP7_75t_L g323 ( 
.A1(n_309),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_323)
);

AOI21xp5_ASAP7_75t_L g310 ( 
.A1(n_304),
.A2(n_11),
.B(n_15),
.Y(n_310)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_310),
.Y(n_319)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_311),
.Y(n_326)
);

OAI21xp5_ASAP7_75t_SL g312 ( 
.A1(n_305),
.A2(n_7),
.B(n_12),
.Y(n_312)
);

AOI21xp5_ASAP7_75t_L g322 ( 
.A1(n_312),
.A2(n_315),
.B(n_316),
.Y(n_322)
);

OAI21xp5_ASAP7_75t_L g315 ( 
.A1(n_297),
.A2(n_7),
.B(n_11),
.Y(n_315)
);

AND2x2_ASAP7_75t_L g316 ( 
.A(n_298),
.B(n_6),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_318),
.B(n_314),
.C(n_298),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_320),
.B(n_316),
.C(n_5),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_L g321 ( 
.A1(n_317),
.A2(n_307),
.B1(n_296),
.B2(n_6),
.Y(n_321)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_321),
.Y(n_329)
);

OAI21xp5_ASAP7_75t_SL g327 ( 
.A1(n_323),
.A2(n_325),
.B(n_322),
.Y(n_327)
);

OAI21xp5_ASAP7_75t_L g324 ( 
.A1(n_317),
.A2(n_2),
.B(n_3),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_324),
.B(n_4),
.C(n_30),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_SL g325 ( 
.A(n_313),
.B(n_4),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_327),
.B(n_321),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_328),
.B(n_330),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_331),
.B(n_329),
.C(n_326),
.Y(n_333)
);

AOI22xp5_ASAP7_75t_L g334 ( 
.A1(n_333),
.A2(n_319),
.B1(n_332),
.B2(n_38),
.Y(n_334)
);

OAI21xp5_ASAP7_75t_L g335 ( 
.A1(n_334),
.A2(n_38),
.B(n_39),
.Y(n_335)
);

XNOR2xp5_ASAP7_75t_L g336 ( 
.A(n_335),
.B(n_38),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_SL g337 ( 
.A(n_336),
.B(n_39),
.Y(n_337)
);


endmodule