module real_aes_7470_n_99 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_99);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_99;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_503;
wire n_357;
wire n_287;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_364;
wire n_421;
wire n_555;
wire n_319;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_379;
wire n_374;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_178;
wire n_409;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_725;
wire n_504;
wire n_455;
wire n_310;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_417;
wire n_363;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_527;
wire n_434;
wire n_502;
wire n_600;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_713;
wire n_404;
wire n_288;
wire n_598;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_720;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_249;
wire n_623;
wire n_721;
wire n_446;
wire n_221;
wire n_681;
wire n_156;
wire n_456;
wire n_359;
wire n_717;
wire n_712;
wire n_266;
wire n_183;
wire n_312;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_521;
wire n_140;
wire n_418;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_698;
wire n_371;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_719;
wire n_473;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_646;
wire n_710;
wire n_650;
wire n_105;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
NAND3xp33_ASAP7_75t_SL g104 ( .A(n_0), .B(n_85), .C(n_105), .Y(n_104) );
INVx1_ASAP7_75t_L g121 ( .A(n_0), .Y(n_121) );
A2O1A1Ixp33_ASAP7_75t_L g453 ( .A1(n_1), .A2(n_142), .B(n_154), .C(n_454), .Y(n_453) );
INVx1_ASAP7_75t_L g261 ( .A(n_2), .Y(n_261) );
AOI21xp5_ASAP7_75t_L g492 ( .A1(n_3), .A2(n_169), .B(n_493), .Y(n_492) );
NAND2xp5_ASAP7_75t_L g498 ( .A(n_4), .B(n_165), .Y(n_498) );
AOI21xp33_ASAP7_75t_L g168 ( .A1(n_5), .A2(n_169), .B(n_170), .Y(n_168) );
AND2x6_ASAP7_75t_L g142 ( .A(n_6), .B(n_143), .Y(n_142) );
AOI21xp5_ASAP7_75t_L g236 ( .A1(n_7), .A2(n_237), .B(n_238), .Y(n_236) );
NAND2xp5_ASAP7_75t_L g102 ( .A(n_8), .B(n_103), .Y(n_102) );
NOR2xp33_ASAP7_75t_L g122 ( .A(n_8), .B(n_39), .Y(n_122) );
INVx1_ASAP7_75t_L g469 ( .A(n_9), .Y(n_469) );
NAND2xp5_ASAP7_75t_SL g457 ( .A(n_10), .B(n_175), .Y(n_457) );
INVx1_ASAP7_75t_L g177 ( .A(n_11), .Y(n_177) );
NAND2xp5_ASAP7_75t_L g228 ( .A(n_12), .B(n_229), .Y(n_228) );
INVx1_ASAP7_75t_L g139 ( .A(n_13), .Y(n_139) );
INVx1_ASAP7_75t_L g243 ( .A(n_14), .Y(n_243) );
A2O1A1Ixp33_ASAP7_75t_L g477 ( .A1(n_15), .A2(n_178), .B(n_244), .C(n_478), .Y(n_477) );
NAND2xp5_ASAP7_75t_L g480 ( .A(n_16), .B(n_165), .Y(n_480) );
NAND2xp5_ASAP7_75t_L g215 ( .A(n_17), .B(n_188), .Y(n_215) );
NAND2xp5_ASAP7_75t_SL g197 ( .A(n_18), .B(n_169), .Y(n_197) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_19), .B(n_511), .Y(n_510) );
A2O1A1Ixp33_ASAP7_75t_L g485 ( .A1(n_20), .A2(n_145), .B(n_229), .C(n_486), .Y(n_485) );
NAND2xp5_ASAP7_75t_L g191 ( .A(n_21), .B(n_165), .Y(n_191) );
NAND2xp5_ASAP7_75t_SL g532 ( .A(n_22), .B(n_175), .Y(n_532) );
A2O1A1Ixp33_ASAP7_75t_L g240 ( .A1(n_23), .A2(n_241), .B(n_242), .C(n_244), .Y(n_240) );
NAND2xp5_ASAP7_75t_SL g519 ( .A(n_24), .B(n_175), .Y(n_519) );
CKINVDCx16_ASAP7_75t_R g528 ( .A(n_25), .Y(n_528) );
INVx1_ASAP7_75t_L g518 ( .A(n_26), .Y(n_518) );
BUFx6f_ASAP7_75t_L g150 ( .A(n_27), .Y(n_150) );
CKINVDCx20_ASAP7_75t_R g452 ( .A(n_28), .Y(n_452) );
NAND2xp5_ASAP7_75t_L g262 ( .A(n_29), .B(n_175), .Y(n_262) );
INVx1_ASAP7_75t_L g507 ( .A(n_30), .Y(n_507) );
INVx1_ASAP7_75t_L g153 ( .A(n_31), .Y(n_153) );
INVx2_ASAP7_75t_L g147 ( .A(n_32), .Y(n_147) );
CKINVDCx20_ASAP7_75t_R g459 ( .A(n_33), .Y(n_459) );
A2O1A1Ixp33_ASAP7_75t_L g495 ( .A1(n_34), .A2(n_179), .B(n_229), .C(n_496), .Y(n_495) );
INVxp67_ASAP7_75t_L g508 ( .A(n_35), .Y(n_508) );
A2O1A1Ixp33_ASAP7_75t_L g198 ( .A1(n_36), .A2(n_142), .B(n_154), .C(n_199), .Y(n_198) );
CKINVDCx14_ASAP7_75t_R g494 ( .A(n_37), .Y(n_494) );
A2O1A1Ixp33_ASAP7_75t_L g516 ( .A1(n_38), .A2(n_154), .B(n_517), .C(n_521), .Y(n_516) );
INVx1_ASAP7_75t_L g103 ( .A(n_39), .Y(n_103) );
INVx1_ASAP7_75t_L g151 ( .A(n_40), .Y(n_151) );
A2O1A1Ixp33_ASAP7_75t_L g467 ( .A1(n_41), .A2(n_174), .B(n_204), .C(n_468), .Y(n_467) );
NAND2xp5_ASAP7_75t_SL g214 ( .A(n_42), .B(n_175), .Y(n_214) );
CKINVDCx20_ASAP7_75t_R g523 ( .A(n_43), .Y(n_523) );
CKINVDCx20_ASAP7_75t_R g504 ( .A(n_44), .Y(n_504) );
CKINVDCx20_ASAP7_75t_R g123 ( .A(n_45), .Y(n_123) );
INVx1_ASAP7_75t_L g484 ( .A(n_46), .Y(n_484) );
CKINVDCx16_ASAP7_75t_R g157 ( .A(n_47), .Y(n_157) );
NAND2xp5_ASAP7_75t_L g231 ( .A(n_48), .B(n_169), .Y(n_231) );
AOI222xp33_ASAP7_75t_SL g124 ( .A1(n_49), .A2(n_59), .B1(n_125), .B2(n_711), .C1(n_712), .C2(n_716), .Y(n_124) );
AOI22xp33_ASAP7_75t_L g99 ( .A1(n_50), .A2(n_100), .B1(n_108), .B2(n_725), .Y(n_99) );
AOI22xp5_ASAP7_75t_L g144 ( .A1(n_51), .A2(n_145), .B1(n_148), .B2(n_154), .Y(n_144) );
CKINVDCx20_ASAP7_75t_R g208 ( .A(n_52), .Y(n_208) );
CKINVDCx16_ASAP7_75t_R g258 ( .A(n_53), .Y(n_258) );
A2O1A1Ixp33_ASAP7_75t_L g173 ( .A1(n_54), .A2(n_174), .B(n_176), .C(n_179), .Y(n_173) );
CKINVDCx14_ASAP7_75t_R g466 ( .A(n_55), .Y(n_466) );
CKINVDCx20_ASAP7_75t_R g218 ( .A(n_56), .Y(n_218) );
INVx1_ASAP7_75t_L g171 ( .A(n_57), .Y(n_171) );
INVx1_ASAP7_75t_L g143 ( .A(n_58), .Y(n_143) );
CKINVDCx20_ASAP7_75t_R g711 ( .A(n_59), .Y(n_711) );
INVx1_ASAP7_75t_L g138 ( .A(n_60), .Y(n_138) );
INVx1_ASAP7_75t_SL g497 ( .A(n_61), .Y(n_497) );
CKINVDCx20_ASAP7_75t_R g114 ( .A(n_62), .Y(n_114) );
NAND2xp5_ASAP7_75t_L g488 ( .A(n_63), .B(n_165), .Y(n_488) );
OAI22xp5_ASAP7_75t_SL g721 ( .A1(n_64), .A2(n_443), .B1(n_713), .B2(n_722), .Y(n_721) );
CKINVDCx20_ASAP7_75t_R g722 ( .A(n_64), .Y(n_722) );
INVx1_ASAP7_75t_L g531 ( .A(n_65), .Y(n_531) );
A2O1A1Ixp33_ASAP7_75t_SL g187 ( .A1(n_66), .A2(n_179), .B(n_188), .C(n_189), .Y(n_187) );
INVxp67_ASAP7_75t_L g190 ( .A(n_67), .Y(n_190) );
INVx1_ASAP7_75t_L g107 ( .A(n_68), .Y(n_107) );
AOI21xp5_ASAP7_75t_L g464 ( .A1(n_69), .A2(n_169), .B(n_465), .Y(n_464) );
CKINVDCx20_ASAP7_75t_R g535 ( .A(n_70), .Y(n_535) );
CKINVDCx20_ASAP7_75t_R g162 ( .A(n_71), .Y(n_162) );
AOI21xp5_ASAP7_75t_L g474 ( .A1(n_72), .A2(n_169), .B(n_475), .Y(n_474) );
INVx1_ASAP7_75t_L g211 ( .A(n_73), .Y(n_211) );
AOI21xp5_ASAP7_75t_L g502 ( .A1(n_74), .A2(n_237), .B(n_503), .Y(n_502) );
INVx1_ASAP7_75t_L g476 ( .A(n_75), .Y(n_476) );
CKINVDCx16_ASAP7_75t_R g515 ( .A(n_76), .Y(n_515) );
A2O1A1Ixp33_ASAP7_75t_L g212 ( .A1(n_77), .A2(n_142), .B(n_154), .C(n_213), .Y(n_212) );
AOI21xp5_ASAP7_75t_L g482 ( .A1(n_78), .A2(n_169), .B(n_483), .Y(n_482) );
INVx1_ASAP7_75t_L g479 ( .A(n_79), .Y(n_479) );
NAND2xp5_ASAP7_75t_SL g200 ( .A(n_80), .B(n_201), .Y(n_200) );
INVx2_ASAP7_75t_L g136 ( .A(n_81), .Y(n_136) );
INVx1_ASAP7_75t_L g455 ( .A(n_82), .Y(n_455) );
NAND2xp5_ASAP7_75t_L g202 ( .A(n_83), .B(n_188), .Y(n_202) );
A2O1A1Ixp33_ASAP7_75t_L g259 ( .A1(n_84), .A2(n_142), .B(n_154), .C(n_260), .Y(n_259) );
OR2x2_ASAP7_75t_L g118 ( .A(n_85), .B(n_119), .Y(n_118) );
INVx2_ASAP7_75t_L g442 ( .A(n_85), .Y(n_442) );
OR2x2_ASAP7_75t_L g710 ( .A(n_85), .B(n_120), .Y(n_710) );
A2O1A1Ixp33_ASAP7_75t_L g529 ( .A1(n_86), .A2(n_154), .B(n_530), .C(n_533), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g181 ( .A(n_87), .B(n_182), .Y(n_181) );
CKINVDCx20_ASAP7_75t_R g265 ( .A(n_88), .Y(n_265) );
A2O1A1Ixp33_ASAP7_75t_L g225 ( .A1(n_89), .A2(n_142), .B(n_154), .C(n_226), .Y(n_225) );
CKINVDCx20_ASAP7_75t_R g233 ( .A(n_90), .Y(n_233) );
INVx1_ASAP7_75t_L g186 ( .A(n_91), .Y(n_186) );
CKINVDCx16_ASAP7_75t_R g239 ( .A(n_92), .Y(n_239) );
NAND2xp5_ASAP7_75t_SL g227 ( .A(n_93), .B(n_201), .Y(n_227) );
NAND2xp5_ASAP7_75t_L g470 ( .A(n_94), .B(n_167), .Y(n_470) );
NAND2xp5_ASAP7_75t_L g245 ( .A(n_95), .B(n_167), .Y(n_245) );
NAND2xp5_ASAP7_75t_L g106 ( .A(n_96), .B(n_107), .Y(n_106) );
AOI21xp5_ASAP7_75t_L g184 ( .A1(n_97), .A2(n_169), .B(n_185), .Y(n_184) );
INVx2_ASAP7_75t_L g487 ( .A(n_98), .Y(n_487) );
INVx1_ASAP7_75t_L g100 ( .A(n_101), .Y(n_100) );
CKINVDCx6p67_ASAP7_75t_R g726 ( .A(n_101), .Y(n_726) );
OR2x2_ASAP7_75t_L g101 ( .A(n_102), .B(n_104), .Y(n_101) );
INVx1_ASAP7_75t_SL g105 ( .A(n_106), .Y(n_105) );
BUFx2_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
AOI22xp5_ASAP7_75t_L g109 ( .A1(n_110), .A2(n_124), .B1(n_719), .B2(n_720), .Y(n_109) );
NOR2xp33_ASAP7_75t_L g110 ( .A(n_111), .B(n_115), .Y(n_110) );
INVx1_ASAP7_75t_SL g111 ( .A(n_112), .Y(n_111) );
INVx1_ASAP7_75t_SL g719 ( .A(n_112), .Y(n_719) );
BUFx2_ASAP7_75t_L g112 ( .A(n_113), .Y(n_112) );
INVx2_ASAP7_75t_L g113 ( .A(n_114), .Y(n_113) );
AOI21xp5_ASAP7_75t_L g720 ( .A1(n_115), .A2(n_721), .B(n_723), .Y(n_720) );
NOR2xp33_ASAP7_75t_SL g115 ( .A(n_116), .B(n_123), .Y(n_115) );
INVx1_ASAP7_75t_SL g116 ( .A(n_117), .Y(n_116) );
INVx1_ASAP7_75t_SL g117 ( .A(n_118), .Y(n_117) );
INVx1_ASAP7_75t_SL g724 ( .A(n_118), .Y(n_724) );
NOR2x2_ASAP7_75t_L g718 ( .A(n_119), .B(n_442), .Y(n_718) );
INVx2_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
OR2x2_ASAP7_75t_L g441 ( .A(n_120), .B(n_442), .Y(n_441) );
AND2x2_ASAP7_75t_L g120 ( .A(n_121), .B(n_122), .Y(n_120) );
OAI22xp5_ASAP7_75t_SL g125 ( .A1(n_126), .A2(n_439), .B1(n_443), .B2(n_710), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
OAI22xp5_ASAP7_75t_SL g712 ( .A1(n_127), .A2(n_439), .B1(n_713), .B2(n_714), .Y(n_712) );
AND3x1_ASAP7_75t_L g127 ( .A(n_128), .B(n_364), .C(n_413), .Y(n_127) );
NOR3xp33_ASAP7_75t_SL g128 ( .A(n_129), .B(n_271), .C(n_309), .Y(n_128) );
OAI222xp33_ASAP7_75t_L g129 ( .A1(n_130), .A2(n_192), .B1(n_246), .B2(n_252), .C1(n_266), .C2(n_269), .Y(n_129) );
NAND2xp5_ASAP7_75t_L g130 ( .A(n_131), .B(n_163), .Y(n_130) );
NAND2xp5_ASAP7_75t_L g338 ( .A(n_131), .B(n_339), .Y(n_338) );
NAND2xp5_ASAP7_75t_L g405 ( .A(n_131), .B(n_314), .Y(n_405) );
BUFx2_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
OR2x2_ASAP7_75t_L g282 ( .A(n_132), .B(n_183), .Y(n_282) );
NAND2xp5_ASAP7_75t_L g290 ( .A(n_132), .B(n_164), .Y(n_290) );
AND2x2_ASAP7_75t_L g325 ( .A(n_132), .B(n_302), .Y(n_325) );
OR2x2_ASAP7_75t_L g349 ( .A(n_132), .B(n_164), .Y(n_349) );
OR2x2_ASAP7_75t_L g357 ( .A(n_132), .B(n_256), .Y(n_357) );
AND2x2_ASAP7_75t_L g360 ( .A(n_132), .B(n_183), .Y(n_360) );
INVx3_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
OR2x2_ASAP7_75t_L g254 ( .A(n_133), .B(n_255), .Y(n_254) );
AND2x2_ASAP7_75t_L g268 ( .A(n_133), .B(n_183), .Y(n_268) );
AND2x2_ASAP7_75t_L g318 ( .A(n_133), .B(n_256), .Y(n_318) );
AND2x2_ASAP7_75t_L g331 ( .A(n_133), .B(n_164), .Y(n_331) );
NOR2xp33_ASAP7_75t_L g438 ( .A(n_133), .B(n_417), .Y(n_438) );
AO21x2_ASAP7_75t_L g133 ( .A1(n_134), .A2(n_140), .B(n_161), .Y(n_133) );
NOR2xp33_ASAP7_75t_L g161 ( .A(n_134), .B(n_162), .Y(n_161) );
INVx2_ASAP7_75t_L g206 ( .A(n_134), .Y(n_206) );
AO21x2_ASAP7_75t_L g256 ( .A1(n_134), .A2(n_257), .B(n_264), .Y(n_256) );
INVx1_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
BUFx6f_ASAP7_75t_L g167 ( .A(n_135), .Y(n_167) );
AND2x2_ASAP7_75t_L g135 ( .A(n_136), .B(n_137), .Y(n_135) );
AND2x2_ASAP7_75t_SL g182 ( .A(n_136), .B(n_137), .Y(n_182) );
NAND2xp5_ASAP7_75t_L g137 ( .A(n_138), .B(n_139), .Y(n_137) );
OAI22xp33_ASAP7_75t_L g140 ( .A1(n_141), .A2(n_144), .B1(n_157), .B2(n_158), .Y(n_140) );
O2A1O1Ixp33_ASAP7_75t_L g170 ( .A1(n_141), .A2(n_171), .B(n_172), .C(n_173), .Y(n_170) );
O2A1O1Ixp33_ASAP7_75t_L g185 ( .A1(n_141), .A2(n_172), .B(n_186), .C(n_187), .Y(n_185) );
O2A1O1Ixp33_ASAP7_75t_L g238 ( .A1(n_141), .A2(n_172), .B(n_239), .C(n_240), .Y(n_238) );
O2A1O1Ixp33_ASAP7_75t_SL g465 ( .A1(n_141), .A2(n_172), .B(n_466), .C(n_467), .Y(n_465) );
O2A1O1Ixp33_ASAP7_75t_SL g475 ( .A1(n_141), .A2(n_172), .B(n_476), .C(n_477), .Y(n_475) );
O2A1O1Ixp33_ASAP7_75t_SL g483 ( .A1(n_141), .A2(n_172), .B(n_484), .C(n_485), .Y(n_483) );
O2A1O1Ixp33_ASAP7_75t_L g493 ( .A1(n_141), .A2(n_172), .B(n_494), .C(n_495), .Y(n_493) );
O2A1O1Ixp33_ASAP7_75t_SL g503 ( .A1(n_141), .A2(n_172), .B(n_504), .C(n_505), .Y(n_503) );
INVx1_ASAP7_75t_L g533 ( .A(n_141), .Y(n_533) );
INVx4_ASAP7_75t_SL g141 ( .A(n_142), .Y(n_141) );
NAND2x1p5_ASAP7_75t_L g158 ( .A(n_142), .B(n_159), .Y(n_158) );
AND2x4_ASAP7_75t_L g169 ( .A(n_142), .B(n_159), .Y(n_169) );
BUFx3_ASAP7_75t_L g521 ( .A(n_142), .Y(n_521) );
INVx2_ASAP7_75t_L g263 ( .A(n_145), .Y(n_263) );
INVx3_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
INVx1_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
INVx2_ASAP7_75t_L g155 ( .A(n_147), .Y(n_155) );
INVx1_ASAP7_75t_L g160 ( .A(n_147), .Y(n_160) );
OAI22xp5_ASAP7_75t_SL g148 ( .A1(n_149), .A2(n_151), .B1(n_152), .B2(n_153), .Y(n_148) );
INVx2_ASAP7_75t_L g152 ( .A(n_149), .Y(n_152) );
INVx4_ASAP7_75t_L g241 ( .A(n_149), .Y(n_241) );
BUFx6f_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
INVx1_ASAP7_75t_L g156 ( .A(n_150), .Y(n_156) );
AND2x2_ASAP7_75t_L g159 ( .A(n_150), .B(n_160), .Y(n_159) );
BUFx6f_ASAP7_75t_L g175 ( .A(n_150), .Y(n_175) );
INVx3_ASAP7_75t_L g178 ( .A(n_150), .Y(n_178) );
INVx1_ASAP7_75t_L g188 ( .A(n_150), .Y(n_188) );
INVx2_ASAP7_75t_L g456 ( .A(n_152), .Y(n_456) );
INVx5_ASAP7_75t_L g172 ( .A(n_154), .Y(n_172) );
AND2x6_ASAP7_75t_L g154 ( .A(n_155), .B(n_156), .Y(n_154) );
BUFx6f_ASAP7_75t_L g180 ( .A(n_155), .Y(n_180) );
BUFx3_ASAP7_75t_L g205 ( .A(n_155), .Y(n_205) );
OAI21xp5_ASAP7_75t_L g210 ( .A1(n_158), .A2(n_211), .B(n_212), .Y(n_210) );
OAI21xp5_ASAP7_75t_L g257 ( .A1(n_158), .A2(n_258), .B(n_259), .Y(n_257) );
OAI21xp5_ASAP7_75t_L g451 ( .A1(n_158), .A2(n_452), .B(n_453), .Y(n_451) );
O2A1O1Ixp33_ASAP7_75t_L g514 ( .A1(n_158), .A2(n_182), .B(n_515), .C(n_516), .Y(n_514) );
OAI21xp5_ASAP7_75t_L g527 ( .A1(n_158), .A2(n_528), .B(n_529), .Y(n_527) );
INVx1_ASAP7_75t_L g509 ( .A(n_160), .Y(n_509) );
O2A1O1Ixp33_ASAP7_75t_L g356 ( .A1(n_163), .A2(n_357), .B(n_358), .C(n_361), .Y(n_356) );
NAND2xp5_ASAP7_75t_L g385 ( .A(n_163), .B(n_386), .Y(n_385) );
NAND2xp5_ASAP7_75t_L g423 ( .A(n_163), .B(n_301), .Y(n_423) );
AND2x2_ASAP7_75t_L g163 ( .A(n_164), .B(n_183), .Y(n_163) );
AND2x2_ASAP7_75t_SL g267 ( .A(n_164), .B(n_268), .Y(n_267) );
INVx2_ASAP7_75t_L g281 ( .A(n_164), .Y(n_281) );
AND2x2_ASAP7_75t_L g308 ( .A(n_164), .B(n_302), .Y(n_308) );
INVx1_ASAP7_75t_SL g316 ( .A(n_164), .Y(n_316) );
AND2x2_ASAP7_75t_L g339 ( .A(n_164), .B(n_340), .Y(n_339) );
BUFx2_ASAP7_75t_L g417 ( .A(n_164), .Y(n_417) );
OA21x2_ASAP7_75t_L g164 ( .A1(n_165), .A2(n_168), .B(n_181), .Y(n_164) );
INVx3_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
NOR2xp33_ASAP7_75t_SL g207 ( .A(n_166), .B(n_208), .Y(n_207) );
NOR2xp33_ASAP7_75t_L g458 ( .A(n_166), .B(n_459), .Y(n_458) );
NOR2xp33_ASAP7_75t_L g522 ( .A(n_166), .B(n_523), .Y(n_522) );
AO21x2_ASAP7_75t_L g526 ( .A1(n_166), .A2(n_527), .B(n_534), .Y(n_526) );
INVx4_ASAP7_75t_L g166 ( .A(n_167), .Y(n_166) );
OA21x2_ASAP7_75t_L g183 ( .A1(n_167), .A2(n_184), .B(n_191), .Y(n_183) );
HB1xp67_ASAP7_75t_L g473 ( .A(n_167), .Y(n_473) );
BUFx2_ASAP7_75t_L g237 ( .A(n_169), .Y(n_237) );
INVx2_ASAP7_75t_L g174 ( .A(n_175), .Y(n_174) );
INVx4_ASAP7_75t_L g229 ( .A(n_175), .Y(n_229) );
NOR2xp33_ASAP7_75t_L g176 ( .A(n_177), .B(n_178), .Y(n_176) );
NOR2xp33_ASAP7_75t_L g189 ( .A(n_178), .B(n_190), .Y(n_189) );
INVx5_ASAP7_75t_L g201 ( .A(n_178), .Y(n_201) );
NOR2xp33_ASAP7_75t_L g468 ( .A(n_178), .B(n_469), .Y(n_468) );
INVx3_ASAP7_75t_L g179 ( .A(n_180), .Y(n_179) );
HB1xp67_ASAP7_75t_L g230 ( .A(n_180), .Y(n_230) );
INVx1_ASAP7_75t_L g219 ( .A(n_182), .Y(n_219) );
INVx2_ASAP7_75t_L g223 ( .A(n_182), .Y(n_223) );
OA21x2_ASAP7_75t_L g235 ( .A1(n_182), .A2(n_236), .B(n_245), .Y(n_235) );
OA21x2_ASAP7_75t_L g463 ( .A1(n_182), .A2(n_464), .B(n_470), .Y(n_463) );
BUFx2_ASAP7_75t_L g253 ( .A(n_183), .Y(n_253) );
INVx1_ASAP7_75t_L g315 ( .A(n_183), .Y(n_315) );
INVx3_ASAP7_75t_L g340 ( .A(n_183), .Y(n_340) );
NAND2xp5_ASAP7_75t_SL g273 ( .A(n_192), .B(n_274), .Y(n_273) );
OR2x2_ASAP7_75t_L g192 ( .A(n_193), .B(n_220), .Y(n_192) );
INVx1_ASAP7_75t_L g336 ( .A(n_193), .Y(n_336) );
OAI32xp33_ASAP7_75t_L g342 ( .A1(n_193), .A2(n_281), .A3(n_343), .B1(n_344), .B2(n_345), .Y(n_342) );
OAI22xp5_ASAP7_75t_L g346 ( .A1(n_193), .A2(n_347), .B1(n_350), .B2(n_355), .Y(n_346) );
INVx4_ASAP7_75t_L g193 ( .A(n_194), .Y(n_193) );
AND2x2_ASAP7_75t_L g284 ( .A(n_194), .B(n_285), .Y(n_284) );
AND2x2_ASAP7_75t_L g362 ( .A(n_194), .B(n_363), .Y(n_362) );
AND2x2_ASAP7_75t_L g432 ( .A(n_194), .B(n_378), .Y(n_432) );
AND2x2_ASAP7_75t_L g194 ( .A(n_195), .B(n_209), .Y(n_194) );
AND2x2_ASAP7_75t_L g247 ( .A(n_195), .B(n_248), .Y(n_247) );
INVx2_ASAP7_75t_L g277 ( .A(n_195), .Y(n_277) );
INVx1_ASAP7_75t_L g296 ( .A(n_195), .Y(n_296) );
OR2x2_ASAP7_75t_L g304 ( .A(n_195), .B(n_305), .Y(n_304) );
AND2x2_ASAP7_75t_L g311 ( .A(n_195), .B(n_285), .Y(n_311) );
NOR2xp33_ASAP7_75t_L g319 ( .A(n_195), .B(n_320), .Y(n_319) );
AND2x2_ASAP7_75t_L g332 ( .A(n_195), .B(n_250), .Y(n_332) );
INVx3_ASAP7_75t_L g354 ( .A(n_195), .Y(n_354) );
AND2x2_ASAP7_75t_L g379 ( .A(n_195), .B(n_251), .Y(n_379) );
NOR2xp33_ASAP7_75t_L g427 ( .A(n_195), .B(n_344), .Y(n_427) );
OR2x6_ASAP7_75t_L g195 ( .A(n_196), .B(n_207), .Y(n_195) );
AOI21xp5_ASAP7_75t_SL g196 ( .A1(n_197), .A2(n_198), .B(n_206), .Y(n_196) );
AOI21xp5_ASAP7_75t_L g199 ( .A1(n_200), .A2(n_202), .B(n_203), .Y(n_199) );
O2A1O1Ixp33_ASAP7_75t_L g260 ( .A1(n_201), .A2(n_261), .B(n_262), .C(n_263), .Y(n_260) );
OAI22xp33_ASAP7_75t_L g506 ( .A1(n_201), .A2(n_241), .B1(n_507), .B2(n_508), .Y(n_506) );
O2A1O1Ixp33_ASAP7_75t_L g517 ( .A1(n_201), .A2(n_518), .B(n_519), .C(n_520), .Y(n_517) );
AOI21xp5_ASAP7_75t_L g213 ( .A1(n_203), .A2(n_214), .B(n_215), .Y(n_213) );
O2A1O1Ixp5_ASAP7_75t_L g454 ( .A1(n_203), .A2(n_455), .B(n_456), .C(n_457), .Y(n_454) );
O2A1O1Ixp33_ASAP7_75t_L g530 ( .A1(n_203), .A2(n_456), .B(n_531), .C(n_532), .Y(n_530) );
INVx2_ASAP7_75t_L g203 ( .A(n_204), .Y(n_203) );
INVx2_ASAP7_75t_L g204 ( .A(n_205), .Y(n_204) );
INVx1_ASAP7_75t_L g244 ( .A(n_205), .Y(n_244) );
INVx1_ASAP7_75t_L g216 ( .A(n_206), .Y(n_216) );
INVx2_ASAP7_75t_L g251 ( .A(n_209), .Y(n_251) );
AND2x2_ASAP7_75t_L g383 ( .A(n_209), .B(n_221), .Y(n_383) );
AO21x2_ASAP7_75t_L g209 ( .A1(n_210), .A2(n_216), .B(n_217), .Y(n_209) );
INVx1_ASAP7_75t_L g501 ( .A(n_216), .Y(n_501) );
AO21x2_ASAP7_75t_L g553 ( .A1(n_216), .A2(n_554), .B(n_555), .Y(n_553) );
NOR2xp33_ASAP7_75t_L g217 ( .A(n_218), .B(n_219), .Y(n_217) );
NOR2xp33_ASAP7_75t_L g232 ( .A(n_219), .B(n_233), .Y(n_232) );
NOR2xp33_ASAP7_75t_L g264 ( .A(n_219), .B(n_265), .Y(n_264) );
AO21x2_ASAP7_75t_L g450 ( .A1(n_219), .A2(n_451), .B(n_458), .Y(n_450) );
INVx2_ASAP7_75t_L g425 ( .A(n_220), .Y(n_425) );
OR2x2_ASAP7_75t_L g220 ( .A(n_221), .B(n_234), .Y(n_220) );
INVx1_ASAP7_75t_L g270 ( .A(n_221), .Y(n_270) );
AND2x2_ASAP7_75t_L g297 ( .A(n_221), .B(n_298), .Y(n_297) );
NAND2xp5_ASAP7_75t_L g305 ( .A(n_221), .B(n_251), .Y(n_305) );
AND2x2_ASAP7_75t_L g363 ( .A(n_221), .B(n_286), .Y(n_363) );
INVx2_ASAP7_75t_L g221 ( .A(n_222), .Y(n_221) );
INVx1_ASAP7_75t_L g249 ( .A(n_222), .Y(n_249) );
AND2x2_ASAP7_75t_L g276 ( .A(n_222), .B(n_277), .Y(n_276) );
AND2x2_ASAP7_75t_L g285 ( .A(n_222), .B(n_286), .Y(n_285) );
NAND2xp5_ASAP7_75t_L g351 ( .A(n_222), .B(n_251), .Y(n_351) );
AO21x2_ASAP7_75t_L g222 ( .A1(n_223), .A2(n_224), .B(n_232), .Y(n_222) );
INVx1_ASAP7_75t_L g511 ( .A(n_223), .Y(n_511) );
NOR2xp33_ASAP7_75t_L g534 ( .A(n_223), .B(n_535), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g224 ( .A(n_225), .B(n_231), .Y(n_224) );
AOI21xp5_ASAP7_75t_L g226 ( .A1(n_227), .A2(n_228), .B(n_230), .Y(n_226) );
NOR2xp33_ASAP7_75t_L g496 ( .A(n_229), .B(n_497), .Y(n_496) );
NAND2xp5_ASAP7_75t_L g278 ( .A(n_234), .B(n_279), .Y(n_278) );
INVx2_ASAP7_75t_L g298 ( .A(n_234), .Y(n_298) );
NAND2xp5_ASAP7_75t_L g344 ( .A(n_234), .B(n_251), .Y(n_344) );
AND2x2_ASAP7_75t_L g353 ( .A(n_234), .B(n_354), .Y(n_353) );
INVx1_ASAP7_75t_L g378 ( .A(n_234), .Y(n_378) );
INVx2_ASAP7_75t_L g234 ( .A(n_235), .Y(n_234) );
AND2x2_ASAP7_75t_L g250 ( .A(n_235), .B(n_251), .Y(n_250) );
INVx1_ASAP7_75t_L g286 ( .A(n_235), .Y(n_286) );
NOR2xp33_ASAP7_75t_L g242 ( .A(n_241), .B(n_243), .Y(n_242) );
NOR2xp33_ASAP7_75t_L g478 ( .A(n_241), .B(n_479), .Y(n_478) );
NOR2xp33_ASAP7_75t_L g486 ( .A(n_241), .B(n_487), .Y(n_486) );
OAI22xp5_ASAP7_75t_L g414 ( .A1(n_246), .A2(n_256), .B1(n_415), .B2(n_418), .Y(n_414) );
INVx1_ASAP7_75t_SL g246 ( .A(n_247), .Y(n_246) );
OAI21xp5_ASAP7_75t_SL g437 ( .A1(n_248), .A2(n_359), .B(n_438), .Y(n_437) );
AND2x2_ASAP7_75t_L g248 ( .A(n_249), .B(n_250), .Y(n_248) );
NOR2xp33_ASAP7_75t_L g371 ( .A(n_249), .B(n_354), .Y(n_371) );
INVx1_ASAP7_75t_L g396 ( .A(n_249), .Y(n_396) );
NAND2xp5_ASAP7_75t_L g269 ( .A(n_250), .B(n_270), .Y(n_269) );
AND2x2_ASAP7_75t_L g323 ( .A(n_250), .B(n_276), .Y(n_323) );
INVx2_ASAP7_75t_L g279 ( .A(n_251), .Y(n_279) );
INVx1_ASAP7_75t_L g329 ( .A(n_251), .Y(n_329) );
OAI221xp5_ASAP7_75t_L g420 ( .A1(n_252), .A2(n_404), .B1(n_421), .B2(n_424), .C(n_426), .Y(n_420) );
OR2x2_ASAP7_75t_L g252 ( .A(n_253), .B(n_254), .Y(n_252) );
INVx1_ASAP7_75t_L g291 ( .A(n_253), .Y(n_291) );
NAND2xp5_ASAP7_75t_L g343 ( .A(n_253), .B(n_302), .Y(n_343) );
NOR2xp33_ASAP7_75t_L g312 ( .A(n_254), .B(n_313), .Y(n_312) );
OR2x2_ASAP7_75t_L g345 ( .A(n_254), .B(n_291), .Y(n_345) );
INVx3_ASAP7_75t_SL g386 ( .A(n_254), .Y(n_386) );
AND2x2_ASAP7_75t_L g330 ( .A(n_255), .B(n_331), .Y(n_330) );
AND2x2_ASAP7_75t_L g359 ( .A(n_255), .B(n_360), .Y(n_359) );
NAND2xp5_ASAP7_75t_L g374 ( .A(n_255), .B(n_268), .Y(n_374) );
NAND2xp5_ASAP7_75t_L g400 ( .A(n_255), .B(n_314), .Y(n_400) );
INVx3_ASAP7_75t_L g255 ( .A(n_256), .Y(n_255) );
INVx3_ASAP7_75t_L g302 ( .A(n_256), .Y(n_302) );
OAI322xp33_ASAP7_75t_L g397 ( .A1(n_256), .A2(n_328), .A3(n_350), .B1(n_398), .B2(n_400), .C1(n_401), .C2(n_402), .Y(n_397) );
INVx1_ASAP7_75t_L g266 ( .A(n_267), .Y(n_266) );
AOI21xp33_ASAP7_75t_L g421 ( .A1(n_267), .A2(n_270), .B(n_422), .Y(n_421) );
NOR2xp33_ASAP7_75t_SL g347 ( .A(n_268), .B(n_348), .Y(n_347) );
AND2x2_ASAP7_75t_L g369 ( .A(n_268), .B(n_281), .Y(n_369) );
NAND2xp5_ASAP7_75t_L g384 ( .A(n_268), .B(n_308), .Y(n_384) );
INVxp67_ASAP7_75t_L g335 ( .A(n_270), .Y(n_335) );
AOI211xp5_ASAP7_75t_L g341 ( .A1(n_270), .A2(n_342), .B(n_346), .C(n_356), .Y(n_341) );
OAI221xp5_ASAP7_75t_SL g271 ( .A1(n_272), .A2(n_280), .B1(n_283), .B2(n_287), .C(n_292), .Y(n_271) );
INVxp67_ASAP7_75t_L g272 ( .A(n_273), .Y(n_272) );
OR2x2_ASAP7_75t_L g274 ( .A(n_275), .B(n_278), .Y(n_274) );
INVx1_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
AND2x2_ASAP7_75t_L g295 ( .A(n_279), .B(n_296), .Y(n_295) );
INVx1_ASAP7_75t_L g412 ( .A(n_279), .Y(n_412) );
OAI221xp5_ASAP7_75t_L g428 ( .A1(n_280), .A2(n_429), .B1(n_434), .B2(n_435), .C(n_437), .Y(n_428) );
OR2x2_ASAP7_75t_L g280 ( .A(n_281), .B(n_282), .Y(n_280) );
NAND2xp5_ASAP7_75t_L g324 ( .A(n_281), .B(n_325), .Y(n_324) );
INVx1_ASAP7_75t_SL g328 ( .A(n_281), .Y(n_328) );
NAND2xp5_ASAP7_75t_L g366 ( .A(n_281), .B(n_359), .Y(n_366) );
AND2x2_ASAP7_75t_L g408 ( .A(n_281), .B(n_386), .Y(n_408) );
NOR2xp33_ASAP7_75t_L g306 ( .A(n_282), .B(n_307), .Y(n_306) );
OAI22xp33_ASAP7_75t_L g403 ( .A1(n_282), .A2(n_294), .B1(n_404), .B2(n_405), .Y(n_403) );
OR2x2_ASAP7_75t_L g434 ( .A(n_282), .B(n_302), .Y(n_434) );
CKINVDCx16_ASAP7_75t_R g283 ( .A(n_284), .Y(n_283) );
INVx1_ASAP7_75t_L g411 ( .A(n_285), .Y(n_411) );
AND2x2_ASAP7_75t_L g436 ( .A(n_285), .B(n_379), .Y(n_436) );
INVxp67_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
NOR2xp33_ASAP7_75t_SL g288 ( .A(n_289), .B(n_291), .Y(n_288) );
INVx1_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
OR2x2_ASAP7_75t_L g300 ( .A(n_290), .B(n_301), .Y(n_300) );
AOI22xp5_ASAP7_75t_L g292 ( .A1(n_293), .A2(n_299), .B1(n_303), .B2(n_306), .Y(n_292) );
INVx1_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
NAND2xp5_ASAP7_75t_L g294 ( .A(n_295), .B(n_297), .Y(n_294) );
INVx1_ASAP7_75t_L g367 ( .A(n_295), .Y(n_367) );
NAND2xp5_ASAP7_75t_L g402 ( .A(n_295), .B(n_335), .Y(n_402) );
AOI322xp5_ASAP7_75t_L g326 ( .A1(n_297), .A2(n_327), .A3(n_329), .B1(n_330), .B2(n_332), .C1(n_333), .C2(n_337), .Y(n_326) );
INVxp67_ASAP7_75t_L g320 ( .A(n_298), .Y(n_320) );
INVx1_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
OAI22xp5_ASAP7_75t_L g321 ( .A1(n_300), .A2(n_305), .B1(n_322), .B2(n_324), .Y(n_321) );
NAND2xp5_ASAP7_75t_L g401 ( .A(n_301), .B(n_314), .Y(n_401) );
INVx1_ASAP7_75t_SL g301 ( .A(n_302), .Y(n_301) );
NOR2xp33_ASAP7_75t_L g410 ( .A(n_302), .B(n_340), .Y(n_410) );
NOR2xp33_ASAP7_75t_L g416 ( .A(n_302), .B(n_417), .Y(n_416) );
INVx1_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
OR2x2_ASAP7_75t_L g398 ( .A(n_304), .B(n_399), .Y(n_398) );
INVx1_ASAP7_75t_SL g307 ( .A(n_308), .Y(n_307) );
NAND3xp33_ASAP7_75t_SL g309 ( .A(n_310), .B(n_326), .C(n_341), .Y(n_309) );
AOI221xp5_ASAP7_75t_L g310 ( .A1(n_311), .A2(n_312), .B1(n_317), .B2(n_319), .C(n_321), .Y(n_310) );
AND2x2_ASAP7_75t_L g317 ( .A(n_313), .B(n_318), .Y(n_317) );
INVx3_ASAP7_75t_SL g313 ( .A(n_314), .Y(n_313) );
AND2x4_ASAP7_75t_L g314 ( .A(n_315), .B(n_316), .Y(n_314) );
AND2x2_ASAP7_75t_L g327 ( .A(n_318), .B(n_328), .Y(n_327) );
HB1xp67_ASAP7_75t_L g399 ( .A(n_320), .Y(n_399) );
INVx1_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
NAND2xp5_ASAP7_75t_L g355 ( .A(n_325), .B(n_339), .Y(n_355) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_328), .B(n_386), .Y(n_392) );
NOR2xp33_ASAP7_75t_L g388 ( .A(n_329), .B(n_389), .Y(n_388) );
INVx1_ASAP7_75t_SL g404 ( .A(n_332), .Y(n_404) );
AND2x2_ASAP7_75t_L g419 ( .A(n_332), .B(n_396), .Y(n_419) );
INVx1_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
NAND2xp5_ASAP7_75t_L g334 ( .A(n_335), .B(n_336), .Y(n_334) );
INVx1_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
AOI211xp5_ASAP7_75t_L g413 ( .A1(n_343), .A2(n_414), .B(n_420), .C(n_428), .Y(n_413) );
INVx1_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
OR2x2_ASAP7_75t_L g350 ( .A(n_351), .B(n_352), .Y(n_350) );
INVx1_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
AND2x2_ASAP7_75t_L g382 ( .A(n_353), .B(n_383), .Y(n_382) );
NAND2x1_ASAP7_75t_SL g424 ( .A(n_354), .B(n_425), .Y(n_424) );
CKINVDCx16_ASAP7_75t_R g394 ( .A(n_357), .Y(n_394) );
INVx1_ASAP7_75t_SL g358 ( .A(n_359), .Y(n_358) );
INVx1_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
INVx1_ASAP7_75t_L g389 ( .A(n_363), .Y(n_389) );
AND2x2_ASAP7_75t_L g393 ( .A(n_363), .B(n_379), .Y(n_393) );
NOR5xp2_ASAP7_75t_L g364 ( .A(n_365), .B(n_380), .C(n_397), .D(n_403), .E(n_406), .Y(n_364) );
OAI221xp5_ASAP7_75t_L g365 ( .A1(n_366), .A2(n_367), .B1(n_368), .B2(n_370), .C(n_372), .Y(n_365) );
INVx2_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
NAND2xp5_ASAP7_75t_L g426 ( .A(n_369), .B(n_427), .Y(n_426) );
INVxp67_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_373), .B(n_375), .Y(n_372) );
INVx1_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
INVx1_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
NAND2xp5_ASAP7_75t_L g376 ( .A(n_377), .B(n_379), .Y(n_376) );
INVx1_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
AND2x2_ASAP7_75t_L g395 ( .A(n_379), .B(n_396), .Y(n_395) );
OAI221xp5_ASAP7_75t_SL g380 ( .A1(n_381), .A2(n_384), .B1(n_385), .B2(n_387), .C(n_390), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
INVx1_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
AOI22xp33_ASAP7_75t_L g390 ( .A1(n_391), .A2(n_393), .B1(n_394), .B2(n_395), .Y(n_390) );
INVx1_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
INVx1_ASAP7_75t_L g433 ( .A(n_393), .Y(n_433) );
AOI211xp5_ASAP7_75t_SL g406 ( .A1(n_407), .A2(n_409), .B(n_411), .C(n_412), .Y(n_406) );
INVx1_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
INVx1_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
INVx1_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
INVx1_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
INVx1_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
INVxp67_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
NAND2xp5_ASAP7_75t_L g430 ( .A(n_431), .B(n_433), .Y(n_430) );
INVx1_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
CKINVDCx14_ASAP7_75t_R g435 ( .A(n_436), .Y(n_435) );
INVx2_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
INVx2_ASAP7_75t_L g713 ( .A(n_443), .Y(n_713) );
OR2x2_ASAP7_75t_SL g443 ( .A(n_444), .B(n_665), .Y(n_443) );
NAND5xp2_ASAP7_75t_L g444 ( .A(n_445), .B(n_577), .C(n_615), .D(n_636), .E(n_653), .Y(n_444) );
NOR3xp33_ASAP7_75t_L g445 ( .A(n_446), .B(n_549), .C(n_570), .Y(n_445) );
OAI221xp5_ASAP7_75t_SL g446 ( .A1(n_447), .A2(n_489), .B1(n_512), .B2(n_536), .C(n_540), .Y(n_446) );
NAND2xp5_ASAP7_75t_L g447 ( .A(n_448), .B(n_460), .Y(n_447) );
INVx1_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
NAND2xp5_ASAP7_75t_L g557 ( .A(n_449), .B(n_538), .Y(n_557) );
OR2x2_ASAP7_75t_L g584 ( .A(n_449), .B(n_472), .Y(n_584) );
AND2x2_ASAP7_75t_L g598 ( .A(n_449), .B(n_472), .Y(n_598) );
NOR2xp33_ASAP7_75t_L g612 ( .A(n_449), .B(n_463), .Y(n_612) );
AND2x2_ASAP7_75t_L g650 ( .A(n_449), .B(n_614), .Y(n_650) );
AND2x2_ASAP7_75t_L g679 ( .A(n_449), .B(n_589), .Y(n_679) );
NAND2xp5_ASAP7_75t_L g696 ( .A(n_449), .B(n_561), .Y(n_696) );
INVx4_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
AND2x2_ASAP7_75t_L g576 ( .A(n_450), .B(n_471), .Y(n_576) );
BUFx3_ASAP7_75t_L g601 ( .A(n_450), .Y(n_601) );
AND2x2_ASAP7_75t_L g630 ( .A(n_450), .B(n_472), .Y(n_630) );
AND3x2_ASAP7_75t_L g643 ( .A(n_450), .B(n_644), .C(n_645), .Y(n_643) );
INVx1_ASAP7_75t_L g566 ( .A(n_460), .Y(n_566) );
AND2x2_ASAP7_75t_L g460 ( .A(n_461), .B(n_471), .Y(n_460) );
AOI32xp33_ASAP7_75t_L g621 ( .A1(n_461), .A2(n_573), .A3(n_622), .B1(n_625), .B2(n_626), .Y(n_621) );
INVx1_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
AND2x2_ASAP7_75t_L g548 ( .A(n_462), .B(n_471), .Y(n_548) );
NAND2xp5_ASAP7_75t_SL g619 ( .A(n_462), .B(n_576), .Y(n_619) );
AND2x2_ASAP7_75t_L g626 ( .A(n_462), .B(n_598), .Y(n_626) );
OR2x2_ASAP7_75t_L g632 ( .A(n_462), .B(n_633), .Y(n_632) );
NAND2xp5_ASAP7_75t_L g657 ( .A(n_462), .B(n_587), .Y(n_657) );
OR2x2_ASAP7_75t_L g675 ( .A(n_462), .B(n_500), .Y(n_675) );
BUFx3_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
AND2x2_ASAP7_75t_L g539 ( .A(n_463), .B(n_481), .Y(n_539) );
INVx2_ASAP7_75t_L g561 ( .A(n_463), .Y(n_561) );
OR2x2_ASAP7_75t_L g583 ( .A(n_463), .B(n_481), .Y(n_583) );
AND2x2_ASAP7_75t_L g588 ( .A(n_463), .B(n_589), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g639 ( .A(n_463), .B(n_640), .Y(n_639) );
AND2x2_ASAP7_75t_L g644 ( .A(n_463), .B(n_538), .Y(n_644) );
INVx1_ASAP7_75t_SL g695 ( .A(n_471), .Y(n_695) );
AND2x2_ASAP7_75t_L g471 ( .A(n_472), .B(n_481), .Y(n_471) );
INVx1_ASAP7_75t_SL g538 ( .A(n_472), .Y(n_538) );
HB1xp67_ASAP7_75t_L g587 ( .A(n_472), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g623 ( .A(n_472), .B(n_624), .Y(n_623) );
NAND3xp33_ASAP7_75t_L g690 ( .A(n_472), .B(n_561), .C(n_679), .Y(n_690) );
OA21x2_ASAP7_75t_L g472 ( .A1(n_473), .A2(n_474), .B(n_480), .Y(n_472) );
OA21x2_ASAP7_75t_L g481 ( .A1(n_473), .A2(n_482), .B(n_488), .Y(n_481) );
OA21x2_ASAP7_75t_L g491 ( .A1(n_473), .A2(n_492), .B(n_498), .Y(n_491) );
INVx2_ASAP7_75t_L g589 ( .A(n_481), .Y(n_589) );
HB1xp67_ASAP7_75t_L g603 ( .A(n_481), .Y(n_603) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_490), .B(n_499), .Y(n_489) );
INVx1_ASAP7_75t_L g625 ( .A(n_490), .Y(n_625) );
INVx1_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
AND2x2_ASAP7_75t_L g543 ( .A(n_491), .B(n_525), .Y(n_543) );
INVx2_ASAP7_75t_L g560 ( .A(n_491), .Y(n_560) );
AND2x2_ASAP7_75t_L g565 ( .A(n_491), .B(n_526), .Y(n_565) );
AND2x2_ASAP7_75t_L g580 ( .A(n_491), .B(n_513), .Y(n_580) );
AND2x2_ASAP7_75t_L g592 ( .A(n_491), .B(n_564), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g607 ( .A(n_499), .B(n_608), .Y(n_607) );
NAND2x1p5_ASAP7_75t_L g664 ( .A(n_499), .B(n_565), .Y(n_664) );
NAND2xp5_ASAP7_75t_L g683 ( .A(n_499), .B(n_684), .Y(n_683) );
NAND2xp5_ASAP7_75t_L g687 ( .A(n_499), .B(n_559), .Y(n_687) );
BUFx3_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
OR2x2_ASAP7_75t_L g524 ( .A(n_500), .B(n_525), .Y(n_524) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_500), .B(n_543), .Y(n_542) );
AND2x2_ASAP7_75t_L g569 ( .A(n_500), .B(n_513), .Y(n_569) );
AND2x2_ASAP7_75t_L g595 ( .A(n_500), .B(n_525), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g634 ( .A(n_500), .B(n_635), .Y(n_634) );
OA21x2_ASAP7_75t_L g500 ( .A1(n_501), .A2(n_502), .B(n_510), .Y(n_500) );
INVx1_ASAP7_75t_L g554 ( .A(n_502), .Y(n_554) );
NAND2xp5_ASAP7_75t_SL g505 ( .A(n_506), .B(n_509), .Y(n_505) );
INVx2_ASAP7_75t_L g520 ( .A(n_509), .Y(n_520) );
INVx1_ASAP7_75t_L g555 ( .A(n_510), .Y(n_555) );
OR2x2_ASAP7_75t_L g512 ( .A(n_513), .B(n_524), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_513), .B(n_546), .Y(n_545) );
AND2x4_ASAP7_75t_L g559 ( .A(n_513), .B(n_560), .Y(n_559) );
INVx3_ASAP7_75t_SL g564 ( .A(n_513), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g617 ( .A(n_513), .B(n_551), .Y(n_617) );
OR2x2_ASAP7_75t_L g627 ( .A(n_513), .B(n_553), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g655 ( .A(n_513), .B(n_595), .Y(n_655) );
OR2x2_ASAP7_75t_L g685 ( .A(n_513), .B(n_525), .Y(n_685) );
AND2x2_ASAP7_75t_L g689 ( .A(n_513), .B(n_526), .Y(n_689) );
NAND2xp5_ASAP7_75t_SL g702 ( .A(n_513), .B(n_565), .Y(n_702) );
AND2x2_ASAP7_75t_L g709 ( .A(n_513), .B(n_591), .Y(n_709) );
OR2x6_ASAP7_75t_L g513 ( .A(n_514), .B(n_522), .Y(n_513) );
INVx1_ASAP7_75t_SL g652 ( .A(n_524), .Y(n_652) );
AND2x2_ASAP7_75t_L g591 ( .A(n_525), .B(n_553), .Y(n_591) );
AND2x2_ASAP7_75t_L g605 ( .A(n_525), .B(n_560), .Y(n_605) );
AND2x2_ASAP7_75t_L g608 ( .A(n_525), .B(n_564), .Y(n_608) );
INVx1_ASAP7_75t_L g635 ( .A(n_525), .Y(n_635) );
INVx2_ASAP7_75t_SL g525 ( .A(n_526), .Y(n_525) );
BUFx2_ASAP7_75t_L g547 ( .A(n_526), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_537), .B(n_539), .Y(n_536) );
A2O1A1Ixp33_ASAP7_75t_L g706 ( .A1(n_537), .A2(n_583), .B(n_707), .C(n_708), .Y(n_706) );
HB1xp67_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
AND2x2_ASAP7_75t_L g613 ( .A(n_538), .B(n_614), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g571 ( .A(n_539), .B(n_556), .Y(n_571) );
AND2x2_ASAP7_75t_L g597 ( .A(n_539), .B(n_598), .Y(n_597) );
OAI21xp5_ASAP7_75t_SL g540 ( .A1(n_541), .A2(n_544), .B(n_548), .Y(n_540) );
INVx1_ASAP7_75t_L g541 ( .A(n_542), .Y(n_541) );
NOR2xp33_ASAP7_75t_L g641 ( .A(n_542), .B(n_642), .Y(n_641) );
AND2x2_ASAP7_75t_L g568 ( .A(n_543), .B(n_569), .Y(n_568) );
NAND2xp5_ASAP7_75t_L g609 ( .A(n_543), .B(n_564), .Y(n_609) );
AND2x2_ASAP7_75t_L g700 ( .A(n_543), .B(n_551), .Y(n_700) );
INVxp67_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
INVx1_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
AND2x2_ASAP7_75t_L g573 ( .A(n_547), .B(n_560), .Y(n_573) );
OR2x2_ASAP7_75t_L g574 ( .A(n_547), .B(n_558), .Y(n_574) );
OAI322xp33_ASAP7_75t_L g549 ( .A1(n_550), .A2(n_557), .A3(n_558), .B1(n_561), .B2(n_562), .C1(n_566), .C2(n_567), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g550 ( .A(n_551), .B(n_556), .Y(n_550) );
AND2x2_ASAP7_75t_L g661 ( .A(n_551), .B(n_573), .Y(n_661) );
NAND2xp5_ASAP7_75t_L g707 ( .A(n_551), .B(n_625), .Y(n_707) );
INVx2_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
INVx1_ASAP7_75t_SL g552 ( .A(n_553), .Y(n_552) );
AND2x2_ASAP7_75t_L g604 ( .A(n_553), .B(n_605), .Y(n_604) );
INVx1_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
OR2x2_ASAP7_75t_L g670 ( .A(n_557), .B(n_583), .Y(n_670) );
NAND2xp5_ASAP7_75t_L g651 ( .A(n_558), .B(n_652), .Y(n_651) );
INVx3_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g648 ( .A(n_559), .B(n_591), .Y(n_648) );
AND2x2_ASAP7_75t_L g594 ( .A(n_560), .B(n_564), .Y(n_594) );
AND2x2_ASAP7_75t_L g602 ( .A(n_561), .B(n_603), .Y(n_602) );
A2O1A1Ixp33_ASAP7_75t_L g699 ( .A1(n_561), .A2(n_640), .B(n_700), .C(n_701), .Y(n_699) );
AOI21xp33_ASAP7_75t_L g672 ( .A1(n_562), .A2(n_575), .B(n_673), .Y(n_672) );
INVx1_ASAP7_75t_SL g562 ( .A(n_563), .Y(n_562) );
AND2x2_ASAP7_75t_L g563 ( .A(n_564), .B(n_565), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g631 ( .A(n_564), .B(n_591), .Y(n_631) );
AND2x2_ASAP7_75t_L g637 ( .A(n_564), .B(n_605), .Y(n_637) );
AND2x2_ASAP7_75t_L g671 ( .A(n_564), .B(n_573), .Y(n_671) );
NOR2xp33_ASAP7_75t_L g579 ( .A(n_565), .B(n_580), .Y(n_579) );
INVx2_ASAP7_75t_SL g681 ( .A(n_565), .Y(n_681) );
INVx1_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
AOI22xp5_ASAP7_75t_L g596 ( .A1(n_569), .A2(n_597), .B1(n_599), .B2(n_604), .Y(n_596) );
OAI22xp5_ASAP7_75t_SL g570 ( .A1(n_571), .A2(n_572), .B1(n_574), .B2(n_575), .Y(n_570) );
OAI22xp33_ASAP7_75t_L g606 ( .A1(n_571), .A2(n_607), .B1(n_609), .B2(n_610), .Y(n_606) );
INVxp67_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
INVx1_ASAP7_75t_SL g575 ( .A(n_576), .Y(n_575) );
AOI221xp5_ASAP7_75t_L g677 ( .A1(n_576), .A2(n_678), .B1(n_680), .B2(n_682), .C(n_686), .Y(n_677) );
AOI211xp5_ASAP7_75t_L g577 ( .A1(n_578), .A2(n_581), .B(n_585), .C(n_606), .Y(n_577) );
INVxp67_ASAP7_75t_L g578 ( .A(n_579), .Y(n_578) );
INVx1_ASAP7_75t_L g581 ( .A(n_582), .Y(n_581) );
OR2x2_ASAP7_75t_L g582 ( .A(n_583), .B(n_584), .Y(n_582) );
OR2x2_ASAP7_75t_L g647 ( .A(n_583), .B(n_600), .Y(n_647) );
INVx1_ASAP7_75t_L g698 ( .A(n_583), .Y(n_698) );
OAI221xp5_ASAP7_75t_L g585 ( .A1(n_584), .A2(n_586), .B1(n_590), .B2(n_593), .C(n_596), .Y(n_585) );
INVx2_ASAP7_75t_SL g640 ( .A(n_584), .Y(n_640) );
NAND2xp5_ASAP7_75t_L g586 ( .A(n_587), .B(n_588), .Y(n_586) );
INVx1_ASAP7_75t_L g705 ( .A(n_587), .Y(n_705) );
AND2x2_ASAP7_75t_L g629 ( .A(n_588), .B(n_630), .Y(n_629) );
INVx2_ASAP7_75t_L g614 ( .A(n_589), .Y(n_614) );
NAND2xp5_ASAP7_75t_L g590 ( .A(n_591), .B(n_592), .Y(n_590) );
INVx1_ASAP7_75t_L g676 ( .A(n_592), .Y(n_676) );
NAND2xp5_ASAP7_75t_L g593 ( .A(n_594), .B(n_595), .Y(n_593) );
AND2x2_ASAP7_75t_L g599 ( .A(n_600), .B(n_602), .Y(n_599) );
NOR2xp33_ASAP7_75t_L g701 ( .A(n_600), .B(n_702), .Y(n_701) );
CKINVDCx16_ASAP7_75t_R g600 ( .A(n_601), .Y(n_600) );
INVxp67_ASAP7_75t_L g645 ( .A(n_603), .Y(n_645) );
O2A1O1Ixp33_ASAP7_75t_L g615 ( .A1(n_604), .A2(n_616), .B(n_618), .C(n_620), .Y(n_615) );
INVx1_ASAP7_75t_L g693 ( .A(n_607), .Y(n_693) );
INVx1_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
NOR2xp33_ASAP7_75t_L g668 ( .A(n_611), .B(n_669), .Y(n_668) );
AND2x2_ASAP7_75t_L g611 ( .A(n_612), .B(n_613), .Y(n_611) );
INVx2_ASAP7_75t_L g624 ( .A(n_614), .Y(n_624) );
INVx1_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
INVx1_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
OAI222xp33_ASAP7_75t_L g620 ( .A1(n_621), .A2(n_627), .B1(n_628), .B2(n_631), .C1(n_632), .C2(n_634), .Y(n_620) );
INVx1_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
INVx1_ASAP7_75t_SL g660 ( .A(n_624), .Y(n_660) );
NOR2xp33_ASAP7_75t_L g680 ( .A(n_627), .B(n_681), .Y(n_680) );
NAND2xp33_ASAP7_75t_SL g658 ( .A(n_628), .B(n_659), .Y(n_658) );
INVx1_ASAP7_75t_SL g628 ( .A(n_629), .Y(n_628) );
INVx1_ASAP7_75t_SL g633 ( .A(n_630), .Y(n_633) );
AND2x2_ASAP7_75t_L g697 ( .A(n_630), .B(n_698), .Y(n_697) );
OR2x2_ASAP7_75t_L g663 ( .A(n_633), .B(n_660), .Y(n_663) );
INVx1_ASAP7_75t_L g692 ( .A(n_634), .Y(n_692) );
AOI211xp5_ASAP7_75t_L g636 ( .A1(n_637), .A2(n_638), .B(n_641), .C(n_646), .Y(n_636) );
INVx1_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
NAND2xp5_ASAP7_75t_L g659 ( .A(n_640), .B(n_660), .Y(n_659) );
INVx2_ASAP7_75t_SL g642 ( .A(n_643), .Y(n_642) );
AOI322xp5_ASAP7_75t_L g691 ( .A1(n_643), .A2(n_671), .A3(n_676), .B1(n_692), .B2(n_693), .C1(n_694), .C2(n_697), .Y(n_691) );
AND2x2_ASAP7_75t_L g678 ( .A(n_644), .B(n_679), .Y(n_678) );
OAI22xp33_ASAP7_75t_L g646 ( .A1(n_647), .A2(n_648), .B1(n_649), .B2(n_651), .Y(n_646) );
INVxp33_ASAP7_75t_L g649 ( .A(n_650), .Y(n_649) );
AOI221xp5_ASAP7_75t_L g653 ( .A1(n_654), .A2(n_656), .B1(n_658), .B2(n_661), .C(n_662), .Y(n_653) );
INVx1_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
INVx1_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
NOR2xp33_ASAP7_75t_L g662 ( .A(n_663), .B(n_664), .Y(n_662) );
NAND5xp2_ASAP7_75t_L g665 ( .A(n_666), .B(n_677), .C(n_691), .D(n_699), .E(n_703), .Y(n_665) );
AOI21xp5_ASAP7_75t_L g666 ( .A1(n_667), .A2(n_671), .B(n_672), .Y(n_666) );
INVxp67_ASAP7_75t_L g667 ( .A(n_668), .Y(n_667) );
INVx2_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
INVxp33_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
NOR2xp33_ASAP7_75t_L g674 ( .A(n_675), .B(n_676), .Y(n_674) );
A2O1A1Ixp33_ASAP7_75t_L g703 ( .A1(n_679), .A2(n_704), .B(n_705), .C(n_706), .Y(n_703) );
AOI31xp33_ASAP7_75t_L g686 ( .A1(n_681), .A2(n_687), .A3(n_688), .B(n_690), .Y(n_686) );
INVx1_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
INVx1_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
INVx1_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
NOR2xp33_ASAP7_75t_L g694 ( .A(n_695), .B(n_696), .Y(n_694) );
INVx1_ASAP7_75t_L g704 ( .A(n_702), .Y(n_704) );
INVx1_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
INVx1_ASAP7_75t_L g715 ( .A(n_710), .Y(n_715) );
INVx2_ASAP7_75t_L g714 ( .A(n_715), .Y(n_714) );
INVx1_ASAP7_75t_L g716 ( .A(n_717), .Y(n_716) );
INVx2_ASAP7_75t_L g717 ( .A(n_718), .Y(n_717) );
INVx1_ASAP7_75t_SL g723 ( .A(n_724), .Y(n_723) );
INVx2_ASAP7_75t_L g725 ( .A(n_726), .Y(n_725) );
endmodule