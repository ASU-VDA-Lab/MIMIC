module fake_jpeg_13140_n_243 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_243);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_243;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_127;
wire n_76;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_233;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_16),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_9),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_10),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_7),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

INVx11_ASAP7_75t_L g30 ( 
.A(n_16),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

BUFx8_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_7),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_4),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_1),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_19),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_39),
.Y(n_79)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_32),
.Y(n_40)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_40),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_19),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_41),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_19),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_42),
.Y(n_89)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_43),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_38),
.Y(n_44)
);

BUFx2_ASAP7_75t_L g68 ( 
.A(n_44),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_22),
.B(n_15),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_45),
.B(n_46),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_22),
.B(n_13),
.Y(n_46)
);

INVx13_ASAP7_75t_L g47 ( 
.A(n_32),
.Y(n_47)
);

BUFx12_ASAP7_75t_L g72 ( 
.A(n_47),
.Y(n_72)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_34),
.Y(n_48)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_48),
.Y(n_75)
);

CKINVDCx9p33_ASAP7_75t_R g49 ( 
.A(n_32),
.Y(n_49)
);

INVx11_ASAP7_75t_L g81 ( 
.A(n_49),
.Y(n_81)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_32),
.Y(n_50)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_50),
.Y(n_73)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_33),
.Y(n_51)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_51),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

BUFx2_ASAP7_75t_L g98 ( 
.A(n_52),
.Y(n_98)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_33),
.Y(n_53)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_53),
.Y(n_88)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_25),
.Y(n_54)
);

INVx5_ASAP7_75t_L g84 ( 
.A(n_54),
.Y(n_84)
);

CKINVDCx14_ASAP7_75t_R g55 ( 
.A(n_30),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_55),
.B(n_63),
.Y(n_82)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_33),
.Y(n_56)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_56),
.Y(n_85)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_33),
.Y(n_57)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_57),
.Y(n_74)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_58),
.Y(n_93)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_25),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_59),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_35),
.Y(n_60)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_60),
.Y(n_76)
);

INVx11_ASAP7_75t_L g61 ( 
.A(n_30),
.Y(n_61)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_61),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_35),
.Y(n_62)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_62),
.Y(n_71)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_26),
.B(n_0),
.Y(n_63)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_31),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_64),
.A2(n_29),
.B1(n_18),
.B2(n_31),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_63),
.A2(n_24),
.B1(n_21),
.B2(n_17),
.Y(n_66)
);

CKINVDCx16_ASAP7_75t_R g114 ( 
.A(n_66),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_60),
.A2(n_35),
.B1(n_24),
.B2(n_21),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_70),
.A2(n_78),
.B1(n_92),
.B2(n_94),
.Y(n_99)
);

OAI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_43),
.A2(n_18),
.B1(n_17),
.B2(n_28),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_53),
.B(n_28),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_80),
.B(n_95),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_83),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_62),
.A2(n_37),
.B1(n_27),
.B2(n_23),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_L g101 ( 
.A1(n_87),
.A2(n_50),
.B1(n_40),
.B2(n_52),
.Y(n_101)
);

OR2x2_ASAP7_75t_L g91 ( 
.A(n_49),
.B(n_26),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_91),
.B(n_59),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_L g92 ( 
.A1(n_39),
.A2(n_29),
.B1(n_37),
.B2(n_27),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_54),
.A2(n_29),
.B1(n_23),
.B2(n_20),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_61),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_41),
.A2(n_20),
.B1(n_36),
.B2(n_2),
.Y(n_97)
);

OAI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_97),
.A2(n_36),
.B1(n_1),
.B2(n_3),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_96),
.B(n_57),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_100),
.B(n_110),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_101),
.A2(n_115),
.B1(n_90),
.B2(n_10),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_67),
.B(n_44),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_102),
.B(n_125),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_79),
.Y(n_103)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_103),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_72),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_104),
.B(n_109),
.Y(n_148)
);

CKINVDCx14_ASAP7_75t_R g132 ( 
.A(n_106),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_91),
.A2(n_64),
.B1(n_47),
.B2(n_42),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_107),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_108),
.A2(n_84),
.B1(n_98),
.B2(n_68),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_72),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_82),
.B(n_13),
.Y(n_110)
);

AND2x2_ASAP7_75t_L g111 ( 
.A(n_75),
.B(n_0),
.Y(n_111)
);

INVx1_ASAP7_75t_SL g129 ( 
.A(n_111),
.Y(n_129)
);

AO22x1_ASAP7_75t_L g112 ( 
.A1(n_81),
.A2(n_0),
.B1(n_1),
.B2(n_5),
.Y(n_112)
);

AOI21xp5_ASAP7_75t_SL g137 ( 
.A1(n_112),
.A2(n_94),
.B(n_83),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_L g115 ( 
.A1(n_92),
.A2(n_6),
.B1(n_8),
.B2(n_9),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_93),
.Y(n_116)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_116),
.Y(n_136)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_74),
.Y(n_117)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_117),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_77),
.B(n_12),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_118),
.Y(n_143)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_71),
.Y(n_119)
);

AND2x2_ASAP7_75t_L g133 ( 
.A(n_119),
.B(n_120),
.Y(n_133)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_69),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_85),
.B(n_74),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_121),
.B(n_123),
.Y(n_150)
);

INVx4_ASAP7_75t_L g122 ( 
.A(n_88),
.Y(n_122)
);

INVx13_ASAP7_75t_L g145 ( 
.A(n_122),
.Y(n_145)
);

NAND3xp33_ASAP7_75t_L g123 ( 
.A(n_81),
.B(n_11),
.C(n_8),
.Y(n_123)
);

INVxp33_ASAP7_75t_L g124 ( 
.A(n_72),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_124),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_79),
.Y(n_125)
);

INVx5_ASAP7_75t_L g126 ( 
.A(n_65),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_126),
.B(n_128),
.Y(n_142)
);

AND2x2_ASAP7_75t_L g127 ( 
.A(n_73),
.B(n_6),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_127),
.B(n_65),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_86),
.Y(n_128)
);

AND2x2_ASAP7_75t_L g166 ( 
.A(n_137),
.B(n_147),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_105),
.A2(n_78),
.B1(n_89),
.B2(n_86),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_140),
.B(n_144),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_141),
.A2(n_149),
.B1(n_109),
.B2(n_104),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_111),
.B(n_76),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_111),
.B(n_76),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_146),
.B(n_151),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_L g149 ( 
.A1(n_105),
.A2(n_98),
.B1(n_68),
.B2(n_89),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_102),
.B(n_6),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_127),
.B(n_8),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_152),
.B(n_112),
.Y(n_157)
);

AO21x1_ASAP7_75t_L g173 ( 
.A1(n_153),
.A2(n_9),
.B(n_11),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g154 ( 
.A(n_129),
.B(n_99),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_154),
.B(n_162),
.C(n_165),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_132),
.B(n_113),
.Y(n_156)
);

INVxp67_ASAP7_75t_L g192 ( 
.A(n_156),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_157),
.B(n_158),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_148),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_136),
.Y(n_159)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_159),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_131),
.B(n_114),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_160),
.B(n_164),
.Y(n_183)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_136),
.Y(n_161)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_161),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_129),
.B(n_116),
.C(n_120),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_133),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_135),
.B(n_134),
.C(n_147),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_137),
.A2(n_119),
.B1(n_128),
.B2(n_103),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_167),
.B(n_170),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_133),
.Y(n_168)
);

OAI21xp33_ASAP7_75t_L g184 ( 
.A1(n_168),
.A2(n_146),
.B(n_139),
.Y(n_184)
);

CKINVDCx14_ASAP7_75t_R g191 ( 
.A(n_169),
.Y(n_191)
);

OAI22xp33_ASAP7_75t_SL g170 ( 
.A1(n_134),
.A2(n_112),
.B1(n_122),
.B2(n_124),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_135),
.A2(n_125),
.B1(n_127),
.B2(n_90),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_171),
.B(n_174),
.Y(n_177)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_133),
.Y(n_172)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_172),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_173),
.A2(n_141),
.B1(n_150),
.B2(n_152),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_143),
.B(n_117),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_142),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_175),
.B(n_168),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_178),
.B(n_188),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_SL g179 ( 
.A1(n_166),
.A2(n_139),
.B(n_144),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_179),
.B(n_189),
.Y(n_198)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_184),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_L g186 ( 
.A1(n_166),
.A2(n_140),
.B(n_151),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_186),
.B(n_171),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_SL g189 ( 
.A1(n_166),
.A2(n_165),
.B(n_158),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_154),
.B(n_142),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_190),
.B(n_162),
.C(n_163),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_193),
.B(n_205),
.C(n_187),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_181),
.B(n_143),
.Y(n_195)
);

OAI21x1_ASAP7_75t_L g213 ( 
.A1(n_195),
.A2(n_200),
.B(n_202),
.Y(n_213)
);

NAND3xp33_ASAP7_75t_L g196 ( 
.A(n_183),
.B(n_163),
.C(n_172),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_196),
.B(n_199),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_188),
.B(n_175),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_185),
.B(n_164),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_180),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_201),
.B(n_204),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_181),
.B(n_130),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_203),
.B(n_190),
.Y(n_208)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_180),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_187),
.B(n_155),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_182),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_206),
.A2(n_182),
.B1(n_161),
.B2(n_159),
.Y(n_207)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_207),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_208),
.B(n_209),
.C(n_211),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_205),
.B(n_189),
.C(n_192),
.Y(n_211)
);

O2A1O1Ixp33_ASAP7_75t_L g214 ( 
.A1(n_197),
.A2(n_176),
.B(n_191),
.C(n_177),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_L g224 ( 
.A1(n_214),
.A2(n_200),
.B(n_186),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_194),
.A2(n_191),
.B1(n_178),
.B2(n_167),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_L g217 ( 
.A1(n_215),
.A2(n_194),
.B1(n_176),
.B2(n_177),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_193),
.B(n_179),
.C(n_185),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_216),
.B(n_198),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_217),
.B(n_221),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_218),
.B(n_219),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_212),
.B(n_183),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_213),
.B(n_199),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_210),
.B(n_206),
.Y(n_223)
);

AOI21xp5_ASAP7_75t_L g226 ( 
.A1(n_223),
.A2(n_224),
.B(n_203),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_222),
.B(n_209),
.C(n_218),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_225),
.B(n_229),
.C(n_230),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_226),
.B(n_130),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_222),
.B(n_216),
.C(n_208),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_SL g230 ( 
.A(n_221),
.B(n_214),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_SL g232 ( 
.A1(n_227),
.A2(n_224),
.B(n_220),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_SL g236 ( 
.A(n_232),
.B(n_233),
.Y(n_236)
);

AOI21xp5_ASAP7_75t_L g233 ( 
.A1(n_228),
.A2(n_155),
.B(n_173),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_234),
.A2(n_228),
.B1(n_230),
.B2(n_153),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_235),
.B(n_237),
.Y(n_238)
);

NOR2x1_ASAP7_75t_R g237 ( 
.A(n_231),
.B(n_138),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_237),
.B(n_138),
.C(n_145),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_239),
.B(n_126),
.Y(n_240)
);

NOR3xp33_ASAP7_75t_L g241 ( 
.A(n_240),
.B(n_238),
.C(n_236),
.Y(n_241)
);

AOI21xp5_ASAP7_75t_SL g242 ( 
.A1(n_241),
.A2(n_145),
.B(n_11),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_242),
.B(n_145),
.Y(n_243)
);


endmodule