module fake_ariane_250_n_1761 (n_83, n_8, n_56, n_60, n_64, n_119, n_124, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_149, n_34, n_69, n_95, n_92, n_143, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_152, n_120, n_106, n_12, n_53, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_49, n_20, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_11, n_129, n_126, n_137, n_122, n_148, n_52, n_135, n_73, n_77, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_151, n_136, n_28, n_80, n_146, n_97, n_154, n_142, n_14, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_127, n_35, n_54, n_25, n_1761);

input n_83;
input n_8;
input n_56;
input n_60;
input n_64;
input n_119;
input n_124;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_149;
input n_34;
input n_69;
input n_95;
input n_92;
input n_143;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_152;
input n_120;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_52;
input n_135;
input n_73;
input n_77;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_151;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_154;
input n_142;
input n_14;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1761;

wire n_913;
wire n_1681;
wire n_1486;
wire n_1507;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_610;
wire n_245;
wire n_1713;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_187;
wire n_1463;
wire n_1238;
wire n_1515;
wire n_817;
wire n_924;
wire n_781;
wire n_1566;
wire n_189;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_524;
wire n_1214;
wire n_634;
wire n_1246;
wire n_1138;
wire n_214;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_232;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1457;
wire n_377;
wire n_1682;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_945;
wire n_958;
wire n_813;
wire n_419;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1184;
wire n_202;
wire n_1535;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1277;
wire n_1746;
wire n_829;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_672;
wire n_740;
wire n_1283;
wire n_167;
wire n_1736;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_242;
wire n_645;
wire n_331;
wire n_559;
wire n_495;
wire n_267;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_200;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_620;
wire n_1074;
wire n_859;
wire n_587;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_206;
wire n_352;
wire n_899;
wire n_1703;
wire n_611;
wire n_1295;
wire n_365;
wire n_238;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_192;
wire n_661;
wire n_1751;
wire n_300;
wire n_533;
wire n_438;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_376;
wire n_512;
wire n_1597;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1213;
wire n_237;
wire n_780;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_209;
wire n_490;
wire n_1461;
wire n_1391;
wire n_225;
wire n_1599;
wire n_1006;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_1594;
wire n_680;
wire n_287;
wire n_1716;
wire n_302;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_212;
wire n_444;
wire n_851;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_182;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_460;
wire n_1555;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_992;
wire n_966;
wire n_955;
wire n_1182;
wire n_794;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_179;
wire n_1292;
wire n_1178;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_306;
wire n_203;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_1717;
wire n_824;
wire n_428;
wire n_159;
wire n_892;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_990;
wire n_1623;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1680;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_1731;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_155;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_698;
wire n_1674;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_172;
wire n_1058;
wire n_347;
wire n_1042;
wire n_183;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_205;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_1728;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_348;
wire n_552;
wire n_670;
wire n_379;
wire n_162;
wire n_264;
wire n_441;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_1743;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_194;
wire n_1163;
wire n_186;
wire n_1384;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1648;
wire n_1413;
wire n_855;
wire n_158;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_647;
wire n_1423;
wire n_600;
wire n_481;
wire n_1053;
wire n_1609;
wire n_529;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_1105;
wire n_547;
wire n_439;
wire n_604;
wire n_677;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_699;
wire n_727;
wire n_301;
wire n_1726;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_325;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_163;
wire n_1693;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_221;
wire n_321;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_845;
wire n_888;
wire n_1649;
wire n_1677;
wire n_1297;
wire n_178;
wire n_551;
wire n_417;
wire n_1708;
wire n_343;
wire n_1222;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_534;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_451;
wire n_745;
wire n_1741;
wire n_1572;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_769;
wire n_1753;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_982;
wire n_915;
wire n_215;
wire n_1075;
wire n_454;
wire n_298;
wire n_1331;
wire n_1529;
wire n_1227;
wire n_655;
wire n_1734;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_509;
wire n_666;
wire n_1747;
wire n_430;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1338;
wire n_1342;
wire n_456;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_873;
wire n_1301;
wire n_1748;
wire n_1243;
wire n_1400;
wire n_342;
wire n_1466;
wire n_1513;
wire n_1527;
wire n_358;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1668;
wire n_1605;
wire n_1078;
wire n_266;
wire n_157;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_480;
wire n_1327;
wire n_1475;
wire n_211;
wire n_642;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_1757;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_1632;
wire n_474;
wire n_805;
wire n_295;
wire n_1658;
wire n_190;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_180;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1258;
wire n_197;
wire n_640;
wire n_463;
wire n_1476;
wire n_1524;
wire n_1733;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_283;
wire n_806;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_682;
wire n_1616;
wire n_819;
wire n_586;
wire n_1324;
wire n_1429;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1759;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_198;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_169;
wire n_1201;
wire n_1288;
wire n_173;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_1367;
wire n_166;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1023;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_467;
wire n_1511;
wire n_1422;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_168;
wire n_538;
wire n_1517;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_810;
wire n_1290;
wire n_181;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_414;
wire n_571;
wire n_1521;
wire n_1694;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_409;
wire n_171;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1444;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_1739;
wire n_161;
wire n_532;
wire n_763;
wire n_540;
wire n_216;
wire n_692;
wire n_984;
wire n_1687;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_1756;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_493;
wire n_1311;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1335;
wire n_1715;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_792;
wire n_1262;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1183;
wire n_1326;
wire n_981;
wire n_1110;
wire n_1758;
wire n_243;
wire n_1407;
wire n_185;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_164;
wire n_184;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_1054;
wire n_508;
wire n_1679;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_191;
wire n_978;
wire n_1011;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_170;
wire n_1536;
wire n_1471;
wire n_160;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_176;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_541;
wire n_499;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_1663;
wire n_1625;
wire n_318;
wire n_1458;
wire n_244;
wire n_679;
wire n_1630;
wire n_220;
wire n_663;
wire n_1720;
wire n_443;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_1735;
wire n_391;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_765;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_857;
wire n_898;
wire n_363;
wire n_1067;
wire n_968;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_1755;
wire n_1285;
wire n_193;
wire n_761;
wire n_733;
wire n_731;
wire n_336;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1106;
wire n_784;
wire n_648;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_701;
wire n_1003;
wire n_1125;
wire n_1710;
wire n_309;
wire n_1344;
wire n_1390;
wire n_401;
wire n_485;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_567;
wire n_369;
wire n_240;
wire n_1727;
wire n_1575;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_188;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_1696;
wire n_498;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1497;
wire n_459;
wire n_1136;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1316;
wire n_175;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_709;
wire n_809;
wire n_1686;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_199;
wire n_217;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_308;
wire n_1223;
wire n_201;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_948;
wire n_922;
wire n_1004;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_196;
wire n_1337;
wire n_774;
wire n_933;
wire n_596;
wire n_954;
wire n_1168;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_664;
wire n_252;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1732;
wire n_415;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1126;
wire n_195;
wire n_938;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_946;
wire n_757;
wire n_375;
wire n_1655;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_265;
wire n_1583;
wire n_1604;
wire n_208;
wire n_1631;
wire n_1702;
wire n_156;
wire n_174;
wire n_275;
wire n_1375;
wire n_204;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_866;
wire n_246;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_165;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_1569;
wire n_289;
wire n_548;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_177;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1228;
wire n_1244;
wire n_411;
wire n_484;
wire n_849;
wire n_357;
wire n_412;
wire n_1251;
wire n_447;
wire n_1421;
wire n_1233;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

INVx1_ASAP7_75t_L g155 ( 
.A(n_150),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_105),
.Y(n_156)
);

INVx3_ASAP7_75t_L g157 ( 
.A(n_37),
.Y(n_157)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_135),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_15),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_88),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_79),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_35),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_104),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_96),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_72),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_8),
.Y(n_166)
);

CKINVDCx16_ASAP7_75t_R g167 ( 
.A(n_12),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_127),
.Y(n_168)
);

CKINVDCx16_ASAP7_75t_R g169 ( 
.A(n_37),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_61),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_129),
.Y(n_171)
);

INVxp67_ASAP7_75t_SL g172 ( 
.A(n_66),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_149),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_20),
.Y(n_174)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_131),
.Y(n_175)
);

BUFx3_ASAP7_75t_L g176 ( 
.A(n_45),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_121),
.Y(n_177)
);

INVx1_ASAP7_75t_SL g178 ( 
.A(n_77),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_12),
.Y(n_179)
);

CKINVDCx16_ASAP7_75t_R g180 ( 
.A(n_94),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_143),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_0),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_84),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_69),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_95),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_32),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_90),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_85),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_82),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_41),
.Y(n_190)
);

BUFx10_ASAP7_75t_L g191 ( 
.A(n_50),
.Y(n_191)
);

INVx1_ASAP7_75t_SL g192 ( 
.A(n_39),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_0),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_38),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_112),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_27),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_89),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_126),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_139),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_32),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_49),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_116),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_114),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_106),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_128),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_67),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_26),
.Y(n_207)
);

BUFx2_ASAP7_75t_L g208 ( 
.A(n_29),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_10),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_22),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_36),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_98),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_51),
.Y(n_213)
);

INVx2_ASAP7_75t_SL g214 ( 
.A(n_41),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_44),
.Y(n_215)
);

BUFx2_ASAP7_75t_SL g216 ( 
.A(n_130),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_53),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_47),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_70),
.Y(n_219)
);

CKINVDCx14_ASAP7_75t_R g220 ( 
.A(n_50),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_39),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_132),
.Y(n_222)
);

BUFx6f_ASAP7_75t_L g223 ( 
.A(n_15),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_29),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_33),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_87),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_6),
.Y(n_227)
);

BUFx6f_ASAP7_75t_L g228 ( 
.A(n_115),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_11),
.Y(n_229)
);

BUFx8_ASAP7_75t_SL g230 ( 
.A(n_99),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_2),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_2),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_65),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_75),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_26),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_137),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_81),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_59),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_117),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_57),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_147),
.Y(n_241)
);

INVx1_ASAP7_75t_SL g242 ( 
.A(n_20),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_101),
.Y(n_243)
);

CKINVDCx14_ASAP7_75t_R g244 ( 
.A(n_3),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_48),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_109),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_107),
.Y(n_247)
);

BUFx10_ASAP7_75t_L g248 ( 
.A(n_142),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_7),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_136),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_45),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_4),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_92),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_108),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_47),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_18),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_71),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_6),
.Y(n_258)
);

INVx1_ASAP7_75t_SL g259 ( 
.A(n_111),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_140),
.Y(n_260)
);

BUFx3_ASAP7_75t_L g261 ( 
.A(n_36),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_24),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_73),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_19),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_13),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_125),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_123),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_118),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_56),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_38),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_51),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_14),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_14),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_133),
.Y(n_274)
);

INVx1_ASAP7_75t_SL g275 ( 
.A(n_100),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_62),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_63),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_7),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_60),
.Y(n_279)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_35),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_22),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_93),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_16),
.Y(n_283)
);

BUFx3_ASAP7_75t_L g284 ( 
.A(n_31),
.Y(n_284)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_134),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_52),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_53),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_13),
.Y(n_288)
);

INVxp67_ASAP7_75t_L g289 ( 
.A(n_10),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_19),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_48),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_148),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_11),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_58),
.Y(n_294)
);

BUFx3_ASAP7_75t_L g295 ( 
.A(n_21),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_31),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_110),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_4),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_46),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_154),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_27),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_83),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_28),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_18),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_44),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_144),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_40),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_17),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_55),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_157),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_157),
.Y(n_311)
);

INVxp67_ASAP7_75t_SL g312 ( 
.A(n_157),
.Y(n_312)
);

NAND2xp33_ASAP7_75t_R g313 ( 
.A(n_160),
.B(n_64),
.Y(n_313)
);

OR2x2_ASAP7_75t_L g314 ( 
.A(n_208),
.B(n_1),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_230),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_171),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_183),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_155),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_155),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_156),
.Y(n_320)
);

HB1xp67_ASAP7_75t_L g321 ( 
.A(n_208),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_156),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_220),
.Y(n_323)
);

INVxp67_ASAP7_75t_L g324 ( 
.A(n_174),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_199),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_244),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_170),
.B(n_1),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_170),
.B(n_3),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_203),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_206),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_181),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_247),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_181),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_257),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_263),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_274),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_302),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_167),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_167),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_184),
.B(n_5),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_184),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_179),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_188),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g344 ( 
.A(n_215),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_188),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_197),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_197),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_198),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_198),
.Y(n_349)
);

CKINVDCx20_ASAP7_75t_R g350 ( 
.A(n_221),
.Y(n_350)
);

CKINVDCx20_ASAP7_75t_R g351 ( 
.A(n_286),
.Y(n_351)
);

INVxp67_ASAP7_75t_SL g352 ( 
.A(n_176),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_205),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_169),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_169),
.Y(n_355)
);

INVxp67_ASAP7_75t_L g356 ( 
.A(n_174),
.Y(n_356)
);

HB1xp67_ASAP7_75t_L g357 ( 
.A(n_176),
.Y(n_357)
);

CKINVDCx20_ASAP7_75t_R g358 ( 
.A(n_301),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_162),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g360 ( 
.A(n_180),
.Y(n_360)
);

INVxp33_ASAP7_75t_L g361 ( 
.A(n_193),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_205),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_212),
.B(n_5),
.Y(n_363)
);

INVx2_ASAP7_75t_L g364 ( 
.A(n_159),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_166),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_212),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_182),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_236),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_186),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_190),
.Y(n_370)
);

AND2x4_ASAP7_75t_L g371 ( 
.A(n_261),
.B(n_8),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_236),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_194),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_196),
.Y(n_374)
);

INVxp67_ASAP7_75t_L g375 ( 
.A(n_193),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_200),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_239),
.Y(n_377)
);

INVxp67_ASAP7_75t_L g378 ( 
.A(n_201),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_209),
.Y(n_379)
);

INVxp67_ASAP7_75t_L g380 ( 
.A(n_201),
.Y(n_380)
);

INVxp67_ASAP7_75t_L g381 ( 
.A(n_214),
.Y(n_381)
);

CKINVDCx6p67_ASAP7_75t_R g382 ( 
.A(n_323),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_364),
.Y(n_383)
);

INVx1_ASAP7_75t_SL g384 ( 
.A(n_360),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_364),
.Y(n_385)
);

INVx2_ASAP7_75t_L g386 ( 
.A(n_364),
.Y(n_386)
);

HB1xp67_ASAP7_75t_L g387 ( 
.A(n_338),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_318),
.Y(n_388)
);

INVx2_ASAP7_75t_L g389 ( 
.A(n_310),
.Y(n_389)
);

AND2x2_ASAP7_75t_L g390 ( 
.A(n_318),
.B(n_180),
.Y(n_390)
);

AND2x4_ASAP7_75t_L g391 ( 
.A(n_371),
.B(n_261),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_319),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_319),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_320),
.Y(n_394)
);

BUFx8_ASAP7_75t_L g395 ( 
.A(n_371),
.Y(n_395)
);

AND2x2_ASAP7_75t_SL g396 ( 
.A(n_371),
.B(n_158),
.Y(n_396)
);

AND2x2_ASAP7_75t_L g397 ( 
.A(n_320),
.B(n_284),
.Y(n_397)
);

AND2x2_ASAP7_75t_L g398 ( 
.A(n_322),
.B(n_284),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_322),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_316),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_331),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_312),
.B(n_239),
.Y(n_402)
);

AND2x2_ASAP7_75t_L g403 ( 
.A(n_331),
.B(n_295),
.Y(n_403)
);

AND2x2_ASAP7_75t_L g404 ( 
.A(n_333),
.B(n_295),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_310),
.B(n_241),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_333),
.Y(n_406)
);

BUFx6f_ASAP7_75t_L g407 ( 
.A(n_341),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_341),
.Y(n_408)
);

INVx2_ASAP7_75t_L g409 ( 
.A(n_311),
.Y(n_409)
);

OAI22xp5_ASAP7_75t_L g410 ( 
.A1(n_314),
.A2(n_192),
.B1(n_242),
.B2(n_214),
.Y(n_410)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_311),
.Y(n_411)
);

HB1xp67_ASAP7_75t_L g412 ( 
.A(n_339),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_343),
.Y(n_413)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_343),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_345),
.Y(n_415)
);

BUFx8_ASAP7_75t_L g416 ( 
.A(n_371),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_345),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_346),
.Y(n_418)
);

BUFx6f_ASAP7_75t_L g419 ( 
.A(n_346),
.Y(n_419)
);

AND2x2_ASAP7_75t_L g420 ( 
.A(n_347),
.B(n_280),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_347),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_348),
.Y(n_422)
);

NOR2xp33_ASAP7_75t_L g423 ( 
.A(n_352),
.B(n_241),
.Y(n_423)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_348),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_349),
.Y(n_425)
);

INVx2_ASAP7_75t_L g426 ( 
.A(n_349),
.Y(n_426)
);

BUFx3_ASAP7_75t_L g427 ( 
.A(n_353),
.Y(n_427)
);

INVx4_ASAP7_75t_L g428 ( 
.A(n_353),
.Y(n_428)
);

BUFx6f_ASAP7_75t_L g429 ( 
.A(n_362),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_362),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_366),
.B(n_368),
.Y(n_431)
);

INVx6_ASAP7_75t_L g432 ( 
.A(n_314),
.Y(n_432)
);

INVx2_ASAP7_75t_L g433 ( 
.A(n_366),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_368),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_372),
.Y(n_435)
);

BUFx6f_ASAP7_75t_L g436 ( 
.A(n_372),
.Y(n_436)
);

INVx2_ASAP7_75t_L g437 ( 
.A(n_377),
.Y(n_437)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_377),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_328),
.Y(n_439)
);

INVx2_ASAP7_75t_L g440 ( 
.A(n_328),
.Y(n_440)
);

AND2x2_ASAP7_75t_L g441 ( 
.A(n_361),
.B(n_280),
.Y(n_441)
);

INVx2_ASAP7_75t_L g442 ( 
.A(n_327),
.Y(n_442)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_340),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_363),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_324),
.Y(n_445)
);

NAND2xp33_ASAP7_75t_R g446 ( 
.A(n_354),
.B(n_210),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_SL g447 ( 
.A(n_395),
.B(n_359),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_SL g448 ( 
.A(n_395),
.B(n_365),
.Y(n_448)
);

INVx2_ASAP7_75t_L g449 ( 
.A(n_386),
.Y(n_449)
);

AND2x2_ASAP7_75t_L g450 ( 
.A(n_390),
.B(n_357),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_407),
.Y(n_451)
);

INVx2_ASAP7_75t_L g452 ( 
.A(n_386),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_SL g453 ( 
.A(n_395),
.B(n_367),
.Y(n_453)
);

INVxp67_ASAP7_75t_SL g454 ( 
.A(n_395),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_407),
.Y(n_455)
);

NAND2xp33_ASAP7_75t_L g456 ( 
.A(n_439),
.B(n_369),
.Y(n_456)
);

INVx3_ASAP7_75t_L g457 ( 
.A(n_407),
.Y(n_457)
);

INVx2_ASAP7_75t_L g458 ( 
.A(n_386),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_SL g459 ( 
.A(n_395),
.B(n_370),
.Y(n_459)
);

INVxp33_ASAP7_75t_L g460 ( 
.A(n_387),
.Y(n_460)
);

INVx2_ASAP7_75t_SL g461 ( 
.A(n_395),
.Y(n_461)
);

NOR2xp33_ASAP7_75t_L g462 ( 
.A(n_440),
.B(n_373),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_407),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_SL g464 ( 
.A(n_416),
.B(n_374),
.Y(n_464)
);

INVxp33_ASAP7_75t_L g465 ( 
.A(n_387),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_440),
.B(n_376),
.Y(n_466)
);

AOI22xp33_ASAP7_75t_L g467 ( 
.A1(n_396),
.A2(n_321),
.B1(n_227),
.B2(n_217),
.Y(n_467)
);

BUFx8_ASAP7_75t_SL g468 ( 
.A(n_400),
.Y(n_468)
);

BUFx3_ASAP7_75t_L g469 ( 
.A(n_427),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_SL g470 ( 
.A(n_416),
.B(n_379),
.Y(n_470)
);

INVx2_ASAP7_75t_L g471 ( 
.A(n_386),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_SL g472 ( 
.A(n_416),
.B(n_355),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_440),
.B(n_439),
.Y(n_473)
);

NAND2xp33_ASAP7_75t_L g474 ( 
.A(n_439),
.B(n_159),
.Y(n_474)
);

NOR2xp33_ASAP7_75t_L g475 ( 
.A(n_440),
.B(n_326),
.Y(n_475)
);

AND2x2_ASAP7_75t_L g476 ( 
.A(n_390),
.B(n_381),
.Y(n_476)
);

INVx3_ASAP7_75t_L g477 ( 
.A(n_407),
.Y(n_477)
);

NOR2xp33_ASAP7_75t_L g478 ( 
.A(n_442),
.B(n_381),
.Y(n_478)
);

INVx2_ASAP7_75t_L g479 ( 
.A(n_407),
.Y(n_479)
);

AOI22xp33_ASAP7_75t_L g480 ( 
.A1(n_396),
.A2(n_264),
.B1(n_207),
.B2(n_227),
.Y(n_480)
);

INVx2_ASAP7_75t_L g481 ( 
.A(n_407),
.Y(n_481)
);

INVx2_ASAP7_75t_L g482 ( 
.A(n_407),
.Y(n_482)
);

NAND3xp33_ASAP7_75t_L g483 ( 
.A(n_428),
.B(n_313),
.C(n_223),
.Y(n_483)
);

INVx5_ASAP7_75t_L g484 ( 
.A(n_407),
.Y(n_484)
);

INVx2_ASAP7_75t_L g485 ( 
.A(n_419),
.Y(n_485)
);

INVx2_ASAP7_75t_L g486 ( 
.A(n_419),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_442),
.B(n_356),
.Y(n_487)
);

INVx3_ASAP7_75t_L g488 ( 
.A(n_419),
.Y(n_488)
);

INVx2_ASAP7_75t_L g489 ( 
.A(n_419),
.Y(n_489)
);

INVxp67_ASAP7_75t_L g490 ( 
.A(n_446),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_442),
.B(n_375),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_419),
.Y(n_492)
);

INVx4_ASAP7_75t_SL g493 ( 
.A(n_419),
.Y(n_493)
);

INVx2_ASAP7_75t_L g494 ( 
.A(n_419),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_419),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_419),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_429),
.Y(n_497)
);

INVx4_ASAP7_75t_L g498 ( 
.A(n_429),
.Y(n_498)
);

INVx3_ASAP7_75t_L g499 ( 
.A(n_429),
.Y(n_499)
);

NAND3xp33_ASAP7_75t_L g500 ( 
.A(n_428),
.B(n_223),
.C(n_159),
.Y(n_500)
);

BUFx3_ASAP7_75t_L g501 ( 
.A(n_427),
.Y(n_501)
);

AND2x2_ASAP7_75t_L g502 ( 
.A(n_390),
.B(n_378),
.Y(n_502)
);

AND2x2_ASAP7_75t_L g503 ( 
.A(n_441),
.B(n_380),
.Y(n_503)
);

INVx2_ASAP7_75t_L g504 ( 
.A(n_429),
.Y(n_504)
);

INVx2_ASAP7_75t_L g505 ( 
.A(n_429),
.Y(n_505)
);

NOR2xp33_ASAP7_75t_L g506 ( 
.A(n_442),
.B(n_317),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_429),
.Y(n_507)
);

INVx5_ASAP7_75t_L g508 ( 
.A(n_429),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_SL g509 ( 
.A(n_416),
.B(n_315),
.Y(n_509)
);

AND3x2_ASAP7_75t_L g510 ( 
.A(n_412),
.B(n_289),
.C(n_217),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_429),
.Y(n_511)
);

BUFx3_ASAP7_75t_L g512 ( 
.A(n_427),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_429),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_436),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_436),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_443),
.B(n_444),
.Y(n_516)
);

INVx3_ASAP7_75t_L g517 ( 
.A(n_436),
.Y(n_517)
);

OAI22xp5_ASAP7_75t_L g518 ( 
.A1(n_432),
.A2(n_231),
.B1(n_262),
.B2(n_256),
.Y(n_518)
);

NOR2xp33_ASAP7_75t_L g519 ( 
.A(n_443),
.B(n_325),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_443),
.B(n_178),
.Y(n_520)
);

BUFx6f_ASAP7_75t_L g521 ( 
.A(n_436),
.Y(n_521)
);

INVx3_ASAP7_75t_L g522 ( 
.A(n_436),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_SL g523 ( 
.A(n_416),
.B(n_329),
.Y(n_523)
);

NAND3xp33_ASAP7_75t_L g524 ( 
.A(n_428),
.B(n_223),
.C(n_159),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_443),
.B(n_259),
.Y(n_525)
);

INVx3_ASAP7_75t_L g526 ( 
.A(n_436),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_436),
.Y(n_527)
);

INVx2_ASAP7_75t_L g528 ( 
.A(n_436),
.Y(n_528)
);

INVx2_ASAP7_75t_SL g529 ( 
.A(n_416),
.Y(n_529)
);

AOI22xp33_ASAP7_75t_L g530 ( 
.A1(n_396),
.A2(n_410),
.B1(n_444),
.B2(n_432),
.Y(n_530)
);

BUFx4f_ASAP7_75t_L g531 ( 
.A(n_396),
.Y(n_531)
);

INVx2_ASAP7_75t_L g532 ( 
.A(n_436),
.Y(n_532)
);

INVxp67_ASAP7_75t_SL g533 ( 
.A(n_431),
.Y(n_533)
);

CKINVDCx5p33_ASAP7_75t_R g534 ( 
.A(n_400),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_388),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_388),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_SL g537 ( 
.A(n_445),
.B(n_330),
.Y(n_537)
);

CKINVDCx6p67_ASAP7_75t_R g538 ( 
.A(n_382),
.Y(n_538)
);

INVx1_ASAP7_75t_SL g539 ( 
.A(n_384),
.Y(n_539)
);

INVx2_ASAP7_75t_L g540 ( 
.A(n_383),
.Y(n_540)
);

INVx4_ASAP7_75t_L g541 ( 
.A(n_428),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_388),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_SL g543 ( 
.A(n_445),
.B(n_332),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_392),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_392),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_392),
.Y(n_546)
);

INVx3_ASAP7_75t_L g547 ( 
.A(n_428),
.Y(n_547)
);

OR2x6_ASAP7_75t_L g548 ( 
.A(n_391),
.B(n_216),
.Y(n_548)
);

OR2x6_ASAP7_75t_L g549 ( 
.A(n_391),
.B(n_432),
.Y(n_549)
);

INVx2_ASAP7_75t_L g550 ( 
.A(n_383),
.Y(n_550)
);

INVx3_ASAP7_75t_L g551 ( 
.A(n_428),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_393),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_393),
.Y(n_553)
);

INVx2_ASAP7_75t_L g554 ( 
.A(n_383),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_393),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_394),
.Y(n_556)
);

INVx2_ASAP7_75t_L g557 ( 
.A(n_385),
.Y(n_557)
);

INVx4_ASAP7_75t_L g558 ( 
.A(n_427),
.Y(n_558)
);

AND2x2_ASAP7_75t_L g559 ( 
.A(n_441),
.B(n_191),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_SL g560 ( 
.A(n_445),
.B(n_334),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_394),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_SL g562 ( 
.A(n_441),
.B(n_335),
.Y(n_562)
);

INVx2_ASAP7_75t_SL g563 ( 
.A(n_432),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_394),
.Y(n_564)
);

INVxp33_ASAP7_75t_L g565 ( 
.A(n_412),
.Y(n_565)
);

OR2x6_ASAP7_75t_L g566 ( 
.A(n_391),
.B(n_216),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_399),
.Y(n_567)
);

NOR2xp33_ASAP7_75t_L g568 ( 
.A(n_444),
.B(n_336),
.Y(n_568)
);

BUFx3_ASAP7_75t_L g569 ( 
.A(n_399),
.Y(n_569)
);

AOI22xp33_ASAP7_75t_L g570 ( 
.A1(n_410),
.A2(n_270),
.B1(n_278),
.B2(n_309),
.Y(n_570)
);

NOR2xp33_ASAP7_75t_L g571 ( 
.A(n_432),
.B(n_337),
.Y(n_571)
);

INVx2_ASAP7_75t_L g572 ( 
.A(n_385),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_385),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_399),
.Y(n_574)
);

BUFx3_ASAP7_75t_L g575 ( 
.A(n_401),
.Y(n_575)
);

AOI22xp33_ASAP7_75t_L g576 ( 
.A1(n_432),
.A2(n_229),
.B1(n_309),
.B2(n_287),
.Y(n_576)
);

BUFx3_ASAP7_75t_L g577 ( 
.A(n_401),
.Y(n_577)
);

INVx3_ASAP7_75t_L g578 ( 
.A(n_414),
.Y(n_578)
);

CKINVDCx5p33_ASAP7_75t_R g579 ( 
.A(n_382),
.Y(n_579)
);

BUFx6f_ASAP7_75t_L g580 ( 
.A(n_389),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_L g581 ( 
.A(n_391),
.B(n_275),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_401),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_SL g583 ( 
.A(n_423),
.B(n_402),
.Y(n_583)
);

INVx4_ASAP7_75t_L g584 ( 
.A(n_414),
.Y(n_584)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_414),
.Y(n_585)
);

BUFx3_ASAP7_75t_L g586 ( 
.A(n_406),
.Y(n_586)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_414),
.Y(n_587)
);

NAND2xp33_ASAP7_75t_L g588 ( 
.A(n_431),
.B(n_159),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_406),
.Y(n_589)
);

INVx2_ASAP7_75t_L g590 ( 
.A(n_424),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_406),
.Y(n_591)
);

INVx2_ASAP7_75t_SL g592 ( 
.A(n_432),
.Y(n_592)
);

AOI22xp33_ASAP7_75t_L g593 ( 
.A1(n_423),
.A2(n_287),
.B1(n_270),
.B2(n_245),
.Y(n_593)
);

OR2x6_ASAP7_75t_L g594 ( 
.A(n_391),
.B(n_207),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_L g595 ( 
.A(n_462),
.B(n_402),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_L g596 ( 
.A(n_533),
.B(n_391),
.Y(n_596)
);

AND2x2_ASAP7_75t_L g597 ( 
.A(n_503),
.B(n_384),
.Y(n_597)
);

INVx2_ASAP7_75t_L g598 ( 
.A(n_584),
.Y(n_598)
);

INVx2_ASAP7_75t_L g599 ( 
.A(n_584),
.Y(n_599)
);

AND2x2_ASAP7_75t_L g600 ( 
.A(n_503),
.B(n_382),
.Y(n_600)
);

INVx2_ASAP7_75t_SL g601 ( 
.A(n_539),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_569),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_L g603 ( 
.A(n_478),
.B(n_408),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_L g604 ( 
.A(n_506),
.B(n_408),
.Y(n_604)
);

BUFx5_ASAP7_75t_L g605 ( 
.A(n_451),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g606 ( 
.A(n_519),
.B(n_408),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_569),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_520),
.B(n_413),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_L g609 ( 
.A(n_525),
.B(n_413),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_L g610 ( 
.A(n_466),
.B(n_413),
.Y(n_610)
);

INVx2_ASAP7_75t_L g611 ( 
.A(n_584),
.Y(n_611)
);

AND2x2_ASAP7_75t_L g612 ( 
.A(n_502),
.B(n_382),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_569),
.Y(n_613)
);

AOI21xp5_ASAP7_75t_L g614 ( 
.A1(n_473),
.A2(n_516),
.B(n_583),
.Y(n_614)
);

AND2x2_ASAP7_75t_L g615 ( 
.A(n_502),
.B(n_397),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_575),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_L g617 ( 
.A(n_530),
.B(n_415),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_575),
.Y(n_618)
);

INVxp33_ASAP7_75t_L g619 ( 
.A(n_475),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_L g620 ( 
.A(n_487),
.B(n_415),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_L g621 ( 
.A(n_491),
.B(n_415),
.Y(n_621)
);

INVx3_ASAP7_75t_L g622 ( 
.A(n_469),
.Y(n_622)
);

INVx4_ASAP7_75t_L g623 ( 
.A(n_549),
.Y(n_623)
);

NOR2xp33_ASAP7_75t_L g624 ( 
.A(n_490),
.B(n_417),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_568),
.B(n_417),
.Y(n_625)
);

AND2x2_ASAP7_75t_L g626 ( 
.A(n_476),
.B(n_397),
.Y(n_626)
);

NOR2xp33_ASAP7_75t_R g627 ( 
.A(n_534),
.B(n_446),
.Y(n_627)
);

NAND2x1p5_ASAP7_75t_L g628 ( 
.A(n_531),
.B(n_461),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_SL g629 ( 
.A(n_531),
.B(n_417),
.Y(n_629)
);

AND2x2_ASAP7_75t_L g630 ( 
.A(n_476),
.B(n_397),
.Y(n_630)
);

BUFx6f_ASAP7_75t_L g631 ( 
.A(n_461),
.Y(n_631)
);

AND2x2_ASAP7_75t_L g632 ( 
.A(n_559),
.B(n_398),
.Y(n_632)
);

AOI22xp5_ASAP7_75t_L g633 ( 
.A1(n_531),
.A2(n_418),
.B1(n_421),
.B2(n_435),
.Y(n_633)
);

BUFx6f_ASAP7_75t_SL g634 ( 
.A(n_468),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_575),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_L g636 ( 
.A(n_559),
.B(n_418),
.Y(n_636)
);

HB1xp67_ASAP7_75t_L g637 ( 
.A(n_549),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_577),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_SL g639 ( 
.A(n_531),
.B(n_418),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_L g640 ( 
.A(n_577),
.B(n_421),
.Y(n_640)
);

OR2x2_ASAP7_75t_L g641 ( 
.A(n_450),
.B(n_398),
.Y(n_641)
);

INVx2_ASAP7_75t_SL g642 ( 
.A(n_450),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_L g643 ( 
.A(n_577),
.B(n_421),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_586),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_586),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_586),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_535),
.Y(n_647)
);

INVx3_ASAP7_75t_L g648 ( 
.A(n_469),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_480),
.B(n_422),
.Y(n_649)
);

OR2x2_ASAP7_75t_L g650 ( 
.A(n_460),
.B(n_398),
.Y(n_650)
);

INVx2_ASAP7_75t_L g651 ( 
.A(n_584),
.Y(n_651)
);

CKINVDCx5p33_ASAP7_75t_R g652 ( 
.A(n_538),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_535),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_L g654 ( 
.A(n_456),
.B(n_422),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_536),
.Y(n_655)
);

BUFx6f_ASAP7_75t_L g656 ( 
.A(n_529),
.Y(n_656)
);

INVx2_ASAP7_75t_L g657 ( 
.A(n_578),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_L g658 ( 
.A(n_563),
.B(n_422),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_536),
.Y(n_659)
);

AND2x4_ASAP7_75t_L g660 ( 
.A(n_549),
.B(n_398),
.Y(n_660)
);

NOR2xp67_ASAP7_75t_L g661 ( 
.A(n_579),
.B(n_424),
.Y(n_661)
);

NOR3xp33_ASAP7_75t_L g662 ( 
.A(n_571),
.B(n_235),
.C(n_229),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_SL g663 ( 
.A(n_529),
.B(n_425),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_563),
.B(n_592),
.Y(n_664)
);

AOI22xp5_ASAP7_75t_L g665 ( 
.A1(n_549),
.A2(n_425),
.B1(n_435),
.B2(n_434),
.Y(n_665)
);

INVx2_ASAP7_75t_L g666 ( 
.A(n_578),
.Y(n_666)
);

AND2x2_ASAP7_75t_L g667 ( 
.A(n_465),
.B(n_403),
.Y(n_667)
);

OAI221xp5_ASAP7_75t_L g668 ( 
.A1(n_593),
.A2(n_235),
.B1(n_245),
.B2(n_258),
.C(n_264),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_SL g669 ( 
.A(n_592),
.B(n_425),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_542),
.Y(n_670)
);

NOR2xp33_ASAP7_75t_L g671 ( 
.A(n_541),
.B(n_430),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_581),
.B(n_430),
.Y(n_672)
);

NOR2xp67_ASAP7_75t_L g673 ( 
.A(n_483),
.B(n_424),
.Y(n_673)
);

NOR2xp33_ASAP7_75t_L g674 ( 
.A(n_541),
.B(n_430),
.Y(n_674)
);

NOR3xp33_ASAP7_75t_L g675 ( 
.A(n_537),
.B(n_265),
.C(n_258),
.Y(n_675)
);

HB1xp67_ASAP7_75t_L g676 ( 
.A(n_549),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_547),
.B(n_434),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_L g678 ( 
.A(n_547),
.B(n_434),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_L g679 ( 
.A(n_547),
.B(n_435),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_542),
.Y(n_680)
);

AND2x2_ASAP7_75t_L g681 ( 
.A(n_565),
.B(n_403),
.Y(n_681)
);

AND2x2_ASAP7_75t_L g682 ( 
.A(n_538),
.B(n_403),
.Y(n_682)
);

OR2x6_ASAP7_75t_L g683 ( 
.A(n_594),
.B(n_420),
.Y(n_683)
);

AOI22xp5_ASAP7_75t_L g684 ( 
.A1(n_447),
.A2(n_420),
.B1(n_404),
.B2(n_403),
.Y(n_684)
);

AOI22x1_ASAP7_75t_L g685 ( 
.A1(n_544),
.A2(n_409),
.B1(n_389),
.B2(n_411),
.Y(n_685)
);

INVx2_ASAP7_75t_L g686 ( 
.A(n_578),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_547),
.B(n_551),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_SL g688 ( 
.A(n_541),
.B(n_424),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_L g689 ( 
.A(n_551),
.B(n_404),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_545),
.Y(n_690)
);

NOR3xp33_ASAP7_75t_L g691 ( 
.A(n_543),
.B(n_271),
.C(n_265),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_L g692 ( 
.A(n_551),
.B(n_404),
.Y(n_692)
);

AND2x4_ASAP7_75t_L g693 ( 
.A(n_594),
.B(n_404),
.Y(n_693)
);

NAND3xp33_ASAP7_75t_L g694 ( 
.A(n_518),
.B(n_405),
.C(n_426),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_551),
.B(n_467),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_L g696 ( 
.A(n_545),
.B(n_426),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_SL g697 ( 
.A(n_541),
.B(n_521),
.Y(n_697)
);

BUFx3_ASAP7_75t_L g698 ( 
.A(n_469),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_SL g699 ( 
.A(n_521),
.B(n_426),
.Y(n_699)
);

INVxp33_ASAP7_75t_L g700 ( 
.A(n_562),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_SL g701 ( 
.A(n_521),
.B(n_426),
.Y(n_701)
);

AND2x6_ASAP7_75t_SL g702 ( 
.A(n_594),
.B(n_271),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_L g703 ( 
.A(n_546),
.B(n_433),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_546),
.Y(n_704)
);

NOR2xp67_ASAP7_75t_L g705 ( 
.A(n_483),
.B(n_433),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_SL g706 ( 
.A(n_521),
.B(n_433),
.Y(n_706)
);

BUFx6f_ASAP7_75t_L g707 ( 
.A(n_580),
.Y(n_707)
);

CKINVDCx5p33_ASAP7_75t_R g708 ( 
.A(n_560),
.Y(n_708)
);

OR2x6_ASAP7_75t_L g709 ( 
.A(n_594),
.B(n_420),
.Y(n_709)
);

NOR3xp33_ASAP7_75t_L g710 ( 
.A(n_448),
.B(n_296),
.C(n_278),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_L g711 ( 
.A(n_552),
.B(n_553),
.Y(n_711)
);

INVx4_ASAP7_75t_L g712 ( 
.A(n_548),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_552),
.Y(n_713)
);

NOR2xp33_ASAP7_75t_L g714 ( 
.A(n_472),
.B(n_433),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_L g715 ( 
.A(n_553),
.B(n_437),
.Y(n_715)
);

INVx2_ASAP7_75t_L g716 ( 
.A(n_578),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_L g717 ( 
.A(n_555),
.B(n_437),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_L g718 ( 
.A(n_555),
.B(n_437),
.Y(n_718)
);

AOI22xp33_ASAP7_75t_L g719 ( 
.A1(n_570),
.A2(n_438),
.B1(n_437),
.B2(n_411),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_SL g720 ( 
.A(n_521),
.B(n_438),
.Y(n_720)
);

BUFx6f_ASAP7_75t_L g721 ( 
.A(n_580),
.Y(n_721)
);

NOR2xp33_ASAP7_75t_SL g722 ( 
.A(n_454),
.B(n_342),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_SL g723 ( 
.A(n_521),
.B(n_438),
.Y(n_723)
);

NAND3xp33_ASAP7_75t_L g724 ( 
.A(n_576),
.B(n_405),
.C(n_438),
.Y(n_724)
);

AOI22xp5_ASAP7_75t_L g725 ( 
.A1(n_453),
.A2(n_420),
.B1(n_172),
.B2(n_277),
.Y(n_725)
);

HB1xp67_ASAP7_75t_L g726 ( 
.A(n_594),
.Y(n_726)
);

NOR2xp33_ASAP7_75t_L g727 ( 
.A(n_558),
.B(n_389),
.Y(n_727)
);

AOI22xp33_ASAP7_75t_L g728 ( 
.A1(n_548),
.A2(n_411),
.B1(n_409),
.B2(n_389),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_556),
.Y(n_729)
);

NOR2xp33_ASAP7_75t_L g730 ( 
.A(n_558),
.B(n_409),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_556),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_561),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_L g733 ( 
.A(n_561),
.B(n_409),
.Y(n_733)
);

AND2x2_ASAP7_75t_L g734 ( 
.A(n_548),
.B(n_344),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_564),
.Y(n_735)
);

AND2x4_ASAP7_75t_L g736 ( 
.A(n_548),
.B(n_411),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_L g737 ( 
.A(n_564),
.B(n_254),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_567),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_567),
.B(n_254),
.Y(n_739)
);

INVx2_ASAP7_75t_L g740 ( 
.A(n_585),
.Y(n_740)
);

AOI22xp5_ASAP7_75t_L g741 ( 
.A1(n_459),
.A2(n_268),
.B1(n_277),
.B2(n_297),
.Y(n_741)
);

CKINVDCx16_ASAP7_75t_R g742 ( 
.A(n_548),
.Y(n_742)
);

AND2x2_ASAP7_75t_SL g743 ( 
.A(n_558),
.B(n_158),
.Y(n_743)
);

INVx3_ASAP7_75t_L g744 ( 
.A(n_501),
.Y(n_744)
);

BUFx2_ASAP7_75t_L g745 ( 
.A(n_566),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_574),
.Y(n_746)
);

OAI22xp5_ASAP7_75t_L g747 ( 
.A1(n_566),
.A2(n_211),
.B1(n_308),
.B2(n_307),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_574),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_SL g749 ( 
.A(n_558),
.B(n_268),
.Y(n_749)
);

AOI22xp5_ASAP7_75t_L g750 ( 
.A1(n_464),
.A2(n_297),
.B1(n_306),
.B2(n_226),
.Y(n_750)
);

NOR3xp33_ASAP7_75t_L g751 ( 
.A(n_470),
.B(n_509),
.C(n_523),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_582),
.Y(n_752)
);

INVx4_ASAP7_75t_L g753 ( 
.A(n_566),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_582),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_589),
.Y(n_755)
);

INVx2_ASAP7_75t_L g756 ( 
.A(n_587),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_589),
.B(n_296),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_L g758 ( 
.A(n_591),
.B(n_304),
.Y(n_758)
);

INVx1_ASAP7_75t_SL g759 ( 
.A(n_510),
.Y(n_759)
);

NOR2x1p5_ASAP7_75t_L g760 ( 
.A(n_500),
.B(n_213),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_SL g761 ( 
.A(n_580),
.B(n_175),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_SL g762 ( 
.A(n_580),
.B(n_175),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_SL g763 ( 
.A(n_580),
.B(n_285),
.Y(n_763)
);

OR2x2_ASAP7_75t_L g764 ( 
.A(n_597),
.B(n_350),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_L g765 ( 
.A(n_595),
.B(n_591),
.Y(n_765)
);

OAI21xp5_ASAP7_75t_L g766 ( 
.A1(n_614),
.A2(n_455),
.B(n_451),
.Y(n_766)
);

AOI21xp5_ASAP7_75t_L g767 ( 
.A1(n_687),
.A2(n_566),
.B(n_463),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_L g768 ( 
.A(n_625),
.B(n_501),
.Y(n_768)
);

AOI21xp5_ASAP7_75t_L g769 ( 
.A1(n_711),
.A2(n_566),
.B(n_463),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_647),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_604),
.B(n_587),
.Y(n_771)
);

AOI21xp5_ASAP7_75t_L g772 ( 
.A1(n_606),
.A2(n_492),
.B(n_455),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_610),
.B(n_587),
.Y(n_773)
);

AO21x1_ASAP7_75t_L g774 ( 
.A1(n_714),
.A2(n_498),
.B(n_495),
.Y(n_774)
);

BUFx12f_ASAP7_75t_L g775 ( 
.A(n_601),
.Y(n_775)
);

NOR3xp33_ASAP7_75t_L g776 ( 
.A(n_612),
.B(n_304),
.C(n_224),
.Y(n_776)
);

O2A1O1Ixp33_ASAP7_75t_L g777 ( 
.A1(n_596),
.A2(n_590),
.B(n_501),
.C(n_512),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_L g778 ( 
.A(n_624),
.B(n_590),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_653),
.Y(n_779)
);

INVx3_ASAP7_75t_L g780 ( 
.A(n_623),
.Y(n_780)
);

AND2x2_ASAP7_75t_L g781 ( 
.A(n_667),
.B(n_681),
.Y(n_781)
);

AOI21xp5_ASAP7_75t_L g782 ( 
.A1(n_671),
.A2(n_495),
.B(n_492),
.Y(n_782)
);

O2A1O1Ixp5_ASAP7_75t_SL g783 ( 
.A1(n_761),
.A2(n_497),
.B(n_515),
.C(n_514),
.Y(n_783)
);

OAI21xp33_ASAP7_75t_L g784 ( 
.A1(n_619),
.A2(n_627),
.B(n_636),
.Y(n_784)
);

O2A1O1Ixp33_ASAP7_75t_L g785 ( 
.A1(n_689),
.A2(n_590),
.B(n_512),
.C(n_474),
.Y(n_785)
);

OR2x6_ASAP7_75t_L g786 ( 
.A(n_623),
.B(n_512),
.Y(n_786)
);

O2A1O1Ixp33_ASAP7_75t_L g787 ( 
.A1(n_692),
.A2(n_540),
.B(n_573),
.C(n_572),
.Y(n_787)
);

CKINVDCx5p33_ASAP7_75t_R g788 ( 
.A(n_627),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_655),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_SL g790 ( 
.A(n_619),
.B(n_580),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_L g791 ( 
.A(n_632),
.B(n_624),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_659),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_L g793 ( 
.A(n_615),
.B(n_540),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_L g794 ( 
.A(n_626),
.B(n_540),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_SL g795 ( 
.A(n_660),
.B(n_498),
.Y(n_795)
);

NOR2xp33_ASAP7_75t_L g796 ( 
.A(n_700),
.B(n_351),
.Y(n_796)
);

CKINVDCx10_ASAP7_75t_R g797 ( 
.A(n_634),
.Y(n_797)
);

AOI21xp5_ASAP7_75t_L g798 ( 
.A1(n_671),
.A2(n_497),
.B(n_496),
.Y(n_798)
);

NOR2x1_ASAP7_75t_L g799 ( 
.A(n_661),
.B(n_498),
.Y(n_799)
);

BUFx2_ASAP7_75t_L g800 ( 
.A(n_600),
.Y(n_800)
);

BUFx6f_ASAP7_75t_L g801 ( 
.A(n_707),
.Y(n_801)
);

OAI22xp5_ASAP7_75t_L g802 ( 
.A1(n_743),
.A2(n_550),
.B1(n_573),
.B2(n_572),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_L g803 ( 
.A(n_630),
.B(n_550),
.Y(n_803)
);

OAI21xp5_ASAP7_75t_L g804 ( 
.A1(n_673),
.A2(n_507),
.B(n_496),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_SL g805 ( 
.A(n_660),
.B(n_743),
.Y(n_805)
);

AND2x4_ASAP7_75t_L g806 ( 
.A(n_660),
.B(n_493),
.Y(n_806)
);

AOI21xp33_ASAP7_75t_L g807 ( 
.A1(n_674),
.A2(n_588),
.B(n_554),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_SL g808 ( 
.A(n_693),
.B(n_498),
.Y(n_808)
);

INVxp67_ASAP7_75t_L g809 ( 
.A(n_650),
.Y(n_809)
);

NOR3xp33_ASAP7_75t_L g810 ( 
.A(n_642),
.B(n_225),
.C(n_218),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_670),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_L g812 ( 
.A(n_684),
.B(n_550),
.Y(n_812)
);

BUFx8_ASAP7_75t_SL g813 ( 
.A(n_634),
.Y(n_813)
);

BUFx4f_ASAP7_75t_L g814 ( 
.A(n_682),
.Y(n_814)
);

AND2x4_ASAP7_75t_L g815 ( 
.A(n_637),
.B(n_493),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_603),
.B(n_620),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_L g817 ( 
.A(n_621),
.B(n_554),
.Y(n_817)
);

AND2x2_ASAP7_75t_L g818 ( 
.A(n_641),
.B(n_358),
.Y(n_818)
);

OAI21xp5_ASAP7_75t_L g819 ( 
.A1(n_705),
.A2(n_511),
.B(n_507),
.Y(n_819)
);

BUFx3_ASAP7_75t_L g820 ( 
.A(n_652),
.Y(n_820)
);

NOR3xp33_ASAP7_75t_L g821 ( 
.A(n_747),
.B(n_668),
.C(n_662),
.Y(n_821)
);

A2O1A1Ixp33_ASAP7_75t_L g822 ( 
.A1(n_674),
.A2(n_573),
.B(n_572),
.C(n_557),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_680),
.Y(n_823)
);

AOI21xp5_ASAP7_75t_L g824 ( 
.A1(n_608),
.A2(n_513),
.B(n_511),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_L g825 ( 
.A(n_609),
.B(n_554),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_L g826 ( 
.A(n_693),
.B(n_557),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_L g827 ( 
.A(n_693),
.B(n_557),
.Y(n_827)
);

AND2x2_ASAP7_75t_L g828 ( 
.A(n_734),
.B(n_191),
.Y(n_828)
);

NOR2xp33_ASAP7_75t_L g829 ( 
.A(n_700),
.B(n_457),
.Y(n_829)
);

AND2x2_ASAP7_75t_L g830 ( 
.A(n_722),
.B(n_191),
.Y(n_830)
);

AOI21xp33_ASAP7_75t_L g831 ( 
.A1(n_617),
.A2(n_695),
.B(n_714),
.Y(n_831)
);

AOI22xp5_ASAP7_75t_L g832 ( 
.A1(n_637),
.A2(n_513),
.B1(n_514),
.B2(n_527),
.Y(n_832)
);

BUFx6f_ASAP7_75t_L g833 ( 
.A(n_707),
.Y(n_833)
);

AOI21xp5_ASAP7_75t_L g834 ( 
.A1(n_677),
.A2(n_515),
.B(n_527),
.Y(n_834)
);

BUFx6f_ASAP7_75t_L g835 ( 
.A(n_707),
.Y(n_835)
);

AOI21xp5_ASAP7_75t_L g836 ( 
.A1(n_678),
.A2(n_532),
.B(n_528),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_L g837 ( 
.A(n_672),
.B(n_676),
.Y(n_837)
);

AOI21xp5_ASAP7_75t_L g838 ( 
.A1(n_679),
.A2(n_532),
.B(n_528),
.Y(n_838)
);

AOI22xp5_ASAP7_75t_L g839 ( 
.A1(n_676),
.A2(n_499),
.B1(n_488),
.B2(n_526),
.Y(n_839)
);

BUFx6f_ASAP7_75t_L g840 ( 
.A(n_707),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_L g841 ( 
.A(n_690),
.B(n_457),
.Y(n_841)
);

INVx3_ASAP7_75t_L g842 ( 
.A(n_712),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_704),
.B(n_457),
.Y(n_843)
);

INVx3_ASAP7_75t_L g844 ( 
.A(n_712),
.Y(n_844)
);

OAI22xp5_ASAP7_75t_L g845 ( 
.A1(n_665),
.A2(n_713),
.B1(n_731),
.B2(n_729),
.Y(n_845)
);

AND2x2_ASAP7_75t_L g846 ( 
.A(n_708),
.B(n_191),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_L g847 ( 
.A(n_732),
.B(n_449),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_L g848 ( 
.A(n_735),
.B(n_449),
.Y(n_848)
);

AOI21xp5_ASAP7_75t_L g849 ( 
.A1(n_629),
.A2(n_532),
.B(n_528),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_738),
.B(n_449),
.Y(n_850)
);

BUFx12f_ASAP7_75t_L g851 ( 
.A(n_702),
.Y(n_851)
);

O2A1O1Ixp33_ASAP7_75t_L g852 ( 
.A1(n_629),
.A2(n_479),
.B(n_481),
.C(n_482),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_L g853 ( 
.A(n_746),
.B(n_748),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_752),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_754),
.Y(n_855)
);

AOI21xp5_ASAP7_75t_L g856 ( 
.A1(n_639),
.A2(n_479),
.B(n_481),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_755),
.B(n_452),
.Y(n_857)
);

AOI22xp5_ASAP7_75t_L g858 ( 
.A1(n_683),
.A2(n_526),
.B1(n_457),
.B2(n_522),
.Y(n_858)
);

AOI21xp5_ASAP7_75t_L g859 ( 
.A1(n_639),
.A2(n_479),
.B(n_481),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_SL g860 ( 
.A(n_726),
.B(n_477),
.Y(n_860)
);

INVx2_ASAP7_75t_L g861 ( 
.A(n_740),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_SL g862 ( 
.A(n_726),
.B(n_742),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_L g863 ( 
.A(n_657),
.B(n_452),
.Y(n_863)
);

AOI21xp5_ASAP7_75t_L g864 ( 
.A1(n_697),
.A2(n_482),
.B(n_486),
.Y(n_864)
);

INVxp33_ASAP7_75t_SL g865 ( 
.A(n_750),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_657),
.Y(n_866)
);

BUFx3_ASAP7_75t_L g867 ( 
.A(n_759),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_666),
.B(n_452),
.Y(n_868)
);

HB1xp67_ASAP7_75t_L g869 ( 
.A(n_683),
.Y(n_869)
);

INVx3_ASAP7_75t_L g870 ( 
.A(n_753),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_L g871 ( 
.A(n_666),
.B(n_458),
.Y(n_871)
);

INVx3_ASAP7_75t_L g872 ( 
.A(n_753),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_649),
.B(n_477),
.Y(n_873)
);

AND2x6_ASAP7_75t_L g874 ( 
.A(n_631),
.B(n_482),
.Y(n_874)
);

HB1xp67_ASAP7_75t_L g875 ( 
.A(n_683),
.Y(n_875)
);

AO21x1_ASAP7_75t_L g876 ( 
.A1(n_761),
.A2(n_504),
.B(n_486),
.Y(n_876)
);

CKINVDCx5p33_ASAP7_75t_R g877 ( 
.A(n_709),
.Y(n_877)
);

NOR2xp33_ASAP7_75t_L g878 ( 
.A(n_709),
.B(n_477),
.Y(n_878)
);

NOR2x1_ASAP7_75t_R g879 ( 
.A(n_745),
.B(n_232),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_686),
.Y(n_880)
);

INVx2_ASAP7_75t_L g881 ( 
.A(n_756),
.Y(n_881)
);

AOI22xp5_ASAP7_75t_L g882 ( 
.A1(n_709),
.A2(n_751),
.B1(n_710),
.B2(n_736),
.Y(n_882)
);

AOI21xp5_ASAP7_75t_L g883 ( 
.A1(n_697),
.A2(n_494),
.B(n_485),
.Y(n_883)
);

AOI21xp5_ASAP7_75t_L g884 ( 
.A1(n_688),
.A2(n_494),
.B(n_485),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_686),
.Y(n_885)
);

NOR2xp33_ASAP7_75t_L g886 ( 
.A(n_725),
.B(n_477),
.Y(n_886)
);

OAI22xp5_ASAP7_75t_L g887 ( 
.A1(n_633),
.A2(n_485),
.B1(n_486),
.B2(n_489),
.Y(n_887)
);

A2O1A1Ixp33_ASAP7_75t_L g888 ( 
.A1(n_654),
.A2(n_526),
.B(n_488),
.C(n_522),
.Y(n_888)
);

AOI21xp5_ASAP7_75t_L g889 ( 
.A1(n_688),
.A2(n_701),
.B(n_699),
.Y(n_889)
);

AOI22xp33_ASAP7_75t_L g890 ( 
.A1(n_736),
.A2(n_458),
.B1(n_471),
.B2(n_248),
.Y(n_890)
);

BUFx4f_ASAP7_75t_L g891 ( 
.A(n_631),
.Y(n_891)
);

AOI21xp5_ASAP7_75t_L g892 ( 
.A1(n_699),
.A2(n_505),
.B(n_494),
.Y(n_892)
);

AOI21xp5_ASAP7_75t_L g893 ( 
.A1(n_701),
.A2(n_505),
.B(n_504),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_L g894 ( 
.A(n_716),
.B(n_458),
.Y(n_894)
);

AO21x1_ASAP7_75t_L g895 ( 
.A1(n_762),
.A2(n_504),
.B(n_489),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_L g896 ( 
.A(n_716),
.B(n_471),
.Y(n_896)
);

AOI21xp5_ASAP7_75t_L g897 ( 
.A1(n_706),
.A2(n_489),
.B(n_505),
.Y(n_897)
);

NOR2xp33_ASAP7_75t_L g898 ( 
.A(n_602),
.B(n_488),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_L g899 ( 
.A(n_640),
.B(n_488),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_757),
.Y(n_900)
);

AOI21xp5_ASAP7_75t_L g901 ( 
.A1(n_706),
.A2(n_526),
.B(n_499),
.Y(n_901)
);

AOI21xp5_ASAP7_75t_L g902 ( 
.A1(n_720),
.A2(n_522),
.B(n_517),
.Y(n_902)
);

OAI22xp5_ASAP7_75t_L g903 ( 
.A1(n_728),
.A2(n_499),
.B1(n_522),
.B2(n_517),
.Y(n_903)
);

NOR2xp33_ASAP7_75t_L g904 ( 
.A(n_607),
.B(n_499),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_SL g905 ( 
.A(n_698),
.B(n_517),
.Y(n_905)
);

AOI21xp5_ASAP7_75t_L g906 ( 
.A1(n_720),
.A2(n_517),
.B(n_508),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_L g907 ( 
.A(n_643),
.B(n_471),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_758),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_696),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_703),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_L g911 ( 
.A(n_598),
.B(n_493),
.Y(n_911)
);

BUFx6f_ASAP7_75t_L g912 ( 
.A(n_721),
.Y(n_912)
);

AOI21xp5_ASAP7_75t_L g913 ( 
.A1(n_723),
.A2(n_508),
.B(n_484),
.Y(n_913)
);

O2A1O1Ixp5_ASAP7_75t_L g914 ( 
.A1(n_669),
.A2(n_524),
.B(n_500),
.C(n_285),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_L g915 ( 
.A(n_598),
.B(n_599),
.Y(n_915)
);

AND2x4_ASAP7_75t_SL g916 ( 
.A(n_631),
.B(n_248),
.Y(n_916)
);

AOI21xp5_ASAP7_75t_L g917 ( 
.A1(n_723),
.A2(n_508),
.B(n_484),
.Y(n_917)
);

NOR2x1p5_ASAP7_75t_SL g918 ( 
.A(n_605),
.B(n_493),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_SL g919 ( 
.A(n_698),
.B(n_493),
.Y(n_919)
);

BUFx6f_ASAP7_75t_L g920 ( 
.A(n_721),
.Y(n_920)
);

O2A1O1Ixp33_ASAP7_75t_L g921 ( 
.A1(n_669),
.A2(n_524),
.B(n_305),
.C(n_303),
.Y(n_921)
);

INVx5_ASAP7_75t_L g922 ( 
.A(n_631),
.Y(n_922)
);

AOI21xp5_ASAP7_75t_L g923 ( 
.A1(n_664),
.A2(n_508),
.B(n_484),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_L g924 ( 
.A(n_611),
.B(n_484),
.Y(n_924)
);

NOR2xp33_ASAP7_75t_L g925 ( 
.A(n_613),
.B(n_249),
.Y(n_925)
);

NOR3xp33_ASAP7_75t_L g926 ( 
.A(n_675),
.B(n_252),
.C(n_251),
.Y(n_926)
);

AOI21xp5_ASAP7_75t_L g927 ( 
.A1(n_715),
.A2(n_508),
.B(n_484),
.Y(n_927)
);

INVx2_ASAP7_75t_L g928 ( 
.A(n_651),
.Y(n_928)
);

INVx2_ASAP7_75t_L g929 ( 
.A(n_651),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_717),
.B(n_484),
.Y(n_930)
);

NOR2xp33_ASAP7_75t_L g931 ( 
.A(n_616),
.B(n_255),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_L g932 ( 
.A(n_718),
.B(n_508),
.Y(n_932)
);

INVx1_ASAP7_75t_SL g933 ( 
.A(n_737),
.Y(n_933)
);

AO21x1_ASAP7_75t_L g934 ( 
.A1(n_762),
.A2(n_248),
.B(n_228),
.Y(n_934)
);

AOI21xp5_ASAP7_75t_L g935 ( 
.A1(n_733),
.A2(n_164),
.B(n_294),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_L g936 ( 
.A(n_618),
.B(n_223),
.Y(n_936)
);

AO21x1_ASAP7_75t_L g937 ( 
.A1(n_763),
.A2(n_248),
.B(n_228),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_L g938 ( 
.A(n_635),
.B(n_223),
.Y(n_938)
);

AOI21xp5_ASAP7_75t_L g939 ( 
.A1(n_727),
.A2(n_161),
.B(n_292),
.Y(n_939)
);

AOI22xp5_ASAP7_75t_L g940 ( 
.A1(n_741),
.A2(n_290),
.B1(n_299),
.B2(n_298),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_L g941 ( 
.A(n_638),
.B(n_272),
.Y(n_941)
);

AOI21xp5_ASAP7_75t_L g942 ( 
.A1(n_727),
.A2(n_300),
.B(n_163),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_L g943 ( 
.A(n_644),
.B(n_645),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_L g944 ( 
.A(n_933),
.B(n_691),
.Y(n_944)
);

AND2x4_ASAP7_75t_L g945 ( 
.A(n_806),
.B(n_815),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_SL g946 ( 
.A(n_784),
.B(n_656),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_SL g947 ( 
.A(n_865),
.B(n_656),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_L g948 ( 
.A(n_791),
.B(n_719),
.Y(n_948)
);

AOI21xp5_ASAP7_75t_L g949 ( 
.A1(n_765),
.A2(n_730),
.B(n_658),
.Y(n_949)
);

AOI21xp5_ASAP7_75t_L g950 ( 
.A1(n_765),
.A2(n_730),
.B(n_663),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_770),
.Y(n_951)
);

AOI21xp5_ASAP7_75t_L g952 ( 
.A1(n_816),
.A2(n_663),
.B(n_721),
.Y(n_952)
);

INVx1_ASAP7_75t_SL g953 ( 
.A(n_800),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_L g954 ( 
.A(n_781),
.B(n_719),
.Y(n_954)
);

NOR2xp33_ASAP7_75t_L g955 ( 
.A(n_764),
.B(n_749),
.Y(n_955)
);

OAI22xp5_ASAP7_75t_L g956 ( 
.A1(n_853),
.A2(n_646),
.B1(n_728),
.B2(n_622),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_L g957 ( 
.A(n_837),
.B(n_739),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_SL g958 ( 
.A(n_788),
.B(n_814),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_779),
.Y(n_959)
);

AOI21xp33_ASAP7_75t_L g960 ( 
.A1(n_796),
.A2(n_749),
.B(n_724),
.Y(n_960)
);

INVx1_ASAP7_75t_SL g961 ( 
.A(n_867),
.Y(n_961)
);

BUFx5_ASAP7_75t_L g962 ( 
.A(n_874),
.Y(n_962)
);

INVx4_ASAP7_75t_L g963 ( 
.A(n_806),
.Y(n_963)
);

INVx1_ASAP7_75t_L g964 ( 
.A(n_789),
.Y(n_964)
);

BUFx2_ASAP7_75t_L g965 ( 
.A(n_775),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_792),
.Y(n_966)
);

OAI22xp5_ASAP7_75t_L g967 ( 
.A1(n_853),
.A2(n_694),
.B1(n_622),
.B2(n_744),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_811),
.Y(n_968)
);

AND2x2_ASAP7_75t_L g969 ( 
.A(n_818),
.B(n_760),
.Y(n_969)
);

BUFx6f_ASAP7_75t_L g970 ( 
.A(n_801),
.Y(n_970)
);

O2A1O1Ixp33_ASAP7_75t_L g971 ( 
.A1(n_821),
.A2(n_744),
.B(n_648),
.C(n_763),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_L g972 ( 
.A(n_900),
.B(n_908),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_SL g973 ( 
.A(n_891),
.B(n_656),
.Y(n_973)
);

BUFx6f_ASAP7_75t_L g974 ( 
.A(n_801),
.Y(n_974)
);

AOI21xp5_ASAP7_75t_L g975 ( 
.A1(n_771),
.A2(n_721),
.B(n_648),
.Y(n_975)
);

AOI21xp5_ASAP7_75t_L g976 ( 
.A1(n_771),
.A2(n_773),
.B(n_768),
.Y(n_976)
);

AOI22xp33_ASAP7_75t_L g977 ( 
.A1(n_828),
.A2(n_628),
.B1(n_291),
.B2(n_293),
.Y(n_977)
);

NOR2xp33_ASAP7_75t_R g978 ( 
.A(n_797),
.B(n_605),
.Y(n_978)
);

AOI21xp5_ASAP7_75t_L g979 ( 
.A1(n_773),
.A2(n_628),
.B(n_685),
.Y(n_979)
);

A2O1A1Ixp33_ASAP7_75t_SL g980 ( 
.A1(n_766),
.A2(n_605),
.B(n_288),
.C(n_283),
.Y(n_980)
);

INVxp67_ASAP7_75t_L g981 ( 
.A(n_846),
.Y(n_981)
);

AOI21xp5_ASAP7_75t_L g982 ( 
.A1(n_817),
.A2(n_605),
.B(n_282),
.Y(n_982)
);

BUFx6f_ASAP7_75t_L g983 ( 
.A(n_801),
.Y(n_983)
);

AOI21xp5_ASAP7_75t_L g984 ( 
.A1(n_778),
.A2(n_605),
.B(n_237),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_823),
.Y(n_985)
);

OAI22xp5_ASAP7_75t_SL g986 ( 
.A1(n_851),
.A2(n_273),
.B1(n_281),
.B2(n_187),
.Y(n_986)
);

INVx3_ASAP7_75t_L g987 ( 
.A(n_815),
.Y(n_987)
);

A2O1A1Ixp33_ASAP7_75t_L g988 ( 
.A1(n_769),
.A2(n_886),
.B(n_767),
.C(n_831),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_SL g989 ( 
.A(n_891),
.B(n_780),
.Y(n_989)
);

BUFx3_ASAP7_75t_L g990 ( 
.A(n_820),
.Y(n_990)
);

BUFx3_ASAP7_75t_L g991 ( 
.A(n_813),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_L g992 ( 
.A(n_809),
.B(n_605),
.Y(n_992)
);

BUFx8_ASAP7_75t_L g993 ( 
.A(n_830),
.Y(n_993)
);

AND2x2_ASAP7_75t_L g994 ( 
.A(n_877),
.B(n_869),
.Y(n_994)
);

O2A1O1Ixp33_ASAP7_75t_L g995 ( 
.A1(n_776),
.A2(n_9),
.B(n_16),
.C(n_17),
.Y(n_995)
);

AOI22xp33_ASAP7_75t_L g996 ( 
.A1(n_805),
.A2(n_875),
.B1(n_862),
.B2(n_926),
.Y(n_996)
);

OAI21x1_ASAP7_75t_L g997 ( 
.A1(n_892),
.A2(n_228),
.B(n_138),
.Y(n_997)
);

AOI22xp33_ASAP7_75t_L g998 ( 
.A1(n_940),
.A2(n_279),
.B1(n_276),
.B2(n_269),
.Y(n_998)
);

AOI21xp5_ASAP7_75t_L g999 ( 
.A1(n_778),
.A2(n_267),
.B(n_266),
.Y(n_999)
);

NOR2xp33_ASAP7_75t_L g1000 ( 
.A(n_829),
.B(n_260),
.Y(n_1000)
);

OR2x6_ASAP7_75t_SL g1001 ( 
.A(n_941),
.B(n_253),
.Y(n_1001)
);

NAND2xp33_ASAP7_75t_SL g1002 ( 
.A(n_793),
.B(n_794),
.Y(n_1002)
);

INVx1_ASAP7_75t_L g1003 ( 
.A(n_854),
.Y(n_1003)
);

OAI22xp5_ASAP7_75t_L g1004 ( 
.A1(n_845),
.A2(n_250),
.B1(n_246),
.B2(n_243),
.Y(n_1004)
);

NOR2xp33_ASAP7_75t_L g1005 ( 
.A(n_882),
.B(n_240),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_855),
.Y(n_1006)
);

OAI22x1_ASAP7_75t_L g1007 ( 
.A1(n_925),
.A2(n_238),
.B1(n_234),
.B2(n_233),
.Y(n_1007)
);

AOI21xp5_ASAP7_75t_L g1008 ( 
.A1(n_825),
.A2(n_189),
.B(n_222),
.Y(n_1008)
);

INVx3_ASAP7_75t_L g1009 ( 
.A(n_786),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_L g1010 ( 
.A(n_909),
.B(n_9),
.Y(n_1010)
);

NOR2xp33_ASAP7_75t_L g1011 ( 
.A(n_879),
.B(n_165),
.Y(n_1011)
);

NAND3xp33_ASAP7_75t_SL g1012 ( 
.A(n_810),
.B(n_168),
.C(n_173),
.Y(n_1012)
);

INVx1_ASAP7_75t_L g1013 ( 
.A(n_943),
.Y(n_1013)
);

OR2x2_ASAP7_75t_L g1014 ( 
.A(n_941),
.B(n_21),
.Y(n_1014)
);

AO21x1_ASAP7_75t_L g1015 ( 
.A1(n_802),
.A2(n_228),
.B(n_97),
.Y(n_1015)
);

HB1xp67_ASAP7_75t_L g1016 ( 
.A(n_826),
.Y(n_1016)
);

AND2x4_ASAP7_75t_L g1017 ( 
.A(n_780),
.B(n_786),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_L g1018 ( 
.A(n_910),
.B(n_23),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_L g1019 ( 
.A(n_803),
.B(n_23),
.Y(n_1019)
);

O2A1O1Ixp33_ASAP7_75t_L g1020 ( 
.A1(n_845),
.A2(n_24),
.B(n_25),
.C(n_28),
.Y(n_1020)
);

OAI22xp5_ASAP7_75t_L g1021 ( 
.A1(n_802),
.A2(n_219),
.B1(n_204),
.B2(n_202),
.Y(n_1021)
);

NAND2xp5_ASAP7_75t_L g1022 ( 
.A(n_827),
.B(n_931),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_L g1023 ( 
.A(n_916),
.B(n_25),
.Y(n_1023)
);

OAI22xp5_ASAP7_75t_L g1024 ( 
.A1(n_812),
.A2(n_195),
.B1(n_185),
.B2(n_177),
.Y(n_1024)
);

NAND3xp33_ASAP7_75t_L g1025 ( 
.A(n_822),
.B(n_228),
.C(n_33),
.Y(n_1025)
);

INVx4_ASAP7_75t_L g1026 ( 
.A(n_786),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_943),
.Y(n_1027)
);

O2A1O1Ixp33_ASAP7_75t_SL g1028 ( 
.A1(n_888),
.A2(n_30),
.B(n_34),
.C(n_40),
.Y(n_1028)
);

INVx3_ASAP7_75t_L g1029 ( 
.A(n_842),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_L g1030 ( 
.A(n_878),
.B(n_30),
.Y(n_1030)
);

INVx1_ASAP7_75t_L g1031 ( 
.A(n_866),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_L g1032 ( 
.A(n_831),
.B(n_34),
.Y(n_1032)
);

NAND2xp5_ASAP7_75t_SL g1033 ( 
.A(n_922),
.B(n_42),
.Y(n_1033)
);

INVx5_ASAP7_75t_L g1034 ( 
.A(n_874),
.Y(n_1034)
);

INVx1_ASAP7_75t_L g1035 ( 
.A(n_880),
.Y(n_1035)
);

NOR2xp33_ASAP7_75t_SL g1036 ( 
.A(n_922),
.B(n_42),
.Y(n_1036)
);

INVxp67_ASAP7_75t_L g1037 ( 
.A(n_860),
.Y(n_1037)
);

NAND2x1p5_ASAP7_75t_L g1038 ( 
.A(n_922),
.B(n_842),
.Y(n_1038)
);

AOI21xp5_ASAP7_75t_L g1039 ( 
.A1(n_782),
.A2(n_102),
.B(n_152),
.Y(n_1039)
);

A2O1A1Ixp33_ASAP7_75t_L g1040 ( 
.A1(n_807),
.A2(n_43),
.B(n_46),
.C(n_49),
.Y(n_1040)
);

AND2x4_ASAP7_75t_L g1041 ( 
.A(n_844),
.B(n_43),
.Y(n_1041)
);

O2A1O1Ixp33_ASAP7_75t_L g1042 ( 
.A1(n_807),
.A2(n_52),
.B(n_54),
.C(n_55),
.Y(n_1042)
);

A2O1A1Ixp33_ASAP7_75t_L g1043 ( 
.A1(n_777),
.A2(n_54),
.B(n_68),
.C(n_74),
.Y(n_1043)
);

NOR2xp33_ASAP7_75t_L g1044 ( 
.A(n_795),
.B(n_76),
.Y(n_1044)
);

BUFx12f_ASAP7_75t_L g1045 ( 
.A(n_833),
.Y(n_1045)
);

NOR2xp33_ASAP7_75t_L g1046 ( 
.A(n_808),
.B(n_78),
.Y(n_1046)
);

NOR2xp33_ASAP7_75t_SL g1047 ( 
.A(n_922),
.B(n_80),
.Y(n_1047)
);

INVx2_ASAP7_75t_L g1048 ( 
.A(n_861),
.Y(n_1048)
);

CKINVDCx20_ASAP7_75t_R g1049 ( 
.A(n_833),
.Y(n_1049)
);

NOR2xp33_ASAP7_75t_R g1050 ( 
.A(n_833),
.B(n_86),
.Y(n_1050)
);

A2O1A1Ixp33_ASAP7_75t_L g1051 ( 
.A1(n_787),
.A2(n_91),
.B(n_103),
.C(n_113),
.Y(n_1051)
);

AOI21xp5_ASAP7_75t_L g1052 ( 
.A1(n_798),
.A2(n_119),
.B(n_120),
.Y(n_1052)
);

AOI21xp5_ASAP7_75t_L g1053 ( 
.A1(n_907),
.A2(n_122),
.B(n_124),
.Y(n_1053)
);

NOR2xp33_ASAP7_75t_SL g1054 ( 
.A(n_874),
.B(n_141),
.Y(n_1054)
);

NOR3xp33_ASAP7_75t_L g1055 ( 
.A(n_790),
.B(n_145),
.C(n_146),
.Y(n_1055)
);

OA22x2_ASAP7_75t_L g1056 ( 
.A1(n_832),
.A2(n_151),
.B1(n_153),
.B2(n_885),
.Y(n_1056)
);

AOI21xp5_ASAP7_75t_L g1057 ( 
.A1(n_930),
.A2(n_932),
.B(n_772),
.Y(n_1057)
);

O2A1O1Ixp33_ASAP7_75t_L g1058 ( 
.A1(n_785),
.A2(n_857),
.B(n_850),
.C(n_848),
.Y(n_1058)
);

BUFx12f_ASAP7_75t_L g1059 ( 
.A(n_835),
.Y(n_1059)
);

BUFx6f_ASAP7_75t_L g1060 ( 
.A(n_840),
.Y(n_1060)
);

NAND2x1p5_ASAP7_75t_L g1061 ( 
.A(n_844),
.B(n_870),
.Y(n_1061)
);

OAI22xp5_ASAP7_75t_L g1062 ( 
.A1(n_858),
.A2(n_850),
.B1(n_857),
.B2(n_847),
.Y(n_1062)
);

AOI21xp5_ASAP7_75t_L g1063 ( 
.A1(n_930),
.A2(n_932),
.B(n_838),
.Y(n_1063)
);

BUFx6f_ASAP7_75t_L g1064 ( 
.A(n_840),
.Y(n_1064)
);

INVx1_ASAP7_75t_L g1065 ( 
.A(n_881),
.Y(n_1065)
);

OR2x6_ASAP7_75t_L g1066 ( 
.A(n_870),
.B(n_872),
.Y(n_1066)
);

NAND2xp5_ASAP7_75t_L g1067 ( 
.A(n_872),
.B(n_847),
.Y(n_1067)
);

INVx3_ASAP7_75t_L g1068 ( 
.A(n_840),
.Y(n_1068)
);

NAND2xp5_ASAP7_75t_L g1069 ( 
.A(n_848),
.B(n_928),
.Y(n_1069)
);

AOI22xp5_ASAP7_75t_L g1070 ( 
.A1(n_874),
.A2(n_839),
.B1(n_903),
.B2(n_890),
.Y(n_1070)
);

O2A1O1Ixp33_ASAP7_75t_L g1071 ( 
.A1(n_905),
.A2(n_903),
.B(n_843),
.C(n_841),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_SL g1072 ( 
.A(n_912),
.B(n_920),
.Y(n_1072)
);

OAI22x1_ASAP7_75t_L g1073 ( 
.A1(n_929),
.A2(n_919),
.B1(n_904),
.B2(n_898),
.Y(n_1073)
);

NOR2xp33_ASAP7_75t_L g1074 ( 
.A(n_912),
.B(n_920),
.Y(n_1074)
);

O2A1O1Ixp33_ASAP7_75t_L g1075 ( 
.A1(n_939),
.A2(n_942),
.B(n_887),
.C(n_889),
.Y(n_1075)
);

INVx4_ASAP7_75t_L g1076 ( 
.A(n_874),
.Y(n_1076)
);

INVx1_ASAP7_75t_L g1077 ( 
.A(n_936),
.Y(n_1077)
);

A2O1A1Ixp33_ASAP7_75t_L g1078 ( 
.A1(n_804),
.A2(n_819),
.B(n_921),
.C(n_918),
.Y(n_1078)
);

INVx1_ASAP7_75t_L g1079 ( 
.A(n_936),
.Y(n_1079)
);

OAI21xp5_ASAP7_75t_L g1080 ( 
.A1(n_783),
.A2(n_824),
.B(n_836),
.Y(n_1080)
);

AOI21xp5_ASAP7_75t_L g1081 ( 
.A1(n_915),
.A2(n_883),
.B(n_864),
.Y(n_1081)
);

NOR2xp67_ASAP7_75t_L g1082 ( 
.A(n_1034),
.B(n_1076),
.Y(n_1082)
);

AOI21xp5_ASAP7_75t_L g1083 ( 
.A1(n_976),
.A2(n_899),
.B(n_873),
.Y(n_1083)
);

AO31x2_ASAP7_75t_L g1084 ( 
.A1(n_988),
.A2(n_774),
.A3(n_895),
.B(n_876),
.Y(n_1084)
);

INVx2_ASAP7_75t_SL g1085 ( 
.A(n_990),
.Y(n_1085)
);

OAI21x1_ASAP7_75t_L g1086 ( 
.A1(n_1081),
.A2(n_893),
.B(n_897),
.Y(n_1086)
);

AOI21xp5_ASAP7_75t_L g1087 ( 
.A1(n_949),
.A2(n_834),
.B(n_887),
.Y(n_1087)
);

INVx1_ASAP7_75t_L g1088 ( 
.A(n_951),
.Y(n_1088)
);

NAND2xp5_ASAP7_75t_L g1089 ( 
.A(n_972),
.B(n_912),
.Y(n_1089)
);

NAND2xp33_ASAP7_75t_SL g1090 ( 
.A(n_978),
.B(n_920),
.Y(n_1090)
);

OAI22xp5_ASAP7_75t_L g1091 ( 
.A1(n_1022),
.A2(n_924),
.B1(n_896),
.B2(n_868),
.Y(n_1091)
);

NOR2xp67_ASAP7_75t_R g1092 ( 
.A(n_1034),
.B(n_799),
.Y(n_1092)
);

AOI221xp5_ASAP7_75t_SL g1093 ( 
.A1(n_1020),
.A2(n_1042),
.B1(n_1040),
.B2(n_995),
.C(n_1032),
.Y(n_1093)
);

NAND3xp33_ASAP7_75t_L g1094 ( 
.A(n_1025),
.B(n_938),
.C(n_935),
.Y(n_1094)
);

OAI21x1_ASAP7_75t_SL g1095 ( 
.A1(n_1015),
.A2(n_852),
.B(n_849),
.Y(n_1095)
);

INVx1_ASAP7_75t_L g1096 ( 
.A(n_959),
.Y(n_1096)
);

AOI221xp5_ASAP7_75t_L g1097 ( 
.A1(n_955),
.A2(n_938),
.B1(n_863),
.B2(n_868),
.C(n_871),
.Y(n_1097)
);

AND2x4_ASAP7_75t_L g1098 ( 
.A(n_945),
.B(n_863),
.Y(n_1098)
);

AOI22xp5_ASAP7_75t_L g1099 ( 
.A1(n_1005),
.A2(n_871),
.B1(n_894),
.B2(n_896),
.Y(n_1099)
);

INVxp67_ASAP7_75t_L g1100 ( 
.A(n_953),
.Y(n_1100)
);

OAI21x1_ASAP7_75t_L g1101 ( 
.A1(n_1063),
.A2(n_856),
.B(n_859),
.Y(n_1101)
);

AOI21xp5_ASAP7_75t_L g1102 ( 
.A1(n_1057),
.A2(n_894),
.B(n_911),
.Y(n_1102)
);

AOI22xp5_ASAP7_75t_L g1103 ( 
.A1(n_981),
.A2(n_934),
.B1(n_937),
.B2(n_884),
.Y(n_1103)
);

AOI21xp5_ASAP7_75t_L g1104 ( 
.A1(n_1002),
.A2(n_927),
.B(n_923),
.Y(n_1104)
);

OR2x2_ASAP7_75t_L g1105 ( 
.A(n_953),
.B(n_901),
.Y(n_1105)
);

AOI21xp5_ASAP7_75t_L g1106 ( 
.A1(n_1062),
.A2(n_902),
.B(n_906),
.Y(n_1106)
);

AO31x2_ASAP7_75t_L g1107 ( 
.A1(n_1078),
.A2(n_913),
.A3(n_917),
.B(n_914),
.Y(n_1107)
);

NAND2xp5_ASAP7_75t_L g1108 ( 
.A(n_1013),
.B(n_1027),
.Y(n_1108)
);

OAI21x1_ASAP7_75t_L g1109 ( 
.A1(n_997),
.A2(n_979),
.B(n_1080),
.Y(n_1109)
);

OAI21x1_ASAP7_75t_L g1110 ( 
.A1(n_1080),
.A2(n_1075),
.B(n_975),
.Y(n_1110)
);

BUFx3_ASAP7_75t_L g1111 ( 
.A(n_965),
.Y(n_1111)
);

NOR2xp33_ASAP7_75t_L g1112 ( 
.A(n_1049),
.B(n_963),
.Y(n_1112)
);

OAI21x1_ASAP7_75t_L g1113 ( 
.A1(n_1058),
.A2(n_1079),
.B(n_1077),
.Y(n_1113)
);

A2O1A1Ixp33_ASAP7_75t_L g1114 ( 
.A1(n_960),
.A2(n_1000),
.B(n_1025),
.C(n_957),
.Y(n_1114)
);

BUFx2_ASAP7_75t_R g1115 ( 
.A(n_991),
.Y(n_1115)
);

A2O1A1Ixp33_ASAP7_75t_L g1116 ( 
.A1(n_1014),
.A2(n_1070),
.B(n_948),
.C(n_1030),
.Y(n_1116)
);

INVxp67_ASAP7_75t_SL g1117 ( 
.A(n_945),
.Y(n_1117)
);

AND2x2_ASAP7_75t_L g1118 ( 
.A(n_994),
.B(n_969),
.Y(n_1118)
);

NAND2xp5_ASAP7_75t_SL g1119 ( 
.A(n_1034),
.B(n_1036),
.Y(n_1119)
);

INVx1_ASAP7_75t_L g1120 ( 
.A(n_964),
.Y(n_1120)
);

AND2x4_ASAP7_75t_L g1121 ( 
.A(n_963),
.B(n_987),
.Y(n_1121)
);

OAI21x1_ASAP7_75t_L g1122 ( 
.A1(n_952),
.A2(n_1039),
.B(n_1052),
.Y(n_1122)
);

NOR2xp67_ASAP7_75t_L g1123 ( 
.A(n_1076),
.B(n_1068),
.Y(n_1123)
);

AND2x2_ASAP7_75t_L g1124 ( 
.A(n_944),
.B(n_961),
.Y(n_1124)
);

BUFx2_ASAP7_75t_L g1125 ( 
.A(n_1045),
.Y(n_1125)
);

NAND2xp5_ASAP7_75t_L g1126 ( 
.A(n_961),
.B(n_1016),
.Y(n_1126)
);

OAI22x1_ASAP7_75t_L g1127 ( 
.A1(n_1041),
.A2(n_947),
.B1(n_1023),
.B2(n_985),
.Y(n_1127)
);

AO31x2_ASAP7_75t_L g1128 ( 
.A1(n_1073),
.A2(n_984),
.A3(n_982),
.B(n_967),
.Y(n_1128)
);

NOR2xp33_ASAP7_75t_L g1129 ( 
.A(n_958),
.B(n_1001),
.Y(n_1129)
);

O2A1O1Ixp5_ASAP7_75t_SL g1130 ( 
.A1(n_946),
.A2(n_1033),
.B(n_1035),
.C(n_1031),
.Y(n_1130)
);

OA21x2_ASAP7_75t_L g1131 ( 
.A1(n_950),
.A2(n_1043),
.B(n_1051),
.Y(n_1131)
);

AOI21xp5_ASAP7_75t_L g1132 ( 
.A1(n_967),
.A2(n_1071),
.B(n_1067),
.Y(n_1132)
);

NAND2x1p5_ASAP7_75t_L g1133 ( 
.A(n_987),
.B(n_1026),
.Y(n_1133)
);

OAI21x1_ASAP7_75t_L g1134 ( 
.A1(n_971),
.A2(n_1053),
.B(n_1069),
.Y(n_1134)
);

NOR2xp67_ASAP7_75t_SL g1135 ( 
.A(n_1059),
.B(n_1060),
.Y(n_1135)
);

AO21x2_ASAP7_75t_L g1136 ( 
.A1(n_980),
.A2(n_956),
.B(n_954),
.Y(n_1136)
);

O2A1O1Ixp33_ASAP7_75t_L g1137 ( 
.A1(n_1004),
.A2(n_1028),
.B(n_1010),
.C(n_1018),
.Y(n_1137)
);

INVx3_ASAP7_75t_L g1138 ( 
.A(n_1017),
.Y(n_1138)
);

CKINVDCx5p33_ASAP7_75t_R g1139 ( 
.A(n_993),
.Y(n_1139)
);

NOR2xp67_ASAP7_75t_L g1140 ( 
.A(n_1068),
.B(n_1029),
.Y(n_1140)
);

O2A1O1Ixp5_ASAP7_75t_L g1141 ( 
.A1(n_1021),
.A2(n_1024),
.B(n_1044),
.C(n_1046),
.Y(n_1141)
);

BUFx10_ASAP7_75t_L g1142 ( 
.A(n_1011),
.Y(n_1142)
);

OAI21x1_ASAP7_75t_SL g1143 ( 
.A1(n_992),
.A2(n_1019),
.B(n_1026),
.Y(n_1143)
);

AOI221x1_ASAP7_75t_L g1144 ( 
.A1(n_1021),
.A2(n_1055),
.B1(n_1024),
.B2(n_1007),
.C(n_1041),
.Y(n_1144)
);

NOR2x1_ASAP7_75t_R g1145 ( 
.A(n_1017),
.B(n_989),
.Y(n_1145)
);

AND2x6_ASAP7_75t_L g1146 ( 
.A(n_1009),
.B(n_1029),
.Y(n_1146)
);

AOI21xp5_ASAP7_75t_L g1147 ( 
.A1(n_1054),
.A2(n_1047),
.B(n_1036),
.Y(n_1147)
);

NAND3x1_ASAP7_75t_L g1148 ( 
.A(n_966),
.B(n_1006),
.C(n_968),
.Y(n_1148)
);

AOI22xp5_ASAP7_75t_L g1149 ( 
.A1(n_1056),
.A2(n_1054),
.B1(n_977),
.B2(n_996),
.Y(n_1149)
);

AOI21xp5_ASAP7_75t_L g1150 ( 
.A1(n_1047),
.A2(n_973),
.B(n_1066),
.Y(n_1150)
);

OAI21xp5_ASAP7_75t_L g1151 ( 
.A1(n_999),
.A2(n_1008),
.B(n_1037),
.Y(n_1151)
);

INVx1_ASAP7_75t_L g1152 ( 
.A(n_1003),
.Y(n_1152)
);

AOI21xp5_ASAP7_75t_L g1153 ( 
.A1(n_1066),
.A2(n_1072),
.B(n_1074),
.Y(n_1153)
);

AOI22xp33_ASAP7_75t_L g1154 ( 
.A1(n_1048),
.A2(n_1065),
.B1(n_998),
.B2(n_986),
.Y(n_1154)
);

A2O1A1Ixp33_ASAP7_75t_L g1155 ( 
.A1(n_1012),
.A2(n_1064),
.B(n_970),
.C(n_974),
.Y(n_1155)
);

INVx2_ASAP7_75t_L g1156 ( 
.A(n_970),
.Y(n_1156)
);

INVx1_ASAP7_75t_L g1157 ( 
.A(n_970),
.Y(n_1157)
);

BUFx10_ASAP7_75t_L g1158 ( 
.A(n_974),
.Y(n_1158)
);

INVx4_ASAP7_75t_L g1159 ( 
.A(n_974),
.Y(n_1159)
);

BUFx6f_ASAP7_75t_L g1160 ( 
.A(n_983),
.Y(n_1160)
);

BUFx3_ASAP7_75t_L g1161 ( 
.A(n_983),
.Y(n_1161)
);

AOI22xp5_ASAP7_75t_L g1162 ( 
.A1(n_962),
.A2(n_1061),
.B1(n_1038),
.B2(n_1060),
.Y(n_1162)
);

INVx5_ASAP7_75t_L g1163 ( 
.A(n_983),
.Y(n_1163)
);

INVx1_ASAP7_75t_L g1164 ( 
.A(n_1060),
.Y(n_1164)
);

AOI21xp5_ASAP7_75t_L g1165 ( 
.A1(n_1061),
.A2(n_1038),
.B(n_1064),
.Y(n_1165)
);

OAI21xp5_ASAP7_75t_L g1166 ( 
.A1(n_962),
.A2(n_950),
.B(n_1032),
.Y(n_1166)
);

AOI221x1_ASAP7_75t_L g1167 ( 
.A1(n_1050),
.A2(n_1040),
.B1(n_1002),
.B2(n_1025),
.C(n_821),
.Y(n_1167)
);

INVx2_ASAP7_75t_SL g1168 ( 
.A(n_962),
.Y(n_1168)
);

AOI21xp5_ASAP7_75t_L g1169 ( 
.A1(n_962),
.A2(n_976),
.B(n_949),
.Y(n_1169)
);

OA21x2_ASAP7_75t_L g1170 ( 
.A1(n_962),
.A2(n_1080),
.B(n_988),
.Y(n_1170)
);

AO31x2_ASAP7_75t_L g1171 ( 
.A1(n_988),
.A2(n_774),
.A3(n_895),
.B(n_876),
.Y(n_1171)
);

HB1xp67_ASAP7_75t_L g1172 ( 
.A(n_953),
.Y(n_1172)
);

AOI21xp5_ASAP7_75t_L g1173 ( 
.A1(n_976),
.A2(n_949),
.B(n_765),
.Y(n_1173)
);

OAI21x1_ASAP7_75t_L g1174 ( 
.A1(n_1081),
.A2(n_1063),
.B(n_997),
.Y(n_1174)
);

OAI22xp33_ASAP7_75t_L g1175 ( 
.A1(n_1036),
.A2(n_619),
.B1(n_865),
.B2(n_400),
.Y(n_1175)
);

OAI21x1_ASAP7_75t_L g1176 ( 
.A1(n_1081),
.A2(n_1063),
.B(n_997),
.Y(n_1176)
);

AO31x2_ASAP7_75t_L g1177 ( 
.A1(n_988),
.A2(n_774),
.A3(n_895),
.B(n_876),
.Y(n_1177)
);

INVx1_ASAP7_75t_L g1178 ( 
.A(n_951),
.Y(n_1178)
);

AOI21xp5_ASAP7_75t_L g1179 ( 
.A1(n_976),
.A2(n_949),
.B(n_765),
.Y(n_1179)
);

AO21x1_ASAP7_75t_L g1180 ( 
.A1(n_1002),
.A2(n_1032),
.B(n_946),
.Y(n_1180)
);

AOI21xp5_ASAP7_75t_L g1181 ( 
.A1(n_976),
.A2(n_949),
.B(n_765),
.Y(n_1181)
);

AOI21xp5_ASAP7_75t_L g1182 ( 
.A1(n_976),
.A2(n_949),
.B(n_765),
.Y(n_1182)
);

AOI21xp5_ASAP7_75t_SL g1183 ( 
.A1(n_1076),
.A2(n_765),
.B(n_802),
.Y(n_1183)
);

BUFx10_ASAP7_75t_L g1184 ( 
.A(n_1011),
.Y(n_1184)
);

NAND2xp5_ASAP7_75t_L g1185 ( 
.A(n_972),
.B(n_597),
.Y(n_1185)
);

AOI21xp5_ASAP7_75t_L g1186 ( 
.A1(n_976),
.A2(n_949),
.B(n_765),
.Y(n_1186)
);

OR2x2_ASAP7_75t_L g1187 ( 
.A(n_953),
.B(n_764),
.Y(n_1187)
);

INVx1_ASAP7_75t_SL g1188 ( 
.A(n_953),
.Y(n_1188)
);

AND2x2_ASAP7_75t_L g1189 ( 
.A(n_953),
.B(n_818),
.Y(n_1189)
);

INVx1_ASAP7_75t_SL g1190 ( 
.A(n_953),
.Y(n_1190)
);

INVxp67_ASAP7_75t_L g1191 ( 
.A(n_953),
.Y(n_1191)
);

OAI22x1_ASAP7_75t_L g1192 ( 
.A1(n_1005),
.A2(n_400),
.B1(n_534),
.B2(n_955),
.Y(n_1192)
);

NAND2xp5_ASAP7_75t_L g1193 ( 
.A(n_972),
.B(n_597),
.Y(n_1193)
);

AO31x2_ASAP7_75t_L g1194 ( 
.A1(n_988),
.A2(n_774),
.A3(n_895),
.B(n_876),
.Y(n_1194)
);

INVx1_ASAP7_75t_SL g1195 ( 
.A(n_953),
.Y(n_1195)
);

NAND2x1p5_ASAP7_75t_L g1196 ( 
.A(n_963),
.B(n_1034),
.Y(n_1196)
);

AOI22xp5_ASAP7_75t_L g1197 ( 
.A1(n_955),
.A2(n_865),
.B1(n_821),
.B2(n_568),
.Y(n_1197)
);

INVx3_ASAP7_75t_SL g1198 ( 
.A(n_991),
.Y(n_1198)
);

O2A1O1Ixp33_ASAP7_75t_L g1199 ( 
.A1(n_995),
.A2(n_568),
.B(n_519),
.C(n_506),
.Y(n_1199)
);

OAI21x1_ASAP7_75t_L g1200 ( 
.A1(n_1081),
.A2(n_1063),
.B(n_997),
.Y(n_1200)
);

AOI21xp5_ASAP7_75t_L g1201 ( 
.A1(n_976),
.A2(n_949),
.B(n_765),
.Y(n_1201)
);

AOI21xp5_ASAP7_75t_L g1202 ( 
.A1(n_976),
.A2(n_949),
.B(n_765),
.Y(n_1202)
);

OAI21xp5_ASAP7_75t_SL g1203 ( 
.A1(n_1020),
.A2(n_568),
.B(n_995),
.Y(n_1203)
);

OR2x2_ASAP7_75t_L g1204 ( 
.A(n_953),
.B(n_764),
.Y(n_1204)
);

AOI21xp5_ASAP7_75t_L g1205 ( 
.A1(n_976),
.A2(n_949),
.B(n_765),
.Y(n_1205)
);

AO31x2_ASAP7_75t_L g1206 ( 
.A1(n_988),
.A2(n_774),
.A3(n_895),
.B(n_876),
.Y(n_1206)
);

O2A1O1Ixp33_ASAP7_75t_L g1207 ( 
.A1(n_995),
.A2(n_568),
.B(n_519),
.C(n_506),
.Y(n_1207)
);

OAI21xp5_ASAP7_75t_L g1208 ( 
.A1(n_950),
.A2(n_1032),
.B(n_949),
.Y(n_1208)
);

NOR2xp67_ASAP7_75t_SL g1209 ( 
.A(n_991),
.B(n_534),
.Y(n_1209)
);

OAI21x1_ASAP7_75t_L g1210 ( 
.A1(n_1081),
.A2(n_1063),
.B(n_997),
.Y(n_1210)
);

INVx5_ASAP7_75t_L g1211 ( 
.A(n_1034),
.Y(n_1211)
);

OA21x2_ASAP7_75t_L g1212 ( 
.A1(n_1080),
.A2(n_988),
.B(n_1063),
.Y(n_1212)
);

AO31x2_ASAP7_75t_L g1213 ( 
.A1(n_988),
.A2(n_774),
.A3(n_895),
.B(n_876),
.Y(n_1213)
);

CKINVDCx5p33_ASAP7_75t_R g1214 ( 
.A(n_991),
.Y(n_1214)
);

INVxp67_ASAP7_75t_L g1215 ( 
.A(n_953),
.Y(n_1215)
);

INVx1_ASAP7_75t_L g1216 ( 
.A(n_951),
.Y(n_1216)
);

INVx2_ASAP7_75t_SL g1217 ( 
.A(n_990),
.Y(n_1217)
);

OAI21x1_ASAP7_75t_L g1218 ( 
.A1(n_1081),
.A2(n_1063),
.B(n_997),
.Y(n_1218)
);

AOI22xp33_ASAP7_75t_L g1219 ( 
.A1(n_1005),
.A2(n_818),
.B1(n_360),
.B2(n_337),
.Y(n_1219)
);

BUFx12f_ASAP7_75t_L g1220 ( 
.A(n_1139),
.Y(n_1220)
);

AND2x2_ASAP7_75t_L g1221 ( 
.A(n_1124),
.B(n_1189),
.Y(n_1221)
);

AOI22xp33_ASAP7_75t_L g1222 ( 
.A1(n_1197),
.A2(n_1149),
.B1(n_1219),
.B2(n_1175),
.Y(n_1222)
);

INVx1_ASAP7_75t_L g1223 ( 
.A(n_1088),
.Y(n_1223)
);

INVx1_ASAP7_75t_L g1224 ( 
.A(n_1096),
.Y(n_1224)
);

OAI22xp5_ASAP7_75t_SL g1225 ( 
.A1(n_1197),
.A2(n_1192),
.B1(n_1129),
.B2(n_1149),
.Y(n_1225)
);

BUFx12f_ASAP7_75t_L g1226 ( 
.A(n_1214),
.Y(n_1226)
);

AOI22xp33_ASAP7_75t_L g1227 ( 
.A1(n_1147),
.A2(n_1204),
.B1(n_1187),
.B2(n_1193),
.Y(n_1227)
);

BUFx12f_ASAP7_75t_L g1228 ( 
.A(n_1142),
.Y(n_1228)
);

INVx1_ASAP7_75t_L g1229 ( 
.A(n_1120),
.Y(n_1229)
);

NAND2xp5_ASAP7_75t_L g1230 ( 
.A(n_1185),
.B(n_1108),
.Y(n_1230)
);

INVx8_ASAP7_75t_L g1231 ( 
.A(n_1146),
.Y(n_1231)
);

BUFx12f_ASAP7_75t_L g1232 ( 
.A(n_1142),
.Y(n_1232)
);

AND2x2_ASAP7_75t_L g1233 ( 
.A(n_1118),
.B(n_1188),
.Y(n_1233)
);

BUFx4f_ASAP7_75t_SL g1234 ( 
.A(n_1198),
.Y(n_1234)
);

BUFx2_ASAP7_75t_L g1235 ( 
.A(n_1172),
.Y(n_1235)
);

BUFx8_ASAP7_75t_L g1236 ( 
.A(n_1125),
.Y(n_1236)
);

INVx1_ASAP7_75t_SL g1237 ( 
.A(n_1188),
.Y(n_1237)
);

CKINVDCx5p33_ASAP7_75t_R g1238 ( 
.A(n_1115),
.Y(n_1238)
);

AND2x2_ASAP7_75t_L g1239 ( 
.A(n_1190),
.B(n_1195),
.Y(n_1239)
);

OAI22xp5_ASAP7_75t_L g1240 ( 
.A1(n_1199),
.A2(n_1207),
.B1(n_1203),
.B2(n_1114),
.Y(n_1240)
);

AND2x2_ASAP7_75t_L g1241 ( 
.A(n_1190),
.B(n_1195),
.Y(n_1241)
);

AOI22xp33_ASAP7_75t_L g1242 ( 
.A1(n_1127),
.A2(n_1097),
.B1(n_1152),
.B2(n_1178),
.Y(n_1242)
);

CKINVDCx6p67_ASAP7_75t_R g1243 ( 
.A(n_1111),
.Y(n_1243)
);

OAI22xp5_ASAP7_75t_L g1244 ( 
.A1(n_1203),
.A2(n_1116),
.B1(n_1137),
.B2(n_1183),
.Y(n_1244)
);

INVx2_ASAP7_75t_SL g1245 ( 
.A(n_1085),
.Y(n_1245)
);

BUFx5_ASAP7_75t_L g1246 ( 
.A(n_1146),
.Y(n_1246)
);

NAND2x1p5_ASAP7_75t_L g1247 ( 
.A(n_1211),
.B(n_1082),
.Y(n_1247)
);

INVx6_ASAP7_75t_L g1248 ( 
.A(n_1163),
.Y(n_1248)
);

CKINVDCx6p67_ASAP7_75t_R g1249 ( 
.A(n_1184),
.Y(n_1249)
);

INVx1_ASAP7_75t_L g1250 ( 
.A(n_1216),
.Y(n_1250)
);

BUFx2_ASAP7_75t_SL g1251 ( 
.A(n_1217),
.Y(n_1251)
);

BUFx8_ASAP7_75t_L g1252 ( 
.A(n_1160),
.Y(n_1252)
);

INVx4_ASAP7_75t_L g1253 ( 
.A(n_1211),
.Y(n_1253)
);

CKINVDCx11_ASAP7_75t_R g1254 ( 
.A(n_1184),
.Y(n_1254)
);

CKINVDCx11_ASAP7_75t_R g1255 ( 
.A(n_1158),
.Y(n_1255)
);

OAI22xp5_ASAP7_75t_L g1256 ( 
.A1(n_1154),
.A2(n_1132),
.B1(n_1099),
.B2(n_1148),
.Y(n_1256)
);

NAND2x1p5_ASAP7_75t_L g1257 ( 
.A(n_1211),
.B(n_1082),
.Y(n_1257)
);

INVx4_ASAP7_75t_L g1258 ( 
.A(n_1160),
.Y(n_1258)
);

AOI22xp33_ASAP7_75t_L g1259 ( 
.A1(n_1098),
.A2(n_1100),
.B1(n_1215),
.B2(n_1191),
.Y(n_1259)
);

CKINVDCx11_ASAP7_75t_R g1260 ( 
.A(n_1158),
.Y(n_1260)
);

CKINVDCx12_ASAP7_75t_R g1261 ( 
.A(n_1145),
.Y(n_1261)
);

BUFx4f_ASAP7_75t_L g1262 ( 
.A(n_1146),
.Y(n_1262)
);

CKINVDCx11_ASAP7_75t_R g1263 ( 
.A(n_1161),
.Y(n_1263)
);

CKINVDCx11_ASAP7_75t_R g1264 ( 
.A(n_1156),
.Y(n_1264)
);

AOI22xp33_ASAP7_75t_L g1265 ( 
.A1(n_1098),
.A2(n_1099),
.B1(n_1126),
.B2(n_1180),
.Y(n_1265)
);

AOI22xp33_ASAP7_75t_L g1266 ( 
.A1(n_1208),
.A2(n_1091),
.B1(n_1117),
.B2(n_1119),
.Y(n_1266)
);

AOI22xp33_ASAP7_75t_SL g1267 ( 
.A1(n_1131),
.A2(n_1208),
.B1(n_1166),
.B2(n_1141),
.Y(n_1267)
);

AOI22xp33_ASAP7_75t_L g1268 ( 
.A1(n_1105),
.A2(n_1131),
.B1(n_1136),
.B2(n_1094),
.Y(n_1268)
);

INVx1_ASAP7_75t_L g1269 ( 
.A(n_1089),
.Y(n_1269)
);

CKINVDCx20_ASAP7_75t_R g1270 ( 
.A(n_1090),
.Y(n_1270)
);

BUFx6f_ASAP7_75t_L g1271 ( 
.A(n_1121),
.Y(n_1271)
);

AND2x2_ASAP7_75t_L g1272 ( 
.A(n_1112),
.B(n_1138),
.Y(n_1272)
);

AOI22xp33_ASAP7_75t_L g1273 ( 
.A1(n_1136),
.A2(n_1094),
.B1(n_1166),
.B2(n_1146),
.Y(n_1273)
);

AOI22xp33_ASAP7_75t_SL g1274 ( 
.A1(n_1167),
.A2(n_1170),
.B1(n_1144),
.B2(n_1093),
.Y(n_1274)
);

INVx2_ASAP7_75t_L g1275 ( 
.A(n_1157),
.Y(n_1275)
);

INVx1_ASAP7_75t_L g1276 ( 
.A(n_1164),
.Y(n_1276)
);

INVx1_ASAP7_75t_L g1277 ( 
.A(n_1113),
.Y(n_1277)
);

INVx1_ASAP7_75t_SL g1278 ( 
.A(n_1121),
.Y(n_1278)
);

CKINVDCx11_ASAP7_75t_R g1279 ( 
.A(n_1209),
.Y(n_1279)
);

CKINVDCx5p33_ASAP7_75t_R g1280 ( 
.A(n_1159),
.Y(n_1280)
);

INVxp33_ASAP7_75t_SL g1281 ( 
.A(n_1135),
.Y(n_1281)
);

AOI22xp33_ASAP7_75t_SL g1282 ( 
.A1(n_1170),
.A2(n_1093),
.B1(n_1138),
.B2(n_1212),
.Y(n_1282)
);

BUFx3_ASAP7_75t_L g1283 ( 
.A(n_1133),
.Y(n_1283)
);

AOI22xp33_ASAP7_75t_L g1284 ( 
.A1(n_1151),
.A2(n_1179),
.B1(n_1201),
.B2(n_1181),
.Y(n_1284)
);

INVxp67_ASAP7_75t_SL g1285 ( 
.A(n_1212),
.Y(n_1285)
);

BUFx4_ASAP7_75t_SL g1286 ( 
.A(n_1145),
.Y(n_1286)
);

INVx6_ASAP7_75t_L g1287 ( 
.A(n_1159),
.Y(n_1287)
);

INVx3_ASAP7_75t_SL g1288 ( 
.A(n_1168),
.Y(n_1288)
);

CKINVDCx20_ASAP7_75t_R g1289 ( 
.A(n_1162),
.Y(n_1289)
);

INVx1_ASAP7_75t_L g1290 ( 
.A(n_1143),
.Y(n_1290)
);

AOI22xp33_ASAP7_75t_SL g1291 ( 
.A1(n_1151),
.A2(n_1150),
.B1(n_1205),
.B2(n_1202),
.Y(n_1291)
);

AOI22xp5_ASAP7_75t_L g1292 ( 
.A1(n_1140),
.A2(n_1123),
.B1(n_1162),
.B2(n_1153),
.Y(n_1292)
);

AOI21xp33_ASAP7_75t_L g1293 ( 
.A1(n_1103),
.A2(n_1095),
.B(n_1134),
.Y(n_1293)
);

CKINVDCx16_ASAP7_75t_R g1294 ( 
.A(n_1103),
.Y(n_1294)
);

INVx1_ASAP7_75t_L g1295 ( 
.A(n_1140),
.Y(n_1295)
);

INVx1_ASAP7_75t_L g1296 ( 
.A(n_1084),
.Y(n_1296)
);

INVx6_ASAP7_75t_L g1297 ( 
.A(n_1196),
.Y(n_1297)
);

INVx4_ASAP7_75t_L g1298 ( 
.A(n_1155),
.Y(n_1298)
);

BUFx2_ASAP7_75t_L g1299 ( 
.A(n_1128),
.Y(n_1299)
);

NAND2xp5_ASAP7_75t_L g1300 ( 
.A(n_1173),
.B(n_1186),
.Y(n_1300)
);

CKINVDCx11_ASAP7_75t_R g1301 ( 
.A(n_1092),
.Y(n_1301)
);

OAI22x1_ASAP7_75t_L g1302 ( 
.A1(n_1130),
.A2(n_1092),
.B1(n_1128),
.B2(n_1165),
.Y(n_1302)
);

BUFx8_ASAP7_75t_L g1303 ( 
.A(n_1123),
.Y(n_1303)
);

INVx6_ASAP7_75t_L g1304 ( 
.A(n_1110),
.Y(n_1304)
);

AOI22xp33_ASAP7_75t_L g1305 ( 
.A1(n_1182),
.A2(n_1087),
.B1(n_1083),
.B2(n_1169),
.Y(n_1305)
);

CKINVDCx20_ASAP7_75t_R g1306 ( 
.A(n_1106),
.Y(n_1306)
);

BUFx2_ASAP7_75t_SL g1307 ( 
.A(n_1104),
.Y(n_1307)
);

AOI22xp33_ASAP7_75t_SL g1308 ( 
.A1(n_1122),
.A2(n_1109),
.B1(n_1102),
.B2(n_1218),
.Y(n_1308)
);

INVx1_ASAP7_75t_L g1309 ( 
.A(n_1171),
.Y(n_1309)
);

INVx3_ASAP7_75t_SL g1310 ( 
.A(n_1177),
.Y(n_1310)
);

CKINVDCx5p33_ASAP7_75t_R g1311 ( 
.A(n_1177),
.Y(n_1311)
);

AOI22xp33_ASAP7_75t_SL g1312 ( 
.A1(n_1174),
.A2(n_1210),
.B1(n_1200),
.B2(n_1176),
.Y(n_1312)
);

OAI22xp33_ASAP7_75t_L g1313 ( 
.A1(n_1194),
.A2(n_1206),
.B1(n_1213),
.B2(n_1107),
.Y(n_1313)
);

AOI22xp33_ASAP7_75t_L g1314 ( 
.A1(n_1101),
.A2(n_1086),
.B1(n_1194),
.B2(n_1206),
.Y(n_1314)
);

INVx3_ASAP7_75t_L g1315 ( 
.A(n_1194),
.Y(n_1315)
);

INVx1_ASAP7_75t_L g1316 ( 
.A(n_1213),
.Y(n_1316)
);

OAI22xp33_ASAP7_75t_L g1317 ( 
.A1(n_1206),
.A2(n_1197),
.B1(n_1149),
.B2(n_1147),
.Y(n_1317)
);

INVx1_ASAP7_75t_L g1318 ( 
.A(n_1107),
.Y(n_1318)
);

CKINVDCx20_ASAP7_75t_R g1319 ( 
.A(n_1107),
.Y(n_1319)
);

AOI22xp33_ASAP7_75t_L g1320 ( 
.A1(n_1197),
.A2(n_821),
.B1(n_662),
.B2(n_1149),
.Y(n_1320)
);

NAND2x1p5_ASAP7_75t_L g1321 ( 
.A(n_1211),
.B(n_1034),
.Y(n_1321)
);

AOI22x1_ASAP7_75t_SL g1322 ( 
.A1(n_1139),
.A2(n_1214),
.B1(n_534),
.B2(n_215),
.Y(n_1322)
);

AOI22xp33_ASAP7_75t_L g1323 ( 
.A1(n_1197),
.A2(n_821),
.B1(n_662),
.B2(n_1149),
.Y(n_1323)
);

OAI22xp5_ASAP7_75t_L g1324 ( 
.A1(n_1197),
.A2(n_1147),
.B1(n_1207),
.B2(n_1199),
.Y(n_1324)
);

OAI22xp5_ASAP7_75t_L g1325 ( 
.A1(n_1197),
.A2(n_1147),
.B1(n_1207),
.B2(n_1199),
.Y(n_1325)
);

OAI22xp5_ASAP7_75t_SL g1326 ( 
.A1(n_1197),
.A2(n_1192),
.B1(n_1219),
.B2(n_534),
.Y(n_1326)
);

AOI22xp33_ASAP7_75t_SL g1327 ( 
.A1(n_1147),
.A2(n_337),
.B1(n_344),
.B2(n_342),
.Y(n_1327)
);

AOI22xp33_ASAP7_75t_L g1328 ( 
.A1(n_1197),
.A2(n_821),
.B1(n_662),
.B2(n_1149),
.Y(n_1328)
);

HB1xp67_ASAP7_75t_SL g1329 ( 
.A(n_1111),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_1088),
.Y(n_1330)
);

NAND2xp5_ASAP7_75t_L g1331 ( 
.A(n_1185),
.B(n_1193),
.Y(n_1331)
);

AOI22xp33_ASAP7_75t_L g1332 ( 
.A1(n_1197),
.A2(n_821),
.B1(n_662),
.B2(n_1149),
.Y(n_1332)
);

INVx1_ASAP7_75t_L g1333 ( 
.A(n_1088),
.Y(n_1333)
);

AOI22xp33_ASAP7_75t_L g1334 ( 
.A1(n_1197),
.A2(n_821),
.B1(n_662),
.B2(n_1149),
.Y(n_1334)
);

OAI22xp5_ASAP7_75t_L g1335 ( 
.A1(n_1197),
.A2(n_1147),
.B1(n_1207),
.B2(n_1199),
.Y(n_1335)
);

INVx1_ASAP7_75t_L g1336 ( 
.A(n_1088),
.Y(n_1336)
);

AOI22xp33_ASAP7_75t_L g1337 ( 
.A1(n_1197),
.A2(n_821),
.B1(n_662),
.B2(n_1149),
.Y(n_1337)
);

INVx1_ASAP7_75t_L g1338 ( 
.A(n_1296),
.Y(n_1338)
);

NAND2xp5_ASAP7_75t_L g1339 ( 
.A(n_1230),
.B(n_1294),
.Y(n_1339)
);

HB1xp67_ASAP7_75t_L g1340 ( 
.A(n_1318),
.Y(n_1340)
);

INVx1_ASAP7_75t_L g1341 ( 
.A(n_1309),
.Y(n_1341)
);

BUFx2_ASAP7_75t_L g1342 ( 
.A(n_1304),
.Y(n_1342)
);

AND2x2_ASAP7_75t_L g1343 ( 
.A(n_1223),
.B(n_1224),
.Y(n_1343)
);

HB1xp67_ASAP7_75t_L g1344 ( 
.A(n_1300),
.Y(n_1344)
);

INVx1_ASAP7_75t_L g1345 ( 
.A(n_1316),
.Y(n_1345)
);

INVx2_ASAP7_75t_SL g1346 ( 
.A(n_1304),
.Y(n_1346)
);

INVx3_ASAP7_75t_L g1347 ( 
.A(n_1304),
.Y(n_1347)
);

AND2x2_ASAP7_75t_L g1348 ( 
.A(n_1229),
.B(n_1250),
.Y(n_1348)
);

AND2x2_ASAP7_75t_L g1349 ( 
.A(n_1330),
.B(n_1333),
.Y(n_1349)
);

OR2x2_ASAP7_75t_L g1350 ( 
.A(n_1235),
.B(n_1311),
.Y(n_1350)
);

INVx1_ASAP7_75t_L g1351 ( 
.A(n_1277),
.Y(n_1351)
);

INVx1_ASAP7_75t_L g1352 ( 
.A(n_1336),
.Y(n_1352)
);

INVx6_ASAP7_75t_L g1353 ( 
.A(n_1231),
.Y(n_1353)
);

AND2x2_ASAP7_75t_L g1354 ( 
.A(n_1233),
.B(n_1221),
.Y(n_1354)
);

INVx2_ASAP7_75t_SL g1355 ( 
.A(n_1290),
.Y(n_1355)
);

INVxp67_ASAP7_75t_L g1356 ( 
.A(n_1302),
.Y(n_1356)
);

OAI21xp5_ASAP7_75t_L g1357 ( 
.A1(n_1337),
.A2(n_1323),
.B(n_1320),
.Y(n_1357)
);

INVx1_ASAP7_75t_L g1358 ( 
.A(n_1315),
.Y(n_1358)
);

INVx1_ASAP7_75t_L g1359 ( 
.A(n_1299),
.Y(n_1359)
);

HB1xp67_ASAP7_75t_L g1360 ( 
.A(n_1285),
.Y(n_1360)
);

AND2x2_ASAP7_75t_L g1361 ( 
.A(n_1285),
.B(n_1267),
.Y(n_1361)
);

OAI21x1_ASAP7_75t_L g1362 ( 
.A1(n_1305),
.A2(n_1284),
.B(n_1314),
.Y(n_1362)
);

INVx1_ASAP7_75t_L g1363 ( 
.A(n_1269),
.Y(n_1363)
);

BUFx2_ASAP7_75t_L g1364 ( 
.A(n_1306),
.Y(n_1364)
);

AOI21xp5_ASAP7_75t_L g1365 ( 
.A1(n_1305),
.A2(n_1284),
.B(n_1240),
.Y(n_1365)
);

INVx2_ASAP7_75t_L g1366 ( 
.A(n_1310),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_1313),
.Y(n_1367)
);

INVx1_ASAP7_75t_L g1368 ( 
.A(n_1313),
.Y(n_1368)
);

INVx4_ASAP7_75t_L g1369 ( 
.A(n_1262),
.Y(n_1369)
);

NAND2xp5_ASAP7_75t_L g1370 ( 
.A(n_1317),
.B(n_1265),
.Y(n_1370)
);

INVx1_ASAP7_75t_L g1371 ( 
.A(n_1319),
.Y(n_1371)
);

AOI22xp33_ASAP7_75t_SL g1372 ( 
.A1(n_1225),
.A2(n_1256),
.B1(n_1335),
.B2(n_1325),
.Y(n_1372)
);

HB1xp67_ASAP7_75t_L g1373 ( 
.A(n_1314),
.Y(n_1373)
);

INVx2_ASAP7_75t_L g1374 ( 
.A(n_1310),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_1276),
.Y(n_1375)
);

NAND2xp5_ASAP7_75t_L g1376 ( 
.A(n_1317),
.B(n_1265),
.Y(n_1376)
);

INVx1_ASAP7_75t_L g1377 ( 
.A(n_1282),
.Y(n_1377)
);

INVx1_ASAP7_75t_L g1378 ( 
.A(n_1282),
.Y(n_1378)
);

INVx4_ASAP7_75t_L g1379 ( 
.A(n_1231),
.Y(n_1379)
);

BUFx3_ASAP7_75t_L g1380 ( 
.A(n_1246),
.Y(n_1380)
);

OAI21x1_ASAP7_75t_L g1381 ( 
.A1(n_1268),
.A2(n_1273),
.B(n_1244),
.Y(n_1381)
);

AND2x4_ASAP7_75t_L g1382 ( 
.A(n_1292),
.B(n_1295),
.Y(n_1382)
);

AOI22xp33_ASAP7_75t_L g1383 ( 
.A1(n_1222),
.A2(n_1327),
.B1(n_1334),
.B2(n_1332),
.Y(n_1383)
);

HB1xp67_ASAP7_75t_L g1384 ( 
.A(n_1239),
.Y(n_1384)
);

BUFx2_ASAP7_75t_L g1385 ( 
.A(n_1288),
.Y(n_1385)
);

AND2x4_ASAP7_75t_L g1386 ( 
.A(n_1273),
.B(n_1298),
.Y(n_1386)
);

OAI21x1_ASAP7_75t_L g1387 ( 
.A1(n_1268),
.A2(n_1324),
.B(n_1266),
.Y(n_1387)
);

INVx1_ASAP7_75t_L g1388 ( 
.A(n_1267),
.Y(n_1388)
);

OA21x2_ASAP7_75t_L g1389 ( 
.A1(n_1293),
.A2(n_1266),
.B(n_1242),
.Y(n_1389)
);

AND2x2_ASAP7_75t_L g1390 ( 
.A(n_1241),
.B(n_1274),
.Y(n_1390)
);

BUFx2_ASAP7_75t_L g1391 ( 
.A(n_1288),
.Y(n_1391)
);

HB1xp67_ASAP7_75t_L g1392 ( 
.A(n_1307),
.Y(n_1392)
);

OAI21x1_ASAP7_75t_L g1393 ( 
.A1(n_1242),
.A2(n_1321),
.B(n_1257),
.Y(n_1393)
);

NAND2xp5_ASAP7_75t_L g1394 ( 
.A(n_1331),
.B(n_1227),
.Y(n_1394)
);

OR2x2_ASAP7_75t_L g1395 ( 
.A(n_1227),
.B(n_1237),
.Y(n_1395)
);

INVx1_ASAP7_75t_L g1396 ( 
.A(n_1275),
.Y(n_1396)
);

INVx1_ASAP7_75t_L g1397 ( 
.A(n_1291),
.Y(n_1397)
);

AND2x2_ASAP7_75t_L g1398 ( 
.A(n_1274),
.B(n_1272),
.Y(n_1398)
);

INVx1_ASAP7_75t_L g1399 ( 
.A(n_1291),
.Y(n_1399)
);

INVx1_ASAP7_75t_L g1400 ( 
.A(n_1308),
.Y(n_1400)
);

INVx1_ASAP7_75t_L g1401 ( 
.A(n_1308),
.Y(n_1401)
);

OA21x2_ASAP7_75t_L g1402 ( 
.A1(n_1320),
.A2(n_1337),
.B(n_1323),
.Y(n_1402)
);

OR2x2_ASAP7_75t_L g1403 ( 
.A(n_1328),
.B(n_1332),
.Y(n_1403)
);

INVx1_ASAP7_75t_L g1404 ( 
.A(n_1298),
.Y(n_1404)
);

INVx1_ASAP7_75t_L g1405 ( 
.A(n_1312),
.Y(n_1405)
);

NAND2xp5_ASAP7_75t_L g1406 ( 
.A(n_1328),
.B(n_1334),
.Y(n_1406)
);

INVx1_ASAP7_75t_L g1407 ( 
.A(n_1312),
.Y(n_1407)
);

INVx3_ASAP7_75t_L g1408 ( 
.A(n_1253),
.Y(n_1408)
);

BUFx2_ASAP7_75t_L g1409 ( 
.A(n_1258),
.Y(n_1409)
);

AND2x2_ASAP7_75t_L g1410 ( 
.A(n_1259),
.B(n_1222),
.Y(n_1410)
);

NOR2xp33_ASAP7_75t_L g1411 ( 
.A(n_1322),
.B(n_1326),
.Y(n_1411)
);

OR2x6_ASAP7_75t_L g1412 ( 
.A(n_1321),
.B(n_1247),
.Y(n_1412)
);

HB1xp67_ASAP7_75t_L g1413 ( 
.A(n_1278),
.Y(n_1413)
);

INVx2_ASAP7_75t_L g1414 ( 
.A(n_1289),
.Y(n_1414)
);

OA21x2_ASAP7_75t_L g1415 ( 
.A1(n_1259),
.A2(n_1280),
.B(n_1245),
.Y(n_1415)
);

AND2x2_ASAP7_75t_L g1416 ( 
.A(n_1271),
.B(n_1251),
.Y(n_1416)
);

AO21x2_ASAP7_75t_L g1417 ( 
.A1(n_1370),
.A2(n_1261),
.B(n_1327),
.Y(n_1417)
);

OA21x2_ASAP7_75t_L g1418 ( 
.A1(n_1362),
.A2(n_1301),
.B(n_1297),
.Y(n_1418)
);

NAND2x1p5_ASAP7_75t_L g1419 ( 
.A(n_1404),
.B(n_1369),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_1352),
.Y(n_1420)
);

OR2x2_ASAP7_75t_L g1421 ( 
.A(n_1384),
.B(n_1243),
.Y(n_1421)
);

AO32x2_ASAP7_75t_L g1422 ( 
.A1(n_1355),
.A2(n_1329),
.A3(n_1264),
.B1(n_1249),
.B2(n_1263),
.Y(n_1422)
);

AND2x2_ASAP7_75t_L g1423 ( 
.A(n_1364),
.B(n_1271),
.Y(n_1423)
);

AO21x1_ASAP7_75t_L g1424 ( 
.A1(n_1406),
.A2(n_1329),
.B(n_1286),
.Y(n_1424)
);

OR2x6_ASAP7_75t_L g1425 ( 
.A(n_1393),
.B(n_1248),
.Y(n_1425)
);

OAI21xp5_ASAP7_75t_L g1426 ( 
.A1(n_1357),
.A2(n_1281),
.B(n_1270),
.Y(n_1426)
);

NOR2x1_ASAP7_75t_L g1427 ( 
.A(n_1404),
.B(n_1283),
.Y(n_1427)
);

AND2x2_ASAP7_75t_L g1428 ( 
.A(n_1364),
.B(n_1238),
.Y(n_1428)
);

INVxp67_ASAP7_75t_L g1429 ( 
.A(n_1344),
.Y(n_1429)
);

CKINVDCx20_ASAP7_75t_R g1430 ( 
.A(n_1385),
.Y(n_1430)
);

AND2x2_ASAP7_75t_L g1431 ( 
.A(n_1354),
.B(n_1254),
.Y(n_1431)
);

AND2x2_ASAP7_75t_L g1432 ( 
.A(n_1354),
.B(n_1279),
.Y(n_1432)
);

AND2x4_ASAP7_75t_L g1433 ( 
.A(n_1350),
.B(n_1234),
.Y(n_1433)
);

INVx1_ASAP7_75t_L g1434 ( 
.A(n_1375),
.Y(n_1434)
);

A2O1A1Ixp33_ASAP7_75t_L g1435 ( 
.A1(n_1357),
.A2(n_1383),
.B(n_1403),
.C(n_1372),
.Y(n_1435)
);

A2O1A1Ixp33_ASAP7_75t_L g1436 ( 
.A1(n_1403),
.A2(n_1303),
.B(n_1252),
.C(n_1248),
.Y(n_1436)
);

AND2x2_ASAP7_75t_L g1437 ( 
.A(n_1390),
.B(n_1260),
.Y(n_1437)
);

NOR2x1_ASAP7_75t_SL g1438 ( 
.A(n_1412),
.B(n_1228),
.Y(n_1438)
);

NAND2xp5_ASAP7_75t_L g1439 ( 
.A(n_1344),
.B(n_1252),
.Y(n_1439)
);

OAI21xp5_ASAP7_75t_L g1440 ( 
.A1(n_1406),
.A2(n_1232),
.B(n_1255),
.Y(n_1440)
);

INVx4_ASAP7_75t_L g1441 ( 
.A(n_1385),
.Y(n_1441)
);

AND2x2_ASAP7_75t_L g1442 ( 
.A(n_1390),
.B(n_1287),
.Y(n_1442)
);

AOI221xp5_ASAP7_75t_L g1443 ( 
.A1(n_1372),
.A2(n_1236),
.B1(n_1234),
.B2(n_1220),
.C(n_1226),
.Y(n_1443)
);

BUFx3_ASAP7_75t_L g1444 ( 
.A(n_1391),
.Y(n_1444)
);

NAND4xp25_ASAP7_75t_L g1445 ( 
.A(n_1365),
.B(n_1236),
.C(n_1287),
.D(n_1397),
.Y(n_1445)
);

OAI211xp5_ASAP7_75t_L g1446 ( 
.A1(n_1402),
.A2(n_1365),
.B(n_1397),
.C(n_1399),
.Y(n_1446)
);

AND2x2_ASAP7_75t_L g1447 ( 
.A(n_1398),
.B(n_1343),
.Y(n_1447)
);

AO32x1_ASAP7_75t_L g1448 ( 
.A1(n_1355),
.A2(n_1410),
.A3(n_1378),
.B1(n_1377),
.B2(n_1388),
.Y(n_1448)
);

AND2x2_ASAP7_75t_L g1449 ( 
.A(n_1398),
.B(n_1343),
.Y(n_1449)
);

OA21x2_ASAP7_75t_L g1450 ( 
.A1(n_1356),
.A2(n_1381),
.B(n_1400),
.Y(n_1450)
);

AO32x1_ASAP7_75t_L g1451 ( 
.A1(n_1355),
.A2(n_1410),
.A3(n_1377),
.B1(n_1378),
.B2(n_1388),
.Y(n_1451)
);

OR2x2_ASAP7_75t_L g1452 ( 
.A(n_1339),
.B(n_1395),
.Y(n_1452)
);

NAND3xp33_ASAP7_75t_L g1453 ( 
.A(n_1402),
.B(n_1399),
.C(n_1356),
.Y(n_1453)
);

AOI21xp5_ASAP7_75t_L g1454 ( 
.A1(n_1402),
.A2(n_1360),
.B(n_1387),
.Y(n_1454)
);

AO32x1_ASAP7_75t_L g1455 ( 
.A1(n_1405),
.A2(n_1407),
.A3(n_1346),
.B1(n_1401),
.B2(n_1400),
.Y(n_1455)
);

AO21x2_ASAP7_75t_L g1456 ( 
.A1(n_1376),
.A2(n_1401),
.B(n_1407),
.Y(n_1456)
);

NAND2xp5_ASAP7_75t_L g1457 ( 
.A(n_1394),
.B(n_1348),
.Y(n_1457)
);

CKINVDCx5p33_ASAP7_75t_R g1458 ( 
.A(n_1391),
.Y(n_1458)
);

OAI21xp5_ASAP7_75t_L g1459 ( 
.A1(n_1402),
.A2(n_1387),
.B(n_1376),
.Y(n_1459)
);

OR2x6_ASAP7_75t_L g1460 ( 
.A(n_1393),
.B(n_1386),
.Y(n_1460)
);

AND2x4_ASAP7_75t_L g1461 ( 
.A(n_1382),
.B(n_1380),
.Y(n_1461)
);

AND2x2_ASAP7_75t_L g1462 ( 
.A(n_1348),
.B(n_1349),
.Y(n_1462)
);

NOR2xp33_ASAP7_75t_L g1463 ( 
.A(n_1402),
.B(n_1339),
.Y(n_1463)
);

OAI221xp5_ASAP7_75t_SL g1464 ( 
.A1(n_1361),
.A2(n_1394),
.B1(n_1411),
.B2(n_1395),
.C(n_1405),
.Y(n_1464)
);

OR2x2_ASAP7_75t_L g1465 ( 
.A(n_1349),
.B(n_1371),
.Y(n_1465)
);

AND2x2_ASAP7_75t_L g1466 ( 
.A(n_1371),
.B(n_1416),
.Y(n_1466)
);

OAI22xp5_ASAP7_75t_L g1467 ( 
.A1(n_1386),
.A2(n_1389),
.B1(n_1368),
.B2(n_1367),
.Y(n_1467)
);

OR2x2_ASAP7_75t_L g1468 ( 
.A(n_1363),
.B(n_1413),
.Y(n_1468)
);

OR2x2_ASAP7_75t_L g1469 ( 
.A(n_1363),
.B(n_1367),
.Y(n_1469)
);

AND2x4_ASAP7_75t_L g1470 ( 
.A(n_1382),
.B(n_1380),
.Y(n_1470)
);

OAI22xp5_ASAP7_75t_L g1471 ( 
.A1(n_1386),
.A2(n_1389),
.B1(n_1368),
.B2(n_1379),
.Y(n_1471)
);

OAI22xp5_ASAP7_75t_L g1472 ( 
.A1(n_1389),
.A2(n_1379),
.B1(n_1353),
.B2(n_1369),
.Y(n_1472)
);

AOI221xp5_ASAP7_75t_L g1473 ( 
.A1(n_1373),
.A2(n_1382),
.B1(n_1360),
.B2(n_1351),
.C(n_1359),
.Y(n_1473)
);

NAND2xp5_ASAP7_75t_L g1474 ( 
.A(n_1389),
.B(n_1392),
.Y(n_1474)
);

OR2x2_ASAP7_75t_L g1475 ( 
.A(n_1457),
.B(n_1452),
.Y(n_1475)
);

AOI22xp33_ASAP7_75t_L g1476 ( 
.A1(n_1417),
.A2(n_1373),
.B1(n_1389),
.B2(n_1415),
.Y(n_1476)
);

INVx1_ASAP7_75t_L g1477 ( 
.A(n_1420),
.Y(n_1477)
);

NOR2xp33_ASAP7_75t_L g1478 ( 
.A(n_1458),
.B(n_1433),
.Y(n_1478)
);

AND2x4_ASAP7_75t_L g1479 ( 
.A(n_1461),
.B(n_1380),
.Y(n_1479)
);

INVxp67_ASAP7_75t_L g1480 ( 
.A(n_1474),
.Y(n_1480)
);

NOR2xp67_ASAP7_75t_L g1481 ( 
.A(n_1474),
.B(n_1392),
.Y(n_1481)
);

OR2x2_ASAP7_75t_L g1482 ( 
.A(n_1457),
.B(n_1359),
.Y(n_1482)
);

BUFx2_ASAP7_75t_L g1483 ( 
.A(n_1429),
.Y(n_1483)
);

NAND2xp5_ASAP7_75t_L g1484 ( 
.A(n_1429),
.B(n_1351),
.Y(n_1484)
);

INVxp67_ASAP7_75t_SL g1485 ( 
.A(n_1463),
.Y(n_1485)
);

AOI22xp33_ASAP7_75t_SL g1486 ( 
.A1(n_1446),
.A2(n_1415),
.B1(n_1387),
.B2(n_1381),
.Y(n_1486)
);

AND2x2_ASAP7_75t_L g1487 ( 
.A(n_1462),
.B(n_1342),
.Y(n_1487)
);

INVx2_ASAP7_75t_L g1488 ( 
.A(n_1434),
.Y(n_1488)
);

NOR2xp33_ASAP7_75t_L g1489 ( 
.A(n_1433),
.B(n_1409),
.Y(n_1489)
);

INVxp67_ASAP7_75t_L g1490 ( 
.A(n_1463),
.Y(n_1490)
);

INVxp67_ASAP7_75t_L g1491 ( 
.A(n_1468),
.Y(n_1491)
);

NAND2xp5_ASAP7_75t_L g1492 ( 
.A(n_1454),
.B(n_1381),
.Y(n_1492)
);

OR2x2_ASAP7_75t_L g1493 ( 
.A(n_1465),
.B(n_1340),
.Y(n_1493)
);

NAND2xp5_ASAP7_75t_L g1494 ( 
.A(n_1454),
.B(n_1340),
.Y(n_1494)
);

AND2x2_ASAP7_75t_L g1495 ( 
.A(n_1447),
.B(n_1346),
.Y(n_1495)
);

AOI22xp33_ASAP7_75t_L g1496 ( 
.A1(n_1417),
.A2(n_1415),
.B1(n_1374),
.B2(n_1366),
.Y(n_1496)
);

AND2x2_ASAP7_75t_L g1497 ( 
.A(n_1449),
.B(n_1346),
.Y(n_1497)
);

INVxp67_ASAP7_75t_SL g1498 ( 
.A(n_1471),
.Y(n_1498)
);

AOI22xp33_ASAP7_75t_L g1499 ( 
.A1(n_1453),
.A2(n_1415),
.B1(n_1374),
.B2(n_1366),
.Y(n_1499)
);

AND2x2_ASAP7_75t_L g1500 ( 
.A(n_1466),
.B(n_1347),
.Y(n_1500)
);

INVx1_ASAP7_75t_L g1501 ( 
.A(n_1469),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_1450),
.Y(n_1502)
);

NAND2xp5_ASAP7_75t_L g1503 ( 
.A(n_1459),
.B(n_1338),
.Y(n_1503)
);

INVx1_ASAP7_75t_L g1504 ( 
.A(n_1450),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_1467),
.Y(n_1505)
);

INVx1_ASAP7_75t_L g1506 ( 
.A(n_1467),
.Y(n_1506)
);

AND2x2_ASAP7_75t_L g1507 ( 
.A(n_1461),
.B(n_1415),
.Y(n_1507)
);

INVx1_ASAP7_75t_L g1508 ( 
.A(n_1456),
.Y(n_1508)
);

AND2x2_ASAP7_75t_L g1509 ( 
.A(n_1470),
.B(n_1358),
.Y(n_1509)
);

INVx4_ASAP7_75t_L g1510 ( 
.A(n_1419),
.Y(n_1510)
);

INVx2_ASAP7_75t_SL g1511 ( 
.A(n_1488),
.Y(n_1511)
);

NAND2xp5_ASAP7_75t_L g1512 ( 
.A(n_1490),
.B(n_1459),
.Y(n_1512)
);

AO21x2_ASAP7_75t_L g1513 ( 
.A1(n_1492),
.A2(n_1446),
.B(n_1471),
.Y(n_1513)
);

NOR2x1_ASAP7_75t_L g1514 ( 
.A(n_1481),
.B(n_1430),
.Y(n_1514)
);

INVx2_ASAP7_75t_L g1515 ( 
.A(n_1502),
.Y(n_1515)
);

AND2x4_ASAP7_75t_L g1516 ( 
.A(n_1481),
.B(n_1470),
.Y(n_1516)
);

NAND4xp25_ASAP7_75t_L g1517 ( 
.A(n_1486),
.B(n_1435),
.C(n_1443),
.D(n_1464),
.Y(n_1517)
);

INVx2_ASAP7_75t_L g1518 ( 
.A(n_1502),
.Y(n_1518)
);

AND2x2_ASAP7_75t_L g1519 ( 
.A(n_1498),
.B(n_1444),
.Y(n_1519)
);

NOR2x1_ASAP7_75t_L g1520 ( 
.A(n_1483),
.B(n_1430),
.Y(n_1520)
);

NAND2xp33_ASAP7_75t_SL g1521 ( 
.A(n_1510),
.B(n_1441),
.Y(n_1521)
);

AND2x4_ASAP7_75t_L g1522 ( 
.A(n_1507),
.B(n_1460),
.Y(n_1522)
);

AOI21xp33_ASAP7_75t_SL g1523 ( 
.A1(n_1478),
.A2(n_1435),
.B(n_1432),
.Y(n_1523)
);

AND2x2_ASAP7_75t_L g1524 ( 
.A(n_1490),
.B(n_1444),
.Y(n_1524)
);

NAND2xp5_ASAP7_75t_L g1525 ( 
.A(n_1485),
.B(n_1473),
.Y(n_1525)
);

BUFx2_ASAP7_75t_L g1526 ( 
.A(n_1483),
.Y(n_1526)
);

INVx2_ASAP7_75t_L g1527 ( 
.A(n_1504),
.Y(n_1527)
);

INVxp67_ASAP7_75t_SL g1528 ( 
.A(n_1480),
.Y(n_1528)
);

INVx1_ASAP7_75t_L g1529 ( 
.A(n_1488),
.Y(n_1529)
);

INVx2_ASAP7_75t_SL g1530 ( 
.A(n_1488),
.Y(n_1530)
);

INVx1_ASAP7_75t_L g1531 ( 
.A(n_1484),
.Y(n_1531)
);

BUFx2_ASAP7_75t_L g1532 ( 
.A(n_1479),
.Y(n_1532)
);

BUFx3_ASAP7_75t_L g1533 ( 
.A(n_1479),
.Y(n_1533)
);

NAND2xp5_ASAP7_75t_L g1534 ( 
.A(n_1505),
.B(n_1473),
.Y(n_1534)
);

AOI221x1_ASAP7_75t_L g1535 ( 
.A1(n_1508),
.A2(n_1439),
.B1(n_1440),
.B2(n_1445),
.C(n_1472),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_1484),
.Y(n_1536)
);

AOI221xp5_ASAP7_75t_L g1537 ( 
.A1(n_1505),
.A2(n_1464),
.B1(n_1443),
.B2(n_1472),
.C(n_1426),
.Y(n_1537)
);

OAI33xp33_ASAP7_75t_L g1538 ( 
.A1(n_1506),
.A2(n_1439),
.A3(n_1421),
.B1(n_1396),
.B2(n_1341),
.B3(n_1345),
.Y(n_1538)
);

INVx2_ASAP7_75t_L g1539 ( 
.A(n_1504),
.Y(n_1539)
);

OAI211xp5_ASAP7_75t_L g1540 ( 
.A1(n_1486),
.A2(n_1426),
.B(n_1440),
.C(n_1437),
.Y(n_1540)
);

AND2x2_ASAP7_75t_L g1541 ( 
.A(n_1487),
.B(n_1441),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_1477),
.Y(n_1542)
);

OAI222xp33_ASAP7_75t_L g1543 ( 
.A1(n_1476),
.A2(n_1460),
.B1(n_1414),
.B2(n_1448),
.C1(n_1451),
.C2(n_1455),
.Y(n_1543)
);

INVx1_ASAP7_75t_L g1544 ( 
.A(n_1477),
.Y(n_1544)
);

BUFx2_ASAP7_75t_L g1545 ( 
.A(n_1479),
.Y(n_1545)
);

AOI21xp5_ASAP7_75t_SL g1546 ( 
.A1(n_1494),
.A2(n_1438),
.B(n_1436),
.Y(n_1546)
);

OR2x2_ASAP7_75t_L g1547 ( 
.A(n_1506),
.B(n_1442),
.Y(n_1547)
);

OAI321xp33_ASAP7_75t_L g1548 ( 
.A1(n_1492),
.A2(n_1436),
.A3(n_1451),
.B1(n_1448),
.B2(n_1425),
.C(n_1455),
.Y(n_1548)
);

AND2x2_ASAP7_75t_L g1549 ( 
.A(n_1495),
.B(n_1431),
.Y(n_1549)
);

AOI221xp5_ASAP7_75t_L g1550 ( 
.A1(n_1503),
.A2(n_1424),
.B1(n_1428),
.B2(n_1414),
.C(n_1422),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_1542),
.Y(n_1551)
);

AND2x2_ASAP7_75t_L g1552 ( 
.A(n_1532),
.B(n_1480),
.Y(n_1552)
);

AND2x2_ASAP7_75t_L g1553 ( 
.A(n_1532),
.B(n_1495),
.Y(n_1553)
);

OR2x2_ASAP7_75t_L g1554 ( 
.A(n_1534),
.B(n_1493),
.Y(n_1554)
);

OR2x2_ASAP7_75t_L g1555 ( 
.A(n_1534),
.B(n_1493),
.Y(n_1555)
);

OR2x2_ASAP7_75t_L g1556 ( 
.A(n_1525),
.B(n_1482),
.Y(n_1556)
);

AND2x2_ASAP7_75t_L g1557 ( 
.A(n_1545),
.B(n_1497),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_1542),
.Y(n_1558)
);

NAND2x1_ASAP7_75t_SL g1559 ( 
.A(n_1514),
.B(n_1479),
.Y(n_1559)
);

INVx1_ASAP7_75t_L g1560 ( 
.A(n_1544),
.Y(n_1560)
);

NOR2xp67_ASAP7_75t_L g1561 ( 
.A(n_1540),
.B(n_1494),
.Y(n_1561)
);

AND2x2_ASAP7_75t_L g1562 ( 
.A(n_1545),
.B(n_1497),
.Y(n_1562)
);

INVx2_ASAP7_75t_SL g1563 ( 
.A(n_1516),
.Y(n_1563)
);

INVx2_ASAP7_75t_L g1564 ( 
.A(n_1511),
.Y(n_1564)
);

INVx2_ASAP7_75t_L g1565 ( 
.A(n_1511),
.Y(n_1565)
);

NAND2xp5_ASAP7_75t_L g1566 ( 
.A(n_1531),
.B(n_1501),
.Y(n_1566)
);

AND2x2_ASAP7_75t_L g1567 ( 
.A(n_1514),
.B(n_1491),
.Y(n_1567)
);

NAND2xp5_ASAP7_75t_L g1568 ( 
.A(n_1531),
.B(n_1501),
.Y(n_1568)
);

HB1xp67_ASAP7_75t_L g1569 ( 
.A(n_1536),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_1544),
.Y(n_1570)
);

INVx1_ASAP7_75t_L g1571 ( 
.A(n_1529),
.Y(n_1571)
);

INVx1_ASAP7_75t_L g1572 ( 
.A(n_1529),
.Y(n_1572)
);

AND2x2_ASAP7_75t_L g1573 ( 
.A(n_1519),
.B(n_1491),
.Y(n_1573)
);

INVx1_ASAP7_75t_L g1574 ( 
.A(n_1536),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_1515),
.Y(n_1575)
);

NOR3xp33_ASAP7_75t_SL g1576 ( 
.A(n_1517),
.B(n_1489),
.C(n_1422),
.Y(n_1576)
);

NAND2x1p5_ASAP7_75t_L g1577 ( 
.A(n_1520),
.B(n_1418),
.Y(n_1577)
);

AND2x2_ASAP7_75t_L g1578 ( 
.A(n_1519),
.B(n_1526),
.Y(n_1578)
);

INVx1_ASAP7_75t_L g1579 ( 
.A(n_1515),
.Y(n_1579)
);

AND2x2_ASAP7_75t_L g1580 ( 
.A(n_1526),
.B(n_1500),
.Y(n_1580)
);

INVx2_ASAP7_75t_L g1581 ( 
.A(n_1511),
.Y(n_1581)
);

HB1xp67_ASAP7_75t_L g1582 ( 
.A(n_1547),
.Y(n_1582)
);

AND2x2_ASAP7_75t_L g1583 ( 
.A(n_1520),
.B(n_1500),
.Y(n_1583)
);

OAI22xp5_ASAP7_75t_L g1584 ( 
.A1(n_1537),
.A2(n_1499),
.B1(n_1496),
.B2(n_1475),
.Y(n_1584)
);

HB1xp67_ASAP7_75t_L g1585 ( 
.A(n_1547),
.Y(n_1585)
);

AND2x2_ASAP7_75t_L g1586 ( 
.A(n_1528),
.B(n_1509),
.Y(n_1586)
);

AOI31xp33_ASAP7_75t_L g1587 ( 
.A1(n_1550),
.A2(n_1422),
.A3(n_1419),
.B(n_1427),
.Y(n_1587)
);

CKINVDCx16_ASAP7_75t_R g1588 ( 
.A(n_1549),
.Y(n_1588)
);

INVx1_ASAP7_75t_L g1589 ( 
.A(n_1551),
.Y(n_1589)
);

INVxp67_ASAP7_75t_SL g1590 ( 
.A(n_1561),
.Y(n_1590)
);

OR2x2_ASAP7_75t_L g1591 ( 
.A(n_1554),
.B(n_1512),
.Y(n_1591)
);

AND2x2_ASAP7_75t_L g1592 ( 
.A(n_1588),
.B(n_1533),
.Y(n_1592)
);

INVx2_ASAP7_75t_L g1593 ( 
.A(n_1564),
.Y(n_1593)
);

OR2x2_ASAP7_75t_L g1594 ( 
.A(n_1554),
.B(n_1512),
.Y(n_1594)
);

INVx3_ASAP7_75t_L g1595 ( 
.A(n_1588),
.Y(n_1595)
);

INVx2_ASAP7_75t_L g1596 ( 
.A(n_1564),
.Y(n_1596)
);

NAND2xp5_ASAP7_75t_L g1597 ( 
.A(n_1556),
.B(n_1525),
.Y(n_1597)
);

NOR2xp33_ASAP7_75t_L g1598 ( 
.A(n_1555),
.B(n_1523),
.Y(n_1598)
);

OAI21xp5_ASAP7_75t_L g1599 ( 
.A1(n_1561),
.A2(n_1523),
.B(n_1517),
.Y(n_1599)
);

INVx1_ASAP7_75t_L g1600 ( 
.A(n_1551),
.Y(n_1600)
);

NAND2xp5_ASAP7_75t_L g1601 ( 
.A(n_1556),
.B(n_1530),
.Y(n_1601)
);

INVx1_ASAP7_75t_L g1602 ( 
.A(n_1558),
.Y(n_1602)
);

NAND2xp5_ASAP7_75t_L g1603 ( 
.A(n_1555),
.B(n_1530),
.Y(n_1603)
);

NAND2xp5_ASAP7_75t_L g1604 ( 
.A(n_1569),
.B(n_1530),
.Y(n_1604)
);

INVx1_ASAP7_75t_L g1605 ( 
.A(n_1558),
.Y(n_1605)
);

INVx2_ASAP7_75t_L g1606 ( 
.A(n_1564),
.Y(n_1606)
);

AND2x2_ASAP7_75t_L g1607 ( 
.A(n_1578),
.B(n_1533),
.Y(n_1607)
);

INVx1_ASAP7_75t_SL g1608 ( 
.A(n_1578),
.Y(n_1608)
);

OR2x2_ASAP7_75t_L g1609 ( 
.A(n_1582),
.B(n_1482),
.Y(n_1609)
);

NAND2xp5_ASAP7_75t_L g1610 ( 
.A(n_1574),
.B(n_1515),
.Y(n_1610)
);

NAND3xp33_ASAP7_75t_L g1611 ( 
.A(n_1576),
.B(n_1550),
.C(n_1540),
.Y(n_1611)
);

NAND2xp5_ASAP7_75t_L g1612 ( 
.A(n_1574),
.B(n_1518),
.Y(n_1612)
);

AND2x2_ASAP7_75t_L g1613 ( 
.A(n_1578),
.B(n_1533),
.Y(n_1613)
);

AND2x2_ASAP7_75t_L g1614 ( 
.A(n_1553),
.B(n_1524),
.Y(n_1614)
);

AND2x2_ASAP7_75t_L g1615 ( 
.A(n_1553),
.B(n_1524),
.Y(n_1615)
);

AND2x2_ASAP7_75t_L g1616 ( 
.A(n_1553),
.B(n_1549),
.Y(n_1616)
);

INVx1_ASAP7_75t_L g1617 ( 
.A(n_1560),
.Y(n_1617)
);

HB1xp67_ASAP7_75t_L g1618 ( 
.A(n_1573),
.Y(n_1618)
);

INVx1_ASAP7_75t_L g1619 ( 
.A(n_1560),
.Y(n_1619)
);

INVx2_ASAP7_75t_L g1620 ( 
.A(n_1565),
.Y(n_1620)
);

INVx1_ASAP7_75t_L g1621 ( 
.A(n_1570),
.Y(n_1621)
);

INVx1_ASAP7_75t_L g1622 ( 
.A(n_1570),
.Y(n_1622)
);

NAND2xp5_ASAP7_75t_L g1623 ( 
.A(n_1585),
.B(n_1576),
.Y(n_1623)
);

AND2x2_ASAP7_75t_L g1624 ( 
.A(n_1557),
.B(n_1541),
.Y(n_1624)
);

NAND2xp5_ASAP7_75t_L g1625 ( 
.A(n_1566),
.B(n_1568),
.Y(n_1625)
);

NAND2xp5_ASAP7_75t_L g1626 ( 
.A(n_1566),
.B(n_1568),
.Y(n_1626)
);

INVx2_ASAP7_75t_L g1627 ( 
.A(n_1565),
.Y(n_1627)
);

INVx1_ASAP7_75t_L g1628 ( 
.A(n_1571),
.Y(n_1628)
);

OR2x2_ASAP7_75t_L g1629 ( 
.A(n_1584),
.B(n_1518),
.Y(n_1629)
);

HB1xp67_ASAP7_75t_L g1630 ( 
.A(n_1571),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_1630),
.Y(n_1631)
);

OR2x2_ASAP7_75t_L g1632 ( 
.A(n_1591),
.B(n_1584),
.Y(n_1632)
);

INVx2_ASAP7_75t_L g1633 ( 
.A(n_1595),
.Y(n_1633)
);

AND2x4_ASAP7_75t_L g1634 ( 
.A(n_1595),
.B(n_1563),
.Y(n_1634)
);

NAND2xp5_ASAP7_75t_L g1635 ( 
.A(n_1598),
.B(n_1573),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_1589),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_1589),
.Y(n_1637)
);

INVx1_ASAP7_75t_L g1638 ( 
.A(n_1600),
.Y(n_1638)
);

INVx1_ASAP7_75t_L g1639 ( 
.A(n_1630),
.Y(n_1639)
);

NOR2xp33_ASAP7_75t_L g1640 ( 
.A(n_1597),
.B(n_1590),
.Y(n_1640)
);

AND2x2_ASAP7_75t_L g1641 ( 
.A(n_1592),
.B(n_1563),
.Y(n_1641)
);

OR2x2_ASAP7_75t_L g1642 ( 
.A(n_1591),
.B(n_1587),
.Y(n_1642)
);

OR2x2_ASAP7_75t_L g1643 ( 
.A(n_1594),
.B(n_1587),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_1600),
.Y(n_1644)
);

AND2x2_ASAP7_75t_L g1645 ( 
.A(n_1592),
.B(n_1563),
.Y(n_1645)
);

INVx2_ASAP7_75t_L g1646 ( 
.A(n_1595),
.Y(n_1646)
);

NAND2xp5_ASAP7_75t_L g1647 ( 
.A(n_1599),
.B(n_1573),
.Y(n_1647)
);

NAND2xp5_ASAP7_75t_SL g1648 ( 
.A(n_1611),
.B(n_1567),
.Y(n_1648)
);

NAND2xp5_ASAP7_75t_L g1649 ( 
.A(n_1599),
.B(n_1590),
.Y(n_1649)
);

INVx1_ASAP7_75t_L g1650 ( 
.A(n_1602),
.Y(n_1650)
);

AOI22xp5_ASAP7_75t_L g1651 ( 
.A1(n_1611),
.A2(n_1513),
.B1(n_1537),
.B2(n_1538),
.Y(n_1651)
);

NAND2xp5_ASAP7_75t_L g1652 ( 
.A(n_1597),
.B(n_1552),
.Y(n_1652)
);

AND2x2_ASAP7_75t_L g1653 ( 
.A(n_1595),
.B(n_1567),
.Y(n_1653)
);

AND2x2_ASAP7_75t_L g1654 ( 
.A(n_1616),
.B(n_1567),
.Y(n_1654)
);

NOR2x2_ASAP7_75t_L g1655 ( 
.A(n_1593),
.B(n_1565),
.Y(n_1655)
);

AND2x2_ASAP7_75t_L g1656 ( 
.A(n_1616),
.B(n_1552),
.Y(n_1656)
);

NAND2xp5_ASAP7_75t_L g1657 ( 
.A(n_1618),
.B(n_1552),
.Y(n_1657)
);

AOI32xp33_ASAP7_75t_L g1658 ( 
.A1(n_1623),
.A2(n_1548),
.A3(n_1586),
.B1(n_1583),
.B2(n_1581),
.Y(n_1658)
);

NAND2xp5_ASAP7_75t_L g1659 ( 
.A(n_1608),
.B(n_1586),
.Y(n_1659)
);

NAND2xp5_ASAP7_75t_L g1660 ( 
.A(n_1608),
.B(n_1586),
.Y(n_1660)
);

NOR2xp33_ASAP7_75t_L g1661 ( 
.A(n_1594),
.B(n_1557),
.Y(n_1661)
);

NAND2xp5_ASAP7_75t_L g1662 ( 
.A(n_1623),
.B(n_1557),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_1602),
.Y(n_1663)
);

INVx2_ASAP7_75t_L g1664 ( 
.A(n_1593),
.Y(n_1664)
);

INVx1_ASAP7_75t_L g1665 ( 
.A(n_1605),
.Y(n_1665)
);

AOI22xp5_ASAP7_75t_L g1666 ( 
.A1(n_1651),
.A2(n_1513),
.B1(n_1629),
.B2(n_1577),
.Y(n_1666)
);

AOI21xp5_ASAP7_75t_L g1667 ( 
.A1(n_1648),
.A2(n_1629),
.B(n_1546),
.Y(n_1667)
);

OAI22x1_ASAP7_75t_L g1668 ( 
.A1(n_1648),
.A2(n_1607),
.B1(n_1613),
.B2(n_1577),
.Y(n_1668)
);

AOI22xp5_ASAP7_75t_L g1669 ( 
.A1(n_1649),
.A2(n_1513),
.B1(n_1632),
.B2(n_1642),
.Y(n_1669)
);

AND2x4_ASAP7_75t_L g1670 ( 
.A(n_1641),
.B(n_1614),
.Y(n_1670)
);

INVx2_ASAP7_75t_L g1671 ( 
.A(n_1655),
.Y(n_1671)
);

INVxp67_ASAP7_75t_L g1672 ( 
.A(n_1640),
.Y(n_1672)
);

INVx1_ASAP7_75t_L g1673 ( 
.A(n_1631),
.Y(n_1673)
);

AOI21xp5_ASAP7_75t_L g1674 ( 
.A1(n_1647),
.A2(n_1546),
.B(n_1604),
.Y(n_1674)
);

AOI22xp5_ASAP7_75t_L g1675 ( 
.A1(n_1632),
.A2(n_1513),
.B1(n_1577),
.B2(n_1522),
.Y(n_1675)
);

OR2x2_ASAP7_75t_L g1676 ( 
.A(n_1652),
.B(n_1609),
.Y(n_1676)
);

NAND4xp25_ASAP7_75t_L g1677 ( 
.A(n_1658),
.B(n_1535),
.C(n_1607),
.D(n_1613),
.Y(n_1677)
);

INVx1_ASAP7_75t_SL g1678 ( 
.A(n_1633),
.Y(n_1678)
);

NAND2xp5_ASAP7_75t_L g1679 ( 
.A(n_1661),
.B(n_1614),
.Y(n_1679)
);

AOI21xp33_ASAP7_75t_L g1680 ( 
.A1(n_1642),
.A2(n_1627),
.B(n_1606),
.Y(n_1680)
);

OAI22xp5_ASAP7_75t_L g1681 ( 
.A1(n_1643),
.A2(n_1577),
.B1(n_1615),
.B2(n_1624),
.Y(n_1681)
);

INVx2_ASAP7_75t_L g1682 ( 
.A(n_1655),
.Y(n_1682)
);

INVxp67_ASAP7_75t_SL g1683 ( 
.A(n_1633),
.Y(n_1683)
);

OAI21xp33_ASAP7_75t_SL g1684 ( 
.A1(n_1643),
.A2(n_1615),
.B(n_1559),
.Y(n_1684)
);

NAND2xp5_ASAP7_75t_L g1685 ( 
.A(n_1656),
.B(n_1635),
.Y(n_1685)
);

OR2x2_ASAP7_75t_L g1686 ( 
.A(n_1662),
.B(n_1659),
.Y(n_1686)
);

NAND2xp5_ASAP7_75t_L g1687 ( 
.A(n_1656),
.B(n_1625),
.Y(n_1687)
);

O2A1O1Ixp5_ASAP7_75t_L g1688 ( 
.A1(n_1646),
.A2(n_1606),
.B(n_1627),
.C(n_1593),
.Y(n_1688)
);

INVx1_ASAP7_75t_L g1689 ( 
.A(n_1631),
.Y(n_1689)
);

AOI21xp5_ASAP7_75t_L g1690 ( 
.A1(n_1657),
.A2(n_1604),
.B(n_1625),
.Y(n_1690)
);

INVx2_ASAP7_75t_L g1691 ( 
.A(n_1670),
.Y(n_1691)
);

OAI22xp5_ASAP7_75t_L g1692 ( 
.A1(n_1666),
.A2(n_1660),
.B1(n_1654),
.B2(n_1641),
.Y(n_1692)
);

HB1xp67_ASAP7_75t_L g1693 ( 
.A(n_1678),
.Y(n_1693)
);

OR2x2_ASAP7_75t_L g1694 ( 
.A(n_1687),
.B(n_1601),
.Y(n_1694)
);

NAND4xp25_ASAP7_75t_SL g1695 ( 
.A(n_1684),
.B(n_1654),
.C(n_1653),
.D(n_1645),
.Y(n_1695)
);

AND2x4_ASAP7_75t_L g1696 ( 
.A(n_1670),
.B(n_1645),
.Y(n_1696)
);

A2O1A1Ixp33_ASAP7_75t_L g1697 ( 
.A1(n_1667),
.A2(n_1548),
.B(n_1559),
.C(n_1653),
.Y(n_1697)
);

A2O1A1Ixp33_ASAP7_75t_L g1698 ( 
.A1(n_1677),
.A2(n_1664),
.B(n_1603),
.C(n_1626),
.Y(n_1698)
);

NAND2xp5_ASAP7_75t_L g1699 ( 
.A(n_1672),
.B(n_1639),
.Y(n_1699)
);

OAI32xp33_ASAP7_75t_L g1700 ( 
.A1(n_1677),
.A2(n_1639),
.A3(n_1646),
.B1(n_1603),
.B2(n_1601),
.Y(n_1700)
);

INVx1_ASAP7_75t_L g1701 ( 
.A(n_1673),
.Y(n_1701)
);

AOI22xp33_ASAP7_75t_L g1702 ( 
.A1(n_1671),
.A2(n_1664),
.B1(n_1634),
.B2(n_1620),
.Y(n_1702)
);

AOI322xp5_ASAP7_75t_L g1703 ( 
.A1(n_1669),
.A2(n_1682),
.A3(n_1680),
.B1(n_1675),
.B2(n_1678),
.C1(n_1679),
.C2(n_1683),
.Y(n_1703)
);

OAI22xp5_ASAP7_75t_L g1704 ( 
.A1(n_1674),
.A2(n_1676),
.B1(n_1686),
.B2(n_1685),
.Y(n_1704)
);

NAND2xp5_ASAP7_75t_L g1705 ( 
.A(n_1690),
.B(n_1626),
.Y(n_1705)
);

NAND2xp5_ASAP7_75t_SL g1706 ( 
.A(n_1668),
.B(n_1634),
.Y(n_1706)
);

INVxp67_ASAP7_75t_L g1707 ( 
.A(n_1689),
.Y(n_1707)
);

NAND2xp5_ASAP7_75t_L g1708 ( 
.A(n_1681),
.B(n_1636),
.Y(n_1708)
);

NAND3xp33_ASAP7_75t_L g1709 ( 
.A(n_1688),
.B(n_1634),
.C(n_1663),
.Y(n_1709)
);

INVx1_ASAP7_75t_L g1710 ( 
.A(n_1693),
.Y(n_1710)
);

AND2x2_ASAP7_75t_L g1711 ( 
.A(n_1696),
.B(n_1624),
.Y(n_1711)
);

AND2x2_ASAP7_75t_L g1712 ( 
.A(n_1696),
.B(n_1637),
.Y(n_1712)
);

INVx1_ASAP7_75t_L g1713 ( 
.A(n_1699),
.Y(n_1713)
);

INVx1_ASAP7_75t_L g1714 ( 
.A(n_1701),
.Y(n_1714)
);

NAND2xp5_ASAP7_75t_L g1715 ( 
.A(n_1705),
.B(n_1638),
.Y(n_1715)
);

XNOR2xp5_ASAP7_75t_L g1716 ( 
.A(n_1704),
.B(n_1535),
.Y(n_1716)
);

AOI21xp5_ASAP7_75t_L g1717 ( 
.A1(n_1698),
.A2(n_1665),
.B(n_1650),
.Y(n_1717)
);

AND2x2_ASAP7_75t_L g1718 ( 
.A(n_1691),
.B(n_1644),
.Y(n_1718)
);

INVxp67_ASAP7_75t_L g1719 ( 
.A(n_1708),
.Y(n_1719)
);

OAI22xp5_ASAP7_75t_L g1720 ( 
.A1(n_1697),
.A2(n_1609),
.B1(n_1583),
.B2(n_1622),
.Y(n_1720)
);

INVx1_ASAP7_75t_L g1721 ( 
.A(n_1710),
.Y(n_1721)
);

NOR3xp33_ASAP7_75t_L g1722 ( 
.A(n_1719),
.B(n_1700),
.C(n_1704),
.Y(n_1722)
);

NAND2xp5_ASAP7_75t_L g1723 ( 
.A(n_1711),
.B(n_1703),
.Y(n_1723)
);

NAND2xp33_ASAP7_75t_SL g1724 ( 
.A(n_1711),
.B(n_1706),
.Y(n_1724)
);

OAI322xp33_ASAP7_75t_L g1725 ( 
.A1(n_1716),
.A2(n_1692),
.A3(n_1707),
.B1(n_1709),
.B2(n_1694),
.C1(n_1695),
.C2(n_1702),
.Y(n_1725)
);

INVxp33_ASAP7_75t_L g1726 ( 
.A(n_1712),
.Y(n_1726)
);

NAND2xp5_ASAP7_75t_L g1727 ( 
.A(n_1712),
.B(n_1605),
.Y(n_1727)
);

NAND2xp5_ASAP7_75t_L g1728 ( 
.A(n_1718),
.B(n_1617),
.Y(n_1728)
);

NOR2xp33_ASAP7_75t_L g1729 ( 
.A(n_1715),
.B(n_1617),
.Y(n_1729)
);

OAI321xp33_ASAP7_75t_L g1730 ( 
.A1(n_1720),
.A2(n_1620),
.A3(n_1627),
.B1(n_1596),
.B2(n_1606),
.C(n_1621),
.Y(n_1730)
);

BUFx4f_ASAP7_75t_L g1731 ( 
.A(n_1713),
.Y(n_1731)
);

AOI322xp5_ASAP7_75t_L g1732 ( 
.A1(n_1723),
.A2(n_1714),
.A3(n_1718),
.B1(n_1717),
.B2(n_1620),
.C1(n_1596),
.C2(n_1612),
.Y(n_1732)
);

OAI211xp5_ASAP7_75t_SL g1733 ( 
.A1(n_1722),
.A2(n_1596),
.B(n_1622),
.C(n_1621),
.Y(n_1733)
);

OAI211xp5_ASAP7_75t_L g1734 ( 
.A1(n_1724),
.A2(n_1619),
.B(n_1628),
.C(n_1521),
.Y(n_1734)
);

OAI21xp33_ASAP7_75t_L g1735 ( 
.A1(n_1726),
.A2(n_1619),
.B(n_1628),
.Y(n_1735)
);

OAI221xp5_ASAP7_75t_L g1736 ( 
.A1(n_1731),
.A2(n_1612),
.B1(n_1610),
.B2(n_1575),
.C(n_1579),
.Y(n_1736)
);

AOI221xp5_ASAP7_75t_L g1737 ( 
.A1(n_1733),
.A2(n_1725),
.B1(n_1730),
.B2(n_1729),
.C(n_1731),
.Y(n_1737)
);

AOI22xp5_ASAP7_75t_L g1738 ( 
.A1(n_1736),
.A2(n_1721),
.B1(n_1728),
.B2(n_1727),
.Y(n_1738)
);

AOI221xp5_ASAP7_75t_L g1739 ( 
.A1(n_1735),
.A2(n_1543),
.B1(n_1610),
.B2(n_1527),
.C(n_1518),
.Y(n_1739)
);

AOI22xp5_ASAP7_75t_L g1740 ( 
.A1(n_1734),
.A2(n_1579),
.B1(n_1575),
.B2(n_1527),
.Y(n_1740)
);

AOI21xp5_ASAP7_75t_L g1741 ( 
.A1(n_1732),
.A2(n_1581),
.B(n_1572),
.Y(n_1741)
);

O2A1O1Ixp33_ASAP7_75t_L g1742 ( 
.A1(n_1733),
.A2(n_1543),
.B(n_1581),
.C(n_1527),
.Y(n_1742)
);

INVx2_ASAP7_75t_L g1743 ( 
.A(n_1738),
.Y(n_1743)
);

NAND2xp5_ASAP7_75t_L g1744 ( 
.A(n_1737),
.B(n_1539),
.Y(n_1744)
);

AOI22xp5_ASAP7_75t_L g1745 ( 
.A1(n_1739),
.A2(n_1539),
.B1(n_1516),
.B2(n_1583),
.Y(n_1745)
);

INVx1_ASAP7_75t_L g1746 ( 
.A(n_1741),
.Y(n_1746)
);

INVx2_ASAP7_75t_SL g1747 ( 
.A(n_1740),
.Y(n_1747)
);

AND2x4_ASAP7_75t_L g1748 ( 
.A(n_1747),
.B(n_1580),
.Y(n_1748)
);

NAND3xp33_ASAP7_75t_SL g1749 ( 
.A(n_1743),
.B(n_1742),
.C(n_1422),
.Y(n_1749)
);

XOR2xp5_ASAP7_75t_L g1750 ( 
.A(n_1744),
.B(n_1522),
.Y(n_1750)
);

NOR3xp33_ASAP7_75t_L g1751 ( 
.A(n_1749),
.B(n_1746),
.C(n_1745),
.Y(n_1751)
);

INVx1_ASAP7_75t_L g1752 ( 
.A(n_1751),
.Y(n_1752)
);

INVx1_ASAP7_75t_L g1753 ( 
.A(n_1752),
.Y(n_1753)
);

INVxp67_ASAP7_75t_L g1754 ( 
.A(n_1753),
.Y(n_1754)
);

OAI22xp5_ASAP7_75t_L g1755 ( 
.A1(n_1754),
.A2(n_1748),
.B1(n_1750),
.B2(n_1539),
.Y(n_1755)
);

INVx1_ASAP7_75t_L g1756 ( 
.A(n_1755),
.Y(n_1756)
);

AOI21x1_ASAP7_75t_L g1757 ( 
.A1(n_1756),
.A2(n_1580),
.B(n_1562),
.Y(n_1757)
);

INVxp67_ASAP7_75t_L g1758 ( 
.A(n_1757),
.Y(n_1758)
);

XOR2xp5_ASAP7_75t_L g1759 ( 
.A(n_1757),
.B(n_1423),
.Y(n_1759)
);

OAI221xp5_ASAP7_75t_L g1760 ( 
.A1(n_1758),
.A2(n_1572),
.B1(n_1580),
.B2(n_1562),
.C(n_1408),
.Y(n_1760)
);

AOI211xp5_ASAP7_75t_L g1761 ( 
.A1(n_1760),
.A2(n_1759),
.B(n_1562),
.C(n_1516),
.Y(n_1761)
);


endmodule