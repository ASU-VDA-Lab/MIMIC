module fake_jpeg_30661_n_539 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_539);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_539;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_387;
wire n_270;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_349;
wire n_21;
wire n_288;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx3_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

INVx8_ASAP7_75t_SL g20 ( 
.A(n_1),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_7),
.Y(n_22)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

CKINVDCx16_ASAP7_75t_R g25 ( 
.A(n_16),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_13),
.Y(n_27)
);

INVx13_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

INVx13_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_10),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_2),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_15),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_13),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_8),
.Y(n_38)
);

INVx11_ASAP7_75t_SL g39 ( 
.A(n_16),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_7),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_17),
.Y(n_41)
);

CKINVDCx14_ASAP7_75t_R g42 ( 
.A(n_6),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_3),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_15),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_12),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_1),
.Y(n_46)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_14),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_10),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_11),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_16),
.Y(n_50)
);

BUFx5_ASAP7_75t_L g51 ( 
.A(n_5),
.Y(n_51)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_19),
.Y(n_52)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_52),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_26),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_53),
.Y(n_105)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_19),
.Y(n_54)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_54),
.Y(n_116)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_26),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_55),
.Y(n_123)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_56),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_26),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_57),
.Y(n_125)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_23),
.Y(n_58)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_58),
.Y(n_106)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_19),
.Y(n_59)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_59),
.Y(n_140)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_23),
.Y(n_60)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_60),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_26),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_61),
.Y(n_132)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_51),
.Y(n_62)
);

INVx5_ASAP7_75t_L g122 ( 
.A(n_62),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_32),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_63),
.Y(n_137)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_32),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_64),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_32),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_65),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g66 ( 
.A(n_40),
.B(n_9),
.C(n_1),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g135 ( 
.A(n_66),
.B(n_70),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_32),
.Y(n_67)
);

INVx6_ASAP7_75t_L g117 ( 
.A(n_67),
.Y(n_117)
);

INVx5_ASAP7_75t_L g68 ( 
.A(n_51),
.Y(n_68)
);

INVx5_ASAP7_75t_L g128 ( 
.A(n_68),
.Y(n_128)
);

INVx11_ASAP7_75t_L g69 ( 
.A(n_39),
.Y(n_69)
);

INVx6_ASAP7_75t_L g151 ( 
.A(n_69),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g70 ( 
.A(n_40),
.B(n_9),
.C(n_2),
.Y(n_70)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_47),
.Y(n_71)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_71),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_41),
.Y(n_72)
);

INVx5_ASAP7_75t_L g130 ( 
.A(n_72),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_41),
.Y(n_73)
);

INVx3_ASAP7_75t_L g160 ( 
.A(n_73),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_25),
.B(n_9),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_74),
.B(n_80),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_41),
.Y(n_75)
);

INVx3_ASAP7_75t_L g163 ( 
.A(n_75),
.Y(n_163)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_51),
.Y(n_76)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_76),
.Y(n_109)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_34),
.Y(n_77)
);

INVx4_ASAP7_75t_L g148 ( 
.A(n_77),
.Y(n_148)
);

INVx8_ASAP7_75t_L g78 ( 
.A(n_39),
.Y(n_78)
);

INVx4_ASAP7_75t_L g149 ( 
.A(n_78),
.Y(n_149)
);

BUFx5_ASAP7_75t_L g79 ( 
.A(n_35),
.Y(n_79)
);

INVx4_ASAP7_75t_L g152 ( 
.A(n_79),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_25),
.B(n_10),
.Y(n_80)
);

BUFx12f_ASAP7_75t_L g81 ( 
.A(n_28),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_81),
.B(n_83),
.Y(n_127)
);

INVx13_ASAP7_75t_L g82 ( 
.A(n_20),
.Y(n_82)
);

BUFx12f_ASAP7_75t_L g120 ( 
.A(n_82),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_22),
.B(n_8),
.Y(n_83)
);

BUFx12_ASAP7_75t_L g84 ( 
.A(n_20),
.Y(n_84)
);

CKINVDCx16_ASAP7_75t_R g144 ( 
.A(n_84),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_22),
.B(n_37),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_85),
.B(n_87),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_41),
.Y(n_86)
);

INVx4_ASAP7_75t_L g153 ( 
.A(n_86),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_27),
.B(n_8),
.Y(n_87)
);

BUFx3_ASAP7_75t_L g88 ( 
.A(n_34),
.Y(n_88)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_88),
.Y(n_121)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_47),
.Y(n_89)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_89),
.Y(n_129)
);

HB1xp67_ASAP7_75t_L g90 ( 
.A(n_23),
.Y(n_90)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_90),
.Y(n_131)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_34),
.Y(n_91)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_91),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_27),
.B(n_11),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_92),
.B(n_97),
.Y(n_139)
);

BUFx5_ASAP7_75t_L g93 ( 
.A(n_35),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_93),
.B(n_94),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_33),
.B(n_11),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_48),
.Y(n_95)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_95),
.Y(n_134)
);

INVx8_ASAP7_75t_L g96 ( 
.A(n_48),
.Y(n_96)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_96),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_33),
.B(n_7),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_48),
.Y(n_98)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_98),
.Y(n_143)
);

INVx8_ASAP7_75t_L g99 ( 
.A(n_48),
.Y(n_99)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_99),
.Y(n_147)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_35),
.Y(n_100)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_100),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_37),
.B(n_12),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_101),
.B(n_44),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_50),
.Y(n_102)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_102),
.Y(n_156)
);

BUFx12_ASAP7_75t_L g103 ( 
.A(n_28),
.Y(n_103)
);

BUFx12f_ASAP7_75t_L g126 ( 
.A(n_103),
.Y(n_126)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_47),
.Y(n_104)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_104),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_107),
.B(n_38),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_96),
.A2(n_42),
.B1(n_35),
.B2(n_46),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_110),
.A2(n_157),
.B1(n_29),
.B2(n_69),
.Y(n_214)
);

AOI22xp33_ASAP7_75t_L g111 ( 
.A1(n_55),
.A2(n_31),
.B1(n_50),
.B2(n_46),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_111),
.A2(n_145),
.B1(n_154),
.B2(n_46),
.Y(n_182)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_90),
.Y(n_112)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_112),
.Y(n_183)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_58),
.Y(n_114)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_114),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_77),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_124),
.B(n_103),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_53),
.A2(n_44),
.B1(n_31),
.B2(n_50),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_138),
.A2(n_165),
.B1(n_29),
.B2(n_24),
.Y(n_210)
);

OA22x2_ASAP7_75t_L g142 ( 
.A1(n_64),
.A2(n_31),
.B1(n_49),
.B2(n_36),
.Y(n_142)
);

AO22x1_ASAP7_75t_SL g194 ( 
.A1(n_142),
.A2(n_72),
.B1(n_102),
.B2(n_95),
.Y(n_194)
);

AOI22xp33_ASAP7_75t_L g145 ( 
.A1(n_57),
.A2(n_31),
.B1(n_50),
.B2(n_35),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_L g154 ( 
.A1(n_61),
.A2(n_35),
.B1(n_46),
.B2(n_45),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_60),
.Y(n_155)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_155),
.Y(n_199)
);

AOI22xp33_ASAP7_75t_SL g157 ( 
.A1(n_99),
.A2(n_42),
.B1(n_46),
.B2(n_45),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_78),
.A2(n_38),
.B1(n_21),
.B2(n_45),
.Y(n_158)
);

AND2x2_ASAP7_75t_L g207 ( 
.A(n_158),
.B(n_43),
.Y(n_207)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_88),
.Y(n_162)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_162),
.Y(n_167)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_63),
.Y(n_164)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_164),
.Y(n_172)
);

OAI22xp33_ASAP7_75t_SL g165 ( 
.A1(n_65),
.A2(n_49),
.B1(n_24),
.B2(n_43),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g168 ( 
.A(n_105),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g274 ( 
.A(n_168),
.Y(n_274)
);

INVx6_ASAP7_75t_L g169 ( 
.A(n_105),
.Y(n_169)
);

INVx6_ASAP7_75t_L g244 ( 
.A(n_169),
.Y(n_244)
);

AND2x2_ASAP7_75t_SL g170 ( 
.A(n_139),
.B(n_135),
.Y(n_170)
);

AND2x2_ASAP7_75t_L g243 ( 
.A(n_170),
.B(n_177),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_171),
.B(n_175),
.Y(n_228)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_115),
.Y(n_173)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_173),
.Y(n_242)
);

INVx3_ASAP7_75t_L g174 ( 
.A(n_151),
.Y(n_174)
);

INVx3_ASAP7_75t_L g227 ( 
.A(n_174),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_161),
.B(n_21),
.Y(n_175)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_119),
.Y(n_176)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_176),
.Y(n_261)
);

AOI22x1_ASAP7_75t_L g177 ( 
.A1(n_135),
.A2(n_62),
.B1(n_76),
.B2(n_98),
.Y(n_177)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_129),
.Y(n_178)
);

INVx3_ASAP7_75t_L g247 ( 
.A(n_178),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_161),
.B(n_36),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_179),
.B(n_185),
.Y(n_237)
);

INVx3_ASAP7_75t_L g180 ( 
.A(n_151),
.Y(n_180)
);

INVx6_ASAP7_75t_L g250 ( 
.A(n_180),
.Y(n_250)
);

BUFx6f_ASAP7_75t_L g181 ( 
.A(n_125),
.Y(n_181)
);

INVx11_ASAP7_75t_L g262 ( 
.A(n_181),
.Y(n_262)
);

AND2x2_ASAP7_75t_L g253 ( 
.A(n_182),
.B(n_207),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_184),
.B(n_202),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_118),
.B(n_127),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_118),
.B(n_127),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_186),
.B(n_213),
.Y(n_231)
);

AOI21xp33_ASAP7_75t_L g187 ( 
.A1(n_166),
.A2(n_36),
.B(n_49),
.Y(n_187)
);

OR2x2_ASAP7_75t_L g235 ( 
.A(n_187),
.B(n_211),
.Y(n_235)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_159),
.Y(n_189)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_189),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_166),
.B(n_144),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_SL g275 ( 
.A(n_190),
.B(n_200),
.Y(n_275)
);

BUFx6f_ASAP7_75t_L g191 ( 
.A(n_125),
.Y(n_191)
);

CKINVDCx6p67_ASAP7_75t_R g265 ( 
.A(n_191),
.Y(n_265)
);

INVx8_ASAP7_75t_L g192 ( 
.A(n_132),
.Y(n_192)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_192),
.Y(n_239)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_150),
.Y(n_193)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_193),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_194),
.A2(n_205),
.B1(n_215),
.B2(n_221),
.Y(n_259)
);

BUFx10_ASAP7_75t_L g195 ( 
.A(n_126),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_195),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_145),
.A2(n_67),
.B1(n_86),
.B2(n_75),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_196),
.A2(n_146),
.B1(n_123),
.B2(n_141),
.Y(n_230)
);

AOI22xp33_ASAP7_75t_SL g197 ( 
.A1(n_128),
.A2(n_81),
.B1(n_46),
.B2(n_73),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g229 ( 
.A1(n_197),
.A2(n_210),
.B1(n_157),
.B2(n_207),
.Y(n_229)
);

INVx4_ASAP7_75t_L g198 ( 
.A(n_121),
.Y(n_198)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_198),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_120),
.B(n_84),
.Y(n_200)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_131),
.Y(n_201)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_201),
.Y(n_246)
);

CKINVDCx16_ASAP7_75t_R g202 ( 
.A(n_142),
.Y(n_202)
);

BUFx8_ASAP7_75t_L g203 ( 
.A(n_126),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_203),
.Y(n_260)
);

INVx4_ASAP7_75t_SL g204 ( 
.A(n_152),
.Y(n_204)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_204),
.Y(n_248)
);

AOI22xp33_ASAP7_75t_L g205 ( 
.A1(n_117),
.A2(n_43),
.B1(n_29),
.B2(n_24),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_133),
.Y(n_206)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_206),
.Y(n_255)
);

BUFx6f_ASAP7_75t_L g208 ( 
.A(n_132),
.Y(n_208)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_208),
.Y(n_267)
);

INVx3_ASAP7_75t_L g209 ( 
.A(n_120),
.Y(n_209)
);

INVxp67_ASAP7_75t_L g270 ( 
.A(n_209),
.Y(n_270)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_136),
.Y(n_211)
);

INVx6_ASAP7_75t_L g212 ( 
.A(n_137),
.Y(n_212)
);

AOI22xp33_ASAP7_75t_SL g256 ( 
.A1(n_212),
.A2(n_217),
.B1(n_218),
.B2(n_219),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_165),
.B(n_142),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_214),
.A2(n_143),
.B1(n_140),
.B2(n_116),
.Y(n_249)
);

AOI22xp33_ASAP7_75t_L g215 ( 
.A1(n_117),
.A2(n_81),
.B1(n_30),
.B2(n_28),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_106),
.B(n_15),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_216),
.B(n_226),
.Y(n_233)
);

INVx3_ASAP7_75t_L g217 ( 
.A(n_149),
.Y(n_217)
);

INVx4_ASAP7_75t_SL g218 ( 
.A(n_122),
.Y(n_218)
);

BUFx6f_ASAP7_75t_L g219 ( 
.A(n_137),
.Y(n_219)
);

OAI21xp33_ASAP7_75t_SL g220 ( 
.A1(n_110),
.A2(n_103),
.B(n_84),
.Y(n_220)
);

AOI32xp33_ASAP7_75t_L g236 ( 
.A1(n_220),
.A2(n_153),
.A3(n_109),
.B1(n_163),
.B2(n_160),
.Y(n_236)
);

AOI22xp33_ASAP7_75t_L g221 ( 
.A1(n_134),
.A2(n_30),
.B1(n_28),
.B2(n_82),
.Y(n_221)
);

INVx5_ASAP7_75t_L g222 ( 
.A(n_130),
.Y(n_222)
);

AOI22xp33_ASAP7_75t_SL g263 ( 
.A1(n_222),
.A2(n_223),
.B1(n_224),
.B2(n_225),
.Y(n_263)
);

HB1xp67_ASAP7_75t_L g223 ( 
.A(n_113),
.Y(n_223)
);

INVx3_ASAP7_75t_L g224 ( 
.A(n_147),
.Y(n_224)
);

INVx4_ASAP7_75t_L g225 ( 
.A(n_148),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_108),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_229),
.A2(n_238),
.B1(n_258),
.B2(n_264),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_L g279 ( 
.A1(n_230),
.A2(n_212),
.B1(n_208),
.B2(n_219),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_170),
.B(n_194),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_234),
.B(n_252),
.Y(n_284)
);

NAND2x1_ASAP7_75t_L g309 ( 
.A(n_236),
.B(n_17),
.Y(n_309)
);

OAI22xp33_ASAP7_75t_SL g238 ( 
.A1(n_177),
.A2(n_123),
.B1(n_141),
.B2(n_156),
.Y(n_238)
);

OA22x2_ASAP7_75t_L g302 ( 
.A1(n_249),
.A2(n_251),
.B1(n_254),
.B2(n_230),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_220),
.A2(n_146),
.B1(n_111),
.B2(n_154),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_251),
.A2(n_271),
.B1(n_168),
.B2(n_191),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_183),
.B(n_0),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_197),
.A2(n_30),
.B1(n_2),
.B2(n_3),
.Y(n_254)
);

INVxp67_ASAP7_75t_L g288 ( 
.A(n_254),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_188),
.B(n_0),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_257),
.B(n_272),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_L g258 ( 
.A1(n_169),
.A2(n_30),
.B1(n_3),
.B2(n_4),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_205),
.A2(n_0),
.B1(n_3),
.B2(n_4),
.Y(n_264)
);

AOI21xp5_ASAP7_75t_SL g266 ( 
.A1(n_199),
.A2(n_14),
.B(n_4),
.Y(n_266)
);

INVxp67_ASAP7_75t_L g289 ( 
.A(n_266),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_215),
.A2(n_0),
.B1(n_4),
.B2(n_5),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_268),
.A2(n_14),
.B1(n_17),
.B2(n_18),
.Y(n_308)
);

OAI21xp5_ASAP7_75t_SL g269 ( 
.A1(n_221),
.A2(n_14),
.B(n_5),
.Y(n_269)
);

AOI21xp5_ASAP7_75t_L g293 ( 
.A1(n_269),
.A2(n_6),
.B(n_12),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_172),
.A2(n_18),
.B1(n_5),
.B2(n_6),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_167),
.B(n_0),
.Y(n_272)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_255),
.Y(n_277)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_277),
.Y(n_324)
);

INVx3_ASAP7_75t_L g278 ( 
.A(n_250),
.Y(n_278)
);

INVx4_ASAP7_75t_L g330 ( 
.A(n_278),
.Y(n_330)
);

AOI22xp5_ASAP7_75t_L g356 ( 
.A1(n_279),
.A2(n_299),
.B1(n_267),
.B2(n_239),
.Y(n_356)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_265),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_280),
.B(n_283),
.Y(n_321)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_231),
.B(n_198),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_SL g325 ( 
.A(n_281),
.B(n_285),
.Y(n_325)
);

BUFx6f_ASAP7_75t_L g282 ( 
.A(n_274),
.Y(n_282)
);

INVx4_ASAP7_75t_L g343 ( 
.A(n_282),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_SL g283 ( 
.A(n_231),
.B(n_228),
.Y(n_283)
);

MAJx2_ASAP7_75t_L g285 ( 
.A(n_243),
.B(n_218),
.C(n_204),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_233),
.B(n_224),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_287),
.B(n_294),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_SL g290 ( 
.A(n_237),
.B(n_209),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_290),
.B(n_295),
.Y(n_336)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_255),
.Y(n_291)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_291),
.Y(n_359)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_232),
.Y(n_292)
);

INVx1_ASAP7_75t_SL g333 ( 
.A(n_292),
.Y(n_333)
);

OAI21xp5_ASAP7_75t_SL g348 ( 
.A1(n_293),
.A2(n_318),
.B(n_289),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_233),
.B(n_225),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_275),
.B(n_203),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_234),
.B(n_180),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_296),
.B(n_298),
.Y(n_342)
);

NOR2xp67_ASAP7_75t_SL g297 ( 
.A(n_273),
.B(n_195),
.Y(n_297)
);

INVxp67_ASAP7_75t_L g322 ( 
.A(n_297),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_252),
.B(n_192),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g300 ( 
.A(n_235),
.B(n_222),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g347 ( 
.A(n_300),
.B(n_301),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_241),
.B(n_203),
.Y(n_301)
);

AND2x2_ASAP7_75t_L g328 ( 
.A(n_302),
.B(n_308),
.Y(n_328)
);

INVx3_ASAP7_75t_L g303 ( 
.A(n_250),
.Y(n_303)
);

INVx8_ASAP7_75t_L g360 ( 
.A(n_303),
.Y(n_360)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_232),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_304),
.B(n_305),
.Y(n_351)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_246),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_257),
.B(n_181),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_306),
.B(n_311),
.Y(n_355)
);

O2A1O1Ixp33_ASAP7_75t_L g307 ( 
.A1(n_269),
.A2(n_195),
.B(n_15),
.C(n_16),
.Y(n_307)
);

OAI21xp5_ASAP7_75t_L g326 ( 
.A1(n_307),
.A2(n_271),
.B(n_248),
.Y(n_326)
);

AND2x2_ASAP7_75t_L g337 ( 
.A(n_309),
.B(n_316),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_265),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_310),
.Y(n_323)
);

INVxp67_ASAP7_75t_L g311 ( 
.A(n_260),
.Y(n_311)
);

INVx2_ASAP7_75t_L g312 ( 
.A(n_242),
.Y(n_312)
);

INVx3_ASAP7_75t_L g345 ( 
.A(n_312),
.Y(n_345)
);

AOI22xp33_ASAP7_75t_SL g313 ( 
.A1(n_265),
.A2(n_17),
.B1(n_18),
.B2(n_248),
.Y(n_313)
);

INVxp67_ASAP7_75t_L g346 ( 
.A(n_313),
.Y(n_346)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_243),
.B(n_18),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_SL g339 ( 
.A(n_314),
.B(n_264),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_272),
.B(n_235),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_315),
.B(n_259),
.Y(n_358)
);

OA21x2_ASAP7_75t_L g316 ( 
.A1(n_243),
.A2(n_253),
.B(n_249),
.Y(n_316)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_242),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_317),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_R g318 ( 
.A(n_253),
.B(n_266),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_246),
.Y(n_319)
);

AND2x2_ASAP7_75t_L g341 ( 
.A(n_319),
.B(n_245),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_265),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_320),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_326),
.B(n_358),
.Y(n_370)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_296),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g369 ( 
.A(n_331),
.B(n_332),
.Y(n_369)
);

CKINVDCx20_ASAP7_75t_R g332 ( 
.A(n_312),
.Y(n_332)
);

AOI21xp5_ASAP7_75t_SL g334 ( 
.A1(n_318),
.A2(n_253),
.B(n_263),
.Y(n_334)
);

OAI21xp5_ASAP7_75t_L g365 ( 
.A1(n_334),
.A2(n_354),
.B(n_316),
.Y(n_365)
);

BUFx24_ASAP7_75t_SL g335 ( 
.A(n_315),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g364 ( 
.A(n_335),
.B(n_350),
.Y(n_364)
);

XNOR2xp5_ASAP7_75t_L g361 ( 
.A(n_339),
.B(n_349),
.Y(n_361)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_317),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g371 ( 
.A(n_340),
.B(n_344),
.Y(n_371)
);

CKINVDCx16_ASAP7_75t_R g390 ( 
.A(n_341),
.Y(n_390)
);

CKINVDCx20_ASAP7_75t_R g344 ( 
.A(n_287),
.Y(n_344)
);

AOI21xp5_ASAP7_75t_L g386 ( 
.A1(n_348),
.A2(n_354),
.B(n_337),
.Y(n_386)
);

XNOR2xp5_ASAP7_75t_SL g349 ( 
.A(n_281),
.B(n_259),
.Y(n_349)
);

INVxp67_ASAP7_75t_L g350 ( 
.A(n_307),
.Y(n_350)
);

INVxp67_ASAP7_75t_L g352 ( 
.A(n_294),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_L g375 ( 
.A(n_352),
.B(n_353),
.Y(n_375)
);

INVxp67_ASAP7_75t_L g353 ( 
.A(n_293),
.Y(n_353)
);

OAI21xp5_ASAP7_75t_L g354 ( 
.A1(n_289),
.A2(n_241),
.B(n_260),
.Y(n_354)
);

OAI22xp5_ASAP7_75t_SL g373 ( 
.A1(n_356),
.A2(n_357),
.B1(n_276),
.B2(n_358),
.Y(n_373)
);

AOI22xp5_ASAP7_75t_L g357 ( 
.A1(n_299),
.A2(n_288),
.B1(n_276),
.B2(n_302),
.Y(n_357)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_351),
.Y(n_362)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_362),
.Y(n_397)
);

AOI22xp5_ASAP7_75t_L g363 ( 
.A1(n_328),
.A2(n_288),
.B1(n_302),
.B2(n_309),
.Y(n_363)
);

OAI22xp5_ASAP7_75t_SL g399 ( 
.A1(n_363),
.A2(n_383),
.B1(n_395),
.B2(n_346),
.Y(n_399)
);

OAI21xp5_ASAP7_75t_L g408 ( 
.A1(n_365),
.A2(n_367),
.B(n_394),
.Y(n_408)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_351),
.Y(n_366)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_366),
.Y(n_398)
);

OAI21xp5_ASAP7_75t_L g367 ( 
.A1(n_334),
.A2(n_316),
.B(n_284),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_324),
.Y(n_368)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_368),
.Y(n_409)
);

MAJIxp5_ASAP7_75t_L g372 ( 
.A(n_325),
.B(n_285),
.C(n_284),
.Y(n_372)
);

MAJIxp5_ASAP7_75t_L g410 ( 
.A(n_372),
.B(n_382),
.C(n_348),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_373),
.B(n_374),
.Y(n_403)
);

OAI22xp5_ASAP7_75t_L g374 ( 
.A1(n_357),
.A2(n_302),
.B1(n_298),
.B2(n_309),
.Y(n_374)
);

CKINVDCx20_ASAP7_75t_R g376 ( 
.A(n_341),
.Y(n_376)
);

CKINVDCx20_ASAP7_75t_R g407 ( 
.A(n_376),
.Y(n_407)
);

OAI22xp5_ASAP7_75t_L g377 ( 
.A1(n_331),
.A2(n_306),
.B1(n_308),
.B2(n_286),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_377),
.B(n_378),
.Y(n_406)
);

OAI22xp5_ASAP7_75t_SL g378 ( 
.A1(n_344),
.A2(n_286),
.B1(n_311),
.B2(n_256),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_324),
.Y(n_379)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_379),
.Y(n_411)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_359),
.Y(n_380)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_380),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_338),
.B(n_277),
.Y(n_381)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_381),
.Y(n_419)
);

MAJIxp5_ASAP7_75t_L g382 ( 
.A(n_325),
.B(n_349),
.C(n_342),
.Y(n_382)
);

AOI22xp5_ASAP7_75t_L g383 ( 
.A1(n_328),
.A2(n_314),
.B1(n_268),
.B2(n_303),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_338),
.B(n_319),
.Y(n_384)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_384),
.Y(n_421)
);

NOR2xp33_ASAP7_75t_SL g385 ( 
.A(n_336),
.B(n_347),
.Y(n_385)
);

NAND3xp33_ASAP7_75t_L g422 ( 
.A(n_385),
.B(n_327),
.C(n_340),
.Y(n_422)
);

OAI21xp5_ASAP7_75t_SL g423 ( 
.A1(n_386),
.A2(n_330),
.B(n_345),
.Y(n_423)
);

AOI22xp5_ASAP7_75t_SL g387 ( 
.A1(n_328),
.A2(n_278),
.B1(n_292),
.B2(n_304),
.Y(n_387)
);

AOI21xp5_ASAP7_75t_L g404 ( 
.A1(n_387),
.A2(n_326),
.B(n_322),
.Y(n_404)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_359),
.Y(n_388)
);

INVxp67_ASAP7_75t_L g401 ( 
.A(n_388),
.Y(n_401)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_355),
.Y(n_389)
);

NOR2xp33_ASAP7_75t_L g413 ( 
.A(n_389),
.B(n_355),
.Y(n_413)
);

OAI22xp5_ASAP7_75t_L g391 ( 
.A1(n_356),
.A2(n_267),
.B1(n_282),
.B2(n_239),
.Y(n_391)
);

OAI22xp5_ASAP7_75t_L g396 ( 
.A1(n_391),
.A2(n_376),
.B1(n_393),
.B2(n_389),
.Y(n_396)
);

XNOR2xp5_ASAP7_75t_L g392 ( 
.A(n_342),
.B(n_240),
.Y(n_392)
);

XNOR2xp5_ASAP7_75t_L g402 ( 
.A(n_392),
.B(n_339),
.Y(n_402)
);

CKINVDCx20_ASAP7_75t_R g393 ( 
.A(n_341),
.Y(n_393)
);

CKINVDCx20_ASAP7_75t_R g425 ( 
.A(n_393),
.Y(n_425)
);

OAI21xp5_ASAP7_75t_L g394 ( 
.A1(n_334),
.A2(n_245),
.B(n_240),
.Y(n_394)
);

AOI22xp5_ASAP7_75t_L g395 ( 
.A1(n_337),
.A2(n_244),
.B1(n_274),
.B2(n_227),
.Y(n_395)
);

AOI22xp5_ASAP7_75t_L g438 ( 
.A1(n_396),
.A2(n_414),
.B1(n_390),
.B2(n_374),
.Y(n_438)
);

AOI22xp5_ASAP7_75t_SL g451 ( 
.A1(n_399),
.A2(n_378),
.B1(n_391),
.B2(n_377),
.Y(n_451)
);

XOR2xp5_ASAP7_75t_L g400 ( 
.A(n_361),
.B(n_337),
.Y(n_400)
);

MAJIxp5_ASAP7_75t_L g435 ( 
.A(n_400),
.B(n_417),
.C(n_418),
.Y(n_435)
);

XNOR2xp5_ASAP7_75t_L g444 ( 
.A(n_402),
.B(n_410),
.Y(n_444)
);

INVxp67_ASAP7_75t_L g441 ( 
.A(n_404),
.Y(n_441)
);

AOI21xp33_ASAP7_75t_L g405 ( 
.A1(n_375),
.A2(n_347),
.B(n_336),
.Y(n_405)
);

NAND3xp33_ASAP7_75t_L g448 ( 
.A(n_405),
.B(n_415),
.C(n_371),
.Y(n_448)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_413),
.Y(n_428)
);

OAI22xp5_ASAP7_75t_SL g414 ( 
.A1(n_363),
.A2(n_321),
.B1(n_333),
.B2(n_323),
.Y(n_414)
);

NOR2xp33_ASAP7_75t_SL g415 ( 
.A(n_364),
.B(n_321),
.Y(n_415)
);

NOR2xp33_ASAP7_75t_L g416 ( 
.A(n_385),
.B(n_329),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_SL g431 ( 
.A(n_416),
.B(n_424),
.Y(n_431)
);

XNOR2xp5_ASAP7_75t_L g417 ( 
.A(n_372),
.B(n_333),
.Y(n_417)
);

XNOR2xp5_ASAP7_75t_L g418 ( 
.A(n_382),
.B(n_333),
.Y(n_418)
);

OAI22x1_ASAP7_75t_L g420 ( 
.A1(n_365),
.A2(n_329),
.B1(n_323),
.B2(n_360),
.Y(n_420)
);

OAI22xp5_ASAP7_75t_L g440 ( 
.A1(n_420),
.A2(n_387),
.B1(n_394),
.B2(n_390),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_L g446 ( 
.A(n_422),
.B(n_426),
.Y(n_446)
);

CKINVDCx20_ASAP7_75t_R g427 ( 
.A(n_423),
.Y(n_427)
);

MAJIxp5_ASAP7_75t_L g424 ( 
.A(n_361),
.B(n_327),
.C(n_332),
.Y(n_424)
);

HB1xp67_ASAP7_75t_L g426 ( 
.A(n_362),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_397),
.B(n_366),
.Y(n_429)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_429),
.Y(n_455)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_397),
.Y(n_430)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_430),
.Y(n_465)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_398),
.Y(n_432)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_432),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_398),
.B(n_381),
.Y(n_433)
);

CKINVDCx20_ASAP7_75t_R g471 ( 
.A(n_433),
.Y(n_471)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_409),
.Y(n_434)
);

NOR2xp33_ASAP7_75t_L g462 ( 
.A(n_434),
.B(n_436),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_SL g436 ( 
.A(n_424),
.B(n_370),
.Y(n_436)
);

OAI22xp5_ASAP7_75t_SL g437 ( 
.A1(n_403),
.A2(n_370),
.B1(n_383),
.B2(n_367),
.Y(n_437)
);

OAI22xp5_ASAP7_75t_L g463 ( 
.A1(n_437),
.A2(n_442),
.B1(n_443),
.B2(n_447),
.Y(n_463)
);

OAI22xp5_ASAP7_75t_SL g453 ( 
.A1(n_438),
.A2(n_451),
.B1(n_406),
.B2(n_420),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_407),
.B(n_384),
.Y(n_439)
);

HB1xp67_ASAP7_75t_L g474 ( 
.A(n_439),
.Y(n_474)
);

OAI21xp5_ASAP7_75t_SL g459 ( 
.A1(n_440),
.A2(n_404),
.B(n_406),
.Y(n_459)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_409),
.Y(n_442)
);

OAI22xp5_ASAP7_75t_SL g443 ( 
.A1(n_403),
.A2(n_369),
.B1(n_371),
.B2(n_373),
.Y(n_443)
);

NOR2xp33_ASAP7_75t_SL g445 ( 
.A(n_425),
.B(n_369),
.Y(n_445)
);

NOR2xp33_ASAP7_75t_SL g470 ( 
.A(n_445),
.B(n_452),
.Y(n_470)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_411),
.Y(n_447)
);

OAI22xp5_ASAP7_75t_L g473 ( 
.A1(n_448),
.A2(n_449),
.B1(n_450),
.B2(n_388),
.Y(n_473)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_411),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_412),
.Y(n_450)
);

NOR2xp33_ASAP7_75t_L g452 ( 
.A(n_414),
.B(n_392),
.Y(n_452)
);

AOI22xp5_ASAP7_75t_L g483 ( 
.A1(n_453),
.A2(n_467),
.B1(n_428),
.B2(n_432),
.Y(n_483)
);

NAND2x1p5_ASAP7_75t_L g454 ( 
.A(n_427),
.B(n_408),
.Y(n_454)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_454),
.Y(n_479)
);

XNOR2xp5_ASAP7_75t_L g456 ( 
.A(n_444),
.B(n_418),
.Y(n_456)
);

XNOR2xp5_ASAP7_75t_L g480 ( 
.A(n_456),
.B(n_439),
.Y(n_480)
);

AOI21xp5_ASAP7_75t_L g457 ( 
.A1(n_441),
.A2(n_408),
.B(n_423),
.Y(n_457)
);

INVxp67_ASAP7_75t_L g485 ( 
.A(n_457),
.Y(n_485)
);

XOR2xp5_ASAP7_75t_L g458 ( 
.A(n_435),
.B(n_400),
.Y(n_458)
);

XNOR2xp5_ASAP7_75t_SL g486 ( 
.A(n_458),
.B(n_459),
.Y(n_486)
);

MAJIxp5_ASAP7_75t_L g460 ( 
.A(n_431),
.B(n_417),
.C(n_410),
.Y(n_460)
);

MAJIxp5_ASAP7_75t_L g477 ( 
.A(n_460),
.B(n_461),
.C(n_469),
.Y(n_477)
);

MAJIxp5_ASAP7_75t_L g461 ( 
.A(n_444),
.B(n_402),
.C(n_399),
.Y(n_461)
);

XOR2xp5_ASAP7_75t_L g464 ( 
.A(n_435),
.B(n_386),
.Y(n_464)
);

XOR2xp5_ASAP7_75t_L g475 ( 
.A(n_464),
.B(n_443),
.Y(n_475)
);

OAI21xp5_ASAP7_75t_L g466 ( 
.A1(n_441),
.A2(n_421),
.B(n_419),
.Y(n_466)
);

AOI21xp5_ASAP7_75t_L g484 ( 
.A1(n_466),
.A2(n_433),
.B(n_428),
.Y(n_484)
);

OAI22xp5_ASAP7_75t_SL g467 ( 
.A1(n_451),
.A2(n_421),
.B1(n_419),
.B2(n_395),
.Y(n_467)
);

MAJIxp5_ASAP7_75t_L g469 ( 
.A(n_438),
.B(n_401),
.C(n_412),
.Y(n_469)
);

MAJIxp5_ASAP7_75t_L g472 ( 
.A(n_437),
.B(n_401),
.C(n_368),
.Y(n_472)
);

MAJIxp5_ASAP7_75t_L g482 ( 
.A(n_472),
.B(n_427),
.C(n_430),
.Y(n_482)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_473),
.Y(n_481)
);

XOR2xp5_ASAP7_75t_L g502 ( 
.A(n_475),
.B(n_480),
.Y(n_502)
);

XNOR2xp5_ASAP7_75t_L g476 ( 
.A(n_456),
.B(n_446),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_SL g503 ( 
.A(n_476),
.B(n_478),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_470),
.B(n_429),
.Y(n_478)
);

XNOR2xp5_ASAP7_75t_L g497 ( 
.A(n_482),
.B(n_483),
.Y(n_497)
);

XNOR2xp5_ASAP7_75t_L g498 ( 
.A(n_484),
.B(n_488),
.Y(n_498)
);

OAI21xp5_ASAP7_75t_SL g487 ( 
.A1(n_457),
.A2(n_450),
.B(n_449),
.Y(n_487)
);

AOI21xp5_ASAP7_75t_L g492 ( 
.A1(n_487),
.A2(n_466),
.B(n_459),
.Y(n_492)
);

XOR2xp5_ASAP7_75t_L g488 ( 
.A(n_464),
.B(n_447),
.Y(n_488)
);

MAJIxp5_ASAP7_75t_L g489 ( 
.A(n_460),
.B(n_442),
.C(n_434),
.Y(n_489)
);

MAJIxp5_ASAP7_75t_L g499 ( 
.A(n_489),
.B(n_491),
.C(n_468),
.Y(n_499)
);

XNOR2xp5_ASAP7_75t_L g490 ( 
.A(n_461),
.B(n_379),
.Y(n_490)
);

HB1xp67_ASAP7_75t_L g505 ( 
.A(n_490),
.Y(n_505)
);

MAJIxp5_ASAP7_75t_L g491 ( 
.A(n_472),
.B(n_380),
.C(n_330),
.Y(n_491)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_492),
.Y(n_514)
);

AOI22xp5_ASAP7_75t_L g493 ( 
.A1(n_481),
.A2(n_463),
.B1(n_467),
.B2(n_453),
.Y(n_493)
);

OAI22xp5_ASAP7_75t_SL g515 ( 
.A1(n_493),
.A2(n_500),
.B1(n_504),
.B2(n_343),
.Y(n_515)
);

FAx1_ASAP7_75t_SL g494 ( 
.A(n_480),
.B(n_469),
.CI(n_454),
.CON(n_494),
.SN(n_494)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_494),
.Y(n_516)
);

FAx1_ASAP7_75t_SL g495 ( 
.A(n_486),
.B(n_454),
.CI(n_470),
.CON(n_495),
.SN(n_495)
);

NAND2xp5_ASAP7_75t_SL g508 ( 
.A(n_495),
.B(n_499),
.Y(n_508)
);

AOI22xp5_ASAP7_75t_L g496 ( 
.A1(n_475),
.A2(n_455),
.B1(n_471),
.B2(n_474),
.Y(n_496)
);

OAI22xp5_ASAP7_75t_L g509 ( 
.A1(n_496),
.A2(n_491),
.B1(n_489),
.B2(n_486),
.Y(n_509)
);

AOI22xp5_ASAP7_75t_L g500 ( 
.A1(n_485),
.A2(n_455),
.B1(n_471),
.B2(n_462),
.Y(n_500)
);

MAJIxp5_ASAP7_75t_L g501 ( 
.A(n_477),
.B(n_458),
.C(n_468),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_SL g511 ( 
.A(n_501),
.B(n_330),
.Y(n_511)
);

AOI22xp5_ASAP7_75t_L g504 ( 
.A1(n_485),
.A2(n_479),
.B1(n_488),
.B2(n_465),
.Y(n_504)
);

OAI21x1_ASAP7_75t_SL g506 ( 
.A1(n_482),
.A2(n_465),
.B(n_360),
.Y(n_506)
);

AOI21xp5_ASAP7_75t_L g512 ( 
.A1(n_506),
.A2(n_343),
.B(n_345),
.Y(n_512)
);

XNOR2xp5_ASAP7_75t_L g507 ( 
.A(n_502),
.B(n_477),
.Y(n_507)
);

XNOR2xp5_ASAP7_75t_SL g523 ( 
.A(n_507),
.B(n_510),
.Y(n_523)
);

AOI22xp5_ASAP7_75t_L g518 ( 
.A1(n_509),
.A2(n_512),
.B1(n_515),
.B2(n_498),
.Y(n_518)
);

XOR2xp5_ASAP7_75t_L g510 ( 
.A(n_502),
.B(n_360),
.Y(n_510)
);

AOI21xp5_ASAP7_75t_L g519 ( 
.A1(n_511),
.A2(n_513),
.B(n_517),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_SL g513 ( 
.A(n_501),
.B(n_343),
.Y(n_513)
);

XNOR2xp5_ASAP7_75t_L g517 ( 
.A(n_497),
.B(n_227),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_518),
.B(n_524),
.Y(n_528)
);

AOI21x1_ASAP7_75t_L g520 ( 
.A1(n_508),
.A2(n_495),
.B(n_500),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_SL g525 ( 
.A(n_520),
.B(n_522),
.Y(n_525)
);

MAJx2_ASAP7_75t_L g521 ( 
.A(n_516),
.B(n_499),
.C(n_494),
.Y(n_521)
);

NOR2x1_ASAP7_75t_L g527 ( 
.A(n_521),
.B(n_498),
.Y(n_527)
);

MAJIxp5_ASAP7_75t_L g522 ( 
.A(n_507),
.B(n_503),
.C(n_497),
.Y(n_522)
);

INVx1_ASAP7_75t_SL g524 ( 
.A(n_517),
.Y(n_524)
);

AND2x2_ASAP7_75t_L g526 ( 
.A(n_520),
.B(n_514),
.Y(n_526)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_526),
.Y(n_530)
);

AND2x2_ASAP7_75t_L g531 ( 
.A(n_527),
.B(n_504),
.Y(n_531)
);

OAI21xp5_ASAP7_75t_SL g529 ( 
.A1(n_525),
.A2(n_519),
.B(n_523),
.Y(n_529)
);

MAJIxp5_ASAP7_75t_L g532 ( 
.A(n_529),
.B(n_528),
.C(n_510),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_531),
.B(n_515),
.Y(n_533)
);

AO21x1_ASAP7_75t_L g534 ( 
.A1(n_532),
.A2(n_533),
.B(n_530),
.Y(n_534)
);

AOI22xp5_ASAP7_75t_L g535 ( 
.A1(n_534),
.A2(n_505),
.B1(n_493),
.B2(n_244),
.Y(n_535)
);

A2O1A1Ixp33_ASAP7_75t_L g536 ( 
.A1(n_535),
.A2(n_270),
.B(n_262),
.C(n_247),
.Y(n_536)
);

OAI21xp5_ASAP7_75t_SL g537 ( 
.A1(n_536),
.A2(n_270),
.B(n_247),
.Y(n_537)
);

MAJIxp5_ASAP7_75t_L g538 ( 
.A(n_537),
.B(n_261),
.C(n_262),
.Y(n_538)
);

XOR2xp5_ASAP7_75t_L g539 ( 
.A(n_538),
.B(n_261),
.Y(n_539)
);


endmodule