module fake_jpeg_22745_n_319 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_319);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_319;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_145;
wire n_20;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g15 ( 
.A(n_9),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

BUFx5_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_11),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_14),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_10),
.Y(n_25)
);

BUFx2_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_10),
.Y(n_28)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

BUFx24_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_31),
.Y(n_32)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_32),
.Y(n_55)
);

INVx4_ASAP7_75t_SL g33 ( 
.A(n_31),
.Y(n_33)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_33),
.A2(n_29),
.B1(n_19),
.B2(n_17),
.Y(n_47)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_24),
.B(n_27),
.Y(n_36)
);

OR2x2_ASAP7_75t_L g60 ( 
.A(n_36),
.B(n_39),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_31),
.Y(n_37)
);

BUFx2_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_31),
.Y(n_38)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_38),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_24),
.B(n_14),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_26),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_41),
.B(n_29),
.Y(n_54)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_42),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_39),
.B(n_36),
.Y(n_46)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_46),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_47),
.A2(n_50),
.B1(n_35),
.B2(n_33),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_41),
.B(n_21),
.Y(n_49)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_49),
.Y(n_77)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_41),
.B(n_21),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_53),
.B(n_54),
.Y(n_86)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_34),
.Y(n_56)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_56),
.Y(n_74)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_32),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_57),
.B(n_59),
.Y(n_70)
);

BUFx5_ASAP7_75t_L g58 ( 
.A(n_32),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_58),
.Y(n_75)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_32),
.Y(n_59)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_37),
.Y(n_61)
);

INVx4_ASAP7_75t_SL g80 ( 
.A(n_61),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_37),
.Y(n_62)
);

BUFx2_ASAP7_75t_L g85 ( 
.A(n_62),
.Y(n_85)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_37),
.Y(n_63)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_63),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_40),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_64),
.Y(n_87)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_40),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g88 ( 
.A(n_65),
.Y(n_88)
);

OAI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_43),
.A2(n_35),
.B1(n_34),
.B2(n_29),
.Y(n_66)
);

OAI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_66),
.A2(n_82),
.B1(n_42),
.B2(n_40),
.Y(n_108)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_55),
.Y(n_67)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_67),
.Y(n_96)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_65),
.Y(n_68)
);

INVx6_ASAP7_75t_L g90 ( 
.A(n_68),
.Y(n_90)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_58),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_69),
.B(n_78),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_43),
.A2(n_35),
.B1(n_34),
.B2(n_29),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_72),
.A2(n_44),
.B1(n_84),
.B2(n_79),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_73),
.A2(n_81),
.B1(n_33),
.B2(n_42),
.Y(n_98)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_55),
.Y(n_76)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_76),
.Y(n_107)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_64),
.Y(n_78)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_48),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_79),
.B(n_84),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_45),
.A2(n_19),
.B1(n_24),
.B2(n_27),
.Y(n_81)
);

OAI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_48),
.A2(n_19),
.B1(n_18),
.B2(n_33),
.Y(n_82)
);

BUFx12f_ASAP7_75t_L g83 ( 
.A(n_59),
.Y(n_83)
);

BUFx12_ASAP7_75t_L g100 ( 
.A(n_83),
.Y(n_100)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_56),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_71),
.B(n_60),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_92),
.B(n_106),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_83),
.Y(n_93)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_93),
.Y(n_129)
);

BUFx2_ASAP7_75t_L g94 ( 
.A(n_83),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_94),
.Y(n_118)
);

OAI22xp33_ASAP7_75t_L g97 ( 
.A1(n_72),
.A2(n_76),
.B1(n_67),
.B2(n_78),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_97),
.A2(n_99),
.B1(n_108),
.B2(n_109),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_98),
.A2(n_104),
.B1(n_113),
.B2(n_114),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_86),
.A2(n_45),
.B1(n_33),
.B2(n_42),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_87),
.B(n_60),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_101),
.B(n_103),
.Y(n_119)
);

INVx1_ASAP7_75t_SL g102 ( 
.A(n_75),
.Y(n_102)
);

INVx1_ASAP7_75t_SL g135 ( 
.A(n_102),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_74),
.B(n_22),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_74),
.A2(n_27),
.B1(n_44),
.B2(n_50),
.Y(n_104)
);

CKINVDCx14_ASAP7_75t_R g105 ( 
.A(n_70),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_105),
.B(n_80),
.Y(n_137)
);

CKINVDCx16_ASAP7_75t_R g106 ( 
.A(n_85),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_77),
.B(n_30),
.Y(n_110)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_110),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_77),
.B(n_80),
.Y(n_111)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_111),
.Y(n_126)
);

AND2x2_ASAP7_75t_L g112 ( 
.A(n_75),
.B(n_17),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_112),
.B(n_113),
.C(n_96),
.Y(n_130)
);

BUFx12f_ASAP7_75t_SL g113 ( 
.A(n_88),
.Y(n_113)
);

INVx5_ASAP7_75t_L g114 ( 
.A(n_88),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_101),
.A2(n_63),
.B1(n_51),
.B2(n_57),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_115),
.A2(n_123),
.B1(n_106),
.B2(n_90),
.Y(n_145)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_100),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g155 ( 
.A1(n_120),
.A2(n_121),
.B1(n_132),
.B2(n_134),
.Y(n_155)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_100),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_95),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_122),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_103),
.A2(n_61),
.B1(n_51),
.B2(n_89),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_105),
.B(n_89),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_125),
.B(n_127),
.Y(n_148)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_95),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_91),
.B(n_62),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_128),
.B(n_131),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_130),
.B(n_133),
.C(n_123),
.Y(n_147)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_91),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_94),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_99),
.B(n_52),
.C(n_17),
.Y(n_133)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_100),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_94),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_SL g141 ( 
.A1(n_136),
.A2(n_139),
.B(n_107),
.Y(n_141)
);

INVxp33_ASAP7_75t_L g162 ( 
.A(n_137),
.Y(n_162)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_111),
.Y(n_139)
);

A2O1A1Ixp33_ASAP7_75t_SL g140 ( 
.A1(n_109),
.A2(n_23),
.B(n_18),
.C(n_38),
.Y(n_140)
);

AOI21xp5_ASAP7_75t_L g163 ( 
.A1(n_140),
.A2(n_68),
.B(n_69),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_SL g182 ( 
.A1(n_141),
.A2(n_153),
.B(n_157),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_117),
.A2(n_107),
.B1(n_96),
.B2(n_112),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_142),
.A2(n_156),
.B1(n_158),
.B2(n_140),
.Y(n_168)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_128),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_143),
.B(n_146),
.Y(n_176)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_129),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_144),
.Y(n_167)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_145),
.Y(n_170)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_125),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_147),
.B(n_151),
.C(n_160),
.Y(n_173)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_119),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_149),
.B(n_152),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_129),
.Y(n_150)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_150),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_130),
.B(n_119),
.C(n_133),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_115),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_SL g153 ( 
.A1(n_122),
.A2(n_92),
.B(n_112),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g154 ( 
.A(n_117),
.B(n_110),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g175 ( 
.A(n_154),
.B(n_140),
.Y(n_175)
);

OAI32xp33_ASAP7_75t_L g156 ( 
.A1(n_140),
.A2(n_18),
.A3(n_23),
.B1(n_15),
.B2(n_30),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_116),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_138),
.A2(n_90),
.B1(n_23),
.B2(n_15),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_131),
.B(n_102),
.C(n_90),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_SL g189 ( 
.A1(n_163),
.A2(n_165),
.B(n_166),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_L g164 ( 
.A1(n_127),
.A2(n_126),
.B(n_139),
.Y(n_164)
);

AOI21xp5_ASAP7_75t_L g179 ( 
.A1(n_164),
.A2(n_20),
.B(n_28),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_126),
.A2(n_28),
.B1(n_25),
.B2(n_20),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_SL g166 ( 
.A1(n_124),
.A2(n_15),
.B(n_30),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_SL g211 ( 
.A1(n_168),
.A2(n_179),
.B(n_183),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_159),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_169),
.Y(n_196)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_148),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_171),
.B(n_178),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_152),
.A2(n_140),
.B1(n_124),
.B2(n_118),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_174),
.A2(n_177),
.B1(n_180),
.B2(n_192),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_175),
.B(n_173),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_163),
.A2(n_136),
.B1(n_132),
.B2(n_118),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_148),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_149),
.A2(n_145),
.B1(n_147),
.B2(n_153),
.Y(n_180)
);

OR2x2_ASAP7_75t_L g181 ( 
.A(n_159),
.B(n_20),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_181),
.B(n_166),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_157),
.A2(n_134),
.B1(n_121),
.B2(n_120),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_161),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_184),
.B(n_187),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_151),
.B(n_135),
.C(n_114),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_185),
.B(n_144),
.C(n_150),
.Y(n_206)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_161),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_156),
.A2(n_142),
.B1(n_146),
.B2(n_143),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_188),
.B(n_190),
.Y(n_210)
);

INVxp67_ASAP7_75t_L g190 ( 
.A(n_155),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_SL g191 ( 
.A1(n_141),
.A2(n_135),
.B(n_52),
.Y(n_191)
);

AOI21xp5_ASAP7_75t_L g199 ( 
.A1(n_191),
.A2(n_164),
.B(n_160),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_154),
.A2(n_62),
.B1(n_25),
.B2(n_85),
.Y(n_192)
);

CKINVDCx16_ASAP7_75t_R g193 ( 
.A(n_186),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_193),
.B(n_195),
.Y(n_219)
);

INVx3_ASAP7_75t_L g195 ( 
.A(n_177),
.Y(n_195)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_176),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_197),
.B(n_203),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_198),
.B(n_189),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_SL g231 ( 
.A1(n_199),
.A2(n_189),
.B(n_192),
.Y(n_231)
);

XOR2x2_ASAP7_75t_L g200 ( 
.A(n_175),
.B(n_162),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_SL g234 ( 
.A(n_200),
.B(n_201),
.Y(n_234)
);

FAx1_ASAP7_75t_SL g203 ( 
.A(n_180),
.B(n_165),
.CI(n_38),
.CON(n_203),
.SN(n_203)
);

BUFx6f_ASAP7_75t_L g204 ( 
.A(n_172),
.Y(n_204)
);

INVx13_ASAP7_75t_L g217 ( 
.A(n_204),
.Y(n_217)
);

HB1xp67_ASAP7_75t_L g205 ( 
.A(n_167),
.Y(n_205)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_205),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_206),
.B(n_208),
.C(n_216),
.Y(n_223)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_176),
.Y(n_207)
);

AOI22xp33_ASAP7_75t_L g222 ( 
.A1(n_207),
.A2(n_171),
.B1(n_191),
.B2(n_169),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_173),
.B(n_100),
.C(n_93),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_SL g212 ( 
.A(n_168),
.B(n_26),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_212),
.B(n_181),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_170),
.A2(n_93),
.B1(n_22),
.B2(n_16),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_213),
.A2(n_214),
.B1(n_215),
.B2(n_183),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_186),
.A2(n_22),
.B1(n_16),
.B2(n_52),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_174),
.A2(n_184),
.B1(n_187),
.B2(n_178),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_185),
.B(n_26),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_196),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_220),
.Y(n_247)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_222),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_224),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_225),
.A2(n_232),
.B1(n_237),
.B2(n_212),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_198),
.B(n_182),
.Y(n_226)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_226),
.Y(n_244)
);

AOI22xp33_ASAP7_75t_L g227 ( 
.A1(n_199),
.A2(n_167),
.B1(n_182),
.B2(n_179),
.Y(n_227)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_227),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_194),
.Y(n_228)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_228),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_202),
.Y(n_229)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_229),
.Y(n_249)
);

INVxp67_ASAP7_75t_L g230 ( 
.A(n_206),
.Y(n_230)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_230),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_231),
.B(n_211),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_L g232 ( 
.A1(n_195),
.A2(n_215),
.B1(n_209),
.B2(n_210),
.Y(n_232)
);

AOI21xp5_ASAP7_75t_L g233 ( 
.A1(n_211),
.A2(n_188),
.B(n_181),
.Y(n_233)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_233),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_235),
.B(n_26),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_208),
.B(n_201),
.C(n_216),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_236),
.B(n_223),
.C(n_234),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_200),
.A2(n_22),
.B1(n_1),
.B2(n_2),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_240),
.B(n_248),
.C(n_251),
.Y(n_261)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_241),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_L g267 ( 
.A1(n_242),
.A2(n_237),
.B1(n_231),
.B2(n_232),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_SL g243 ( 
.A(n_234),
.B(n_209),
.Y(n_243)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_243),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_223),
.B(n_214),
.C(n_203),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_236),
.B(n_203),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_228),
.B(n_213),
.C(n_204),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_252),
.B(n_255),
.C(n_256),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g257 ( 
.A(n_253),
.B(n_235),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_226),
.B(n_13),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_229),
.B(n_0),
.C(n_1),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_257),
.B(n_258),
.Y(n_277)
);

CKINVDCx16_ASAP7_75t_R g258 ( 
.A(n_252),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_247),
.B(n_220),
.Y(n_260)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_260),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_254),
.A2(n_219),
.B1(n_224),
.B2(n_230),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_262),
.B(n_243),
.Y(n_278)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_256),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_263),
.B(n_271),
.C(n_272),
.Y(n_285)
);

OAI21xp5_ASAP7_75t_SL g265 ( 
.A1(n_244),
.A2(n_233),
.B(n_221),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_265),
.B(n_266),
.C(n_246),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_255),
.B(n_225),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_267),
.A2(n_263),
.B1(n_270),
.B2(n_259),
.Y(n_279)
);

CKINVDCx14_ASAP7_75t_R g268 ( 
.A(n_248),
.Y(n_268)
);

AOI22xp33_ASAP7_75t_L g283 ( 
.A1(n_268),
.A2(n_218),
.B1(n_14),
.B2(n_13),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_239),
.B(n_217),
.Y(n_269)
);

INVxp67_ASAP7_75t_L g273 ( 
.A(n_269),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_250),
.B(n_240),
.C(n_249),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_241),
.Y(n_272)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_274),
.Y(n_286)
);

OAI21xp5_ASAP7_75t_L g276 ( 
.A1(n_271),
.A2(n_245),
.B(n_238),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_276),
.B(n_284),
.Y(n_289)
);

XOR2xp5_ASAP7_75t_L g291 ( 
.A(n_278),
.B(n_280),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_L g293 ( 
.A1(n_279),
.A2(n_281),
.B1(n_283),
.B2(n_0),
.Y(n_293)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_261),
.B(n_251),
.Y(n_280)
);

AOI21xp33_ASAP7_75t_L g281 ( 
.A1(n_259),
.A2(n_218),
.B(n_217),
.Y(n_281)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_261),
.B(n_253),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g295 ( 
.A(n_282),
.B(n_2),
.Y(n_295)
);

NOR3xp33_ASAP7_75t_SL g284 ( 
.A(n_265),
.B(n_12),
.C(n_1),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_280),
.B(n_264),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_287),
.B(n_292),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_284),
.B(n_262),
.Y(n_288)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_288),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_273),
.A2(n_264),
.B1(n_272),
.B2(n_12),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_290),
.B(n_295),
.C(n_278),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_282),
.B(n_0),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_293),
.B(n_294),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_275),
.B(n_0),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_285),
.B(n_2),
.Y(n_296)
);

OR2x2_ASAP7_75t_SL g297 ( 
.A(n_296),
.B(n_273),
.Y(n_297)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_297),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_299),
.B(n_291),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_296),
.B(n_277),
.Y(n_300)
);

OR2x2_ASAP7_75t_L g307 ( 
.A(n_300),
.B(n_295),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_286),
.B(n_285),
.Y(n_301)
);

AOI21xp5_ASAP7_75t_L g305 ( 
.A1(n_301),
.A2(n_304),
.B(n_289),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_291),
.B(n_3),
.C(n_4),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_305),
.B(n_307),
.C(n_308),
.Y(n_311)
);

NOR2xp67_ASAP7_75t_SL g309 ( 
.A(n_303),
.B(n_3),
.Y(n_309)
);

AOI21xp5_ASAP7_75t_SL g312 ( 
.A1(n_309),
.A2(n_310),
.B(n_302),
.Y(n_312)
);

INVxp67_ASAP7_75t_L g310 ( 
.A(n_298),
.Y(n_310)
);

OAI31xp33_ASAP7_75t_L g313 ( 
.A1(n_312),
.A2(n_306),
.A3(n_301),
.B(n_6),
.Y(n_313)
);

OAI21xp5_ASAP7_75t_SL g314 ( 
.A1(n_313),
.A2(n_4),
.B(n_5),
.Y(n_314)
);

AOI322xp5_ASAP7_75t_L g315 ( 
.A1(n_314),
.A2(n_311),
.A3(n_5),
.B1(n_6),
.B2(n_7),
.C1(n_8),
.C2(n_9),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_315),
.B(n_4),
.C(n_5),
.Y(n_316)
);

OAI211xp5_ASAP7_75t_L g317 ( 
.A1(n_316),
.A2(n_4),
.B(n_5),
.C(n_6),
.Y(n_317)
);

A2O1A1O1Ixp25_ASAP7_75t_L g318 ( 
.A1(n_317),
.A2(n_6),
.B(n_7),
.C(n_8),
.D(n_9),
.Y(n_318)
);

AOI21xp5_ASAP7_75t_L g319 ( 
.A1(n_318),
.A2(n_7),
.B(n_314),
.Y(n_319)
);


endmodule