module fake_jpeg_31678_n_165 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_165);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_165;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_93;
wire n_54;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_140;
wire n_82;
wire n_155;
wire n_118;
wire n_96;

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_16),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_19),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_25),
.Y(n_52)
);

BUFx10_ASAP7_75t_L g53 ( 
.A(n_5),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_28),
.Y(n_54)
);

INVx11_ASAP7_75t_L g55 ( 
.A(n_6),
.Y(n_55)
);

OR2x2_ASAP7_75t_L g56 ( 
.A(n_6),
.B(n_38),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_37),
.Y(n_57)
);

CKINVDCx16_ASAP7_75t_R g58 ( 
.A(n_0),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_0),
.B(n_13),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_36),
.Y(n_60)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_34),
.Y(n_61)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_47),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_44),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_9),
.Y(n_64)
);

CKINVDCx16_ASAP7_75t_R g65 ( 
.A(n_3),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_41),
.Y(n_66)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_32),
.Y(n_67)
);

CKINVDCx14_ASAP7_75t_R g68 ( 
.A(n_39),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_24),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_49),
.Y(n_70)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_8),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_10),
.Y(n_72)
);

INVx5_ASAP7_75t_L g73 ( 
.A(n_55),
.Y(n_73)
);

INVx5_ASAP7_75t_L g85 ( 
.A(n_73),
.Y(n_85)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_62),
.Y(n_74)
);

INVx5_ASAP7_75t_L g96 ( 
.A(n_74),
.Y(n_96)
);

INVx8_ASAP7_75t_L g75 ( 
.A(n_67),
.Y(n_75)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_75),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_56),
.B(n_1),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_76),
.B(n_77),
.Y(n_83)
);

INVx3_ASAP7_75t_SL g77 ( 
.A(n_67),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_50),
.Y(n_78)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_78),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_50),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_79),
.B(n_53),
.Y(n_89)
);

OR2x2_ASAP7_75t_L g80 ( 
.A(n_56),
.B(n_1),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_80),
.B(n_81),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_53),
.Y(n_81)
);

A2O1A1Ixp33_ASAP7_75t_L g84 ( 
.A1(n_80),
.A2(n_65),
.B(n_58),
.C(n_57),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_84),
.B(n_2),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_81),
.B(n_64),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_87),
.B(n_93),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g101 ( 
.A(n_89),
.B(n_2),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_77),
.A2(n_71),
.B1(n_62),
.B2(n_61),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_90),
.A2(n_91),
.B1(n_92),
.B2(n_82),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_77),
.A2(n_71),
.B1(n_62),
.B2(n_61),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_74),
.A2(n_72),
.B1(n_68),
.B2(n_53),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_75),
.B(n_59),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_78),
.A2(n_55),
.B1(n_57),
.B2(n_54),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_94),
.A2(n_66),
.B1(n_63),
.B2(n_51),
.Y(n_106)
);

BUFx12_ASAP7_75t_L g95 ( 
.A(n_73),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_95),
.B(n_70),
.Y(n_99)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_88),
.Y(n_97)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_97),
.Y(n_135)
);

OAI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_88),
.A2(n_79),
.B1(n_52),
.B2(n_60),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_98),
.A2(n_107),
.B1(n_8),
.B2(n_9),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_99),
.B(n_102),
.Y(n_116)
);

INVx5_ASAP7_75t_L g100 ( 
.A(n_85),
.Y(n_100)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_100),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_101),
.B(n_106),
.Y(n_121)
);

CKINVDCx16_ASAP7_75t_R g102 ( 
.A(n_94),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_103),
.B(n_111),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_86),
.B(n_69),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_104),
.B(n_112),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_85),
.Y(n_108)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_108),
.Y(n_120)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_82),
.Y(n_109)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_109),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_83),
.B(n_3),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_110),
.B(n_7),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_84),
.B(n_22),
.C(n_46),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_96),
.B(n_4),
.Y(n_112)
);

NOR3xp33_ASAP7_75t_SL g113 ( 
.A(n_95),
.B(n_4),
.C(n_5),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_113),
.B(n_115),
.Y(n_128)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_95),
.Y(n_114)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_114),
.Y(n_132)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_87),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_105),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_117),
.B(n_123),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_101),
.B(n_7),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_125),
.B(n_130),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_126),
.A2(n_12),
.B1(n_17),
.B2(n_18),
.Y(n_139)
);

AOI22x1_ASAP7_75t_L g127 ( 
.A1(n_107),
.A2(n_27),
.B1(n_45),
.B2(n_43),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_127),
.A2(n_20),
.B1(n_30),
.B2(n_31),
.Y(n_143)
);

AOI21xp5_ASAP7_75t_L g129 ( 
.A1(n_110),
.A2(n_23),
.B(n_42),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_L g138 ( 
.A1(n_129),
.A2(n_11),
.B(n_12),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_100),
.B(n_10),
.Y(n_130)
);

AND2x6_ASAP7_75t_L g131 ( 
.A(n_98),
.B(n_26),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_131),
.B(n_133),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_108),
.B(n_11),
.Y(n_133)
);

OAI32xp33_ASAP7_75t_L g134 ( 
.A1(n_102),
.A2(n_21),
.A3(n_40),
.B1(n_14),
.B2(n_15),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_134),
.B(n_33),
.Y(n_147)
);

NAND2x1_ASAP7_75t_SL g136 ( 
.A(n_116),
.B(n_29),
.Y(n_136)
);

NAND3xp33_ASAP7_75t_L g151 ( 
.A(n_136),
.B(n_146),
.C(n_147),
.Y(n_151)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_122),
.Y(n_137)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_137),
.Y(n_154)
);

OR2x2_ASAP7_75t_L g152 ( 
.A(n_138),
.B(n_142),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_139),
.B(n_140),
.Y(n_150)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_132),
.Y(n_140)
);

INVx4_ASAP7_75t_L g142 ( 
.A(n_119),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_143),
.B(n_149),
.C(n_127),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_135),
.Y(n_146)
);

AOI21xp5_ASAP7_75t_SL g148 ( 
.A1(n_121),
.A2(n_35),
.B(n_48),
.Y(n_148)
);

AO22x1_ASAP7_75t_SL g153 ( 
.A1(n_148),
.A2(n_134),
.B1(n_129),
.B2(n_131),
.Y(n_153)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_120),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_153),
.A2(n_126),
.B1(n_145),
.B2(n_144),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_155),
.B(n_139),
.C(n_124),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_156),
.B(n_157),
.C(n_158),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_152),
.B(n_141),
.C(n_150),
.Y(n_157)
);

O2A1O1Ixp33_ASAP7_75t_SL g159 ( 
.A1(n_157),
.A2(n_150),
.B(n_153),
.C(n_151),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_159),
.B(n_138),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_SL g162 ( 
.A1(n_161),
.A2(n_148),
.B(n_136),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_162),
.A2(n_160),
.B1(n_118),
.B2(n_128),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_163),
.B(n_154),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_164),
.B(n_149),
.Y(n_165)
);


endmodule