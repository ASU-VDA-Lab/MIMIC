module fake_jpeg_17962_n_24 (n_3, n_2, n_1, n_0, n_4, n_5, n_24);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_24;

wire n_13;
wire n_21;
wire n_10;
wire n_23;
wire n_6;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_16;
wire n_9;
wire n_11;
wire n_17;
wire n_12;
wire n_8;
wire n_15;
wire n_7;

NOR2xp33_ASAP7_75t_L g6 ( 
.A(n_0),
.B(n_4),
.Y(n_6)
);

BUFx12f_ASAP7_75t_L g7 ( 
.A(n_2),
.Y(n_7)
);

INVx6_ASAP7_75t_L g8 ( 
.A(n_2),
.Y(n_8)
);

AOI22xp33_ASAP7_75t_SL g9 ( 
.A1(n_4),
.A2(n_2),
.B1(n_5),
.B2(n_3),
.Y(n_9)
);

NOR2xp33_ASAP7_75t_L g10 ( 
.A(n_0),
.B(n_5),
.Y(n_10)
);

XOR2xp5_ASAP7_75t_L g11 ( 
.A(n_6),
.B(n_0),
.Y(n_11)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_11),
.B(n_15),
.Y(n_16)
);

OAI22xp5_ASAP7_75t_SL g12 ( 
.A1(n_9),
.A2(n_1),
.B1(n_3),
.B2(n_8),
.Y(n_12)
);

OAI22xp5_ASAP7_75t_L g17 ( 
.A1(n_12),
.A2(n_8),
.B1(n_1),
.B2(n_7),
.Y(n_17)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_7),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_SL g18 ( 
.A(n_13),
.B(n_14),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g14 ( 
.A(n_6),
.B(n_10),
.Y(n_14)
);

XNOR2xp5_ASAP7_75t_L g15 ( 
.A(n_10),
.B(n_1),
.Y(n_15)
);

AOI21xp5_ASAP7_75t_L g21 ( 
.A1(n_17),
.A2(n_19),
.B(n_7),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_11),
.B(n_7),
.C(n_8),
.Y(n_19)
);

AOI22xp33_ASAP7_75t_SL g20 ( 
.A1(n_19),
.A2(n_7),
.B1(n_15),
.B2(n_18),
.Y(n_20)
);

OAI21xp5_ASAP7_75t_L g23 ( 
.A1(n_20),
.A2(n_21),
.B(n_22),
.Y(n_23)
);

AOI21xp5_ASAP7_75t_L g22 ( 
.A1(n_16),
.A2(n_9),
.B(n_11),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_23),
.Y(n_24)
);


endmodule