module fake_jpeg_8488_n_107 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_107);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_107;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_106;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

BUFx3_ASAP7_75t_L g11 ( 
.A(n_0),
.Y(n_11)
);

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_7),
.Y(n_12)
);

BUFx4f_ASAP7_75t_SL g13 ( 
.A(n_5),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_0),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_9),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_7),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_1),
.B(n_8),
.Y(n_17)
);

INVx8_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

BUFx16f_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_17),
.B(n_1),
.Y(n_24)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_24),
.Y(n_45)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_22),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_25),
.B(n_26),
.Y(n_46)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_22),
.Y(n_27)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_27),
.Y(n_39)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_22),
.Y(n_28)
);

INVxp67_ASAP7_75t_L g34 ( 
.A(n_28),
.Y(n_34)
);

BUFx24_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

INVxp67_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_17),
.B(n_2),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_30),
.Y(n_44)
);

INVx1_ASAP7_75t_SL g31 ( 
.A(n_13),
.Y(n_31)
);

AND2x2_ASAP7_75t_L g41 ( 
.A(n_31),
.B(n_14),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

INVx5_ASAP7_75t_L g36 ( 
.A(n_32),
.Y(n_36)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

HB1xp67_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

OAI22xp33_ASAP7_75t_L g35 ( 
.A1(n_33),
.A2(n_19),
.B1(n_12),
.B2(n_23),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_35),
.A2(n_31),
.B1(n_21),
.B2(n_15),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g37 ( 
.A1(n_24),
.A2(n_19),
.B1(n_18),
.B2(n_16),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_L g52 ( 
.A1(n_37),
.A2(n_42),
.B1(n_14),
.B2(n_20),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_41),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_L g42 ( 
.A1(n_26),
.A2(n_18),
.B1(n_20),
.B2(n_23),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_45),
.B(n_27),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_48),
.B(n_49),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_45),
.B(n_27),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_46),
.B(n_16),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_50),
.B(n_56),
.Y(n_65)
);

O2A1O1Ixp33_ASAP7_75t_L g64 ( 
.A1(n_52),
.A2(n_54),
.B(n_34),
.C(n_3),
.Y(n_64)
);

OAI21xp5_ASAP7_75t_SL g53 ( 
.A1(n_41),
.A2(n_21),
.B(n_15),
.Y(n_53)
);

OAI21xp5_ASAP7_75t_L g70 ( 
.A1(n_53),
.A2(n_55),
.B(n_57),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_41),
.B(n_13),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_55),
.B(n_2),
.Y(n_71)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_35),
.Y(n_56)
);

INVxp67_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

INVx1_ASAP7_75t_SL g67 ( 
.A(n_57),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_36),
.A2(n_25),
.B1(n_32),
.B2(n_29),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_58),
.A2(n_59),
.B1(n_40),
.B2(n_39),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_36),
.A2(n_29),
.B1(n_3),
.B2(n_4),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_60),
.B(n_63),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_47),
.A2(n_39),
.B1(n_43),
.B2(n_44),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_62),
.A2(n_51),
.B1(n_59),
.B2(n_58),
.Y(n_77)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_51),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_64),
.B(n_66),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_48),
.Y(n_66)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_49),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_68),
.B(n_69),
.Y(n_76)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_54),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_70),
.B(n_29),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_71),
.B(n_3),
.Y(n_74)
);

XNOR2xp5_ASAP7_75t_L g72 ( 
.A(n_70),
.B(n_53),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_72),
.B(n_74),
.Y(n_87)
);

BUFx12_ASAP7_75t_L g75 ( 
.A(n_67),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_75),
.B(n_77),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_66),
.B(n_34),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_78),
.B(n_80),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_SL g85 ( 
.A1(n_79),
.A2(n_61),
.B(n_62),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_68),
.B(n_4),
.Y(n_80)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_78),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_82),
.A2(n_86),
.B1(n_88),
.B2(n_65),
.Y(n_92)
);

AO22x1_ASAP7_75t_L g84 ( 
.A1(n_73),
.A2(n_64),
.B1(n_69),
.B2(n_60),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_84),
.A2(n_63),
.B1(n_75),
.B2(n_4),
.Y(n_94)
);

XOR2xp5_ASAP7_75t_L g91 ( 
.A(n_85),
.B(n_77),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_76),
.A2(n_65),
.B1(n_63),
.B2(n_67),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_81),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_85),
.B(n_72),
.C(n_87),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_90),
.B(n_91),
.C(n_93),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_92),
.B(n_94),
.Y(n_97)
);

XNOR2xp5_ASAP7_75t_L g93 ( 
.A(n_89),
.B(n_80),
.Y(n_93)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_91),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_95),
.B(n_83),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_90),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_98),
.B(n_75),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_L g102 ( 
.A1(n_99),
.A2(n_100),
.B(n_96),
.Y(n_102)
);

OAI22x1_ASAP7_75t_L g100 ( 
.A1(n_97),
.A2(n_84),
.B1(n_88),
.B2(n_86),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_101),
.B(n_96),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_L g105 ( 
.A1(n_102),
.A2(n_103),
.B(n_38),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_SL g104 ( 
.A1(n_103),
.A2(n_5),
.B(n_6),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_104),
.B(n_105),
.Y(n_106)
);

XNOR2xp5_ASAP7_75t_L g107 ( 
.A(n_106),
.B(n_10),
.Y(n_107)
);


endmodule