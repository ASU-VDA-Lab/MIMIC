module real_jpeg_28933_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_201;
wire n_114;
wire n_68;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_249;
wire n_166;
wire n_176;
wire n_215;
wire n_221;
wire n_194;
wire n_104;
wire n_153;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_237;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_243;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_200;
wire n_48;
wire n_164;
wire n_184;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_155;
wire n_120;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_242;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_238;
wire n_67;
wire n_79;
wire n_178;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_172;
wire n_160;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_222;
wire n_19;
wire n_148;
wire n_118;
wire n_220;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_205;
wire n_117;
wire n_193;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_225;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_97;
wire n_75;
wire n_187;
wire n_34;
wire n_230;
wire n_190;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_202;
wire n_213;
wire n_167;
wire n_244;
wire n_216;
wire n_133;
wire n_179;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_127;
wire n_210;
wire n_206;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_181;
wire n_85;
wire n_101;
wire n_182;
wire n_96;
wire n_89;

INVx5_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

INVx11_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_1),
.A2(n_59),
.B1(n_60),
.B2(n_61),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_1),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_L g62 ( 
.A1(n_1),
.A2(n_55),
.B1(n_56),
.B2(n_59),
.Y(n_62)
);

O2A1O1Ixp33_ASAP7_75t_SL g96 ( 
.A1(n_1),
.A2(n_10),
.B(n_56),
.C(n_97),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_2),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_3),
.A2(n_54),
.B1(n_55),
.B2(n_56),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_3),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_L g152 ( 
.A1(n_3),
.A2(n_54),
.B1(n_60),
.B2(n_61),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_SL g190 ( 
.A1(n_3),
.A2(n_38),
.B1(n_39),
.B2(n_54),
.Y(n_190)
);

AOI22xp33_ASAP7_75t_SL g200 ( 
.A1(n_3),
.A2(n_26),
.B1(n_32),
.B2(n_54),
.Y(n_200)
);

AOI22xp33_ASAP7_75t_L g77 ( 
.A1(n_4),
.A2(n_60),
.B1(n_61),
.B2(n_78),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_4),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_4),
.A2(n_55),
.B1(n_56),
.B2(n_78),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_L g146 ( 
.A1(n_4),
.A2(n_38),
.B1(n_39),
.B2(n_78),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_4),
.A2(n_26),
.B1(n_32),
.B2(n_78),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g30 ( 
.A1(n_5),
.A2(n_26),
.B1(n_31),
.B2(n_32),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_5),
.Y(n_31)
);

AOI22xp33_ASAP7_75t_L g86 ( 
.A1(n_5),
.A2(n_31),
.B1(n_38),
.B2(n_39),
.Y(n_86)
);

BUFx10_ASAP7_75t_L g55 ( 
.A(n_6),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_7),
.A2(n_26),
.B1(n_32),
.B2(n_84),
.Y(n_83)
);

CKINVDCx16_ASAP7_75t_R g84 ( 
.A(n_7),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_L g47 ( 
.A1(n_8),
.A2(n_38),
.B1(n_39),
.B2(n_48),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_8),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_8),
.A2(n_26),
.B1(n_32),
.B2(n_48),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_8),
.A2(n_48),
.B1(n_60),
.B2(n_61),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_L g34 ( 
.A1(n_9),
.A2(n_26),
.B1(n_32),
.B2(n_35),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_9),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_9),
.A2(n_35),
.B1(n_38),
.B2(n_39),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_10),
.Y(n_98)
);

OAI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_10),
.A2(n_55),
.B1(n_56),
.B2(n_98),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_10),
.B(n_58),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_10),
.B(n_38),
.Y(n_180)
);

A2O1A1O1Ixp25_ASAP7_75t_L g182 ( 
.A1(n_10),
.A2(n_38),
.B(n_42),
.C(n_180),
.D(n_183),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_10),
.B(n_69),
.Y(n_187)
);

OAI21xp33_ASAP7_75t_L g211 ( 
.A1(n_10),
.A2(n_25),
.B(n_193),
.Y(n_211)
);

A2O1A1O1Ixp25_ASAP7_75t_L g221 ( 
.A1(n_10),
.A2(n_61),
.B(n_74),
.C(n_110),
.D(n_222),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_10),
.B(n_61),
.Y(n_222)
);

O2A1O1Ixp33_ASAP7_75t_L g42 ( 
.A1(n_11),
.A2(n_38),
.B(n_43),
.C(n_46),
.Y(n_42)
);

INVx11_ASAP7_75t_L g45 ( 
.A(n_11),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g46 ( 
.A1(n_11),
.A2(n_26),
.B1(n_32),
.B2(n_45),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_12),
.A2(n_55),
.B1(n_56),
.B2(n_64),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_12),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_12),
.A2(n_60),
.B1(n_61),
.B2(n_64),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g192 ( 
.A1(n_12),
.A2(n_26),
.B1(n_32),
.B2(n_64),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_12),
.A2(n_38),
.B1(n_39),
.B2(n_64),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g37 ( 
.A1(n_13),
.A2(n_38),
.B1(n_39),
.B2(n_40),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_13),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_13),
.A2(n_40),
.B1(n_60),
.B2(n_61),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_L g168 ( 
.A1(n_13),
.A2(n_26),
.B1(n_32),
.B2(n_40),
.Y(n_168)
);

BUFx24_ASAP7_75t_L g60 ( 
.A(n_14),
.Y(n_60)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_15),
.Y(n_70)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_15),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_15),
.A2(n_60),
.B1(n_61),
.B2(n_72),
.Y(n_75)
);

INVx11_ASAP7_75t_SL g27 ( 
.A(n_16),
.Y(n_27)
);

XNOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_133),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_132),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_111),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_21),
.B(n_111),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_79),
.C(n_87),
.Y(n_21)
);

XNOR2xp5_ASAP7_75t_SL g154 ( 
.A(n_22),
.B(n_79),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_SL g22 ( 
.A(n_23),
.B(n_50),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_23),
.B(n_52),
.C(n_65),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_36),
.Y(n_23)
);

XOR2xp5_ASAP7_75t_L g140 ( 
.A(n_24),
.B(n_36),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_29),
.B1(n_33),
.B2(n_34),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_25),
.A2(n_34),
.B1(n_81),
.B2(n_83),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_25),
.Y(n_101)
);

AOI21xp5_ASAP7_75t_L g119 ( 
.A1(n_25),
.A2(n_81),
.B(n_83),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_25),
.A2(n_81),
.B1(n_103),
.B2(n_168),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_L g191 ( 
.A1(n_25),
.A2(n_192),
.B(n_193),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_25),
.B(n_195),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g25 ( 
.A(n_26),
.B(n_28),
.Y(n_25)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_26),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_26),
.B(n_44),
.Y(n_181)
);

INVx11_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_30),
.Y(n_29)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_30),
.A2(n_82),
.B1(n_101),
.B2(n_102),
.Y(n_100)
);

AOI32xp33_ASAP7_75t_L g179 ( 
.A1(n_32),
.A2(n_39),
.A3(n_45),
.B1(n_180),
.B2(n_181),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_SL g212 ( 
.A(n_32),
.B(n_213),
.Y(n_212)
);

INVx11_ASAP7_75t_L g82 ( 
.A(n_33),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_33),
.B(n_98),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_L g36 ( 
.A1(n_37),
.A2(n_41),
.B1(n_47),
.B2(n_49),
.Y(n_36)
);

OAI21xp5_ASAP7_75t_SL g143 ( 
.A1(n_37),
.A2(n_49),
.B(n_144),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g43 ( 
.A(n_38),
.B(n_44),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_38),
.A2(n_39),
.B1(n_70),
.B2(n_71),
.Y(n_69)
);

AOI32xp33_ASAP7_75t_L g229 ( 
.A1(n_38),
.A2(n_60),
.A3(n_222),
.B1(n_230),
.B2(n_231),
.Y(n_229)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

NAND2xp33_ASAP7_75t_SL g231 ( 
.A(n_39),
.B(n_71),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_41),
.A2(n_47),
.B1(n_49),
.B2(n_86),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_SL g241 ( 
.A1(n_41),
.A2(n_242),
.B(n_243),
.Y(n_241)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_42),
.A2(n_46),
.B1(n_116),
.B2(n_117),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_42),
.B(n_145),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_42),
.A2(n_46),
.B1(n_224),
.B2(n_225),
.Y(n_223)
);

INVx11_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_46),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_49),
.B(n_146),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_L g189 ( 
.A1(n_49),
.A2(n_144),
.B(n_190),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_SL g206 ( 
.A(n_49),
.B(n_98),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_51),
.A2(n_52),
.B1(n_65),
.B2(n_66),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_53),
.A2(n_57),
.B1(n_58),
.B2(n_63),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_53),
.Y(n_91)
);

INVx13_ASAP7_75t_L g56 ( 
.A(n_55),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_57),
.B(n_94),
.Y(n_93)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_57),
.Y(n_125)
);

AOI21xp5_ASAP7_75t_L g147 ( 
.A1(n_57),
.A2(n_148),
.B(n_149),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_SL g57 ( 
.A(n_58),
.B(n_62),
.Y(n_57)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_58),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_58),
.B(n_94),
.Y(n_127)
);

OAI21xp33_ASAP7_75t_L g97 ( 
.A1(n_59),
.A2(n_61),
.B(n_98),
.Y(n_97)
);

INVx5_ASAP7_75t_SL g61 ( 
.A(n_60),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_63),
.Y(n_126)
);

CKINVDCx16_ASAP7_75t_R g65 ( 
.A(n_66),
.Y(n_65)
);

OAI21xp5_ASAP7_75t_L g66 ( 
.A1(n_67),
.A2(n_68),
.B(n_73),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_67),
.A2(n_68),
.B1(n_106),
.B2(n_129),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_68),
.B(n_77),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_L g166 ( 
.A1(n_68),
.A2(n_73),
.B(n_152),
.Y(n_166)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_69),
.B(n_75),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_69),
.A2(n_74),
.B1(n_108),
.B2(n_151),
.Y(n_150)
);

INVx6_ASAP7_75t_L g230 ( 
.A(n_71),
.Y(n_230)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_74),
.B(n_76),
.Y(n_73)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_74),
.Y(n_106)
);

CKINVDCx16_ASAP7_75t_R g76 ( 
.A(n_77),
.Y(n_76)
);

XNOR2xp5_ASAP7_75t_L g79 ( 
.A(n_80),
.B(n_85),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_80),
.B(n_85),
.Y(n_121)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_81),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_SL g207 ( 
.A1(n_81),
.A2(n_200),
.B(n_208),
.Y(n_207)
);

INVx11_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_82),
.B(n_194),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_86),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_87),
.A2(n_88),
.B1(n_154),
.B2(n_155),
.Y(n_153)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_95),
.C(n_104),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_89),
.A2(n_90),
.B1(n_104),
.B2(n_105),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_90),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_L g90 ( 
.A1(n_91),
.A2(n_92),
.B(n_93),
.Y(n_90)
);

XOR2xp5_ASAP7_75t_L g138 ( 
.A(n_95),
.B(n_139),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_99),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_96),
.A2(n_99),
.B1(n_100),
.B2(n_164),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_96),
.Y(n_164)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_101),
.A2(n_199),
.B1(n_201),
.B2(n_202),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_103),
.Y(n_102)
);

CKINVDCx16_ASAP7_75t_R g104 ( 
.A(n_105),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_SL g105 ( 
.A1(n_106),
.A2(n_107),
.B(n_109),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_108),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_L g111 ( 
.A(n_112),
.B(n_131),
.Y(n_111)
);

XNOR2xp5_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_120),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_114),
.A2(n_115),
.B1(n_118),
.B2(n_119),
.Y(n_113)
);

CKINVDCx14_ASAP7_75t_R g114 ( 
.A(n_115),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_119),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_121),
.A2(n_122),
.B1(n_123),
.B2(n_130),
.Y(n_120)
);

CKINVDCx16_ASAP7_75t_R g130 ( 
.A(n_121),
.Y(n_130)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

XNOR2xp5_ASAP7_75t_SL g123 ( 
.A(n_124),
.B(n_128),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_SL g124 ( 
.A1(n_125),
.A2(n_126),
.B(n_127),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_127),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_172),
.Y(n_133)
);

INVxp33_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

AOI21xp5_ASAP7_75t_L g135 ( 
.A1(n_136),
.A2(n_156),
.B(n_171),
.Y(n_135)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_136),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_153),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g171 ( 
.A(n_137),
.B(n_153),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_140),
.C(n_141),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_L g157 ( 
.A(n_138),
.B(n_158),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_140),
.B(n_141),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_147),
.C(n_150),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_142),
.A2(n_143),
.B1(n_150),
.B2(n_162),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_143),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_SL g160 ( 
.A(n_147),
.B(n_161),
.Y(n_160)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_150),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_152),
.Y(n_151)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_154),
.Y(n_155)
);

AND2x2_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_159),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_157),
.B(n_159),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_163),
.C(n_165),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_160),
.B(n_248),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_163),
.B(n_165),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_167),
.C(n_169),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_SL g236 ( 
.A(n_166),
.B(n_237),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_167),
.A2(n_169),
.B1(n_170),
.B2(n_238),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_167),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_168),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_170),
.Y(n_169)
);

NOR3xp33_ASAP7_75t_L g172 ( 
.A(n_173),
.B(n_250),
.C(n_251),
.Y(n_172)
);

AOI21xp5_ASAP7_75t_L g173 ( 
.A1(n_174),
.A2(n_245),
.B(n_249),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_SL g174 ( 
.A1(n_175),
.A2(n_233),
.B(n_244),
.Y(n_174)
);

AOI21xp5_ASAP7_75t_L g175 ( 
.A1(n_176),
.A2(n_217),
.B(n_232),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_SL g176 ( 
.A1(n_177),
.A2(n_196),
.B(n_216),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_184),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_178),
.B(n_184),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_182),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_179),
.B(n_182),
.Y(n_203)
);

CKINVDCx14_ASAP7_75t_R g243 ( 
.A(n_183),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_191),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_186),
.A2(n_187),
.B1(n_188),
.B2(n_189),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_186),
.B(n_189),
.C(n_191),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_187),
.Y(n_186)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_190),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_192),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_195),
.Y(n_194)
);

AOI21xp5_ASAP7_75t_L g196 ( 
.A1(n_197),
.A2(n_204),
.B(n_215),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_203),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_SL g215 ( 
.A(n_198),
.B(n_203),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_200),
.Y(n_199)
);

AOI21xp5_ASAP7_75t_L g227 ( 
.A1(n_202),
.A2(n_209),
.B(n_228),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_SL g204 ( 
.A1(n_205),
.A2(n_210),
.B(n_214),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_207),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_206),
.B(n_207),
.Y(n_214)
);

INVxp67_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_211),
.B(n_212),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_219),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_SL g232 ( 
.A(n_218),
.B(n_219),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_226),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_223),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_221),
.B(n_223),
.C(n_226),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_225),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_SL g226 ( 
.A(n_227),
.B(n_229),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_227),
.B(n_229),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_235),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_234),
.B(n_235),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_239),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_236),
.B(n_240),
.C(n_241),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_241),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_247),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_SL g249 ( 
.A(n_246),
.B(n_247),
.Y(n_249)
);


endmodule