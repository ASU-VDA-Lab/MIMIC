module fake_jpeg_19493_n_37 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_37);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_37;

wire n_21;
wire n_33;
wire n_23;
wire n_27;
wire n_22;
wire n_19;
wire n_20;
wire n_18;
wire n_35;
wire n_34;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_36;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_32;
wire n_15;

INVx3_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

BUFx5_ASAP7_75t_L g16 ( 
.A(n_13),
.Y(n_16)
);

INVx6_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

INVx11_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_15),
.B(n_0),
.Y(n_20)
);

AND2x2_ASAP7_75t_L g27 ( 
.A(n_20),
.B(n_21),
.Y(n_27)
);

A2O1A1Ixp33_ASAP7_75t_L g21 ( 
.A1(n_19),
.A2(n_1),
.B(n_2),
.C(n_3),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_17),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_L g28 ( 
.A1(n_22),
.A2(n_23),
.B1(n_24),
.B2(n_18),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_19),
.B(n_17),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_17),
.B(n_4),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_20),
.Y(n_25)
);

OAI21xp33_ASAP7_75t_L g29 ( 
.A1(n_25),
.A2(n_26),
.B(n_16),
.Y(n_29)
);

AOI22xp33_ASAP7_75t_SL g26 ( 
.A1(n_22),
.A2(n_15),
.B1(n_18),
.B2(n_16),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g30 ( 
.A1(n_28),
.A2(n_18),
.B1(n_8),
.B2(n_9),
.Y(n_30)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_29),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_30),
.Y(n_33)
);

XOR2xp5_ASAP7_75t_L g31 ( 
.A(n_27),
.B(n_7),
.Y(n_31)
);

AOI22xp33_ASAP7_75t_SL g34 ( 
.A1(n_32),
.A2(n_33),
.B1(n_29),
.B2(n_27),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_34),
.Y(n_35)
);

NAND3xp33_ASAP7_75t_L g36 ( 
.A(n_35),
.B(n_31),
.C(n_11),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_L g37 ( 
.A1(n_36),
.A2(n_10),
.B1(n_12),
.B2(n_14),
.Y(n_37)
);


endmodule