module fake_ariane_2061_n_1858 (n_83, n_8, n_56, n_60, n_170, n_160, n_64, n_119, n_124, n_167, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_149, n_34, n_158, n_69, n_95, n_92, n_143, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_152, n_120, n_169, n_106, n_12, n_53, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_166, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_159, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_148, n_164, n_52, n_157, n_135, n_73, n_77, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_151, n_136, n_28, n_80, n_146, n_97, n_154, n_142, n_161, n_14, n_163, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_1858);

input n_83;
input n_8;
input n_56;
input n_60;
input n_170;
input n_160;
input n_64;
input n_119;
input n_124;
input n_167;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_149;
input n_34;
input n_158;
input n_69;
input n_95;
input n_92;
input n_143;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_166;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_159;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_164;
input n_52;
input n_157;
input n_135;
input n_73;
input n_77;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_151;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1858;

wire n_913;
wire n_1681;
wire n_1486;
wire n_1507;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_610;
wire n_245;
wire n_1713;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_187;
wire n_1463;
wire n_1238;
wire n_1515;
wire n_817;
wire n_1837;
wire n_924;
wire n_781;
wire n_1566;
wire n_189;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_524;
wire n_1214;
wire n_634;
wire n_1839;
wire n_1246;
wire n_1138;
wire n_214;
wire n_1853;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_232;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1835;
wire n_1457;
wire n_377;
wire n_1682;
wire n_1836;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_945;
wire n_958;
wire n_813;
wire n_419;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1184;
wire n_202;
wire n_1535;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1277;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_672;
wire n_740;
wire n_1283;
wire n_1736;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_645;
wire n_242;
wire n_331;
wire n_559;
wire n_267;
wire n_495;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_200;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1847;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1851;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_587;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_352;
wire n_206;
wire n_899;
wire n_1703;
wire n_611;
wire n_1295;
wire n_1850;
wire n_365;
wire n_238;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_192;
wire n_661;
wire n_1751;
wire n_300;
wire n_533;
wire n_438;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_1811;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_1840;
wire n_376;
wire n_512;
wire n_1597;
wire n_1771;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_237;
wire n_780;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_209;
wire n_490;
wire n_1461;
wire n_1391;
wire n_225;
wire n_1599;
wire n_1006;
wire n_1830;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_1838;
wire n_1594;
wire n_680;
wire n_287;
wire n_1716;
wire n_302;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_212;
wire n_444;
wire n_851;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_1819;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_182;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_1833;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_460;
wire n_1555;
wire n_1842;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_992;
wire n_966;
wire n_955;
wire n_1182;
wire n_794;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_179;
wire n_1292;
wire n_1178;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_306;
wire n_203;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_437;
wire n_337;
wire n_274;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1787;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_1717;
wire n_1812;
wire n_824;
wire n_428;
wire n_892;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_1855;
wire n_990;
wire n_1623;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_1780;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1825;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1832;
wire n_1841;
wire n_1680;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_1731;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_698;
wire n_1674;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_172;
wire n_1058;
wire n_347;
wire n_1042;
wire n_183;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_205;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_1728;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_1817;
wire n_348;
wire n_552;
wire n_670;
wire n_1826;
wire n_379;
wire n_264;
wire n_441;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_1743;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_194;
wire n_1802;
wire n_1163;
wire n_186;
wire n_1795;
wire n_1384;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1648;
wire n_1413;
wire n_855;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_647;
wire n_1423;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_529;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1828;
wire n_1798;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_1105;
wire n_547;
wire n_439;
wire n_604;
wire n_677;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_699;
wire n_727;
wire n_301;
wire n_1726;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_325;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1693;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1823;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_221;
wire n_321;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_845;
wire n_888;
wire n_1649;
wire n_1677;
wire n_1297;
wire n_178;
wire n_551;
wire n_417;
wire n_1708;
wire n_343;
wire n_1222;
wire n_1844;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_534;
wire n_1791;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_451;
wire n_745;
wire n_1741;
wire n_1572;
wire n_1793;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_769;
wire n_1797;
wire n_1753;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_982;
wire n_1800;
wire n_915;
wire n_215;
wire n_1075;
wire n_454;
wire n_298;
wire n_1331;
wire n_1529;
wire n_1227;
wire n_655;
wire n_1734;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_509;
wire n_1854;
wire n_666;
wire n_1747;
wire n_430;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_456;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_873;
wire n_1301;
wire n_1748;
wire n_1243;
wire n_1400;
wire n_342;
wire n_1466;
wire n_1513;
wire n_1527;
wire n_358;
wire n_1783;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1668;
wire n_1605;
wire n_1078;
wire n_266;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_1786;
wire n_480;
wire n_1327;
wire n_1475;
wire n_211;
wire n_642;
wire n_1804;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_1757;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_1632;
wire n_1769;
wire n_474;
wire n_805;
wire n_295;
wire n_1658;
wire n_190;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_180;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1258;
wire n_197;
wire n_640;
wire n_463;
wire n_1476;
wire n_1524;
wire n_1733;
wire n_1856;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_1807;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_1784;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_283;
wire n_806;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_1824;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_1822;
wire n_682;
wire n_1616;
wire n_819;
wire n_586;
wire n_1429;
wire n_1324;
wire n_1778;
wire n_1776;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1759;
wire n_1829;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_1815;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_198;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_1852;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_1288;
wire n_1201;
wire n_173;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_1367;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1023;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_467;
wire n_1511;
wire n_1422;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_538;
wire n_1517;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1773;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_810;
wire n_1290;
wire n_181;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_236;
wire n_683;
wire n_601;
wire n_565;
wire n_628;
wire n_1300;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_414;
wire n_571;
wire n_1521;
wire n_1694;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_409;
wire n_171;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1444;
wire n_1803;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_1739;
wire n_1814;
wire n_532;
wire n_1789;
wire n_763;
wire n_540;
wire n_216;
wire n_692;
wire n_1857;
wire n_984;
wire n_1687;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_1816;
wire n_1756;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_1772;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_493;
wire n_1311;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1335;
wire n_1715;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_1785;
wire n_792;
wire n_1262;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1183;
wire n_1326;
wire n_1805;
wire n_981;
wire n_1110;
wire n_1758;
wire n_243;
wire n_1407;
wire n_185;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_184;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_1054;
wire n_508;
wire n_1679;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_191;
wire n_1834;
wire n_978;
wire n_1011;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_1536;
wire n_1471;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_176;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_541;
wire n_499;
wire n_1775;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_1663;
wire n_1625;
wire n_318;
wire n_1458;
wire n_244;
wire n_679;
wire n_1630;
wire n_220;
wire n_663;
wire n_1720;
wire n_443;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_1735;
wire n_1788;
wire n_391;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_765;
wire n_1809;
wire n_1843;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_898;
wire n_857;
wire n_363;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_1755;
wire n_1285;
wire n_193;
wire n_733;
wire n_761;
wire n_731;
wire n_336;
wire n_1813;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1106;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_1770;
wire n_701;
wire n_1003;
wire n_1125;
wire n_1710;
wire n_309;
wire n_1344;
wire n_1390;
wire n_401;
wire n_485;
wire n_1792;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_567;
wire n_369;
wire n_240;
wire n_1727;
wire n_1575;
wire n_1848;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_188;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_1845;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1806;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_1696;
wire n_498;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1831;
wire n_1497;
wire n_459;
wire n_1136;
wire n_1782;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1316;
wire n_175;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_1781;
wire n_709;
wire n_809;
wire n_1686;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_199;
wire n_217;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_308;
wire n_1223;
wire n_201;
wire n_1768;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_948;
wire n_922;
wire n_1004;
wire n_1810;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_1764;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_196;
wire n_1337;
wire n_774;
wire n_933;
wire n_1779;
wire n_596;
wire n_954;
wire n_1168;
wire n_1821;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_252;
wire n_664;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1732;
wire n_415;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1799;
wire n_1126;
wire n_195;
wire n_1846;
wire n_938;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_946;
wire n_757;
wire n_375;
wire n_1655;
wire n_1818;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_265;
wire n_1583;
wire n_1604;
wire n_208;
wire n_1631;
wire n_1702;
wire n_174;
wire n_275;
wire n_1794;
wire n_1375;
wire n_204;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_1827;
wire n_866;
wire n_246;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_1569;
wire n_548;
wire n_289;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_177;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1228;
wire n_1244;
wire n_1796;
wire n_411;
wire n_484;
wire n_849;
wire n_1820;
wire n_357;
wire n_412;
wire n_1251;
wire n_447;
wire n_1421;
wire n_1762;
wire n_1233;
wire n_1808;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_4),
.Y(n_171)
);

BUFx10_ASAP7_75t_L g172 ( 
.A(n_60),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_9),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_151),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_159),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_136),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_75),
.Y(n_177)
);

INVx1_ASAP7_75t_SL g178 ( 
.A(n_78),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_169),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_30),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_18),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_1),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_120),
.Y(n_183)
);

INVx1_ASAP7_75t_SL g184 ( 
.A(n_13),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_150),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_60),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_43),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_143),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_163),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_145),
.Y(n_190)
);

BUFx10_ASAP7_75t_L g191 ( 
.A(n_98),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_119),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_144),
.Y(n_193)
);

INVx1_ASAP7_75t_SL g194 ( 
.A(n_8),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_94),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_18),
.Y(n_196)
);

BUFx2_ASAP7_75t_L g197 ( 
.A(n_11),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_29),
.Y(n_198)
);

INVx1_ASAP7_75t_SL g199 ( 
.A(n_106),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_95),
.Y(n_200)
);

BUFx3_ASAP7_75t_L g201 ( 
.A(n_147),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_5),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_24),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_2),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_122),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_81),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_63),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_14),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_110),
.Y(n_209)
);

BUFx8_ASAP7_75t_SL g210 ( 
.A(n_166),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_142),
.Y(n_211)
);

BUFx3_ASAP7_75t_L g212 ( 
.A(n_30),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_149),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_54),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_108),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_115),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_160),
.Y(n_217)
);

BUFx10_ASAP7_75t_L g218 ( 
.A(n_1),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_39),
.Y(n_219)
);

BUFx2_ASAP7_75t_L g220 ( 
.A(n_0),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_31),
.Y(n_221)
);

CKINVDCx16_ASAP7_75t_R g222 ( 
.A(n_58),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_85),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_4),
.Y(n_224)
);

INVxp67_ASAP7_75t_L g225 ( 
.A(n_128),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_26),
.Y(n_226)
);

BUFx6f_ASAP7_75t_L g227 ( 
.A(n_113),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_15),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_116),
.Y(n_229)
);

BUFx3_ASAP7_75t_L g230 ( 
.A(n_13),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_45),
.Y(n_231)
);

BUFx2_ASAP7_75t_SL g232 ( 
.A(n_101),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_86),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_126),
.Y(n_234)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_140),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_33),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_7),
.Y(n_237)
);

BUFx3_ASAP7_75t_L g238 ( 
.A(n_158),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_5),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_92),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_114),
.Y(n_241)
);

BUFx6f_ASAP7_75t_L g242 ( 
.A(n_82),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_3),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_31),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_58),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_168),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_28),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_56),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_14),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_8),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_44),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_12),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_19),
.Y(n_253)
);

BUFx3_ASAP7_75t_L g254 ( 
.A(n_131),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_111),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_52),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_91),
.Y(n_257)
);

INVx2_ASAP7_75t_SL g258 ( 
.A(n_134),
.Y(n_258)
);

BUFx10_ASAP7_75t_L g259 ( 
.A(n_56),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_42),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_103),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_21),
.Y(n_262)
);

INVx1_ASAP7_75t_SL g263 ( 
.A(n_148),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_69),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_50),
.Y(n_265)
);

INVx1_ASAP7_75t_SL g266 ( 
.A(n_42),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_15),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_132),
.Y(n_268)
);

BUFx6f_ASAP7_75t_L g269 ( 
.A(n_123),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_80),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_133),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_76),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_25),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_89),
.Y(n_274)
);

BUFx8_ASAP7_75t_SL g275 ( 
.A(n_57),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_47),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_9),
.Y(n_277)
);

INVxp33_ASAP7_75t_SL g278 ( 
.A(n_36),
.Y(n_278)
);

BUFx10_ASAP7_75t_L g279 ( 
.A(n_61),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_170),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_104),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_139),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_71),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_167),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_127),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_34),
.Y(n_286)
);

CKINVDCx11_ASAP7_75t_R g287 ( 
.A(n_37),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_55),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_157),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_50),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_96),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_97),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_65),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_79),
.Y(n_294)
);

BUFx6f_ASAP7_75t_L g295 ( 
.A(n_74),
.Y(n_295)
);

BUFx6f_ASAP7_75t_L g296 ( 
.A(n_125),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_25),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_107),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_68),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_32),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_20),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_0),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_155),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_162),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_129),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_64),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_88),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_45),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_44),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_7),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_36),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_102),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_20),
.Y(n_313)
);

BUFx5_ASAP7_75t_L g314 ( 
.A(n_29),
.Y(n_314)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_164),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_93),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_100),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_109),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_17),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_40),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_28),
.Y(n_321)
);

CKINVDCx16_ASAP7_75t_R g322 ( 
.A(n_146),
.Y(n_322)
);

CKINVDCx16_ASAP7_75t_R g323 ( 
.A(n_54),
.Y(n_323)
);

INVx2_ASAP7_75t_L g324 ( 
.A(n_6),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_66),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_32),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_40),
.Y(n_327)
);

INVx2_ASAP7_75t_SL g328 ( 
.A(n_154),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_49),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_67),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_55),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_124),
.Y(n_332)
);

BUFx3_ASAP7_75t_L g333 ( 
.A(n_156),
.Y(n_333)
);

INVx2_ASAP7_75t_SL g334 ( 
.A(n_38),
.Y(n_334)
);

INVx2_ASAP7_75t_L g335 ( 
.A(n_3),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_17),
.Y(n_336)
);

INVx1_ASAP7_75t_SL g337 ( 
.A(n_70),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_152),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g339 ( 
.A(n_19),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_16),
.Y(n_340)
);

INVxp33_ASAP7_75t_SL g341 ( 
.A(n_287),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_275),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_314),
.Y(n_343)
);

INVxp67_ASAP7_75t_SL g344 ( 
.A(n_212),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_210),
.Y(n_345)
);

CKINVDCx20_ASAP7_75t_R g346 ( 
.A(n_216),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_222),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_314),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_278),
.B(n_2),
.Y(n_349)
);

CKINVDCx20_ASAP7_75t_R g350 ( 
.A(n_231),
.Y(n_350)
);

INVxp67_ASAP7_75t_SL g351 ( 
.A(n_212),
.Y(n_351)
);

HB1xp67_ASAP7_75t_L g352 ( 
.A(n_197),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_323),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_314),
.Y(n_354)
);

CKINVDCx16_ASAP7_75t_R g355 ( 
.A(n_322),
.Y(n_355)
);

INVxp33_ASAP7_75t_SL g356 ( 
.A(n_220),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_334),
.B(n_6),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_314),
.Y(n_358)
);

INVx2_ASAP7_75t_L g359 ( 
.A(n_314),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_219),
.Y(n_360)
);

BUFx2_ASAP7_75t_L g361 ( 
.A(n_230),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_236),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_314),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g364 ( 
.A(n_311),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_243),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_314),
.Y(n_366)
);

INVxp33_ASAP7_75t_L g367 ( 
.A(n_196),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_314),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_324),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_244),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_245),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_324),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_L g373 ( 
.A(n_334),
.B(n_10),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_335),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_335),
.Y(n_375)
);

HB1xp67_ASAP7_75t_L g376 ( 
.A(n_171),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_249),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_235),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_235),
.Y(n_379)
);

INVx2_ASAP7_75t_L g380 ( 
.A(n_201),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_L g381 ( 
.A(n_230),
.B(n_174),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_315),
.Y(n_382)
);

CKINVDCx16_ASAP7_75t_R g383 ( 
.A(n_191),
.Y(n_383)
);

CKINVDCx20_ASAP7_75t_R g384 ( 
.A(n_331),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_251),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_253),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_262),
.Y(n_387)
);

HB1xp67_ASAP7_75t_L g388 ( 
.A(n_171),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_315),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_202),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_265),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_214),
.Y(n_392)
);

NOR2xp67_ASAP7_75t_L g393 ( 
.A(n_221),
.B(n_10),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_224),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_267),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_276),
.Y(n_396)
);

NOR2xp67_ASAP7_75t_L g397 ( 
.A(n_226),
.B(n_11),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_277),
.Y(n_398)
);

INVxp67_ASAP7_75t_L g399 ( 
.A(n_228),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_288),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_237),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_290),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_173),
.Y(n_403)
);

INVxp67_ASAP7_75t_L g404 ( 
.A(n_239),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_247),
.Y(n_405)
);

INVxp67_ASAP7_75t_SL g406 ( 
.A(n_248),
.Y(n_406)
);

INVxp33_ASAP7_75t_L g407 ( 
.A(n_250),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_256),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_260),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_273),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_286),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_297),
.Y(n_412)
);

BUFx3_ASAP7_75t_L g413 ( 
.A(n_201),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_300),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_301),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_173),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_302),
.Y(n_417)
);

AND2x4_ASAP7_75t_L g418 ( 
.A(n_258),
.B(n_12),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_309),
.Y(n_419)
);

BUFx10_ASAP7_75t_L g420 ( 
.A(n_258),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_180),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_180),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_321),
.Y(n_423)
);

OAI22xp5_ASAP7_75t_L g424 ( 
.A1(n_356),
.A2(n_339),
.B1(n_208),
.B2(n_336),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_380),
.B(n_176),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_343),
.Y(n_426)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_359),
.Y(n_427)
);

HB1xp67_ASAP7_75t_L g428 ( 
.A(n_352),
.Y(n_428)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_359),
.Y(n_429)
);

BUFx6f_ASAP7_75t_L g430 ( 
.A(n_359),
.Y(n_430)
);

AOI22xp5_ASAP7_75t_L g431 ( 
.A1(n_383),
.A2(n_184),
.B1(n_194),
.B2(n_266),
.Y(n_431)
);

BUFx6f_ASAP7_75t_L g432 ( 
.A(n_343),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_348),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_348),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_354),
.Y(n_435)
);

AOI22xp5_ASAP7_75t_L g436 ( 
.A1(n_383),
.A2(n_320),
.B1(n_252),
.B2(n_181),
.Y(n_436)
);

INVx2_ASAP7_75t_L g437 ( 
.A(n_354),
.Y(n_437)
);

BUFx2_ASAP7_75t_L g438 ( 
.A(n_347),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_380),
.B(n_189),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_358),
.Y(n_440)
);

INVx2_ASAP7_75t_SL g441 ( 
.A(n_420),
.Y(n_441)
);

AND2x4_ASAP7_75t_L g442 ( 
.A(n_418),
.B(n_328),
.Y(n_442)
);

AND2x6_ASAP7_75t_L g443 ( 
.A(n_418),
.B(n_227),
.Y(n_443)
);

BUFx6f_ASAP7_75t_L g444 ( 
.A(n_358),
.Y(n_444)
);

NOR2xp33_ASAP7_75t_L g445 ( 
.A(n_413),
.B(n_225),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_380),
.B(n_193),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_363),
.Y(n_447)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_363),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_366),
.B(n_205),
.Y(n_449)
);

BUFx6f_ASAP7_75t_L g450 ( 
.A(n_366),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_368),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_368),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_413),
.B(n_209),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_378),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_378),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_379),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_345),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_379),
.Y(n_458)
);

BUFx6f_ASAP7_75t_L g459 ( 
.A(n_382),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_413),
.B(n_217),
.Y(n_460)
);

BUFx6f_ASAP7_75t_L g461 ( 
.A(n_382),
.Y(n_461)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_389),
.Y(n_462)
);

INVx3_ASAP7_75t_L g463 ( 
.A(n_418),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_389),
.Y(n_464)
);

NAND3xp33_ASAP7_75t_L g465 ( 
.A(n_357),
.B(n_340),
.C(n_327),
.Y(n_465)
);

INVx2_ASAP7_75t_L g466 ( 
.A(n_369),
.Y(n_466)
);

BUFx2_ASAP7_75t_L g467 ( 
.A(n_353),
.Y(n_467)
);

INVx2_ASAP7_75t_L g468 ( 
.A(n_369),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_372),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_372),
.Y(n_470)
);

INVx2_ASAP7_75t_L g471 ( 
.A(n_374),
.Y(n_471)
);

INVx2_ASAP7_75t_L g472 ( 
.A(n_374),
.Y(n_472)
);

INVx3_ASAP7_75t_L g473 ( 
.A(n_418),
.Y(n_473)
);

AND2x2_ASAP7_75t_L g474 ( 
.A(n_361),
.B(n_191),
.Y(n_474)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_375),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_375),
.Y(n_476)
);

NOR2xp33_ASAP7_75t_L g477 ( 
.A(n_420),
.B(n_344),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_390),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_390),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_392),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_392),
.Y(n_481)
);

HB1xp67_ASAP7_75t_L g482 ( 
.A(n_403),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_394),
.Y(n_483)
);

BUFx6f_ASAP7_75t_L g484 ( 
.A(n_394),
.Y(n_484)
);

HB1xp67_ASAP7_75t_L g485 ( 
.A(n_416),
.Y(n_485)
);

AND2x4_ASAP7_75t_L g486 ( 
.A(n_351),
.B(n_328),
.Y(n_486)
);

INVx2_ASAP7_75t_L g487 ( 
.A(n_401),
.Y(n_487)
);

BUFx2_ASAP7_75t_L g488 ( 
.A(n_421),
.Y(n_488)
);

AND2x2_ASAP7_75t_L g489 ( 
.A(n_361),
.B(n_191),
.Y(n_489)
);

HB1xp67_ASAP7_75t_L g490 ( 
.A(n_422),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_401),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_405),
.Y(n_492)
);

INVx2_ASAP7_75t_L g493 ( 
.A(n_405),
.Y(n_493)
);

INVx5_ASAP7_75t_L g494 ( 
.A(n_420),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_381),
.B(n_223),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_408),
.Y(n_496)
);

INVx3_ASAP7_75t_L g497 ( 
.A(n_408),
.Y(n_497)
);

INVx6_ASAP7_75t_L g498 ( 
.A(n_420),
.Y(n_498)
);

INVx2_ASAP7_75t_L g499 ( 
.A(n_409),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_437),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_437),
.Y(n_501)
);

INVx2_ASAP7_75t_L g502 ( 
.A(n_427),
.Y(n_502)
);

INVx2_ASAP7_75t_L g503 ( 
.A(n_427),
.Y(n_503)
);

NOR2xp33_ASAP7_75t_L g504 ( 
.A(n_441),
.B(n_355),
.Y(n_504)
);

AOI22xp33_ASAP7_75t_L g505 ( 
.A1(n_465),
.A2(n_373),
.B1(n_349),
.B2(n_407),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_441),
.B(n_355),
.Y(n_506)
);

AND3x2_ASAP7_75t_L g507 ( 
.A(n_467),
.B(n_388),
.C(n_376),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_SL g508 ( 
.A(n_441),
.B(n_477),
.Y(n_508)
);

INVx4_ASAP7_75t_L g509 ( 
.A(n_443),
.Y(n_509)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_427),
.Y(n_510)
);

OAI22xp5_ASAP7_75t_L g511 ( 
.A1(n_442),
.A2(n_326),
.B1(n_204),
.B2(n_203),
.Y(n_511)
);

INVxp67_ASAP7_75t_SL g512 ( 
.A(n_463),
.Y(n_512)
);

HB1xp67_ASAP7_75t_L g513 ( 
.A(n_428),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_SL g514 ( 
.A(n_477),
.B(n_360),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_437),
.Y(n_515)
);

INVx2_ASAP7_75t_L g516 ( 
.A(n_429),
.Y(n_516)
);

AND2x2_ASAP7_75t_L g517 ( 
.A(n_474),
.B(n_367),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_448),
.Y(n_518)
);

INVx2_ASAP7_75t_L g519 ( 
.A(n_429),
.Y(n_519)
);

AND2x2_ASAP7_75t_L g520 ( 
.A(n_474),
.B(n_489),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_448),
.Y(n_521)
);

NAND2xp33_ASAP7_75t_SL g522 ( 
.A(n_488),
.B(n_362),
.Y(n_522)
);

NAND3xp33_ASAP7_75t_L g523 ( 
.A(n_426),
.B(n_397),
.C(n_393),
.Y(n_523)
);

AND2x2_ASAP7_75t_L g524 ( 
.A(n_474),
.B(n_406),
.Y(n_524)
);

INVx1_ASAP7_75t_SL g525 ( 
.A(n_438),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_448),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_429),
.Y(n_527)
);

INVx3_ASAP7_75t_L g528 ( 
.A(n_432),
.Y(n_528)
);

BUFx6f_ASAP7_75t_SL g529 ( 
.A(n_486),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_426),
.Y(n_530)
);

BUFx4f_ASAP7_75t_L g531 ( 
.A(n_443),
.Y(n_531)
);

HB1xp67_ASAP7_75t_L g532 ( 
.A(n_428),
.Y(n_532)
);

INVx2_ASAP7_75t_SL g533 ( 
.A(n_489),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_L g534 ( 
.A(n_486),
.B(n_365),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_433),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_L g536 ( 
.A(n_486),
.B(n_370),
.Y(n_536)
);

AOI22xp33_ASAP7_75t_L g537 ( 
.A1(n_465),
.A2(n_397),
.B1(n_393),
.B2(n_399),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g538 ( 
.A(n_486),
.B(n_371),
.Y(n_538)
);

INVx3_ASAP7_75t_L g539 ( 
.A(n_432),
.Y(n_539)
);

INVx2_ASAP7_75t_SL g540 ( 
.A(n_489),
.Y(n_540)
);

INVx4_ASAP7_75t_L g541 ( 
.A(n_443),
.Y(n_541)
);

BUFx3_ASAP7_75t_L g542 ( 
.A(n_433),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_486),
.B(n_377),
.Y(n_543)
);

NOR2xp33_ASAP7_75t_L g544 ( 
.A(n_498),
.B(n_385),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_434),
.Y(n_545)
);

INVx2_ASAP7_75t_L g546 ( 
.A(n_432),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_434),
.Y(n_547)
);

INVxp67_ASAP7_75t_R g548 ( 
.A(n_482),
.Y(n_548)
);

INVx4_ASAP7_75t_L g549 ( 
.A(n_443),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_435),
.Y(n_550)
);

INVx2_ASAP7_75t_L g551 ( 
.A(n_432),
.Y(n_551)
);

AND2x2_ASAP7_75t_L g552 ( 
.A(n_478),
.B(n_409),
.Y(n_552)
);

INVx4_ASAP7_75t_L g553 ( 
.A(n_443),
.Y(n_553)
);

INVx4_ASAP7_75t_L g554 ( 
.A(n_443),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_L g555 ( 
.A(n_463),
.B(n_473),
.Y(n_555)
);

AND2x4_ASAP7_75t_L g556 ( 
.A(n_463),
.B(n_399),
.Y(n_556)
);

INVx3_ASAP7_75t_L g557 ( 
.A(n_432),
.Y(n_557)
);

NAND3xp33_ASAP7_75t_SL g558 ( 
.A(n_436),
.B(n_387),
.C(n_386),
.Y(n_558)
);

INVx1_ASAP7_75t_SL g559 ( 
.A(n_438),
.Y(n_559)
);

OAI22xp5_ASAP7_75t_L g560 ( 
.A1(n_442),
.A2(n_436),
.B1(n_473),
.B2(n_463),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_SL g561 ( 
.A(n_488),
.B(n_391),
.Y(n_561)
);

INVx2_ASAP7_75t_SL g562 ( 
.A(n_498),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_L g563 ( 
.A(n_463),
.B(n_395),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_440),
.Y(n_564)
);

NAND2xp33_ASAP7_75t_SL g565 ( 
.A(n_482),
.B(n_396),
.Y(n_565)
);

INVx3_ASAP7_75t_L g566 ( 
.A(n_432),
.Y(n_566)
);

INVx2_ASAP7_75t_SL g567 ( 
.A(n_498),
.Y(n_567)
);

BUFx2_ASAP7_75t_L g568 ( 
.A(n_467),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_SL g569 ( 
.A(n_485),
.B(n_398),
.Y(n_569)
);

BUFx6f_ASAP7_75t_L g570 ( 
.A(n_430),
.Y(n_570)
);

AND2x2_ASAP7_75t_L g571 ( 
.A(n_478),
.B(n_410),
.Y(n_571)
);

NOR2xp33_ASAP7_75t_L g572 ( 
.A(n_498),
.B(n_400),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_432),
.Y(n_573)
);

AND2x2_ASAP7_75t_L g574 ( 
.A(n_479),
.B(n_410),
.Y(n_574)
);

NOR2x1p5_ASAP7_75t_L g575 ( 
.A(n_457),
.B(n_402),
.Y(n_575)
);

INVx4_ASAP7_75t_L g576 ( 
.A(n_443),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_440),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_L g578 ( 
.A(n_473),
.B(n_411),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_SL g579 ( 
.A(n_485),
.B(n_175),
.Y(n_579)
);

BUFx10_ASAP7_75t_L g580 ( 
.A(n_498),
.Y(n_580)
);

INVx2_ASAP7_75t_SL g581 ( 
.A(n_498),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_L g582 ( 
.A(n_473),
.B(n_411),
.Y(n_582)
);

AND2x2_ASAP7_75t_SL g583 ( 
.A(n_442),
.B(n_227),
.Y(n_583)
);

AND2x6_ASAP7_75t_L g584 ( 
.A(n_473),
.B(n_238),
.Y(n_584)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_444),
.Y(n_585)
);

AOI22xp33_ASAP7_75t_L g586 ( 
.A1(n_442),
.A2(n_404),
.B1(n_279),
.B2(n_259),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_447),
.Y(n_587)
);

BUFx10_ASAP7_75t_L g588 ( 
.A(n_445),
.Y(n_588)
);

OAI22xp5_ASAP7_75t_L g589 ( 
.A1(n_442),
.A2(n_252),
.B1(n_198),
.B2(n_208),
.Y(n_589)
);

BUFx3_ASAP7_75t_L g590 ( 
.A(n_447),
.Y(n_590)
);

INVx3_ASAP7_75t_L g591 ( 
.A(n_444),
.Y(n_591)
);

CKINVDCx5p33_ASAP7_75t_R g592 ( 
.A(n_467),
.Y(n_592)
);

INVx2_ASAP7_75t_SL g593 ( 
.A(n_443),
.Y(n_593)
);

INVxp67_ASAP7_75t_SL g594 ( 
.A(n_430),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_451),
.Y(n_595)
);

NOR2xp33_ASAP7_75t_L g596 ( 
.A(n_445),
.B(n_495),
.Y(n_596)
);

AND2x2_ASAP7_75t_L g597 ( 
.A(n_479),
.B(n_412),
.Y(n_597)
);

NOR2xp33_ASAP7_75t_L g598 ( 
.A(n_495),
.B(n_341),
.Y(n_598)
);

AND2x2_ASAP7_75t_L g599 ( 
.A(n_480),
.B(n_412),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_451),
.Y(n_600)
);

NAND2xp33_ASAP7_75t_L g601 ( 
.A(n_443),
.B(n_175),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_SL g602 ( 
.A(n_490),
.B(n_494),
.Y(n_602)
);

OR2x2_ASAP7_75t_L g603 ( 
.A(n_424),
.B(n_404),
.Y(n_603)
);

INVx2_ASAP7_75t_L g604 ( 
.A(n_444),
.Y(n_604)
);

NOR2x1p5_ASAP7_75t_L g605 ( 
.A(n_424),
.B(n_181),
.Y(n_605)
);

OR2x6_ASAP7_75t_L g606 ( 
.A(n_487),
.B(n_493),
.Y(n_606)
);

AOI22xp33_ASAP7_75t_L g607 ( 
.A1(n_431),
.A2(n_279),
.B1(n_259),
.B2(n_218),
.Y(n_607)
);

INVx2_ASAP7_75t_L g608 ( 
.A(n_444),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_452),
.Y(n_609)
);

AOI22xp33_ASAP7_75t_L g610 ( 
.A1(n_431),
.A2(n_480),
.B1(n_481),
.B2(n_496),
.Y(n_610)
);

CKINVDCx20_ASAP7_75t_R g611 ( 
.A(n_490),
.Y(n_611)
);

INVx2_ASAP7_75t_L g612 ( 
.A(n_444),
.Y(n_612)
);

INVx4_ASAP7_75t_L g613 ( 
.A(n_494),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_SL g614 ( 
.A(n_494),
.B(n_177),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_L g615 ( 
.A(n_494),
.B(n_414),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_452),
.Y(n_616)
);

BUFx2_ASAP7_75t_L g617 ( 
.A(n_497),
.Y(n_617)
);

OR2x6_ASAP7_75t_L g618 ( 
.A(n_487),
.B(n_414),
.Y(n_618)
);

INVx2_ASAP7_75t_SL g619 ( 
.A(n_453),
.Y(n_619)
);

AOI22xp33_ASAP7_75t_L g620 ( 
.A1(n_481),
.A2(n_279),
.B1(n_259),
.B2(n_218),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_SL g621 ( 
.A(n_494),
.B(n_177),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_459),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_459),
.Y(n_623)
);

BUFx3_ASAP7_75t_L g624 ( 
.A(n_444),
.Y(n_624)
);

OR2x2_ASAP7_75t_L g625 ( 
.A(n_497),
.B(n_423),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_459),
.Y(n_626)
);

INVx4_ASAP7_75t_L g627 ( 
.A(n_494),
.Y(n_627)
);

OR2x6_ASAP7_75t_L g628 ( 
.A(n_487),
.B(n_415),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_SL g629 ( 
.A(n_494),
.B(n_179),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_L g630 ( 
.A(n_494),
.B(n_415),
.Y(n_630)
);

CKINVDCx20_ASAP7_75t_R g631 ( 
.A(n_453),
.Y(n_631)
);

INVx2_ASAP7_75t_L g632 ( 
.A(n_444),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_459),
.Y(n_633)
);

INVx2_ASAP7_75t_L g634 ( 
.A(n_450),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_SL g635 ( 
.A(n_497),
.B(n_179),
.Y(n_635)
);

INVx2_ASAP7_75t_L g636 ( 
.A(n_450),
.Y(n_636)
);

INVxp33_ASAP7_75t_L g637 ( 
.A(n_460),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_459),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_SL g639 ( 
.A(n_497),
.B(n_183),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_SL g640 ( 
.A(n_497),
.B(n_183),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_SL g641 ( 
.A(n_484),
.B(n_185),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_L g642 ( 
.A(n_483),
.B(n_417),
.Y(n_642)
);

NOR2xp33_ASAP7_75t_L g643 ( 
.A(n_460),
.B(n_417),
.Y(n_643)
);

OAI22xp33_ASAP7_75t_L g644 ( 
.A1(n_483),
.A2(n_336),
.B1(n_319),
.B2(n_187),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_459),
.Y(n_645)
);

INVx3_ASAP7_75t_L g646 ( 
.A(n_450),
.Y(n_646)
);

AOI22xp5_ASAP7_75t_L g647 ( 
.A1(n_491),
.A2(n_308),
.B1(n_329),
.B2(n_326),
.Y(n_647)
);

INVx2_ASAP7_75t_L g648 ( 
.A(n_450),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_459),
.Y(n_649)
);

INVx2_ASAP7_75t_L g650 ( 
.A(n_450),
.Y(n_650)
);

INVx4_ASAP7_75t_L g651 ( 
.A(n_450),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_596),
.B(n_491),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_542),
.Y(n_653)
);

INVx2_ASAP7_75t_L g654 ( 
.A(n_502),
.Y(n_654)
);

NOR2xp33_ASAP7_75t_L g655 ( 
.A(n_637),
.B(n_449),
.Y(n_655)
);

AOI22xp5_ASAP7_75t_L g656 ( 
.A1(n_520),
.A2(n_496),
.B1(n_492),
.B2(n_449),
.Y(n_656)
);

AOI22xp33_ASAP7_75t_L g657 ( 
.A1(n_583),
.A2(n_484),
.B1(n_492),
.B2(n_493),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_SL g658 ( 
.A(n_580),
.B(n_450),
.Y(n_658)
);

INVx5_ASAP7_75t_L g659 ( 
.A(n_509),
.Y(n_659)
);

NAND2xp33_ASAP7_75t_L g660 ( 
.A(n_562),
.B(n_430),
.Y(n_660)
);

INVxp67_ASAP7_75t_L g661 ( 
.A(n_525),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_542),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_SL g663 ( 
.A(n_580),
.B(n_430),
.Y(n_663)
);

INVxp67_ASAP7_75t_L g664 ( 
.A(n_559),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_L g665 ( 
.A(n_619),
.B(n_484),
.Y(n_665)
);

AOI22xp33_ASAP7_75t_L g666 ( 
.A1(n_583),
.A2(n_603),
.B1(n_605),
.B2(n_529),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_590),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_SL g668 ( 
.A(n_580),
.B(n_509),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_SL g669 ( 
.A(n_580),
.B(n_430),
.Y(n_669)
);

INVx2_ASAP7_75t_L g670 ( 
.A(n_502),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_590),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_617),
.Y(n_672)
);

INVx2_ASAP7_75t_SL g673 ( 
.A(n_517),
.Y(n_673)
);

INVx2_ASAP7_75t_L g674 ( 
.A(n_503),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_619),
.B(n_484),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_SL g676 ( 
.A(n_509),
.B(n_430),
.Y(n_676)
);

AOI22xp33_ASAP7_75t_L g677 ( 
.A1(n_583),
.A2(n_484),
.B1(n_493),
.B2(n_499),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_L g678 ( 
.A(n_556),
.B(n_484),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_530),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_556),
.B(n_484),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_L g681 ( 
.A(n_556),
.B(n_499),
.Y(n_681)
);

BUFx6f_ASAP7_75t_L g682 ( 
.A(n_531),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_530),
.Y(n_683)
);

O2A1O1Ixp33_ASAP7_75t_L g684 ( 
.A1(n_560),
.A2(n_499),
.B(n_458),
.C(n_454),
.Y(n_684)
);

CKINVDCx5p33_ASAP7_75t_R g685 ( 
.A(n_592),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_L g686 ( 
.A(n_556),
.B(n_425),
.Y(n_686)
);

BUFx6f_ASAP7_75t_SL g687 ( 
.A(n_533),
.Y(n_687)
);

AND2x2_ASAP7_75t_L g688 ( 
.A(n_517),
.B(n_346),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_SL g689 ( 
.A(n_541),
.B(n_549),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_643),
.B(n_425),
.Y(n_690)
);

BUFx3_ASAP7_75t_L g691 ( 
.A(n_531),
.Y(n_691)
);

NOR2xp33_ASAP7_75t_L g692 ( 
.A(n_533),
.B(n_439),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_L g693 ( 
.A(n_544),
.B(n_439),
.Y(n_693)
);

BUFx6f_ASAP7_75t_L g694 ( 
.A(n_531),
.Y(n_694)
);

CKINVDCx5p33_ASAP7_75t_R g695 ( 
.A(n_592),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_SL g696 ( 
.A(n_541),
.B(n_430),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_535),
.Y(n_697)
);

INVx8_ASAP7_75t_L g698 ( 
.A(n_529),
.Y(n_698)
);

AOI22xp5_ASAP7_75t_L g699 ( 
.A1(n_520),
.A2(n_454),
.B1(n_455),
.B2(n_456),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_SL g700 ( 
.A(n_541),
.B(n_461),
.Y(n_700)
);

INVx1_ASAP7_75t_SL g701 ( 
.A(n_568),
.Y(n_701)
);

INVx5_ASAP7_75t_L g702 ( 
.A(n_549),
.Y(n_702)
);

OR2x6_ASAP7_75t_L g703 ( 
.A(n_606),
.B(n_455),
.Y(n_703)
);

INVx2_ASAP7_75t_L g704 ( 
.A(n_503),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_L g705 ( 
.A(n_572),
.B(n_446),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_L g706 ( 
.A(n_504),
.B(n_446),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_512),
.B(n_456),
.Y(n_707)
);

NOR2xp33_ASAP7_75t_L g708 ( 
.A(n_540),
.B(n_458),
.Y(n_708)
);

AOI22xp5_ASAP7_75t_L g709 ( 
.A1(n_529),
.A2(n_464),
.B1(n_185),
.B2(n_305),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_L g710 ( 
.A(n_524),
.B(n_464),
.Y(n_710)
);

INVx2_ASAP7_75t_L g711 ( 
.A(n_510),
.Y(n_711)
);

INVx2_ASAP7_75t_L g712 ( 
.A(n_510),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_545),
.Y(n_713)
);

INVxp67_ASAP7_75t_L g714 ( 
.A(n_568),
.Y(n_714)
);

INVx2_ASAP7_75t_SL g715 ( 
.A(n_513),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_545),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_SL g717 ( 
.A(n_549),
.B(n_461),
.Y(n_717)
);

INVx2_ASAP7_75t_L g718 ( 
.A(n_516),
.Y(n_718)
);

INVx3_ASAP7_75t_L g719 ( 
.A(n_553),
.Y(n_719)
);

INVx2_ASAP7_75t_L g720 ( 
.A(n_516),
.Y(n_720)
);

BUFx6f_ASAP7_75t_L g721 ( 
.A(n_553),
.Y(n_721)
);

NOR3xp33_ASAP7_75t_L g722 ( 
.A(n_558),
.B(n_186),
.C(n_182),
.Y(n_722)
);

OR2x2_ASAP7_75t_L g723 ( 
.A(n_603),
.B(n_350),
.Y(n_723)
);

INVx3_ASAP7_75t_L g724 ( 
.A(n_553),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_L g725 ( 
.A(n_563),
.B(n_469),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_547),
.Y(n_726)
);

INVx2_ASAP7_75t_L g727 ( 
.A(n_519),
.Y(n_727)
);

INVx2_ASAP7_75t_SL g728 ( 
.A(n_532),
.Y(n_728)
);

NOR2xp33_ASAP7_75t_L g729 ( 
.A(n_540),
.B(n_470),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_508),
.B(n_470),
.Y(n_730)
);

AO22x2_ASAP7_75t_L g731 ( 
.A1(n_523),
.A2(n_476),
.B1(n_419),
.B2(n_423),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_552),
.B(n_476),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_547),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_550),
.Y(n_734)
);

BUFx3_ASAP7_75t_L g735 ( 
.A(n_606),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_L g736 ( 
.A(n_552),
.B(n_462),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_L g737 ( 
.A(n_571),
.B(n_462),
.Y(n_737)
);

INVx2_ASAP7_75t_SL g738 ( 
.A(n_625),
.Y(n_738)
);

AND2x2_ASAP7_75t_L g739 ( 
.A(n_548),
.B(n_364),
.Y(n_739)
);

NOR2x1p5_ASAP7_75t_L g740 ( 
.A(n_506),
.B(n_534),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_L g741 ( 
.A(n_571),
.B(n_462),
.Y(n_741)
);

INVx3_ASAP7_75t_L g742 ( 
.A(n_554),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_SL g743 ( 
.A(n_554),
.B(n_461),
.Y(n_743)
);

OR2x2_ASAP7_75t_L g744 ( 
.A(n_598),
.B(n_384),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_SL g745 ( 
.A(n_554),
.B(n_461),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_SL g746 ( 
.A(n_576),
.B(n_461),
.Y(n_746)
);

INVx2_ASAP7_75t_SL g747 ( 
.A(n_625),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_574),
.B(n_597),
.Y(n_748)
);

AND2x2_ASAP7_75t_L g749 ( 
.A(n_548),
.B(n_419),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_550),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_L g751 ( 
.A(n_574),
.B(n_466),
.Y(n_751)
);

AOI22xp5_ASAP7_75t_L g752 ( 
.A1(n_536),
.A2(n_195),
.B1(n_192),
.B2(n_188),
.Y(n_752)
);

NOR2xp33_ASAP7_75t_L g753 ( 
.A(n_538),
.B(n_543),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_SL g754 ( 
.A(n_576),
.B(n_588),
.Y(n_754)
);

AOI221xp5_ASAP7_75t_L g755 ( 
.A1(n_644),
.A2(n_198),
.B1(n_310),
.B2(n_308),
.C(n_319),
.Y(n_755)
);

INVx2_ASAP7_75t_L g756 ( 
.A(n_519),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_597),
.B(n_466),
.Y(n_757)
);

INVx1_ASAP7_75t_SL g758 ( 
.A(n_611),
.Y(n_758)
);

NAND2xp33_ASAP7_75t_L g759 ( 
.A(n_562),
.B(n_182),
.Y(n_759)
);

INVx2_ASAP7_75t_L g760 ( 
.A(n_527),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_599),
.B(n_466),
.Y(n_761)
);

AOI22xp33_ASAP7_75t_L g762 ( 
.A1(n_605),
.A2(n_461),
.B1(n_475),
.B2(n_471),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_599),
.B(n_468),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_L g764 ( 
.A(n_610),
.B(n_468),
.Y(n_764)
);

O2A1O1Ixp5_ASAP7_75t_L g765 ( 
.A1(n_641),
.A2(n_475),
.B(n_472),
.C(n_471),
.Y(n_765)
);

INVxp67_ASAP7_75t_L g766 ( 
.A(n_522),
.Y(n_766)
);

NOR2xp33_ASAP7_75t_L g767 ( 
.A(n_514),
.B(n_461),
.Y(n_767)
);

INVx2_ASAP7_75t_L g768 ( 
.A(n_527),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_L g769 ( 
.A(n_588),
.B(n_468),
.Y(n_769)
);

BUFx6f_ASAP7_75t_L g770 ( 
.A(n_576),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_588),
.B(n_471),
.Y(n_771)
);

INVx2_ASAP7_75t_L g772 ( 
.A(n_500),
.Y(n_772)
);

NOR2x1p5_ASAP7_75t_L g773 ( 
.A(n_507),
.B(n_342),
.Y(n_773)
);

O2A1O1Ixp33_ASAP7_75t_L g774 ( 
.A1(n_555),
.A2(n_475),
.B(n_472),
.C(n_274),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_578),
.B(n_472),
.Y(n_775)
);

INVx2_ASAP7_75t_L g776 ( 
.A(n_500),
.Y(n_776)
);

NOR3xp33_ASAP7_75t_L g777 ( 
.A(n_561),
.B(n_186),
.C(n_329),
.Y(n_777)
);

INVx2_ASAP7_75t_L g778 ( 
.A(n_501),
.Y(n_778)
);

AND2x2_ASAP7_75t_L g779 ( 
.A(n_647),
.B(n_172),
.Y(n_779)
);

INVx2_ASAP7_75t_L g780 ( 
.A(n_501),
.Y(n_780)
);

O2A1O1Ixp33_ASAP7_75t_L g781 ( 
.A1(n_582),
.A2(n_280),
.B(n_332),
.C(n_233),
.Y(n_781)
);

NOR2xp33_ASAP7_75t_L g782 ( 
.A(n_631),
.B(n_187),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_L g783 ( 
.A(n_618),
.B(n_628),
.Y(n_783)
);

INVx3_ASAP7_75t_L g784 ( 
.A(n_593),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_564),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_L g786 ( 
.A(n_618),
.B(n_178),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_564),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_L g788 ( 
.A(n_618),
.B(n_199),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_577),
.Y(n_789)
);

INVx2_ASAP7_75t_L g790 ( 
.A(n_515),
.Y(n_790)
);

INVx2_ASAP7_75t_L g791 ( 
.A(n_515),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_618),
.B(n_263),
.Y(n_792)
);

A2O1A1Ixp33_ASAP7_75t_L g793 ( 
.A1(n_505),
.A2(n_313),
.B(n_310),
.C(n_203),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_L g794 ( 
.A(n_618),
.B(n_337),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_L g795 ( 
.A(n_628),
.B(n_188),
.Y(n_795)
);

INVx4_ASAP7_75t_L g796 ( 
.A(n_606),
.Y(n_796)
);

AND2x2_ASAP7_75t_L g797 ( 
.A(n_647),
.B(n_172),
.Y(n_797)
);

NOR2xp67_ASAP7_75t_SL g798 ( 
.A(n_567),
.B(n_204),
.Y(n_798)
);

INVx2_ASAP7_75t_L g799 ( 
.A(n_518),
.Y(n_799)
);

AOI22xp33_ASAP7_75t_L g800 ( 
.A1(n_607),
.A2(n_172),
.B1(n_218),
.B2(n_333),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_SL g801 ( 
.A(n_593),
.B(n_190),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_L g802 ( 
.A(n_628),
.B(n_190),
.Y(n_802)
);

AND2x2_ASAP7_75t_L g803 ( 
.A(n_575),
.B(n_313),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_577),
.Y(n_804)
);

HB1xp67_ASAP7_75t_L g805 ( 
.A(n_628),
.Y(n_805)
);

INVx2_ASAP7_75t_L g806 ( 
.A(n_518),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_L g807 ( 
.A(n_628),
.B(n_192),
.Y(n_807)
);

INVx2_ASAP7_75t_L g808 ( 
.A(n_521),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_L g809 ( 
.A(n_587),
.B(n_195),
.Y(n_809)
);

INVx2_ASAP7_75t_L g810 ( 
.A(n_521),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_587),
.Y(n_811)
);

AOI22xp5_ASAP7_75t_L g812 ( 
.A1(n_584),
.A2(n_211),
.B1(n_330),
.B2(n_325),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_L g813 ( 
.A(n_595),
.B(n_200),
.Y(n_813)
);

NOR2xp33_ASAP7_75t_SL g814 ( 
.A(n_584),
.B(n_320),
.Y(n_814)
);

AOI22xp5_ASAP7_75t_L g815 ( 
.A1(n_584),
.A2(n_207),
.B1(n_330),
.B2(n_325),
.Y(n_815)
);

INVx4_ASAP7_75t_L g816 ( 
.A(n_606),
.Y(n_816)
);

AND2x4_ASAP7_75t_L g817 ( 
.A(n_606),
.B(n_238),
.Y(n_817)
);

A2O1A1Ixp33_ASAP7_75t_L g818 ( 
.A1(n_595),
.A2(n_283),
.B(n_312),
.C(n_304),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_SL g819 ( 
.A(n_570),
.B(n_200),
.Y(n_819)
);

NOR2xp33_ASAP7_75t_SL g820 ( 
.A(n_661),
.B(n_584),
.Y(n_820)
);

AO22x1_ASAP7_75t_L g821 ( 
.A1(n_685),
.A2(n_584),
.B1(n_511),
.B2(n_589),
.Y(n_821)
);

O2A1O1Ixp33_ASAP7_75t_L g822 ( 
.A1(n_793),
.A2(n_569),
.B(n_579),
.C(n_639),
.Y(n_822)
);

BUFx6f_ASAP7_75t_L g823 ( 
.A(n_682),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_L g824 ( 
.A(n_655),
.B(n_586),
.Y(n_824)
);

INVx2_ASAP7_75t_L g825 ( 
.A(n_654),
.Y(n_825)
);

INVx1_ASAP7_75t_SL g826 ( 
.A(n_701),
.Y(n_826)
);

NAND2xp33_ASAP7_75t_L g827 ( 
.A(n_721),
.B(n_567),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_L g828 ( 
.A(n_655),
.B(n_642),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_L g829 ( 
.A(n_753),
.B(n_584),
.Y(n_829)
);

INVx2_ASAP7_75t_L g830 ( 
.A(n_654),
.Y(n_830)
);

AOI21xp5_ASAP7_75t_L g831 ( 
.A1(n_693),
.A2(n_581),
.B(n_594),
.Y(n_831)
);

BUFx6f_ASAP7_75t_L g832 ( 
.A(n_682),
.Y(n_832)
);

AOI21xp5_ASAP7_75t_L g833 ( 
.A1(n_705),
.A2(n_581),
.B(n_652),
.Y(n_833)
);

OR2x2_ASAP7_75t_SL g834 ( 
.A(n_744),
.B(n_523),
.Y(n_834)
);

INVx2_ASAP7_75t_L g835 ( 
.A(n_670),
.Y(n_835)
);

INVx1_ASAP7_75t_SL g836 ( 
.A(n_758),
.Y(n_836)
);

AOI21xp5_ASAP7_75t_L g837 ( 
.A1(n_690),
.A2(n_602),
.B(n_614),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_753),
.B(n_706),
.Y(n_838)
);

AOI21xp5_ASAP7_75t_L g839 ( 
.A1(n_660),
.A2(n_629),
.B(n_621),
.Y(n_839)
);

AOI21xp5_ASAP7_75t_L g840 ( 
.A1(n_660),
.A2(n_627),
.B(n_613),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_L g841 ( 
.A(n_692),
.B(n_584),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_679),
.Y(n_842)
);

AOI21xp5_ASAP7_75t_L g843 ( 
.A1(n_725),
.A2(n_627),
.B(n_613),
.Y(n_843)
);

AND2x2_ASAP7_75t_L g844 ( 
.A(n_664),
.B(n_575),
.Y(n_844)
);

OAI321xp33_ASAP7_75t_L g845 ( 
.A1(n_779),
.A2(n_537),
.A3(n_620),
.B1(n_616),
.B2(n_609),
.C(n_600),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_SL g846 ( 
.A(n_721),
.B(n_770),
.Y(n_846)
);

AOI21xp5_ASAP7_75t_L g847 ( 
.A1(n_658),
.A2(n_627),
.B(n_613),
.Y(n_847)
);

INVx4_ASAP7_75t_L g848 ( 
.A(n_698),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_692),
.B(n_600),
.Y(n_849)
);

OAI22xp5_ASAP7_75t_L g850 ( 
.A1(n_748),
.A2(n_609),
.B1(n_616),
.B2(n_635),
.Y(n_850)
);

OAI21xp5_ASAP7_75t_L g851 ( 
.A1(n_765),
.A2(n_526),
.B(n_650),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_L g852 ( 
.A(n_738),
.B(n_526),
.Y(n_852)
);

OAI21xp5_ASAP7_75t_L g853 ( 
.A1(n_676),
.A2(n_634),
.B(n_650),
.Y(n_853)
);

OAI21xp33_ASAP7_75t_L g854 ( 
.A1(n_755),
.A2(n_640),
.B(n_615),
.Y(n_854)
);

NOR2xp33_ASAP7_75t_L g855 ( 
.A(n_673),
.B(n_565),
.Y(n_855)
);

INVxp67_ASAP7_75t_L g856 ( 
.A(n_749),
.Y(n_856)
);

BUFx6f_ASAP7_75t_L g857 ( 
.A(n_682),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_L g858 ( 
.A(n_747),
.B(n_686),
.Y(n_858)
);

BUFx6f_ASAP7_75t_L g859 ( 
.A(n_682),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_L g860 ( 
.A(n_708),
.B(n_528),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_L g861 ( 
.A(n_708),
.B(n_528),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_683),
.Y(n_862)
);

INVx2_ASAP7_75t_SL g863 ( 
.A(n_685),
.Y(n_863)
);

A2O1A1Ixp33_ASAP7_75t_L g864 ( 
.A1(n_697),
.A2(n_645),
.B(n_649),
.C(n_622),
.Y(n_864)
);

INVx2_ASAP7_75t_L g865 ( 
.A(n_674),
.Y(n_865)
);

AOI21xp5_ASAP7_75t_L g866 ( 
.A1(n_658),
.A2(n_608),
.B(n_612),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_713),
.Y(n_867)
);

AOI21xp5_ASAP7_75t_L g868 ( 
.A1(n_663),
.A2(n_608),
.B(n_612),
.Y(n_868)
);

AOI21xp5_ASAP7_75t_L g869 ( 
.A1(n_663),
.A2(n_585),
.B(n_604),
.Y(n_869)
);

AOI22xp33_ASAP7_75t_L g870 ( 
.A1(n_797),
.A2(n_601),
.B1(n_649),
.B2(n_623),
.Y(n_870)
);

O2A1O1Ixp33_ASAP7_75t_L g871 ( 
.A1(n_793),
.A2(n_630),
.B(n_646),
.C(n_591),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_729),
.B(n_710),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_729),
.B(n_528),
.Y(n_873)
);

OAI21xp5_ASAP7_75t_L g874 ( 
.A1(n_676),
.A2(n_551),
.B(n_648),
.Y(n_874)
);

BUFx6f_ASAP7_75t_L g875 ( 
.A(n_694),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_656),
.B(n_539),
.Y(n_876)
);

AND2x2_ASAP7_75t_L g877 ( 
.A(n_688),
.B(n_714),
.Y(n_877)
);

AOI21xp5_ASAP7_75t_L g878 ( 
.A1(n_669),
.A2(n_573),
.B(n_648),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_740),
.B(n_539),
.Y(n_879)
);

NOR2xp33_ASAP7_75t_R g880 ( 
.A(n_695),
.B(n_557),
.Y(n_880)
);

AOI21x1_ASAP7_75t_L g881 ( 
.A1(n_696),
.A2(n_717),
.B(n_700),
.Y(n_881)
);

AOI21x1_ASAP7_75t_L g882 ( 
.A1(n_696),
.A2(n_622),
.B(n_623),
.Y(n_882)
);

O2A1O1Ixp33_ASAP7_75t_L g883 ( 
.A1(n_681),
.A2(n_646),
.B(n_566),
.C(n_591),
.Y(n_883)
);

OAI21xp5_ASAP7_75t_L g884 ( 
.A1(n_700),
.A2(n_551),
.B(n_573),
.Y(n_884)
);

INVx2_ASAP7_75t_L g885 ( 
.A(n_704),
.Y(n_885)
);

O2A1O1Ixp33_ASAP7_75t_L g886 ( 
.A1(n_769),
.A2(n_591),
.B(n_646),
.C(n_566),
.Y(n_886)
);

OAI21xp33_ASAP7_75t_L g887 ( 
.A1(n_752),
.A2(n_557),
.B(n_566),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_SL g888 ( 
.A(n_721),
.B(n_570),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_716),
.Y(n_889)
);

AOI21xp5_ASAP7_75t_L g890 ( 
.A1(n_669),
.A2(n_546),
.B(n_585),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_726),
.Y(n_891)
);

A2O1A1Ixp33_ASAP7_75t_L g892 ( 
.A1(n_733),
.A2(n_633),
.B(n_645),
.C(n_638),
.Y(n_892)
);

NOR2xp33_ASAP7_75t_L g893 ( 
.A(n_672),
.B(n_651),
.Y(n_893)
);

AOI21xp5_ASAP7_75t_L g894 ( 
.A1(n_668),
.A2(n_546),
.B(n_636),
.Y(n_894)
);

OAI21xp5_ASAP7_75t_L g895 ( 
.A1(n_717),
.A2(n_604),
.B(n_632),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_L g896 ( 
.A(n_732),
.B(n_557),
.Y(n_896)
);

INVx2_ASAP7_75t_SL g897 ( 
.A(n_695),
.Y(n_897)
);

BUFx3_ASAP7_75t_L g898 ( 
.A(n_715),
.Y(n_898)
);

O2A1O1Ixp33_ASAP7_75t_L g899 ( 
.A1(n_771),
.A2(n_638),
.B(n_633),
.C(n_626),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_SL g900 ( 
.A(n_721),
.B(n_570),
.Y(n_900)
);

AOI22xp5_ASAP7_75t_L g901 ( 
.A1(n_666),
.A2(n_651),
.B1(n_626),
.B2(n_624),
.Y(n_901)
);

AOI22xp5_ASAP7_75t_L g902 ( 
.A1(n_703),
.A2(n_624),
.B1(n_634),
.B2(n_632),
.Y(n_902)
);

AOI21xp5_ASAP7_75t_L g903 ( 
.A1(n_668),
.A2(n_636),
.B(n_570),
.Y(n_903)
);

INVx2_ASAP7_75t_L g904 ( 
.A(n_704),
.Y(n_904)
);

AOI21xp5_ASAP7_75t_L g905 ( 
.A1(n_775),
.A2(n_570),
.B(n_338),
.Y(n_905)
);

BUFx6f_ASAP7_75t_L g906 ( 
.A(n_694),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_L g907 ( 
.A(n_699),
.B(n_206),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_SL g908 ( 
.A(n_770),
.B(n_206),
.Y(n_908)
);

OAI21x1_ASAP7_75t_L g909 ( 
.A1(n_684),
.A2(n_257),
.B(n_303),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_L g910 ( 
.A(n_734),
.B(n_207),
.Y(n_910)
);

INVx2_ASAP7_75t_L g911 ( 
.A(n_711),
.Y(n_911)
);

AOI21xp5_ASAP7_75t_L g912 ( 
.A1(n_665),
.A2(n_338),
.B(n_211),
.Y(n_912)
);

AOI21xp5_ASAP7_75t_L g913 ( 
.A1(n_675),
.A2(n_305),
.B(n_318),
.Y(n_913)
);

INVx2_ASAP7_75t_L g914 ( 
.A(n_712),
.Y(n_914)
);

OR2x2_ASAP7_75t_L g915 ( 
.A(n_723),
.B(n_16),
.Y(n_915)
);

AOI21xp5_ASAP7_75t_L g916 ( 
.A1(n_743),
.A2(n_306),
.B(n_318),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_750),
.Y(n_917)
);

AOI21xp5_ASAP7_75t_L g918 ( 
.A1(n_743),
.A2(n_307),
.B(n_317),
.Y(n_918)
);

CKINVDCx5p33_ASAP7_75t_R g919 ( 
.A(n_687),
.Y(n_919)
);

INVx2_ASAP7_75t_L g920 ( 
.A(n_718),
.Y(n_920)
);

INVx2_ASAP7_75t_L g921 ( 
.A(n_718),
.Y(n_921)
);

AOI21xp5_ASAP7_75t_L g922 ( 
.A1(n_745),
.A2(n_307),
.B(n_317),
.Y(n_922)
);

INVx2_ASAP7_75t_L g923 ( 
.A(n_720),
.Y(n_923)
);

NOR2xp67_ASAP7_75t_L g924 ( 
.A(n_766),
.B(n_316),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_L g925 ( 
.A(n_785),
.B(n_787),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_L g926 ( 
.A(n_789),
.B(n_255),
.Y(n_926)
);

AND2x2_ASAP7_75t_SL g927 ( 
.A(n_814),
.B(n_268),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_804),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_L g929 ( 
.A(n_811),
.B(n_284),
.Y(n_929)
);

INVx2_ASAP7_75t_L g930 ( 
.A(n_720),
.Y(n_930)
);

INVx2_ASAP7_75t_L g931 ( 
.A(n_727),
.Y(n_931)
);

OR2x6_ASAP7_75t_SL g932 ( 
.A(n_795),
.B(n_213),
.Y(n_932)
);

NAND2x1_ASAP7_75t_L g933 ( 
.A(n_770),
.B(n_227),
.Y(n_933)
);

AOI21xp5_ASAP7_75t_L g934 ( 
.A1(n_745),
.A2(n_746),
.B(n_754),
.Y(n_934)
);

INVx2_ASAP7_75t_L g935 ( 
.A(n_727),
.Y(n_935)
);

A2O1A1Ixp33_ASAP7_75t_L g936 ( 
.A1(n_736),
.A2(n_333),
.B(n_254),
.C(n_232),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_737),
.Y(n_937)
);

AOI21xp5_ASAP7_75t_L g938 ( 
.A1(n_746),
.A2(n_299),
.B(n_298),
.Y(n_938)
);

A2O1A1Ixp33_ASAP7_75t_L g939 ( 
.A1(n_741),
.A2(n_254),
.B(n_296),
.C(n_227),
.Y(n_939)
);

INVx2_ASAP7_75t_L g940 ( 
.A(n_756),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_L g941 ( 
.A(n_653),
.B(n_215),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_L g942 ( 
.A(n_662),
.B(n_229),
.Y(n_942)
);

BUFx6f_ASAP7_75t_L g943 ( 
.A(n_694),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_L g944 ( 
.A(n_667),
.B(n_234),
.Y(n_944)
);

INVxp67_ASAP7_75t_R g945 ( 
.A(n_739),
.Y(n_945)
);

AOI21xp5_ASAP7_75t_L g946 ( 
.A1(n_754),
.A2(n_272),
.B(n_240),
.Y(n_946)
);

OAI21xp5_ASAP7_75t_L g947 ( 
.A1(n_678),
.A2(n_281),
.B(n_241),
.Y(n_947)
);

A2O1A1Ixp33_ASAP7_75t_L g948 ( 
.A1(n_751),
.A2(n_296),
.B(n_295),
.C(n_242),
.Y(n_948)
);

OAI21xp5_ASAP7_75t_L g949 ( 
.A1(n_680),
.A2(n_282),
.B(n_246),
.Y(n_949)
);

BUFx4f_ASAP7_75t_L g950 ( 
.A(n_698),
.Y(n_950)
);

INVx3_ASAP7_75t_L g951 ( 
.A(n_796),
.Y(n_951)
);

OAI321xp33_ASAP7_75t_L g952 ( 
.A1(n_800),
.A2(n_296),
.A3(n_295),
.B1(n_269),
.B2(n_242),
.C(n_227),
.Y(n_952)
);

INVx2_ASAP7_75t_L g953 ( 
.A(n_756),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_SL g954 ( 
.A(n_770),
.B(n_296),
.Y(n_954)
);

OAI21xp5_ASAP7_75t_L g955 ( 
.A1(n_760),
.A2(n_285),
.B(n_261),
.Y(n_955)
);

OAI21xp5_ASAP7_75t_L g956 ( 
.A1(n_760),
.A2(n_289),
.B(n_264),
.Y(n_956)
);

AOI22xp5_ASAP7_75t_L g957 ( 
.A1(n_703),
.A2(n_291),
.B1(n_270),
.B2(n_294),
.Y(n_957)
);

OAI22xp5_ASAP7_75t_L g958 ( 
.A1(n_757),
.A2(n_293),
.B1(n_292),
.B2(n_271),
.Y(n_958)
);

INVx2_ASAP7_75t_L g959 ( 
.A(n_768),
.Y(n_959)
);

BUFx6f_ASAP7_75t_L g960 ( 
.A(n_694),
.Y(n_960)
);

INVx4_ASAP7_75t_L g961 ( 
.A(n_698),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_761),
.Y(n_962)
);

AOI21xp5_ASAP7_75t_L g963 ( 
.A1(n_707),
.A2(n_296),
.B(n_295),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_SL g964 ( 
.A(n_659),
.B(n_295),
.Y(n_964)
);

CKINVDCx12_ASAP7_75t_R g965 ( 
.A(n_803),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_L g966 ( 
.A(n_671),
.B(n_21),
.Y(n_966)
);

OAI22xp5_ASAP7_75t_L g967 ( 
.A1(n_763),
.A2(n_295),
.B1(n_269),
.B2(n_242),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_772),
.Y(n_968)
);

INVx4_ASAP7_75t_L g969 ( 
.A(n_698),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_L g970 ( 
.A(n_786),
.B(n_22),
.Y(n_970)
);

AOI22xp5_ASAP7_75t_L g971 ( 
.A1(n_703),
.A2(n_242),
.B1(n_269),
.B2(n_24),
.Y(n_971)
);

O2A1O1Ixp33_ASAP7_75t_L g972 ( 
.A1(n_759),
.A2(n_22),
.B(n_23),
.C(n_26),
.Y(n_972)
);

A2O1A1Ixp33_ASAP7_75t_L g973 ( 
.A1(n_818),
.A2(n_722),
.B(n_780),
.C(n_778),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_L g974 ( 
.A(n_788),
.B(n_792),
.Y(n_974)
);

NOR2xp33_ASAP7_75t_L g975 ( 
.A(n_805),
.B(n_735),
.Y(n_975)
);

AOI22xp33_ASAP7_75t_L g976 ( 
.A1(n_731),
.A2(n_269),
.B1(n_242),
.B2(n_33),
.Y(n_976)
);

INVx3_ASAP7_75t_L g977 ( 
.A(n_796),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_SL g978 ( 
.A(n_659),
.B(n_269),
.Y(n_978)
);

OAI21xp5_ASAP7_75t_L g979 ( 
.A1(n_768),
.A2(n_72),
.B(n_161),
.Y(n_979)
);

INVx1_ASAP7_75t_L g980 ( 
.A(n_772),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_L g981 ( 
.A(n_794),
.B(n_23),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_SL g982 ( 
.A(n_659),
.B(n_27),
.Y(n_982)
);

AOI21xp5_ASAP7_75t_L g983 ( 
.A1(n_689),
.A2(n_73),
.B(n_153),
.Y(n_983)
);

NOR2xp33_ASAP7_75t_L g984 ( 
.A(n_735),
.B(n_27),
.Y(n_984)
);

O2A1O1Ixp33_ASAP7_75t_L g985 ( 
.A1(n_759),
.A2(n_34),
.B(n_35),
.C(n_37),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_SL g986 ( 
.A(n_659),
.B(n_35),
.Y(n_986)
);

NAND2xp5_ASAP7_75t_L g987 ( 
.A(n_809),
.B(n_38),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_SL g988 ( 
.A(n_702),
.B(n_719),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_SL g989 ( 
.A(n_702),
.B(n_39),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_L g990 ( 
.A(n_813),
.B(n_41),
.Y(n_990)
);

OAI21xp33_ASAP7_75t_L g991 ( 
.A1(n_782),
.A2(n_41),
.B(n_43),
.Y(n_991)
);

INVx4_ASAP7_75t_L g992 ( 
.A(n_703),
.Y(n_992)
);

OAI21xp5_ASAP7_75t_L g993 ( 
.A1(n_776),
.A2(n_87),
.B(n_141),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_SL g994 ( 
.A(n_702),
.B(n_46),
.Y(n_994)
);

AOI22xp5_ASAP7_75t_L g995 ( 
.A1(n_687),
.A2(n_816),
.B1(n_796),
.B2(n_782),
.Y(n_995)
);

AND2x2_ASAP7_75t_SL g996 ( 
.A(n_816),
.B(n_46),
.Y(n_996)
);

NOR2x1_ASAP7_75t_R g997 ( 
.A(n_728),
.B(n_47),
.Y(n_997)
);

AOI22xp5_ASAP7_75t_L g998 ( 
.A1(n_816),
.A2(n_48),
.B1(n_49),
.B2(n_51),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_L g999 ( 
.A(n_730),
.B(n_48),
.Y(n_999)
);

INVx1_ASAP7_75t_L g1000 ( 
.A(n_776),
.Y(n_1000)
);

NOR2xp33_ASAP7_75t_L g1001 ( 
.A(n_783),
.B(n_51),
.Y(n_1001)
);

CKINVDCx14_ASAP7_75t_R g1002 ( 
.A(n_709),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_L g1003 ( 
.A(n_731),
.B(n_762),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_L g1004 ( 
.A(n_838),
.B(n_731),
.Y(n_1004)
);

OAI22xp5_ASAP7_75t_L g1005 ( 
.A1(n_872),
.A2(n_812),
.B1(n_815),
.B2(n_719),
.Y(n_1005)
);

A2O1A1Ixp33_ASAP7_75t_L g1006 ( 
.A1(n_822),
.A2(n_767),
.B(n_781),
.C(n_818),
.Y(n_1006)
);

O2A1O1Ixp5_ASAP7_75t_SL g1007 ( 
.A1(n_982),
.A2(n_819),
.B(n_801),
.C(n_764),
.Y(n_1007)
);

AOI22x1_ASAP7_75t_L g1008 ( 
.A1(n_833),
.A2(n_780),
.B1(n_778),
.B2(n_810),
.Y(n_1008)
);

BUFx6f_ASAP7_75t_L g1009 ( 
.A(n_950),
.Y(n_1009)
);

O2A1O1Ixp33_ASAP7_75t_L g1010 ( 
.A1(n_991),
.A2(n_774),
.B(n_799),
.C(n_810),
.Y(n_1010)
);

O2A1O1Ixp33_ASAP7_75t_L g1011 ( 
.A1(n_828),
.A2(n_799),
.B(n_808),
.C(n_806),
.Y(n_1011)
);

OAI21x1_ASAP7_75t_L g1012 ( 
.A1(n_851),
.A2(n_808),
.B(n_806),
.Y(n_1012)
);

BUFx6f_ASAP7_75t_L g1013 ( 
.A(n_950),
.Y(n_1013)
);

O2A1O1Ixp5_ASAP7_75t_L g1014 ( 
.A1(n_982),
.A2(n_819),
.B(n_801),
.C(n_767),
.Y(n_1014)
);

OAI22xp5_ASAP7_75t_L g1015 ( 
.A1(n_849),
.A2(n_927),
.B1(n_925),
.B2(n_858),
.Y(n_1015)
);

AOI221xp5_ASAP7_75t_L g1016 ( 
.A1(n_824),
.A2(n_777),
.B1(n_807),
.B2(n_802),
.C(n_791),
.Y(n_1016)
);

INVx2_ASAP7_75t_L g1017 ( 
.A(n_959),
.Y(n_1017)
);

NOR2xp67_ASAP7_75t_L g1018 ( 
.A(n_863),
.B(n_817),
.Y(n_1018)
);

NAND3xp33_ASAP7_75t_L g1019 ( 
.A(n_972),
.B(n_798),
.C(n_657),
.Y(n_1019)
);

NOR2xp33_ASAP7_75t_SL g1020 ( 
.A(n_927),
.B(n_826),
.Y(n_1020)
);

OAI21xp5_ASAP7_75t_L g1021 ( 
.A1(n_841),
.A2(n_791),
.B(n_790),
.Y(n_1021)
);

A2O1A1Ixp33_ASAP7_75t_L g1022 ( 
.A1(n_1001),
.A2(n_790),
.B(n_724),
.C(n_742),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_L g1023 ( 
.A(n_856),
.B(n_817),
.Y(n_1023)
);

AOI21xp5_ASAP7_75t_L g1024 ( 
.A1(n_829),
.A2(n_742),
.B(n_724),
.Y(n_1024)
);

NAND2xp5_ASAP7_75t_SL g1025 ( 
.A(n_898),
.B(n_702),
.Y(n_1025)
);

NOR2xp33_ASAP7_75t_L g1026 ( 
.A(n_856),
.B(n_784),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_842),
.Y(n_1027)
);

INVx1_ASAP7_75t_L g1028 ( 
.A(n_862),
.Y(n_1028)
);

INVx1_ASAP7_75t_SL g1029 ( 
.A(n_836),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_L g1030 ( 
.A(n_937),
.B(n_677),
.Y(n_1030)
);

OAI22xp5_ASAP7_75t_L g1031 ( 
.A1(n_962),
.A2(n_742),
.B1(n_724),
.B2(n_719),
.Y(n_1031)
);

BUFx8_ASAP7_75t_L g1032 ( 
.A(n_897),
.Y(n_1032)
);

INVx2_ASAP7_75t_L g1033 ( 
.A(n_825),
.Y(n_1033)
);

AOI21xp5_ASAP7_75t_L g1034 ( 
.A1(n_831),
.A2(n_784),
.B(n_691),
.Y(n_1034)
);

AOI21xp5_ASAP7_75t_L g1035 ( 
.A1(n_860),
.A2(n_52),
.B(n_53),
.Y(n_1035)
);

AND2x4_ASAP7_75t_L g1036 ( 
.A(n_992),
.B(n_773),
.Y(n_1036)
);

INVx2_ASAP7_75t_L g1037 ( 
.A(n_830),
.Y(n_1037)
);

INVx2_ASAP7_75t_L g1038 ( 
.A(n_835),
.Y(n_1038)
);

CKINVDCx6p67_ASAP7_75t_R g1039 ( 
.A(n_965),
.Y(n_1039)
);

NAND2xp5_ASAP7_75t_L g1040 ( 
.A(n_974),
.B(n_975),
.Y(n_1040)
);

BUFx3_ASAP7_75t_L g1041 ( 
.A(n_844),
.Y(n_1041)
);

AOI21x1_ASAP7_75t_L g1042 ( 
.A1(n_882),
.A2(n_105),
.B(n_138),
.Y(n_1042)
);

AOI21xp5_ASAP7_75t_L g1043 ( 
.A1(n_861),
.A2(n_873),
.B(n_837),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_L g1044 ( 
.A(n_975),
.B(n_53),
.Y(n_1044)
);

INVx1_ASAP7_75t_L g1045 ( 
.A(n_867),
.Y(n_1045)
);

NOR3xp33_ASAP7_75t_L g1046 ( 
.A(n_821),
.B(n_57),
.C(n_59),
.Y(n_1046)
);

NOR2x1_ASAP7_75t_L g1047 ( 
.A(n_848),
.B(n_961),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_L g1048 ( 
.A(n_877),
.B(n_889),
.Y(n_1048)
);

AOI33xp33_ASAP7_75t_L g1049 ( 
.A1(n_985),
.A2(n_59),
.A3(n_61),
.B1(n_62),
.B2(n_77),
.B3(n_83),
.Y(n_1049)
);

O2A1O1Ixp33_ASAP7_75t_L g1050 ( 
.A1(n_973),
.A2(n_84),
.B(n_90),
.C(n_99),
.Y(n_1050)
);

AOI21xp5_ASAP7_75t_L g1051 ( 
.A1(n_934),
.A2(n_112),
.B(n_117),
.Y(n_1051)
);

INVx2_ASAP7_75t_L g1052 ( 
.A(n_865),
.Y(n_1052)
);

O2A1O1Ixp33_ASAP7_75t_L g1053 ( 
.A1(n_973),
.A2(n_118),
.B(n_121),
.C(n_130),
.Y(n_1053)
);

NOR2xp33_ASAP7_75t_L g1054 ( 
.A(n_834),
.B(n_135),
.Y(n_1054)
);

OAI22xp5_ASAP7_75t_L g1055 ( 
.A1(n_907),
.A2(n_137),
.B1(n_165),
.B2(n_870),
.Y(n_1055)
);

CKINVDCx5p33_ASAP7_75t_R g1056 ( 
.A(n_880),
.Y(n_1056)
);

NAND2xp5_ASAP7_75t_L g1057 ( 
.A(n_891),
.B(n_917),
.Y(n_1057)
);

OAI22xp5_ASAP7_75t_L g1058 ( 
.A1(n_870),
.A2(n_928),
.B1(n_893),
.B2(n_852),
.Y(n_1058)
);

AOI21x1_ASAP7_75t_L g1059 ( 
.A1(n_954),
.A2(n_909),
.B(n_964),
.Y(n_1059)
);

INVx1_ASAP7_75t_L g1060 ( 
.A(n_968),
.Y(n_1060)
);

AND2x2_ASAP7_75t_L g1061 ( 
.A(n_945),
.B(n_1002),
.Y(n_1061)
);

NOR2xp33_ASAP7_75t_L g1062 ( 
.A(n_1002),
.B(n_845),
.Y(n_1062)
);

O2A1O1Ixp33_ASAP7_75t_L g1063 ( 
.A1(n_987),
.A2(n_990),
.B(n_999),
.C(n_850),
.Y(n_1063)
);

INVx4_ASAP7_75t_L g1064 ( 
.A(n_848),
.Y(n_1064)
);

NAND2xp5_ASAP7_75t_L g1065 ( 
.A(n_855),
.B(n_984),
.Y(n_1065)
);

NAND2xp5_ASAP7_75t_L g1066 ( 
.A(n_855),
.B(n_984),
.Y(n_1066)
);

NAND2xp5_ASAP7_75t_L g1067 ( 
.A(n_980),
.B(n_1000),
.Y(n_1067)
);

INVx1_ASAP7_75t_L g1068 ( 
.A(n_885),
.Y(n_1068)
);

A2O1A1Ixp33_ASAP7_75t_L g1069 ( 
.A1(n_854),
.A2(n_971),
.B(n_981),
.C(n_970),
.Y(n_1069)
);

INVx1_ASAP7_75t_L g1070 ( 
.A(n_904),
.Y(n_1070)
);

INVx2_ASAP7_75t_L g1071 ( 
.A(n_911),
.Y(n_1071)
);

INVx3_ASAP7_75t_L g1072 ( 
.A(n_969),
.Y(n_1072)
);

AOI22xp5_ASAP7_75t_L g1073 ( 
.A1(n_996),
.A2(n_820),
.B1(n_976),
.B2(n_924),
.Y(n_1073)
);

AOI21xp5_ASAP7_75t_L g1074 ( 
.A1(n_886),
.A2(n_896),
.B(n_878),
.Y(n_1074)
);

OAI22xp5_ASAP7_75t_L g1075 ( 
.A1(n_893),
.A2(n_976),
.B1(n_876),
.B2(n_910),
.Y(n_1075)
);

AOI221xp5_ASAP7_75t_L g1076 ( 
.A1(n_915),
.A2(n_936),
.B1(n_956),
.B2(n_955),
.C(n_958),
.Y(n_1076)
);

INVx1_ASAP7_75t_L g1077 ( 
.A(n_914),
.Y(n_1077)
);

AND2x4_ASAP7_75t_L g1078 ( 
.A(n_992),
.B(n_951),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_L g1079 ( 
.A(n_977),
.B(n_926),
.Y(n_1079)
);

OAI22xp33_ASAP7_75t_L g1080 ( 
.A1(n_998),
.A2(n_952),
.B1(n_957),
.B2(n_929),
.Y(n_1080)
);

BUFx6f_ASAP7_75t_L g1081 ( 
.A(n_823),
.Y(n_1081)
);

AOI21xp5_ASAP7_75t_L g1082 ( 
.A1(n_868),
.A2(n_869),
.B(n_890),
.Y(n_1082)
);

NAND2xp5_ASAP7_75t_L g1083 ( 
.A(n_977),
.B(n_1003),
.Y(n_1083)
);

INVxp67_ASAP7_75t_L g1084 ( 
.A(n_966),
.Y(n_1084)
);

AOI21xp5_ASAP7_75t_L g1085 ( 
.A1(n_827),
.A2(n_866),
.B(n_883),
.Y(n_1085)
);

OAI22xp5_ASAP7_75t_L g1086 ( 
.A1(n_947),
.A2(n_949),
.B1(n_902),
.B2(n_879),
.Y(n_1086)
);

BUFx2_ASAP7_75t_L g1087 ( 
.A(n_932),
.Y(n_1087)
);

CKINVDCx6p67_ASAP7_75t_R g1088 ( 
.A(n_986),
.Y(n_1088)
);

AOI21x1_ASAP7_75t_L g1089 ( 
.A1(n_954),
.A2(n_964),
.B(n_978),
.Y(n_1089)
);

O2A1O1Ixp5_ASAP7_75t_L g1090 ( 
.A1(n_986),
.A2(n_994),
.B(n_989),
.C(n_908),
.Y(n_1090)
);

BUFx2_ASAP7_75t_L g1091 ( 
.A(n_997),
.Y(n_1091)
);

INVx2_ASAP7_75t_L g1092 ( 
.A(n_920),
.Y(n_1092)
);

AOI33xp33_ASAP7_75t_L g1093 ( 
.A1(n_871),
.A2(n_899),
.A3(n_901),
.B1(n_953),
.B2(n_940),
.B3(n_921),
.Y(n_1093)
);

AOI21xp5_ASAP7_75t_L g1094 ( 
.A1(n_894),
.A2(n_843),
.B(n_903),
.Y(n_1094)
);

INVx1_ASAP7_75t_L g1095 ( 
.A(n_923),
.Y(n_1095)
);

BUFx6f_ASAP7_75t_L g1096 ( 
.A(n_823),
.Y(n_1096)
);

NAND2xp5_ASAP7_75t_L g1097 ( 
.A(n_930),
.B(n_931),
.Y(n_1097)
);

HB1xp67_ASAP7_75t_L g1098 ( 
.A(n_823),
.Y(n_1098)
);

AND2x2_ASAP7_75t_L g1099 ( 
.A(n_941),
.B(n_942),
.Y(n_1099)
);

NOR2xp33_ASAP7_75t_L g1100 ( 
.A(n_944),
.B(n_908),
.Y(n_1100)
);

INVx3_ASAP7_75t_L g1101 ( 
.A(n_823),
.Y(n_1101)
);

INVx1_ASAP7_75t_L g1102 ( 
.A(n_935),
.Y(n_1102)
);

NOR3xp33_ASAP7_75t_SL g1103 ( 
.A(n_912),
.B(n_913),
.C(n_989),
.Y(n_1103)
);

NOR2xp67_ASAP7_75t_L g1104 ( 
.A(n_916),
.B(n_922),
.Y(n_1104)
);

AOI22xp5_ASAP7_75t_L g1105 ( 
.A1(n_994),
.A2(n_846),
.B1(n_988),
.B2(n_887),
.Y(n_1105)
);

OR2x6_ASAP7_75t_L g1106 ( 
.A(n_832),
.B(n_906),
.Y(n_1106)
);

BUFx12f_ASAP7_75t_L g1107 ( 
.A(n_832),
.Y(n_1107)
);

AND2x4_ASAP7_75t_L g1108 ( 
.A(n_832),
.B(n_906),
.Y(n_1108)
);

INVx2_ASAP7_75t_L g1109 ( 
.A(n_881),
.Y(n_1109)
);

AOI21xp5_ASAP7_75t_L g1110 ( 
.A1(n_864),
.A2(n_892),
.B(n_988),
.Y(n_1110)
);

AOI22xp33_ASAP7_75t_L g1111 ( 
.A1(n_979),
.A2(n_993),
.B1(n_918),
.B2(n_832),
.Y(n_1111)
);

INVx2_ASAP7_75t_L g1112 ( 
.A(n_857),
.Y(n_1112)
);

INVx1_ASAP7_75t_L g1113 ( 
.A(n_864),
.Y(n_1113)
);

HB1xp67_ASAP7_75t_L g1114 ( 
.A(n_857),
.Y(n_1114)
);

NAND2xp5_ASAP7_75t_L g1115 ( 
.A(n_857),
.B(n_859),
.Y(n_1115)
);

CKINVDCx11_ASAP7_75t_R g1116 ( 
.A(n_859),
.Y(n_1116)
);

BUFx6f_ASAP7_75t_L g1117 ( 
.A(n_859),
.Y(n_1117)
);

AOI21xp5_ASAP7_75t_L g1118 ( 
.A1(n_892),
.A2(n_900),
.B(n_888),
.Y(n_1118)
);

INVx2_ASAP7_75t_L g1119 ( 
.A(n_859),
.Y(n_1119)
);

BUFx6f_ASAP7_75t_L g1120 ( 
.A(n_875),
.Y(n_1120)
);

NAND2xp5_ASAP7_75t_SL g1121 ( 
.A(n_875),
.B(n_943),
.Y(n_1121)
);

INVx2_ASAP7_75t_L g1122 ( 
.A(n_875),
.Y(n_1122)
);

AOI21xp5_ASAP7_75t_L g1123 ( 
.A1(n_888),
.A2(n_900),
.B(n_839),
.Y(n_1123)
);

INVx1_ASAP7_75t_L g1124 ( 
.A(n_936),
.Y(n_1124)
);

INVx2_ASAP7_75t_L g1125 ( 
.A(n_875),
.Y(n_1125)
);

NAND2xp5_ASAP7_75t_SL g1126 ( 
.A(n_906),
.B(n_943),
.Y(n_1126)
);

AND2x4_ASAP7_75t_L g1127 ( 
.A(n_943),
.B(n_960),
.Y(n_1127)
);

O2A1O1Ixp33_ASAP7_75t_L g1128 ( 
.A1(n_939),
.A2(n_905),
.B(n_948),
.C(n_895),
.Y(n_1128)
);

AND2x4_ASAP7_75t_L g1129 ( 
.A(n_943),
.B(n_960),
.Y(n_1129)
);

HB1xp67_ASAP7_75t_L g1130 ( 
.A(n_960),
.Y(n_1130)
);

A2O1A1Ixp33_ASAP7_75t_L g1131 ( 
.A1(n_983),
.A2(n_939),
.B(n_963),
.C(n_884),
.Y(n_1131)
);

AOI21xp5_ASAP7_75t_L g1132 ( 
.A1(n_840),
.A2(n_847),
.B(n_846),
.Y(n_1132)
);

AND2x2_ASAP7_75t_L g1133 ( 
.A(n_946),
.B(n_960),
.Y(n_1133)
);

INVx2_ASAP7_75t_L g1134 ( 
.A(n_933),
.Y(n_1134)
);

INVx1_ASAP7_75t_L g1135 ( 
.A(n_853),
.Y(n_1135)
);

NOR2xp33_ASAP7_75t_SL g1136 ( 
.A(n_938),
.B(n_948),
.Y(n_1136)
);

AO32x2_ASAP7_75t_L g1137 ( 
.A1(n_967),
.A2(n_850),
.A3(n_992),
.B1(n_560),
.B2(n_619),
.Y(n_1137)
);

O2A1O1Ixp33_ASAP7_75t_L g1138 ( 
.A1(n_874),
.A2(n_838),
.B(n_596),
.C(n_872),
.Y(n_1138)
);

INVx2_ASAP7_75t_L g1139 ( 
.A(n_978),
.Y(n_1139)
);

NOR2xp67_ASAP7_75t_L g1140 ( 
.A(n_863),
.B(n_661),
.Y(n_1140)
);

BUFx16f_ASAP7_75t_R g1141 ( 
.A(n_1002),
.Y(n_1141)
);

NAND2xp5_ASAP7_75t_SL g1142 ( 
.A(n_826),
.B(n_701),
.Y(n_1142)
);

INVx1_ASAP7_75t_SL g1143 ( 
.A(n_826),
.Y(n_1143)
);

AND2x2_ASAP7_75t_L g1144 ( 
.A(n_877),
.B(n_517),
.Y(n_1144)
);

BUFx12f_ASAP7_75t_L g1145 ( 
.A(n_919),
.Y(n_1145)
);

AOI21xp5_ASAP7_75t_L g1146 ( 
.A1(n_838),
.A2(n_872),
.B(n_833),
.Y(n_1146)
);

NOR2xp33_ASAP7_75t_L g1147 ( 
.A(n_838),
.B(n_744),
.Y(n_1147)
);

OAI22x1_ASAP7_75t_L g1148 ( 
.A1(n_995),
.A2(n_605),
.B1(n_436),
.B2(n_431),
.Y(n_1148)
);

INVx2_ASAP7_75t_L g1149 ( 
.A(n_959),
.Y(n_1149)
);

NAND2xp5_ASAP7_75t_L g1150 ( 
.A(n_838),
.B(n_655),
.Y(n_1150)
);

A2O1A1Ixp33_ASAP7_75t_L g1151 ( 
.A1(n_838),
.A2(n_753),
.B(n_872),
.C(n_822),
.Y(n_1151)
);

INVx3_ASAP7_75t_L g1152 ( 
.A(n_848),
.Y(n_1152)
);

O2A1O1Ixp33_ASAP7_75t_L g1153 ( 
.A1(n_838),
.A2(n_596),
.B(n_872),
.C(n_991),
.Y(n_1153)
);

AOI21xp5_ASAP7_75t_L g1154 ( 
.A1(n_1146),
.A2(n_1151),
.B(n_1138),
.Y(n_1154)
);

AOI21xp5_ASAP7_75t_L g1155 ( 
.A1(n_1146),
.A2(n_1138),
.B(n_1153),
.Y(n_1155)
);

OR2x2_ASAP7_75t_L g1156 ( 
.A(n_1147),
.B(n_1143),
.Y(n_1156)
);

A2O1A1Ixp33_ASAP7_75t_L g1157 ( 
.A1(n_1153),
.A2(n_1100),
.B(n_1076),
.C(n_1054),
.Y(n_1157)
);

O2A1O1Ixp5_ASAP7_75t_L g1158 ( 
.A1(n_1069),
.A2(n_1055),
.B(n_1090),
.C(n_1014),
.Y(n_1158)
);

INVx2_ASAP7_75t_L g1159 ( 
.A(n_1017),
.Y(n_1159)
);

O2A1O1Ixp33_ASAP7_75t_SL g1160 ( 
.A1(n_1150),
.A2(n_1065),
.B(n_1066),
.C(n_1022),
.Y(n_1160)
);

AND2x2_ASAP7_75t_L g1161 ( 
.A(n_1144),
.B(n_1061),
.Y(n_1161)
);

NAND3x1_ASAP7_75t_L g1162 ( 
.A(n_1054),
.B(n_1062),
.C(n_1046),
.Y(n_1162)
);

INVx3_ASAP7_75t_L g1163 ( 
.A(n_1009),
.Y(n_1163)
);

A2O1A1Ixp33_ASAP7_75t_L g1164 ( 
.A1(n_1100),
.A2(n_1063),
.B(n_1073),
.C(n_1090),
.Y(n_1164)
);

OAI22xp5_ASAP7_75t_L g1165 ( 
.A1(n_1015),
.A2(n_1075),
.B1(n_1057),
.B2(n_1004),
.Y(n_1165)
);

OAI21xp5_ASAP7_75t_L g1166 ( 
.A1(n_1110),
.A2(n_1007),
.B(n_1014),
.Y(n_1166)
);

INVx1_ASAP7_75t_L g1167 ( 
.A(n_1027),
.Y(n_1167)
);

O2A1O1Ixp33_ASAP7_75t_SL g1168 ( 
.A1(n_1063),
.A2(n_1006),
.B(n_1005),
.C(n_1079),
.Y(n_1168)
);

INVx3_ASAP7_75t_L g1169 ( 
.A(n_1009),
.Y(n_1169)
);

OR2x2_ASAP7_75t_L g1170 ( 
.A(n_1048),
.B(n_1040),
.Y(n_1170)
);

A2O1A1Ixp33_ASAP7_75t_L g1171 ( 
.A1(n_1046),
.A2(n_1053),
.B(n_1050),
.C(n_1099),
.Y(n_1171)
);

NAND2xp5_ASAP7_75t_L g1172 ( 
.A(n_1030),
.B(n_1058),
.Y(n_1172)
);

OAI22xp5_ASAP7_75t_L g1173 ( 
.A1(n_1044),
.A2(n_1088),
.B1(n_1080),
.B2(n_1111),
.Y(n_1173)
);

INVx4_ASAP7_75t_L g1174 ( 
.A(n_1009),
.Y(n_1174)
);

AOI21xp5_ASAP7_75t_L g1175 ( 
.A1(n_1043),
.A2(n_1024),
.B(n_1094),
.Y(n_1175)
);

O2A1O1Ixp33_ASAP7_75t_SL g1176 ( 
.A1(n_1086),
.A2(n_1084),
.B(n_1031),
.C(n_1025),
.Y(n_1176)
);

BUFx2_ASAP7_75t_SL g1177 ( 
.A(n_1140),
.Y(n_1177)
);

OAI22xp5_ASAP7_75t_L g1178 ( 
.A1(n_1080),
.A2(n_1111),
.B1(n_1019),
.B2(n_1113),
.Y(n_1178)
);

AOI21xp5_ASAP7_75t_L g1179 ( 
.A1(n_1043),
.A2(n_1024),
.B(n_1094),
.Y(n_1179)
);

NAND2xp5_ASAP7_75t_SL g1180 ( 
.A(n_1020),
.B(n_1078),
.Y(n_1180)
);

INVx2_ASAP7_75t_SL g1181 ( 
.A(n_1032),
.Y(n_1181)
);

NAND2xp5_ASAP7_75t_L g1182 ( 
.A(n_1029),
.B(n_1142),
.Y(n_1182)
);

CKINVDCx11_ASAP7_75t_R g1183 ( 
.A(n_1145),
.Y(n_1183)
);

NAND2xp5_ASAP7_75t_L g1184 ( 
.A(n_1023),
.B(n_1028),
.Y(n_1184)
);

OAI21x1_ASAP7_75t_L g1185 ( 
.A1(n_1132),
.A2(n_1008),
.B(n_1082),
.Y(n_1185)
);

AOI21xp5_ASAP7_75t_L g1186 ( 
.A1(n_1082),
.A2(n_1132),
.B(n_1011),
.Y(n_1186)
);

BUFx12f_ASAP7_75t_L g1187 ( 
.A(n_1032),
.Y(n_1187)
);

INVx4_ASAP7_75t_L g1188 ( 
.A(n_1013),
.Y(n_1188)
);

INVxp67_ASAP7_75t_SL g1189 ( 
.A(n_1026),
.Y(n_1189)
);

AO32x1_ASAP7_75t_L g1190 ( 
.A1(n_1109),
.A2(n_1124),
.A3(n_1135),
.B1(n_1139),
.B2(n_1060),
.Y(n_1190)
);

NAND2xp5_ASAP7_75t_L g1191 ( 
.A(n_1045),
.B(n_1148),
.Y(n_1191)
);

OAI21xp5_ASAP7_75t_L g1192 ( 
.A1(n_1110),
.A2(n_1118),
.B(n_1128),
.Y(n_1192)
);

NOR2xp33_ASAP7_75t_L g1193 ( 
.A(n_1041),
.B(n_1084),
.Y(n_1193)
);

CKINVDCx20_ASAP7_75t_R g1194 ( 
.A(n_1039),
.Y(n_1194)
);

CKINVDCx20_ASAP7_75t_R g1195 ( 
.A(n_1116),
.Y(n_1195)
);

A2O1A1Ixp33_ASAP7_75t_L g1196 ( 
.A1(n_1050),
.A2(n_1053),
.B(n_1016),
.C(n_1011),
.Y(n_1196)
);

OAI21x1_ASAP7_75t_L g1197 ( 
.A1(n_1123),
.A2(n_1012),
.B(n_1085),
.Y(n_1197)
);

AO31x2_ASAP7_75t_L g1198 ( 
.A1(n_1131),
.A2(n_1118),
.A3(n_1074),
.B(n_1085),
.Y(n_1198)
);

AOI21xp5_ASAP7_75t_L g1199 ( 
.A1(n_1074),
.A2(n_1034),
.B(n_1123),
.Y(n_1199)
);

INVx2_ASAP7_75t_L g1200 ( 
.A(n_1149),
.Y(n_1200)
);

NAND2xp5_ASAP7_75t_L g1201 ( 
.A(n_1067),
.B(n_1078),
.Y(n_1201)
);

A2O1A1Ixp33_ASAP7_75t_L g1202 ( 
.A1(n_1049),
.A2(n_1010),
.B(n_1105),
.C(n_1035),
.Y(n_1202)
);

AO31x2_ASAP7_75t_L g1203 ( 
.A1(n_1034),
.A2(n_1083),
.A3(n_1051),
.B(n_1052),
.Y(n_1203)
);

NAND2xp5_ASAP7_75t_L g1204 ( 
.A(n_1068),
.B(n_1070),
.Y(n_1204)
);

AOI21xp5_ASAP7_75t_L g1205 ( 
.A1(n_1021),
.A2(n_1051),
.B(n_1128),
.Y(n_1205)
);

AND2x4_ASAP7_75t_L g1206 ( 
.A(n_1036),
.B(n_1013),
.Y(n_1206)
);

OR2x2_ASAP7_75t_L g1207 ( 
.A(n_1036),
.B(n_1077),
.Y(n_1207)
);

O2A1O1Ixp33_ASAP7_75t_SL g1208 ( 
.A1(n_1121),
.A2(n_1126),
.B(n_1115),
.C(n_1035),
.Y(n_1208)
);

OAI21xp5_ASAP7_75t_L g1209 ( 
.A1(n_1010),
.A2(n_1104),
.B(n_1103),
.Y(n_1209)
);

O2A1O1Ixp33_ASAP7_75t_L g1210 ( 
.A1(n_1136),
.A2(n_1103),
.B(n_1087),
.C(n_1091),
.Y(n_1210)
);

HB1xp67_ASAP7_75t_L g1211 ( 
.A(n_1018),
.Y(n_1211)
);

BUFx8_ASAP7_75t_L g1212 ( 
.A(n_1107),
.Y(n_1212)
);

OAI21x1_ASAP7_75t_L g1213 ( 
.A1(n_1059),
.A2(n_1042),
.B(n_1089),
.Y(n_1213)
);

OAI21x1_ASAP7_75t_L g1214 ( 
.A1(n_1133),
.A2(n_1134),
.B(n_1101),
.Y(n_1214)
);

NAND2xp5_ASAP7_75t_L g1215 ( 
.A(n_1095),
.B(n_1102),
.Y(n_1215)
);

AO22x2_ASAP7_75t_L g1216 ( 
.A1(n_1033),
.A2(n_1037),
.B1(n_1038),
.B2(n_1092),
.Y(n_1216)
);

BUFx3_ASAP7_75t_L g1217 ( 
.A(n_1108),
.Y(n_1217)
);

BUFx2_ASAP7_75t_L g1218 ( 
.A(n_1106),
.Y(n_1218)
);

HB1xp67_ASAP7_75t_L g1219 ( 
.A(n_1098),
.Y(n_1219)
);

NOR2xp33_ASAP7_75t_L g1220 ( 
.A(n_1141),
.B(n_1114),
.Y(n_1220)
);

INVx2_ASAP7_75t_L g1221 ( 
.A(n_1071),
.Y(n_1221)
);

AOI221x1_ASAP7_75t_L g1222 ( 
.A1(n_1097),
.A2(n_1101),
.B1(n_1127),
.B2(n_1108),
.C(n_1129),
.Y(n_1222)
);

INVx3_ASAP7_75t_L g1223 ( 
.A(n_1064),
.Y(n_1223)
);

CKINVDCx8_ASAP7_75t_R g1224 ( 
.A(n_1127),
.Y(n_1224)
);

NOR2xp33_ASAP7_75t_L g1225 ( 
.A(n_1098),
.B(n_1130),
.Y(n_1225)
);

OAI22x1_ASAP7_75t_L g1226 ( 
.A1(n_1112),
.A2(n_1119),
.B1(n_1122),
.B2(n_1125),
.Y(n_1226)
);

INVx1_ASAP7_75t_L g1227 ( 
.A(n_1114),
.Y(n_1227)
);

OAI21xp5_ASAP7_75t_L g1228 ( 
.A1(n_1093),
.A2(n_1130),
.B(n_1129),
.Y(n_1228)
);

INVx2_ASAP7_75t_SL g1229 ( 
.A(n_1106),
.Y(n_1229)
);

INVxp67_ASAP7_75t_SL g1230 ( 
.A(n_1081),
.Y(n_1230)
);

INVx2_ASAP7_75t_SL g1231 ( 
.A(n_1064),
.Y(n_1231)
);

O2A1O1Ixp33_ASAP7_75t_SL g1232 ( 
.A1(n_1072),
.A2(n_1152),
.B(n_1047),
.C(n_1137),
.Y(n_1232)
);

OAI21xp5_ASAP7_75t_L g1233 ( 
.A1(n_1152),
.A2(n_1072),
.B(n_1137),
.Y(n_1233)
);

NAND3xp33_ASAP7_75t_L g1234 ( 
.A(n_1081),
.B(n_1096),
.C(n_1117),
.Y(n_1234)
);

BUFx3_ASAP7_75t_L g1235 ( 
.A(n_1081),
.Y(n_1235)
);

OAI21x1_ASAP7_75t_L g1236 ( 
.A1(n_1137),
.A2(n_1096),
.B(n_1117),
.Y(n_1236)
);

AOI31xp67_ASAP7_75t_L g1237 ( 
.A1(n_1137),
.A2(n_1096),
.A3(n_1117),
.B(n_1120),
.Y(n_1237)
);

AOI21xp5_ASAP7_75t_L g1238 ( 
.A1(n_1120),
.A2(n_1146),
.B(n_1151),
.Y(n_1238)
);

AOI21x1_ASAP7_75t_L g1239 ( 
.A1(n_1120),
.A2(n_1085),
.B(n_1074),
.Y(n_1239)
);

AO31x2_ASAP7_75t_L g1240 ( 
.A1(n_1131),
.A2(n_1109),
.A3(n_1110),
.B(n_1069),
.Y(n_1240)
);

OA21x2_ASAP7_75t_L g1241 ( 
.A1(n_1094),
.A2(n_1082),
.B(n_1043),
.Y(n_1241)
);

AOI21xp5_ASAP7_75t_L g1242 ( 
.A1(n_1146),
.A2(n_1151),
.B(n_838),
.Y(n_1242)
);

AOI21xp5_ASAP7_75t_L g1243 ( 
.A1(n_1146),
.A2(n_1151),
.B(n_838),
.Y(n_1243)
);

CKINVDCx5p33_ASAP7_75t_R g1244 ( 
.A(n_1145),
.Y(n_1244)
);

O2A1O1Ixp33_ASAP7_75t_SL g1245 ( 
.A1(n_1151),
.A2(n_838),
.B(n_1153),
.C(n_1150),
.Y(n_1245)
);

AOI221xp5_ASAP7_75t_SL g1246 ( 
.A1(n_1153),
.A2(n_991),
.B1(n_1151),
.B2(n_793),
.C(n_1035),
.Y(n_1246)
);

CKINVDCx5p33_ASAP7_75t_R g1247 ( 
.A(n_1145),
.Y(n_1247)
);

INVx5_ASAP7_75t_L g1248 ( 
.A(n_1009),
.Y(n_1248)
);

OAI22xp5_ASAP7_75t_L g1249 ( 
.A1(n_1151),
.A2(n_838),
.B1(n_872),
.B2(n_1065),
.Y(n_1249)
);

BUFx6f_ASAP7_75t_L g1250 ( 
.A(n_1116),
.Y(n_1250)
);

OAI21x1_ASAP7_75t_L g1251 ( 
.A1(n_1132),
.A2(n_1008),
.B(n_1094),
.Y(n_1251)
);

AOI21xp5_ASAP7_75t_L g1252 ( 
.A1(n_1146),
.A2(n_1151),
.B(n_838),
.Y(n_1252)
);

AND2x2_ASAP7_75t_L g1253 ( 
.A(n_1147),
.B(n_517),
.Y(n_1253)
);

AOI21xp5_ASAP7_75t_L g1254 ( 
.A1(n_1146),
.A2(n_1151),
.B(n_838),
.Y(n_1254)
);

INVx1_ASAP7_75t_L g1255 ( 
.A(n_1027),
.Y(n_1255)
);

AOI21xp5_ASAP7_75t_L g1256 ( 
.A1(n_1146),
.A2(n_1151),
.B(n_838),
.Y(n_1256)
);

O2A1O1Ixp33_ASAP7_75t_L g1257 ( 
.A1(n_1065),
.A2(n_1066),
.B(n_1147),
.C(n_1151),
.Y(n_1257)
);

INVx1_ASAP7_75t_L g1258 ( 
.A(n_1027),
.Y(n_1258)
);

INVx1_ASAP7_75t_L g1259 ( 
.A(n_1027),
.Y(n_1259)
);

INVx2_ASAP7_75t_SL g1260 ( 
.A(n_1032),
.Y(n_1260)
);

INVx3_ASAP7_75t_L g1261 ( 
.A(n_1009),
.Y(n_1261)
);

A2O1A1Ixp33_ASAP7_75t_L g1262 ( 
.A1(n_1153),
.A2(n_838),
.B(n_1147),
.C(n_1100),
.Y(n_1262)
);

AOI21xp5_ASAP7_75t_L g1263 ( 
.A1(n_1146),
.A2(n_1151),
.B(n_838),
.Y(n_1263)
);

OAI21x1_ASAP7_75t_L g1264 ( 
.A1(n_1132),
.A2(n_1008),
.B(n_1094),
.Y(n_1264)
);

AOI21xp5_ASAP7_75t_L g1265 ( 
.A1(n_1146),
.A2(n_1151),
.B(n_838),
.Y(n_1265)
);

AOI21xp5_ASAP7_75t_L g1266 ( 
.A1(n_1146),
.A2(n_1151),
.B(n_838),
.Y(n_1266)
);

AO31x2_ASAP7_75t_L g1267 ( 
.A1(n_1131),
.A2(n_1109),
.A3(n_1110),
.B(n_1069),
.Y(n_1267)
);

BUFx4f_ASAP7_75t_L g1268 ( 
.A(n_1009),
.Y(n_1268)
);

AOI21xp5_ASAP7_75t_L g1269 ( 
.A1(n_1146),
.A2(n_1151),
.B(n_838),
.Y(n_1269)
);

BUFx2_ASAP7_75t_L g1270 ( 
.A(n_1041),
.Y(n_1270)
);

INVx1_ASAP7_75t_L g1271 ( 
.A(n_1027),
.Y(n_1271)
);

O2A1O1Ixp33_ASAP7_75t_L g1272 ( 
.A1(n_1065),
.A2(n_1066),
.B(n_1147),
.C(n_1151),
.Y(n_1272)
);

AOI21xp5_ASAP7_75t_L g1273 ( 
.A1(n_1146),
.A2(n_1151),
.B(n_838),
.Y(n_1273)
);

OR2x2_ASAP7_75t_L g1274 ( 
.A(n_1147),
.B(n_701),
.Y(n_1274)
);

AOI22xp5_ASAP7_75t_L g1275 ( 
.A1(n_1147),
.A2(n_685),
.B1(n_695),
.B2(n_592),
.Y(n_1275)
);

CKINVDCx20_ASAP7_75t_R g1276 ( 
.A(n_1039),
.Y(n_1276)
);

AND2x4_ASAP7_75t_L g1277 ( 
.A(n_1036),
.B(n_992),
.Y(n_1277)
);

OAI21x1_ASAP7_75t_L g1278 ( 
.A1(n_1132),
.A2(n_1008),
.B(n_1094),
.Y(n_1278)
);

OAI21x1_ASAP7_75t_L g1279 ( 
.A1(n_1132),
.A2(n_1008),
.B(n_1094),
.Y(n_1279)
);

INVx1_ASAP7_75t_L g1280 ( 
.A(n_1027),
.Y(n_1280)
);

AOI21xp5_ASAP7_75t_L g1281 ( 
.A1(n_1146),
.A2(n_1151),
.B(n_838),
.Y(n_1281)
);

INVxp33_ASAP7_75t_L g1282 ( 
.A(n_1140),
.Y(n_1282)
);

O2A1O1Ixp33_ASAP7_75t_L g1283 ( 
.A1(n_1065),
.A2(n_1066),
.B(n_1147),
.C(n_1151),
.Y(n_1283)
);

NOR2xp67_ASAP7_75t_L g1284 ( 
.A(n_1056),
.B(n_661),
.Y(n_1284)
);

OAI21xp5_ASAP7_75t_L g1285 ( 
.A1(n_1151),
.A2(n_838),
.B(n_1138),
.Y(n_1285)
);

NAND2xp5_ASAP7_75t_L g1286 ( 
.A(n_1150),
.B(n_838),
.Y(n_1286)
);

A2O1A1Ixp33_ASAP7_75t_L g1287 ( 
.A1(n_1153),
.A2(n_838),
.B(n_1147),
.C(n_1100),
.Y(n_1287)
);

AND2x2_ASAP7_75t_L g1288 ( 
.A(n_1147),
.B(n_517),
.Y(n_1288)
);

INVx2_ASAP7_75t_L g1289 ( 
.A(n_1017),
.Y(n_1289)
);

HB1xp67_ASAP7_75t_L g1290 ( 
.A(n_1143),
.Y(n_1290)
);

OAI21xp5_ASAP7_75t_L g1291 ( 
.A1(n_1151),
.A2(n_838),
.B(n_1138),
.Y(n_1291)
);

NAND2x1p5_ASAP7_75t_L g1292 ( 
.A(n_1078),
.B(n_992),
.Y(n_1292)
);

AOI21xp5_ASAP7_75t_L g1293 ( 
.A1(n_1146),
.A2(n_1151),
.B(n_838),
.Y(n_1293)
);

AND2x4_ASAP7_75t_L g1294 ( 
.A(n_1036),
.B(n_992),
.Y(n_1294)
);

AOI21xp5_ASAP7_75t_SL g1295 ( 
.A1(n_1151),
.A2(n_872),
.B(n_1015),
.Y(n_1295)
);

INVx1_ASAP7_75t_L g1296 ( 
.A(n_1027),
.Y(n_1296)
);

A2O1A1Ixp33_ASAP7_75t_L g1297 ( 
.A1(n_1153),
.A2(n_838),
.B(n_1147),
.C(n_1100),
.Y(n_1297)
);

AO31x2_ASAP7_75t_L g1298 ( 
.A1(n_1131),
.A2(n_1109),
.A3(n_1110),
.B(n_1069),
.Y(n_1298)
);

O2A1O1Ixp33_ASAP7_75t_L g1299 ( 
.A1(n_1065),
.A2(n_1066),
.B(n_1147),
.C(n_1151),
.Y(n_1299)
);

INVx1_ASAP7_75t_L g1300 ( 
.A(n_1027),
.Y(n_1300)
);

NOR2xp33_ASAP7_75t_SL g1301 ( 
.A(n_1020),
.B(n_927),
.Y(n_1301)
);

BUFx2_ASAP7_75t_L g1302 ( 
.A(n_1041),
.Y(n_1302)
);

AOI21xp5_ASAP7_75t_L g1303 ( 
.A1(n_1146),
.A2(n_1151),
.B(n_838),
.Y(n_1303)
);

INVx1_ASAP7_75t_L g1304 ( 
.A(n_1027),
.Y(n_1304)
);

OAI21x1_ASAP7_75t_L g1305 ( 
.A1(n_1132),
.A2(n_1008),
.B(n_1094),
.Y(n_1305)
);

INVx2_ASAP7_75t_L g1306 ( 
.A(n_1017),
.Y(n_1306)
);

OAI21x1_ASAP7_75t_L g1307 ( 
.A1(n_1132),
.A2(n_1008),
.B(n_1094),
.Y(n_1307)
);

AND2x2_ASAP7_75t_L g1308 ( 
.A(n_1147),
.B(n_517),
.Y(n_1308)
);

OAI21xp5_ASAP7_75t_L g1309 ( 
.A1(n_1151),
.A2(n_838),
.B(n_1138),
.Y(n_1309)
);

OAI21xp5_ASAP7_75t_L g1310 ( 
.A1(n_1151),
.A2(n_838),
.B(n_1138),
.Y(n_1310)
);

AOI21x1_ASAP7_75t_L g1311 ( 
.A1(n_1085),
.A2(n_1074),
.B(n_1043),
.Y(n_1311)
);

AOI21xp5_ASAP7_75t_L g1312 ( 
.A1(n_1146),
.A2(n_1151),
.B(n_838),
.Y(n_1312)
);

A2O1A1Ixp33_ASAP7_75t_L g1313 ( 
.A1(n_1153),
.A2(n_838),
.B(n_1147),
.C(n_1100),
.Y(n_1313)
);

NAND2xp5_ASAP7_75t_L g1314 ( 
.A(n_1286),
.B(n_1170),
.Y(n_1314)
);

OAI22xp5_ASAP7_75t_L g1315 ( 
.A1(n_1262),
.A2(n_1313),
.B1(n_1287),
.B2(n_1297),
.Y(n_1315)
);

AOI22xp33_ASAP7_75t_L g1316 ( 
.A1(n_1301),
.A2(n_1173),
.B1(n_1178),
.B2(n_1165),
.Y(n_1316)
);

AOI22xp33_ASAP7_75t_SL g1317 ( 
.A1(n_1301),
.A2(n_1173),
.B1(n_1178),
.B2(n_1165),
.Y(n_1317)
);

CKINVDCx11_ASAP7_75t_R g1318 ( 
.A(n_1183),
.Y(n_1318)
);

AOI22xp33_ASAP7_75t_L g1319 ( 
.A1(n_1253),
.A2(n_1308),
.B1(n_1288),
.B2(n_1249),
.Y(n_1319)
);

BUFx8_ASAP7_75t_L g1320 ( 
.A(n_1187),
.Y(n_1320)
);

AOI22xp5_ASAP7_75t_L g1321 ( 
.A1(n_1162),
.A2(n_1275),
.B1(n_1193),
.B2(n_1274),
.Y(n_1321)
);

INVx2_ASAP7_75t_SL g1322 ( 
.A(n_1212),
.Y(n_1322)
);

INVx1_ASAP7_75t_L g1323 ( 
.A(n_1167),
.Y(n_1323)
);

CKINVDCx20_ASAP7_75t_R g1324 ( 
.A(n_1195),
.Y(n_1324)
);

AOI22xp33_ASAP7_75t_L g1325 ( 
.A1(n_1249),
.A2(n_1172),
.B1(n_1286),
.B2(n_1191),
.Y(n_1325)
);

INVx6_ASAP7_75t_L g1326 ( 
.A(n_1212),
.Y(n_1326)
);

AOI22xp33_ASAP7_75t_L g1327 ( 
.A1(n_1172),
.A2(n_1291),
.B1(n_1285),
.B2(n_1309),
.Y(n_1327)
);

AOI22xp33_ASAP7_75t_L g1328 ( 
.A1(n_1285),
.A2(n_1291),
.B1(n_1310),
.B2(n_1309),
.Y(n_1328)
);

AND2x2_ASAP7_75t_L g1329 ( 
.A(n_1161),
.B(n_1156),
.Y(n_1329)
);

INVx3_ASAP7_75t_L g1330 ( 
.A(n_1235),
.Y(n_1330)
);

AOI22xp33_ASAP7_75t_L g1331 ( 
.A1(n_1310),
.A2(n_1180),
.B1(n_1192),
.B2(n_1255),
.Y(n_1331)
);

BUFx12f_ASAP7_75t_L g1332 ( 
.A(n_1244),
.Y(n_1332)
);

OAI22xp33_ASAP7_75t_L g1333 ( 
.A1(n_1189),
.A2(n_1282),
.B1(n_1250),
.B2(n_1302),
.Y(n_1333)
);

CKINVDCx11_ASAP7_75t_R g1334 ( 
.A(n_1194),
.Y(n_1334)
);

HB1xp67_ASAP7_75t_L g1335 ( 
.A(n_1219),
.Y(n_1335)
);

INVx6_ASAP7_75t_L g1336 ( 
.A(n_1248),
.Y(n_1336)
);

INVx2_ASAP7_75t_L g1337 ( 
.A(n_1214),
.Y(n_1337)
);

INVx1_ASAP7_75t_L g1338 ( 
.A(n_1258),
.Y(n_1338)
);

AOI22xp33_ASAP7_75t_L g1339 ( 
.A1(n_1192),
.A2(n_1259),
.B1(n_1280),
.B2(n_1296),
.Y(n_1339)
);

AOI22xp33_ASAP7_75t_L g1340 ( 
.A1(n_1271),
.A2(n_1300),
.B1(n_1304),
.B2(n_1184),
.Y(n_1340)
);

INVx1_ASAP7_75t_L g1341 ( 
.A(n_1204),
.Y(n_1341)
);

CKINVDCx20_ASAP7_75t_R g1342 ( 
.A(n_1276),
.Y(n_1342)
);

AOI22xp33_ASAP7_75t_SL g1343 ( 
.A1(n_1211),
.A2(n_1177),
.B1(n_1207),
.B2(n_1209),
.Y(n_1343)
);

NAND2xp5_ASAP7_75t_L g1344 ( 
.A(n_1257),
.B(n_1272),
.Y(n_1344)
);

AOI22xp33_ASAP7_75t_SL g1345 ( 
.A1(n_1209),
.A2(n_1220),
.B1(n_1270),
.B2(n_1201),
.Y(n_1345)
);

INVx1_ASAP7_75t_L g1346 ( 
.A(n_1204),
.Y(n_1346)
);

INVx1_ASAP7_75t_L g1347 ( 
.A(n_1215),
.Y(n_1347)
);

AOI22xp33_ASAP7_75t_L g1348 ( 
.A1(n_1201),
.A2(n_1200),
.B1(n_1221),
.B2(n_1306),
.Y(n_1348)
);

BUFx12f_ASAP7_75t_L g1349 ( 
.A(n_1247),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_1159),
.Y(n_1350)
);

AOI22xp5_ASAP7_75t_L g1351 ( 
.A1(n_1157),
.A2(n_1284),
.B1(n_1171),
.B2(n_1246),
.Y(n_1351)
);

BUFx2_ASAP7_75t_L g1352 ( 
.A(n_1217),
.Y(n_1352)
);

BUFx2_ASAP7_75t_L g1353 ( 
.A(n_1230),
.Y(n_1353)
);

BUFx12f_ASAP7_75t_L g1354 ( 
.A(n_1250),
.Y(n_1354)
);

OAI22xp5_ASAP7_75t_L g1355 ( 
.A1(n_1283),
.A2(n_1299),
.B1(n_1164),
.B2(n_1196),
.Y(n_1355)
);

CKINVDCx16_ASAP7_75t_R g1356 ( 
.A(n_1250),
.Y(n_1356)
);

AOI22xp33_ASAP7_75t_L g1357 ( 
.A1(n_1289),
.A2(n_1290),
.B1(n_1277),
.B2(n_1294),
.Y(n_1357)
);

INVx1_ASAP7_75t_L g1358 ( 
.A(n_1227),
.Y(n_1358)
);

INVx1_ASAP7_75t_L g1359 ( 
.A(n_1225),
.Y(n_1359)
);

BUFx2_ASAP7_75t_L g1360 ( 
.A(n_1206),
.Y(n_1360)
);

CKINVDCx20_ASAP7_75t_R g1361 ( 
.A(n_1181),
.Y(n_1361)
);

INVx1_ASAP7_75t_L g1362 ( 
.A(n_1228),
.Y(n_1362)
);

AOI22xp33_ASAP7_75t_L g1363 ( 
.A1(n_1277),
.A2(n_1294),
.B1(n_1312),
.B2(n_1303),
.Y(n_1363)
);

INVx2_ASAP7_75t_SL g1364 ( 
.A(n_1268),
.Y(n_1364)
);

AOI22xp33_ASAP7_75t_L g1365 ( 
.A1(n_1242),
.A2(n_1256),
.B1(n_1254),
.B2(n_1252),
.Y(n_1365)
);

OAI21xp5_ASAP7_75t_SL g1366 ( 
.A1(n_1210),
.A2(n_1202),
.B(n_1273),
.Y(n_1366)
);

AOI22xp33_ASAP7_75t_L g1367 ( 
.A1(n_1243),
.A2(n_1269),
.B1(n_1265),
.B2(n_1293),
.Y(n_1367)
);

BUFx3_ASAP7_75t_L g1368 ( 
.A(n_1268),
.Y(n_1368)
);

OAI22xp5_ASAP7_75t_L g1369 ( 
.A1(n_1295),
.A2(n_1281),
.B1(n_1266),
.B2(n_1263),
.Y(n_1369)
);

BUFx12f_ASAP7_75t_L g1370 ( 
.A(n_1260),
.Y(n_1370)
);

INVx1_ASAP7_75t_L g1371 ( 
.A(n_1228),
.Y(n_1371)
);

INVx2_ASAP7_75t_L g1372 ( 
.A(n_1203),
.Y(n_1372)
);

NAND2xp5_ASAP7_75t_L g1373 ( 
.A(n_1182),
.B(n_1245),
.Y(n_1373)
);

NAND2xp5_ASAP7_75t_SL g1374 ( 
.A(n_1246),
.B(n_1233),
.Y(n_1374)
);

NAND2xp5_ASAP7_75t_L g1375 ( 
.A(n_1206),
.B(n_1248),
.Y(n_1375)
);

AOI22xp33_ASAP7_75t_L g1376 ( 
.A1(n_1166),
.A2(n_1205),
.B1(n_1155),
.B2(n_1154),
.Y(n_1376)
);

AOI22xp33_ASAP7_75t_L g1377 ( 
.A1(n_1166),
.A2(n_1233),
.B1(n_1218),
.B2(n_1229),
.Y(n_1377)
);

INVx1_ASAP7_75t_L g1378 ( 
.A(n_1226),
.Y(n_1378)
);

INVx1_ASAP7_75t_L g1379 ( 
.A(n_1222),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_1234),
.Y(n_1380)
);

BUFx12f_ASAP7_75t_L g1381 ( 
.A(n_1174),
.Y(n_1381)
);

INVx2_ASAP7_75t_L g1382 ( 
.A(n_1237),
.Y(n_1382)
);

CKINVDCx11_ASAP7_75t_R g1383 ( 
.A(n_1224),
.Y(n_1383)
);

INVx1_ASAP7_75t_L g1384 ( 
.A(n_1234),
.Y(n_1384)
);

INVx6_ASAP7_75t_L g1385 ( 
.A(n_1174),
.Y(n_1385)
);

NAND2xp5_ASAP7_75t_L g1386 ( 
.A(n_1163),
.B(n_1261),
.Y(n_1386)
);

INVx1_ASAP7_75t_L g1387 ( 
.A(n_1236),
.Y(n_1387)
);

NAND2x1p5_ASAP7_75t_L g1388 ( 
.A(n_1188),
.B(n_1169),
.Y(n_1388)
);

CKINVDCx5p33_ASAP7_75t_R g1389 ( 
.A(n_1231),
.Y(n_1389)
);

NAND2x1p5_ASAP7_75t_L g1390 ( 
.A(n_1223),
.B(n_1238),
.Y(n_1390)
);

AOI22xp33_ASAP7_75t_SL g1391 ( 
.A1(n_1292),
.A2(n_1176),
.B1(n_1158),
.B2(n_1168),
.Y(n_1391)
);

INVx4_ASAP7_75t_L g1392 ( 
.A(n_1223),
.Y(n_1392)
);

INVx1_ASAP7_75t_SL g1393 ( 
.A(n_1241),
.Y(n_1393)
);

INVx3_ASAP7_75t_L g1394 ( 
.A(n_1239),
.Y(n_1394)
);

OAI22xp5_ASAP7_75t_L g1395 ( 
.A1(n_1186),
.A2(n_1199),
.B1(n_1311),
.B2(n_1179),
.Y(n_1395)
);

OAI22xp33_ASAP7_75t_L g1396 ( 
.A1(n_1160),
.A2(n_1232),
.B1(n_1175),
.B2(n_1241),
.Y(n_1396)
);

CKINVDCx11_ASAP7_75t_R g1397 ( 
.A(n_1190),
.Y(n_1397)
);

AOI22xp33_ASAP7_75t_SL g1398 ( 
.A1(n_1185),
.A2(n_1190),
.B1(n_1307),
.B2(n_1264),
.Y(n_1398)
);

AOI22xp33_ASAP7_75t_L g1399 ( 
.A1(n_1190),
.A2(n_1213),
.B1(n_1197),
.B2(n_1305),
.Y(n_1399)
);

BUFx12f_ASAP7_75t_L g1400 ( 
.A(n_1208),
.Y(n_1400)
);

CKINVDCx20_ASAP7_75t_R g1401 ( 
.A(n_1240),
.Y(n_1401)
);

BUFx4f_ASAP7_75t_L g1402 ( 
.A(n_1267),
.Y(n_1402)
);

BUFx6f_ASAP7_75t_L g1403 ( 
.A(n_1251),
.Y(n_1403)
);

BUFx12f_ASAP7_75t_L g1404 ( 
.A(n_1267),
.Y(n_1404)
);

BUFx2_ASAP7_75t_L g1405 ( 
.A(n_1298),
.Y(n_1405)
);

NAND2x1p5_ASAP7_75t_L g1406 ( 
.A(n_1278),
.B(n_1279),
.Y(n_1406)
);

BUFx12f_ASAP7_75t_L g1407 ( 
.A(n_1198),
.Y(n_1407)
);

BUFx3_ASAP7_75t_L g1408 ( 
.A(n_1198),
.Y(n_1408)
);

HB1xp67_ASAP7_75t_L g1409 ( 
.A(n_1198),
.Y(n_1409)
);

INVx2_ASAP7_75t_L g1410 ( 
.A(n_1216),
.Y(n_1410)
);

AOI22xp33_ASAP7_75t_L g1411 ( 
.A1(n_1301),
.A2(n_1062),
.B1(n_1148),
.B2(n_927),
.Y(n_1411)
);

BUFx2_ASAP7_75t_SL g1412 ( 
.A(n_1195),
.Y(n_1412)
);

CKINVDCx20_ASAP7_75t_R g1413 ( 
.A(n_1183),
.Y(n_1413)
);

CKINVDCx5p33_ASAP7_75t_R g1414 ( 
.A(n_1183),
.Y(n_1414)
);

OAI22xp5_ASAP7_75t_L g1415 ( 
.A1(n_1262),
.A2(n_838),
.B1(n_1313),
.B2(n_1297),
.Y(n_1415)
);

CKINVDCx5p33_ASAP7_75t_R g1416 ( 
.A(n_1183),
.Y(n_1416)
);

INVx1_ASAP7_75t_L g1417 ( 
.A(n_1167),
.Y(n_1417)
);

AOI22xp33_ASAP7_75t_L g1418 ( 
.A1(n_1301),
.A2(n_1062),
.B1(n_1148),
.B2(n_927),
.Y(n_1418)
);

AND2x2_ASAP7_75t_L g1419 ( 
.A(n_1253),
.B(n_1288),
.Y(n_1419)
);

BUFx6f_ASAP7_75t_L g1420 ( 
.A(n_1277),
.Y(n_1420)
);

NAND2xp5_ASAP7_75t_L g1421 ( 
.A(n_1286),
.B(n_1170),
.Y(n_1421)
);

BUFx12f_ASAP7_75t_L g1422 ( 
.A(n_1183),
.Y(n_1422)
);

AOI22xp33_ASAP7_75t_L g1423 ( 
.A1(n_1301),
.A2(n_1062),
.B1(n_1148),
.B2(n_927),
.Y(n_1423)
);

OAI22xp5_ASAP7_75t_L g1424 ( 
.A1(n_1262),
.A2(n_838),
.B1(n_1313),
.B2(n_1297),
.Y(n_1424)
);

OAI22xp33_ASAP7_75t_L g1425 ( 
.A1(n_1301),
.A2(n_1020),
.B1(n_1073),
.B2(n_1275),
.Y(n_1425)
);

CKINVDCx11_ASAP7_75t_R g1426 ( 
.A(n_1183),
.Y(n_1426)
);

BUFx4f_ASAP7_75t_SL g1427 ( 
.A(n_1187),
.Y(n_1427)
);

OAI22xp5_ASAP7_75t_L g1428 ( 
.A1(n_1262),
.A2(n_838),
.B1(n_1313),
.B2(n_1297),
.Y(n_1428)
);

INVx1_ASAP7_75t_L g1429 ( 
.A(n_1167),
.Y(n_1429)
);

INVx1_ASAP7_75t_L g1430 ( 
.A(n_1167),
.Y(n_1430)
);

BUFx2_ASAP7_75t_L g1431 ( 
.A(n_1270),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_1167),
.Y(n_1432)
);

CKINVDCx11_ASAP7_75t_R g1433 ( 
.A(n_1183),
.Y(n_1433)
);

OAI22xp33_ASAP7_75t_L g1434 ( 
.A1(n_1301),
.A2(n_1020),
.B1(n_1073),
.B2(n_1275),
.Y(n_1434)
);

INVx1_ASAP7_75t_L g1435 ( 
.A(n_1167),
.Y(n_1435)
);

NAND2xp5_ASAP7_75t_L g1436 ( 
.A(n_1286),
.B(n_1170),
.Y(n_1436)
);

OAI21xp5_ASAP7_75t_SL g1437 ( 
.A1(n_1275),
.A2(n_1157),
.B(n_1257),
.Y(n_1437)
);

NAND2xp5_ASAP7_75t_L g1438 ( 
.A(n_1286),
.B(n_1170),
.Y(n_1438)
);

INVx1_ASAP7_75t_L g1439 ( 
.A(n_1167),
.Y(n_1439)
);

AOI22xp33_ASAP7_75t_L g1440 ( 
.A1(n_1301),
.A2(n_1062),
.B1(n_1148),
.B2(n_927),
.Y(n_1440)
);

AOI22xp33_ASAP7_75t_L g1441 ( 
.A1(n_1301),
.A2(n_1062),
.B1(n_1148),
.B2(n_927),
.Y(n_1441)
);

OAI22xp33_ASAP7_75t_L g1442 ( 
.A1(n_1301),
.A2(n_1020),
.B1(n_1073),
.B2(n_1275),
.Y(n_1442)
);

INVx1_ASAP7_75t_SL g1443 ( 
.A(n_1156),
.Y(n_1443)
);

INVx1_ASAP7_75t_L g1444 ( 
.A(n_1167),
.Y(n_1444)
);

INVx2_ASAP7_75t_L g1445 ( 
.A(n_1216),
.Y(n_1445)
);

INVx2_ASAP7_75t_L g1446 ( 
.A(n_1216),
.Y(n_1446)
);

BUFx3_ASAP7_75t_L g1447 ( 
.A(n_1353),
.Y(n_1447)
);

INVx1_ASAP7_75t_L g1448 ( 
.A(n_1409),
.Y(n_1448)
);

INVx1_ASAP7_75t_L g1449 ( 
.A(n_1405),
.Y(n_1449)
);

NAND2xp5_ASAP7_75t_L g1450 ( 
.A(n_1325),
.B(n_1327),
.Y(n_1450)
);

OAI21x1_ASAP7_75t_L g1451 ( 
.A1(n_1406),
.A2(n_1395),
.B(n_1369),
.Y(n_1451)
);

AOI222xp33_ASAP7_75t_L g1452 ( 
.A1(n_1316),
.A2(n_1437),
.B1(n_1319),
.B2(n_1442),
.C1(n_1434),
.C2(n_1425),
.Y(n_1452)
);

NAND2x1p5_ASAP7_75t_L g1453 ( 
.A(n_1380),
.B(n_1384),
.Y(n_1453)
);

BUFx2_ASAP7_75t_L g1454 ( 
.A(n_1407),
.Y(n_1454)
);

BUFx3_ASAP7_75t_L g1455 ( 
.A(n_1431),
.Y(n_1455)
);

INVx2_ASAP7_75t_SL g1456 ( 
.A(n_1335),
.Y(n_1456)
);

BUFx6f_ASAP7_75t_L g1457 ( 
.A(n_1400),
.Y(n_1457)
);

AND2x4_ASAP7_75t_L g1458 ( 
.A(n_1408),
.B(n_1387),
.Y(n_1458)
);

INVx1_ASAP7_75t_L g1459 ( 
.A(n_1323),
.Y(n_1459)
);

OAI21x1_ASAP7_75t_L g1460 ( 
.A1(n_1406),
.A2(n_1367),
.B(n_1365),
.Y(n_1460)
);

HB1xp67_ASAP7_75t_L g1461 ( 
.A(n_1359),
.Y(n_1461)
);

BUFx2_ASAP7_75t_L g1462 ( 
.A(n_1407),
.Y(n_1462)
);

INVx1_ASAP7_75t_L g1463 ( 
.A(n_1338),
.Y(n_1463)
);

AO21x2_ASAP7_75t_L g1464 ( 
.A1(n_1396),
.A2(n_1382),
.B(n_1372),
.Y(n_1464)
);

AOI221xp5_ASAP7_75t_L g1465 ( 
.A1(n_1316),
.A2(n_1355),
.B1(n_1424),
.B2(n_1415),
.C(n_1428),
.Y(n_1465)
);

INVx1_ASAP7_75t_L g1466 ( 
.A(n_1417),
.Y(n_1466)
);

AND2x4_ASAP7_75t_L g1467 ( 
.A(n_1408),
.B(n_1401),
.Y(n_1467)
);

AND2x2_ASAP7_75t_L g1468 ( 
.A(n_1328),
.B(n_1429),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_1430),
.Y(n_1469)
);

AND2x2_ASAP7_75t_L g1470 ( 
.A(n_1328),
.B(n_1432),
.Y(n_1470)
);

AO21x1_ASAP7_75t_L g1471 ( 
.A1(n_1315),
.A2(n_1366),
.B(n_1344),
.Y(n_1471)
);

INVx1_ASAP7_75t_L g1472 ( 
.A(n_1435),
.Y(n_1472)
);

HB1xp67_ASAP7_75t_L g1473 ( 
.A(n_1358),
.Y(n_1473)
);

INVx1_ASAP7_75t_L g1474 ( 
.A(n_1439),
.Y(n_1474)
);

INVx1_ASAP7_75t_L g1475 ( 
.A(n_1444),
.Y(n_1475)
);

INVx1_ASAP7_75t_SL g1476 ( 
.A(n_1352),
.Y(n_1476)
);

INVx1_ASAP7_75t_L g1477 ( 
.A(n_1337),
.Y(n_1477)
);

OAI21x1_ASAP7_75t_L g1478 ( 
.A1(n_1365),
.A2(n_1367),
.B(n_1399),
.Y(n_1478)
);

OA21x2_ASAP7_75t_L g1479 ( 
.A1(n_1376),
.A2(n_1399),
.B(n_1382),
.Y(n_1479)
);

INVx1_ASAP7_75t_L g1480 ( 
.A(n_1374),
.Y(n_1480)
);

OAI21x1_ASAP7_75t_L g1481 ( 
.A1(n_1376),
.A2(n_1394),
.B(n_1390),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_1374),
.Y(n_1482)
);

INVx1_ASAP7_75t_L g1483 ( 
.A(n_1341),
.Y(n_1483)
);

HB1xp67_ASAP7_75t_L g1484 ( 
.A(n_1373),
.Y(n_1484)
);

INVx1_ASAP7_75t_L g1485 ( 
.A(n_1346),
.Y(n_1485)
);

AOI22xp33_ASAP7_75t_L g1486 ( 
.A1(n_1411),
.A2(n_1418),
.B1(n_1423),
.B2(n_1440),
.Y(n_1486)
);

OA21x2_ASAP7_75t_L g1487 ( 
.A1(n_1327),
.A2(n_1393),
.B(n_1377),
.Y(n_1487)
);

INVx1_ASAP7_75t_L g1488 ( 
.A(n_1404),
.Y(n_1488)
);

INVx1_ASAP7_75t_L g1489 ( 
.A(n_1404),
.Y(n_1489)
);

INVx1_ASAP7_75t_L g1490 ( 
.A(n_1402),
.Y(n_1490)
);

OAI21xp5_ASAP7_75t_L g1491 ( 
.A1(n_1317),
.A2(n_1351),
.B(n_1391),
.Y(n_1491)
);

AO21x2_ASAP7_75t_L g1492 ( 
.A1(n_1379),
.A2(n_1362),
.B(n_1371),
.Y(n_1492)
);

BUFx3_ASAP7_75t_L g1493 ( 
.A(n_1390),
.Y(n_1493)
);

AND2x2_ASAP7_75t_L g1494 ( 
.A(n_1339),
.B(n_1377),
.Y(n_1494)
);

HB1xp67_ASAP7_75t_L g1495 ( 
.A(n_1329),
.Y(n_1495)
);

INVx1_ASAP7_75t_L g1496 ( 
.A(n_1339),
.Y(n_1496)
);

INVx1_ASAP7_75t_L g1497 ( 
.A(n_1410),
.Y(n_1497)
);

INVx5_ASAP7_75t_SL g1498 ( 
.A(n_1420),
.Y(n_1498)
);

CKINVDCx5p33_ASAP7_75t_R g1499 ( 
.A(n_1334),
.Y(n_1499)
);

AND2x2_ASAP7_75t_L g1500 ( 
.A(n_1419),
.B(n_1325),
.Y(n_1500)
);

HB1xp67_ASAP7_75t_L g1501 ( 
.A(n_1347),
.Y(n_1501)
);

AOI22xp33_ASAP7_75t_L g1502 ( 
.A1(n_1411),
.A2(n_1441),
.B1(n_1423),
.B2(n_1418),
.Y(n_1502)
);

INVx1_ASAP7_75t_SL g1503 ( 
.A(n_1443),
.Y(n_1503)
);

HB1xp67_ASAP7_75t_L g1504 ( 
.A(n_1314),
.Y(n_1504)
);

AND2x4_ASAP7_75t_L g1505 ( 
.A(n_1363),
.B(n_1445),
.Y(n_1505)
);

OA21x2_ASAP7_75t_L g1506 ( 
.A1(n_1331),
.A2(n_1363),
.B(n_1378),
.Y(n_1506)
);

INVx2_ASAP7_75t_L g1507 ( 
.A(n_1446),
.Y(n_1507)
);

HB1xp67_ASAP7_75t_L g1508 ( 
.A(n_1421),
.Y(n_1508)
);

BUFx2_ASAP7_75t_L g1509 ( 
.A(n_1403),
.Y(n_1509)
);

OAI22xp5_ASAP7_75t_L g1510 ( 
.A1(n_1319),
.A2(n_1441),
.B1(n_1440),
.B2(n_1331),
.Y(n_1510)
);

INVx3_ASAP7_75t_L g1511 ( 
.A(n_1403),
.Y(n_1511)
);

OA21x2_ASAP7_75t_L g1512 ( 
.A1(n_1340),
.A2(n_1348),
.B(n_1350),
.Y(n_1512)
);

NAND2xp5_ASAP7_75t_L g1513 ( 
.A(n_1340),
.B(n_1438),
.Y(n_1513)
);

AND2x2_ASAP7_75t_L g1514 ( 
.A(n_1436),
.B(n_1397),
.Y(n_1514)
);

OA21x2_ASAP7_75t_L g1515 ( 
.A1(n_1348),
.A2(n_1357),
.B(n_1398),
.Y(n_1515)
);

OR2x2_ASAP7_75t_L g1516 ( 
.A(n_1321),
.B(n_1333),
.Y(n_1516)
);

INVx3_ASAP7_75t_L g1517 ( 
.A(n_1392),
.Y(n_1517)
);

NAND2xp5_ASAP7_75t_L g1518 ( 
.A(n_1345),
.B(n_1343),
.Y(n_1518)
);

HB1xp67_ASAP7_75t_L g1519 ( 
.A(n_1330),
.Y(n_1519)
);

INVx1_ASAP7_75t_L g1520 ( 
.A(n_1386),
.Y(n_1520)
);

INVx1_ASAP7_75t_L g1521 ( 
.A(n_1392),
.Y(n_1521)
);

OA21x2_ASAP7_75t_L g1522 ( 
.A1(n_1357),
.A2(n_1375),
.B(n_1360),
.Y(n_1522)
);

AND2x2_ASAP7_75t_L g1523 ( 
.A(n_1330),
.B(n_1356),
.Y(n_1523)
);

AOI21x1_ASAP7_75t_L g1524 ( 
.A1(n_1364),
.A2(n_1336),
.B(n_1322),
.Y(n_1524)
);

AOI21xp5_ASAP7_75t_L g1525 ( 
.A1(n_1388),
.A2(n_1368),
.B(n_1389),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_1388),
.Y(n_1526)
);

INVx1_ASAP7_75t_L g1527 ( 
.A(n_1385),
.Y(n_1527)
);

O2A1O1Ixp33_ASAP7_75t_L g1528 ( 
.A1(n_1368),
.A2(n_1361),
.B(n_1342),
.C(n_1324),
.Y(n_1528)
);

AOI22xp5_ASAP7_75t_L g1529 ( 
.A1(n_1452),
.A2(n_1383),
.B1(n_1370),
.B2(n_1326),
.Y(n_1529)
);

OAI22xp5_ASAP7_75t_L g1530 ( 
.A1(n_1465),
.A2(n_1326),
.B1(n_1354),
.B2(n_1413),
.Y(n_1530)
);

OAI22xp5_ASAP7_75t_L g1531 ( 
.A1(n_1465),
.A2(n_1326),
.B1(n_1354),
.B2(n_1422),
.Y(n_1531)
);

AND2x2_ASAP7_75t_L g1532 ( 
.A(n_1455),
.B(n_1412),
.Y(n_1532)
);

AND2x4_ASAP7_75t_L g1533 ( 
.A(n_1447),
.B(n_1414),
.Y(n_1533)
);

OAI21xp5_ASAP7_75t_L g1534 ( 
.A1(n_1491),
.A2(n_1416),
.B(n_1383),
.Y(n_1534)
);

AND2x2_ASAP7_75t_L g1535 ( 
.A(n_1455),
.B(n_1495),
.Y(n_1535)
);

AND2x2_ASAP7_75t_L g1536 ( 
.A(n_1455),
.B(n_1370),
.Y(n_1536)
);

AND2x2_ASAP7_75t_L g1537 ( 
.A(n_1514),
.B(n_1422),
.Y(n_1537)
);

INVx1_ASAP7_75t_L g1538 ( 
.A(n_1473),
.Y(n_1538)
);

AND2x2_ASAP7_75t_L g1539 ( 
.A(n_1514),
.B(n_1349),
.Y(n_1539)
);

AND2x2_ASAP7_75t_L g1540 ( 
.A(n_1523),
.B(n_1349),
.Y(n_1540)
);

AND2x2_ASAP7_75t_L g1541 ( 
.A(n_1523),
.B(n_1456),
.Y(n_1541)
);

NAND3xp33_ASAP7_75t_L g1542 ( 
.A(n_1452),
.B(n_1320),
.C(n_1318),
.Y(n_1542)
);

NAND2xp5_ASAP7_75t_L g1543 ( 
.A(n_1480),
.B(n_1381),
.Y(n_1543)
);

OAI22xp5_ASAP7_75t_L g1544 ( 
.A1(n_1450),
.A2(n_1427),
.B1(n_1332),
.B2(n_1381),
.Y(n_1544)
);

NOR2xp33_ASAP7_75t_L g1545 ( 
.A(n_1499),
.B(n_1528),
.Y(n_1545)
);

A2O1A1Ixp33_ASAP7_75t_L g1546 ( 
.A1(n_1491),
.A2(n_1318),
.B(n_1320),
.C(n_1426),
.Y(n_1546)
);

AOI22xp33_ASAP7_75t_L g1547 ( 
.A1(n_1486),
.A2(n_1433),
.B1(n_1332),
.B2(n_1320),
.Y(n_1547)
);

INVxp67_ASAP7_75t_L g1548 ( 
.A(n_1519),
.Y(n_1548)
);

A2O1A1Ixp33_ASAP7_75t_L g1549 ( 
.A1(n_1510),
.A2(n_1502),
.B(n_1450),
.C(n_1518),
.Y(n_1549)
);

OAI21xp5_ASAP7_75t_L g1550 ( 
.A1(n_1510),
.A2(n_1494),
.B(n_1496),
.Y(n_1550)
);

AND2x4_ASAP7_75t_L g1551 ( 
.A(n_1447),
.B(n_1456),
.Y(n_1551)
);

AOI22xp5_ASAP7_75t_L g1552 ( 
.A1(n_1471),
.A2(n_1494),
.B1(n_1518),
.B2(n_1516),
.Y(n_1552)
);

NOR2xp33_ASAP7_75t_L g1553 ( 
.A(n_1476),
.B(n_1471),
.Y(n_1553)
);

O2A1O1Ixp33_ASAP7_75t_SL g1554 ( 
.A1(n_1461),
.A2(n_1476),
.B(n_1516),
.C(n_1525),
.Y(n_1554)
);

O2A1O1Ixp33_ASAP7_75t_L g1555 ( 
.A1(n_1484),
.A2(n_1496),
.B(n_1480),
.C(n_1482),
.Y(n_1555)
);

INVx1_ASAP7_75t_L g1556 ( 
.A(n_1501),
.Y(n_1556)
);

AND2x4_ASAP7_75t_L g1557 ( 
.A(n_1447),
.B(n_1488),
.Y(n_1557)
);

OR2x2_ASAP7_75t_L g1558 ( 
.A(n_1500),
.B(n_1504),
.Y(n_1558)
);

NAND2xp5_ASAP7_75t_L g1559 ( 
.A(n_1482),
.B(n_1468),
.Y(n_1559)
);

OA21x2_ASAP7_75t_L g1560 ( 
.A1(n_1451),
.A2(n_1478),
.B(n_1460),
.Y(n_1560)
);

OA21x2_ASAP7_75t_L g1561 ( 
.A1(n_1478),
.A2(n_1460),
.B(n_1481),
.Y(n_1561)
);

OR2x2_ASAP7_75t_L g1562 ( 
.A(n_1500),
.B(n_1508),
.Y(n_1562)
);

AND2x2_ASAP7_75t_L g1563 ( 
.A(n_1468),
.B(n_1470),
.Y(n_1563)
);

OAI21xp5_ASAP7_75t_L g1564 ( 
.A1(n_1506),
.A2(n_1487),
.B(n_1470),
.Y(n_1564)
);

INVx1_ASAP7_75t_L g1565 ( 
.A(n_1459),
.Y(n_1565)
);

AND2x2_ASAP7_75t_L g1566 ( 
.A(n_1453),
.B(n_1467),
.Y(n_1566)
);

CKINVDCx5p33_ASAP7_75t_R g1567 ( 
.A(n_1503),
.Y(n_1567)
);

OAI22xp5_ASAP7_75t_L g1568 ( 
.A1(n_1513),
.A2(n_1506),
.B1(n_1487),
.B2(n_1457),
.Y(n_1568)
);

OAI211xp5_ASAP7_75t_L g1569 ( 
.A1(n_1506),
.A2(n_1487),
.B(n_1513),
.C(n_1479),
.Y(n_1569)
);

OAI21x1_ASAP7_75t_SL g1570 ( 
.A1(n_1524),
.A2(n_1521),
.B(n_1472),
.Y(n_1570)
);

O2A1O1Ixp33_ASAP7_75t_L g1571 ( 
.A1(n_1506),
.A2(n_1503),
.B(n_1520),
.C(n_1526),
.Y(n_1571)
);

NAND2xp5_ASAP7_75t_L g1572 ( 
.A(n_1483),
.B(n_1485),
.Y(n_1572)
);

AND2x4_ASAP7_75t_L g1573 ( 
.A(n_1488),
.B(n_1489),
.Y(n_1573)
);

AND2x2_ASAP7_75t_L g1574 ( 
.A(n_1463),
.B(n_1466),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_1463),
.Y(n_1575)
);

AOI211xp5_ASAP7_75t_L g1576 ( 
.A1(n_1505),
.A2(n_1457),
.B(n_1474),
.C(n_1475),
.Y(n_1576)
);

OR2x6_ASAP7_75t_L g1577 ( 
.A(n_1505),
.B(n_1454),
.Y(n_1577)
);

A2O1A1Ixp33_ASAP7_75t_L g1578 ( 
.A1(n_1505),
.A2(n_1489),
.B(n_1462),
.C(n_1454),
.Y(n_1578)
);

BUFx2_ASAP7_75t_L g1579 ( 
.A(n_1527),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_1469),
.Y(n_1580)
);

A2O1A1Ixp33_ASAP7_75t_L g1581 ( 
.A1(n_1462),
.A2(n_1490),
.B(n_1458),
.C(n_1493),
.Y(n_1581)
);

AO32x2_ASAP7_75t_L g1582 ( 
.A1(n_1512),
.A2(n_1492),
.A3(n_1522),
.B1(n_1515),
.B2(n_1507),
.Y(n_1582)
);

AO32x2_ASAP7_75t_L g1583 ( 
.A1(n_1512),
.A2(n_1492),
.A3(n_1522),
.B1(n_1515),
.B2(n_1507),
.Y(n_1583)
);

AND2x6_ASAP7_75t_L g1584 ( 
.A(n_1498),
.B(n_1493),
.Y(n_1584)
);

INVx1_ASAP7_75t_L g1585 ( 
.A(n_1565),
.Y(n_1585)
);

NAND2xp5_ASAP7_75t_L g1586 ( 
.A(n_1559),
.B(n_1492),
.Y(n_1586)
);

INVx2_ASAP7_75t_L g1587 ( 
.A(n_1582),
.Y(n_1587)
);

INVx2_ASAP7_75t_L g1588 ( 
.A(n_1582),
.Y(n_1588)
);

AND2x2_ASAP7_75t_L g1589 ( 
.A(n_1563),
.B(n_1479),
.Y(n_1589)
);

AND2x2_ASAP7_75t_L g1590 ( 
.A(n_1559),
.B(n_1479),
.Y(n_1590)
);

INVx2_ASAP7_75t_L g1591 ( 
.A(n_1582),
.Y(n_1591)
);

NAND2xp5_ASAP7_75t_L g1592 ( 
.A(n_1553),
.B(n_1574),
.Y(n_1592)
);

AND2x2_ASAP7_75t_L g1593 ( 
.A(n_1560),
.B(n_1479),
.Y(n_1593)
);

INVx2_ASAP7_75t_L g1594 ( 
.A(n_1583),
.Y(n_1594)
);

INVx1_ASAP7_75t_L g1595 ( 
.A(n_1575),
.Y(n_1595)
);

OR2x2_ASAP7_75t_L g1596 ( 
.A(n_1558),
.B(n_1562),
.Y(n_1596)
);

OR2x2_ASAP7_75t_L g1597 ( 
.A(n_1538),
.B(n_1464),
.Y(n_1597)
);

INVx2_ASAP7_75t_L g1598 ( 
.A(n_1583),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1580),
.Y(n_1599)
);

INVx2_ASAP7_75t_L g1600 ( 
.A(n_1583),
.Y(n_1600)
);

INVx2_ASAP7_75t_L g1601 ( 
.A(n_1561),
.Y(n_1601)
);

INVx8_ASAP7_75t_L g1602 ( 
.A(n_1584),
.Y(n_1602)
);

AND2x4_ASAP7_75t_SL g1603 ( 
.A(n_1577),
.B(n_1458),
.Y(n_1603)
);

AND2x4_ASAP7_75t_L g1604 ( 
.A(n_1577),
.B(n_1511),
.Y(n_1604)
);

INVx1_ASAP7_75t_L g1605 ( 
.A(n_1572),
.Y(n_1605)
);

INVx1_ASAP7_75t_L g1606 ( 
.A(n_1572),
.Y(n_1606)
);

INVx2_ASAP7_75t_SL g1607 ( 
.A(n_1551),
.Y(n_1607)
);

INVx2_ASAP7_75t_SL g1608 ( 
.A(n_1551),
.Y(n_1608)
);

OAI22xp5_ASAP7_75t_L g1609 ( 
.A1(n_1552),
.A2(n_1515),
.B1(n_1526),
.B2(n_1517),
.Y(n_1609)
);

INVx2_ASAP7_75t_SL g1610 ( 
.A(n_1557),
.Y(n_1610)
);

AND2x2_ASAP7_75t_L g1611 ( 
.A(n_1535),
.B(n_1464),
.Y(n_1611)
);

INVx1_ASAP7_75t_L g1612 ( 
.A(n_1556),
.Y(n_1612)
);

OR2x2_ASAP7_75t_L g1613 ( 
.A(n_1548),
.B(n_1448),
.Y(n_1613)
);

OR2x2_ASAP7_75t_L g1614 ( 
.A(n_1564),
.B(n_1449),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_1570),
.Y(n_1615)
);

OR2x2_ASAP7_75t_L g1616 ( 
.A(n_1564),
.B(n_1509),
.Y(n_1616)
);

AND2x2_ASAP7_75t_L g1617 ( 
.A(n_1541),
.B(n_1509),
.Y(n_1617)
);

BUFx3_ASAP7_75t_L g1618 ( 
.A(n_1612),
.Y(n_1618)
);

AND2x2_ASAP7_75t_L g1619 ( 
.A(n_1607),
.B(n_1608),
.Y(n_1619)
);

INVx1_ASAP7_75t_L g1620 ( 
.A(n_1585),
.Y(n_1620)
);

AND2x2_ASAP7_75t_L g1621 ( 
.A(n_1607),
.B(n_1532),
.Y(n_1621)
);

NAND2xp5_ASAP7_75t_L g1622 ( 
.A(n_1592),
.B(n_1605),
.Y(n_1622)
);

AND2x2_ASAP7_75t_L g1623 ( 
.A(n_1607),
.B(n_1579),
.Y(n_1623)
);

INVx1_ASAP7_75t_L g1624 ( 
.A(n_1585),
.Y(n_1624)
);

INVx1_ASAP7_75t_L g1625 ( 
.A(n_1585),
.Y(n_1625)
);

INVx1_ASAP7_75t_L g1626 ( 
.A(n_1595),
.Y(n_1626)
);

AND2x2_ASAP7_75t_L g1627 ( 
.A(n_1608),
.B(n_1566),
.Y(n_1627)
);

AOI221xp5_ASAP7_75t_L g1628 ( 
.A1(n_1609),
.A2(n_1549),
.B1(n_1550),
.B2(n_1555),
.C(n_1568),
.Y(n_1628)
);

AOI22xp33_ASAP7_75t_L g1629 ( 
.A1(n_1609),
.A2(n_1550),
.B1(n_1542),
.B2(n_1568),
.Y(n_1629)
);

INVx1_ASAP7_75t_L g1630 ( 
.A(n_1595),
.Y(n_1630)
);

INVx3_ASAP7_75t_L g1631 ( 
.A(n_1602),
.Y(n_1631)
);

INVxp67_ASAP7_75t_SL g1632 ( 
.A(n_1586),
.Y(n_1632)
);

INVxp67_ASAP7_75t_L g1633 ( 
.A(n_1592),
.Y(n_1633)
);

OR2x2_ASAP7_75t_L g1634 ( 
.A(n_1596),
.B(n_1569),
.Y(n_1634)
);

OR2x2_ASAP7_75t_L g1635 ( 
.A(n_1596),
.B(n_1569),
.Y(n_1635)
);

OAI33xp33_ASAP7_75t_L g1636 ( 
.A1(n_1586),
.A2(n_1542),
.A3(n_1530),
.B1(n_1531),
.B2(n_1544),
.B3(n_1543),
.Y(n_1636)
);

INVx2_ASAP7_75t_L g1637 ( 
.A(n_1601),
.Y(n_1637)
);

AOI21xp5_ASAP7_75t_L g1638 ( 
.A1(n_1602),
.A2(n_1554),
.B(n_1530),
.Y(n_1638)
);

INVx1_ASAP7_75t_L g1639 ( 
.A(n_1599),
.Y(n_1639)
);

NAND2xp5_ASAP7_75t_L g1640 ( 
.A(n_1605),
.B(n_1567),
.Y(n_1640)
);

BUFx6f_ASAP7_75t_L g1641 ( 
.A(n_1602),
.Y(n_1641)
);

AOI22xp5_ASAP7_75t_L g1642 ( 
.A1(n_1589),
.A2(n_1529),
.B1(n_1531),
.B2(n_1576),
.Y(n_1642)
);

AOI211xp5_ASAP7_75t_L g1643 ( 
.A1(n_1614),
.A2(n_1534),
.B(n_1546),
.C(n_1544),
.Y(n_1643)
);

HB1xp67_ASAP7_75t_L g1644 ( 
.A(n_1613),
.Y(n_1644)
);

OR2x6_ASAP7_75t_L g1645 ( 
.A(n_1602),
.B(n_1571),
.Y(n_1645)
);

AO21x2_ASAP7_75t_L g1646 ( 
.A1(n_1587),
.A2(n_1578),
.B(n_1477),
.Y(n_1646)
);

HB1xp67_ASAP7_75t_SL g1647 ( 
.A(n_1610),
.Y(n_1647)
);

BUFx6f_ASAP7_75t_SL g1648 ( 
.A(n_1604),
.Y(n_1648)
);

AOI222xp33_ASAP7_75t_L g1649 ( 
.A1(n_1590),
.A2(n_1534),
.B1(n_1547),
.B2(n_1537),
.C1(n_1573),
.C2(n_1497),
.Y(n_1649)
);

INVxp67_ASAP7_75t_L g1650 ( 
.A(n_1612),
.Y(n_1650)
);

OR2x6_ASAP7_75t_L g1651 ( 
.A(n_1602),
.B(n_1581),
.Y(n_1651)
);

AND2x2_ASAP7_75t_L g1652 ( 
.A(n_1589),
.B(n_1533),
.Y(n_1652)
);

INVxp67_ASAP7_75t_SL g1653 ( 
.A(n_1616),
.Y(n_1653)
);

INVx1_ASAP7_75t_L g1654 ( 
.A(n_1599),
.Y(n_1654)
);

NAND4xp25_ASAP7_75t_SL g1655 ( 
.A(n_1615),
.B(n_1539),
.C(n_1536),
.D(n_1540),
.Y(n_1655)
);

OR2x2_ASAP7_75t_L g1656 ( 
.A(n_1634),
.B(n_1597),
.Y(n_1656)
);

NAND2xp5_ASAP7_75t_L g1657 ( 
.A(n_1622),
.B(n_1644),
.Y(n_1657)
);

HB1xp67_ASAP7_75t_L g1658 ( 
.A(n_1634),
.Y(n_1658)
);

AND2x2_ASAP7_75t_L g1659 ( 
.A(n_1653),
.B(n_1589),
.Y(n_1659)
);

NOR2xp33_ASAP7_75t_L g1660 ( 
.A(n_1655),
.B(n_1545),
.Y(n_1660)
);

HB1xp67_ASAP7_75t_L g1661 ( 
.A(n_1635),
.Y(n_1661)
);

AND2x2_ASAP7_75t_L g1662 ( 
.A(n_1652),
.B(n_1611),
.Y(n_1662)
);

AOI22xp33_ASAP7_75t_L g1663 ( 
.A1(n_1628),
.A2(n_1629),
.B1(n_1636),
.B2(n_1635),
.Y(n_1663)
);

AND2x2_ASAP7_75t_L g1664 ( 
.A(n_1652),
.B(n_1611),
.Y(n_1664)
);

AND2x2_ASAP7_75t_L g1665 ( 
.A(n_1619),
.B(n_1611),
.Y(n_1665)
);

AND2x2_ASAP7_75t_L g1666 ( 
.A(n_1619),
.B(n_1617),
.Y(n_1666)
);

INVx1_ASAP7_75t_L g1667 ( 
.A(n_1620),
.Y(n_1667)
);

INVx1_ASAP7_75t_L g1668 ( 
.A(n_1624),
.Y(n_1668)
);

NOR2xp33_ASAP7_75t_L g1669 ( 
.A(n_1640),
.B(n_1610),
.Y(n_1669)
);

OAI22xp5_ASAP7_75t_L g1670 ( 
.A1(n_1643),
.A2(n_1642),
.B1(n_1638),
.B2(n_1647),
.Y(n_1670)
);

NAND2xp5_ASAP7_75t_L g1671 ( 
.A(n_1633),
.B(n_1606),
.Y(n_1671)
);

AND2x2_ASAP7_75t_L g1672 ( 
.A(n_1623),
.B(n_1617),
.Y(n_1672)
);

AND2x4_ASAP7_75t_L g1673 ( 
.A(n_1645),
.B(n_1603),
.Y(n_1673)
);

AND2x2_ASAP7_75t_SL g1674 ( 
.A(n_1641),
.B(n_1603),
.Y(n_1674)
);

INVx1_ASAP7_75t_L g1675 ( 
.A(n_1625),
.Y(n_1675)
);

OR2x2_ASAP7_75t_L g1676 ( 
.A(n_1632),
.B(n_1587),
.Y(n_1676)
);

AND2x4_ASAP7_75t_L g1677 ( 
.A(n_1645),
.B(n_1603),
.Y(n_1677)
);

INVx3_ASAP7_75t_L g1678 ( 
.A(n_1648),
.Y(n_1678)
);

INVx1_ASAP7_75t_L g1679 ( 
.A(n_1626),
.Y(n_1679)
);

HB1xp67_ASAP7_75t_L g1680 ( 
.A(n_1630),
.Y(n_1680)
);

INVx2_ASAP7_75t_L g1681 ( 
.A(n_1637),
.Y(n_1681)
);

INVx1_ASAP7_75t_SL g1682 ( 
.A(n_1618),
.Y(n_1682)
);

CKINVDCx20_ASAP7_75t_R g1683 ( 
.A(n_1621),
.Y(n_1683)
);

BUFx2_ASAP7_75t_L g1684 ( 
.A(n_1631),
.Y(n_1684)
);

NAND2xp5_ASAP7_75t_L g1685 ( 
.A(n_1658),
.B(n_1650),
.Y(n_1685)
);

NAND2xp5_ASAP7_75t_L g1686 ( 
.A(n_1658),
.B(n_1639),
.Y(n_1686)
);

AND2x2_ASAP7_75t_L g1687 ( 
.A(n_1662),
.B(n_1621),
.Y(n_1687)
);

AND2x2_ASAP7_75t_L g1688 ( 
.A(n_1662),
.B(n_1627),
.Y(n_1688)
);

NAND2xp5_ASAP7_75t_L g1689 ( 
.A(n_1661),
.B(n_1663),
.Y(n_1689)
);

INVx2_ASAP7_75t_L g1690 ( 
.A(n_1681),
.Y(n_1690)
);

AND2x2_ASAP7_75t_L g1691 ( 
.A(n_1664),
.B(n_1618),
.Y(n_1691)
);

AOI21xp33_ASAP7_75t_SL g1692 ( 
.A1(n_1670),
.A2(n_1649),
.B(n_1631),
.Y(n_1692)
);

INVxp33_ASAP7_75t_L g1693 ( 
.A(n_1661),
.Y(n_1693)
);

INVx2_ASAP7_75t_SL g1694 ( 
.A(n_1674),
.Y(n_1694)
);

AOI32xp33_ASAP7_75t_L g1695 ( 
.A1(n_1663),
.A2(n_1593),
.A3(n_1598),
.B1(n_1594),
.B2(n_1600),
.Y(n_1695)
);

INVx2_ASAP7_75t_L g1696 ( 
.A(n_1681),
.Y(n_1696)
);

INVx1_ASAP7_75t_L g1697 ( 
.A(n_1680),
.Y(n_1697)
);

INVx3_ASAP7_75t_L g1698 ( 
.A(n_1673),
.Y(n_1698)
);

AND2x4_ASAP7_75t_L g1699 ( 
.A(n_1673),
.B(n_1587),
.Y(n_1699)
);

AND2x2_ASAP7_75t_L g1700 ( 
.A(n_1659),
.B(n_1645),
.Y(n_1700)
);

AND2x2_ASAP7_75t_L g1701 ( 
.A(n_1659),
.B(n_1665),
.Y(n_1701)
);

INVx2_ASAP7_75t_L g1702 ( 
.A(n_1681),
.Y(n_1702)
);

INVx2_ASAP7_75t_SL g1703 ( 
.A(n_1674),
.Y(n_1703)
);

AND2x4_ASAP7_75t_L g1704 ( 
.A(n_1673),
.B(n_1587),
.Y(n_1704)
);

AND2x2_ASAP7_75t_L g1705 ( 
.A(n_1659),
.B(n_1645),
.Y(n_1705)
);

AND2x4_ASAP7_75t_L g1706 ( 
.A(n_1673),
.B(n_1677),
.Y(n_1706)
);

HB1xp67_ASAP7_75t_L g1707 ( 
.A(n_1680),
.Y(n_1707)
);

NOR2xp67_ASAP7_75t_L g1708 ( 
.A(n_1678),
.B(n_1631),
.Y(n_1708)
);

INVx1_ASAP7_75t_SL g1709 ( 
.A(n_1682),
.Y(n_1709)
);

INVx2_ASAP7_75t_L g1710 ( 
.A(n_1676),
.Y(n_1710)
);

INVx1_ASAP7_75t_L g1711 ( 
.A(n_1667),
.Y(n_1711)
);

BUFx2_ASAP7_75t_L g1712 ( 
.A(n_1674),
.Y(n_1712)
);

NAND2xp5_ASAP7_75t_L g1713 ( 
.A(n_1671),
.B(n_1654),
.Y(n_1713)
);

INVx1_ASAP7_75t_L g1714 ( 
.A(n_1667),
.Y(n_1714)
);

INVx1_ASAP7_75t_L g1715 ( 
.A(n_1668),
.Y(n_1715)
);

NOR4xp25_ASAP7_75t_L g1716 ( 
.A(n_1670),
.B(n_1591),
.C(n_1598),
.D(n_1600),
.Y(n_1716)
);

INVx1_ASAP7_75t_L g1717 ( 
.A(n_1668),
.Y(n_1717)
);

BUFx2_ASAP7_75t_L g1718 ( 
.A(n_1674),
.Y(n_1718)
);

OR2x2_ASAP7_75t_L g1719 ( 
.A(n_1656),
.B(n_1588),
.Y(n_1719)
);

AND2x4_ASAP7_75t_SL g1720 ( 
.A(n_1683),
.B(n_1641),
.Y(n_1720)
);

INVx2_ASAP7_75t_L g1721 ( 
.A(n_1676),
.Y(n_1721)
);

NAND2xp5_ASAP7_75t_SL g1722 ( 
.A(n_1678),
.B(n_1641),
.Y(n_1722)
);

OR2x2_ASAP7_75t_L g1723 ( 
.A(n_1716),
.B(n_1657),
.Y(n_1723)
);

AND2x2_ASAP7_75t_L g1724 ( 
.A(n_1712),
.B(n_1684),
.Y(n_1724)
);

NOR2x1_ASAP7_75t_L g1725 ( 
.A(n_1709),
.B(n_1678),
.Y(n_1725)
);

INVx2_ASAP7_75t_L g1726 ( 
.A(n_1690),
.Y(n_1726)
);

NAND2xp5_ASAP7_75t_L g1727 ( 
.A(n_1716),
.B(n_1657),
.Y(n_1727)
);

INVxp33_ASAP7_75t_L g1728 ( 
.A(n_1706),
.Y(n_1728)
);

INVx1_ASAP7_75t_L g1729 ( 
.A(n_1711),
.Y(n_1729)
);

AND2x2_ASAP7_75t_L g1730 ( 
.A(n_1712),
.B(n_1684),
.Y(n_1730)
);

NAND2xp5_ASAP7_75t_L g1731 ( 
.A(n_1695),
.B(n_1675),
.Y(n_1731)
);

INVx1_ASAP7_75t_L g1732 ( 
.A(n_1711),
.Y(n_1732)
);

AND2x2_ASAP7_75t_L g1733 ( 
.A(n_1712),
.B(n_1682),
.Y(n_1733)
);

AND2x2_ASAP7_75t_L g1734 ( 
.A(n_1718),
.B(n_1720),
.Y(n_1734)
);

NAND4xp25_ASAP7_75t_L g1735 ( 
.A(n_1689),
.B(n_1660),
.C(n_1669),
.D(n_1666),
.Y(n_1735)
);

AND2x2_ASAP7_75t_L g1736 ( 
.A(n_1718),
.B(n_1666),
.Y(n_1736)
);

OR2x2_ASAP7_75t_L g1737 ( 
.A(n_1685),
.B(n_1671),
.Y(n_1737)
);

INVx2_ASAP7_75t_L g1738 ( 
.A(n_1690),
.Y(n_1738)
);

BUFx2_ASAP7_75t_L g1739 ( 
.A(n_1718),
.Y(n_1739)
);

INVx1_ASAP7_75t_SL g1740 ( 
.A(n_1709),
.Y(n_1740)
);

AND2x2_ASAP7_75t_L g1741 ( 
.A(n_1688),
.B(n_1678),
.Y(n_1741)
);

NOR2xp33_ASAP7_75t_L g1742 ( 
.A(n_1689),
.B(n_1660),
.Y(n_1742)
);

INVx1_ASAP7_75t_L g1743 ( 
.A(n_1711),
.Y(n_1743)
);

INVxp67_ASAP7_75t_L g1744 ( 
.A(n_1707),
.Y(n_1744)
);

INVx1_ASAP7_75t_L g1745 ( 
.A(n_1714),
.Y(n_1745)
);

AND2x2_ASAP7_75t_L g1746 ( 
.A(n_1720),
.B(n_1666),
.Y(n_1746)
);

OR2x2_ASAP7_75t_L g1747 ( 
.A(n_1685),
.B(n_1656),
.Y(n_1747)
);

OR2x2_ASAP7_75t_L g1748 ( 
.A(n_1686),
.B(n_1656),
.Y(n_1748)
);

OR2x2_ASAP7_75t_L g1749 ( 
.A(n_1686),
.B(n_1676),
.Y(n_1749)
);

AND2x2_ASAP7_75t_L g1750 ( 
.A(n_1720),
.B(n_1672),
.Y(n_1750)
);

NAND2xp5_ASAP7_75t_L g1751 ( 
.A(n_1695),
.B(n_1675),
.Y(n_1751)
);

INVx1_ASAP7_75t_L g1752 ( 
.A(n_1714),
.Y(n_1752)
);

AND2x2_ASAP7_75t_L g1753 ( 
.A(n_1720),
.B(n_1672),
.Y(n_1753)
);

AND2x2_ASAP7_75t_L g1754 ( 
.A(n_1687),
.B(n_1672),
.Y(n_1754)
);

NAND2xp5_ASAP7_75t_L g1755 ( 
.A(n_1707),
.B(n_1679),
.Y(n_1755)
);

NOR2xp33_ASAP7_75t_L g1756 ( 
.A(n_1693),
.B(n_1669),
.Y(n_1756)
);

INVx2_ASAP7_75t_L g1757 ( 
.A(n_1690),
.Y(n_1757)
);

INVx2_ASAP7_75t_L g1758 ( 
.A(n_1690),
.Y(n_1758)
);

AND2x2_ASAP7_75t_L g1759 ( 
.A(n_1734),
.B(n_1706),
.Y(n_1759)
);

INVx2_ASAP7_75t_SL g1760 ( 
.A(n_1733),
.Y(n_1760)
);

NOR3xp33_ASAP7_75t_L g1761 ( 
.A(n_1742),
.B(n_1692),
.C(n_1697),
.Y(n_1761)
);

NOR3xp33_ASAP7_75t_L g1762 ( 
.A(n_1742),
.B(n_1692),
.C(n_1697),
.Y(n_1762)
);

OAI21xp5_ASAP7_75t_L g1763 ( 
.A1(n_1723),
.A2(n_1727),
.B(n_1725),
.Y(n_1763)
);

O2A1O1Ixp33_ASAP7_75t_L g1764 ( 
.A1(n_1723),
.A2(n_1693),
.B(n_1697),
.C(n_1721),
.Y(n_1764)
);

AOI22xp5_ASAP7_75t_L g1765 ( 
.A1(n_1727),
.A2(n_1646),
.B1(n_1699),
.B2(n_1704),
.Y(n_1765)
);

OAI211xp5_ASAP7_75t_L g1766 ( 
.A1(n_1735),
.A2(n_1698),
.B(n_1694),
.C(n_1703),
.Y(n_1766)
);

AOI22xp33_ASAP7_75t_L g1767 ( 
.A1(n_1731),
.A2(n_1751),
.B1(n_1735),
.B2(n_1600),
.Y(n_1767)
);

INVx1_ASAP7_75t_L g1768 ( 
.A(n_1729),
.Y(n_1768)
);

NOR2xp33_ASAP7_75t_L g1769 ( 
.A(n_1740),
.B(n_1706),
.Y(n_1769)
);

OAI21xp5_ASAP7_75t_SL g1770 ( 
.A1(n_1756),
.A2(n_1703),
.B(n_1694),
.Y(n_1770)
);

NOR2xp33_ASAP7_75t_L g1771 ( 
.A(n_1740),
.B(n_1706),
.Y(n_1771)
);

NAND2xp5_ASAP7_75t_L g1772 ( 
.A(n_1756),
.B(n_1687),
.Y(n_1772)
);

NOR2xp33_ASAP7_75t_L g1773 ( 
.A(n_1728),
.B(n_1706),
.Y(n_1773)
);

OR2x2_ASAP7_75t_L g1774 ( 
.A(n_1747),
.B(n_1713),
.Y(n_1774)
);

NOR2x1_ASAP7_75t_SL g1775 ( 
.A(n_1734),
.B(n_1722),
.Y(n_1775)
);

NAND2xp5_ASAP7_75t_L g1776 ( 
.A(n_1739),
.B(n_1687),
.Y(n_1776)
);

OAI21xp5_ASAP7_75t_L g1777 ( 
.A1(n_1725),
.A2(n_1722),
.B(n_1708),
.Y(n_1777)
);

OAI22xp5_ASAP7_75t_L g1778 ( 
.A1(n_1731),
.A2(n_1703),
.B1(n_1694),
.B2(n_1698),
.Y(n_1778)
);

NAND2xp5_ASAP7_75t_L g1779 ( 
.A(n_1739),
.B(n_1733),
.Y(n_1779)
);

OAI211xp5_ASAP7_75t_L g1780 ( 
.A1(n_1751),
.A2(n_1744),
.B(n_1724),
.C(n_1730),
.Y(n_1780)
);

NOR2xp33_ASAP7_75t_L g1781 ( 
.A(n_1737),
.B(n_1706),
.Y(n_1781)
);

OAI22xp33_ASAP7_75t_L g1782 ( 
.A1(n_1749),
.A2(n_1614),
.B1(n_1651),
.B2(n_1719),
.Y(n_1782)
);

OAI221xp5_ASAP7_75t_L g1783 ( 
.A1(n_1749),
.A2(n_1719),
.B1(n_1588),
.B2(n_1591),
.C(n_1594),
.Y(n_1783)
);

OAI22xp5_ASAP7_75t_L g1784 ( 
.A1(n_1750),
.A2(n_1698),
.B1(n_1678),
.B2(n_1708),
.Y(n_1784)
);

NOR2xp33_ASAP7_75t_L g1785 ( 
.A(n_1780),
.B(n_1760),
.Y(n_1785)
);

NAND2xp5_ASAP7_75t_SL g1786 ( 
.A(n_1761),
.B(n_1741),
.Y(n_1786)
);

AOI22xp5_ASAP7_75t_L g1787 ( 
.A1(n_1761),
.A2(n_1741),
.B1(n_1757),
.B2(n_1738),
.Y(n_1787)
);

INVx2_ASAP7_75t_L g1788 ( 
.A(n_1759),
.Y(n_1788)
);

NOR2xp33_ASAP7_75t_L g1789 ( 
.A(n_1779),
.B(n_1737),
.Y(n_1789)
);

NAND4xp25_ASAP7_75t_SL g1790 ( 
.A(n_1762),
.B(n_1736),
.C(n_1741),
.D(n_1750),
.Y(n_1790)
);

AOI22xp5_ASAP7_75t_L g1791 ( 
.A1(n_1762),
.A2(n_1758),
.B1(n_1757),
.B2(n_1726),
.Y(n_1791)
);

AND2x2_ASAP7_75t_L g1792 ( 
.A(n_1769),
.B(n_1753),
.Y(n_1792)
);

INVx1_ASAP7_75t_L g1793 ( 
.A(n_1768),
.Y(n_1793)
);

INVx1_ASAP7_75t_L g1794 ( 
.A(n_1776),
.Y(n_1794)
);

NAND2xp5_ASAP7_75t_L g1795 ( 
.A(n_1772),
.B(n_1754),
.Y(n_1795)
);

AOI21xp33_ASAP7_75t_SL g1796 ( 
.A1(n_1764),
.A2(n_1744),
.B(n_1747),
.Y(n_1796)
);

INVxp67_ASAP7_75t_SL g1797 ( 
.A(n_1763),
.Y(n_1797)
);

INVx1_ASAP7_75t_L g1798 ( 
.A(n_1774),
.Y(n_1798)
);

AOI221xp5_ASAP7_75t_L g1799 ( 
.A1(n_1767),
.A2(n_1721),
.B1(n_1710),
.B2(n_1729),
.C(n_1732),
.Y(n_1799)
);

NOR2xp33_ASAP7_75t_L g1800 ( 
.A(n_1771),
.B(n_1698),
.Y(n_1800)
);

INVx1_ASAP7_75t_L g1801 ( 
.A(n_1781),
.Y(n_1801)
);

INVx1_ASAP7_75t_L g1802 ( 
.A(n_1773),
.Y(n_1802)
);

AOI21xp33_ASAP7_75t_L g1803 ( 
.A1(n_1778),
.A2(n_1738),
.B(n_1726),
.Y(n_1803)
);

INVx2_ASAP7_75t_SL g1804 ( 
.A(n_1784),
.Y(n_1804)
);

AOI21xp33_ASAP7_75t_L g1805 ( 
.A1(n_1797),
.A2(n_1766),
.B(n_1765),
.Y(n_1805)
);

AOI21xp33_ASAP7_75t_SL g1806 ( 
.A1(n_1786),
.A2(n_1785),
.B(n_1804),
.Y(n_1806)
);

INVx1_ASAP7_75t_L g1807 ( 
.A(n_1791),
.Y(n_1807)
);

NAND2xp5_ASAP7_75t_L g1808 ( 
.A(n_1789),
.B(n_1754),
.Y(n_1808)
);

OR2x2_ASAP7_75t_L g1809 ( 
.A(n_1795),
.B(n_1748),
.Y(n_1809)
);

AOI21xp5_ASAP7_75t_L g1810 ( 
.A1(n_1797),
.A2(n_1775),
.B(n_1777),
.Y(n_1810)
);

INVxp67_ASAP7_75t_L g1811 ( 
.A(n_1785),
.Y(n_1811)
);

NOR2xp33_ASAP7_75t_L g1812 ( 
.A(n_1790),
.B(n_1770),
.Y(n_1812)
);

INVx1_ASAP7_75t_L g1813 ( 
.A(n_1793),
.Y(n_1813)
);

NAND2xp5_ASAP7_75t_L g1814 ( 
.A(n_1798),
.B(n_1736),
.Y(n_1814)
);

NAND2xp5_ASAP7_75t_L g1815 ( 
.A(n_1801),
.B(n_1724),
.Y(n_1815)
);

NOR4xp25_ASAP7_75t_L g1816 ( 
.A(n_1802),
.B(n_1783),
.C(n_1730),
.D(n_1782),
.Y(n_1816)
);

NOR2xp33_ASAP7_75t_L g1817 ( 
.A(n_1811),
.B(n_1796),
.Y(n_1817)
);

OAI21xp5_ASAP7_75t_L g1818 ( 
.A1(n_1816),
.A2(n_1787),
.B(n_1799),
.Y(n_1818)
);

NAND2xp5_ASAP7_75t_L g1819 ( 
.A(n_1808),
.B(n_1788),
.Y(n_1819)
);

INVx1_ASAP7_75t_L g1820 ( 
.A(n_1814),
.Y(n_1820)
);

NAND4xp25_ASAP7_75t_L g1821 ( 
.A(n_1812),
.B(n_1800),
.C(n_1794),
.D(n_1792),
.Y(n_1821)
);

INVx1_ASAP7_75t_L g1822 ( 
.A(n_1809),
.Y(n_1822)
);

OAI321xp33_ASAP7_75t_L g1823 ( 
.A1(n_1807),
.A2(n_1800),
.A3(n_1758),
.B1(n_1757),
.B2(n_1726),
.C(n_1738),
.Y(n_1823)
);

NAND2xp5_ASAP7_75t_L g1824 ( 
.A(n_1806),
.B(n_1803),
.Y(n_1824)
);

OR2x2_ASAP7_75t_L g1825 ( 
.A(n_1815),
.B(n_1748),
.Y(n_1825)
);

NAND2xp5_ASAP7_75t_L g1826 ( 
.A(n_1813),
.B(n_1688),
.Y(n_1826)
);

OAI221xp5_ASAP7_75t_SL g1827 ( 
.A1(n_1824),
.A2(n_1810),
.B1(n_1805),
.B2(n_1710),
.C(n_1721),
.Y(n_1827)
);

OAI31xp33_ASAP7_75t_L g1828 ( 
.A1(n_1817),
.A2(n_1710),
.A3(n_1721),
.B(n_1758),
.Y(n_1828)
);

OAI21xp33_ASAP7_75t_L g1829 ( 
.A1(n_1818),
.A2(n_1755),
.B(n_1743),
.Y(n_1829)
);

NAND2xp5_ASAP7_75t_L g1830 ( 
.A(n_1822),
.B(n_1753),
.Y(n_1830)
);

AOI221xp5_ASAP7_75t_L g1831 ( 
.A1(n_1823),
.A2(n_1821),
.B1(n_1820),
.B2(n_1826),
.C(n_1819),
.Y(n_1831)
);

OAI222xp33_ASAP7_75t_L g1832 ( 
.A1(n_1827),
.A2(n_1825),
.B1(n_1710),
.B2(n_1752),
.C1(n_1743),
.C2(n_1732),
.Y(n_1832)
);

AOI21xp5_ASAP7_75t_L g1833 ( 
.A1(n_1829),
.A2(n_1755),
.B(n_1752),
.Y(n_1833)
);

OAI211xp5_ASAP7_75t_SL g1834 ( 
.A1(n_1831),
.A2(n_1698),
.B(n_1745),
.C(n_1719),
.Y(n_1834)
);

OAI221xp5_ASAP7_75t_L g1835 ( 
.A1(n_1828),
.A2(n_1745),
.B1(n_1702),
.B2(n_1696),
.C(n_1705),
.Y(n_1835)
);

AOI22xp33_ASAP7_75t_L g1836 ( 
.A1(n_1830),
.A2(n_1702),
.B1(n_1696),
.B2(n_1699),
.Y(n_1836)
);

AOI211xp5_ASAP7_75t_L g1837 ( 
.A1(n_1827),
.A2(n_1705),
.B(n_1700),
.C(n_1699),
.Y(n_1837)
);

HB1xp67_ASAP7_75t_L g1838 ( 
.A(n_1832),
.Y(n_1838)
);

AND2x2_ASAP7_75t_L g1839 ( 
.A(n_1837),
.B(n_1746),
.Y(n_1839)
);

NOR2x1p5_ASAP7_75t_L g1840 ( 
.A(n_1834),
.B(n_1746),
.Y(n_1840)
);

AOI22xp5_ASAP7_75t_L g1841 ( 
.A1(n_1836),
.A2(n_1704),
.B1(n_1699),
.B2(n_1705),
.Y(n_1841)
);

NAND4xp75_ASAP7_75t_L g1842 ( 
.A(n_1833),
.B(n_1700),
.C(n_1701),
.D(n_1691),
.Y(n_1842)
);

NOR3xp33_ASAP7_75t_L g1843 ( 
.A(n_1838),
.B(n_1835),
.C(n_1702),
.Y(n_1843)
);

O2A1O1Ixp33_ASAP7_75t_L g1844 ( 
.A1(n_1839),
.A2(n_1700),
.B(n_1704),
.C(n_1699),
.Y(n_1844)
);

AOI221xp5_ASAP7_75t_L g1845 ( 
.A1(n_1841),
.A2(n_1699),
.B1(n_1704),
.B2(n_1696),
.C(n_1702),
.Y(n_1845)
);

OAI21xp5_ASAP7_75t_L g1846 ( 
.A1(n_1843),
.A2(n_1842),
.B(n_1840),
.Y(n_1846)
);

INVx1_ASAP7_75t_L g1847 ( 
.A(n_1846),
.Y(n_1847)
);

INVx2_ASAP7_75t_L g1848 ( 
.A(n_1847),
.Y(n_1848)
);

NAND2xp5_ASAP7_75t_SL g1849 ( 
.A(n_1847),
.B(n_1844),
.Y(n_1849)
);

AOI22xp5_ASAP7_75t_L g1850 ( 
.A1(n_1848),
.A2(n_1845),
.B1(n_1704),
.B2(n_1696),
.Y(n_1850)
);

INVx1_ASAP7_75t_L g1851 ( 
.A(n_1849),
.Y(n_1851)
);

NAND2xp5_ASAP7_75t_L g1852 ( 
.A(n_1851),
.B(n_1850),
.Y(n_1852)
);

AOI22xp5_ASAP7_75t_L g1853 ( 
.A1(n_1851),
.A2(n_1704),
.B1(n_1701),
.B2(n_1715),
.Y(n_1853)
);

OAI22xp5_ASAP7_75t_L g1854 ( 
.A1(n_1853),
.A2(n_1717),
.B1(n_1715),
.B2(n_1714),
.Y(n_1854)
);

AOI21xp5_ASAP7_75t_L g1855 ( 
.A1(n_1854),
.A2(n_1852),
.B(n_1717),
.Y(n_1855)
);

HB1xp67_ASAP7_75t_L g1856 ( 
.A(n_1855),
.Y(n_1856)
);

OAI221xp5_ASAP7_75t_L g1857 ( 
.A1(n_1856),
.A2(n_1717),
.B1(n_1715),
.B2(n_1701),
.C(n_1713),
.Y(n_1857)
);

AOI211xp5_ASAP7_75t_L g1858 ( 
.A1(n_1857),
.A2(n_1691),
.B(n_1673),
.C(n_1677),
.Y(n_1858)
);


endmodule