module fake_jpeg_28383_n_357 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_357);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_357;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

BUFx4f_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

INVx4_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_8),
.Y(n_21)
);

HB1xp67_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_16),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_11),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_8),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

BUFx4f_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_1),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_14),
.Y(n_32)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_15),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_10),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_8),
.Y(n_36)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_17),
.Y(n_37)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_38),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_26),
.Y(n_39)
);

INVx6_ASAP7_75t_L g81 ( 
.A(n_39),
.Y(n_81)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_17),
.Y(n_40)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_40),
.Y(n_62)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_18),
.Y(n_41)
);

INVx6_ASAP7_75t_L g91 ( 
.A(n_41),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_25),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_42),
.B(n_45),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_17),
.Y(n_43)
);

INVx5_ASAP7_75t_SL g83 ( 
.A(n_43),
.Y(n_83)
);

BUFx12_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_44),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_25),
.Y(n_45)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_46),
.Y(n_67)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_17),
.Y(n_47)
);

INVx8_ASAP7_75t_L g90 ( 
.A(n_47),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_26),
.Y(n_48)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_48),
.Y(n_84)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_20),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_49),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_32),
.B(n_16),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_50),
.B(n_53),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_26),
.Y(n_51)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_51),
.Y(n_93)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_52),
.Y(n_88)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_20),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_31),
.B(n_0),
.Y(n_54)
);

AND2x2_ASAP7_75t_L g64 ( 
.A(n_54),
.B(n_19),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_20),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_55),
.Y(n_70)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_29),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_56),
.Y(n_74)
);

NOR2x1_ASAP7_75t_L g60 ( 
.A(n_42),
.B(n_32),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_60),
.B(n_61),
.Y(n_106)
);

CKINVDCx14_ASAP7_75t_R g61 ( 
.A(n_54),
.Y(n_61)
);

CKINVDCx16_ASAP7_75t_R g63 ( 
.A(n_44),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_63),
.B(n_64),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_45),
.B(n_34),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g121 ( 
.A(n_65),
.B(n_79),
.Y(n_121)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_49),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_66),
.B(n_86),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_39),
.B(n_31),
.C(n_36),
.Y(n_68)
);

XNOR2xp5_ASAP7_75t_L g122 ( 
.A(n_68),
.B(n_73),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_38),
.A2(n_33),
.B1(n_24),
.B2(n_28),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_71),
.A2(n_75),
.B1(n_23),
.B2(n_36),
.Y(n_130)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_49),
.B(n_19),
.Y(n_72)
);

INVx1_ASAP7_75t_SL g115 ( 
.A(n_72),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_41),
.A2(n_34),
.B1(n_33),
.B2(n_30),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_40),
.A2(n_33),
.B1(n_21),
.B2(n_27),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_43),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_78),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_53),
.B(n_21),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_46),
.A2(n_27),
.B1(n_30),
.B2(n_24),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_80),
.A2(n_85),
.B1(n_29),
.B2(n_35),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_55),
.B(n_28),
.Y(n_82)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_82),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_L g85 ( 
.A1(n_40),
.A2(n_52),
.B1(n_37),
.B2(n_56),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_44),
.B(n_19),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_43),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_87),
.Y(n_112)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_55),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_89),
.Y(n_126)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_56),
.Y(n_92)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_92),
.Y(n_98)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_84),
.Y(n_94)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_94),
.Y(n_133)
);

CKINVDCx12_ASAP7_75t_R g95 ( 
.A(n_57),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_95),
.B(n_102),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_L g96 ( 
.A1(n_81),
.A2(n_52),
.B1(n_19),
.B2(n_18),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_96),
.A2(n_101),
.B1(n_110),
.B2(n_119),
.Y(n_154)
);

INVx8_ASAP7_75t_L g97 ( 
.A(n_90),
.Y(n_97)
);

INVx4_ASAP7_75t_SL g148 ( 
.A(n_97),
.Y(n_148)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_71),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_99),
.B(n_100),
.Y(n_140)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_72),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_77),
.A2(n_19),
.B1(n_18),
.B2(n_23),
.Y(n_101)
);

INVx5_ASAP7_75t_L g102 ( 
.A(n_90),
.Y(n_102)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_84),
.Y(n_103)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_103),
.Y(n_143)
);

BUFx12_ASAP7_75t_L g104 ( 
.A(n_57),
.Y(n_104)
);

BUFx10_ASAP7_75t_L g135 ( 
.A(n_104),
.Y(n_135)
);

INVx5_ASAP7_75t_L g105 ( 
.A(n_78),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_105),
.B(n_113),
.Y(n_147)
);

O2A1O1Ixp33_ASAP7_75t_L g107 ( 
.A1(n_73),
.A2(n_51),
.B(n_48),
.C(n_39),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_107),
.A2(n_131),
.B1(n_58),
.B2(n_93),
.Y(n_142)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_72),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_108),
.B(n_120),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_109),
.A2(n_117),
.B1(n_29),
.B2(n_22),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_77),
.A2(n_23),
.B1(n_11),
.B2(n_12),
.Y(n_110)
);

BUFx3_ASAP7_75t_L g113 ( 
.A(n_93),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_64),
.A2(n_68),
.B1(n_76),
.B2(n_60),
.Y(n_117)
);

OR2x6_ASAP7_75t_L g118 ( 
.A(n_64),
.B(n_29),
.Y(n_118)
);

NAND2x1_ASAP7_75t_SL g150 ( 
.A(n_118),
.B(n_129),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_91),
.A2(n_23),
.B1(n_11),
.B2(n_12),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_59),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_91),
.A2(n_81),
.B1(n_83),
.B2(n_88),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_L g161 ( 
.A1(n_123),
.A2(n_127),
.B1(n_115),
.B2(n_102),
.Y(n_161)
);

BUFx8_ASAP7_75t_L g124 ( 
.A(n_83),
.Y(n_124)
);

INVx3_ASAP7_75t_L g155 ( 
.A(n_124),
.Y(n_155)
);

INVx8_ASAP7_75t_L g127 ( 
.A(n_74),
.Y(n_127)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_127),
.Y(n_144)
);

BUFx12f_ASAP7_75t_L g128 ( 
.A(n_87),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_128),
.Y(n_136)
);

OA22x2_ASAP7_75t_L g129 ( 
.A1(n_62),
.A2(n_88),
.B1(n_89),
.B2(n_48),
.Y(n_129)
);

AND2x2_ASAP7_75t_L g137 ( 
.A(n_129),
.B(n_130),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_62),
.A2(n_51),
.B1(n_47),
.B2(n_43),
.Y(n_131)
);

AND2x2_ASAP7_75t_SL g132 ( 
.A(n_74),
.B(n_36),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_132),
.B(n_70),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_122),
.B(n_58),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_134),
.B(n_145),
.Y(n_173)
);

FAx1_ASAP7_75t_SL g138 ( 
.A(n_114),
.B(n_22),
.CI(n_44),
.CON(n_138),
.SN(n_138)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_138),
.B(n_121),
.Y(n_172)
);

AND2x2_ASAP7_75t_L g171 ( 
.A(n_139),
.B(n_150),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_142),
.A2(n_105),
.B1(n_97),
.B2(n_125),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_122),
.B(n_70),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_126),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_149),
.Y(n_166)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_129),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_151),
.B(n_159),
.Y(n_182)
);

AND2x2_ASAP7_75t_L g192 ( 
.A(n_152),
.B(n_153),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_118),
.B(n_100),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_118),
.B(n_115),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_156),
.B(n_160),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_99),
.A2(n_130),
.B1(n_107),
.B2(n_118),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_157),
.A2(n_94),
.B1(n_103),
.B2(n_98),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_126),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_158),
.Y(n_175)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_129),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_118),
.B(n_29),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_161),
.A2(n_128),
.B1(n_104),
.B2(n_2),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_106),
.B(n_67),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_SL g168 ( 
.A(n_162),
.B(n_120),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_108),
.B(n_47),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_163),
.B(n_164),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_116),
.B(n_69),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_132),
.A2(n_69),
.B1(n_47),
.B2(n_67),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_165),
.A2(n_104),
.B1(n_1),
.B2(n_2),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_SL g167 ( 
.A1(n_156),
.A2(n_132),
.B(n_98),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_SL g220 ( 
.A1(n_167),
.A2(n_158),
.B(n_136),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_SL g211 ( 
.A(n_168),
.B(n_172),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_169),
.A2(n_174),
.B1(n_178),
.B2(n_180),
.Y(n_214)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_147),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_170),
.B(n_181),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_137),
.A2(n_157),
.B1(n_151),
.B2(n_159),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_176),
.A2(n_185),
.B1(n_178),
.B2(n_184),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_137),
.A2(n_131),
.B1(n_113),
.B2(n_112),
.Y(n_178)
);

BUFx2_ASAP7_75t_L g179 ( 
.A(n_149),
.Y(n_179)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_179),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_137),
.A2(n_112),
.B1(n_111),
.B2(n_124),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_139),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_140),
.B(n_145),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_183),
.B(n_193),
.Y(n_203)
);

CKINVDCx16_ASAP7_75t_R g184 ( 
.A(n_164),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_184),
.B(n_197),
.Y(n_205)
);

AOI22xp33_ASAP7_75t_L g185 ( 
.A1(n_160),
.A2(n_111),
.B1(n_124),
.B2(n_128),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_165),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_186),
.B(n_187),
.Y(n_221)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_140),
.Y(n_187)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_146),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_189),
.B(n_191),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_190),
.A2(n_195),
.B1(n_155),
.B2(n_148),
.Y(n_229)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_142),
.Y(n_191)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_133),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_133),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_194),
.B(n_196),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_134),
.B(n_0),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_162),
.B(n_15),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_141),
.B(n_16),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_198),
.B(n_200),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_154),
.A2(n_13),
.B1(n_12),
.B2(n_2),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_199),
.A2(n_186),
.B1(n_191),
.B2(n_180),
.Y(n_222)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_143),
.Y(n_200)
);

NOR2x1_ASAP7_75t_L g201 ( 
.A(n_150),
.B(n_0),
.Y(n_201)
);

AO21x1_ASAP7_75t_L g213 ( 
.A1(n_201),
.A2(n_138),
.B(n_144),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_179),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_202),
.Y(n_237)
);

NOR3xp33_ASAP7_75t_L g206 ( 
.A(n_187),
.B(n_141),
.C(n_154),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_206),
.B(n_215),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_L g207 ( 
.A1(n_192),
.A2(n_163),
.B(n_150),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_L g236 ( 
.A1(n_207),
.A2(n_212),
.B(n_220),
.Y(n_236)
);

OAI22x1_ASAP7_75t_L g209 ( 
.A1(n_176),
.A2(n_138),
.B1(n_153),
.B2(n_152),
.Y(n_209)
);

AOI22xp33_ASAP7_75t_L g255 ( 
.A1(n_209),
.A2(n_229),
.B1(n_234),
.B2(n_223),
.Y(n_255)
);

AOI21xp5_ASAP7_75t_L g212 ( 
.A1(n_192),
.A2(n_136),
.B(n_144),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_213),
.B(n_230),
.Y(n_242)
);

INVxp67_ASAP7_75t_L g215 ( 
.A(n_201),
.Y(n_215)
);

INVx1_ASAP7_75t_SL g216 ( 
.A(n_171),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_216),
.B(n_218),
.Y(n_243)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_179),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_217),
.B(n_226),
.Y(n_262)
);

NAND3xp33_ASAP7_75t_L g218 ( 
.A(n_168),
.B(n_13),
.C(n_1),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_222),
.A2(n_233),
.B1(n_235),
.B2(n_166),
.Y(n_260)
);

AOI21xp5_ASAP7_75t_L g223 ( 
.A1(n_192),
.A2(n_148),
.B(n_155),
.Y(n_223)
);

INVxp67_ASAP7_75t_L g261 ( 
.A(n_223),
.Y(n_261)
);

AND2x2_ASAP7_75t_L g224 ( 
.A(n_182),
.B(n_143),
.Y(n_224)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_224),
.Y(n_252)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_182),
.Y(n_226)
);

AND2x2_ASAP7_75t_L g227 ( 
.A(n_177),
.B(n_148),
.Y(n_227)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_227),
.Y(n_254)
);

CKINVDCx16_ASAP7_75t_R g228 ( 
.A(n_188),
.Y(n_228)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_228),
.Y(n_256)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_169),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_171),
.A2(n_135),
.B1(n_13),
.B2(n_3),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_231),
.A2(n_199),
.B1(n_188),
.B2(n_170),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_195),
.A2(n_135),
.B1(n_1),
.B2(n_3),
.Y(n_232)
);

CKINVDCx14_ASAP7_75t_R g251 ( 
.A(n_232),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_174),
.A2(n_0),
.B1(n_3),
.B2(n_4),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_177),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_207),
.B(n_173),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_238),
.B(n_247),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_216),
.B(n_173),
.C(n_183),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_239),
.B(n_250),
.C(n_219),
.Y(n_266)
);

BUFx12f_ASAP7_75t_SL g240 ( 
.A(n_209),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_SL g279 ( 
.A1(n_240),
.A2(n_215),
.B(n_224),
.Y(n_279)
);

BUFx24_ASAP7_75t_SL g244 ( 
.A(n_211),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_244),
.B(n_245),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_230),
.A2(n_181),
.B1(n_171),
.B2(n_167),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_246),
.A2(n_233),
.B1(n_235),
.B2(n_217),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_212),
.B(n_196),
.Y(n_247)
);

A2O1A1O1Ixp25_ASAP7_75t_L g248 ( 
.A1(n_213),
.A2(n_201),
.B(n_190),
.C(n_189),
.D(n_166),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_248),
.B(n_257),
.Y(n_271)
);

CKINVDCx16_ASAP7_75t_R g249 ( 
.A(n_225),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_249),
.B(n_253),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_203),
.B(n_220),
.C(n_228),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_202),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_L g277 ( 
.A1(n_255),
.A2(n_260),
.B1(n_232),
.B2(n_234),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_203),
.B(n_175),
.Y(n_257)
);

CKINVDCx16_ASAP7_75t_R g258 ( 
.A(n_225),
.Y(n_258)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_258),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_204),
.B(n_175),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_259),
.B(n_231),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_238),
.B(n_204),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_263),
.B(n_265),
.Y(n_290)
);

CKINVDCx16_ASAP7_75t_R g264 ( 
.A(n_262),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_264),
.B(n_267),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_259),
.B(n_213),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_266),
.B(n_274),
.Y(n_292)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_237),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_239),
.B(n_219),
.C(n_227),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_269),
.B(n_278),
.C(n_280),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_250),
.A2(n_221),
.B1(n_229),
.B2(n_226),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_270),
.A2(n_281),
.B1(n_246),
.B2(n_245),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_257),
.B(n_221),
.Y(n_273)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_273),
.Y(n_302)
);

OAI21xp5_ASAP7_75t_SL g303 ( 
.A1(n_277),
.A2(n_279),
.B(n_241),
.Y(n_303)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_236),
.B(n_214),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_247),
.B(n_227),
.C(n_224),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_260),
.A2(n_214),
.B1(n_222),
.B2(n_205),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_L g299 ( 
.A1(n_282),
.A2(n_251),
.B1(n_242),
.B2(n_252),
.Y(n_299)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_262),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_283),
.B(n_285),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_256),
.B(n_210),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_284),
.B(n_256),
.Y(n_291)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_237),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_SL g286 ( 
.A(n_272),
.B(n_211),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_286),
.B(n_293),
.Y(n_306)
);

INVx2_ASAP7_75t_SL g287 ( 
.A(n_267),
.Y(n_287)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_287),
.Y(n_307)
);

HB1xp67_ASAP7_75t_L g288 ( 
.A(n_276),
.Y(n_288)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_288),
.Y(n_313)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_291),
.Y(n_315)
);

HB1xp67_ASAP7_75t_L g293 ( 
.A(n_273),
.Y(n_293)
);

AND2x2_ASAP7_75t_L g294 ( 
.A(n_278),
.B(n_240),
.Y(n_294)
);

AOI21xp5_ASAP7_75t_L g318 ( 
.A1(n_294),
.A2(n_296),
.B(n_303),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_284),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_295),
.B(n_304),
.Y(n_311)
);

AO21x1_ASAP7_75t_L g296 ( 
.A1(n_279),
.A2(n_236),
.B(n_242),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_SL g319 ( 
.A1(n_298),
.A2(n_254),
.B1(n_261),
.B2(n_248),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_L g305 ( 
.A1(n_299),
.A2(n_282),
.B1(n_280),
.B2(n_252),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_266),
.B(n_268),
.C(n_269),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_301),
.B(n_268),
.C(n_274),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_275),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g324 ( 
.A1(n_305),
.A2(n_319),
.B1(n_294),
.B2(n_261),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_308),
.B(n_309),
.C(n_310),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_301),
.B(n_270),
.C(n_263),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_289),
.B(n_271),
.C(n_265),
.Y(n_310)
);

XOR2xp5_ASAP7_75t_L g312 ( 
.A(n_290),
.B(n_271),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g327 ( 
.A(n_312),
.B(n_314),
.Y(n_327)
);

XNOR2xp5_ASAP7_75t_SL g314 ( 
.A(n_290),
.B(n_281),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_289),
.B(n_254),
.C(n_208),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_316),
.B(n_291),
.C(n_298),
.Y(n_330)
);

XNOR2xp5_ASAP7_75t_SL g317 ( 
.A(n_292),
.B(n_243),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_L g322 ( 
.A(n_317),
.B(n_292),
.Y(n_322)
);

AOI21xp5_ASAP7_75t_SL g320 ( 
.A1(n_318),
.A2(n_296),
.B(n_303),
.Y(n_320)
);

OAI21xp5_ASAP7_75t_SL g339 ( 
.A1(n_320),
.A2(n_194),
.B(n_193),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_SL g321 ( 
.A(n_306),
.B(n_300),
.Y(n_321)
);

AOI21xp5_ASAP7_75t_L g334 ( 
.A1(n_321),
.A2(n_322),
.B(n_326),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_L g340 ( 
.A1(n_324),
.A2(n_325),
.B1(n_329),
.B2(n_331),
.Y(n_340)
);

AOI22xp5_ASAP7_75t_L g325 ( 
.A1(n_311),
.A2(n_287),
.B1(n_294),
.B2(n_302),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_319),
.Y(n_326)
);

INVxp67_ASAP7_75t_L g328 ( 
.A(n_318),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_SL g336 ( 
.A1(n_328),
.A2(n_309),
.B1(n_317),
.B2(n_310),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_313),
.B(n_297),
.Y(n_329)
);

OAI21x1_ASAP7_75t_L g335 ( 
.A1(n_330),
.A2(n_316),
.B(n_314),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_315),
.B(n_208),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_307),
.Y(n_332)
);

AOI22xp5_ASAP7_75t_L g333 ( 
.A1(n_332),
.A2(n_287),
.B1(n_304),
.B2(n_200),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_333),
.B(n_4),
.Y(n_346)
);

XNOR2xp5_ASAP7_75t_L g342 ( 
.A(n_335),
.B(n_341),
.Y(n_342)
);

INVxp67_ASAP7_75t_L g344 ( 
.A(n_336),
.Y(n_344)
);

NOR2xp67_ASAP7_75t_L g337 ( 
.A(n_320),
.B(n_312),
.Y(n_337)
);

OAI21xp5_ASAP7_75t_L g347 ( 
.A1(n_337),
.A2(n_338),
.B(n_339),
.Y(n_347)
);

NOR2xp67_ASAP7_75t_SL g338 ( 
.A(n_330),
.B(n_308),
.Y(n_338)
);

AOI22xp5_ASAP7_75t_SL g341 ( 
.A1(n_328),
.A2(n_135),
.B1(n_5),
.B2(n_6),
.Y(n_341)
);

AOI22xp5_ASAP7_75t_SL g343 ( 
.A1(n_334),
.A2(n_336),
.B1(n_327),
.B2(n_340),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_343),
.B(n_346),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_341),
.B(n_323),
.C(n_322),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_345),
.B(n_348),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_SL g348 ( 
.A(n_340),
.B(n_323),
.Y(n_348)
);

AOI21xp5_ASAP7_75t_L g349 ( 
.A1(n_347),
.A2(n_135),
.B(n_6),
.Y(n_349)
);

AOI322xp5_ASAP7_75t_L g354 ( 
.A1(n_349),
.A2(n_350),
.A3(n_5),
.B1(n_7),
.B2(n_9),
.C1(n_10),
.C2(n_351),
.Y(n_354)
);

NOR4xp25_ASAP7_75t_L g350 ( 
.A(n_344),
.B(n_345),
.C(n_342),
.D(n_135),
.Y(n_350)
);

AOI22xp5_ASAP7_75t_SL g353 ( 
.A1(n_352),
.A2(n_344),
.B1(n_7),
.B2(n_8),
.Y(n_353)
);

AOI21xp5_ASAP7_75t_SL g355 ( 
.A1(n_353),
.A2(n_354),
.B(n_7),
.Y(n_355)
);

XOR2x2_ASAP7_75t_L g356 ( 
.A(n_355),
.B(n_9),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_356),
.B(n_10),
.Y(n_357)
);


endmodule