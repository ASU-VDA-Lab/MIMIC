module fake_jpeg_990_n_335 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_335);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_335;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx12f_ASAP7_75t_L g15 ( 
.A(n_2),
.Y(n_15)
);

INVx4_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_8),
.Y(n_17)
);

INVx6_ASAP7_75t_SL g18 ( 
.A(n_2),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_3),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_0),
.B(n_10),
.Y(n_24)
);

BUFx12_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

BUFx24_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

INVxp67_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_12),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_0),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_11),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_5),
.Y(n_35)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_12),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_9),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_9),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_33),
.Y(n_39)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_39),
.Y(n_72)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_16),
.Y(n_40)
);

INVx2_ASAP7_75t_SL g71 ( 
.A(n_40),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_16),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_41),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_24),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_42),
.B(n_44),
.Y(n_98)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_15),
.Y(n_43)
);

INVx5_ASAP7_75t_L g106 ( 
.A(n_43),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_24),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_27),
.B(n_14),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_45),
.B(n_60),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_16),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_46),
.Y(n_87)
);

CKINVDCx14_ASAP7_75t_R g47 ( 
.A(n_18),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_47),
.B(n_53),
.Y(n_70)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_33),
.Y(n_48)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_48),
.Y(n_77)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_15),
.Y(n_49)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_49),
.Y(n_100)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_19),
.Y(n_50)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_50),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_28),
.B(n_14),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_51),
.B(n_52),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_20),
.B(n_0),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_18),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_15),
.Y(n_54)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_54),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_20),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_55),
.B(n_61),
.Y(n_73)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_15),
.Y(n_56)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_56),
.Y(n_113)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_15),
.Y(n_57)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_57),
.Y(n_86)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_20),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g110 ( 
.A(n_58),
.Y(n_110)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_21),
.Y(n_59)
);

BUFx2_ASAP7_75t_L g80 ( 
.A(n_59),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_28),
.B(n_9),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_22),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_22),
.A2(n_29),
.B1(n_37),
.B2(n_19),
.Y(n_62)
);

OA22x2_ASAP7_75t_L g95 ( 
.A1(n_62),
.A2(n_66),
.B1(n_59),
.B2(n_49),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_38),
.B(n_13),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_63),
.B(n_68),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_22),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_64),
.B(n_67),
.Y(n_81)
);

BUFx12_ASAP7_75t_L g65 ( 
.A(n_26),
.Y(n_65)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_65),
.Y(n_78)
);

INVx5_ASAP7_75t_L g66 ( 
.A(n_21),
.Y(n_66)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_66),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_29),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_29),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_52),
.B(n_32),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_69),
.B(n_88),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_42),
.A2(n_21),
.B1(n_35),
.B2(n_37),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_75),
.A2(n_89),
.B1(n_90),
.B2(n_92),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_44),
.A2(n_31),
.B1(n_32),
.B2(n_34),
.Y(n_76)
);

OA22x2_ASAP7_75t_L g117 ( 
.A1(n_76),
.A2(n_95),
.B1(n_104),
.B2(n_65),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_41),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_84),
.B(n_112),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_62),
.A2(n_35),
.B1(n_21),
.B2(n_38),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_85),
.A2(n_94),
.B1(n_99),
.B2(n_54),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_60),
.B(n_34),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_55),
.A2(n_35),
.B1(n_21),
.B2(n_31),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_61),
.A2(n_35),
.B1(n_30),
.B2(n_23),
.Y(n_90)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_39),
.Y(n_91)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_91),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_64),
.A2(n_35),
.B1(n_30),
.B2(n_23),
.Y(n_92)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_48),
.Y(n_93)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_93),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_67),
.A2(n_17),
.B1(n_26),
.B2(n_36),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_63),
.B(n_17),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g147 ( 
.A(n_96),
.B(n_108),
.Y(n_147)
);

OAI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_68),
.A2(n_36),
.B1(n_26),
.B2(n_13),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_L g102 ( 
.A1(n_50),
.A2(n_26),
.B1(n_36),
.B2(n_25),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_102),
.A2(n_25),
.B1(n_3),
.B2(n_4),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_40),
.A2(n_26),
.B1(n_25),
.B2(n_2),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_103),
.A2(n_65),
.B1(n_43),
.B2(n_54),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_45),
.A2(n_25),
.B1(n_1),
.B2(n_2),
.Y(n_104)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_57),
.Y(n_107)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_107),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_53),
.B(n_0),
.Y(n_108)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_41),
.Y(n_109)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_109),
.Y(n_121)
);

INVx6_ASAP7_75t_L g111 ( 
.A(n_58),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_111),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_46),
.Y(n_112)
);

INVx6_ASAP7_75t_L g114 ( 
.A(n_46),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_114),
.Y(n_138)
);

O2A1O1Ixp33_ASAP7_75t_L g115 ( 
.A1(n_95),
.A2(n_65),
.B(n_43),
.C(n_56),
.Y(n_115)
);

AOI21xp5_ASAP7_75t_L g164 ( 
.A1(n_115),
.A2(n_83),
.B(n_114),
.Y(n_164)
);

AND2x2_ASAP7_75t_L g157 ( 
.A(n_117),
.B(n_148),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_118),
.A2(n_124),
.B1(n_130),
.B2(n_131),
.Y(n_191)
);

INVx11_ASAP7_75t_L g120 ( 
.A(n_78),
.Y(n_120)
);

INVx4_ASAP7_75t_L g176 ( 
.A(n_120),
.Y(n_176)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_91),
.Y(n_122)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_122),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_97),
.B(n_1),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_126),
.B(n_145),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_127),
.A2(n_134),
.B1(n_136),
.B2(n_71),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_70),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_129),
.B(n_153),
.Y(n_188)
);

AOI22xp33_ASAP7_75t_L g130 ( 
.A1(n_105),
.A2(n_25),
.B1(n_4),
.B2(n_5),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_L g131 ( 
.A1(n_69),
.A2(n_1),
.B1(n_4),
.B2(n_5),
.Y(n_131)
);

BUFx2_ASAP7_75t_L g132 ( 
.A(n_80),
.Y(n_132)
);

BUFx2_ASAP7_75t_L g167 ( 
.A(n_132),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_101),
.A2(n_4),
.B1(n_6),
.B2(n_7),
.Y(n_134)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_106),
.Y(n_135)
);

BUFx12f_ASAP7_75t_L g180 ( 
.A(n_135),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_85),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_136)
);

HB1xp67_ASAP7_75t_L g139 ( 
.A(n_71),
.Y(n_139)
);

INVx1_ASAP7_75t_SL g170 ( 
.A(n_139),
.Y(n_170)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_93),
.Y(n_140)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_140),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_L g141 ( 
.A1(n_72),
.A2(n_8),
.B1(n_6),
.B2(n_7),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_141),
.A2(n_144),
.B1(n_133),
.B2(n_125),
.Y(n_186)
);

INVx4_ASAP7_75t_L g142 ( 
.A(n_106),
.Y(n_142)
);

INVx3_ASAP7_75t_L g165 ( 
.A(n_142),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_94),
.A2(n_77),
.B1(n_95),
.B2(n_73),
.Y(n_143)
);

AOI21xp33_ASAP7_75t_L g160 ( 
.A1(n_143),
.A2(n_104),
.B(n_109),
.Y(n_160)
);

AND2x2_ASAP7_75t_L g144 ( 
.A(n_71),
.B(n_6),
.Y(n_144)
);

NAND2x1_ASAP7_75t_L g184 ( 
.A(n_144),
.B(n_134),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_98),
.B(n_8),
.Y(n_145)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_83),
.Y(n_146)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_146),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_79),
.B(n_86),
.C(n_107),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_88),
.B(n_96),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_149),
.B(n_154),
.Y(n_166)
);

INVx6_ASAP7_75t_L g150 ( 
.A(n_82),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g181 ( 
.A(n_150),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_81),
.B(n_113),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_151),
.B(n_155),
.Y(n_178)
);

INVx11_ASAP7_75t_L g152 ( 
.A(n_78),
.Y(n_152)
);

INVx5_ASAP7_75t_SL g174 ( 
.A(n_152),
.Y(n_174)
);

CKINVDCx16_ASAP7_75t_R g153 ( 
.A(n_80),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g154 ( 
.A(n_76),
.B(n_95),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_113),
.B(n_100),
.Y(n_155)
);

AND2x2_ASAP7_75t_L g197 ( 
.A(n_158),
.B(n_164),
.Y(n_197)
);

AOI21xp5_ASAP7_75t_SL g201 ( 
.A1(n_160),
.A2(n_191),
.B(n_178),
.Y(n_201)
);

AOI22xp33_ASAP7_75t_L g161 ( 
.A1(n_154),
.A2(n_100),
.B1(n_82),
.B2(n_87),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_161),
.A2(n_168),
.B1(n_172),
.B2(n_182),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_124),
.A2(n_86),
.B1(n_87),
.B2(n_110),
.Y(n_168)
);

AOI21xp33_ASAP7_75t_L g169 ( 
.A1(n_147),
.A2(n_110),
.B(n_111),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_SL g222 ( 
.A(n_169),
.B(n_186),
.Y(n_222)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_122),
.Y(n_171)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_171),
.Y(n_199)
);

AOI22xp33_ASAP7_75t_L g172 ( 
.A1(n_115),
.A2(n_74),
.B1(n_151),
.B2(n_140),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_129),
.B(n_74),
.Y(n_173)
);

CKINVDCx14_ASAP7_75t_R g226 ( 
.A(n_173),
.Y(n_226)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_123),
.Y(n_175)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_175),
.Y(n_204)
);

INVx13_ASAP7_75t_L g177 ( 
.A(n_120),
.Y(n_177)
);

INVx1_ASAP7_75t_SL g214 ( 
.A(n_177),
.Y(n_214)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_123),
.Y(n_179)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_179),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_136),
.A2(n_127),
.B1(n_117),
.B2(n_128),
.Y(n_182)
);

INVx13_ASAP7_75t_L g183 ( 
.A(n_152),
.Y(n_183)
);

CKINVDCx16_ASAP7_75t_R g206 ( 
.A(n_183),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_184),
.B(n_132),
.Y(n_203)
);

AND2x6_ASAP7_75t_L g185 ( 
.A(n_128),
.B(n_147),
.Y(n_185)
);

AND2x6_ASAP7_75t_L g224 ( 
.A(n_185),
.B(n_187),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_186),
.A2(n_138),
.B1(n_119),
.B2(n_150),
.Y(n_213)
);

AND2x6_ASAP7_75t_L g187 ( 
.A(n_117),
.B(n_116),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_148),
.B(n_155),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_189),
.B(n_146),
.Y(n_195)
);

INVx13_ASAP7_75t_L g190 ( 
.A(n_153),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_190),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_132),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_192),
.B(n_138),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_SL g193 ( 
.A1(n_157),
.A2(n_117),
.B(n_133),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_SL g232 ( 
.A1(n_193),
.A2(n_198),
.B(n_201),
.Y(n_232)
);

MAJx2_ASAP7_75t_L g194 ( 
.A(n_157),
.B(n_144),
.C(n_137),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_194),
.B(n_200),
.C(n_207),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_195),
.B(n_200),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_178),
.B(n_121),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_196),
.B(n_202),
.Y(n_233)
);

NOR2x1_ASAP7_75t_L g198 ( 
.A(n_166),
.B(n_121),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_157),
.B(n_137),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_184),
.B(n_135),
.Y(n_202)
);

OAI21xp33_ASAP7_75t_L g240 ( 
.A1(n_203),
.A2(n_221),
.B(n_222),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_188),
.B(n_142),
.C(n_119),
.Y(n_207)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_156),
.Y(n_210)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_210),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_182),
.B(n_119),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_211),
.B(n_180),
.C(n_197),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_167),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_212),
.B(n_223),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_213),
.A2(n_192),
.B1(n_167),
.B2(n_181),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_163),
.B(n_138),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_SL g248 ( 
.A(n_215),
.B(n_219),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_187),
.A2(n_168),
.B1(n_158),
.B2(n_164),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_216),
.A2(n_174),
.B1(n_181),
.B2(n_176),
.Y(n_236)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_217),
.Y(n_238)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_156),
.Y(n_218)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_218),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_170),
.B(n_162),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_SL g220 ( 
.A1(n_185),
.A2(n_184),
.B(n_159),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_SL g235 ( 
.A1(n_220),
.A2(n_225),
.B(n_190),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_170),
.B(n_162),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_165),
.B(n_175),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_SL g225 ( 
.A1(n_159),
.A2(n_171),
.B(n_179),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_221),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_227),
.B(n_230),
.Y(n_258)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_228),
.Y(n_262)
);

CKINVDCx16_ASAP7_75t_R g230 ( 
.A(n_217),
.Y(n_230)
);

AOI21xp5_ASAP7_75t_L g234 ( 
.A1(n_193),
.A2(n_165),
.B(n_176),
.Y(n_234)
);

OAI21xp5_ASAP7_75t_SL g266 ( 
.A1(n_234),
.A2(n_235),
.B(n_239),
.Y(n_266)
);

OAI22xp33_ASAP7_75t_SL g272 ( 
.A1(n_236),
.A2(n_214),
.B1(n_234),
.B2(n_238),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_237),
.B(n_207),
.Y(n_254)
);

AO21x1_ASAP7_75t_L g239 ( 
.A1(n_220),
.A2(n_177),
.B(n_183),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_194),
.B(n_174),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_242),
.B(n_247),
.C(n_225),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_244),
.B(n_229),
.Y(n_275)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_199),
.Y(n_245)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_245),
.Y(n_273)
);

BUFx2_ASAP7_75t_L g246 ( 
.A(n_204),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_246),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_196),
.B(n_180),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_SL g249 ( 
.A1(n_201),
.A2(n_180),
.B(n_198),
.Y(n_249)
);

OAI21xp5_ASAP7_75t_L g261 ( 
.A1(n_249),
.A2(n_252),
.B(n_208),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_226),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_250),
.B(n_251),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_197),
.A2(n_180),
.B1(n_211),
.B2(n_216),
.Y(n_251)
);

AOI21xp5_ASAP7_75t_L g252 ( 
.A1(n_197),
.A2(n_222),
.B(n_203),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_L g253 ( 
.A1(n_213),
.A2(n_202),
.B1(n_209),
.B2(n_198),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_253),
.B(n_218),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_254),
.B(n_256),
.Y(n_279)
);

INVx4_ASAP7_75t_L g255 ( 
.A(n_239),
.Y(n_255)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_255),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_L g259 ( 
.A1(n_236),
.A2(n_209),
.B1(n_224),
.B2(n_208),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_259),
.A2(n_263),
.B1(n_270),
.B2(n_271),
.Y(n_283)
);

OA22x2_ASAP7_75t_L g260 ( 
.A1(n_238),
.A2(n_224),
.B1(n_199),
.B2(n_210),
.Y(n_260)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_260),
.Y(n_277)
);

AOI21xp5_ASAP7_75t_L g278 ( 
.A1(n_261),
.A2(n_274),
.B(n_232),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_227),
.B(n_204),
.Y(n_265)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_265),
.Y(n_280)
);

INVx4_ASAP7_75t_L g267 ( 
.A(n_239),
.Y(n_267)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_267),
.Y(n_287)
);

INVx4_ASAP7_75t_L g268 ( 
.A(n_250),
.Y(n_268)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_268),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_SL g269 ( 
.A(n_248),
.B(n_205),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_SL g284 ( 
.A(n_269),
.B(n_248),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_252),
.A2(n_205),
.B1(n_212),
.B2(n_206),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_L g271 ( 
.A1(n_244),
.A2(n_206),
.B1(n_214),
.B2(n_233),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_272),
.A2(n_270),
.B1(n_255),
.B2(n_267),
.Y(n_286)
);

OAI21xp5_ASAP7_75t_L g274 ( 
.A1(n_249),
.A2(n_240),
.B(n_232),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_275),
.B(n_229),
.C(n_237),
.Y(n_281)
);

AOI21xp5_ASAP7_75t_L g296 ( 
.A1(n_278),
.A2(n_261),
.B(n_274),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_281),
.B(n_275),
.C(n_254),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_265),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_SL g295 ( 
.A(n_282),
.B(n_284),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_268),
.B(n_235),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_SL g297 ( 
.A(n_285),
.B(n_288),
.Y(n_297)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_286),
.Y(n_292)
);

CKINVDCx16_ASAP7_75t_R g288 ( 
.A(n_258),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_263),
.A2(n_251),
.B1(n_233),
.B2(n_242),
.Y(n_289)
);

BUFx2_ASAP7_75t_L g304 ( 
.A(n_289),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_257),
.A2(n_231),
.B1(n_243),
.B2(n_245),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_291),
.B(n_258),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g311 ( 
.A(n_293),
.B(n_300),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_291),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_294),
.B(n_298),
.Y(n_306)
);

AOI21xp5_ASAP7_75t_L g307 ( 
.A1(n_296),
.A2(n_299),
.B(n_266),
.Y(n_307)
);

AO221x1_ASAP7_75t_L g299 ( 
.A1(n_283),
.A2(n_286),
.B1(n_289),
.B2(n_260),
.C(n_269),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_281),
.B(n_256),
.C(n_271),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_279),
.B(n_247),
.C(n_260),
.Y(n_301)
);

INVxp67_ASAP7_75t_L g305 ( 
.A(n_301),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_279),
.B(n_260),
.C(n_259),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_302),
.B(n_277),
.Y(n_312)
);

AOI322xp5_ASAP7_75t_SL g303 ( 
.A1(n_278),
.A2(n_257),
.A3(n_241),
.B1(n_264),
.B2(n_266),
.C1(n_231),
.C2(n_243),
.Y(n_303)
);

OR2x2_ASAP7_75t_L g313 ( 
.A(n_303),
.B(n_277),
.Y(n_313)
);

OR2x2_ASAP7_75t_L g320 ( 
.A(n_307),
.B(n_314),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_SL g308 ( 
.A(n_293),
.B(n_283),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_L g317 ( 
.A(n_308),
.B(n_301),
.Y(n_317)
);

HB1xp67_ASAP7_75t_L g309 ( 
.A(n_297),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_309),
.B(n_310),
.Y(n_319)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_295),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_312),
.B(n_290),
.C(n_292),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_L g315 ( 
.A1(n_313),
.A2(n_280),
.B1(n_302),
.B2(n_304),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_292),
.A2(n_276),
.B1(n_287),
.B2(n_290),
.Y(n_314)
);

OR2x2_ASAP7_75t_L g324 ( 
.A(n_315),
.B(n_316),
.Y(n_324)
);

XOR2xp5_ASAP7_75t_L g325 ( 
.A(n_317),
.B(n_296),
.Y(n_325)
);

BUFx4f_ASAP7_75t_SL g318 ( 
.A(n_309),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_318),
.B(n_280),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_311),
.B(n_300),
.C(n_304),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_321),
.B(n_306),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_321),
.B(n_305),
.C(n_312),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_322),
.B(n_323),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_SL g329 ( 
.A(n_325),
.B(n_276),
.Y(n_329)
);

OAI21xp5_ASAP7_75t_L g327 ( 
.A1(n_326),
.A2(n_320),
.B(n_319),
.Y(n_327)
);

AOI322xp5_ASAP7_75t_L g330 ( 
.A1(n_327),
.A2(n_329),
.A3(n_318),
.B1(n_326),
.B2(n_287),
.C1(n_324),
.C2(n_320),
.Y(n_330)
);

INVxp67_ASAP7_75t_L g332 ( 
.A(n_330),
.Y(n_332)
);

AOI322xp5_ASAP7_75t_L g331 ( 
.A1(n_328),
.A2(n_246),
.A3(n_262),
.B1(n_264),
.B2(n_273),
.C1(n_318),
.C2(n_327),
.Y(n_331)
);

BUFx24_ASAP7_75t_SL g333 ( 
.A(n_332),
.Y(n_333)
);

OAI21xp5_ASAP7_75t_L g334 ( 
.A1(n_333),
.A2(n_331),
.B(n_262),
.Y(n_334)
);

XNOR2xp5_ASAP7_75t_L g335 ( 
.A(n_334),
.B(n_273),
.Y(n_335)
);


endmodule