module fake_ariane_367_n_2250 (n_83, n_8, n_56, n_60, n_170, n_190, n_160, n_64, n_179, n_180, n_119, n_124, n_167, n_90, n_195, n_38, n_213, n_47, n_110, n_153, n_18, n_197, n_221, n_86, n_75, n_89, n_67, n_176, n_149, n_34, n_158, n_172, n_69, n_95, n_175, n_92, n_143, n_183, n_203, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_181, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_115, n_133, n_66, n_205, n_71, n_24, n_7, n_109, n_208, n_96, n_156, n_209, n_49, n_20, n_174, n_100, n_17, n_50, n_187, n_132, n_62, n_210, n_147, n_204, n_200, n_51, n_166, n_76, n_218, n_103, n_79, n_26, n_3, n_46, n_220, n_0, n_84, n_36, n_199, n_91, n_159, n_107, n_189, n_72, n_105, n_128, n_217, n_44, n_30, n_82, n_178, n_31, n_42, n_57, n_131, n_201, n_70, n_222, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_214, n_48, n_94, n_101, n_4, n_134, n_188, n_185, n_2, n_32, n_37, n_58, n_65, n_123, n_212, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_198, n_148, n_164, n_52, n_157, n_184, n_177, n_135, n_73, n_77, n_171, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_182, n_196, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_206, n_13, n_27, n_207, n_29, n_41, n_219, n_140, n_55, n_191, n_151, n_136, n_192, n_28, n_80, n_146, n_211, n_194, n_97, n_154, n_215, n_142, n_161, n_14, n_163, n_88, n_186, n_141, n_68, n_116, n_104, n_202, n_145, n_78, n_193, n_39, n_59, n_63, n_99, n_216, n_16, n_5, n_155, n_127, n_223, n_35, n_54, n_25, n_2250);

input n_83;
input n_8;
input n_56;
input n_60;
input n_170;
input n_190;
input n_160;
input n_64;
input n_179;
input n_180;
input n_119;
input n_124;
input n_167;
input n_90;
input n_195;
input n_38;
input n_213;
input n_47;
input n_110;
input n_153;
input n_18;
input n_197;
input n_221;
input n_86;
input n_75;
input n_89;
input n_67;
input n_176;
input n_149;
input n_34;
input n_158;
input n_172;
input n_69;
input n_95;
input n_175;
input n_92;
input n_143;
input n_183;
input n_203;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_181;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_205;
input n_71;
input n_24;
input n_7;
input n_109;
input n_208;
input n_96;
input n_156;
input n_209;
input n_49;
input n_20;
input n_174;
input n_100;
input n_17;
input n_50;
input n_187;
input n_132;
input n_62;
input n_210;
input n_147;
input n_204;
input n_200;
input n_51;
input n_166;
input n_76;
input n_218;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_220;
input n_0;
input n_84;
input n_36;
input n_199;
input n_91;
input n_159;
input n_107;
input n_189;
input n_72;
input n_105;
input n_128;
input n_217;
input n_44;
input n_30;
input n_82;
input n_178;
input n_31;
input n_42;
input n_57;
input n_131;
input n_201;
input n_70;
input n_222;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_214;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_188;
input n_185;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_212;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_198;
input n_148;
input n_164;
input n_52;
input n_157;
input n_184;
input n_177;
input n_135;
input n_73;
input n_77;
input n_171;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_182;
input n_196;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_206;
input n_13;
input n_27;
input n_207;
input n_29;
input n_41;
input n_219;
input n_140;
input n_55;
input n_191;
input n_151;
input n_136;
input n_192;
input n_28;
input n_80;
input n_146;
input n_211;
input n_194;
input n_97;
input n_154;
input n_215;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_186;
input n_141;
input n_68;
input n_116;
input n_104;
input n_202;
input n_145;
input n_78;
input n_193;
input n_39;
input n_59;
input n_63;
input n_99;
input n_216;
input n_16;
input n_5;
input n_155;
input n_127;
input n_223;
input n_35;
input n_54;
input n_25;

output n_2250;

wire n_913;
wire n_1681;
wire n_2163;
wire n_1486;
wire n_1507;
wire n_1938;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_2131;
wire n_423;
wire n_1383;
wire n_2182;
wire n_603;
wire n_373;
wire n_2135;
wire n_1250;
wire n_2030;
wire n_1169;
wire n_789;
wire n_850;
wire n_1916;
wire n_610;
wire n_245;
wire n_1713;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_2002;
wire n_1463;
wire n_2243;
wire n_1238;
wire n_2011;
wire n_1515;
wire n_817;
wire n_1837;
wire n_924;
wire n_781;
wire n_2013;
wire n_1566;
wire n_717;
wire n_2006;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_2207;
wire n_524;
wire n_1214;
wire n_634;
wire n_1839;
wire n_1246;
wire n_1138;
wire n_2042;
wire n_2123;
wire n_1853;
wire n_764;
wire n_1503;
wire n_2238;
wire n_462;
wire n_1196;
wire n_1181;
wire n_1999;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_232;
wire n_2084;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1835;
wire n_1457;
wire n_377;
wire n_1682;
wire n_1836;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_945;
wire n_958;
wire n_2248;
wire n_813;
wire n_419;
wire n_1985;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1909;
wire n_2156;
wire n_1184;
wire n_1961;
wire n_1535;
wire n_500;
wire n_754;
wire n_665;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1979;
wire n_1277;
wire n_2107;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_2221;
wire n_672;
wire n_740;
wire n_1283;
wire n_1974;
wire n_1736;
wire n_1018;
wire n_2200;
wire n_259;
wire n_953;
wire n_1364;
wire n_1888;
wire n_1224;
wire n_2109;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_242;
wire n_645;
wire n_1944;
wire n_331;
wire n_559;
wire n_2233;
wire n_495;
wire n_267;
wire n_1988;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_1936;
wire n_2149;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_2078;
wire n_1145;
wire n_971;
wire n_2201;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_2049;
wire n_1522;
wire n_518;
wire n_1207;
wire n_786;
wire n_1404;
wire n_868;
wire n_2232;
wire n_1847;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_2227;
wire n_1539;
wire n_884;
wire n_1851;
wire n_2162;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_2192;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_1900;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_1889;
wire n_587;
wire n_1977;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_352;
wire n_899;
wire n_1703;
wire n_611;
wire n_1295;
wire n_2060;
wire n_1850;
wire n_365;
wire n_238;
wire n_2004;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_661;
wire n_2098;
wire n_1751;
wire n_300;
wire n_533;
wire n_1917;
wire n_1924;
wire n_438;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_1811;
wire n_2045;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_1840;
wire n_376;
wire n_512;
wire n_1597;
wire n_1771;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_2061;
wire n_2094;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_237;
wire n_2043;
wire n_780;
wire n_1918;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1949;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_2077;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_490;
wire n_1461;
wire n_1391;
wire n_1947;
wire n_225;
wire n_1599;
wire n_1876;
wire n_1006;
wire n_1830;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_2038;
wire n_2116;
wire n_2145;
wire n_1838;
wire n_1594;
wire n_680;
wire n_1935;
wire n_287;
wire n_1716;
wire n_302;
wire n_1872;
wire n_380;
wire n_1585;
wire n_1432;
wire n_2245;
wire n_249;
wire n_1108;
wire n_851;
wire n_444;
wire n_355;
wire n_1590;
wire n_1351;
wire n_2216;
wire n_1274;
wire n_257;
wire n_652;
wire n_1819;
wire n_475;
wire n_947;
wire n_2134;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_1833;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_1884;
wire n_460;
wire n_1555;
wire n_1842;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_2166;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_2185;
wire n_1376;
wire n_513;
wire n_288;
wire n_1292;
wire n_1178;
wire n_1972;
wire n_2015;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_2202;
wire n_2072;
wire n_306;
wire n_436;
wire n_324;
wire n_2087;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_967;
wire n_1083;
wire n_2161;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1787;
wire n_1389;
wire n_2155;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_1717;
wire n_1812;
wire n_824;
wire n_428;
wire n_2172;
wire n_892;
wire n_1880;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_2219;
wire n_1855;
wire n_2100;
wire n_990;
wire n_1623;
wire n_1903;
wire n_867;
wire n_2147;
wire n_1226;
wire n_2224;
wire n_944;
wire n_749;
wire n_1932;
wire n_1780;
wire n_1970;
wire n_1920;
wire n_2083;
wire n_815;
wire n_542;
wire n_2167;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1911;
wire n_1825;
wire n_1908;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1832;
wire n_1841;
wire n_1680;
wire n_2066;
wire n_964;
wire n_1627;
wire n_2220;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_1731;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_1914;
wire n_934;
wire n_2213;
wire n_1447;
wire n_1220;
wire n_356;
wire n_2019;
wire n_698;
wire n_2130;
wire n_1674;
wire n_2021;
wire n_2025;
wire n_2160;
wire n_1992;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_2142;
wire n_1633;
wire n_404;
wire n_1913;
wire n_2069;
wire n_1058;
wire n_347;
wire n_1042;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_2223;
wire n_1279;
wire n_2144;
wire n_564;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_1728;
wire n_370;
wire n_706;
wire n_2120;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_2041;
wire n_2113;
wire n_1933;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_1817;
wire n_2168;
wire n_552;
wire n_348;
wire n_670;
wire n_1826;
wire n_379;
wire n_264;
wire n_441;
wire n_1951;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_2132;
wire n_980;
wire n_1618;
wire n_1869;
wire n_1743;
wire n_905;
wire n_720;
wire n_926;
wire n_1943;
wire n_1802;
wire n_2178;
wire n_2112;
wire n_1163;
wire n_1795;
wire n_1384;
wire n_2237;
wire n_2146;
wire n_1868;
wire n_1501;
wire n_2241;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_2099;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1879;
wire n_1886;
wire n_1648;
wire n_2187;
wire n_1413;
wire n_2129;
wire n_855;
wire n_808;
wire n_1365;
wire n_553;
wire n_2059;
wire n_1439;
wire n_814;
wire n_578;
wire n_2074;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_2122;
wire n_320;
wire n_1414;
wire n_1134;
wire n_2067;
wire n_1484;
wire n_1901;
wire n_647;
wire n_2055;
wire n_2027;
wire n_1423;
wire n_2117;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_1939;
wire n_2242;
wire n_1906;
wire n_529;
wire n_1899;
wire n_2195;
wire n_502;
wire n_2194;
wire n_1467;
wire n_247;
wire n_1828;
wire n_2159;
wire n_1798;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_1105;
wire n_547;
wire n_604;
wire n_677;
wire n_439;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_2102;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_2023;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_699;
wire n_727;
wire n_301;
wire n_1726;
wire n_2075;
wire n_1945;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_2031;
wire n_2118;
wire n_325;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_2225;
wire n_986;
wire n_1104;
wire n_1963;
wire n_887;
wire n_729;
wire n_2057;
wire n_2218;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1693;
wire n_2125;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_2184;
wire n_314;
wire n_1823;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_2033;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_2217;
wire n_321;
wire n_2226;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1863;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_2214;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_1859;
wire n_262;
wire n_1502;
wire n_1523;
wire n_2190;
wire n_1478;
wire n_1883;
wire n_1969;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_845;
wire n_888;
wire n_1649;
wire n_1677;
wire n_1927;
wire n_1297;
wire n_551;
wire n_417;
wire n_1708;
wire n_343;
wire n_1222;
wire n_1844;
wire n_582;
wire n_1957;
wire n_1953;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_1919;
wire n_534;
wire n_1791;
wire n_2124;
wire n_1894;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_1898;
wire n_451;
wire n_745;
wire n_1741;
wire n_1572;
wire n_1907;
wire n_1793;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1975;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_2119;
wire n_769;
wire n_1797;
wire n_1753;
wire n_1990;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_1895;
wire n_982;
wire n_1800;
wire n_915;
wire n_1075;
wire n_2008;
wire n_454;
wire n_298;
wire n_1331;
wire n_1890;
wire n_1529;
wire n_1227;
wire n_2127;
wire n_655;
wire n_1860;
wire n_1734;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_2211;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_509;
wire n_1854;
wire n_666;
wire n_1747;
wire n_2071;
wire n_430;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_2082;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_456;
wire n_1867;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_2140;
wire n_873;
wire n_1301;
wire n_1748;
wire n_2157;
wire n_1966;
wire n_1243;
wire n_2171;
wire n_1400;
wire n_342;
wire n_2035;
wire n_1466;
wire n_1527;
wire n_1513;
wire n_358;
wire n_1783;
wire n_608;
wire n_1538;
wire n_2128;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1993;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1954;
wire n_1668;
wire n_1878;
wire n_1605;
wire n_1078;
wire n_266;
wire n_1897;
wire n_2137;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_2026;
wire n_1786;
wire n_480;
wire n_1327;
wire n_1475;
wire n_642;
wire n_1804;
wire n_2106;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_1757;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_2091;
wire n_393;
wire n_1632;
wire n_1769;
wire n_474;
wire n_1929;
wire n_1950;
wire n_805;
wire n_2032;
wire n_2090;
wire n_295;
wire n_1658;
wire n_2249;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1997;
wire n_1137;
wire n_1873;
wire n_1258;
wire n_640;
wire n_463;
wire n_1476;
wire n_1524;
wire n_1733;
wire n_1856;
wire n_2016;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1874;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_1807;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_1784;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_283;
wire n_806;
wire n_1984;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_1824;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_1822;
wire n_682;
wire n_1616;
wire n_819;
wire n_1971;
wire n_586;
wire n_1429;
wire n_1324;
wire n_2064;
wire n_1778;
wire n_1776;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1759;
wire n_1829;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_2022;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_1815;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_1864;
wire n_1887;
wire n_1208;
wire n_1987;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_2170;
wire n_790;
wire n_2244;
wire n_2143;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_2198;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_1852;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_2222;
wire n_1995;
wire n_1877;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_2076;
wire n_2133;
wire n_2203;
wire n_833;
wire n_1426;
wire n_2247;
wire n_2230;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_2001;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_2158;
wire n_1201;
wire n_1288;
wire n_858;
wire n_1185;
wire n_2173;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_2070;
wire n_2136;
wire n_426;
wire n_433;
wire n_398;
wire n_1090;
wire n_1367;
wire n_2044;
wire n_928;
wire n_253;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_420;
wire n_1291;
wire n_562;
wire n_2020;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1882;
wire n_1976;
wire n_1023;
wire n_1881;
wire n_988;
wire n_914;
wire n_330;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_1958;
wire n_467;
wire n_1511;
wire n_2177;
wire n_1422;
wire n_1965;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_538;
wire n_1517;
wire n_2036;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_2003;
wire n_2210;
wire n_1307;
wire n_1128;
wire n_2053;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1921;
wire n_1356;
wire n_1341;
wire n_2234;
wire n_1504;
wire n_1955;
wire n_2110;
wire n_1773;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_1948;
wire n_810;
wire n_1290;
wire n_1959;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_2121;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_1960;
wire n_2068;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_1968;
wire n_1885;
wire n_639;
wire n_452;
wire n_673;
wire n_2196;
wire n_1038;
wire n_1978;
wire n_414;
wire n_571;
wire n_1521;
wire n_1694;
wire n_1940;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_409;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_2007;
wire n_526;
wire n_1994;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1973;
wire n_1444;
wire n_1803;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_1739;
wire n_1814;
wire n_532;
wire n_2154;
wire n_2236;
wire n_1789;
wire n_763;
wire n_1986;
wire n_2174;
wire n_540;
wire n_692;
wire n_2054;
wire n_1857;
wire n_984;
wire n_1687;
wire n_2073;
wire n_2150;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_2046;
wire n_1816;
wire n_1910;
wire n_1756;
wire n_1606;
wire n_2189;
wire n_395;
wire n_621;
wire n_1587;
wire n_2093;
wire n_2018;
wire n_1772;
wire n_1014;
wire n_724;
wire n_2204;
wire n_1427;
wire n_1481;
wire n_2040;
wire n_493;
wire n_1311;
wire n_2199;
wire n_1956;
wire n_1589;
wire n_2151;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_2231;
wire n_697;
wire n_622;
wire n_1626;
wire n_1962;
wire n_1335;
wire n_1715;
wire n_296;
wire n_880;
wire n_793;
wire n_2114;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_1785;
wire n_792;
wire n_1262;
wire n_1942;
wire n_2180;
wire n_580;
wire n_1579;
wire n_494;
wire n_2181;
wire n_434;
wire n_2014;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1893;
wire n_1183;
wire n_1326;
wire n_1805;
wire n_981;
wire n_2141;
wire n_1110;
wire n_1758;
wire n_243;
wire n_1407;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_2010;
wire n_1054;
wire n_508;
wire n_1679;
wire n_2126;
wire n_1952;
wire n_1858;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_1834;
wire n_978;
wire n_1011;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_2050;
wire n_2197;
wire n_783;
wire n_556;
wire n_1127;
wire n_1536;
wire n_1471;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_1980;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_1998;
wire n_2165;
wire n_541;
wire n_499;
wire n_1775;
wire n_788;
wire n_908;
wire n_1036;
wire n_2169;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_2028;
wire n_919;
wire n_1663;
wire n_2092;
wire n_2175;
wire n_1625;
wire n_2086;
wire n_1926;
wire n_318;
wire n_1458;
wire n_244;
wire n_679;
wire n_1630;
wire n_663;
wire n_1720;
wire n_443;
wire n_2176;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_1922;
wire n_1735;
wire n_1788;
wire n_391;
wire n_940;
wire n_1537;
wire n_2138;
wire n_2065;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_1930;
wire n_765;
wire n_1809;
wire n_1904;
wire n_1843;
wire n_2000;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_2096;
wire n_2186;
wire n_1530;
wire n_2215;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_898;
wire n_857;
wire n_363;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1937;
wire n_2012;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_2039;
wire n_1755;
wire n_1285;
wire n_733;
wire n_761;
wire n_2212;
wire n_731;
wire n_336;
wire n_1813;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_2111;
wire n_1996;
wire n_1106;
wire n_2009;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_2024;
wire n_1348;
wire n_753;
wire n_1770;
wire n_701;
wire n_1003;
wire n_1125;
wire n_2103;
wire n_1710;
wire n_1865;
wire n_309;
wire n_1344;
wire n_1390;
wire n_485;
wire n_401;
wire n_1792;
wire n_504;
wire n_2062;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_2153;
wire n_1510;
wire n_2139;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_567;
wire n_369;
wire n_240;
wire n_1727;
wire n_2235;
wire n_1991;
wire n_1575;
wire n_1848;
wire n_1892;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_1902;
wire n_997;
wire n_635;
wire n_2206;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_2034;
wire n_1845;
wire n_1934;
wire n_2101;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_2104;
wire n_1265;
wire n_1576;
wire n_2105;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1806;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_2088;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_2005;
wire n_2048;
wire n_1696;
wire n_498;
wire n_1875;
wire n_1059;
wire n_684;
wire n_2108;
wire n_1039;
wire n_2246;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1831;
wire n_2191;
wire n_1497;
wire n_1866;
wire n_2056;
wire n_459;
wire n_1136;
wire n_1782;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_838;
wire n_383;
wire n_1558;
wire n_1941;
wire n_1316;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_1915;
wire n_723;
wire n_1393;
wire n_2240;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_1781;
wire n_709;
wire n_809;
wire n_2085;
wire n_1686;
wire n_1964;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_2188;
wire n_1982;
wire n_2097;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_308;
wire n_1223;
wire n_1768;
wire n_2193;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1983;
wire n_1041;
wire n_2115;
wire n_993;
wire n_1862;
wire n_948;
wire n_2017;
wire n_922;
wire n_1004;
wire n_1810;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_1923;
wire n_1764;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_1337;
wire n_774;
wire n_1946;
wire n_2148;
wire n_933;
wire n_1779;
wire n_596;
wire n_954;
wire n_2051;
wire n_1168;
wire n_1821;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_664;
wire n_252;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1896;
wire n_2164;
wire n_1732;
wire n_415;
wire n_1967;
wire n_2179;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_2052;
wire n_537;
wire n_1063;
wire n_991;
wire n_2183;
wire n_2205;
wire n_389;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1799;
wire n_2080;
wire n_2058;
wire n_1126;
wire n_2029;
wire n_1846;
wire n_1912;
wire n_938;
wire n_1891;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_2209;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_1928;
wire n_946;
wire n_757;
wire n_2047;
wire n_375;
wire n_1655;
wire n_1818;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_2081;
wire n_265;
wire n_1583;
wire n_1604;
wire n_1631;
wire n_1702;
wire n_275;
wire n_1794;
wire n_1375;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_1827;
wire n_866;
wire n_246;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_1115;
wire n_2229;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_2239;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_1871;
wire n_718;
wire n_329;
wire n_1434;
wire n_340;
wire n_1905;
wire n_1569;
wire n_548;
wire n_289;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_1870;
wire n_2063;
wire n_1925;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1861;
wire n_2079;
wire n_1228;
wire n_2152;
wire n_1931;
wire n_1244;
wire n_1796;
wire n_411;
wire n_484;
wire n_849;
wire n_2095;
wire n_1820;
wire n_357;
wire n_412;
wire n_1251;
wire n_1989;
wire n_447;
wire n_1421;
wire n_2208;
wire n_1762;
wire n_1233;
wire n_1808;
wire n_1574;
wire n_1672;
wire n_2228;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_1981;
wire n_2037;
wire n_359;
wire n_1308;
wire n_796;
wire n_573;
wire n_531;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_2089;
wire n_1487;
wire n_675;

BUFx3_ASAP7_75t_L g224 ( 
.A(n_73),
.Y(n_224)
);

BUFx6f_ASAP7_75t_L g225 ( 
.A(n_201),
.Y(n_225)
);

BUFx3_ASAP7_75t_L g226 ( 
.A(n_197),
.Y(n_226)
);

BUFx6f_ASAP7_75t_L g227 ( 
.A(n_52),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_118),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_141),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_110),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_184),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_162),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_198),
.Y(n_233)
);

BUFx3_ASAP7_75t_L g234 ( 
.A(n_30),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_48),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_111),
.Y(n_236)
);

BUFx10_ASAP7_75t_L g237 ( 
.A(n_101),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_169),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_116),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_129),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_109),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_121),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_83),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_119),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_68),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_138),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_193),
.Y(n_247)
);

BUFx3_ASAP7_75t_L g248 ( 
.A(n_170),
.Y(n_248)
);

BUFx6f_ASAP7_75t_L g249 ( 
.A(n_165),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_149),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_0),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_123),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_194),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_148),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_220),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_108),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_156),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_66),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_78),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_37),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_63),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_161),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_79),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_43),
.Y(n_264)
);

BUFx10_ASAP7_75t_L g265 ( 
.A(n_58),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_30),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_207),
.Y(n_267)
);

BUFx10_ASAP7_75t_L g268 ( 
.A(n_221),
.Y(n_268)
);

BUFx10_ASAP7_75t_L g269 ( 
.A(n_185),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_7),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_208),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_144),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_23),
.Y(n_273)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_152),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_18),
.Y(n_275)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_179),
.Y(n_276)
);

INVx1_ASAP7_75t_SL g277 ( 
.A(n_130),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_142),
.Y(n_278)
);

INVx2_ASAP7_75t_SL g279 ( 
.A(n_143),
.Y(n_279)
);

BUFx10_ASAP7_75t_L g280 ( 
.A(n_171),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_55),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_1),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_217),
.Y(n_283)
);

BUFx2_ASAP7_75t_L g284 ( 
.A(n_146),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_15),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_47),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_134),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_3),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_173),
.Y(n_289)
);

INVxp67_ASAP7_75t_SL g290 ( 
.A(n_206),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_124),
.Y(n_291)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_140),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_43),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_91),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_53),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_137),
.Y(n_296)
);

BUFx2_ASAP7_75t_L g297 ( 
.A(n_81),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_98),
.Y(n_298)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_34),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_223),
.Y(n_300)
);

INVx1_ASAP7_75t_SL g301 ( 
.A(n_209),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_106),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_33),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_136),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_71),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_10),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_77),
.Y(n_307)
);

BUFx2_ASAP7_75t_L g308 ( 
.A(n_4),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_139),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_150),
.Y(n_310)
);

INVx1_ASAP7_75t_SL g311 ( 
.A(n_20),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_29),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_222),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_89),
.Y(n_314)
);

BUFx8_ASAP7_75t_SL g315 ( 
.A(n_15),
.Y(n_315)
);

CKINVDCx16_ASAP7_75t_R g316 ( 
.A(n_5),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_40),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_107),
.Y(n_318)
);

BUFx8_ASAP7_75t_SL g319 ( 
.A(n_211),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_55),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_177),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_153),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_159),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_70),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_213),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_164),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_40),
.Y(n_327)
);

INVx1_ASAP7_75t_SL g328 ( 
.A(n_114),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_176),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_202),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_166),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_48),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_188),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_126),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_127),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_37),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_19),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_216),
.Y(n_338)
);

BUFx6f_ASAP7_75t_L g339 ( 
.A(n_44),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_163),
.Y(n_340)
);

INVx2_ASAP7_75t_SL g341 ( 
.A(n_80),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_135),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_113),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_26),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g345 ( 
.A(n_24),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_2),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_47),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_74),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_29),
.Y(n_349)
);

BUFx3_ASAP7_75t_L g350 ( 
.A(n_192),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_19),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_31),
.Y(n_352)
);

INVxp33_ASAP7_75t_SL g353 ( 
.A(n_39),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_103),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_105),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_87),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_181),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_196),
.Y(n_358)
);

HB1xp67_ASAP7_75t_L g359 ( 
.A(n_38),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_125),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_21),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_63),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_50),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_112),
.Y(n_364)
);

CKINVDCx20_ASAP7_75t_R g365 ( 
.A(n_25),
.Y(n_365)
);

BUFx10_ASAP7_75t_L g366 ( 
.A(n_46),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_4),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_52),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_41),
.Y(n_369)
);

BUFx6f_ASAP7_75t_L g370 ( 
.A(n_151),
.Y(n_370)
);

INVx1_ASAP7_75t_SL g371 ( 
.A(n_183),
.Y(n_371)
);

CKINVDCx20_ASAP7_75t_R g372 ( 
.A(n_174),
.Y(n_372)
);

BUFx5_ASAP7_75t_L g373 ( 
.A(n_104),
.Y(n_373)
);

INVx2_ASAP7_75t_SL g374 ( 
.A(n_45),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_57),
.Y(n_375)
);

HB1xp67_ASAP7_75t_L g376 ( 
.A(n_195),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_26),
.Y(n_377)
);

INVxp67_ASAP7_75t_L g378 ( 
.A(n_131),
.Y(n_378)
);

CKINVDCx20_ASAP7_75t_R g379 ( 
.A(n_12),
.Y(n_379)
);

INVx1_ASAP7_75t_SL g380 ( 
.A(n_36),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_76),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_39),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_90),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_60),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_168),
.Y(n_385)
);

BUFx6f_ASAP7_75t_L g386 ( 
.A(n_186),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_56),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_175),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_24),
.Y(n_389)
);

CKINVDCx20_ASAP7_75t_R g390 ( 
.A(n_42),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_210),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_6),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_84),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_99),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_60),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_191),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_117),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_69),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_203),
.Y(n_399)
);

CKINVDCx20_ASAP7_75t_R g400 ( 
.A(n_158),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_0),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_67),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_86),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_11),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_120),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_215),
.Y(n_406)
);

CKINVDCx14_ASAP7_75t_R g407 ( 
.A(n_200),
.Y(n_407)
);

INVx1_ASAP7_75t_SL g408 ( 
.A(n_23),
.Y(n_408)
);

CKINVDCx20_ASAP7_75t_R g409 ( 
.A(n_212),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_65),
.Y(n_410)
);

BUFx3_ASAP7_75t_L g411 ( 
.A(n_218),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_58),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_44),
.Y(n_413)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_189),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_93),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_92),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_28),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_12),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_82),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_75),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_100),
.Y(n_421)
);

BUFx2_ASAP7_75t_SL g422 ( 
.A(n_41),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_122),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_69),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_3),
.Y(n_425)
);

INVx1_ASAP7_75t_SL g426 ( 
.A(n_96),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_172),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_204),
.Y(n_428)
);

INVxp33_ASAP7_75t_L g429 ( 
.A(n_190),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_72),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_18),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_85),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_94),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_145),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_21),
.Y(n_435)
);

HB1xp67_ASAP7_75t_L g436 ( 
.A(n_10),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_51),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_54),
.Y(n_438)
);

INVx1_ASAP7_75t_SL g439 ( 
.A(n_147),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_13),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_157),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_187),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_315),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_319),
.Y(n_444)
);

INVxp67_ASAP7_75t_SL g445 ( 
.A(n_234),
.Y(n_445)
);

CKINVDCx20_ASAP7_75t_R g446 ( 
.A(n_287),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_316),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_227),
.Y(n_448)
);

CKINVDCx20_ASAP7_75t_R g449 ( 
.A(n_300),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_309),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_227),
.Y(n_451)
);

INVx2_ASAP7_75t_L g452 ( 
.A(n_227),
.Y(n_452)
);

INVxp33_ASAP7_75t_L g453 ( 
.A(n_359),
.Y(n_453)
);

CKINVDCx20_ASAP7_75t_R g454 ( 
.A(n_321),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_227),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_227),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_339),
.Y(n_457)
);

HB1xp67_ASAP7_75t_L g458 ( 
.A(n_436),
.Y(n_458)
);

HB1xp67_ASAP7_75t_L g459 ( 
.A(n_308),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_372),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_339),
.Y(n_461)
);

INVxp67_ASAP7_75t_SL g462 ( 
.A(n_234),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_339),
.Y(n_463)
);

CKINVDCx5p33_ASAP7_75t_R g464 ( 
.A(n_400),
.Y(n_464)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_339),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_339),
.Y(n_466)
);

CKINVDCx16_ASAP7_75t_R g467 ( 
.A(n_407),
.Y(n_467)
);

HB1xp67_ASAP7_75t_L g468 ( 
.A(n_245),
.Y(n_468)
);

INVxp67_ASAP7_75t_L g469 ( 
.A(n_422),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_299),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_299),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_274),
.Y(n_472)
);

HB1xp67_ASAP7_75t_L g473 ( 
.A(n_245),
.Y(n_473)
);

CKINVDCx5p33_ASAP7_75t_R g474 ( 
.A(n_409),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_274),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_276),
.Y(n_476)
);

CKINVDCx5p33_ASAP7_75t_R g477 ( 
.A(n_266),
.Y(n_477)
);

INVxp67_ASAP7_75t_L g478 ( 
.A(n_374),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_276),
.Y(n_479)
);

CKINVDCx20_ASAP7_75t_R g480 ( 
.A(n_312),
.Y(n_480)
);

CKINVDCx16_ASAP7_75t_R g481 ( 
.A(n_237),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_292),
.Y(n_482)
);

CKINVDCx20_ASAP7_75t_R g483 ( 
.A(n_320),
.Y(n_483)
);

BUFx3_ASAP7_75t_L g484 ( 
.A(n_224),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_292),
.Y(n_485)
);

CKINVDCx5p33_ASAP7_75t_R g486 ( 
.A(n_270),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_414),
.Y(n_487)
);

CKINVDCx20_ASAP7_75t_R g488 ( 
.A(n_345),
.Y(n_488)
);

INVxp67_ASAP7_75t_SL g489 ( 
.A(n_235),
.Y(n_489)
);

CKINVDCx16_ASAP7_75t_R g490 ( 
.A(n_265),
.Y(n_490)
);

CKINVDCx20_ASAP7_75t_R g491 ( 
.A(n_365),
.Y(n_491)
);

CKINVDCx5p33_ASAP7_75t_R g492 ( 
.A(n_281),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_414),
.Y(n_493)
);

CKINVDCx20_ASAP7_75t_R g494 ( 
.A(n_379),
.Y(n_494)
);

BUFx6f_ASAP7_75t_L g495 ( 
.A(n_225),
.Y(n_495)
);

INVxp67_ASAP7_75t_SL g496 ( 
.A(n_260),
.Y(n_496)
);

INVxp33_ASAP7_75t_L g497 ( 
.A(n_261),
.Y(n_497)
);

CKINVDCx16_ASAP7_75t_R g498 ( 
.A(n_265),
.Y(n_498)
);

INVxp67_ASAP7_75t_SL g499 ( 
.A(n_264),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_273),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_275),
.Y(n_501)
);

INVx1_ASAP7_75t_SL g502 ( 
.A(n_390),
.Y(n_502)
);

HB1xp67_ASAP7_75t_L g503 ( 
.A(n_251),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_282),
.Y(n_504)
);

INVx3_ASAP7_75t_L g505 ( 
.A(n_237),
.Y(n_505)
);

BUFx3_ASAP7_75t_L g506 ( 
.A(n_224),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_286),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_226),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_332),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_337),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_346),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_347),
.Y(n_512)
);

INVxp67_ASAP7_75t_SL g513 ( 
.A(n_361),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_362),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_367),
.Y(n_515)
);

CKINVDCx5p33_ASAP7_75t_R g516 ( 
.A(n_285),
.Y(n_516)
);

CKINVDCx20_ASAP7_75t_R g517 ( 
.A(n_237),
.Y(n_517)
);

CKINVDCx5p33_ASAP7_75t_R g518 ( 
.A(n_288),
.Y(n_518)
);

INVx2_ASAP7_75t_L g519 ( 
.A(n_226),
.Y(n_519)
);

CKINVDCx5p33_ASAP7_75t_R g520 ( 
.A(n_293),
.Y(n_520)
);

INVxp33_ASAP7_75t_L g521 ( 
.A(n_369),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_377),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_384),
.Y(n_523)
);

CKINVDCx5p33_ASAP7_75t_R g524 ( 
.A(n_295),
.Y(n_524)
);

CKINVDCx20_ASAP7_75t_R g525 ( 
.A(n_268),
.Y(n_525)
);

CKINVDCx20_ASAP7_75t_R g526 ( 
.A(n_268),
.Y(n_526)
);

CKINVDCx5p33_ASAP7_75t_R g527 ( 
.A(n_303),
.Y(n_527)
);

INVxp67_ASAP7_75t_SL g528 ( 
.A(n_404),
.Y(n_528)
);

HB1xp67_ASAP7_75t_L g529 ( 
.A(n_251),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_410),
.Y(n_530)
);

CKINVDCx5p33_ASAP7_75t_R g531 ( 
.A(n_306),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_412),
.Y(n_532)
);

BUFx3_ASAP7_75t_L g533 ( 
.A(n_248),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_418),
.Y(n_534)
);

CKINVDCx5p33_ASAP7_75t_R g535 ( 
.A(n_317),
.Y(n_535)
);

CKINVDCx5p33_ASAP7_75t_R g536 ( 
.A(n_327),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_425),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_435),
.Y(n_538)
);

CKINVDCx5p33_ASAP7_75t_R g539 ( 
.A(n_336),
.Y(n_539)
);

INVx2_ASAP7_75t_L g540 ( 
.A(n_248),
.Y(n_540)
);

INVxp67_ASAP7_75t_SL g541 ( 
.A(n_440),
.Y(n_541)
);

CKINVDCx20_ASAP7_75t_R g542 ( 
.A(n_268),
.Y(n_542)
);

CKINVDCx20_ASAP7_75t_R g543 ( 
.A(n_269),
.Y(n_543)
);

BUFx3_ASAP7_75t_L g544 ( 
.A(n_350),
.Y(n_544)
);

CKINVDCx16_ASAP7_75t_R g545 ( 
.A(n_269),
.Y(n_545)
);

CKINVDCx20_ASAP7_75t_R g546 ( 
.A(n_269),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_229),
.Y(n_547)
);

CKINVDCx20_ASAP7_75t_R g548 ( 
.A(n_280),
.Y(n_548)
);

BUFx3_ASAP7_75t_L g549 ( 
.A(n_350),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_230),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_236),
.Y(n_551)
);

CKINVDCx5p33_ASAP7_75t_R g552 ( 
.A(n_344),
.Y(n_552)
);

CKINVDCx20_ASAP7_75t_R g553 ( 
.A(n_280),
.Y(n_553)
);

CKINVDCx5p33_ASAP7_75t_R g554 ( 
.A(n_349),
.Y(n_554)
);

INVx2_ASAP7_75t_L g555 ( 
.A(n_411),
.Y(n_555)
);

INVxp33_ASAP7_75t_SL g556 ( 
.A(n_258),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_241),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_244),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_247),
.Y(n_559)
);

CKINVDCx5p33_ASAP7_75t_R g560 ( 
.A(n_351),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_263),
.Y(n_561)
);

AND2x2_ASAP7_75t_L g562 ( 
.A(n_547),
.B(n_284),
.Y(n_562)
);

CKINVDCx5p33_ASAP7_75t_R g563 ( 
.A(n_450),
.Y(n_563)
);

AND2x2_ASAP7_75t_L g564 ( 
.A(n_547),
.B(n_297),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_L g565 ( 
.A(n_508),
.B(n_519),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_448),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_448),
.Y(n_567)
);

AND2x4_ASAP7_75t_L g568 ( 
.A(n_505),
.B(n_484),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_451),
.Y(n_569)
);

NAND2xp33_ASAP7_75t_L g570 ( 
.A(n_477),
.B(n_352),
.Y(n_570)
);

OA21x2_ASAP7_75t_L g571 ( 
.A1(n_451),
.A2(n_278),
.B(n_272),
.Y(n_571)
);

AND2x2_ASAP7_75t_L g572 ( 
.A(n_550),
.B(n_376),
.Y(n_572)
);

INVx3_ASAP7_75t_L g573 ( 
.A(n_452),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_495),
.Y(n_574)
);

INVx2_ASAP7_75t_L g575 ( 
.A(n_495),
.Y(n_575)
);

AND2x2_ASAP7_75t_L g576 ( 
.A(n_550),
.B(n_429),
.Y(n_576)
);

CKINVDCx20_ASAP7_75t_R g577 ( 
.A(n_480),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_495),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_455),
.Y(n_579)
);

INVx3_ASAP7_75t_L g580 ( 
.A(n_452),
.Y(n_580)
);

AOI22xp5_ASAP7_75t_L g581 ( 
.A1(n_517),
.A2(n_353),
.B1(n_311),
.B2(n_380),
.Y(n_581)
);

BUFx6f_ASAP7_75t_L g582 ( 
.A(n_495),
.Y(n_582)
);

CKINVDCx5p33_ASAP7_75t_R g583 ( 
.A(n_460),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_455),
.Y(n_584)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_495),
.Y(n_585)
);

AND2x4_ASAP7_75t_L g586 ( 
.A(n_551),
.B(n_279),
.Y(n_586)
);

OA21x2_ASAP7_75t_L g587 ( 
.A1(n_456),
.A2(n_461),
.B(n_457),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_456),
.Y(n_588)
);

AND2x4_ASAP7_75t_L g589 ( 
.A(n_505),
.B(n_411),
.Y(n_589)
);

OAI21x1_ASAP7_75t_L g590 ( 
.A1(n_465),
.A2(n_298),
.B(n_294),
.Y(n_590)
);

NOR2xp33_ASAP7_75t_L g591 ( 
.A(n_505),
.B(n_378),
.Y(n_591)
);

INVx3_ASAP7_75t_L g592 ( 
.A(n_465),
.Y(n_592)
);

NOR2xp67_ASAP7_75t_L g593 ( 
.A(n_551),
.B(n_279),
.Y(n_593)
);

BUFx12f_ASAP7_75t_L g594 ( 
.A(n_444),
.Y(n_594)
);

BUFx6f_ASAP7_75t_L g595 ( 
.A(n_457),
.Y(n_595)
);

AOI22xp5_ASAP7_75t_L g596 ( 
.A1(n_525),
.A2(n_542),
.B1(n_543),
.B2(n_526),
.Y(n_596)
);

INVx2_ASAP7_75t_L g597 ( 
.A(n_461),
.Y(n_597)
);

INVx2_ASAP7_75t_L g598 ( 
.A(n_463),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_463),
.Y(n_599)
);

INVx2_ASAP7_75t_L g600 ( 
.A(n_466),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_466),
.Y(n_601)
);

AND2x6_ASAP7_75t_L g602 ( 
.A(n_561),
.B(n_225),
.Y(n_602)
);

CKINVDCx5p33_ASAP7_75t_R g603 ( 
.A(n_464),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_472),
.Y(n_604)
);

BUFx6f_ASAP7_75t_L g605 ( 
.A(n_472),
.Y(n_605)
);

CKINVDCx5p33_ASAP7_75t_R g606 ( 
.A(n_474),
.Y(n_606)
);

INVx2_ASAP7_75t_L g607 ( 
.A(n_475),
.Y(n_607)
);

AND2x2_ASAP7_75t_L g608 ( 
.A(n_557),
.B(n_265),
.Y(n_608)
);

INVx2_ASAP7_75t_L g609 ( 
.A(n_475),
.Y(n_609)
);

INVxp67_ASAP7_75t_L g610 ( 
.A(n_468),
.Y(n_610)
);

HB1xp67_ASAP7_75t_L g611 ( 
.A(n_459),
.Y(n_611)
);

INVx3_ASAP7_75t_L g612 ( 
.A(n_476),
.Y(n_612)
);

BUFx6f_ASAP7_75t_L g613 ( 
.A(n_476),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_L g614 ( 
.A(n_508),
.B(n_302),
.Y(n_614)
);

INVx2_ASAP7_75t_L g615 ( 
.A(n_479),
.Y(n_615)
);

INVx3_ASAP7_75t_L g616 ( 
.A(n_479),
.Y(n_616)
);

BUFx6f_ASAP7_75t_L g617 ( 
.A(n_482),
.Y(n_617)
);

BUFx3_ASAP7_75t_L g618 ( 
.A(n_484),
.Y(n_618)
);

INVx2_ASAP7_75t_L g619 ( 
.A(n_482),
.Y(n_619)
);

INVx6_ASAP7_75t_L g620 ( 
.A(n_506),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_485),
.Y(n_621)
);

INVx2_ASAP7_75t_L g622 ( 
.A(n_485),
.Y(n_622)
);

HB1xp67_ASAP7_75t_L g623 ( 
.A(n_447),
.Y(n_623)
);

BUFx3_ASAP7_75t_L g624 ( 
.A(n_506),
.Y(n_624)
);

NOR2xp33_ASAP7_75t_L g625 ( 
.A(n_467),
.B(n_341),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_487),
.Y(n_626)
);

AND2x4_ASAP7_75t_L g627 ( 
.A(n_557),
.B(n_341),
.Y(n_627)
);

OAI22xp5_ASAP7_75t_L g628 ( 
.A1(n_453),
.A2(n_497),
.B1(n_521),
.B2(n_458),
.Y(n_628)
);

BUFx2_ASAP7_75t_L g629 ( 
.A(n_486),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_487),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_493),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_493),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_558),
.Y(n_633)
);

AND2x2_ASAP7_75t_SL g634 ( 
.A(n_481),
.B(n_225),
.Y(n_634)
);

CKINVDCx16_ASAP7_75t_R g635 ( 
.A(n_481),
.Y(n_635)
);

INVx3_ASAP7_75t_L g636 ( 
.A(n_519),
.Y(n_636)
);

AND2x2_ASAP7_75t_L g637 ( 
.A(n_558),
.B(n_366),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_559),
.Y(n_638)
);

BUFx2_ASAP7_75t_L g639 ( 
.A(n_492),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_559),
.Y(n_640)
);

INVx2_ASAP7_75t_L g641 ( 
.A(n_470),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_L g642 ( 
.A(n_540),
.B(n_305),
.Y(n_642)
);

CKINVDCx20_ASAP7_75t_R g643 ( 
.A(n_483),
.Y(n_643)
);

INVx2_ASAP7_75t_L g644 ( 
.A(n_470),
.Y(n_644)
);

INVx2_ASAP7_75t_L g645 ( 
.A(n_471),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_561),
.Y(n_646)
);

BUFx3_ASAP7_75t_L g647 ( 
.A(n_533),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_471),
.Y(n_648)
);

CKINVDCx5p33_ASAP7_75t_R g649 ( 
.A(n_446),
.Y(n_649)
);

BUFx6f_ASAP7_75t_L g650 ( 
.A(n_540),
.Y(n_650)
);

BUFx6f_ASAP7_75t_L g651 ( 
.A(n_555),
.Y(n_651)
);

CKINVDCx5p33_ASAP7_75t_R g652 ( 
.A(n_449),
.Y(n_652)
);

INVx3_ASAP7_75t_L g653 ( 
.A(n_555),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_L g654 ( 
.A(n_533),
.B(n_307),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_500),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_544),
.B(n_310),
.Y(n_656)
);

INVx2_ASAP7_75t_L g657 ( 
.A(n_587),
.Y(n_657)
);

INVx3_ASAP7_75t_L g658 ( 
.A(n_650),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_L g659 ( 
.A(n_591),
.B(n_467),
.Y(n_659)
);

INVx2_ASAP7_75t_L g660 ( 
.A(n_587),
.Y(n_660)
);

INVx2_ASAP7_75t_L g661 ( 
.A(n_587),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_SL g662 ( 
.A(n_634),
.B(n_516),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_566),
.Y(n_663)
);

BUFx10_ASAP7_75t_L g664 ( 
.A(n_625),
.Y(n_664)
);

INVxp67_ASAP7_75t_SL g665 ( 
.A(n_618),
.Y(n_665)
);

NOR2x1p5_ASAP7_75t_L g666 ( 
.A(n_594),
.B(n_443),
.Y(n_666)
);

NOR2xp33_ASAP7_75t_L g667 ( 
.A(n_618),
.B(n_545),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_566),
.Y(n_668)
);

AND2x2_ASAP7_75t_L g669 ( 
.A(n_608),
.B(n_445),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_SL g670 ( 
.A(n_634),
.B(n_518),
.Y(n_670)
);

INVx2_ASAP7_75t_L g671 ( 
.A(n_587),
.Y(n_671)
);

CKINVDCx5p33_ASAP7_75t_R g672 ( 
.A(n_563),
.Y(n_672)
);

INVx2_ASAP7_75t_L g673 ( 
.A(n_587),
.Y(n_673)
);

AOI22xp5_ASAP7_75t_L g674 ( 
.A1(n_634),
.A2(n_353),
.B1(n_408),
.B2(n_387),
.Y(n_674)
);

BUFx3_ASAP7_75t_L g675 ( 
.A(n_620),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_567),
.Y(n_676)
);

AOI22xp33_ASAP7_75t_SL g677 ( 
.A1(n_628),
.A2(n_545),
.B1(n_548),
.B2(n_546),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_567),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_SL g679 ( 
.A(n_608),
.B(n_520),
.Y(n_679)
);

BUFx3_ASAP7_75t_L g680 ( 
.A(n_620),
.Y(n_680)
);

BUFx10_ASAP7_75t_L g681 ( 
.A(n_568),
.Y(n_681)
);

BUFx6f_ASAP7_75t_L g682 ( 
.A(n_650),
.Y(n_682)
);

INVx2_ASAP7_75t_L g683 ( 
.A(n_597),
.Y(n_683)
);

INVxp67_ASAP7_75t_L g684 ( 
.A(n_629),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_569),
.Y(n_685)
);

INVx2_ASAP7_75t_L g686 ( 
.A(n_598),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_569),
.Y(n_687)
);

INVx2_ASAP7_75t_SL g688 ( 
.A(n_618),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_579),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_579),
.Y(n_690)
);

AOI22xp33_ASAP7_75t_L g691 ( 
.A1(n_586),
.A2(n_627),
.B1(n_562),
.B2(n_564),
.Y(n_691)
);

INVx2_ASAP7_75t_L g692 ( 
.A(n_598),
.Y(n_692)
);

INVx2_ASAP7_75t_L g693 ( 
.A(n_600),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_SL g694 ( 
.A(n_608),
.B(n_524),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_584),
.Y(n_695)
);

OA22x2_ASAP7_75t_L g696 ( 
.A1(n_581),
.A2(n_489),
.B1(n_499),
.B2(n_496),
.Y(n_696)
);

INVx2_ASAP7_75t_L g697 ( 
.A(n_600),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_L g698 ( 
.A(n_589),
.B(n_544),
.Y(n_698)
);

BUFx2_ASAP7_75t_L g699 ( 
.A(n_629),
.Y(n_699)
);

INVx2_ASAP7_75t_SL g700 ( 
.A(n_624),
.Y(n_700)
);

INVx2_ASAP7_75t_L g701 ( 
.A(n_600),
.Y(n_701)
);

BUFx6f_ASAP7_75t_L g702 ( 
.A(n_650),
.Y(n_702)
);

INVx2_ASAP7_75t_L g703 ( 
.A(n_605),
.Y(n_703)
);

BUFx10_ASAP7_75t_L g704 ( 
.A(n_568),
.Y(n_704)
);

CKINVDCx5p33_ASAP7_75t_R g705 ( 
.A(n_583),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_SL g706 ( 
.A(n_637),
.B(n_527),
.Y(n_706)
);

INVx2_ASAP7_75t_L g707 ( 
.A(n_605),
.Y(n_707)
);

INVx2_ASAP7_75t_L g708 ( 
.A(n_605),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_584),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_SL g710 ( 
.A(n_637),
.B(n_531),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_588),
.Y(n_711)
);

INVxp67_ASAP7_75t_L g712 ( 
.A(n_639),
.Y(n_712)
);

AND2x4_ASAP7_75t_L g713 ( 
.A(n_637),
.B(n_513),
.Y(n_713)
);

INVx2_ASAP7_75t_SL g714 ( 
.A(n_624),
.Y(n_714)
);

AOI22xp33_ASAP7_75t_L g715 ( 
.A1(n_586),
.A2(n_556),
.B1(n_503),
.B2(n_529),
.Y(n_715)
);

BUFx6f_ASAP7_75t_L g716 ( 
.A(n_650),
.Y(n_716)
);

INVx2_ASAP7_75t_L g717 ( 
.A(n_605),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_588),
.Y(n_718)
);

INVx3_ASAP7_75t_L g719 ( 
.A(n_650),
.Y(n_719)
);

INVx2_ASAP7_75t_L g720 ( 
.A(n_605),
.Y(n_720)
);

INVx3_ASAP7_75t_L g721 ( 
.A(n_650),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_599),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_599),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_601),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_601),
.Y(n_725)
);

BUFx6f_ASAP7_75t_L g726 ( 
.A(n_650),
.Y(n_726)
);

CKINVDCx5p33_ASAP7_75t_R g727 ( 
.A(n_603),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_SL g728 ( 
.A(n_568),
.B(n_535),
.Y(n_728)
);

INVx2_ASAP7_75t_L g729 ( 
.A(n_605),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_SL g730 ( 
.A(n_568),
.B(n_536),
.Y(n_730)
);

AND2x2_ASAP7_75t_L g731 ( 
.A(n_576),
.B(n_462),
.Y(n_731)
);

INVx2_ASAP7_75t_L g732 ( 
.A(n_605),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_613),
.Y(n_733)
);

BUFx3_ASAP7_75t_L g734 ( 
.A(n_620),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_613),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_613),
.Y(n_736)
);

INVx2_ASAP7_75t_L g737 ( 
.A(n_613),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_613),
.Y(n_738)
);

INVx2_ASAP7_75t_L g739 ( 
.A(n_613),
.Y(n_739)
);

NOR2xp33_ASAP7_75t_SL g740 ( 
.A(n_635),
.B(n_277),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_613),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_SL g742 ( 
.A(n_639),
.B(n_539),
.Y(n_742)
);

AOI22xp33_ASAP7_75t_L g743 ( 
.A1(n_586),
.A2(n_473),
.B1(n_541),
.B2(n_528),
.Y(n_743)
);

INVx2_ASAP7_75t_L g744 ( 
.A(n_617),
.Y(n_744)
);

BUFx6f_ASAP7_75t_L g745 ( 
.A(n_651),
.Y(n_745)
);

BUFx2_ASAP7_75t_L g746 ( 
.A(n_611),
.Y(n_746)
);

INVx2_ASAP7_75t_L g747 ( 
.A(n_617),
.Y(n_747)
);

INVx3_ASAP7_75t_L g748 ( 
.A(n_651),
.Y(n_748)
);

INVx4_ASAP7_75t_L g749 ( 
.A(n_651),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_L g750 ( 
.A(n_589),
.B(n_549),
.Y(n_750)
);

INVx4_ASAP7_75t_L g751 ( 
.A(n_651),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_617),
.Y(n_752)
);

CKINVDCx5p33_ASAP7_75t_R g753 ( 
.A(n_606),
.Y(n_753)
);

AND3x1_ASAP7_75t_L g754 ( 
.A(n_581),
.B(n_501),
.C(n_500),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_L g755 ( 
.A(n_589),
.B(n_552),
.Y(n_755)
);

INVx1_ASAP7_75t_SL g756 ( 
.A(n_577),
.Y(n_756)
);

OAI21xp33_ASAP7_75t_SL g757 ( 
.A1(n_562),
.A2(n_504),
.B(n_501),
.Y(n_757)
);

INVx3_ASAP7_75t_L g758 ( 
.A(n_651),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_617),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_SL g760 ( 
.A(n_576),
.B(n_554),
.Y(n_760)
);

INVx2_ASAP7_75t_L g761 ( 
.A(n_617),
.Y(n_761)
);

BUFx6f_ASAP7_75t_L g762 ( 
.A(n_651),
.Y(n_762)
);

INVx4_ASAP7_75t_L g763 ( 
.A(n_651),
.Y(n_763)
);

OR2x6_ASAP7_75t_L g764 ( 
.A(n_594),
.B(n_504),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_617),
.Y(n_765)
);

NOR2xp33_ASAP7_75t_L g766 ( 
.A(n_624),
.B(n_560),
.Y(n_766)
);

INVx2_ASAP7_75t_SL g767 ( 
.A(n_647),
.Y(n_767)
);

INVxp67_ASAP7_75t_L g768 ( 
.A(n_628),
.Y(n_768)
);

NOR2xp33_ASAP7_75t_L g769 ( 
.A(n_647),
.B(n_490),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_617),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_607),
.Y(n_771)
);

INVx2_ASAP7_75t_L g772 ( 
.A(n_595),
.Y(n_772)
);

BUFx4f_ASAP7_75t_L g773 ( 
.A(n_602),
.Y(n_773)
);

AND2x6_ASAP7_75t_L g774 ( 
.A(n_562),
.B(n_225),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_589),
.B(n_469),
.Y(n_775)
);

INVx2_ASAP7_75t_L g776 ( 
.A(n_595),
.Y(n_776)
);

OAI21xp5_ASAP7_75t_L g777 ( 
.A1(n_590),
.A2(n_325),
.B(n_323),
.Y(n_777)
);

INVx2_ASAP7_75t_SL g778 ( 
.A(n_647),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_607),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_586),
.B(n_498),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_607),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_SL g782 ( 
.A(n_576),
.B(n_228),
.Y(n_782)
);

INVx3_ASAP7_75t_L g783 ( 
.A(n_595),
.Y(n_783)
);

INVx2_ASAP7_75t_L g784 ( 
.A(n_595),
.Y(n_784)
);

INVx4_ASAP7_75t_L g785 ( 
.A(n_602),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_SL g786 ( 
.A(n_564),
.B(n_228),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_609),
.Y(n_787)
);

BUFx6f_ASAP7_75t_L g788 ( 
.A(n_595),
.Y(n_788)
);

AOI22xp5_ASAP7_75t_L g789 ( 
.A1(n_564),
.A2(n_387),
.B1(n_389),
.B2(n_258),
.Y(n_789)
);

CKINVDCx5p33_ASAP7_75t_R g790 ( 
.A(n_649),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_L g791 ( 
.A(n_627),
.B(n_507),
.Y(n_791)
);

INVx3_ASAP7_75t_L g792 ( 
.A(n_595),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_609),
.Y(n_793)
);

AND3x2_ASAP7_75t_L g794 ( 
.A(n_623),
.B(n_478),
.C(n_290),
.Y(n_794)
);

INVx2_ASAP7_75t_L g795 ( 
.A(n_595),
.Y(n_795)
);

INVx3_ASAP7_75t_L g796 ( 
.A(n_612),
.Y(n_796)
);

INVx2_ASAP7_75t_L g797 ( 
.A(n_609),
.Y(n_797)
);

INVx3_ASAP7_75t_L g798 ( 
.A(n_612),
.Y(n_798)
);

INVx2_ASAP7_75t_L g799 ( 
.A(n_615),
.Y(n_799)
);

INVx2_ASAP7_75t_L g800 ( 
.A(n_615),
.Y(n_800)
);

AND2x2_ASAP7_75t_L g801 ( 
.A(n_572),
.B(n_507),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_SL g802 ( 
.A(n_610),
.B(n_231),
.Y(n_802)
);

INVx2_ASAP7_75t_L g803 ( 
.A(n_615),
.Y(n_803)
);

INVx3_ASAP7_75t_L g804 ( 
.A(n_612),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_619),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_619),
.Y(n_806)
);

INVx2_ASAP7_75t_L g807 ( 
.A(n_619),
.Y(n_807)
);

INVx5_ASAP7_75t_L g808 ( 
.A(n_602),
.Y(n_808)
);

INVx2_ASAP7_75t_L g809 ( 
.A(n_622),
.Y(n_809)
);

INVx2_ASAP7_75t_L g810 ( 
.A(n_622),
.Y(n_810)
);

INVx2_ASAP7_75t_L g811 ( 
.A(n_622),
.Y(n_811)
);

BUFx6f_ASAP7_75t_SL g812 ( 
.A(n_627),
.Y(n_812)
);

AOI22xp33_ASAP7_75t_L g813 ( 
.A1(n_627),
.A2(n_553),
.B1(n_366),
.B2(n_537),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_L g814 ( 
.A(n_713),
.B(n_572),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_SL g815 ( 
.A(n_713),
.B(n_610),
.Y(n_815)
);

NOR2xp33_ASAP7_75t_L g816 ( 
.A(n_659),
.B(n_620),
.Y(n_816)
);

NAND2xp33_ASAP7_75t_SL g817 ( 
.A(n_672),
.B(n_623),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_L g818 ( 
.A(n_713),
.B(n_572),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_663),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_SL g820 ( 
.A(n_713),
.B(n_635),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_L g821 ( 
.A(n_669),
.B(n_627),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_L g822 ( 
.A(n_669),
.B(n_633),
.Y(n_822)
);

INVx3_ASAP7_75t_L g823 ( 
.A(n_681),
.Y(n_823)
);

NOR2xp33_ASAP7_75t_L g824 ( 
.A(n_662),
.B(n_620),
.Y(n_824)
);

AO22x2_ASAP7_75t_L g825 ( 
.A1(n_768),
.A2(n_502),
.B1(n_621),
.B2(n_604),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_663),
.Y(n_826)
);

NOR2xp33_ASAP7_75t_L g827 ( 
.A(n_670),
.B(n_570),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_668),
.Y(n_828)
);

INVx8_ASAP7_75t_L g829 ( 
.A(n_764),
.Y(n_829)
);

AND2x2_ASAP7_75t_L g830 ( 
.A(n_699),
.B(n_684),
.Y(n_830)
);

AND2x4_ASAP7_75t_L g831 ( 
.A(n_764),
.B(n_633),
.Y(n_831)
);

OAI22xp33_ASAP7_75t_L g832 ( 
.A1(n_674),
.A2(n_640),
.B1(n_646),
.B2(n_638),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_SL g833 ( 
.A(n_681),
.B(n_638),
.Y(n_833)
);

CKINVDCx5p33_ASAP7_75t_R g834 ( 
.A(n_672),
.Y(n_834)
);

OAI22xp5_ASAP7_75t_L g835 ( 
.A1(n_674),
.A2(n_646),
.B1(n_640),
.B2(n_655),
.Y(n_835)
);

INVxp67_ASAP7_75t_L g836 ( 
.A(n_746),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_676),
.Y(n_837)
);

OAI221xp5_ASAP7_75t_L g838 ( 
.A1(n_691),
.A2(n_656),
.B1(n_654),
.B2(n_655),
.C(n_401),
.Y(n_838)
);

BUFx6f_ASAP7_75t_L g839 ( 
.A(n_675),
.Y(n_839)
);

INVx2_ASAP7_75t_SL g840 ( 
.A(n_746),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_676),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_SL g842 ( 
.A(n_681),
.B(n_612),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_766),
.B(n_654),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_678),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_678),
.Y(n_845)
);

AOI22xp5_ASAP7_75t_L g846 ( 
.A1(n_812),
.A2(n_593),
.B1(n_656),
.B2(n_616),
.Y(n_846)
);

NAND2xp33_ASAP7_75t_L g847 ( 
.A(n_796),
.B(n_602),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_685),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_SL g849 ( 
.A(n_664),
.B(n_593),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_731),
.B(n_636),
.Y(n_850)
);

BUFx12f_ASAP7_75t_L g851 ( 
.A(n_790),
.Y(n_851)
);

INVx2_ASAP7_75t_L g852 ( 
.A(n_683),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_685),
.Y(n_853)
);

INVx2_ASAP7_75t_L g854 ( 
.A(n_683),
.Y(n_854)
);

AOI22xp5_ASAP7_75t_L g855 ( 
.A1(n_812),
.A2(n_616),
.B1(n_621),
.B2(n_604),
.Y(n_855)
);

NAND2xp33_ASAP7_75t_SL g856 ( 
.A(n_705),
.B(n_389),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_SL g857 ( 
.A(n_664),
.B(n_594),
.Y(n_857)
);

INVx4_ASAP7_75t_L g858 ( 
.A(n_681),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_687),
.Y(n_859)
);

NOR2xp33_ASAP7_75t_L g860 ( 
.A(n_664),
.B(n_565),
.Y(n_860)
);

NOR2xp33_ASAP7_75t_L g861 ( 
.A(n_664),
.B(n_565),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_731),
.B(n_796),
.Y(n_862)
);

NOR2xp33_ASAP7_75t_L g863 ( 
.A(n_755),
.B(n_614),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_796),
.B(n_636),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_798),
.B(n_636),
.Y(n_865)
);

BUFx2_ASAP7_75t_L g866 ( 
.A(n_790),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_687),
.Y(n_867)
);

O2A1O1Ixp33_ASAP7_75t_L g868 ( 
.A1(n_757),
.A2(n_616),
.B(n_630),
.C(n_626),
.Y(n_868)
);

NAND2xp33_ASAP7_75t_L g869 ( 
.A(n_798),
.B(n_602),
.Y(n_869)
);

OAI221xp5_ASAP7_75t_L g870 ( 
.A1(n_757),
.A2(n_401),
.B1(n_438),
.B2(n_398),
.C(n_395),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_SL g871 ( 
.A(n_704),
.B(n_798),
.Y(n_871)
);

INVx3_ASAP7_75t_L g872 ( 
.A(n_704),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_804),
.B(n_636),
.Y(n_873)
);

BUFx2_ASAP7_75t_L g874 ( 
.A(n_756),
.Y(n_874)
);

NOR2xp33_ASAP7_75t_L g875 ( 
.A(n_760),
.B(n_614),
.Y(n_875)
);

INVx8_ASAP7_75t_L g876 ( 
.A(n_764),
.Y(n_876)
);

NOR2xp33_ASAP7_75t_L g877 ( 
.A(n_679),
.B(n_694),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_804),
.B(n_653),
.Y(n_878)
);

AO22x2_ASAP7_75t_L g879 ( 
.A1(n_754),
.A2(n_626),
.B1(n_631),
.B2(n_630),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_SL g880 ( 
.A(n_704),
.B(n_231),
.Y(n_880)
);

INVx2_ASAP7_75t_L g881 ( 
.A(n_686),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_SL g882 ( 
.A(n_704),
.B(n_232),
.Y(n_882)
);

AND2x6_ASAP7_75t_SL g883 ( 
.A(n_764),
.B(n_705),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_SL g884 ( 
.A(n_804),
.B(n_616),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_L g885 ( 
.A(n_801),
.B(n_653),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_L g886 ( 
.A(n_801),
.B(n_653),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_689),
.Y(n_887)
);

AOI22xp5_ASAP7_75t_L g888 ( 
.A1(n_812),
.A2(n_632),
.B1(n_631),
.B2(n_232),
.Y(n_888)
);

AOI22xp33_ASAP7_75t_L g889 ( 
.A1(n_696),
.A2(n_571),
.B1(n_632),
.B2(n_641),
.Y(n_889)
);

INVx2_ASAP7_75t_L g890 ( 
.A(n_686),
.Y(n_890)
);

INVxp67_ASAP7_75t_L g891 ( 
.A(n_667),
.Y(n_891)
);

INVxp67_ASAP7_75t_L g892 ( 
.A(n_740),
.Y(n_892)
);

NOR2xp67_ASAP7_75t_L g893 ( 
.A(n_727),
.B(n_653),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_L g894 ( 
.A(n_774),
.B(n_642),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_SL g895 ( 
.A(n_788),
.B(n_233),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_SL g896 ( 
.A(n_712),
.B(n_233),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_L g897 ( 
.A(n_774),
.B(n_642),
.Y(n_897)
);

NOR2x1p5_ASAP7_75t_L g898 ( 
.A(n_727),
.B(n_652),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_SL g899 ( 
.A(n_780),
.B(n_238),
.Y(n_899)
);

AND2x2_ASAP7_75t_L g900 ( 
.A(n_789),
.B(n_596),
.Y(n_900)
);

AND2x4_ASAP7_75t_L g901 ( 
.A(n_764),
.B(n_728),
.Y(n_901)
);

BUFx6f_ASAP7_75t_SL g902 ( 
.A(n_774),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_689),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_774),
.B(n_648),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_690),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_L g906 ( 
.A(n_774),
.B(n_648),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_SL g907 ( 
.A(n_775),
.B(n_238),
.Y(n_907)
);

AOI22xp5_ASAP7_75t_L g908 ( 
.A1(n_774),
.A2(n_239),
.B1(n_242),
.B2(n_240),
.Y(n_908)
);

AND2x2_ASAP7_75t_L g909 ( 
.A(n_789),
.B(n_596),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_L g910 ( 
.A(n_774),
.B(n_641),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_L g911 ( 
.A(n_698),
.B(n_641),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_SL g912 ( 
.A(n_769),
.B(n_239),
.Y(n_912)
);

NAND2xp33_ASAP7_75t_SL g913 ( 
.A(n_753),
.B(n_392),
.Y(n_913)
);

OR2x2_ASAP7_75t_L g914 ( 
.A(n_753),
.B(n_643),
.Y(n_914)
);

CKINVDCx5p33_ASAP7_75t_R g915 ( 
.A(n_666),
.Y(n_915)
);

AO22x2_ASAP7_75t_L g916 ( 
.A1(n_754),
.A2(n_454),
.B1(n_510),
.B2(n_509),
.Y(n_916)
);

INVx2_ASAP7_75t_SL g917 ( 
.A(n_794),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_690),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_L g919 ( 
.A(n_750),
.B(n_644),
.Y(n_919)
);

NOR2xp33_ASAP7_75t_L g920 ( 
.A(n_706),
.B(n_363),
.Y(n_920)
);

NOR2xp33_ASAP7_75t_L g921 ( 
.A(n_710),
.B(n_368),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_L g922 ( 
.A(n_791),
.B(n_644),
.Y(n_922)
);

BUFx6f_ASAP7_75t_L g923 ( 
.A(n_675),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_695),
.Y(n_924)
);

A2O1A1Ixp33_ASAP7_75t_L g925 ( 
.A1(n_777),
.A2(n_590),
.B(n_645),
.C(n_644),
.Y(n_925)
);

NOR2xp33_ASAP7_75t_L g926 ( 
.A(n_782),
.B(n_375),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_L g927 ( 
.A(n_688),
.B(n_645),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_L g928 ( 
.A(n_688),
.B(n_645),
.Y(n_928)
);

INVx2_ASAP7_75t_L g929 ( 
.A(n_692),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_700),
.B(n_573),
.Y(n_930)
);

CKINVDCx5p33_ASAP7_75t_R g931 ( 
.A(n_666),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_695),
.Y(n_932)
);

INVxp67_ASAP7_75t_L g933 ( 
.A(n_740),
.Y(n_933)
);

BUFx3_ASAP7_75t_L g934 ( 
.A(n_700),
.Y(n_934)
);

NOR2xp33_ASAP7_75t_L g935 ( 
.A(n_730),
.B(n_382),
.Y(n_935)
);

INVx3_ASAP7_75t_L g936 ( 
.A(n_675),
.Y(n_936)
);

NOR2xp33_ASAP7_75t_L g937 ( 
.A(n_786),
.B(n_802),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_SL g938 ( 
.A(n_743),
.B(n_242),
.Y(n_938)
);

INVx2_ASAP7_75t_L g939 ( 
.A(n_693),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_SL g940 ( 
.A(n_788),
.B(n_243),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_709),
.Y(n_941)
);

A2O1A1Ixp33_ASAP7_75t_L g942 ( 
.A1(n_709),
.A2(n_590),
.B(n_423),
.C(n_420),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_L g943 ( 
.A(n_714),
.B(n_573),
.Y(n_943)
);

AND2x2_ASAP7_75t_L g944 ( 
.A(n_715),
.B(n_488),
.Y(n_944)
);

AND2x2_ASAP7_75t_L g945 ( 
.A(n_677),
.B(n_491),
.Y(n_945)
);

INVx2_ASAP7_75t_L g946 ( 
.A(n_693),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_L g947 ( 
.A(n_714),
.B(n_573),
.Y(n_947)
);

NAND2x1p5_ASAP7_75t_L g948 ( 
.A(n_785),
.B(n_571),
.Y(n_948)
);

OAI22xp33_ASAP7_75t_L g949 ( 
.A1(n_696),
.A2(n_438),
.B1(n_392),
.B2(n_395),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_L g950 ( 
.A(n_767),
.B(n_573),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_711),
.Y(n_951)
);

INVx1_ASAP7_75t_SL g952 ( 
.A(n_742),
.Y(n_952)
);

INVx8_ASAP7_75t_L g953 ( 
.A(n_808),
.Y(n_953)
);

NOR3xp33_ASAP7_75t_L g954 ( 
.A(n_718),
.B(n_398),
.C(n_402),
.Y(n_954)
);

INVx1_ASAP7_75t_L g955 ( 
.A(n_718),
.Y(n_955)
);

NOR2xp33_ASAP7_75t_L g956 ( 
.A(n_665),
.B(n_413),
.Y(n_956)
);

NOR2xp33_ASAP7_75t_L g957 ( 
.A(n_767),
.B(n_417),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_L g958 ( 
.A(n_778),
.B(n_580),
.Y(n_958)
);

AOI22xp33_ASAP7_75t_L g959 ( 
.A1(n_696),
.A2(n_571),
.B1(n_602),
.B2(n_366),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_722),
.Y(n_960)
);

INVx3_ASAP7_75t_L g961 ( 
.A(n_680),
.Y(n_961)
);

AND2x2_ASAP7_75t_SL g962 ( 
.A(n_773),
.B(n_571),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_SL g963 ( 
.A(n_778),
.B(n_243),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_L g964 ( 
.A(n_771),
.B(n_580),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_SL g965 ( 
.A(n_813),
.B(n_246),
.Y(n_965)
);

INVx2_ASAP7_75t_L g966 ( 
.A(n_697),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_L g967 ( 
.A(n_771),
.B(n_580),
.Y(n_967)
);

BUFx3_ASAP7_75t_L g968 ( 
.A(n_779),
.Y(n_968)
);

OAI221xp5_ASAP7_75t_L g969 ( 
.A1(n_722),
.A2(n_424),
.B1(n_431),
.B2(n_437),
.C(n_509),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_SL g970 ( 
.A(n_788),
.B(n_682),
.Y(n_970)
);

AO22x2_ASAP7_75t_L g971 ( 
.A1(n_657),
.A2(n_538),
.B1(n_515),
.B2(n_514),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_L g972 ( 
.A(n_779),
.B(n_580),
.Y(n_972)
);

AND2x2_ASAP7_75t_L g973 ( 
.A(n_781),
.B(n_494),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_723),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_L g975 ( 
.A(n_781),
.B(n_592),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_L g976 ( 
.A(n_787),
.B(n_592),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_723),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_819),
.Y(n_978)
);

OAI22x1_ASAP7_75t_L g979 ( 
.A1(n_900),
.A2(n_511),
.B1(n_512),
.B2(n_510),
.Y(n_979)
);

AND2x2_ASAP7_75t_L g980 ( 
.A(n_830),
.B(n_511),
.Y(n_980)
);

INVx1_ASAP7_75t_L g981 ( 
.A(n_826),
.Y(n_981)
);

NOR2xp33_ASAP7_75t_L g982 ( 
.A(n_891),
.B(n_724),
.Y(n_982)
);

CKINVDCx14_ASAP7_75t_R g983 ( 
.A(n_834),
.Y(n_983)
);

INVx5_ASAP7_75t_L g984 ( 
.A(n_953),
.Y(n_984)
);

INVx8_ASAP7_75t_L g985 ( 
.A(n_829),
.Y(n_985)
);

AND2x6_ASAP7_75t_SL g986 ( 
.A(n_909),
.B(n_512),
.Y(n_986)
);

OAI21xp5_ASAP7_75t_L g987 ( 
.A1(n_925),
.A2(n_660),
.B(n_657),
.Y(n_987)
);

OAI21xp5_ASAP7_75t_L g988 ( 
.A1(n_942),
.A2(n_661),
.B(n_660),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_L g989 ( 
.A(n_863),
.B(n_787),
.Y(n_989)
);

CKINVDCx5p33_ASAP7_75t_R g990 ( 
.A(n_851),
.Y(n_990)
);

INVx1_ASAP7_75t_L g991 ( 
.A(n_828),
.Y(n_991)
);

BUFx6f_ASAP7_75t_L g992 ( 
.A(n_839),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_L g993 ( 
.A(n_863),
.B(n_793),
.Y(n_993)
);

AOI221xp5_ASAP7_75t_L g994 ( 
.A1(n_832),
.A2(n_514),
.B1(n_515),
.B2(n_522),
.C(n_523),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_L g995 ( 
.A(n_843),
.B(n_793),
.Y(n_995)
);

INVx2_ASAP7_75t_L g996 ( 
.A(n_968),
.Y(n_996)
);

CKINVDCx5p33_ASAP7_75t_R g997 ( 
.A(n_866),
.Y(n_997)
);

BUFx8_ASAP7_75t_L g998 ( 
.A(n_874),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_L g999 ( 
.A(n_862),
.B(n_805),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_L g1000 ( 
.A(n_837),
.B(n_805),
.Y(n_1000)
);

INVx1_ASAP7_75t_L g1001 ( 
.A(n_841),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_L g1002 ( 
.A(n_844),
.B(n_806),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_L g1003 ( 
.A(n_845),
.B(n_806),
.Y(n_1003)
);

OR2x2_ASAP7_75t_L g1004 ( 
.A(n_840),
.B(n_522),
.Y(n_1004)
);

INVx2_ASAP7_75t_SL g1005 ( 
.A(n_914),
.Y(n_1005)
);

O2A1O1Ixp33_ASAP7_75t_L g1006 ( 
.A1(n_822),
.A2(n_725),
.B(n_724),
.C(n_797),
.Y(n_1006)
);

HB1xp67_ASAP7_75t_L g1007 ( 
.A(n_836),
.Y(n_1007)
);

CKINVDCx11_ASAP7_75t_R g1008 ( 
.A(n_883),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_SL g1009 ( 
.A(n_831),
.B(n_891),
.Y(n_1009)
);

INVx5_ASAP7_75t_L g1010 ( 
.A(n_953),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_L g1011 ( 
.A(n_848),
.B(n_797),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_SL g1012 ( 
.A(n_831),
.B(n_788),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_SL g1013 ( 
.A(n_832),
.B(n_788),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_L g1014 ( 
.A(n_853),
.B(n_799),
.Y(n_1014)
);

NOR2xp33_ASAP7_75t_L g1015 ( 
.A(n_836),
.B(n_725),
.Y(n_1015)
);

CKINVDCx20_ASAP7_75t_R g1016 ( 
.A(n_817),
.Y(n_1016)
);

INVx1_ASAP7_75t_L g1017 ( 
.A(n_859),
.Y(n_1017)
);

INVx5_ASAP7_75t_L g1018 ( 
.A(n_953),
.Y(n_1018)
);

NOR2x1p5_ASAP7_75t_L g1019 ( 
.A(n_915),
.B(n_523),
.Y(n_1019)
);

INVx1_ASAP7_75t_L g1020 ( 
.A(n_867),
.Y(n_1020)
);

INVx3_ASAP7_75t_L g1021 ( 
.A(n_858),
.Y(n_1021)
);

INVx2_ASAP7_75t_SL g1022 ( 
.A(n_973),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_L g1023 ( 
.A(n_887),
.B(n_799),
.Y(n_1023)
);

NOR2x2_ASAP7_75t_L g1024 ( 
.A(n_856),
.B(n_800),
.Y(n_1024)
);

NAND2x1_ASAP7_75t_L g1025 ( 
.A(n_858),
.B(n_783),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_SL g1026 ( 
.A(n_827),
.B(n_682),
.Y(n_1026)
);

AND2x2_ASAP7_75t_L g1027 ( 
.A(n_814),
.B(n_530),
.Y(n_1027)
);

AOI22xp5_ASAP7_75t_L g1028 ( 
.A1(n_877),
.A2(n_735),
.B1(n_736),
.B2(n_733),
.Y(n_1028)
);

BUFx8_ASAP7_75t_SL g1029 ( 
.A(n_931),
.Y(n_1029)
);

AND2x2_ASAP7_75t_L g1030 ( 
.A(n_818),
.B(n_530),
.Y(n_1030)
);

CKINVDCx20_ASAP7_75t_R g1031 ( 
.A(n_913),
.Y(n_1031)
);

BUFx3_ASAP7_75t_L g1032 ( 
.A(n_917),
.Y(n_1032)
);

BUFx2_ASAP7_75t_L g1033 ( 
.A(n_892),
.Y(n_1033)
);

INVx1_ASAP7_75t_L g1034 ( 
.A(n_903),
.Y(n_1034)
);

HB1xp67_ASAP7_75t_L g1035 ( 
.A(n_892),
.Y(n_1035)
);

INVx2_ASAP7_75t_SL g1036 ( 
.A(n_898),
.Y(n_1036)
);

AND2x2_ASAP7_75t_L g1037 ( 
.A(n_815),
.B(n_532),
.Y(n_1037)
);

INVx1_ASAP7_75t_L g1038 ( 
.A(n_905),
.Y(n_1038)
);

AOI21xp5_ASAP7_75t_L g1039 ( 
.A1(n_970),
.A2(n_735),
.B(n_733),
.Y(n_1039)
);

INVx2_ASAP7_75t_SL g1040 ( 
.A(n_829),
.Y(n_1040)
);

BUFx6f_ASAP7_75t_L g1041 ( 
.A(n_839),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_918),
.Y(n_1042)
);

NAND2xp5_ASAP7_75t_L g1043 ( 
.A(n_924),
.B(n_800),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_L g1044 ( 
.A(n_932),
.B(n_803),
.Y(n_1044)
);

BUFx2_ASAP7_75t_L g1045 ( 
.A(n_933),
.Y(n_1045)
);

INVx3_ASAP7_75t_L g1046 ( 
.A(n_823),
.Y(n_1046)
);

BUFx3_ASAP7_75t_L g1047 ( 
.A(n_944),
.Y(n_1047)
);

NOR2xp33_ASAP7_75t_L g1048 ( 
.A(n_933),
.B(n_749),
.Y(n_1048)
);

NOR2xp67_ASAP7_75t_L g1049 ( 
.A(n_857),
.B(n_803),
.Y(n_1049)
);

BUFx3_ASAP7_75t_L g1050 ( 
.A(n_952),
.Y(n_1050)
);

NAND2xp5_ASAP7_75t_SL g1051 ( 
.A(n_827),
.B(n_682),
.Y(n_1051)
);

NOR3xp33_ASAP7_75t_SL g1052 ( 
.A(n_870),
.B(n_250),
.C(n_246),
.Y(n_1052)
);

INVx1_ASAP7_75t_L g1053 ( 
.A(n_941),
.Y(n_1053)
);

INVx5_ASAP7_75t_L g1054 ( 
.A(n_823),
.Y(n_1054)
);

BUFx6f_ASAP7_75t_L g1055 ( 
.A(n_839),
.Y(n_1055)
);

BUFx6f_ASAP7_75t_L g1056 ( 
.A(n_839),
.Y(n_1056)
);

INVx4_ASAP7_75t_L g1057 ( 
.A(n_829),
.Y(n_1057)
);

AOI22xp33_ASAP7_75t_L g1058 ( 
.A1(n_916),
.A2(n_809),
.B1(n_810),
.B2(n_807),
.Y(n_1058)
);

AOI22xp33_ASAP7_75t_L g1059 ( 
.A1(n_916),
.A2(n_809),
.B1(n_810),
.B2(n_807),
.Y(n_1059)
);

AOI22xp5_ASAP7_75t_L g1060 ( 
.A1(n_877),
.A2(n_738),
.B1(n_741),
.B2(n_736),
.Y(n_1060)
);

NOR2xp67_ASAP7_75t_L g1061 ( 
.A(n_956),
.B(n_811),
.Y(n_1061)
);

AOI22xp5_ASAP7_75t_L g1062 ( 
.A1(n_901),
.A2(n_741),
.B1(n_752),
.B2(n_738),
.Y(n_1062)
);

AND2x4_ASAP7_75t_L g1063 ( 
.A(n_901),
.B(n_680),
.Y(n_1063)
);

AOI22xp33_ASAP7_75t_L g1064 ( 
.A1(n_916),
.A2(n_811),
.B1(n_661),
.B2(n_673),
.Y(n_1064)
);

NAND2xp5_ASAP7_75t_L g1065 ( 
.A(n_951),
.B(n_671),
.Y(n_1065)
);

INVx1_ASAP7_75t_L g1066 ( 
.A(n_955),
.Y(n_1066)
);

INVx1_ASAP7_75t_L g1067 ( 
.A(n_960),
.Y(n_1067)
);

NOR2x2_ASAP7_75t_L g1068 ( 
.A(n_954),
.B(n_703),
.Y(n_1068)
);

NAND2xp5_ASAP7_75t_L g1069 ( 
.A(n_974),
.B(n_671),
.Y(n_1069)
);

INVx1_ASAP7_75t_L g1070 ( 
.A(n_977),
.Y(n_1070)
);

INVx1_ASAP7_75t_L g1071 ( 
.A(n_885),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_SL g1072 ( 
.A(n_860),
.B(n_682),
.Y(n_1072)
);

NAND2xp5_ASAP7_75t_SL g1073 ( 
.A(n_860),
.B(n_682),
.Y(n_1073)
);

BUFx6f_ASAP7_75t_L g1074 ( 
.A(n_923),
.Y(n_1074)
);

NAND2xp5_ASAP7_75t_SL g1075 ( 
.A(n_861),
.B(n_702),
.Y(n_1075)
);

AND2x2_ASAP7_75t_L g1076 ( 
.A(n_945),
.B(n_532),
.Y(n_1076)
);

INVx5_ASAP7_75t_L g1077 ( 
.A(n_872),
.Y(n_1077)
);

OAI22xp5_ASAP7_75t_SL g1078 ( 
.A1(n_920),
.A2(n_537),
.B1(n_538),
.B2(n_534),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_L g1079 ( 
.A(n_861),
.B(n_821),
.Y(n_1079)
);

AND2x6_ASAP7_75t_L g1080 ( 
.A(n_872),
.B(n_673),
.Y(n_1080)
);

INVx1_ASAP7_75t_L g1081 ( 
.A(n_886),
.Y(n_1081)
);

INVx1_ASAP7_75t_L g1082 ( 
.A(n_850),
.Y(n_1082)
);

INVx1_ASAP7_75t_L g1083 ( 
.A(n_864),
.Y(n_1083)
);

NAND2xp5_ASAP7_75t_L g1084 ( 
.A(n_875),
.B(n_697),
.Y(n_1084)
);

INVx1_ASAP7_75t_L g1085 ( 
.A(n_865),
.Y(n_1085)
);

NAND2xp5_ASAP7_75t_L g1086 ( 
.A(n_875),
.B(n_701),
.Y(n_1086)
);

NAND2xp5_ASAP7_75t_SL g1087 ( 
.A(n_888),
.B(n_702),
.Y(n_1087)
);

INVx1_ASAP7_75t_L g1088 ( 
.A(n_873),
.Y(n_1088)
);

NAND2xp33_ASAP7_75t_SL g1089 ( 
.A(n_912),
.B(n_783),
.Y(n_1089)
);

AOI22xp33_ASAP7_75t_SL g1090 ( 
.A1(n_879),
.A2(n_534),
.B1(n_439),
.B2(n_371),
.Y(n_1090)
);

NAND2xp5_ASAP7_75t_L g1091 ( 
.A(n_816),
.B(n_701),
.Y(n_1091)
);

AND2x2_ASAP7_75t_L g1092 ( 
.A(n_820),
.B(n_571),
.Y(n_1092)
);

BUFx6f_ASAP7_75t_L g1093 ( 
.A(n_923),
.Y(n_1093)
);

INVx1_ASAP7_75t_L g1094 ( 
.A(n_878),
.Y(n_1094)
);

NAND2xp5_ASAP7_75t_L g1095 ( 
.A(n_816),
.B(n_752),
.Y(n_1095)
);

AND2x4_ASAP7_75t_L g1096 ( 
.A(n_893),
.B(n_680),
.Y(n_1096)
);

INVx2_ASAP7_75t_L g1097 ( 
.A(n_852),
.Y(n_1097)
);

INVx2_ASAP7_75t_SL g1098 ( 
.A(n_876),
.Y(n_1098)
);

NAND2xp5_ASAP7_75t_L g1099 ( 
.A(n_922),
.B(n_759),
.Y(n_1099)
);

CKINVDCx20_ASAP7_75t_R g1100 ( 
.A(n_876),
.Y(n_1100)
);

OR2x2_ASAP7_75t_SL g1101 ( 
.A(n_965),
.B(n_326),
.Y(n_1101)
);

INVx1_ASAP7_75t_L g1102 ( 
.A(n_964),
.Y(n_1102)
);

INVx3_ASAP7_75t_L g1103 ( 
.A(n_923),
.Y(n_1103)
);

INVx1_ASAP7_75t_L g1104 ( 
.A(n_967),
.Y(n_1104)
);

NAND2xp5_ASAP7_75t_L g1105 ( 
.A(n_879),
.B(n_759),
.Y(n_1105)
);

INVx2_ASAP7_75t_L g1106 ( 
.A(n_854),
.Y(n_1106)
);

INVx3_ASAP7_75t_L g1107 ( 
.A(n_923),
.Y(n_1107)
);

INVx1_ASAP7_75t_L g1108 ( 
.A(n_972),
.Y(n_1108)
);

INVx1_ASAP7_75t_L g1109 ( 
.A(n_975),
.Y(n_1109)
);

AND2x2_ASAP7_75t_L g1110 ( 
.A(n_825),
.B(n_592),
.Y(n_1110)
);

BUFx6f_ASAP7_75t_L g1111 ( 
.A(n_876),
.Y(n_1111)
);

NAND2xp5_ASAP7_75t_SL g1112 ( 
.A(n_934),
.B(n_702),
.Y(n_1112)
);

INVx3_ASAP7_75t_L g1113 ( 
.A(n_936),
.Y(n_1113)
);

NAND2xp5_ASAP7_75t_L g1114 ( 
.A(n_879),
.B(n_765),
.Y(n_1114)
);

NAND2xp5_ASAP7_75t_SL g1115 ( 
.A(n_937),
.B(n_702),
.Y(n_1115)
);

BUFx12f_ASAP7_75t_L g1116 ( 
.A(n_962),
.Y(n_1116)
);

AOI22xp5_ASAP7_75t_L g1117 ( 
.A1(n_937),
.A2(n_765),
.B1(n_770),
.B2(n_703),
.Y(n_1117)
);

INVx1_ASAP7_75t_L g1118 ( 
.A(n_976),
.Y(n_1118)
);

INVx1_ASAP7_75t_L g1119 ( 
.A(n_868),
.Y(n_1119)
);

INVx2_ASAP7_75t_SL g1120 ( 
.A(n_825),
.Y(n_1120)
);

NOR3xp33_ASAP7_75t_L g1121 ( 
.A(n_969),
.B(n_792),
.C(n_783),
.Y(n_1121)
);

INVx2_ASAP7_75t_SL g1122 ( 
.A(n_825),
.Y(n_1122)
);

INVx3_ASAP7_75t_L g1123 ( 
.A(n_936),
.Y(n_1123)
);

INVx2_ASAP7_75t_L g1124 ( 
.A(n_881),
.Y(n_1124)
);

BUFx12f_ASAP7_75t_SL g1125 ( 
.A(n_896),
.Y(n_1125)
);

INVx3_ASAP7_75t_SL g1126 ( 
.A(n_971),
.Y(n_1126)
);

HB1xp67_ASAP7_75t_L g1127 ( 
.A(n_971),
.Y(n_1127)
);

INVx2_ASAP7_75t_L g1128 ( 
.A(n_890),
.Y(n_1128)
);

INVx3_ASAP7_75t_L g1129 ( 
.A(n_961),
.Y(n_1129)
);

AND2x4_ASAP7_75t_L g1130 ( 
.A(n_871),
.B(n_734),
.Y(n_1130)
);

NAND2xp5_ASAP7_75t_L g1131 ( 
.A(n_835),
.B(n_770),
.Y(n_1131)
);

AND2x4_ASAP7_75t_L g1132 ( 
.A(n_871),
.B(n_734),
.Y(n_1132)
);

NAND2xp5_ASAP7_75t_L g1133 ( 
.A(n_911),
.B(n_707),
.Y(n_1133)
);

OAI21xp5_ASAP7_75t_L g1134 ( 
.A1(n_884),
.A2(n_708),
.B(n_707),
.Y(n_1134)
);

INVx4_ASAP7_75t_L g1135 ( 
.A(n_902),
.Y(n_1135)
);

HB1xp67_ASAP7_75t_L g1136 ( 
.A(n_971),
.Y(n_1136)
);

HB1xp67_ASAP7_75t_L g1137 ( 
.A(n_956),
.Y(n_1137)
);

NAND2xp5_ASAP7_75t_L g1138 ( 
.A(n_919),
.B(n_708),
.Y(n_1138)
);

NAND2xp5_ASAP7_75t_SL g1139 ( 
.A(n_957),
.B(n_702),
.Y(n_1139)
);

AND2x6_ASAP7_75t_L g1140 ( 
.A(n_855),
.B(n_717),
.Y(n_1140)
);

BUFx3_ASAP7_75t_L g1141 ( 
.A(n_920),
.Y(n_1141)
);

NAND2xp5_ASAP7_75t_L g1142 ( 
.A(n_884),
.B(n_717),
.Y(n_1142)
);

AND2x4_ASAP7_75t_L g1143 ( 
.A(n_833),
.B(n_734),
.Y(n_1143)
);

AOI22xp5_ASAP7_75t_L g1144 ( 
.A1(n_957),
.A2(n_926),
.B1(n_921),
.B2(n_838),
.Y(n_1144)
);

INVx2_ASAP7_75t_L g1145 ( 
.A(n_929),
.Y(n_1145)
);

AND3x1_ASAP7_75t_L g1146 ( 
.A(n_954),
.B(n_792),
.C(n_729),
.Y(n_1146)
);

HB1xp67_ASAP7_75t_L g1147 ( 
.A(n_938),
.Y(n_1147)
);

BUFx3_ASAP7_75t_L g1148 ( 
.A(n_921),
.Y(n_1148)
);

NAND2xp5_ASAP7_75t_L g1149 ( 
.A(n_939),
.B(n_946),
.Y(n_1149)
);

INVx1_ASAP7_75t_L g1150 ( 
.A(n_966),
.Y(n_1150)
);

AND2x4_ASAP7_75t_L g1151 ( 
.A(n_833),
.B(n_785),
.Y(n_1151)
);

AND2x2_ASAP7_75t_L g1152 ( 
.A(n_926),
.B(n_592),
.Y(n_1152)
);

NAND2xp5_ASAP7_75t_L g1153 ( 
.A(n_889),
.B(n_720),
.Y(n_1153)
);

INVx1_ASAP7_75t_L g1154 ( 
.A(n_927),
.Y(n_1154)
);

NOR2x2_ASAP7_75t_L g1155 ( 
.A(n_949),
.B(n_720),
.Y(n_1155)
);

NAND2xp5_ASAP7_75t_L g1156 ( 
.A(n_889),
.B(n_729),
.Y(n_1156)
);

INVx2_ASAP7_75t_L g1157 ( 
.A(n_928),
.Y(n_1157)
);

INVx1_ASAP7_75t_L g1158 ( 
.A(n_930),
.Y(n_1158)
);

NAND2xp5_ASAP7_75t_L g1159 ( 
.A(n_949),
.B(n_732),
.Y(n_1159)
);

NAND2xp5_ASAP7_75t_L g1160 ( 
.A(n_962),
.B(n_732),
.Y(n_1160)
);

NAND2xp5_ASAP7_75t_L g1161 ( 
.A(n_959),
.B(n_737),
.Y(n_1161)
);

INVx1_ASAP7_75t_L g1162 ( 
.A(n_943),
.Y(n_1162)
);

AOI21xp5_ASAP7_75t_L g1163 ( 
.A1(n_989),
.A2(n_970),
.B(n_849),
.Y(n_1163)
);

O2A1O1Ixp33_ASAP7_75t_L g1164 ( 
.A1(n_1137),
.A2(n_899),
.B(n_907),
.C(n_935),
.Y(n_1164)
);

BUFx12f_ASAP7_75t_L g1165 ( 
.A(n_998),
.Y(n_1165)
);

NAND2xp5_ASAP7_75t_L g1166 ( 
.A(n_982),
.B(n_935),
.Y(n_1166)
);

AOI22xp33_ASAP7_75t_L g1167 ( 
.A1(n_1090),
.A2(n_959),
.B1(n_897),
.B2(n_894),
.Y(n_1167)
);

AOI21xp5_ASAP7_75t_L g1168 ( 
.A1(n_989),
.A2(n_842),
.B(n_880),
.Y(n_1168)
);

OAI22x1_ASAP7_75t_L g1169 ( 
.A1(n_1144),
.A2(n_846),
.B1(n_882),
.B2(n_908),
.Y(n_1169)
);

INVx3_ASAP7_75t_L g1170 ( 
.A(n_984),
.Y(n_1170)
);

NAND2xp5_ASAP7_75t_L g1171 ( 
.A(n_1015),
.B(n_824),
.Y(n_1171)
);

AND2x2_ASAP7_75t_L g1172 ( 
.A(n_1076),
.B(n_963),
.Y(n_1172)
);

A2O1A1Ixp33_ASAP7_75t_SL g1173 ( 
.A1(n_1121),
.A2(n_824),
.B(n_961),
.C(n_792),
.Y(n_1173)
);

AOI222xp33_ASAP7_75t_L g1174 ( 
.A1(n_1078),
.A2(n_940),
.B1(n_895),
.B2(n_902),
.C1(n_426),
.C2(n_301),
.Y(n_1174)
);

NOR2xp33_ASAP7_75t_SL g1175 ( 
.A(n_990),
.B(n_785),
.Y(n_1175)
);

A2O1A1Ixp33_ASAP7_75t_L g1176 ( 
.A1(n_1079),
.A2(n_842),
.B(n_906),
.C(n_904),
.Y(n_1176)
);

NAND2xp5_ASAP7_75t_L g1177 ( 
.A(n_980),
.B(n_895),
.Y(n_1177)
);

NAND2xp5_ASAP7_75t_L g1178 ( 
.A(n_1027),
.B(n_940),
.Y(n_1178)
);

AND2x2_ASAP7_75t_L g1179 ( 
.A(n_1007),
.B(n_737),
.Y(n_1179)
);

AOI21xp5_ASAP7_75t_L g1180 ( 
.A1(n_993),
.A2(n_950),
.B(n_947),
.Y(n_1180)
);

AOI21xp5_ASAP7_75t_L g1181 ( 
.A1(n_993),
.A2(n_995),
.B(n_1079),
.Y(n_1181)
);

AOI21x1_ASAP7_75t_SL g1182 ( 
.A1(n_1095),
.A2(n_958),
.B(n_910),
.Y(n_1182)
);

NAND2xp5_ASAP7_75t_SL g1183 ( 
.A(n_1141),
.B(n_785),
.Y(n_1183)
);

NAND2xp5_ASAP7_75t_L g1184 ( 
.A(n_1030),
.B(n_739),
.Y(n_1184)
);

O2A1O1Ixp33_ASAP7_75t_L g1185 ( 
.A1(n_995),
.A2(n_869),
.B(n_847),
.C(n_739),
.Y(n_1185)
);

A2O1A1Ixp33_ASAP7_75t_L g1186 ( 
.A1(n_1148),
.A2(n_1061),
.B(n_1006),
.C(n_1048),
.Y(n_1186)
);

NOR2xp33_ASAP7_75t_L g1187 ( 
.A(n_1009),
.B(n_749),
.Y(n_1187)
);

INVx1_ASAP7_75t_L g1188 ( 
.A(n_978),
.Y(n_1188)
);

AOI21xp5_ASAP7_75t_L g1189 ( 
.A1(n_1095),
.A2(n_751),
.B(n_749),
.Y(n_1189)
);

AND2x4_ASAP7_75t_L g1190 ( 
.A(n_1057),
.B(n_744),
.Y(n_1190)
);

OAI21x1_ASAP7_75t_L g1191 ( 
.A1(n_987),
.A2(n_948),
.B(n_719),
.Y(n_1191)
);

NOR2xp33_ASAP7_75t_L g1192 ( 
.A(n_997),
.B(n_749),
.Y(n_1192)
);

NAND2xp5_ASAP7_75t_L g1193 ( 
.A(n_1082),
.B(n_744),
.Y(n_1193)
);

INVx1_ASAP7_75t_SL g1194 ( 
.A(n_1050),
.Y(n_1194)
);

BUFx6f_ASAP7_75t_SL g1195 ( 
.A(n_1005),
.Y(n_1195)
);

AOI21xp5_ASAP7_75t_L g1196 ( 
.A1(n_1091),
.A2(n_763),
.B(n_751),
.Y(n_1196)
);

INVx1_ASAP7_75t_SL g1197 ( 
.A(n_1033),
.Y(n_1197)
);

HB1xp67_ASAP7_75t_L g1198 ( 
.A(n_1127),
.Y(n_1198)
);

HB1xp67_ASAP7_75t_L g1199 ( 
.A(n_1136),
.Y(n_1199)
);

NAND2x1p5_ASAP7_75t_L g1200 ( 
.A(n_984),
.B(n_773),
.Y(n_1200)
);

INVx1_ASAP7_75t_L g1201 ( 
.A(n_981),
.Y(n_1201)
);

NOR2x1_ASAP7_75t_R g1202 ( 
.A(n_1008),
.B(n_250),
.Y(n_1202)
);

NAND2xp5_ASAP7_75t_L g1203 ( 
.A(n_1071),
.B(n_747),
.Y(n_1203)
);

INVx1_ASAP7_75t_SL g1204 ( 
.A(n_1045),
.Y(n_1204)
);

CKINVDCx5p33_ASAP7_75t_R g1205 ( 
.A(n_1029),
.Y(n_1205)
);

INVx2_ASAP7_75t_L g1206 ( 
.A(n_1097),
.Y(n_1206)
);

AOI22x1_ASAP7_75t_L g1207 ( 
.A1(n_1046),
.A2(n_761),
.B1(n_763),
.B2(n_751),
.Y(n_1207)
);

AOI21x1_ASAP7_75t_L g1208 ( 
.A1(n_1139),
.A2(n_761),
.B(n_772),
.Y(n_1208)
);

O2A1O1Ixp5_ASAP7_75t_SL g1209 ( 
.A1(n_1026),
.A2(n_658),
.B(n_719),
.C(n_721),
.Y(n_1209)
);

BUFx2_ASAP7_75t_L g1210 ( 
.A(n_998),
.Y(n_1210)
);

O2A1O1Ixp33_ASAP7_75t_L g1211 ( 
.A1(n_1119),
.A2(n_338),
.B(n_381),
.C(n_388),
.Y(n_1211)
);

AOI22xp33_ASAP7_75t_L g1212 ( 
.A1(n_1090),
.A2(n_948),
.B1(n_340),
.B2(n_403),
.Y(n_1212)
);

AOI21xp5_ASAP7_75t_L g1213 ( 
.A1(n_1091),
.A2(n_1099),
.B(n_1069),
.Y(n_1213)
);

O2A1O1Ixp5_ASAP7_75t_L g1214 ( 
.A1(n_1051),
.A2(n_751),
.B(n_763),
.C(n_719),
.Y(n_1214)
);

NOR2xp67_ASAP7_75t_L g1215 ( 
.A(n_1036),
.B(n_772),
.Y(n_1215)
);

INVx2_ASAP7_75t_L g1216 ( 
.A(n_1106),
.Y(n_1216)
);

BUFx3_ASAP7_75t_L g1217 ( 
.A(n_1032),
.Y(n_1217)
);

AOI21xp5_ASAP7_75t_L g1218 ( 
.A1(n_1099),
.A2(n_763),
.B(n_721),
.Y(n_1218)
);

NOR2xp33_ASAP7_75t_L g1219 ( 
.A(n_1022),
.B(n_658),
.Y(n_1219)
);

NAND2xp5_ASAP7_75t_SL g1220 ( 
.A(n_984),
.B(n_716),
.Y(n_1220)
);

OAI22xp33_ASAP7_75t_L g1221 ( 
.A1(n_994),
.A2(n_259),
.B1(n_335),
.B2(n_391),
.Y(n_1221)
);

BUFx3_ASAP7_75t_L g1222 ( 
.A(n_1100),
.Y(n_1222)
);

OAI22xp5_ASAP7_75t_L g1223 ( 
.A1(n_1131),
.A2(n_658),
.B1(n_721),
.B2(n_758),
.Y(n_1223)
);

NAND3xp33_ASAP7_75t_SL g1224 ( 
.A(n_994),
.B(n_253),
.C(n_252),
.Y(n_1224)
);

BUFx2_ASAP7_75t_L g1225 ( 
.A(n_1125),
.Y(n_1225)
);

OR2x6_ASAP7_75t_L g1226 ( 
.A(n_985),
.B(n_776),
.Y(n_1226)
);

NOR2xp33_ASAP7_75t_L g1227 ( 
.A(n_986),
.B(n_748),
.Y(n_1227)
);

BUFx6f_ASAP7_75t_L g1228 ( 
.A(n_985),
.Y(n_1228)
);

AOI21xp5_ASAP7_75t_L g1229 ( 
.A1(n_1065),
.A2(n_758),
.B(n_748),
.Y(n_1229)
);

AOI22xp33_ASAP7_75t_L g1230 ( 
.A1(n_1120),
.A2(n_393),
.B1(n_330),
.B2(n_421),
.Y(n_1230)
);

BUFx4f_ASAP7_75t_L g1231 ( 
.A(n_1111),
.Y(n_1231)
);

INVxp67_ASAP7_75t_L g1232 ( 
.A(n_1035),
.Y(n_1232)
);

INVx1_ASAP7_75t_L g1233 ( 
.A(n_991),
.Y(n_1233)
);

NAND2xp5_ASAP7_75t_L g1234 ( 
.A(n_1081),
.B(n_748),
.Y(n_1234)
);

NOR2xp33_ASAP7_75t_SL g1235 ( 
.A(n_1057),
.B(n_252),
.Y(n_1235)
);

OAI21xp5_ASAP7_75t_L g1236 ( 
.A1(n_1065),
.A2(n_758),
.B(n_776),
.Y(n_1236)
);

BUFx12f_ASAP7_75t_L g1237 ( 
.A(n_1019),
.Y(n_1237)
);

INVx1_ASAP7_75t_L g1238 ( 
.A(n_1001),
.Y(n_1238)
);

CKINVDCx6p67_ASAP7_75t_R g1239 ( 
.A(n_1031),
.Y(n_1239)
);

INVx1_ASAP7_75t_L g1240 ( 
.A(n_1017),
.Y(n_1240)
);

AOI21xp5_ASAP7_75t_L g1241 ( 
.A1(n_1069),
.A2(n_726),
.B(n_716),
.Y(n_1241)
);

AOI21xp5_ASAP7_75t_L g1242 ( 
.A1(n_1131),
.A2(n_726),
.B(n_716),
.Y(n_1242)
);

NAND2xp5_ASAP7_75t_SL g1243 ( 
.A(n_1010),
.B(n_716),
.Y(n_1243)
);

AOI21xp5_ASAP7_75t_L g1244 ( 
.A1(n_999),
.A2(n_1006),
.B(n_1084),
.Y(n_1244)
);

NAND3xp33_ASAP7_75t_L g1245 ( 
.A(n_1052),
.B(n_357),
.C(n_343),
.Y(n_1245)
);

NOR2xp33_ASAP7_75t_SL g1246 ( 
.A(n_1135),
.B(n_253),
.Y(n_1246)
);

AOI21xp5_ASAP7_75t_L g1247 ( 
.A1(n_999),
.A2(n_726),
.B(n_716),
.Y(n_1247)
);

NAND3xp33_ASAP7_75t_SL g1248 ( 
.A(n_1016),
.B(n_1004),
.C(n_1013),
.Y(n_1248)
);

BUFx12f_ASAP7_75t_L g1249 ( 
.A(n_1135),
.Y(n_1249)
);

NAND2xp5_ASAP7_75t_SL g1250 ( 
.A(n_1010),
.B(n_726),
.Y(n_1250)
);

NOR2xp33_ASAP7_75t_L g1251 ( 
.A(n_1147),
.B(n_996),
.Y(n_1251)
);

OAI22xp5_ASAP7_75t_L g1252 ( 
.A1(n_1000),
.A2(n_784),
.B1(n_795),
.B2(n_255),
.Y(n_1252)
);

AOI22xp33_ASAP7_75t_L g1253 ( 
.A1(n_1122),
.A2(n_406),
.B1(n_602),
.B2(n_328),
.Y(n_1253)
);

NAND2xp5_ASAP7_75t_L g1254 ( 
.A(n_1037),
.B(n_784),
.Y(n_1254)
);

OAI22xp5_ASAP7_75t_L g1255 ( 
.A1(n_1000),
.A2(n_795),
.B1(n_254),
.B2(n_259),
.Y(n_1255)
);

NOR2xp33_ASAP7_75t_L g1256 ( 
.A(n_1154),
.B(n_726),
.Y(n_1256)
);

NAND2xp5_ASAP7_75t_L g1257 ( 
.A(n_1020),
.B(n_745),
.Y(n_1257)
);

NAND2xp5_ASAP7_75t_L g1258 ( 
.A(n_1034),
.B(n_745),
.Y(n_1258)
);

O2A1O1Ixp33_ASAP7_75t_L g1259 ( 
.A1(n_1002),
.A2(n_585),
.B(n_578),
.C(n_575),
.Y(n_1259)
);

NAND2xp5_ASAP7_75t_SL g1260 ( 
.A(n_1010),
.B(n_745),
.Y(n_1260)
);

BUFx3_ASAP7_75t_L g1261 ( 
.A(n_985),
.Y(n_1261)
);

AOI21xp5_ASAP7_75t_L g1262 ( 
.A1(n_1084),
.A2(n_762),
.B(n_745),
.Y(n_1262)
);

OAI21xp33_ASAP7_75t_SL g1263 ( 
.A1(n_1038),
.A2(n_1),
.B(n_2),
.Y(n_1263)
);

NOR3xp33_ASAP7_75t_L g1264 ( 
.A(n_983),
.B(n_441),
.C(n_442),
.Y(n_1264)
);

OR2x2_ASAP7_75t_L g1265 ( 
.A(n_1101),
.B(n_745),
.Y(n_1265)
);

A2O1A1Ixp33_ASAP7_75t_L g1266 ( 
.A1(n_1086),
.A2(n_762),
.B(n_257),
.C(n_256),
.Y(n_1266)
);

NOR2xp33_ASAP7_75t_R g1267 ( 
.A(n_1111),
.B(n_254),
.Y(n_1267)
);

NAND2xp5_ASAP7_75t_SL g1268 ( 
.A(n_1010),
.B(n_762),
.Y(n_1268)
);

NAND2xp5_ASAP7_75t_L g1269 ( 
.A(n_1042),
.B(n_762),
.Y(n_1269)
);

OAI22xp5_ASAP7_75t_L g1270 ( 
.A1(n_1002),
.A2(n_255),
.B1(n_399),
.B2(n_256),
.Y(n_1270)
);

AOI21xp5_ASAP7_75t_L g1271 ( 
.A1(n_1086),
.A2(n_1138),
.B(n_1133),
.Y(n_1271)
);

AOI21xp5_ASAP7_75t_L g1272 ( 
.A1(n_1133),
.A2(n_762),
.B(n_364),
.Y(n_1272)
);

NAND2xp5_ASAP7_75t_L g1273 ( 
.A(n_1053),
.B(n_257),
.Y(n_1273)
);

AND2x4_ASAP7_75t_SL g1274 ( 
.A(n_1111),
.B(n_225),
.Y(n_1274)
);

OAI22xp5_ASAP7_75t_L g1275 ( 
.A1(n_1003),
.A2(n_335),
.B1(n_391),
.B2(n_394),
.Y(n_1275)
);

INVx2_ASAP7_75t_L g1276 ( 
.A(n_1124),
.Y(n_1276)
);

NOR3xp33_ASAP7_75t_L g1277 ( 
.A(n_1089),
.B(n_442),
.C(n_394),
.Y(n_1277)
);

INVx2_ASAP7_75t_L g1278 ( 
.A(n_1128),
.Y(n_1278)
);

AOI21xp5_ASAP7_75t_L g1279 ( 
.A1(n_1072),
.A2(n_360),
.B(n_289),
.Y(n_1279)
);

INVxp67_ASAP7_75t_SL g1280 ( 
.A(n_987),
.Y(n_1280)
);

AOI21xp5_ASAP7_75t_L g1281 ( 
.A1(n_1073),
.A2(n_385),
.B(n_291),
.Y(n_1281)
);

AND2x2_ASAP7_75t_L g1282 ( 
.A(n_979),
.B(n_5),
.Y(n_1282)
);

HB1xp67_ASAP7_75t_L g1283 ( 
.A(n_1160),
.Y(n_1283)
);

AOI22xp33_ASAP7_75t_L g1284 ( 
.A1(n_1126),
.A2(n_1059),
.B1(n_1058),
.B2(n_1110),
.Y(n_1284)
);

BUFx6f_ASAP7_75t_L g1285 ( 
.A(n_1018),
.Y(n_1285)
);

INVx1_ASAP7_75t_L g1286 ( 
.A(n_1066),
.Y(n_1286)
);

NOR2xp33_ASAP7_75t_SL g1287 ( 
.A(n_1116),
.B(n_396),
.Y(n_1287)
);

AOI22xp5_ASAP7_75t_L g1288 ( 
.A1(n_1146),
.A2(n_397),
.B1(n_396),
.B2(n_399),
.Y(n_1288)
);

INVx1_ASAP7_75t_L g1289 ( 
.A(n_1067),
.Y(n_1289)
);

OR2x6_ASAP7_75t_SL g1290 ( 
.A(n_1024),
.B(n_397),
.Y(n_1290)
);

NOR2xp33_ASAP7_75t_R g1291 ( 
.A(n_1018),
.B(n_441),
.Y(n_1291)
);

INVx2_ASAP7_75t_L g1292 ( 
.A(n_1145),
.Y(n_1292)
);

AND2x2_ASAP7_75t_L g1293 ( 
.A(n_1070),
.B(n_6),
.Y(n_1293)
);

O2A1O1Ixp5_ASAP7_75t_SL g1294 ( 
.A1(n_1115),
.A2(n_602),
.B(n_574),
.C(n_575),
.Y(n_1294)
);

NOR2xp33_ASAP7_75t_R g1295 ( 
.A(n_1018),
.B(n_262),
.Y(n_1295)
);

INVx2_ASAP7_75t_SL g1296 ( 
.A(n_1040),
.Y(n_1296)
);

INVx2_ASAP7_75t_SL g1297 ( 
.A(n_1098),
.Y(n_1297)
);

INVx6_ASAP7_75t_L g1298 ( 
.A(n_1018),
.Y(n_1298)
);

AOI21xp5_ASAP7_75t_L g1299 ( 
.A1(n_1075),
.A2(n_356),
.B(n_304),
.Y(n_1299)
);

INVx4_ASAP7_75t_L g1300 ( 
.A(n_1054),
.Y(n_1300)
);

OAI21xp5_ASAP7_75t_L g1301 ( 
.A1(n_1028),
.A2(n_585),
.B(n_578),
.Y(n_1301)
);

BUFx2_ASAP7_75t_L g1302 ( 
.A(n_1063),
.Y(n_1302)
);

HB1xp67_ASAP7_75t_L g1303 ( 
.A(n_1160),
.Y(n_1303)
);

NOR2xp33_ASAP7_75t_L g1304 ( 
.A(n_1063),
.B(n_1158),
.Y(n_1304)
);

AOI21xp5_ASAP7_75t_L g1305 ( 
.A1(n_1003),
.A2(n_358),
.B(n_313),
.Y(n_1305)
);

INVx1_ASAP7_75t_L g1306 ( 
.A(n_1150),
.Y(n_1306)
);

O2A1O1Ixp33_ASAP7_75t_L g1307 ( 
.A1(n_1102),
.A2(n_578),
.B(n_575),
.C(n_585),
.Y(n_1307)
);

NOR2xp33_ASAP7_75t_L g1308 ( 
.A(n_1162),
.B(n_1012),
.Y(n_1308)
);

BUFx12f_ASAP7_75t_L g1309 ( 
.A(n_992),
.Y(n_1309)
);

BUFx6f_ASAP7_75t_L g1310 ( 
.A(n_992),
.Y(n_1310)
);

BUFx3_ASAP7_75t_L g1311 ( 
.A(n_992),
.Y(n_1311)
);

NAND2xp5_ASAP7_75t_L g1312 ( 
.A(n_1157),
.B(n_7),
.Y(n_1312)
);

O2A1O1Ixp33_ASAP7_75t_L g1313 ( 
.A1(n_1104),
.A2(n_574),
.B(n_9),
.C(n_11),
.Y(n_1313)
);

BUFx12f_ASAP7_75t_L g1314 ( 
.A(n_1041),
.Y(n_1314)
);

INVx1_ASAP7_75t_SL g1315 ( 
.A(n_1068),
.Y(n_1315)
);

O2A1O1Ixp33_ASAP7_75t_SL g1316 ( 
.A1(n_1025),
.A2(n_574),
.B(n_9),
.C(n_13),
.Y(n_1316)
);

NAND2xp5_ASAP7_75t_L g1317 ( 
.A(n_1108),
.B(n_8),
.Y(n_1317)
);

NOR2xp33_ASAP7_75t_L g1318 ( 
.A(n_1083),
.B(n_8),
.Y(n_1318)
);

OAI21x1_ASAP7_75t_L g1319 ( 
.A1(n_1242),
.A2(n_988),
.B(n_1039),
.Y(n_1319)
);

NAND2xp5_ASAP7_75t_SL g1320 ( 
.A(n_1166),
.B(n_1054),
.Y(n_1320)
);

AO22x2_ASAP7_75t_L g1321 ( 
.A1(n_1248),
.A2(n_1105),
.B1(n_1114),
.B2(n_1155),
.Y(n_1321)
);

OAI21x1_ASAP7_75t_L g1322 ( 
.A1(n_1182),
.A2(n_988),
.B(n_1039),
.Y(n_1322)
);

AO31x2_ASAP7_75t_L g1323 ( 
.A1(n_1271),
.A2(n_1156),
.A3(n_1153),
.B(n_1105),
.Y(n_1323)
);

AND2x4_ASAP7_75t_L g1324 ( 
.A(n_1261),
.B(n_1054),
.Y(n_1324)
);

OAI21x1_ASAP7_75t_L g1325 ( 
.A1(n_1182),
.A2(n_1134),
.B(n_1142),
.Y(n_1325)
);

AO32x2_ASAP7_75t_L g1326 ( 
.A1(n_1223),
.A2(n_1114),
.A3(n_1064),
.B1(n_1159),
.B2(n_1153),
.Y(n_1326)
);

HB1xp67_ASAP7_75t_L g1327 ( 
.A(n_1197),
.Y(n_1327)
);

INVx1_ASAP7_75t_L g1328 ( 
.A(n_1188),
.Y(n_1328)
);

NOR2xp33_ASAP7_75t_SL g1329 ( 
.A(n_1224),
.B(n_1077),
.Y(n_1329)
);

AOI21xp5_ASAP7_75t_L g1330 ( 
.A1(n_1181),
.A2(n_1014),
.B(n_1011),
.Y(n_1330)
);

INVx1_ASAP7_75t_L g1331 ( 
.A(n_1201),
.Y(n_1331)
);

BUFx6f_ASAP7_75t_L g1332 ( 
.A(n_1228),
.Y(n_1332)
);

NAND2xp5_ASAP7_75t_L g1333 ( 
.A(n_1171),
.B(n_1109),
.Y(n_1333)
);

BUFx2_ASAP7_75t_L g1334 ( 
.A(n_1217),
.Y(n_1334)
);

NAND2xp5_ASAP7_75t_L g1335 ( 
.A(n_1283),
.B(n_1118),
.Y(n_1335)
);

AOI221xp5_ASAP7_75t_SL g1336 ( 
.A1(n_1221),
.A2(n_1094),
.B1(n_1088),
.B2(n_1085),
.C(n_1014),
.Y(n_1336)
);

NAND2xp5_ASAP7_75t_L g1337 ( 
.A(n_1283),
.B(n_1011),
.Y(n_1337)
);

AOI21xp5_ASAP7_75t_L g1338 ( 
.A1(n_1213),
.A2(n_1044),
.B(n_1043),
.Y(n_1338)
);

AOI21xp5_ASAP7_75t_L g1339 ( 
.A1(n_1244),
.A2(n_1044),
.B(n_1043),
.Y(n_1339)
);

AOI21xp5_ASAP7_75t_L g1340 ( 
.A1(n_1180),
.A2(n_1023),
.B(n_1142),
.Y(n_1340)
);

INVx1_ASAP7_75t_L g1341 ( 
.A(n_1233),
.Y(n_1341)
);

NAND2xp5_ASAP7_75t_L g1342 ( 
.A(n_1204),
.B(n_1152),
.Y(n_1342)
);

NOR2xp33_ASAP7_75t_L g1343 ( 
.A(n_1315),
.B(n_1046),
.Y(n_1343)
);

AOI21xp5_ASAP7_75t_L g1344 ( 
.A1(n_1247),
.A2(n_1023),
.B(n_1087),
.Y(n_1344)
);

INVx1_ASAP7_75t_L g1345 ( 
.A(n_1238),
.Y(n_1345)
);

AOI21xp5_ASAP7_75t_L g1346 ( 
.A1(n_1262),
.A2(n_1134),
.B(n_1112),
.Y(n_1346)
);

NAND3xp33_ASAP7_75t_L g1347 ( 
.A(n_1211),
.B(n_1060),
.C(n_1117),
.Y(n_1347)
);

AOI21xp5_ASAP7_75t_SL g1348 ( 
.A1(n_1186),
.A2(n_1151),
.B(n_1143),
.Y(n_1348)
);

OAI21xp5_ASAP7_75t_L g1349 ( 
.A1(n_1280),
.A2(n_1151),
.B(n_1140),
.Y(n_1349)
);

OAI21xp5_ASAP7_75t_L g1350 ( 
.A1(n_1280),
.A2(n_1140),
.B(n_1159),
.Y(n_1350)
);

NAND2xp5_ASAP7_75t_L g1351 ( 
.A(n_1304),
.B(n_1092),
.Y(n_1351)
);

OAI21xp5_ASAP7_75t_L g1352 ( 
.A1(n_1168),
.A2(n_1140),
.B(n_1080),
.Y(n_1352)
);

AOI21xp5_ASAP7_75t_L g1353 ( 
.A1(n_1241),
.A2(n_1021),
.B(n_1123),
.Y(n_1353)
);

OAI21x1_ASAP7_75t_L g1354 ( 
.A1(n_1191),
.A2(n_1156),
.B(n_1149),
.Y(n_1354)
);

OAI21xp5_ASAP7_75t_L g1355 ( 
.A1(n_1176),
.A2(n_1140),
.B(n_1080),
.Y(n_1355)
);

AOI221xp5_ASAP7_75t_L g1356 ( 
.A1(n_1221),
.A2(n_1132),
.B1(n_1130),
.B2(n_1143),
.C(n_1062),
.Y(n_1356)
);

AOI21xp5_ASAP7_75t_SL g1357 ( 
.A1(n_1211),
.A2(n_1161),
.B(n_1130),
.Y(n_1357)
);

OAI21x1_ASAP7_75t_L g1358 ( 
.A1(n_1208),
.A2(n_1149),
.B(n_1103),
.Y(n_1358)
);

INVxp67_ASAP7_75t_L g1359 ( 
.A(n_1251),
.Y(n_1359)
);

NAND2xp5_ASAP7_75t_SL g1360 ( 
.A(n_1174),
.B(n_1077),
.Y(n_1360)
);

AOI21xp5_ASAP7_75t_L g1361 ( 
.A1(n_1185),
.A2(n_1021),
.B(n_1113),
.Y(n_1361)
);

BUFx4_ASAP7_75t_SL g1362 ( 
.A(n_1205),
.Y(n_1362)
);

NAND2xp5_ASAP7_75t_L g1363 ( 
.A(n_1172),
.B(n_1049),
.Y(n_1363)
);

NAND3x1_ASAP7_75t_L g1364 ( 
.A(n_1264),
.B(n_1107),
.C(n_1129),
.Y(n_1364)
);

AOI221x1_ASAP7_75t_L g1365 ( 
.A1(n_1169),
.A2(n_1161),
.B1(n_1107),
.B2(n_1132),
.C(n_1129),
.Y(n_1365)
);

BUFx6f_ASAP7_75t_L g1366 ( 
.A(n_1228),
.Y(n_1366)
);

NOR3xp33_ASAP7_75t_SL g1367 ( 
.A(n_1263),
.B(n_322),
.C(n_318),
.Y(n_1367)
);

AO21x2_ASAP7_75t_L g1368 ( 
.A1(n_1259),
.A2(n_1096),
.B(n_1140),
.Y(n_1368)
);

OAI21x1_ASAP7_75t_L g1369 ( 
.A1(n_1294),
.A2(n_1113),
.B(n_1123),
.Y(n_1369)
);

NAND2xp5_ASAP7_75t_SL g1370 ( 
.A(n_1287),
.B(n_1192),
.Y(n_1370)
);

OAI21x1_ASAP7_75t_L g1371 ( 
.A1(n_1209),
.A2(n_1080),
.B(n_1077),
.Y(n_1371)
);

HB1xp67_ASAP7_75t_L g1372 ( 
.A(n_1232),
.Y(n_1372)
);

AOI221xp5_ASAP7_75t_L g1373 ( 
.A1(n_1224),
.A2(n_1096),
.B1(n_1093),
.B2(n_1041),
.C(n_1074),
.Y(n_1373)
);

INVx2_ASAP7_75t_SL g1374 ( 
.A(n_1231),
.Y(n_1374)
);

BUFx10_ASAP7_75t_L g1375 ( 
.A(n_1195),
.Y(n_1375)
);

BUFx2_ASAP7_75t_L g1376 ( 
.A(n_1225),
.Y(n_1376)
);

AOI21xp5_ASAP7_75t_L g1377 ( 
.A1(n_1185),
.A2(n_1077),
.B(n_1093),
.Y(n_1377)
);

AOI21xp5_ASAP7_75t_L g1378 ( 
.A1(n_1189),
.A2(n_1093),
.B(n_1074),
.Y(n_1378)
);

INVx1_ASAP7_75t_L g1379 ( 
.A(n_1240),
.Y(n_1379)
);

OA21x2_ASAP7_75t_L g1380 ( 
.A1(n_1214),
.A2(n_1080),
.B(n_383),
.Y(n_1380)
);

NAND2xp5_ASAP7_75t_L g1381 ( 
.A(n_1194),
.B(n_1055),
.Y(n_1381)
);

AO31x2_ASAP7_75t_L g1382 ( 
.A1(n_1163),
.A2(n_1080),
.A3(n_1074),
.B(n_1056),
.Y(n_1382)
);

NAND2xp5_ASAP7_75t_L g1383 ( 
.A(n_1302),
.B(n_1055),
.Y(n_1383)
);

A2O1A1Ixp33_ASAP7_75t_L g1384 ( 
.A1(n_1164),
.A2(n_1056),
.B(n_1055),
.C(n_267),
.Y(n_1384)
);

AOI21x1_ASAP7_75t_L g1385 ( 
.A1(n_1196),
.A2(n_1056),
.B(n_602),
.Y(n_1385)
);

OAI21x1_ASAP7_75t_L g1386 ( 
.A1(n_1214),
.A2(n_373),
.B(n_582),
.Y(n_1386)
);

AND2x2_ASAP7_75t_L g1387 ( 
.A(n_1282),
.B(n_14),
.Y(n_1387)
);

OA21x2_ASAP7_75t_L g1388 ( 
.A1(n_1236),
.A2(n_271),
.B(n_314),
.Y(n_1388)
);

OAI22x1_ASAP7_75t_L g1389 ( 
.A1(n_1227),
.A2(n_283),
.B1(n_296),
.B2(n_324),
.Y(n_1389)
);

NAND2xp5_ASAP7_75t_L g1390 ( 
.A(n_1179),
.B(n_14),
.Y(n_1390)
);

BUFx3_ASAP7_75t_L g1391 ( 
.A(n_1249),
.Y(n_1391)
);

NAND2xp5_ASAP7_75t_SL g1392 ( 
.A(n_1235),
.B(n_329),
.Y(n_1392)
);

INVxp67_ASAP7_75t_SL g1393 ( 
.A(n_1303),
.Y(n_1393)
);

OAI22xp5_ASAP7_75t_L g1394 ( 
.A1(n_1318),
.A2(n_16),
.B1(n_17),
.B2(n_20),
.Y(n_1394)
);

INVx3_ASAP7_75t_L g1395 ( 
.A(n_1285),
.Y(n_1395)
);

AND2x2_ASAP7_75t_L g1396 ( 
.A(n_1293),
.B(n_17),
.Y(n_1396)
);

AOI21xp5_ASAP7_75t_L g1397 ( 
.A1(n_1218),
.A2(n_249),
.B(n_370),
.Y(n_1397)
);

OAI21xp5_ASAP7_75t_L g1398 ( 
.A1(n_1229),
.A2(n_1307),
.B(n_1259),
.Y(n_1398)
);

OAI21x1_ASAP7_75t_L g1399 ( 
.A1(n_1207),
.A2(n_373),
.B(n_582),
.Y(n_1399)
);

OR2x2_ASAP7_75t_L g1400 ( 
.A(n_1222),
.B(n_22),
.Y(n_1400)
);

INVx2_ASAP7_75t_L g1401 ( 
.A(n_1206),
.Y(n_1401)
);

CKINVDCx20_ASAP7_75t_R g1402 ( 
.A(n_1239),
.Y(n_1402)
);

INVx5_ASAP7_75t_L g1403 ( 
.A(n_1226),
.Y(n_1403)
);

AO32x2_ASAP7_75t_L g1404 ( 
.A1(n_1252),
.A2(n_22),
.A3(n_25),
.B1(n_27),
.B2(n_28),
.Y(n_1404)
);

AOI21x1_ASAP7_75t_L g1405 ( 
.A1(n_1272),
.A2(n_582),
.B(n_373),
.Y(n_1405)
);

NAND2xp5_ASAP7_75t_L g1406 ( 
.A(n_1303),
.B(n_27),
.Y(n_1406)
);

A2O1A1Ixp33_ASAP7_75t_L g1407 ( 
.A1(n_1164),
.A2(n_405),
.B(n_331),
.C(n_434),
.Y(n_1407)
);

OAI22xp5_ASAP7_75t_L g1408 ( 
.A1(n_1318),
.A2(n_31),
.B1(n_32),
.B2(n_33),
.Y(n_1408)
);

OAI21x1_ASAP7_75t_SL g1409 ( 
.A1(n_1178),
.A2(n_32),
.B(n_34),
.Y(n_1409)
);

CKINVDCx16_ASAP7_75t_R g1410 ( 
.A(n_1165),
.Y(n_1410)
);

OAI21x1_ASAP7_75t_L g1411 ( 
.A1(n_1307),
.A2(n_373),
.B(n_582),
.Y(n_1411)
);

NAND2xp5_ASAP7_75t_L g1412 ( 
.A(n_1167),
.B(n_35),
.Y(n_1412)
);

NAND2xp5_ASAP7_75t_L g1413 ( 
.A(n_1198),
.B(n_1199),
.Y(n_1413)
);

OAI21x1_ASAP7_75t_L g1414 ( 
.A1(n_1301),
.A2(n_373),
.B(n_582),
.Y(n_1414)
);

NAND3xp33_ASAP7_75t_L g1415 ( 
.A(n_1313),
.B(n_249),
.C(n_370),
.Y(n_1415)
);

BUFx2_ASAP7_75t_L g1416 ( 
.A(n_1267),
.Y(n_1416)
);

AOI21xp5_ASAP7_75t_L g1417 ( 
.A1(n_1173),
.A2(n_249),
.B(n_370),
.Y(n_1417)
);

OAI21x1_ASAP7_75t_L g1418 ( 
.A1(n_1193),
.A2(n_373),
.B(n_582),
.Y(n_1418)
);

BUFx3_ASAP7_75t_L g1419 ( 
.A(n_1210),
.Y(n_1419)
);

AOI211x1_ASAP7_75t_L g1420 ( 
.A1(n_1177),
.A2(n_36),
.B(n_38),
.C(n_42),
.Y(n_1420)
);

OAI21xp5_ASAP7_75t_L g1421 ( 
.A1(n_1317),
.A2(n_416),
.B(n_334),
.Y(n_1421)
);

AOI21x1_ASAP7_75t_L g1422 ( 
.A1(n_1220),
.A2(n_582),
.B(n_373),
.Y(n_1422)
);

INVx3_ASAP7_75t_L g1423 ( 
.A(n_1285),
.Y(n_1423)
);

AOI221xp5_ASAP7_75t_L g1424 ( 
.A1(n_1313),
.A2(n_433),
.B1(n_333),
.B2(n_342),
.C(n_348),
.Y(n_1424)
);

NAND2xp5_ASAP7_75t_L g1425 ( 
.A(n_1167),
.B(n_46),
.Y(n_1425)
);

AOI21xp5_ASAP7_75t_L g1426 ( 
.A1(n_1257),
.A2(n_249),
.B(n_370),
.Y(n_1426)
);

AOI21xp5_ASAP7_75t_L g1427 ( 
.A1(n_1258),
.A2(n_1269),
.B(n_1256),
.Y(n_1427)
);

OAI21x1_ASAP7_75t_L g1428 ( 
.A1(n_1203),
.A2(n_373),
.B(n_178),
.Y(n_1428)
);

AOI21xp5_ASAP7_75t_L g1429 ( 
.A1(n_1256),
.A2(n_249),
.B(n_370),
.Y(n_1429)
);

AOI21xp5_ASAP7_75t_L g1430 ( 
.A1(n_1234),
.A2(n_1184),
.B(n_1268),
.Y(n_1430)
);

OAI21x1_ASAP7_75t_L g1431 ( 
.A1(n_1243),
.A2(n_132),
.B(n_128),
.Y(n_1431)
);

INVx3_ASAP7_75t_L g1432 ( 
.A(n_1285),
.Y(n_1432)
);

BUFx10_ASAP7_75t_L g1433 ( 
.A(n_1195),
.Y(n_1433)
);

INVx3_ASAP7_75t_L g1434 ( 
.A(n_1285),
.Y(n_1434)
);

AND2x2_ASAP7_75t_L g1435 ( 
.A(n_1199),
.B(n_49),
.Y(n_1435)
);

AOI21xp5_ASAP7_75t_L g1436 ( 
.A1(n_1250),
.A2(n_386),
.B(n_432),
.Y(n_1436)
);

OA21x2_ASAP7_75t_L g1437 ( 
.A1(n_1266),
.A2(n_419),
.B(n_430),
.Y(n_1437)
);

AOI21xp5_ASAP7_75t_L g1438 ( 
.A1(n_1260),
.A2(n_386),
.B(n_428),
.Y(n_1438)
);

BUFx4_ASAP7_75t_SL g1439 ( 
.A(n_1311),
.Y(n_1439)
);

BUFx6f_ASAP7_75t_L g1440 ( 
.A(n_1228),
.Y(n_1440)
);

AOI22xp5_ASAP7_75t_L g1441 ( 
.A1(n_1248),
.A2(n_427),
.B1(n_415),
.B2(n_355),
.Y(n_1441)
);

INVx4_ASAP7_75t_L g1442 ( 
.A(n_1228),
.Y(n_1442)
);

NAND2xp5_ASAP7_75t_L g1443 ( 
.A(n_1308),
.B(n_49),
.Y(n_1443)
);

NAND2xp5_ASAP7_75t_SL g1444 ( 
.A(n_1246),
.B(n_354),
.Y(n_1444)
);

NAND2xp5_ASAP7_75t_L g1445 ( 
.A(n_1286),
.B(n_50),
.Y(n_1445)
);

AO31x2_ASAP7_75t_L g1446 ( 
.A1(n_1306),
.A2(n_386),
.A3(n_808),
.B(n_102),
.Y(n_1446)
);

NAND2xp5_ASAP7_75t_L g1447 ( 
.A(n_1289),
.B(n_51),
.Y(n_1447)
);

AOI21xp5_ASAP7_75t_L g1448 ( 
.A1(n_1255),
.A2(n_386),
.B(n_808),
.Y(n_1448)
);

NOR2xp33_ASAP7_75t_L g1449 ( 
.A(n_1290),
.B(n_1237),
.Y(n_1449)
);

OAI21xp5_ASAP7_75t_L g1450 ( 
.A1(n_1312),
.A2(n_808),
.B(n_54),
.Y(n_1450)
);

BUFx6f_ASAP7_75t_L g1451 ( 
.A(n_1231),
.Y(n_1451)
);

AOI21xp5_ASAP7_75t_L g1452 ( 
.A1(n_1183),
.A2(n_808),
.B(n_115),
.Y(n_1452)
);

OAI21xp5_ASAP7_75t_L g1453 ( 
.A1(n_1245),
.A2(n_53),
.B(n_56),
.Y(n_1453)
);

O2A1O1Ixp33_ASAP7_75t_L g1454 ( 
.A1(n_1264),
.A2(n_57),
.B(n_59),
.C(n_61),
.Y(n_1454)
);

A2O1A1Ixp33_ASAP7_75t_L g1455 ( 
.A1(n_1212),
.A2(n_61),
.B(n_62),
.C(n_64),
.Y(n_1455)
);

HB1xp67_ASAP7_75t_L g1456 ( 
.A(n_1309),
.Y(n_1456)
);

OR2x6_ASAP7_75t_L g1457 ( 
.A(n_1226),
.B(n_1314),
.Y(n_1457)
);

OAI21xp5_ASAP7_75t_L g1458 ( 
.A1(n_1187),
.A2(n_62),
.B(n_64),
.Y(n_1458)
);

AO31x2_ASAP7_75t_L g1459 ( 
.A1(n_1216),
.A2(n_155),
.A3(n_214),
.B(n_205),
.Y(n_1459)
);

AOI21x1_ASAP7_75t_L g1460 ( 
.A1(n_1305),
.A2(n_133),
.B(n_199),
.Y(n_1460)
);

NAND2xp5_ASAP7_75t_L g1461 ( 
.A(n_1212),
.B(n_65),
.Y(n_1461)
);

OAI22xp5_ASAP7_75t_L g1462 ( 
.A1(n_1288),
.A2(n_1284),
.B1(n_1230),
.B2(n_1273),
.Y(n_1462)
);

OAI21xp5_ASAP7_75t_L g1463 ( 
.A1(n_1254),
.A2(n_66),
.B(n_67),
.Y(n_1463)
);

INVx2_ASAP7_75t_L g1464 ( 
.A(n_1276),
.Y(n_1464)
);

AO21x1_ASAP7_75t_L g1465 ( 
.A1(n_1277),
.A2(n_68),
.B(n_88),
.Y(n_1465)
);

NOR2xp67_ASAP7_75t_SL g1466 ( 
.A(n_1300),
.B(n_95),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_1278),
.Y(n_1467)
);

AO21x2_ASAP7_75t_L g1468 ( 
.A1(n_1277),
.A2(n_97),
.B(n_154),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_1292),
.Y(n_1469)
);

OAI21x1_ASAP7_75t_L g1470 ( 
.A1(n_1200),
.A2(n_160),
.B(n_167),
.Y(n_1470)
);

INVx2_ASAP7_75t_L g1471 ( 
.A(n_1265),
.Y(n_1471)
);

AOI21x1_ASAP7_75t_SL g1472 ( 
.A1(n_1190),
.A2(n_180),
.B(n_182),
.Y(n_1472)
);

NAND2xp5_ASAP7_75t_L g1473 ( 
.A(n_1219),
.B(n_219),
.Y(n_1473)
);

CKINVDCx5p33_ASAP7_75t_R g1474 ( 
.A(n_1291),
.Y(n_1474)
);

NOR2xp33_ASAP7_75t_R g1475 ( 
.A(n_1175),
.B(n_1298),
.Y(n_1475)
);

NAND2xp5_ASAP7_75t_L g1476 ( 
.A(n_1284),
.B(n_1270),
.Y(n_1476)
);

INVx4_ASAP7_75t_L g1477 ( 
.A(n_1298),
.Y(n_1477)
);

OR2x2_ASAP7_75t_L g1478 ( 
.A(n_1275),
.B(n_1296),
.Y(n_1478)
);

OAI21xp5_ASAP7_75t_L g1479 ( 
.A1(n_1279),
.A2(n_1281),
.B(n_1299),
.Y(n_1479)
);

INVx1_ASAP7_75t_L g1480 ( 
.A(n_1297),
.Y(n_1480)
);

NOR2xp33_ASAP7_75t_SL g1481 ( 
.A(n_1274),
.B(n_1300),
.Y(n_1481)
);

OAI21x1_ASAP7_75t_L g1482 ( 
.A1(n_1200),
.A2(n_1170),
.B(n_1230),
.Y(n_1482)
);

INVxp67_ASAP7_75t_L g1483 ( 
.A(n_1202),
.Y(n_1483)
);

AO32x2_ASAP7_75t_L g1484 ( 
.A1(n_1316),
.A2(n_1253),
.A3(n_1310),
.B1(n_1215),
.B2(n_1295),
.Y(n_1484)
);

NAND2xp5_ASAP7_75t_L g1485 ( 
.A(n_1190),
.B(n_1310),
.Y(n_1485)
);

OAI21x1_ASAP7_75t_L g1486 ( 
.A1(n_1170),
.A2(n_1253),
.B(n_1310),
.Y(n_1486)
);

OAI22xp5_ASAP7_75t_L g1487 ( 
.A1(n_1298),
.A2(n_1166),
.B1(n_1144),
.B2(n_1171),
.Y(n_1487)
);

OA21x2_ASAP7_75t_L g1488 ( 
.A1(n_1365),
.A2(n_1310),
.B(n_1319),
.Y(n_1488)
);

OAI21x1_ASAP7_75t_L g1489 ( 
.A1(n_1418),
.A2(n_1414),
.B(n_1344),
.Y(n_1489)
);

AO21x2_ASAP7_75t_L g1490 ( 
.A1(n_1398),
.A2(n_1350),
.B(n_1338),
.Y(n_1490)
);

AOI22xp33_ASAP7_75t_L g1491 ( 
.A1(n_1462),
.A2(n_1476),
.B1(n_1360),
.B2(n_1347),
.Y(n_1491)
);

OAI21x1_ASAP7_75t_L g1492 ( 
.A1(n_1322),
.A2(n_1346),
.B(n_1340),
.Y(n_1492)
);

INVx2_ASAP7_75t_L g1493 ( 
.A(n_1323),
.Y(n_1493)
);

AOI22xp33_ASAP7_75t_L g1494 ( 
.A1(n_1462),
.A2(n_1347),
.B1(n_1425),
.B2(n_1412),
.Y(n_1494)
);

INVx3_ASAP7_75t_L g1495 ( 
.A(n_1382),
.Y(n_1495)
);

AND2x2_ASAP7_75t_L g1496 ( 
.A(n_1349),
.B(n_1350),
.Y(n_1496)
);

INVx3_ASAP7_75t_L g1497 ( 
.A(n_1382),
.Y(n_1497)
);

OAI21x1_ASAP7_75t_L g1498 ( 
.A1(n_1411),
.A2(n_1339),
.B(n_1385),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_1328),
.Y(n_1499)
);

AO21x2_ASAP7_75t_L g1500 ( 
.A1(n_1398),
.A2(n_1415),
.B(n_1330),
.Y(n_1500)
);

INVx1_ASAP7_75t_L g1501 ( 
.A(n_1331),
.Y(n_1501)
);

OAI21x1_ASAP7_75t_L g1502 ( 
.A1(n_1405),
.A2(n_1325),
.B(n_1352),
.Y(n_1502)
);

OAI21x1_ASAP7_75t_L g1503 ( 
.A1(n_1352),
.A2(n_1397),
.B(n_1354),
.Y(n_1503)
);

OAI21x1_ASAP7_75t_L g1504 ( 
.A1(n_1358),
.A2(n_1428),
.B(n_1386),
.Y(n_1504)
);

OAI21xp5_ASAP7_75t_L g1505 ( 
.A1(n_1415),
.A2(n_1487),
.B(n_1425),
.Y(n_1505)
);

OAI21x1_ASAP7_75t_L g1506 ( 
.A1(n_1355),
.A2(n_1472),
.B(n_1378),
.Y(n_1506)
);

CKINVDCx8_ASAP7_75t_R g1507 ( 
.A(n_1410),
.Y(n_1507)
);

AND2x4_ASAP7_75t_L g1508 ( 
.A(n_1403),
.B(n_1457),
.Y(n_1508)
);

OAI21x1_ASAP7_75t_L g1509 ( 
.A1(n_1355),
.A2(n_1422),
.B(n_1353),
.Y(n_1509)
);

BUFx8_ASAP7_75t_L g1510 ( 
.A(n_1416),
.Y(n_1510)
);

INVx1_ASAP7_75t_L g1511 ( 
.A(n_1341),
.Y(n_1511)
);

OAI21x1_ASAP7_75t_L g1512 ( 
.A1(n_1371),
.A2(n_1399),
.B(n_1361),
.Y(n_1512)
);

OAI21x1_ASAP7_75t_L g1513 ( 
.A1(n_1369),
.A2(n_1377),
.B(n_1426),
.Y(n_1513)
);

BUFx4f_ASAP7_75t_L g1514 ( 
.A(n_1451),
.Y(n_1514)
);

NAND2xp5_ASAP7_75t_L g1515 ( 
.A(n_1359),
.B(n_1333),
.Y(n_1515)
);

NAND2xp5_ASAP7_75t_L g1516 ( 
.A(n_1333),
.B(n_1327),
.Y(n_1516)
);

HB1xp67_ASAP7_75t_L g1517 ( 
.A(n_1372),
.Y(n_1517)
);

OAI21xp5_ASAP7_75t_L g1518 ( 
.A1(n_1487),
.A2(n_1412),
.B(n_1450),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_1345),
.Y(n_1519)
);

OAI21x1_ASAP7_75t_L g1520 ( 
.A1(n_1427),
.A2(n_1417),
.B(n_1429),
.Y(n_1520)
);

OAI21x1_ASAP7_75t_L g1521 ( 
.A1(n_1430),
.A2(n_1349),
.B(n_1460),
.Y(n_1521)
);

OAI21x1_ASAP7_75t_L g1522 ( 
.A1(n_1482),
.A2(n_1486),
.B(n_1431),
.Y(n_1522)
);

BUFx2_ASAP7_75t_L g1523 ( 
.A(n_1334),
.Y(n_1523)
);

NAND2x1p5_ASAP7_75t_L g1524 ( 
.A(n_1403),
.B(n_1477),
.Y(n_1524)
);

AO21x2_ASAP7_75t_L g1525 ( 
.A1(n_1368),
.A2(n_1450),
.B(n_1357),
.Y(n_1525)
);

OR2x2_ASAP7_75t_L g1526 ( 
.A(n_1413),
.B(n_1393),
.Y(n_1526)
);

INVx2_ASAP7_75t_L g1527 ( 
.A(n_1323),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_1379),
.Y(n_1528)
);

AOI22xp33_ASAP7_75t_L g1529 ( 
.A1(n_1321),
.A2(n_1461),
.B1(n_1471),
.B2(n_1394),
.Y(n_1529)
);

OAI22xp5_ASAP7_75t_L g1530 ( 
.A1(n_1443),
.A2(n_1478),
.B1(n_1421),
.B2(n_1458),
.Y(n_1530)
);

OAI21x1_ASAP7_75t_L g1531 ( 
.A1(n_1380),
.A2(n_1470),
.B(n_1479),
.Y(n_1531)
);

BUFx2_ASAP7_75t_R g1532 ( 
.A(n_1474),
.Y(n_1532)
);

AOI21xp5_ASAP7_75t_L g1533 ( 
.A1(n_1348),
.A2(n_1329),
.B(n_1320),
.Y(n_1533)
);

OAI21x1_ASAP7_75t_L g1534 ( 
.A1(n_1380),
.A2(n_1479),
.B(n_1448),
.Y(n_1534)
);

INVx1_ASAP7_75t_L g1535 ( 
.A(n_1467),
.Y(n_1535)
);

OAI21x1_ASAP7_75t_SL g1536 ( 
.A1(n_1458),
.A2(n_1463),
.B(n_1409),
.Y(n_1536)
);

CKINVDCx5p33_ASAP7_75t_R g1537 ( 
.A(n_1362),
.Y(n_1537)
);

OA21x2_ASAP7_75t_L g1538 ( 
.A1(n_1336),
.A2(n_1463),
.B(n_1337),
.Y(n_1538)
);

OA21x2_ASAP7_75t_L g1539 ( 
.A1(n_1336),
.A2(n_1337),
.B(n_1384),
.Y(n_1539)
);

OAI21x1_ASAP7_75t_L g1540 ( 
.A1(n_1452),
.A2(n_1335),
.B(n_1364),
.Y(n_1540)
);

BUFx12f_ASAP7_75t_L g1541 ( 
.A(n_1375),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_1469),
.Y(n_1542)
);

NOR2xp33_ASAP7_75t_L g1543 ( 
.A(n_1370),
.B(n_1342),
.Y(n_1543)
);

OAI21x1_ASAP7_75t_L g1544 ( 
.A1(n_1335),
.A2(n_1388),
.B(n_1473),
.Y(n_1544)
);

OAI21x1_ASAP7_75t_L g1545 ( 
.A1(n_1388),
.A2(n_1434),
.B(n_1395),
.Y(n_1545)
);

OAI21x1_ASAP7_75t_L g1546 ( 
.A1(n_1395),
.A2(n_1434),
.B(n_1423),
.Y(n_1546)
);

AO22x2_ASAP7_75t_L g1547 ( 
.A1(n_1420),
.A2(n_1394),
.B1(n_1408),
.B2(n_1351),
.Y(n_1547)
);

CKINVDCx16_ASAP7_75t_R g1548 ( 
.A(n_1402),
.Y(n_1548)
);

OAI21x1_ASAP7_75t_L g1549 ( 
.A1(n_1423),
.A2(n_1432),
.B(n_1438),
.Y(n_1549)
);

OA21x2_ASAP7_75t_L g1550 ( 
.A1(n_1465),
.A2(n_1407),
.B(n_1453),
.Y(n_1550)
);

AOI22xp5_ASAP7_75t_L g1551 ( 
.A1(n_1329),
.A2(n_1408),
.B1(n_1441),
.B2(n_1343),
.Y(n_1551)
);

BUFx2_ASAP7_75t_L g1552 ( 
.A(n_1457),
.Y(n_1552)
);

OAI21x1_ASAP7_75t_L g1553 ( 
.A1(n_1432),
.A2(n_1436),
.B(n_1437),
.Y(n_1553)
);

OAI21x1_ASAP7_75t_L g1554 ( 
.A1(n_1437),
.A2(n_1485),
.B(n_1406),
.Y(n_1554)
);

OAI21x1_ASAP7_75t_L g1555 ( 
.A1(n_1363),
.A2(n_1447),
.B(n_1445),
.Y(n_1555)
);

BUFx2_ASAP7_75t_L g1556 ( 
.A(n_1457),
.Y(n_1556)
);

INVx2_ASAP7_75t_L g1557 ( 
.A(n_1401),
.Y(n_1557)
);

CKINVDCx20_ASAP7_75t_R g1558 ( 
.A(n_1391),
.Y(n_1558)
);

OAI21x1_ASAP7_75t_L g1559 ( 
.A1(n_1373),
.A2(n_1356),
.B(n_1390),
.Y(n_1559)
);

BUFx2_ASAP7_75t_L g1560 ( 
.A(n_1419),
.Y(n_1560)
);

INVx3_ASAP7_75t_L g1561 ( 
.A(n_1368),
.Y(n_1561)
);

OAI21x1_ASAP7_75t_L g1562 ( 
.A1(n_1383),
.A2(n_1464),
.B(n_1454),
.Y(n_1562)
);

OA21x2_ASAP7_75t_L g1563 ( 
.A1(n_1455),
.A2(n_1421),
.B(n_1424),
.Y(n_1563)
);

INVx1_ASAP7_75t_L g1564 ( 
.A(n_1435),
.Y(n_1564)
);

OAI21x1_ASAP7_75t_L g1565 ( 
.A1(n_1446),
.A2(n_1381),
.B(n_1480),
.Y(n_1565)
);

AOI21x1_ASAP7_75t_L g1566 ( 
.A1(n_1466),
.A2(n_1392),
.B(n_1444),
.Y(n_1566)
);

NAND2xp5_ASAP7_75t_L g1567 ( 
.A(n_1396),
.B(n_1376),
.Y(n_1567)
);

NAND2xp5_ASAP7_75t_L g1568 ( 
.A(n_1387),
.B(n_1451),
.Y(n_1568)
);

NAND3xp33_ASAP7_75t_L g1569 ( 
.A(n_1367),
.B(n_1400),
.C(n_1449),
.Y(n_1569)
);

OAI21x1_ASAP7_75t_L g1570 ( 
.A1(n_1446),
.A2(n_1484),
.B(n_1459),
.Y(n_1570)
);

OA21x2_ASAP7_75t_L g1571 ( 
.A1(n_1446),
.A2(n_1326),
.B(n_1321),
.Y(n_1571)
);

OR2x2_ASAP7_75t_L g1572 ( 
.A(n_1456),
.B(n_1440),
.Y(n_1572)
);

OAI21x1_ASAP7_75t_L g1573 ( 
.A1(n_1484),
.A2(n_1459),
.B(n_1326),
.Y(n_1573)
);

OAI21x1_ASAP7_75t_SL g1574 ( 
.A1(n_1442),
.A2(n_1477),
.B(n_1374),
.Y(n_1574)
);

NOR2x1_ASAP7_75t_R g1575 ( 
.A(n_1451),
.B(n_1442),
.Y(n_1575)
);

AND2x2_ASAP7_75t_L g1576 ( 
.A(n_1326),
.B(n_1404),
.Y(n_1576)
);

NAND2xp5_ASAP7_75t_L g1577 ( 
.A(n_1324),
.B(n_1332),
.Y(n_1577)
);

OAI21x1_ASAP7_75t_L g1578 ( 
.A1(n_1484),
.A2(n_1459),
.B(n_1468),
.Y(n_1578)
);

INVx1_ASAP7_75t_SL g1579 ( 
.A(n_1439),
.Y(n_1579)
);

AOI21xp5_ASAP7_75t_L g1580 ( 
.A1(n_1481),
.A2(n_1468),
.B(n_1403),
.Y(n_1580)
);

OAI21x1_ASAP7_75t_L g1581 ( 
.A1(n_1481),
.A2(n_1404),
.B(n_1475),
.Y(n_1581)
);

OAI21x1_ASAP7_75t_L g1582 ( 
.A1(n_1404),
.A2(n_1332),
.B(n_1366),
.Y(n_1582)
);

AOI22xp33_ASAP7_75t_SL g1583 ( 
.A1(n_1324),
.A2(n_1375),
.B1(n_1433),
.B2(n_1332),
.Y(n_1583)
);

AOI22xp33_ASAP7_75t_L g1584 ( 
.A1(n_1389),
.A2(n_1433),
.B1(n_1483),
.B2(n_1440),
.Y(n_1584)
);

INVx2_ASAP7_75t_SL g1585 ( 
.A(n_1366),
.Y(n_1585)
);

INVx1_ASAP7_75t_L g1586 ( 
.A(n_1366),
.Y(n_1586)
);

AND2x2_ASAP7_75t_L g1587 ( 
.A(n_1440),
.B(n_1349),
.Y(n_1587)
);

OAI22xp5_ASAP7_75t_L g1588 ( 
.A1(n_1476),
.A2(n_1166),
.B1(n_1144),
.B2(n_1137),
.Y(n_1588)
);

INVx2_ASAP7_75t_SL g1589 ( 
.A(n_1403),
.Y(n_1589)
);

INVx2_ASAP7_75t_L g1590 ( 
.A(n_1323),
.Y(n_1590)
);

OAI21x1_ASAP7_75t_L g1591 ( 
.A1(n_1418),
.A2(n_1414),
.B(n_1319),
.Y(n_1591)
);

OAI21x1_ASAP7_75t_L g1592 ( 
.A1(n_1418),
.A2(n_1414),
.B(n_1319),
.Y(n_1592)
);

INVx3_ASAP7_75t_L g1593 ( 
.A(n_1382),
.Y(n_1593)
);

OAI21x1_ASAP7_75t_L g1594 ( 
.A1(n_1418),
.A2(n_1414),
.B(n_1319),
.Y(n_1594)
);

OA21x2_ASAP7_75t_L g1595 ( 
.A1(n_1365),
.A2(n_1319),
.B(n_1398),
.Y(n_1595)
);

INVx2_ASAP7_75t_L g1596 ( 
.A(n_1323),
.Y(n_1596)
);

BUFx3_ASAP7_75t_L g1597 ( 
.A(n_1451),
.Y(n_1597)
);

OAI21x1_ASAP7_75t_L g1598 ( 
.A1(n_1418),
.A2(n_1414),
.B(n_1319),
.Y(n_1598)
);

NOR2xp33_ASAP7_75t_L g1599 ( 
.A(n_1487),
.B(n_1166),
.Y(n_1599)
);

AOI21xp5_ASAP7_75t_L g1600 ( 
.A1(n_1339),
.A2(n_1181),
.B(n_1338),
.Y(n_1600)
);

OAI21x1_ASAP7_75t_L g1601 ( 
.A1(n_1418),
.A2(n_1414),
.B(n_1319),
.Y(n_1601)
);

HB1xp67_ASAP7_75t_L g1602 ( 
.A(n_1372),
.Y(n_1602)
);

AOI22xp33_ASAP7_75t_L g1603 ( 
.A1(n_1462),
.A2(n_945),
.B1(n_1047),
.B2(n_900),
.Y(n_1603)
);

O2A1O1Ixp33_ASAP7_75t_SL g1604 ( 
.A1(n_1458),
.A2(n_1166),
.B(n_1171),
.C(n_1407),
.Y(n_1604)
);

NAND2xp5_ASAP7_75t_L g1605 ( 
.A(n_1359),
.B(n_1333),
.Y(n_1605)
);

A2O1A1Ixp33_ASAP7_75t_L g1606 ( 
.A1(n_1458),
.A2(n_1144),
.B(n_1166),
.C(n_1211),
.Y(n_1606)
);

OAI21xp5_ASAP7_75t_L g1607 ( 
.A1(n_1415),
.A2(n_1144),
.B(n_1166),
.Y(n_1607)
);

OAI21x1_ASAP7_75t_L g1608 ( 
.A1(n_1418),
.A2(n_1414),
.B(n_1319),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_1328),
.Y(n_1609)
);

AO31x2_ASAP7_75t_L g1610 ( 
.A1(n_1365),
.A2(n_1338),
.A3(n_1330),
.B(n_1340),
.Y(n_1610)
);

AOI21xp5_ASAP7_75t_L g1611 ( 
.A1(n_1339),
.A2(n_1181),
.B(n_1338),
.Y(n_1611)
);

INVx1_ASAP7_75t_L g1612 ( 
.A(n_1328),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1328),
.Y(n_1613)
);

NAND2xp5_ASAP7_75t_L g1614 ( 
.A(n_1359),
.B(n_1333),
.Y(n_1614)
);

OAI22xp5_ASAP7_75t_L g1615 ( 
.A1(n_1476),
.A2(n_1166),
.B1(n_1144),
.B2(n_1137),
.Y(n_1615)
);

OAI22xp33_ASAP7_75t_L g1616 ( 
.A1(n_1476),
.A2(n_1144),
.B1(n_1166),
.B2(n_674),
.Y(n_1616)
);

AO21x2_ASAP7_75t_L g1617 ( 
.A1(n_1398),
.A2(n_1350),
.B(n_1338),
.Y(n_1617)
);

NAND3xp33_ASAP7_75t_L g1618 ( 
.A(n_1394),
.B(n_1144),
.C(n_1408),
.Y(n_1618)
);

BUFx6f_ASAP7_75t_L g1619 ( 
.A(n_1403),
.Y(n_1619)
);

BUFx2_ASAP7_75t_SL g1620 ( 
.A(n_1402),
.Y(n_1620)
);

OA21x2_ASAP7_75t_L g1621 ( 
.A1(n_1365),
.A2(n_1319),
.B(n_1398),
.Y(n_1621)
);

OAI21x1_ASAP7_75t_L g1622 ( 
.A1(n_1418),
.A2(n_1414),
.B(n_1319),
.Y(n_1622)
);

OAI22xp33_ASAP7_75t_L g1623 ( 
.A1(n_1476),
.A2(n_1144),
.B1(n_1166),
.B2(n_674),
.Y(n_1623)
);

OAI21x1_ASAP7_75t_L g1624 ( 
.A1(n_1418),
.A2(n_1414),
.B(n_1319),
.Y(n_1624)
);

AO21x2_ASAP7_75t_L g1625 ( 
.A1(n_1398),
.A2(n_1338),
.B(n_1415),
.Y(n_1625)
);

NOR2xp33_ASAP7_75t_L g1626 ( 
.A(n_1487),
.B(n_1166),
.Y(n_1626)
);

AND2x2_ASAP7_75t_L g1627 ( 
.A(n_1349),
.B(n_1350),
.Y(n_1627)
);

HB1xp67_ASAP7_75t_L g1628 ( 
.A(n_1372),
.Y(n_1628)
);

CKINVDCx5p33_ASAP7_75t_R g1629 ( 
.A(n_1362),
.Y(n_1629)
);

BUFx2_ASAP7_75t_L g1630 ( 
.A(n_1327),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_1328),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_1328),
.Y(n_1632)
);

INVx2_ASAP7_75t_L g1633 ( 
.A(n_1323),
.Y(n_1633)
);

AND2x4_ASAP7_75t_L g1634 ( 
.A(n_1403),
.B(n_1457),
.Y(n_1634)
);

INVx3_ASAP7_75t_L g1635 ( 
.A(n_1382),
.Y(n_1635)
);

INVx2_ASAP7_75t_L g1636 ( 
.A(n_1323),
.Y(n_1636)
);

BUFx3_ASAP7_75t_L g1637 ( 
.A(n_1451),
.Y(n_1637)
);

INVx1_ASAP7_75t_SL g1638 ( 
.A(n_1334),
.Y(n_1638)
);

NAND2xp5_ASAP7_75t_L g1639 ( 
.A(n_1359),
.B(n_1333),
.Y(n_1639)
);

INVx2_ASAP7_75t_L g1640 ( 
.A(n_1323),
.Y(n_1640)
);

INVx2_ASAP7_75t_L g1641 ( 
.A(n_1323),
.Y(n_1641)
);

OAI21x1_ASAP7_75t_L g1642 ( 
.A1(n_1418),
.A2(n_1414),
.B(n_1319),
.Y(n_1642)
);

AO32x2_ASAP7_75t_L g1643 ( 
.A1(n_1394),
.A2(n_1122),
.A3(n_1120),
.B1(n_1408),
.B2(n_1487),
.Y(n_1643)
);

INVx1_ASAP7_75t_SL g1644 ( 
.A(n_1334),
.Y(n_1644)
);

BUFx2_ASAP7_75t_SL g1645 ( 
.A(n_1402),
.Y(n_1645)
);

OAI21x1_ASAP7_75t_L g1646 ( 
.A1(n_1418),
.A2(n_1414),
.B(n_1319),
.Y(n_1646)
);

AND2x2_ASAP7_75t_L g1647 ( 
.A(n_1349),
.B(n_1350),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_1328),
.Y(n_1648)
);

OAI21x1_ASAP7_75t_L g1649 ( 
.A1(n_1418),
.A2(n_1414),
.B(n_1319),
.Y(n_1649)
);

INVx2_ASAP7_75t_L g1650 ( 
.A(n_1323),
.Y(n_1650)
);

OAI211xp5_ASAP7_75t_L g1651 ( 
.A1(n_1458),
.A2(n_1166),
.B(n_1144),
.C(n_1454),
.Y(n_1651)
);

OAI21x1_ASAP7_75t_L g1652 ( 
.A1(n_1418),
.A2(n_1414),
.B(n_1319),
.Y(n_1652)
);

INVx3_ASAP7_75t_L g1653 ( 
.A(n_1382),
.Y(n_1653)
);

INVx2_ASAP7_75t_L g1654 ( 
.A(n_1323),
.Y(n_1654)
);

OAI22xp5_ASAP7_75t_L g1655 ( 
.A1(n_1476),
.A2(n_1166),
.B1(n_1144),
.B2(n_1137),
.Y(n_1655)
);

AO21x1_ASAP7_75t_L g1656 ( 
.A1(n_1412),
.A2(n_1425),
.B(n_1211),
.Y(n_1656)
);

NAND2xp5_ASAP7_75t_L g1657 ( 
.A(n_1359),
.B(n_1333),
.Y(n_1657)
);

AOI22xp33_ASAP7_75t_SL g1658 ( 
.A1(n_1462),
.A2(n_916),
.B1(n_825),
.B2(n_909),
.Y(n_1658)
);

NOR3xp33_ASAP7_75t_L g1659 ( 
.A(n_1394),
.B(n_1408),
.C(n_1454),
.Y(n_1659)
);

OAI21xp5_ASAP7_75t_L g1660 ( 
.A1(n_1415),
.A2(n_1144),
.B(n_1166),
.Y(n_1660)
);

OAI21x1_ASAP7_75t_L g1661 ( 
.A1(n_1418),
.A2(n_1414),
.B(n_1319),
.Y(n_1661)
);

OR2x6_ASAP7_75t_L g1662 ( 
.A(n_1348),
.B(n_1349),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_1328),
.Y(n_1663)
);

INVx2_ASAP7_75t_L g1664 ( 
.A(n_1323),
.Y(n_1664)
);

O2A1O1Ixp33_ASAP7_75t_L g1665 ( 
.A1(n_1394),
.A2(n_1166),
.B(n_1408),
.C(n_1137),
.Y(n_1665)
);

OAI21x1_ASAP7_75t_L g1666 ( 
.A1(n_1418),
.A2(n_1414),
.B(n_1319),
.Y(n_1666)
);

CKINVDCx16_ASAP7_75t_R g1667 ( 
.A(n_1410),
.Y(n_1667)
);

A2O1A1Ixp33_ASAP7_75t_L g1668 ( 
.A1(n_1458),
.A2(n_1144),
.B(n_1166),
.C(n_1211),
.Y(n_1668)
);

BUFx2_ASAP7_75t_SL g1669 ( 
.A(n_1402),
.Y(n_1669)
);

AND2x4_ASAP7_75t_L g1670 ( 
.A(n_1403),
.B(n_1457),
.Y(n_1670)
);

INVx2_ASAP7_75t_L g1671 ( 
.A(n_1323),
.Y(n_1671)
);

AOI21xp5_ASAP7_75t_L g1672 ( 
.A1(n_1599),
.A2(n_1626),
.B(n_1606),
.Y(n_1672)
);

OR2x2_ASAP7_75t_L g1673 ( 
.A(n_1526),
.B(n_1516),
.Y(n_1673)
);

INVx1_ASAP7_75t_L g1674 ( 
.A(n_1499),
.Y(n_1674)
);

INVx1_ASAP7_75t_L g1675 ( 
.A(n_1501),
.Y(n_1675)
);

BUFx3_ASAP7_75t_L g1676 ( 
.A(n_1510),
.Y(n_1676)
);

CKINVDCx6p67_ASAP7_75t_R g1677 ( 
.A(n_1667),
.Y(n_1677)
);

OAI22xp5_ASAP7_75t_L g1678 ( 
.A1(n_1618),
.A2(n_1599),
.B1(n_1626),
.B2(n_1606),
.Y(n_1678)
);

AOI221xp5_ASAP7_75t_L g1679 ( 
.A1(n_1616),
.A2(n_1623),
.B1(n_1615),
.B2(n_1588),
.C(n_1655),
.Y(n_1679)
);

O2A1O1Ixp33_ASAP7_75t_L g1680 ( 
.A1(n_1668),
.A2(n_1530),
.B(n_1665),
.C(n_1659),
.Y(n_1680)
);

AOI21xp5_ASAP7_75t_L g1681 ( 
.A1(n_1668),
.A2(n_1611),
.B(n_1600),
.Y(n_1681)
);

O2A1O1Ixp5_ASAP7_75t_L g1682 ( 
.A1(n_1651),
.A2(n_1656),
.B(n_1518),
.C(n_1505),
.Y(n_1682)
);

AND2x2_ASAP7_75t_L g1683 ( 
.A(n_1564),
.B(n_1630),
.Y(n_1683)
);

INVx3_ASAP7_75t_L g1684 ( 
.A(n_1508),
.Y(n_1684)
);

OR2x2_ASAP7_75t_L g1685 ( 
.A(n_1517),
.B(n_1602),
.Y(n_1685)
);

AND2x2_ASAP7_75t_L g1686 ( 
.A(n_1628),
.B(n_1543),
.Y(n_1686)
);

BUFx2_ASAP7_75t_L g1687 ( 
.A(n_1523),
.Y(n_1687)
);

BUFx2_ASAP7_75t_L g1688 ( 
.A(n_1560),
.Y(n_1688)
);

NAND2xp5_ASAP7_75t_L g1689 ( 
.A(n_1515),
.B(n_1605),
.Y(n_1689)
);

O2A1O1Ixp33_ASAP7_75t_L g1690 ( 
.A1(n_1604),
.A2(n_1607),
.B(n_1660),
.C(n_1536),
.Y(n_1690)
);

AND2x2_ASAP7_75t_L g1691 ( 
.A(n_1543),
.B(n_1567),
.Y(n_1691)
);

AND2x2_ASAP7_75t_L g1692 ( 
.A(n_1614),
.B(n_1639),
.Y(n_1692)
);

NAND2xp5_ASAP7_75t_L g1693 ( 
.A(n_1657),
.B(n_1576),
.Y(n_1693)
);

OAI22xp5_ASAP7_75t_L g1694 ( 
.A1(n_1494),
.A2(n_1491),
.B1(n_1551),
.B2(n_1603),
.Y(n_1694)
);

AOI21xp5_ASAP7_75t_L g1695 ( 
.A1(n_1500),
.A2(n_1625),
.B(n_1617),
.Y(n_1695)
);

AND2x2_ASAP7_75t_L g1696 ( 
.A(n_1568),
.B(n_1638),
.Y(n_1696)
);

OAI22xp5_ASAP7_75t_L g1697 ( 
.A1(n_1658),
.A2(n_1547),
.B1(n_1662),
.B2(n_1563),
.Y(n_1697)
);

AND2x2_ASAP7_75t_L g1698 ( 
.A(n_1644),
.B(n_1511),
.Y(n_1698)
);

AOI211xp5_ASAP7_75t_L g1699 ( 
.A1(n_1604),
.A2(n_1569),
.B(n_1576),
.C(n_1555),
.Y(n_1699)
);

NAND2xp5_ASAP7_75t_L g1700 ( 
.A(n_1519),
.B(n_1528),
.Y(n_1700)
);

OAI22xp5_ASAP7_75t_L g1701 ( 
.A1(n_1547),
.A2(n_1662),
.B1(n_1563),
.B2(n_1529),
.Y(n_1701)
);

BUFx4f_ASAP7_75t_SL g1702 ( 
.A(n_1558),
.Y(n_1702)
);

AOI21x1_ASAP7_75t_SL g1703 ( 
.A1(n_1577),
.A2(n_1670),
.B(n_1634),
.Y(n_1703)
);

AND2x4_ASAP7_75t_SL g1704 ( 
.A(n_1558),
.B(n_1634),
.Y(n_1704)
);

INVx1_ASAP7_75t_SL g1705 ( 
.A(n_1552),
.Y(n_1705)
);

CKINVDCx5p33_ASAP7_75t_R g1706 ( 
.A(n_1537),
.Y(n_1706)
);

NAND2xp5_ASAP7_75t_L g1707 ( 
.A(n_1609),
.B(n_1612),
.Y(n_1707)
);

AND2x2_ASAP7_75t_L g1708 ( 
.A(n_1613),
.B(n_1631),
.Y(n_1708)
);

CKINVDCx5p33_ASAP7_75t_R g1709 ( 
.A(n_1537),
.Y(n_1709)
);

OA21x2_ASAP7_75t_L g1710 ( 
.A1(n_1578),
.A2(n_1570),
.B(n_1573),
.Y(n_1710)
);

OAI22xp5_ASAP7_75t_L g1711 ( 
.A1(n_1547),
.A2(n_1662),
.B1(n_1550),
.B2(n_1627),
.Y(n_1711)
);

BUFx3_ASAP7_75t_L g1712 ( 
.A(n_1510),
.Y(n_1712)
);

AOI21xp5_ASAP7_75t_L g1713 ( 
.A1(n_1500),
.A2(n_1625),
.B(n_1490),
.Y(n_1713)
);

NAND2xp5_ASAP7_75t_L g1714 ( 
.A(n_1632),
.B(n_1648),
.Y(n_1714)
);

AND2x2_ASAP7_75t_L g1715 ( 
.A(n_1663),
.B(n_1643),
.Y(n_1715)
);

AND2x4_ASAP7_75t_L g1716 ( 
.A(n_1670),
.B(n_1556),
.Y(n_1716)
);

AND2x4_ASAP7_75t_L g1717 ( 
.A(n_1662),
.B(n_1589),
.Y(n_1717)
);

OAI22xp5_ASAP7_75t_SL g1718 ( 
.A1(n_1507),
.A2(n_1548),
.B1(n_1579),
.B2(n_1645),
.Y(n_1718)
);

INVxp67_ASAP7_75t_L g1719 ( 
.A(n_1572),
.Y(n_1719)
);

OA21x2_ASAP7_75t_L g1720 ( 
.A1(n_1578),
.A2(n_1570),
.B(n_1573),
.Y(n_1720)
);

AND2x2_ASAP7_75t_L g1721 ( 
.A(n_1643),
.B(n_1496),
.Y(n_1721)
);

AND2x2_ASAP7_75t_L g1722 ( 
.A(n_1643),
.B(n_1496),
.Y(n_1722)
);

CKINVDCx16_ASAP7_75t_R g1723 ( 
.A(n_1620),
.Y(n_1723)
);

AOI21xp5_ASAP7_75t_SL g1724 ( 
.A1(n_1580),
.A2(n_1550),
.B(n_1533),
.Y(n_1724)
);

OAI22x1_ASAP7_75t_L g1725 ( 
.A1(n_1535),
.A2(n_1542),
.B1(n_1538),
.B2(n_1571),
.Y(n_1725)
);

OAI22xp5_ASAP7_75t_L g1726 ( 
.A1(n_1627),
.A2(n_1647),
.B1(n_1538),
.B2(n_1507),
.Y(n_1726)
);

NAND2xp5_ASAP7_75t_L g1727 ( 
.A(n_1538),
.B(n_1647),
.Y(n_1727)
);

NAND2xp5_ASAP7_75t_L g1728 ( 
.A(n_1539),
.B(n_1490),
.Y(n_1728)
);

OA21x2_ASAP7_75t_L g1729 ( 
.A1(n_1531),
.A2(n_1534),
.B(n_1492),
.Y(n_1729)
);

O2A1O1Ixp33_ASAP7_75t_L g1730 ( 
.A1(n_1539),
.A2(n_1574),
.B(n_1500),
.C(n_1586),
.Y(n_1730)
);

NAND2xp5_ASAP7_75t_L g1731 ( 
.A(n_1539),
.B(n_1490),
.Y(n_1731)
);

AND2x2_ASAP7_75t_L g1732 ( 
.A(n_1643),
.B(n_1581),
.Y(n_1732)
);

AND2x2_ASAP7_75t_SL g1733 ( 
.A(n_1619),
.B(n_1571),
.Y(n_1733)
);

BUFx3_ASAP7_75t_L g1734 ( 
.A(n_1510),
.Y(n_1734)
);

NAND2xp5_ASAP7_75t_L g1735 ( 
.A(n_1617),
.B(n_1555),
.Y(n_1735)
);

OA21x2_ASAP7_75t_L g1736 ( 
.A1(n_1531),
.A2(n_1534),
.B(n_1492),
.Y(n_1736)
);

O2A1O1Ixp33_ASAP7_75t_L g1737 ( 
.A1(n_1584),
.A2(n_1525),
.B(n_1617),
.C(n_1585),
.Y(n_1737)
);

NAND2xp5_ASAP7_75t_L g1738 ( 
.A(n_1565),
.B(n_1525),
.Y(n_1738)
);

AND2x2_ASAP7_75t_L g1739 ( 
.A(n_1581),
.B(n_1585),
.Y(n_1739)
);

O2A1O1Ixp5_ASAP7_75t_L g1740 ( 
.A1(n_1566),
.A2(n_1561),
.B(n_1514),
.C(n_1593),
.Y(n_1740)
);

AND2x2_ASAP7_75t_L g1741 ( 
.A(n_1554),
.B(n_1546),
.Y(n_1741)
);

AOI21xp5_ASAP7_75t_SL g1742 ( 
.A1(n_1575),
.A2(n_1525),
.B(n_1524),
.Y(n_1742)
);

NAND2x1p5_ASAP7_75t_L g1743 ( 
.A(n_1619),
.B(n_1540),
.Y(n_1743)
);

INVxp67_ASAP7_75t_L g1744 ( 
.A(n_1669),
.Y(n_1744)
);

AOI21xp5_ASAP7_75t_SL g1745 ( 
.A1(n_1524),
.A2(n_1637),
.B(n_1597),
.Y(n_1745)
);

O2A1O1Ixp33_ASAP7_75t_L g1746 ( 
.A1(n_1595),
.A2(n_1621),
.B(n_1637),
.C(n_1597),
.Y(n_1746)
);

NAND2xp5_ASAP7_75t_L g1747 ( 
.A(n_1565),
.B(n_1544),
.Y(n_1747)
);

AND2x2_ASAP7_75t_L g1748 ( 
.A(n_1546),
.B(n_1582),
.Y(n_1748)
);

INVx2_ASAP7_75t_SL g1749 ( 
.A(n_1541),
.Y(n_1749)
);

AND2x2_ASAP7_75t_L g1750 ( 
.A(n_1582),
.B(n_1562),
.Y(n_1750)
);

INVx5_ASAP7_75t_L g1751 ( 
.A(n_1619),
.Y(n_1751)
);

NAND2xp5_ASAP7_75t_L g1752 ( 
.A(n_1544),
.B(n_1493),
.Y(n_1752)
);

OAI22xp5_ASAP7_75t_L g1753 ( 
.A1(n_1595),
.A2(n_1621),
.B1(n_1583),
.B2(n_1571),
.Y(n_1753)
);

OR2x2_ASAP7_75t_L g1754 ( 
.A(n_1557),
.B(n_1595),
.Y(n_1754)
);

OAI22xp5_ASAP7_75t_L g1755 ( 
.A1(n_1514),
.A2(n_1488),
.B1(n_1532),
.B2(n_1629),
.Y(n_1755)
);

INVx1_ASAP7_75t_L g1756 ( 
.A(n_1671),
.Y(n_1756)
);

INVx1_ASAP7_75t_L g1757 ( 
.A(n_1671),
.Y(n_1757)
);

AOI21xp5_ASAP7_75t_SL g1758 ( 
.A1(n_1488),
.A2(n_1633),
.B(n_1493),
.Y(n_1758)
);

AND2x4_ASAP7_75t_L g1759 ( 
.A(n_1495),
.B(n_1593),
.Y(n_1759)
);

BUFx3_ASAP7_75t_L g1760 ( 
.A(n_1629),
.Y(n_1760)
);

AOI221xp5_ASAP7_75t_L g1761 ( 
.A1(n_1561),
.A2(n_1527),
.B1(n_1664),
.B2(n_1636),
.C(n_1640),
.Y(n_1761)
);

O2A1O1Ixp33_ASAP7_75t_L g1762 ( 
.A1(n_1561),
.A2(n_1488),
.B(n_1664),
.C(n_1650),
.Y(n_1762)
);

O2A1O1Ixp5_ASAP7_75t_L g1763 ( 
.A1(n_1514),
.A2(n_1635),
.B(n_1495),
.C(n_1497),
.Y(n_1763)
);

OAI22xp5_ASAP7_75t_SL g1764 ( 
.A1(n_1559),
.A2(n_1633),
.B1(n_1590),
.B2(n_1527),
.Y(n_1764)
);

O2A1O1Ixp33_ASAP7_75t_L g1765 ( 
.A1(n_1590),
.A2(n_1654),
.B(n_1650),
.C(n_1641),
.Y(n_1765)
);

OA21x2_ASAP7_75t_L g1766 ( 
.A1(n_1521),
.A2(n_1520),
.B(n_1513),
.Y(n_1766)
);

NAND2xp5_ASAP7_75t_L g1767 ( 
.A(n_1596),
.B(n_1636),
.Y(n_1767)
);

AND2x4_ASAP7_75t_L g1768 ( 
.A(n_1495),
.B(n_1653),
.Y(n_1768)
);

AND2x2_ASAP7_75t_L g1769 ( 
.A(n_1559),
.B(n_1545),
.Y(n_1769)
);

AOI221x1_ASAP7_75t_SL g1770 ( 
.A1(n_1610),
.A2(n_1506),
.B1(n_1502),
.B2(n_1553),
.C(n_1503),
.Y(n_1770)
);

AND2x2_ASAP7_75t_L g1771 ( 
.A(n_1549),
.B(n_1653),
.Y(n_1771)
);

NAND2xp5_ASAP7_75t_L g1772 ( 
.A(n_1497),
.B(n_1653),
.Y(n_1772)
);

CKINVDCx20_ASAP7_75t_R g1773 ( 
.A(n_1635),
.Y(n_1773)
);

INVx3_ASAP7_75t_L g1774 ( 
.A(n_1549),
.Y(n_1774)
);

BUFx12f_ASAP7_75t_L g1775 ( 
.A(n_1522),
.Y(n_1775)
);

NAND2xp5_ASAP7_75t_L g1776 ( 
.A(n_1503),
.B(n_1522),
.Y(n_1776)
);

OAI22xp5_ASAP7_75t_L g1777 ( 
.A1(n_1509),
.A2(n_1502),
.B1(n_1498),
.B2(n_1512),
.Y(n_1777)
);

HB1xp67_ASAP7_75t_L g1778 ( 
.A(n_1509),
.Y(n_1778)
);

A2O1A1Ixp33_ASAP7_75t_L g1779 ( 
.A1(n_1498),
.A2(n_1504),
.B(n_1512),
.C(n_1622),
.Y(n_1779)
);

AND2x2_ASAP7_75t_L g1780 ( 
.A(n_1504),
.B(n_1624),
.Y(n_1780)
);

AND2x2_ASAP7_75t_L g1781 ( 
.A(n_1591),
.B(n_1624),
.Y(n_1781)
);

OR2x2_ASAP7_75t_L g1782 ( 
.A(n_1592),
.B(n_1642),
.Y(n_1782)
);

HB1xp67_ASAP7_75t_L g1783 ( 
.A(n_1592),
.Y(n_1783)
);

A2O1A1Ixp33_ASAP7_75t_L g1784 ( 
.A1(n_1594),
.A2(n_1646),
.B(n_1598),
.C(n_1601),
.Y(n_1784)
);

O2A1O1Ixp33_ASAP7_75t_L g1785 ( 
.A1(n_1594),
.A2(n_1646),
.B(n_1598),
.C(n_1601),
.Y(n_1785)
);

NAND2xp5_ASAP7_75t_L g1786 ( 
.A(n_1608),
.B(n_1622),
.Y(n_1786)
);

BUFx3_ASAP7_75t_L g1787 ( 
.A(n_1649),
.Y(n_1787)
);

INVx1_ASAP7_75t_L g1788 ( 
.A(n_1652),
.Y(n_1788)
);

NOR2xp67_ASAP7_75t_L g1789 ( 
.A(n_1652),
.B(n_1661),
.Y(n_1789)
);

OAI22xp5_ASAP7_75t_L g1790 ( 
.A1(n_1661),
.A2(n_1618),
.B1(n_1626),
.B2(n_1599),
.Y(n_1790)
);

INVx1_ASAP7_75t_L g1791 ( 
.A(n_1666),
.Y(n_1791)
);

AOI21xp5_ASAP7_75t_L g1792 ( 
.A1(n_1489),
.A2(n_1626),
.B(n_1599),
.Y(n_1792)
);

NOR2xp67_ASAP7_75t_L g1793 ( 
.A(n_1666),
.B(n_1489),
.Y(n_1793)
);

OAI22xp5_ASAP7_75t_L g1794 ( 
.A1(n_1618),
.A2(n_1626),
.B1(n_1599),
.B2(n_1606),
.Y(n_1794)
);

NAND2xp5_ASAP7_75t_L g1795 ( 
.A(n_1599),
.B(n_1626),
.Y(n_1795)
);

AND2x2_ASAP7_75t_L g1796 ( 
.A(n_1564),
.B(n_1630),
.Y(n_1796)
);

AND2x2_ASAP7_75t_L g1797 ( 
.A(n_1564),
.B(n_1630),
.Y(n_1797)
);

AOI21x1_ASAP7_75t_SL g1798 ( 
.A1(n_1567),
.A2(n_1166),
.B(n_1443),
.Y(n_1798)
);

AOI21xp5_ASAP7_75t_L g1799 ( 
.A1(n_1600),
.A2(n_1611),
.B(n_1599),
.Y(n_1799)
);

AOI21xp5_ASAP7_75t_SL g1800 ( 
.A1(n_1606),
.A2(n_1668),
.B(n_1530),
.Y(n_1800)
);

AOI21xp5_ASAP7_75t_L g1801 ( 
.A1(n_1599),
.A2(n_1626),
.B(n_1606),
.Y(n_1801)
);

OA21x2_ASAP7_75t_L g1802 ( 
.A1(n_1578),
.A2(n_1570),
.B(n_1573),
.Y(n_1802)
);

OR2x2_ASAP7_75t_L g1803 ( 
.A(n_1526),
.B(n_1516),
.Y(n_1803)
);

AND2x2_ASAP7_75t_L g1804 ( 
.A(n_1564),
.B(n_1630),
.Y(n_1804)
);

O2A1O1Ixp5_ASAP7_75t_L g1805 ( 
.A1(n_1651),
.A2(n_1656),
.B(n_1668),
.C(n_1606),
.Y(n_1805)
);

HB1xp67_ASAP7_75t_L g1806 ( 
.A(n_1517),
.Y(n_1806)
);

AOI21xp5_ASAP7_75t_L g1807 ( 
.A1(n_1599),
.A2(n_1626),
.B(n_1606),
.Y(n_1807)
);

AOI21xp5_ASAP7_75t_SL g1808 ( 
.A1(n_1606),
.A2(n_1668),
.B(n_1530),
.Y(n_1808)
);

AOI21xp5_ASAP7_75t_SL g1809 ( 
.A1(n_1606),
.A2(n_1668),
.B(n_1530),
.Y(n_1809)
);

OAI22xp5_ASAP7_75t_L g1810 ( 
.A1(n_1618),
.A2(n_1626),
.B1(n_1599),
.B2(n_1606),
.Y(n_1810)
);

NOR2xp67_ASAP7_75t_L g1811 ( 
.A(n_1569),
.B(n_1359),
.Y(n_1811)
);

O2A1O1Ixp5_ASAP7_75t_L g1812 ( 
.A1(n_1651),
.A2(n_1656),
.B(n_1668),
.C(n_1606),
.Y(n_1812)
);

AOI21x1_ASAP7_75t_SL g1813 ( 
.A1(n_1567),
.A2(n_1166),
.B(n_1443),
.Y(n_1813)
);

CKINVDCx5p33_ASAP7_75t_R g1814 ( 
.A(n_1537),
.Y(n_1814)
);

AND2x4_ASAP7_75t_L g1815 ( 
.A(n_1587),
.B(n_1508),
.Y(n_1815)
);

BUFx2_ASAP7_75t_L g1816 ( 
.A(n_1775),
.Y(n_1816)
);

INVx1_ASAP7_75t_L g1817 ( 
.A(n_1700),
.Y(n_1817)
);

INVx4_ASAP7_75t_L g1818 ( 
.A(n_1751),
.Y(n_1818)
);

OAI21xp5_ASAP7_75t_L g1819 ( 
.A1(n_1672),
.A2(n_1807),
.B(n_1801),
.Y(n_1819)
);

OR2x2_ASAP7_75t_L g1820 ( 
.A(n_1721),
.B(n_1722),
.Y(n_1820)
);

INVx1_ASAP7_75t_L g1821 ( 
.A(n_1700),
.Y(n_1821)
);

AO21x2_ASAP7_75t_L g1822 ( 
.A1(n_1695),
.A2(n_1713),
.B(n_1728),
.Y(n_1822)
);

AND2x2_ASAP7_75t_L g1823 ( 
.A(n_1715),
.B(n_1732),
.Y(n_1823)
);

AO21x2_ASAP7_75t_L g1824 ( 
.A1(n_1695),
.A2(n_1731),
.B(n_1728),
.Y(n_1824)
);

OAI21xp5_ASAP7_75t_L g1825 ( 
.A1(n_1678),
.A2(n_1810),
.B(n_1794),
.Y(n_1825)
);

INVx1_ASAP7_75t_L g1826 ( 
.A(n_1707),
.Y(n_1826)
);

NAND2xp5_ASAP7_75t_L g1827 ( 
.A(n_1795),
.B(n_1692),
.Y(n_1827)
);

OR2x6_ASAP7_75t_L g1828 ( 
.A(n_1724),
.B(n_1742),
.Y(n_1828)
);

NAND3xp33_ASAP7_75t_SL g1829 ( 
.A(n_1679),
.B(n_1680),
.C(n_1805),
.Y(n_1829)
);

INVx1_ASAP7_75t_L g1830 ( 
.A(n_1707),
.Y(n_1830)
);

AND2x2_ASAP7_75t_L g1831 ( 
.A(n_1693),
.B(n_1727),
.Y(n_1831)
);

INVxp67_ASAP7_75t_L g1832 ( 
.A(n_1806),
.Y(n_1832)
);

BUFx3_ASAP7_75t_L g1833 ( 
.A(n_1704),
.Y(n_1833)
);

OR2x6_ASAP7_75t_L g1834 ( 
.A(n_1800),
.B(n_1808),
.Y(n_1834)
);

HB1xp67_ASAP7_75t_L g1835 ( 
.A(n_1685),
.Y(n_1835)
);

AO21x2_ASAP7_75t_L g1836 ( 
.A1(n_1747),
.A2(n_1738),
.B(n_1681),
.Y(n_1836)
);

INVx1_ASAP7_75t_L g1837 ( 
.A(n_1714),
.Y(n_1837)
);

AOI22xp33_ASAP7_75t_L g1838 ( 
.A1(n_1694),
.A2(n_1697),
.B1(n_1679),
.B2(n_1810),
.Y(n_1838)
);

OR2x2_ASAP7_75t_L g1839 ( 
.A(n_1693),
.B(n_1673),
.Y(n_1839)
);

AND2x2_ASAP7_75t_L g1840 ( 
.A(n_1727),
.B(n_1711),
.Y(n_1840)
);

AOI21xp5_ASAP7_75t_L g1841 ( 
.A1(n_1799),
.A2(n_1809),
.B(n_1794),
.Y(n_1841)
);

INVx1_ASAP7_75t_L g1842 ( 
.A(n_1714),
.Y(n_1842)
);

HB1xp67_ASAP7_75t_L g1843 ( 
.A(n_1686),
.Y(n_1843)
);

INVx1_ASAP7_75t_SL g1844 ( 
.A(n_1702),
.Y(n_1844)
);

INVx3_ASAP7_75t_L g1845 ( 
.A(n_1748),
.Y(n_1845)
);

INVx1_ASAP7_75t_L g1846 ( 
.A(n_1674),
.Y(n_1846)
);

INVx2_ASAP7_75t_L g1847 ( 
.A(n_1754),
.Y(n_1847)
);

AND2x2_ASAP7_75t_L g1848 ( 
.A(n_1711),
.B(n_1795),
.Y(n_1848)
);

OR2x6_ASAP7_75t_L g1849 ( 
.A(n_1737),
.B(n_1717),
.Y(n_1849)
);

AOI21x1_ASAP7_75t_L g1850 ( 
.A1(n_1789),
.A2(n_1793),
.B(n_1735),
.Y(n_1850)
);

INVx1_ASAP7_75t_L g1851 ( 
.A(n_1675),
.Y(n_1851)
);

INVx2_ASAP7_75t_SL g1852 ( 
.A(n_1687),
.Y(n_1852)
);

OR2x2_ASAP7_75t_L g1853 ( 
.A(n_1803),
.B(n_1726),
.Y(n_1853)
);

INVxp67_ASAP7_75t_L g1854 ( 
.A(n_1688),
.Y(n_1854)
);

INVxp67_ASAP7_75t_SL g1855 ( 
.A(n_1735),
.Y(n_1855)
);

HB1xp67_ASAP7_75t_L g1856 ( 
.A(n_1698),
.Y(n_1856)
);

HB1xp67_ASAP7_75t_L g1857 ( 
.A(n_1683),
.Y(n_1857)
);

AND2x4_ASAP7_75t_L g1858 ( 
.A(n_1759),
.B(n_1768),
.Y(n_1858)
);

OAI21xp5_ASAP7_75t_L g1859 ( 
.A1(n_1678),
.A2(n_1812),
.B(n_1682),
.Y(n_1859)
);

INVx1_ASAP7_75t_L g1860 ( 
.A(n_1725),
.Y(n_1860)
);

AOI22xp5_ASAP7_75t_L g1861 ( 
.A1(n_1694),
.A2(n_1697),
.B1(n_1701),
.B2(n_1811),
.Y(n_1861)
);

OR2x6_ASAP7_75t_L g1862 ( 
.A(n_1758),
.B(n_1746),
.Y(n_1862)
);

AO21x2_ASAP7_75t_L g1863 ( 
.A1(n_1738),
.A2(n_1752),
.B(n_1784),
.Y(n_1863)
);

AND2x2_ASAP7_75t_L g1864 ( 
.A(n_1726),
.B(n_1708),
.Y(n_1864)
);

HB1xp67_ASAP7_75t_L g1865 ( 
.A(n_1796),
.Y(n_1865)
);

CKINVDCx11_ASAP7_75t_R g1866 ( 
.A(n_1677),
.Y(n_1866)
);

AO21x2_ASAP7_75t_L g1867 ( 
.A1(n_1752),
.A2(n_1753),
.B(n_1779),
.Y(n_1867)
);

OAI21x1_ASAP7_75t_L g1868 ( 
.A1(n_1785),
.A2(n_1777),
.B(n_1799),
.Y(n_1868)
);

INVx1_ASAP7_75t_L g1869 ( 
.A(n_1739),
.Y(n_1869)
);

BUFx4_ASAP7_75t_R g1870 ( 
.A(n_1676),
.Y(n_1870)
);

AND2x2_ASAP7_75t_L g1871 ( 
.A(n_1691),
.B(n_1769),
.Y(n_1871)
);

INVx1_ASAP7_75t_L g1872 ( 
.A(n_1767),
.Y(n_1872)
);

INVx1_ASAP7_75t_L g1873 ( 
.A(n_1767),
.Y(n_1873)
);

INVx1_ASAP7_75t_L g1874 ( 
.A(n_1756),
.Y(n_1874)
);

OR2x6_ASAP7_75t_L g1875 ( 
.A(n_1701),
.B(n_1743),
.Y(n_1875)
);

INVx1_ASAP7_75t_L g1876 ( 
.A(n_1757),
.Y(n_1876)
);

OR2x2_ASAP7_75t_L g1877 ( 
.A(n_1689),
.B(n_1790),
.Y(n_1877)
);

AO21x2_ASAP7_75t_L g1878 ( 
.A1(n_1753),
.A2(n_1776),
.B(n_1762),
.Y(n_1878)
);

OAI21x1_ASAP7_75t_L g1879 ( 
.A1(n_1777),
.A2(n_1786),
.B(n_1730),
.Y(n_1879)
);

BUFx2_ASAP7_75t_L g1880 ( 
.A(n_1750),
.Y(n_1880)
);

INVx2_ASAP7_75t_L g1881 ( 
.A(n_1710),
.Y(n_1881)
);

CKINVDCx20_ASAP7_75t_R g1882 ( 
.A(n_1706),
.Y(n_1882)
);

NAND2xp5_ASAP7_75t_L g1883 ( 
.A(n_1689),
.B(n_1797),
.Y(n_1883)
);

AND2x4_ASAP7_75t_L g1884 ( 
.A(n_1815),
.B(n_1684),
.Y(n_1884)
);

INVx1_ASAP7_75t_L g1885 ( 
.A(n_1733),
.Y(n_1885)
);

BUFx3_ASAP7_75t_L g1886 ( 
.A(n_1712),
.Y(n_1886)
);

NAND2xp5_ASAP7_75t_L g1887 ( 
.A(n_1804),
.B(n_1705),
.Y(n_1887)
);

OA21x2_ASAP7_75t_L g1888 ( 
.A1(n_1792),
.A2(n_1776),
.B(n_1786),
.Y(n_1888)
);

INVx2_ASAP7_75t_L g1889 ( 
.A(n_1720),
.Y(n_1889)
);

AOI22xp33_ASAP7_75t_SL g1890 ( 
.A1(n_1790),
.A2(n_1755),
.B1(n_1773),
.B2(n_1705),
.Y(n_1890)
);

OA21x2_ASAP7_75t_L g1891 ( 
.A1(n_1761),
.A2(n_1788),
.B(n_1791),
.Y(n_1891)
);

AOI21x1_ASAP7_75t_L g1892 ( 
.A1(n_1783),
.A2(n_1778),
.B(n_1780),
.Y(n_1892)
);

AO21x2_ASAP7_75t_L g1893 ( 
.A1(n_1765),
.A2(n_1772),
.B(n_1741),
.Y(n_1893)
);

INVx1_ASAP7_75t_L g1894 ( 
.A(n_1720),
.Y(n_1894)
);

AND2x2_ASAP7_75t_L g1895 ( 
.A(n_1696),
.B(n_1771),
.Y(n_1895)
);

BUFx2_ASAP7_75t_L g1896 ( 
.A(n_1787),
.Y(n_1896)
);

INVx2_ASAP7_75t_L g1897 ( 
.A(n_1802),
.Y(n_1897)
);

INVx2_ASAP7_75t_L g1898 ( 
.A(n_1802),
.Y(n_1898)
);

OR2x2_ASAP7_75t_L g1899 ( 
.A(n_1719),
.B(n_1772),
.Y(n_1899)
);

INVx1_ASAP7_75t_L g1900 ( 
.A(n_1764),
.Y(n_1900)
);

BUFx2_ASAP7_75t_L g1901 ( 
.A(n_1743),
.Y(n_1901)
);

INVx1_ASAP7_75t_L g1902 ( 
.A(n_1846),
.Y(n_1902)
);

INVx2_ASAP7_75t_L g1903 ( 
.A(n_1881),
.Y(n_1903)
);

HB1xp67_ASAP7_75t_L g1904 ( 
.A(n_1894),
.Y(n_1904)
);

AND2x4_ASAP7_75t_L g1905 ( 
.A(n_1845),
.B(n_1759),
.Y(n_1905)
);

INVx1_ASAP7_75t_L g1906 ( 
.A(n_1846),
.Y(n_1906)
);

HB1xp67_ASAP7_75t_L g1907 ( 
.A(n_1894),
.Y(n_1907)
);

NOR4xp25_ASAP7_75t_SL g1908 ( 
.A(n_1816),
.B(n_1860),
.C(n_1901),
.D(n_1896),
.Y(n_1908)
);

OR2x2_ASAP7_75t_L g1909 ( 
.A(n_1877),
.B(n_1782),
.Y(n_1909)
);

INVx3_ASAP7_75t_L g1910 ( 
.A(n_1850),
.Y(n_1910)
);

AND2x2_ASAP7_75t_L g1911 ( 
.A(n_1871),
.B(n_1781),
.Y(n_1911)
);

NAND2xp5_ASAP7_75t_L g1912 ( 
.A(n_1877),
.B(n_1699),
.Y(n_1912)
);

NAND2xp5_ASAP7_75t_L g1913 ( 
.A(n_1831),
.B(n_1848),
.Y(n_1913)
);

AND2x2_ASAP7_75t_L g1914 ( 
.A(n_1840),
.B(n_1848),
.Y(n_1914)
);

AND2x2_ASAP7_75t_L g1915 ( 
.A(n_1840),
.B(n_1729),
.Y(n_1915)
);

INVx2_ASAP7_75t_L g1916 ( 
.A(n_1889),
.Y(n_1916)
);

HB1xp67_ASAP7_75t_L g1917 ( 
.A(n_1897),
.Y(n_1917)
);

INVx1_ASAP7_75t_L g1918 ( 
.A(n_1851),
.Y(n_1918)
);

NAND2xp5_ASAP7_75t_L g1919 ( 
.A(n_1819),
.B(n_1827),
.Y(n_1919)
);

BUFx2_ASAP7_75t_L g1920 ( 
.A(n_1880),
.Y(n_1920)
);

AND2x2_ASAP7_75t_L g1921 ( 
.A(n_1845),
.B(n_1729),
.Y(n_1921)
);

OAI221xp5_ASAP7_75t_L g1922 ( 
.A1(n_1859),
.A2(n_1690),
.B1(n_1755),
.B2(n_1770),
.C(n_1718),
.Y(n_1922)
);

NAND2xp5_ASAP7_75t_L g1923 ( 
.A(n_1855),
.B(n_1774),
.Y(n_1923)
);

AND2x2_ASAP7_75t_L g1924 ( 
.A(n_1823),
.B(n_1736),
.Y(n_1924)
);

OR2x2_ASAP7_75t_L g1925 ( 
.A(n_1820),
.B(n_1774),
.Y(n_1925)
);

INVx3_ASAP7_75t_L g1926 ( 
.A(n_1850),
.Y(n_1926)
);

AOI22xp33_ASAP7_75t_L g1927 ( 
.A1(n_1829),
.A2(n_1838),
.B1(n_1825),
.B2(n_1861),
.Y(n_1927)
);

AOI22xp33_ASAP7_75t_L g1928 ( 
.A1(n_1861),
.A2(n_1716),
.B1(n_1734),
.B2(n_1749),
.Y(n_1928)
);

AND2x2_ASAP7_75t_L g1929 ( 
.A(n_1823),
.B(n_1736),
.Y(n_1929)
);

NAND2xp5_ASAP7_75t_SL g1930 ( 
.A(n_1841),
.B(n_1740),
.Y(n_1930)
);

BUFx2_ASAP7_75t_L g1931 ( 
.A(n_1880),
.Y(n_1931)
);

AND2x2_ASAP7_75t_L g1932 ( 
.A(n_1864),
.B(n_1766),
.Y(n_1932)
);

AND2x2_ASAP7_75t_L g1933 ( 
.A(n_1864),
.B(n_1766),
.Y(n_1933)
);

AOI22xp33_ASAP7_75t_L g1934 ( 
.A1(n_1834),
.A2(n_1716),
.B1(n_1744),
.B2(n_1760),
.Y(n_1934)
);

INVxp67_ASAP7_75t_SL g1935 ( 
.A(n_1898),
.Y(n_1935)
);

NAND2xp5_ASAP7_75t_L g1936 ( 
.A(n_1817),
.B(n_1761),
.Y(n_1936)
);

HB1xp67_ASAP7_75t_L g1937 ( 
.A(n_1860),
.Y(n_1937)
);

BUFx2_ASAP7_75t_L g1938 ( 
.A(n_1896),
.Y(n_1938)
);

NAND2xp5_ASAP7_75t_L g1939 ( 
.A(n_1821),
.B(n_1723),
.Y(n_1939)
);

AND2x2_ASAP7_75t_L g1940 ( 
.A(n_1895),
.B(n_1763),
.Y(n_1940)
);

BUFx3_ASAP7_75t_L g1941 ( 
.A(n_1816),
.Y(n_1941)
);

AND2x2_ASAP7_75t_L g1942 ( 
.A(n_1869),
.B(n_1709),
.Y(n_1942)
);

OR2x2_ASAP7_75t_L g1943 ( 
.A(n_1853),
.B(n_1745),
.Y(n_1943)
);

NAND2xp5_ASAP7_75t_L g1944 ( 
.A(n_1826),
.B(n_1798),
.Y(n_1944)
);

BUFx2_ASAP7_75t_L g1945 ( 
.A(n_1858),
.Y(n_1945)
);

OR2x2_ASAP7_75t_L g1946 ( 
.A(n_1853),
.B(n_1814),
.Y(n_1946)
);

INVx2_ASAP7_75t_L g1947 ( 
.A(n_1874),
.Y(n_1947)
);

INVx1_ASAP7_75t_L g1948 ( 
.A(n_1872),
.Y(n_1948)
);

BUFx3_ASAP7_75t_L g1949 ( 
.A(n_1833),
.Y(n_1949)
);

OR2x2_ASAP7_75t_L g1950 ( 
.A(n_1899),
.B(n_1813),
.Y(n_1950)
);

NAND2xp5_ASAP7_75t_L g1951 ( 
.A(n_1826),
.B(n_1703),
.Y(n_1951)
);

AOI22xp33_ASAP7_75t_SL g1952 ( 
.A1(n_1912),
.A2(n_1834),
.B1(n_1900),
.B2(n_1867),
.Y(n_1952)
);

AO21x2_ASAP7_75t_L g1953 ( 
.A1(n_1912),
.A2(n_1892),
.B(n_1867),
.Y(n_1953)
);

INVx1_ASAP7_75t_L g1954 ( 
.A(n_1902),
.Y(n_1954)
);

INVx1_ASAP7_75t_SL g1955 ( 
.A(n_1949),
.Y(n_1955)
);

OAI221xp5_ASAP7_75t_L g1956 ( 
.A1(n_1927),
.A2(n_1890),
.B1(n_1834),
.B2(n_1900),
.C(n_1849),
.Y(n_1956)
);

AOI211xp5_ASAP7_75t_L g1957 ( 
.A1(n_1922),
.A2(n_1868),
.B(n_1879),
.C(n_1830),
.Y(n_1957)
);

BUFx3_ASAP7_75t_L g1958 ( 
.A(n_1949),
.Y(n_1958)
);

INVx1_ASAP7_75t_L g1959 ( 
.A(n_1902),
.Y(n_1959)
);

HB1xp67_ASAP7_75t_L g1960 ( 
.A(n_1904),
.Y(n_1960)
);

BUFx3_ASAP7_75t_L g1961 ( 
.A(n_1949),
.Y(n_1961)
);

NAND2xp5_ASAP7_75t_L g1962 ( 
.A(n_1919),
.B(n_1914),
.Y(n_1962)
);

NOR4xp25_ASAP7_75t_SL g1963 ( 
.A(n_1930),
.B(n_1901),
.C(n_1870),
.D(n_1885),
.Y(n_1963)
);

BUFx2_ASAP7_75t_L g1964 ( 
.A(n_1941),
.Y(n_1964)
);

AOI221xp5_ASAP7_75t_SL g1965 ( 
.A1(n_1922),
.A2(n_1854),
.B1(n_1832),
.B2(n_1887),
.C(n_1883),
.Y(n_1965)
);

AND2x2_ASAP7_75t_L g1966 ( 
.A(n_1914),
.B(n_1843),
.Y(n_1966)
);

NOR2xp33_ASAP7_75t_R g1967 ( 
.A(n_1941),
.B(n_1882),
.Y(n_1967)
);

AND2x4_ASAP7_75t_L g1968 ( 
.A(n_1914),
.B(n_1858),
.Y(n_1968)
);

OAI33xp33_ASAP7_75t_L g1969 ( 
.A1(n_1944),
.A2(n_1830),
.A3(n_1842),
.B1(n_1837),
.B2(n_1899),
.B3(n_1839),
.Y(n_1969)
);

INVx1_ASAP7_75t_L g1970 ( 
.A(n_1906),
.Y(n_1970)
);

OAI22xp33_ASAP7_75t_L g1971 ( 
.A1(n_1946),
.A2(n_1828),
.B1(n_1862),
.B2(n_1875),
.Y(n_1971)
);

BUFx6f_ASAP7_75t_L g1972 ( 
.A(n_1938),
.Y(n_1972)
);

OAI22xp5_ASAP7_75t_L g1973 ( 
.A1(n_1928),
.A2(n_1862),
.B1(n_1828),
.B2(n_1875),
.Y(n_1973)
);

NOR2x1_ASAP7_75t_L g1974 ( 
.A(n_1950),
.B(n_1886),
.Y(n_1974)
);

NOR2x2_ASAP7_75t_L g1975 ( 
.A(n_1947),
.B(n_1866),
.Y(n_1975)
);

INVx1_ASAP7_75t_L g1976 ( 
.A(n_1906),
.Y(n_1976)
);

BUFx3_ASAP7_75t_L g1977 ( 
.A(n_1942),
.Y(n_1977)
);

AOI222xp33_ASAP7_75t_L g1978 ( 
.A1(n_1936),
.A2(n_1873),
.B1(n_1856),
.B2(n_1847),
.C1(n_1876),
.C2(n_1835),
.Y(n_1978)
);

INVxp67_ASAP7_75t_SL g1979 ( 
.A(n_1917),
.Y(n_1979)
);

NOR2xp33_ASAP7_75t_R g1980 ( 
.A(n_1946),
.B(n_1833),
.Y(n_1980)
);

HB1xp67_ASAP7_75t_L g1981 ( 
.A(n_1904),
.Y(n_1981)
);

NOR2xp33_ASAP7_75t_L g1982 ( 
.A(n_1939),
.B(n_1844),
.Y(n_1982)
);

NOR2xp33_ASAP7_75t_L g1983 ( 
.A(n_1939),
.B(n_1886),
.Y(n_1983)
);

AOI22xp33_ASAP7_75t_SL g1984 ( 
.A1(n_1915),
.A2(n_1867),
.B1(n_1878),
.B2(n_1849),
.Y(n_1984)
);

AO21x1_ASAP7_75t_SL g1985 ( 
.A1(n_1909),
.A2(n_1857),
.B(n_1865),
.Y(n_1985)
);

AND2x6_ASAP7_75t_SL g1986 ( 
.A(n_1942),
.B(n_1828),
.Y(n_1986)
);

INVx1_ASAP7_75t_L g1987 ( 
.A(n_1918),
.Y(n_1987)
);

NAND2xp33_ASAP7_75t_R g1988 ( 
.A(n_1908),
.B(n_1849),
.Y(n_1988)
);

AOI21xp5_ASAP7_75t_SL g1989 ( 
.A1(n_1943),
.A2(n_1878),
.B(n_1818),
.Y(n_1989)
);

AOI21xp5_ASAP7_75t_L g1990 ( 
.A1(n_1908),
.A2(n_1868),
.B(n_1878),
.Y(n_1990)
);

BUFx3_ASAP7_75t_L g1991 ( 
.A(n_1942),
.Y(n_1991)
);

INVx1_ASAP7_75t_L g1992 ( 
.A(n_1918),
.Y(n_1992)
);

AO21x2_ASAP7_75t_L g1993 ( 
.A1(n_1935),
.A2(n_1892),
.B(n_1822),
.Y(n_1993)
);

OR2x6_ASAP7_75t_L g1994 ( 
.A(n_1943),
.B(n_1818),
.Y(n_1994)
);

AND2x2_ASAP7_75t_L g1995 ( 
.A(n_1945),
.B(n_1852),
.Y(n_1995)
);

HB1xp67_ASAP7_75t_L g1996 ( 
.A(n_1907),
.Y(n_1996)
);

NAND3xp33_ASAP7_75t_L g1997 ( 
.A(n_1950),
.B(n_1888),
.C(n_1891),
.Y(n_1997)
);

OAI221xp5_ASAP7_75t_L g1998 ( 
.A1(n_1937),
.A2(n_1951),
.B1(n_1950),
.B2(n_1936),
.C(n_1935),
.Y(n_1998)
);

OAI31xp33_ASAP7_75t_SL g1999 ( 
.A1(n_1915),
.A2(n_1879),
.A3(n_1858),
.B(n_1884),
.Y(n_1999)
);

AOI221xp5_ASAP7_75t_L g2000 ( 
.A1(n_1937),
.A2(n_1893),
.B1(n_1824),
.B2(n_1863),
.C(n_1836),
.Y(n_2000)
);

INVx3_ASAP7_75t_L g2001 ( 
.A(n_1905),
.Y(n_2001)
);

AOI22xp33_ASAP7_75t_L g2002 ( 
.A1(n_1915),
.A2(n_1893),
.B1(n_1822),
.B2(n_1863),
.Y(n_2002)
);

AND2x2_ASAP7_75t_L g2003 ( 
.A(n_1985),
.B(n_1932),
.Y(n_2003)
);

INVx2_ASAP7_75t_L g2004 ( 
.A(n_1993),
.Y(n_2004)
);

OAI21xp5_ASAP7_75t_SL g2005 ( 
.A1(n_1952),
.A2(n_1934),
.B(n_1933),
.Y(n_2005)
);

OA21x2_ASAP7_75t_L g2006 ( 
.A1(n_1990),
.A2(n_1921),
.B(n_1916),
.Y(n_2006)
);

INVx2_ASAP7_75t_L g2007 ( 
.A(n_1993),
.Y(n_2007)
);

BUFx3_ASAP7_75t_L g2008 ( 
.A(n_1953),
.Y(n_2008)
);

INVx1_ASAP7_75t_L g2009 ( 
.A(n_1954),
.Y(n_2009)
);

INVx1_ASAP7_75t_L g2010 ( 
.A(n_1959),
.Y(n_2010)
);

OAI21xp5_ASAP7_75t_L g2011 ( 
.A1(n_1957),
.A2(n_1909),
.B(n_1932),
.Y(n_2011)
);

AND2x4_ASAP7_75t_L g2012 ( 
.A(n_2001),
.B(n_1968),
.Y(n_2012)
);

OAI21x1_ASAP7_75t_L g2013 ( 
.A1(n_1989),
.A2(n_1910),
.B(n_1926),
.Y(n_2013)
);

AND2x2_ASAP7_75t_L g2014 ( 
.A(n_1999),
.B(n_1932),
.Y(n_2014)
);

HB1xp67_ASAP7_75t_L g2015 ( 
.A(n_1960),
.Y(n_2015)
);

INVx1_ASAP7_75t_L g2016 ( 
.A(n_1970),
.Y(n_2016)
);

NAND2xp5_ASAP7_75t_L g2017 ( 
.A(n_1962),
.B(n_1913),
.Y(n_2017)
);

INVx2_ASAP7_75t_L g2018 ( 
.A(n_1953),
.Y(n_2018)
);

INVxp67_ASAP7_75t_SL g2019 ( 
.A(n_1997),
.Y(n_2019)
);

INVx1_ASAP7_75t_L g2020 ( 
.A(n_1976),
.Y(n_2020)
);

INVx1_ASAP7_75t_L g2021 ( 
.A(n_1987),
.Y(n_2021)
);

AND2x2_ASAP7_75t_L g2022 ( 
.A(n_1968),
.B(n_1933),
.Y(n_2022)
);

NAND2xp5_ASAP7_75t_L g2023 ( 
.A(n_1965),
.B(n_1913),
.Y(n_2023)
);

INVx2_ASAP7_75t_L g2024 ( 
.A(n_1960),
.Y(n_2024)
);

INVx1_ASAP7_75t_L g2025 ( 
.A(n_1992),
.Y(n_2025)
);

INVx2_ASAP7_75t_L g2026 ( 
.A(n_1981),
.Y(n_2026)
);

OA21x2_ASAP7_75t_L g2027 ( 
.A1(n_2002),
.A2(n_1921),
.B(n_1903),
.Y(n_2027)
);

AND2x2_ASAP7_75t_L g2028 ( 
.A(n_1966),
.B(n_1933),
.Y(n_2028)
);

BUFx3_ASAP7_75t_L g2029 ( 
.A(n_1972),
.Y(n_2029)
);

INVx4_ASAP7_75t_SL g2030 ( 
.A(n_1958),
.Y(n_2030)
);

INVx4_ASAP7_75t_SL g2031 ( 
.A(n_1961),
.Y(n_2031)
);

OR2x2_ASAP7_75t_L g2032 ( 
.A(n_1996),
.B(n_1909),
.Y(n_2032)
);

INVx3_ASAP7_75t_L g2033 ( 
.A(n_1986),
.Y(n_2033)
);

INVx1_ASAP7_75t_SL g2034 ( 
.A(n_1967),
.Y(n_2034)
);

AND2x2_ASAP7_75t_L g2035 ( 
.A(n_1974),
.B(n_1920),
.Y(n_2035)
);

AND2x2_ASAP7_75t_L g2036 ( 
.A(n_1964),
.B(n_1920),
.Y(n_2036)
);

NAND2xp5_ASAP7_75t_L g2037 ( 
.A(n_1979),
.B(n_1948),
.Y(n_2037)
);

OA21x2_ASAP7_75t_L g2038 ( 
.A1(n_2002),
.A2(n_1921),
.B(n_1903),
.Y(n_2038)
);

NAND2xp5_ASAP7_75t_SL g2039 ( 
.A(n_1980),
.B(n_1931),
.Y(n_2039)
);

INVx2_ASAP7_75t_SL g2040 ( 
.A(n_1972),
.Y(n_2040)
);

HB1xp67_ASAP7_75t_L g2041 ( 
.A(n_1998),
.Y(n_2041)
);

INVx1_ASAP7_75t_L g2042 ( 
.A(n_1978),
.Y(n_2042)
);

INVx1_ASAP7_75t_SL g2043 ( 
.A(n_1955),
.Y(n_2043)
);

NAND2xp33_ASAP7_75t_R g2044 ( 
.A(n_1963),
.B(n_1910),
.Y(n_2044)
);

INVx1_ASAP7_75t_L g2045 ( 
.A(n_2009),
.Y(n_2045)
);

OAI31xp33_ASAP7_75t_L g2046 ( 
.A1(n_2005),
.A2(n_1956),
.A3(n_1971),
.B(n_1973),
.Y(n_2046)
);

INVx1_ASAP7_75t_L g2047 ( 
.A(n_2009),
.Y(n_2047)
);

INVx2_ASAP7_75t_L g2048 ( 
.A(n_2008),
.Y(n_2048)
);

BUFx2_ASAP7_75t_L g2049 ( 
.A(n_2019),
.Y(n_2049)
);

INVx2_ASAP7_75t_SL g2050 ( 
.A(n_2034),
.Y(n_2050)
);

INVx1_ASAP7_75t_L g2051 ( 
.A(n_2010),
.Y(n_2051)
);

AND2x2_ASAP7_75t_L g2052 ( 
.A(n_2003),
.B(n_2014),
.Y(n_2052)
);

AND2x4_ASAP7_75t_L g2053 ( 
.A(n_2030),
.B(n_1994),
.Y(n_2053)
);

AND2x2_ASAP7_75t_L g2054 ( 
.A(n_2003),
.B(n_1977),
.Y(n_2054)
);

INVx1_ASAP7_75t_L g2055 ( 
.A(n_2010),
.Y(n_2055)
);

AND2x2_ASAP7_75t_SL g2056 ( 
.A(n_2041),
.B(n_2033),
.Y(n_2056)
);

AND2x2_ASAP7_75t_L g2057 ( 
.A(n_2014),
.B(n_1991),
.Y(n_2057)
);

INVx6_ASAP7_75t_L g2058 ( 
.A(n_2030),
.Y(n_2058)
);

AND2x2_ASAP7_75t_L g2059 ( 
.A(n_2014),
.B(n_1995),
.Y(n_2059)
);

AND2x2_ASAP7_75t_SL g2060 ( 
.A(n_2041),
.B(n_2000),
.Y(n_2060)
);

AND2x4_ASAP7_75t_SL g2061 ( 
.A(n_2033),
.B(n_1994),
.Y(n_2061)
);

INVx1_ASAP7_75t_L g2062 ( 
.A(n_2016),
.Y(n_2062)
);

INVxp67_ASAP7_75t_L g2063 ( 
.A(n_2034),
.Y(n_2063)
);

INVx2_ASAP7_75t_L g2064 ( 
.A(n_2008),
.Y(n_2064)
);

INVx2_ASAP7_75t_L g2065 ( 
.A(n_2008),
.Y(n_2065)
);

NAND2xp5_ASAP7_75t_L g2066 ( 
.A(n_2019),
.B(n_1952),
.Y(n_2066)
);

OR2x2_ASAP7_75t_L g2067 ( 
.A(n_2023),
.B(n_1925),
.Y(n_2067)
);

NAND2xp33_ASAP7_75t_L g2068 ( 
.A(n_2011),
.B(n_1975),
.Y(n_2068)
);

NAND4xp25_ASAP7_75t_L g2069 ( 
.A(n_2011),
.B(n_1982),
.C(n_1984),
.D(n_1983),
.Y(n_2069)
);

INVx1_ASAP7_75t_L g2070 ( 
.A(n_2020),
.Y(n_2070)
);

INVx1_ASAP7_75t_L g2071 ( 
.A(n_2020),
.Y(n_2071)
);

NAND2xp5_ASAP7_75t_L g2072 ( 
.A(n_2023),
.B(n_1924),
.Y(n_2072)
);

AND2x4_ASAP7_75t_L g2073 ( 
.A(n_2030),
.B(n_1994),
.Y(n_2073)
);

INVxp67_ASAP7_75t_L g2074 ( 
.A(n_2043),
.Y(n_2074)
);

INVxp67_ASAP7_75t_L g2075 ( 
.A(n_2043),
.Y(n_2075)
);

AND2x4_ASAP7_75t_L g2076 ( 
.A(n_2031),
.B(n_1910),
.Y(n_2076)
);

INVx2_ASAP7_75t_L g2077 ( 
.A(n_2008),
.Y(n_2077)
);

AND2x2_ASAP7_75t_L g2078 ( 
.A(n_2031),
.B(n_1929),
.Y(n_2078)
);

AND2x2_ASAP7_75t_L g2079 ( 
.A(n_2031),
.B(n_1911),
.Y(n_2079)
);

INVx2_ASAP7_75t_L g2080 ( 
.A(n_2027),
.Y(n_2080)
);

NAND2xp5_ASAP7_75t_L g2081 ( 
.A(n_2017),
.B(n_1940),
.Y(n_2081)
);

AND2x2_ASAP7_75t_L g2082 ( 
.A(n_2031),
.B(n_1911),
.Y(n_2082)
);

NAND2xp5_ASAP7_75t_L g2083 ( 
.A(n_2017),
.B(n_1940),
.Y(n_2083)
);

NAND2xp5_ASAP7_75t_L g2084 ( 
.A(n_2042),
.B(n_1940),
.Y(n_2084)
);

NAND2xp5_ASAP7_75t_L g2085 ( 
.A(n_2042),
.B(n_2036),
.Y(n_2085)
);

OAI21xp33_ASAP7_75t_L g2086 ( 
.A1(n_2005),
.A2(n_1984),
.B(n_1923),
.Y(n_2086)
);

AND2x4_ASAP7_75t_SL g2087 ( 
.A(n_2033),
.B(n_1905),
.Y(n_2087)
);

AND2x2_ASAP7_75t_L g2088 ( 
.A(n_2057),
.B(n_2022),
.Y(n_2088)
);

AND2x4_ASAP7_75t_L g2089 ( 
.A(n_2087),
.B(n_2033),
.Y(n_2089)
);

INVx2_ASAP7_75t_L g2090 ( 
.A(n_2080),
.Y(n_2090)
);

INVx1_ASAP7_75t_SL g2091 ( 
.A(n_2061),
.Y(n_2091)
);

AND2x2_ASAP7_75t_L g2092 ( 
.A(n_2057),
.B(n_2022),
.Y(n_2092)
);

NAND2xp5_ASAP7_75t_L g2093 ( 
.A(n_2074),
.B(n_2028),
.Y(n_2093)
);

INVx1_ASAP7_75t_L g2094 ( 
.A(n_2045),
.Y(n_2094)
);

AND2x4_ASAP7_75t_L g2095 ( 
.A(n_2087),
.B(n_2033),
.Y(n_2095)
);

AND2x2_ASAP7_75t_L g2096 ( 
.A(n_2052),
.B(n_2012),
.Y(n_2096)
);

NAND2xp5_ASAP7_75t_L g2097 ( 
.A(n_2075),
.B(n_2028),
.Y(n_2097)
);

AND2x2_ASAP7_75t_L g2098 ( 
.A(n_2052),
.B(n_2012),
.Y(n_2098)
);

INVx2_ASAP7_75t_L g2099 ( 
.A(n_2080),
.Y(n_2099)
);

NAND2xp5_ASAP7_75t_L g2100 ( 
.A(n_2049),
.B(n_2050),
.Y(n_2100)
);

OR2x2_ASAP7_75t_L g2101 ( 
.A(n_2085),
.B(n_2032),
.Y(n_2101)
);

INVxp67_ASAP7_75t_L g2102 ( 
.A(n_2050),
.Y(n_2102)
);

INVx1_ASAP7_75t_L g2103 ( 
.A(n_2045),
.Y(n_2103)
);

AOI21xp5_ASAP7_75t_L g2104 ( 
.A1(n_2068),
.A2(n_2039),
.B(n_1969),
.Y(n_2104)
);

AOI22xp5_ASAP7_75t_L g2105 ( 
.A1(n_2060),
.A2(n_2027),
.B1(n_2038),
.B2(n_1969),
.Y(n_2105)
);

AND2x2_ASAP7_75t_L g2106 ( 
.A(n_2053),
.B(n_2012),
.Y(n_2106)
);

NAND2xp5_ASAP7_75t_L g2107 ( 
.A(n_2049),
.B(n_2028),
.Y(n_2107)
);

INVx4_ASAP7_75t_L g2108 ( 
.A(n_2058),
.Y(n_2108)
);

INVx1_ASAP7_75t_L g2109 ( 
.A(n_2047),
.Y(n_2109)
);

NOR2xp33_ASAP7_75t_L g2110 ( 
.A(n_2063),
.B(n_2039),
.Y(n_2110)
);

AND2x4_ASAP7_75t_L g2111 ( 
.A(n_2061),
.B(n_2012),
.Y(n_2111)
);

NAND2xp5_ASAP7_75t_L g2112 ( 
.A(n_2060),
.B(n_2021),
.Y(n_2112)
);

INVx1_ASAP7_75t_L g2113 ( 
.A(n_2047),
.Y(n_2113)
);

INVx1_ASAP7_75t_L g2114 ( 
.A(n_2051),
.Y(n_2114)
);

NAND2xp5_ASAP7_75t_L g2115 ( 
.A(n_2060),
.B(n_2025),
.Y(n_2115)
);

AND2x2_ASAP7_75t_L g2116 ( 
.A(n_2053),
.B(n_2012),
.Y(n_2116)
);

NAND2x1_ASAP7_75t_L g2117 ( 
.A(n_2058),
.B(n_2079),
.Y(n_2117)
);

AND2x2_ASAP7_75t_L g2118 ( 
.A(n_2053),
.B(n_2029),
.Y(n_2118)
);

OR2x2_ASAP7_75t_L g2119 ( 
.A(n_2084),
.B(n_2032),
.Y(n_2119)
);

INVx2_ASAP7_75t_L g2120 ( 
.A(n_2048),
.Y(n_2120)
);

OR2x2_ASAP7_75t_L g2121 ( 
.A(n_2072),
.B(n_2024),
.Y(n_2121)
);

OAI221xp5_ASAP7_75t_L g2122 ( 
.A1(n_2066),
.A2(n_2027),
.B1(n_2038),
.B2(n_2044),
.C(n_2006),
.Y(n_2122)
);

NAND2xp5_ASAP7_75t_L g2123 ( 
.A(n_2056),
.B(n_2025),
.Y(n_2123)
);

AOI21xp33_ASAP7_75t_SL g2124 ( 
.A1(n_2056),
.A2(n_2044),
.B(n_2040),
.Y(n_2124)
);

HB1xp67_ASAP7_75t_L g2125 ( 
.A(n_2051),
.Y(n_2125)
);

OR2x2_ASAP7_75t_L g2126 ( 
.A(n_2067),
.B(n_2037),
.Y(n_2126)
);

OAI21xp33_ASAP7_75t_L g2127 ( 
.A1(n_2086),
.A2(n_2035),
.B(n_2024),
.Y(n_2127)
);

OAI221xp5_ASAP7_75t_L g2128 ( 
.A1(n_2068),
.A2(n_2046),
.B1(n_2069),
.B2(n_2027),
.C(n_2038),
.Y(n_2128)
);

INVx1_ASAP7_75t_SL g2129 ( 
.A(n_2089),
.Y(n_2129)
);

AND2x2_ASAP7_75t_L g2130 ( 
.A(n_2088),
.B(n_2058),
.Y(n_2130)
);

AND2x4_ASAP7_75t_L g2131 ( 
.A(n_2089),
.B(n_2073),
.Y(n_2131)
);

INVx2_ASAP7_75t_L g2132 ( 
.A(n_2096),
.Y(n_2132)
);

OR2x2_ASAP7_75t_L g2133 ( 
.A(n_2119),
.B(n_2067),
.Y(n_2133)
);

INVx1_ASAP7_75t_SL g2134 ( 
.A(n_2089),
.Y(n_2134)
);

AND2x4_ASAP7_75t_L g2135 ( 
.A(n_2095),
.B(n_2073),
.Y(n_2135)
);

AND2x2_ASAP7_75t_L g2136 ( 
.A(n_2088),
.B(n_2058),
.Y(n_2136)
);

NAND2xp5_ASAP7_75t_L g2137 ( 
.A(n_2102),
.B(n_2081),
.Y(n_2137)
);

NOR2x1_ASAP7_75t_L g2138 ( 
.A(n_2100),
.B(n_2073),
.Y(n_2138)
);

INVx1_ASAP7_75t_L g2139 ( 
.A(n_2125),
.Y(n_2139)
);

AND2x4_ASAP7_75t_SL g2140 ( 
.A(n_2095),
.B(n_2054),
.Y(n_2140)
);

INVx1_ASAP7_75t_L g2141 ( 
.A(n_2094),
.Y(n_2141)
);

INVx1_ASAP7_75t_L g2142 ( 
.A(n_2103),
.Y(n_2142)
);

INVx6_ASAP7_75t_L g2143 ( 
.A(n_2108),
.Y(n_2143)
);

INVx1_ASAP7_75t_L g2144 ( 
.A(n_2109),
.Y(n_2144)
);

AOI22xp33_ASAP7_75t_L g2145 ( 
.A1(n_2128),
.A2(n_2038),
.B1(n_2027),
.B2(n_2006),
.Y(n_2145)
);

HB1xp67_ASAP7_75t_L g2146 ( 
.A(n_2110),
.Y(n_2146)
);

OAI22xp33_ASAP7_75t_L g2147 ( 
.A1(n_2105),
.A2(n_1988),
.B1(n_2027),
.B2(n_2038),
.Y(n_2147)
);

INVx2_ASAP7_75t_L g2148 ( 
.A(n_2096),
.Y(n_2148)
);

INVx1_ASAP7_75t_L g2149 ( 
.A(n_2113),
.Y(n_2149)
);

NAND2xp5_ASAP7_75t_L g2150 ( 
.A(n_2112),
.B(n_2083),
.Y(n_2150)
);

INVx1_ASAP7_75t_L g2151 ( 
.A(n_2114),
.Y(n_2151)
);

NAND2xp5_ASAP7_75t_SL g2152 ( 
.A(n_2095),
.B(n_2076),
.Y(n_2152)
);

INVx1_ASAP7_75t_L g2153 ( 
.A(n_2120),
.Y(n_2153)
);

OR2x2_ASAP7_75t_L g2154 ( 
.A(n_2101),
.B(n_2055),
.Y(n_2154)
);

INVx1_ASAP7_75t_L g2155 ( 
.A(n_2120),
.Y(n_2155)
);

AND2x2_ASAP7_75t_L g2156 ( 
.A(n_2092),
.B(n_2079),
.Y(n_2156)
);

INVx1_ASAP7_75t_SL g2157 ( 
.A(n_2091),
.Y(n_2157)
);

AND2x2_ASAP7_75t_L g2158 ( 
.A(n_2092),
.B(n_2082),
.Y(n_2158)
);

AND2x2_ASAP7_75t_L g2159 ( 
.A(n_2140),
.B(n_2108),
.Y(n_2159)
);

INVx1_ASAP7_75t_SL g2160 ( 
.A(n_2146),
.Y(n_2160)
);

AOI22xp5_ASAP7_75t_L g2161 ( 
.A1(n_2145),
.A2(n_2122),
.B1(n_2127),
.B2(n_2104),
.Y(n_2161)
);

INVx2_ASAP7_75t_L g2162 ( 
.A(n_2130),
.Y(n_2162)
);

INVx1_ASAP7_75t_L g2163 ( 
.A(n_2142),
.Y(n_2163)
);

INVx1_ASAP7_75t_L g2164 ( 
.A(n_2142),
.Y(n_2164)
);

NAND2x1_ASAP7_75t_SL g2165 ( 
.A(n_2131),
.B(n_2108),
.Y(n_2165)
);

AOI211xp5_ASAP7_75t_L g2166 ( 
.A1(n_2147),
.A2(n_2124),
.B(n_2115),
.C(n_2110),
.Y(n_2166)
);

INVx1_ASAP7_75t_L g2167 ( 
.A(n_2144),
.Y(n_2167)
);

NAND2xp5_ASAP7_75t_L g2168 ( 
.A(n_2157),
.B(n_2129),
.Y(n_2168)
);

AND2x4_ASAP7_75t_L g2169 ( 
.A(n_2131),
.B(n_2111),
.Y(n_2169)
);

OA21x2_ASAP7_75t_L g2170 ( 
.A1(n_2139),
.A2(n_2064),
.B(n_2048),
.Y(n_2170)
);

OAI221xp5_ASAP7_75t_L g2171 ( 
.A1(n_2138),
.A2(n_2038),
.B1(n_2123),
.B2(n_2006),
.C(n_2090),
.Y(n_2171)
);

INVx1_ASAP7_75t_L g2172 ( 
.A(n_2144),
.Y(n_2172)
);

INVx1_ASAP7_75t_L g2173 ( 
.A(n_2151),
.Y(n_2173)
);

NAND2xp5_ASAP7_75t_L g2174 ( 
.A(n_2134),
.B(n_2093),
.Y(n_2174)
);

INVxp67_ASAP7_75t_L g2175 ( 
.A(n_2131),
.Y(n_2175)
);

OAI22xp5_ASAP7_75t_L g2176 ( 
.A1(n_2133),
.A2(n_2107),
.B1(n_2097),
.B2(n_2121),
.Y(n_2176)
);

AOI21xp33_ASAP7_75t_L g2177 ( 
.A1(n_2139),
.A2(n_2065),
.B(n_2064),
.Y(n_2177)
);

INVx1_ASAP7_75t_L g2178 ( 
.A(n_2151),
.Y(n_2178)
);

INVx1_ASAP7_75t_L g2179 ( 
.A(n_2153),
.Y(n_2179)
);

NAND2xp5_ASAP7_75t_L g2180 ( 
.A(n_2132),
.B(n_2126),
.Y(n_2180)
);

NAND2xp5_ASAP7_75t_L g2181 ( 
.A(n_2132),
.B(n_2090),
.Y(n_2181)
);

INVx3_ASAP7_75t_L g2182 ( 
.A(n_2169),
.Y(n_2182)
);

AND2x2_ASAP7_75t_L g2183 ( 
.A(n_2169),
.B(n_2140),
.Y(n_2183)
);

INVx1_ASAP7_75t_L g2184 ( 
.A(n_2168),
.Y(n_2184)
);

OR2x2_ASAP7_75t_L g2185 ( 
.A(n_2160),
.B(n_2133),
.Y(n_2185)
);

NAND2xp5_ASAP7_75t_L g2186 ( 
.A(n_2160),
.B(n_2148),
.Y(n_2186)
);

NOR2xp67_ASAP7_75t_L g2187 ( 
.A(n_2175),
.B(n_2135),
.Y(n_2187)
);

AOI22xp33_ASAP7_75t_L g2188 ( 
.A1(n_2161),
.A2(n_2099),
.B1(n_2155),
.B2(n_2150),
.Y(n_2188)
);

INVx1_ASAP7_75t_L g2189 ( 
.A(n_2181),
.Y(n_2189)
);

NAND2xp5_ASAP7_75t_L g2190 ( 
.A(n_2162),
.B(n_2148),
.Y(n_2190)
);

INVxp33_ASAP7_75t_L g2191 ( 
.A(n_2165),
.Y(n_2191)
);

NOR2xp33_ASAP7_75t_L g2192 ( 
.A(n_2159),
.B(n_2143),
.Y(n_2192)
);

NAND2xp5_ASAP7_75t_L g2193 ( 
.A(n_2176),
.B(n_2154),
.Y(n_2193)
);

INVx1_ASAP7_75t_L g2194 ( 
.A(n_2163),
.Y(n_2194)
);

AOI22xp33_ASAP7_75t_L g2195 ( 
.A1(n_2171),
.A2(n_2099),
.B1(n_2065),
.B2(n_2077),
.Y(n_2195)
);

INVx1_ASAP7_75t_L g2196 ( 
.A(n_2164),
.Y(n_2196)
);

AND2x2_ASAP7_75t_L g2197 ( 
.A(n_2180),
.B(n_2135),
.Y(n_2197)
);

AOI22xp5_ASAP7_75t_L g2198 ( 
.A1(n_2195),
.A2(n_2188),
.B1(n_2166),
.B2(n_2170),
.Y(n_2198)
);

OAI211xp5_ASAP7_75t_L g2199 ( 
.A1(n_2193),
.A2(n_2188),
.B(n_2195),
.C(n_2187),
.Y(n_2199)
);

AOI21xp5_ASAP7_75t_L g2200 ( 
.A1(n_2191),
.A2(n_2170),
.B(n_2177),
.Y(n_2200)
);

OAI21xp5_ASAP7_75t_L g2201 ( 
.A1(n_2191),
.A2(n_2177),
.B(n_2174),
.Y(n_2201)
);

OAI221xp5_ASAP7_75t_SL g2202 ( 
.A1(n_2185),
.A2(n_2179),
.B1(n_2178),
.B2(n_2167),
.C(n_2173),
.Y(n_2202)
);

OAI22xp33_ASAP7_75t_L g2203 ( 
.A1(n_2186),
.A2(n_2006),
.B1(n_2117),
.B2(n_2121),
.Y(n_2203)
);

AOI21xp5_ASAP7_75t_L g2204 ( 
.A1(n_2190),
.A2(n_2152),
.B(n_2176),
.Y(n_2204)
);

NAND3x1_ASAP7_75t_L g2205 ( 
.A(n_2182),
.B(n_2172),
.C(n_2136),
.Y(n_2205)
);

OAI21xp33_ASAP7_75t_L g2206 ( 
.A1(n_2197),
.A2(n_2136),
.B(n_2130),
.Y(n_2206)
);

NOR2x1_ASAP7_75t_L g2207 ( 
.A(n_2182),
.B(n_2135),
.Y(n_2207)
);

OAI21xp33_ASAP7_75t_L g2208 ( 
.A1(n_2192),
.A2(n_2184),
.B(n_2183),
.Y(n_2208)
);

NAND3xp33_ASAP7_75t_L g2209 ( 
.A(n_2192),
.B(n_2189),
.C(n_2194),
.Y(n_2209)
);

NOR2xp33_ASAP7_75t_L g2210 ( 
.A(n_2196),
.B(n_2143),
.Y(n_2210)
);

OAI221xp5_ASAP7_75t_L g2211 ( 
.A1(n_2198),
.A2(n_2077),
.B1(n_2143),
.B2(n_2137),
.C(n_2154),
.Y(n_2211)
);

BUFx2_ASAP7_75t_L g2212 ( 
.A(n_2207),
.Y(n_2212)
);

OAI22xp33_ASAP7_75t_L g2213 ( 
.A1(n_2200),
.A2(n_2201),
.B1(n_2203),
.B2(n_2204),
.Y(n_2213)
);

CKINVDCx20_ASAP7_75t_R g2214 ( 
.A(n_2208),
.Y(n_2214)
);

AO22x1_ASAP7_75t_L g2215 ( 
.A1(n_2210),
.A2(n_2111),
.B1(n_2149),
.B2(n_2141),
.Y(n_2215)
);

INVxp67_ASAP7_75t_SL g2216 ( 
.A(n_2205),
.Y(n_2216)
);

INVx1_ASAP7_75t_L g2217 ( 
.A(n_2209),
.Y(n_2217)
);

AOI21xp33_ASAP7_75t_R g2218 ( 
.A1(n_2202),
.A2(n_2143),
.B(n_2026),
.Y(n_2218)
);

XNOR2x1_ASAP7_75t_L g2219 ( 
.A(n_2199),
.B(n_2111),
.Y(n_2219)
);

OR2x2_ASAP7_75t_L g2220 ( 
.A(n_2217),
.B(n_2206),
.Y(n_2220)
);

INVx1_ASAP7_75t_L g2221 ( 
.A(n_2212),
.Y(n_2221)
);

AND2x2_ASAP7_75t_L g2222 ( 
.A(n_2216),
.B(n_2156),
.Y(n_2222)
);

INVxp67_ASAP7_75t_SL g2223 ( 
.A(n_2219),
.Y(n_2223)
);

NAND2xp5_ASAP7_75t_L g2224 ( 
.A(n_2218),
.B(n_2215),
.Y(n_2224)
);

INVx1_ASAP7_75t_L g2225 ( 
.A(n_2214),
.Y(n_2225)
);

INVx1_ASAP7_75t_L g2226 ( 
.A(n_2211),
.Y(n_2226)
);

AOI221xp5_ASAP7_75t_L g2227 ( 
.A1(n_2213),
.A2(n_2004),
.B1(n_2007),
.B2(n_2018),
.C(n_2156),
.Y(n_2227)
);

NAND4xp75_ASAP7_75t_L g2228 ( 
.A(n_2221),
.B(n_2118),
.C(n_2158),
.D(n_2116),
.Y(n_2228)
);

NOR3x1_ASAP7_75t_L g2229 ( 
.A(n_2224),
.B(n_2040),
.C(n_2013),
.Y(n_2229)
);

INVx1_ASAP7_75t_L g2230 ( 
.A(n_2222),
.Y(n_2230)
);

NAND2xp5_ASAP7_75t_L g2231 ( 
.A(n_2223),
.B(n_2158),
.Y(n_2231)
);

OAI211xp5_ASAP7_75t_L g2232 ( 
.A1(n_2224),
.A2(n_2118),
.B(n_2106),
.C(n_2116),
.Y(n_2232)
);

INVx1_ASAP7_75t_L g2233 ( 
.A(n_2225),
.Y(n_2233)
);

INVx1_ASAP7_75t_L g2234 ( 
.A(n_2231),
.Y(n_2234)
);

NOR3xp33_ASAP7_75t_L g2235 ( 
.A(n_2230),
.B(n_2226),
.C(n_2220),
.Y(n_2235)
);

INVx1_ASAP7_75t_L g2236 ( 
.A(n_2233),
.Y(n_2236)
);

NOR3xp33_ASAP7_75t_L g2237 ( 
.A(n_2235),
.B(n_2232),
.C(n_2227),
.Y(n_2237)
);

NAND3xp33_ASAP7_75t_L g2238 ( 
.A(n_2237),
.B(n_2234),
.C(n_2236),
.Y(n_2238)
);

INVx2_ASAP7_75t_L g2239 ( 
.A(n_2238),
.Y(n_2239)
);

NOR2xp67_ASAP7_75t_L g2240 ( 
.A(n_2238),
.B(n_2228),
.Y(n_2240)
);

INVx1_ASAP7_75t_L g2241 ( 
.A(n_2239),
.Y(n_2241)
);

AOI21xp5_ASAP7_75t_L g2242 ( 
.A1(n_2240),
.A2(n_2229),
.B(n_2106),
.Y(n_2242)
);

OAI22xp5_ASAP7_75t_L g2243 ( 
.A1(n_2242),
.A2(n_2098),
.B1(n_2059),
.B2(n_2062),
.Y(n_2243)
);

OAI21xp5_ASAP7_75t_L g2244 ( 
.A1(n_2241),
.A2(n_2007),
.B(n_2004),
.Y(n_2244)
);

AOI22xp33_ASAP7_75t_SL g2245 ( 
.A1(n_2243),
.A2(n_2244),
.B1(n_2007),
.B2(n_2004),
.Y(n_2245)
);

OAI21xp5_ASAP7_75t_SL g2246 ( 
.A1(n_2245),
.A2(n_2098),
.B(n_2076),
.Y(n_2246)
);

OR2x6_ASAP7_75t_L g2247 ( 
.A(n_2246),
.B(n_2040),
.Y(n_2247)
);

AOI222xp33_ASAP7_75t_L g2248 ( 
.A1(n_2247),
.A2(n_2018),
.B1(n_2007),
.B2(n_2004),
.C1(n_2076),
.C2(n_2078),
.Y(n_2248)
);

OAI22xp33_ASAP7_75t_L g2249 ( 
.A1(n_2248),
.A2(n_2070),
.B1(n_2071),
.B2(n_2062),
.Y(n_2249)
);

AOI211xp5_ASAP7_75t_L g2250 ( 
.A1(n_2249),
.A2(n_2018),
.B(n_2015),
.C(n_2013),
.Y(n_2250)
);


endmodule