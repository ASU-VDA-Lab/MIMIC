module fake_netlist_5_1678_n_1144 (n_137, n_210, n_168, n_164, n_191, n_91, n_208, n_82, n_122, n_194, n_142, n_176, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_182, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_180, n_184, n_65, n_78, n_74, n_144, n_207, n_114, n_57, n_96, n_37, n_189, n_165, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_177, n_60, n_155, n_152, n_197, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_195, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_203, n_205, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_179, n_125, n_35, n_167, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_202, n_130, n_157, n_29, n_79, n_193, n_131, n_151, n_47, n_173, n_192, n_25, n_53, n_160, n_198, n_188, n_190, n_8, n_201, n_158, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_159, n_163, n_95, n_119, n_183, n_185, n_175, n_169, n_59, n_26, n_133, n_55, n_196, n_99, n_2, n_211, n_181, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_178, n_12, n_67, n_121, n_36, n_76, n_200, n_87, n_150, n_162, n_27, n_170, n_64, n_77, n_102, n_106, n_161, n_209, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_174, n_186, n_199, n_134, n_187, n_32, n_41, n_104, n_172, n_103, n_56, n_51, n_63, n_97, n_141, n_166, n_11, n_206, n_171, n_153, n_7, n_15, n_145, n_48, n_204, n_50, n_52, n_88, n_110, n_1144);

input n_137;
input n_210;
input n_168;
input n_164;
input n_191;
input n_91;
input n_208;
input n_82;
input n_122;
input n_194;
input n_142;
input n_176;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_182;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_180;
input n_184;
input n_65;
input n_78;
input n_74;
input n_144;
input n_207;
input n_114;
input n_57;
input n_96;
input n_37;
input n_189;
input n_165;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_177;
input n_60;
input n_155;
input n_152;
input n_197;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_195;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_203;
input n_205;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_179;
input n_125;
input n_35;
input n_167;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_202;
input n_130;
input n_157;
input n_29;
input n_79;
input n_193;
input n_131;
input n_151;
input n_47;
input n_173;
input n_192;
input n_25;
input n_53;
input n_160;
input n_198;
input n_188;
input n_190;
input n_8;
input n_201;
input n_158;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_159;
input n_163;
input n_95;
input n_119;
input n_183;
input n_185;
input n_175;
input n_169;
input n_59;
input n_26;
input n_133;
input n_55;
input n_196;
input n_99;
input n_2;
input n_211;
input n_181;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_178;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_200;
input n_87;
input n_150;
input n_162;
input n_27;
input n_170;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_209;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_174;
input n_186;
input n_199;
input n_134;
input n_187;
input n_32;
input n_41;
input n_104;
input n_172;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_166;
input n_11;
input n_206;
input n_171;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_204;
input n_50;
input n_52;
input n_88;
input n_110;

output n_1144;

wire n_924;
wire n_676;
wire n_294;
wire n_431;
wire n_318;
wire n_380;
wire n_419;
wire n_977;
wire n_653;
wire n_611;
wire n_444;
wire n_1126;
wire n_642;
wire n_469;
wire n_615;
wire n_851;
wire n_1060;
wire n_1141;
wire n_785;
wire n_316;
wire n_855;
wire n_389;
wire n_843;
wire n_549;
wire n_684;
wire n_850;
wire n_418;
wire n_248;
wire n_315;
wire n_523;
wire n_268;
wire n_451;
wire n_532;
wire n_705;
wire n_619;
wire n_408;
wire n_865;
wire n_913;
wire n_678;
wire n_664;
wire n_376;
wire n_697;
wire n_503;
wire n_967;
wire n_235;
wire n_226;
wire n_605;
wire n_776;
wire n_1139;
wire n_667;
wire n_515;
wire n_790;
wire n_353;
wire n_351;
wire n_367;
wire n_620;
wire n_643;
wire n_1055;
wire n_916;
wire n_452;
wire n_885;
wire n_1081;
wire n_397;
wire n_493;
wire n_525;
wire n_880;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_483;
wire n_544;
wire n_683;
wire n_1007;
wire n_780;
wire n_649;
wire n_552;
wire n_1057;
wire n_1051;
wire n_547;
wire n_1066;
wire n_1085;
wire n_721;
wire n_998;
wire n_841;
wire n_1050;
wire n_1099;
wire n_956;
wire n_564;
wire n_467;
wire n_802;
wire n_423;
wire n_840;
wire n_284;
wire n_245;
wire n_501;
wire n_823;
wire n_725;
wire n_983;
wire n_1128;
wire n_280;
wire n_744;
wire n_1021;
wire n_590;
wire n_629;
wire n_672;
wire n_873;
wire n_378;
wire n_1112;
wire n_551;
wire n_762;
wire n_581;
wire n_688;
wire n_382;
wire n_554;
wire n_800;
wire n_898;
wire n_254;
wire n_690;
wire n_1013;
wire n_583;
wire n_671;
wire n_718;
wire n_819;
wire n_302;
wire n_265;
wire n_1022;
wire n_526;
wire n_915;
wire n_1120;
wire n_719;
wire n_293;
wire n_372;
wire n_443;
wire n_244;
wire n_677;
wire n_859;
wire n_864;
wire n_1110;
wire n_951;
wire n_1121;
wire n_821;
wire n_714;
wire n_447;
wire n_247;
wire n_314;
wire n_433;
wire n_368;
wire n_604;
wire n_321;
wire n_292;
wire n_909;
wire n_625;
wire n_854;
wire n_949;
wire n_621;
wire n_753;
wire n_997;
wire n_455;
wire n_674;
wire n_1008;
wire n_932;
wire n_417;
wire n_946;
wire n_1048;
wire n_612;
wire n_1001;
wire n_212;
wire n_385;
wire n_516;
wire n_498;
wire n_933;
wire n_788;
wire n_507;
wire n_497;
wire n_689;
wire n_738;
wire n_912;
wire n_606;
wire n_559;
wire n_275;
wire n_640;
wire n_968;
wire n_252;
wire n_624;
wire n_825;
wire n_295;
wire n_1010;
wire n_330;
wire n_877;
wire n_508;
wire n_739;
wire n_506;
wire n_737;
wire n_610;
wire n_972;
wire n_692;
wire n_986;
wire n_755;
wire n_1118;
wire n_509;
wire n_568;
wire n_936;
wire n_373;
wire n_820;
wire n_757;
wire n_947;
wire n_1090;
wire n_307;
wire n_633;
wire n_439;
wire n_530;
wire n_1024;
wire n_556;
wire n_1063;
wire n_1107;
wire n_259;
wire n_448;
wire n_758;
wire n_999;
wire n_668;
wire n_733;
wire n_991;
wire n_375;
wire n_301;
wire n_828;
wire n_779;
wire n_576;
wire n_941;
wire n_929;
wire n_981;
wire n_1143;
wire n_804;
wire n_867;
wire n_1124;
wire n_537;
wire n_902;
wire n_587;
wire n_945;
wire n_1104;
wire n_659;
wire n_492;
wire n_792;
wire n_563;
wire n_756;
wire n_878;
wire n_524;
wire n_943;
wire n_399;
wire n_341;
wire n_394;
wire n_250;
wire n_579;
wire n_992;
wire n_1049;
wire n_938;
wire n_1098;
wire n_741;
wire n_548;
wire n_543;
wire n_1068;
wire n_260;
wire n_812;
wire n_842;
wire n_298;
wire n_650;
wire n_984;
wire n_320;
wire n_694;
wire n_518;
wire n_505;
wire n_286;
wire n_883;
wire n_1135;
wire n_282;
wire n_752;
wire n_331;
wire n_905;
wire n_906;
wire n_406;
wire n_519;
wire n_470;
wire n_908;
wire n_782;
wire n_919;
wire n_1108;
wire n_325;
wire n_449;
wire n_1073;
wire n_1100;
wire n_862;
wire n_900;
wire n_724;
wire n_856;
wire n_546;
wire n_1016;
wire n_760;
wire n_658;
wire n_281;
wire n_918;
wire n_240;
wire n_942;
wire n_381;
wire n_220;
wire n_291;
wire n_231;
wire n_257;
wire n_390;
wire n_731;
wire n_456;
wire n_371;
wire n_959;
wire n_1077;
wire n_481;
wire n_535;
wire n_709;
wire n_540;
wire n_317;
wire n_618;
wire n_940;
wire n_896;
wire n_323;
wire n_569;
wire n_769;
wire n_356;
wire n_227;
wire n_592;
wire n_920;
wire n_894;
wire n_1046;
wire n_271;
wire n_934;
wire n_1017;
wire n_831;
wire n_826;
wire n_335;
wire n_886;
wire n_978;
wire n_964;
wire n_1054;
wire n_654;
wire n_370;
wire n_976;
wire n_1095;
wire n_1096;
wire n_234;
wire n_343;
wire n_308;
wire n_379;
wire n_428;
wire n_267;
wire n_514;
wire n_457;
wire n_570;
wire n_833;
wire n_297;
wire n_1045;
wire n_1079;
wire n_853;
wire n_603;
wire n_225;
wire n_377;
wire n_1078;
wire n_751;
wire n_484;
wire n_775;
wire n_219;
wire n_1033;
wire n_988;
wire n_442;
wire n_814;
wire n_636;
wire n_786;
wire n_1083;
wire n_600;
wire n_1142;
wire n_660;
wire n_223;
wire n_1114;
wire n_1129;
wire n_392;
wire n_655;
wire n_704;
wire n_787;
wire n_1009;
wire n_264;
wire n_669;
wire n_472;
wire n_742;
wire n_750;
wire n_454;
wire n_961;
wire n_995;
wire n_955;
wire n_387;
wire n_771;
wire n_374;
wire n_276;
wire n_339;
wire n_882;
wire n_243;
wire n_398;
wire n_396;
wire n_1036;
wire n_635;
wire n_1097;
wire n_347;
wire n_763;
wire n_550;
wire n_522;
wire n_696;
wire n_255;
wire n_1020;
wire n_215;
wire n_350;
wire n_798;
wire n_662;
wire n_459;
wire n_897;
wire n_646;
wire n_1062;
wire n_218;
wire n_400;
wire n_930;
wire n_436;
wire n_962;
wire n_290;
wire n_580;
wire n_221;
wire n_622;
wire n_1040;
wire n_1087;
wire n_723;
wire n_1065;
wire n_1035;
wire n_386;
wire n_578;
wire n_994;
wire n_926;
wire n_287;
wire n_344;
wire n_848;
wire n_555;
wire n_783;
wire n_473;
wire n_422;
wire n_475;
wire n_777;
wire n_1070;
wire n_1030;
wire n_661;
wire n_682;
wire n_415;
wire n_485;
wire n_1043;
wire n_1071;
wire n_496;
wire n_355;
wire n_958;
wire n_849;
wire n_1034;
wire n_486;
wire n_670;
wire n_816;
wire n_336;
wire n_584;
wire n_681;
wire n_591;
wire n_922;
wire n_521;
wire n_614;
wire n_663;
wire n_845;
wire n_337;
wire n_430;
wire n_313;
wire n_631;
wire n_673;
wire n_837;
wire n_479;
wire n_528;
wire n_510;
wire n_216;
wire n_680;
wire n_974;
wire n_395;
wire n_432;
wire n_553;
wire n_727;
wire n_839;
wire n_901;
wire n_311;
wire n_813;
wire n_957;
wire n_830;
wire n_773;
wire n_743;
wire n_214;
wire n_328;
wire n_801;
wire n_299;
wire n_303;
wire n_369;
wire n_675;
wire n_888;
wire n_296;
wire n_613;
wire n_871;
wire n_1119;
wire n_241;
wire n_637;
wire n_357;
wire n_875;
wire n_598;
wire n_685;
wire n_608;
wire n_446;
wire n_445;
wire n_749;
wire n_928;
wire n_858;
wire n_829;
wire n_1064;
wire n_923;
wire n_772;
wire n_691;
wire n_1134;
wire n_881;
wire n_717;
wire n_468;
wire n_499;
wire n_939;
wire n_213;
wire n_342;
wire n_482;
wire n_517;
wire n_1088;
wire n_588;
wire n_361;
wire n_464;
wire n_789;
wire n_363;
wire n_413;
wire n_402;
wire n_734;
wire n_638;
wire n_1086;
wire n_700;
wire n_796;
wire n_573;
wire n_866;
wire n_969;
wire n_236;
wire n_1069;
wire n_1075;
wire n_1132;
wire n_388;
wire n_1127;
wire n_761;
wire n_1012;
wire n_1019;
wire n_1105;
wire n_249;
wire n_903;
wire n_1006;
wire n_740;
wire n_304;
wire n_329;
wire n_274;
wire n_577;
wire n_384;
wire n_582;
wire n_460;
wire n_889;
wire n_973;
wire n_277;
wire n_1061;
wire n_477;
wire n_338;
wire n_571;
wire n_461;
wire n_333;
wire n_693;
wire n_309;
wire n_512;
wire n_836;
wire n_990;
wire n_462;
wire n_975;
wire n_322;
wire n_567;
wire n_258;
wire n_1113;
wire n_652;
wire n_778;
wire n_1111;
wire n_1122;
wire n_306;
wire n_907;
wire n_722;
wire n_1093;
wire n_458;
wire n_288;
wire n_770;
wire n_844;
wire n_1031;
wire n_263;
wire n_471;
wire n_609;
wire n_852;
wire n_989;
wire n_1041;
wire n_1039;
wire n_1102;
wire n_224;
wire n_228;
wire n_283;
wire n_1028;
wire n_383;
wire n_711;
wire n_781;
wire n_834;
wire n_474;
wire n_765;
wire n_542;
wire n_463;
wire n_488;
wire n_595;
wire n_736;
wire n_502;
wire n_893;
wire n_892;
wire n_1015;
wire n_1000;
wire n_891;
wire n_1140;
wire n_239;
wire n_466;
wire n_420;
wire n_630;
wire n_489;
wire n_632;
wire n_699;
wire n_979;
wire n_1002;
wire n_617;
wire n_310;
wire n_593;
wire n_504;
wire n_511;
wire n_846;
wire n_586;
wire n_748;
wire n_1058;
wire n_465;
wire n_838;
wire n_358;
wire n_874;
wire n_362;
wire n_876;
wire n_332;
wire n_1053;
wire n_1101;
wire n_273;
wire n_585;
wire n_349;
wire n_1106;
wire n_270;
wire n_616;
wire n_230;
wire n_953;
wire n_601;
wire n_279;
wire n_917;
wire n_1014;
wire n_966;
wire n_987;
wire n_253;
wire n_261;
wire n_289;
wire n_963;
wire n_745;
wire n_1052;
wire n_954;
wire n_627;
wire n_1116;
wire n_767;
wire n_993;
wire n_217;
wire n_440;
wire n_726;
wire n_478;
wire n_793;
wire n_545;
wire n_982;
wire n_441;
wire n_860;
wire n_1103;
wire n_450;
wire n_648;
wire n_312;
wire n_476;
wire n_818;
wire n_429;
wire n_861;
wire n_534;
wire n_948;
wire n_1076;
wire n_884;
wire n_899;
wire n_345;
wire n_944;
wire n_1091;
wire n_494;
wire n_641;
wire n_628;
wire n_365;
wire n_774;
wire n_729;
wire n_730;
wire n_1059;
wire n_1084;
wire n_1131;
wire n_1133;
wire n_970;
wire n_911;
wire n_557;
wire n_1005;
wire n_354;
wire n_607;
wire n_575;
wire n_480;
wire n_679;
wire n_237;
wire n_425;
wire n_513;
wire n_407;
wire n_527;
wire n_647;
wire n_707;
wire n_710;
wire n_795;
wire n_695;
wire n_832;
wire n_857;
wire n_1072;
wire n_560;
wire n_656;
wire n_340;
wire n_1094;
wire n_561;
wire n_1044;
wire n_346;
wire n_937;
wire n_393;
wire n_229;
wire n_495;
wire n_487;
wire n_602;
wire n_665;
wire n_574;
wire n_437;
wire n_453;
wire n_403;
wire n_421;
wire n_879;
wire n_1130;
wire n_720;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_863;
wire n_910;
wire n_971;
wire n_490;
wire n_805;
wire n_1027;
wire n_326;
wire n_794;
wire n_768;
wire n_921;
wire n_996;
wire n_233;
wire n_404;
wire n_686;
wire n_366;
wire n_572;
wire n_712;
wire n_754;
wire n_847;
wire n_1136;
wire n_815;
wire n_246;
wire n_596;
wire n_1125;
wire n_410;
wire n_1042;
wire n_558;
wire n_708;
wire n_269;
wire n_529;
wire n_735;
wire n_702;
wire n_285;
wire n_822;
wire n_412;
wire n_232;
wire n_327;
wire n_1109;
wire n_657;
wire n_644;
wire n_728;
wire n_895;
wire n_1037;
wire n_1080;
wire n_266;
wire n_272;
wire n_491;
wire n_1074;
wire n_427;
wire n_791;
wire n_732;
wire n_251;
wire n_352;
wire n_566;
wire n_565;
wire n_426;
wire n_520;
wire n_808;
wire n_409;
wire n_797;
wire n_1038;
wire n_1025;
wire n_1082;
wire n_887;
wire n_589;
wire n_716;
wire n_597;
wire n_500;
wire n_562;
wire n_1067;
wire n_300;
wire n_651;
wire n_435;
wire n_809;
wire n_870;
wire n_931;
wire n_334;
wire n_599;
wire n_811;
wire n_766;
wire n_952;
wire n_541;
wire n_807;
wire n_391;
wire n_701;
wire n_434;
wire n_1023;
wire n_645;
wire n_539;
wire n_835;
wire n_538;
wire n_666;
wire n_262;
wire n_803;
wire n_868;
wire n_1092;
wire n_238;
wire n_1117;
wire n_639;
wire n_799;
wire n_914;
wire n_687;
wire n_715;
wire n_411;
wire n_414;
wire n_1026;
wire n_319;
wire n_364;
wire n_965;
wire n_927;
wire n_1089;
wire n_872;
wire n_1138;
wire n_536;
wire n_531;
wire n_935;
wire n_1004;
wire n_242;
wire n_817;
wire n_1032;
wire n_360;
wire n_594;
wire n_764;
wire n_890;
wire n_1056;
wire n_960;
wire n_759;
wire n_1018;
wire n_222;
wire n_438;
wire n_806;
wire n_713;
wire n_1011;
wire n_1123;
wire n_904;
wire n_985;
wire n_1047;
wire n_869;
wire n_324;
wire n_810;
wire n_634;
wire n_416;
wire n_827;
wire n_401;
wire n_348;
wire n_1029;
wire n_626;
wire n_925;
wire n_424;
wire n_1003;
wire n_1137;
wire n_706;
wire n_746;
wire n_256;
wire n_305;
wire n_533;
wire n_950;
wire n_747;
wire n_278;
wire n_784;

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_198),
.Y(n_212)
);

BUFx6f_ASAP7_75t_L g213 ( 
.A(n_50),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_91),
.Y(n_214)
);

CKINVDCx14_ASAP7_75t_R g215 ( 
.A(n_201),
.Y(n_215)
);

INVxp33_ASAP7_75t_R g216 ( 
.A(n_87),
.Y(n_216)
);

INVx2_ASAP7_75t_SL g217 ( 
.A(n_120),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_147),
.Y(n_218)
);

BUFx2_ASAP7_75t_SL g219 ( 
.A(n_161),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_72),
.Y(n_220)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_159),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_158),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_76),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_165),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_81),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_24),
.Y(n_226)
);

BUFx10_ASAP7_75t_L g227 ( 
.A(n_42),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_171),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_144),
.Y(n_229)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_188),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_69),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_75),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_105),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_199),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_189),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_149),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_90),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_155),
.Y(n_238)
);

INVx1_ASAP7_75t_SL g239 ( 
.A(n_39),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_179),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_169),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_127),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_62),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_181),
.Y(n_244)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_160),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_92),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_204),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_38),
.Y(n_248)
);

BUFx3_ASAP7_75t_L g249 ( 
.A(n_167),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_118),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_98),
.Y(n_251)
);

BUFx6f_ASAP7_75t_L g252 ( 
.A(n_141),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_103),
.Y(n_253)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_186),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_84),
.Y(n_255)
);

BUFx3_ASAP7_75t_L g256 ( 
.A(n_196),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_88),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_9),
.Y(n_258)
);

INVxp33_ASAP7_75t_SL g259 ( 
.A(n_83),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_93),
.Y(n_260)
);

INVx2_ASAP7_75t_SL g261 ( 
.A(n_150),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_166),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_173),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_102),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_9),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_78),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_157),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_136),
.Y(n_268)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_14),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_205),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_46),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_11),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_128),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_200),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_126),
.Y(n_275)
);

BUFx8_ASAP7_75t_SL g276 ( 
.A(n_99),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_203),
.Y(n_277)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_184),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_197),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_131),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_193),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_209),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_1),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_258),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_265),
.Y(n_285)
);

BUFx6f_ASAP7_75t_L g286 ( 
.A(n_213),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_226),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_249),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_272),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_249),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_283),
.Y(n_291)
);

INVxp67_ASAP7_75t_SL g292 ( 
.A(n_256),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_256),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_229),
.Y(n_294)
);

BUFx6f_ASAP7_75t_L g295 ( 
.A(n_213),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_235),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_236),
.Y(n_297)
);

INVxp67_ASAP7_75t_SL g298 ( 
.A(n_238),
.Y(n_298)
);

HB1xp67_ASAP7_75t_L g299 ( 
.A(n_269),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_276),
.Y(n_300)
);

NAND2xp33_ASAP7_75t_R g301 ( 
.A(n_212),
.B(n_0),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_240),
.Y(n_302)
);

CKINVDCx16_ASAP7_75t_R g303 ( 
.A(n_215),
.Y(n_303)
);

INVxp67_ASAP7_75t_SL g304 ( 
.A(n_247),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_260),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_214),
.Y(n_306)
);

INVxp67_ASAP7_75t_SL g307 ( 
.A(n_266),
.Y(n_307)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_269),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_273),
.Y(n_309)
);

INVx2_ASAP7_75t_L g310 ( 
.A(n_213),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_275),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_276),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_279),
.Y(n_313)
);

INVxp33_ASAP7_75t_SL g314 ( 
.A(n_219),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_221),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_267),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_221),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_230),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_267),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_230),
.Y(n_320)
);

CKINVDCx16_ASAP7_75t_R g321 ( 
.A(n_215),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_228),
.Y(n_322)
);

INVxp67_ASAP7_75t_SL g323 ( 
.A(n_245),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_218),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_245),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_220),
.Y(n_326)
);

INVxp33_ASAP7_75t_SL g327 ( 
.A(n_222),
.Y(n_327)
);

CKINVDCx16_ASAP7_75t_R g328 ( 
.A(n_234),
.Y(n_328)
);

INVxp67_ASAP7_75t_SL g329 ( 
.A(n_254),
.Y(n_329)
);

INVxp33_ASAP7_75t_SL g330 ( 
.A(n_223),
.Y(n_330)
);

INVxp67_ASAP7_75t_L g331 ( 
.A(n_227),
.Y(n_331)
);

INVxp67_ASAP7_75t_SL g332 ( 
.A(n_254),
.Y(n_332)
);

INVx2_ASAP7_75t_L g333 ( 
.A(n_310),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_299),
.Y(n_334)
);

BUFx6f_ASAP7_75t_L g335 ( 
.A(n_286),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_294),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_296),
.Y(n_337)
);

BUFx2_ASAP7_75t_L g338 ( 
.A(n_300),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_297),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_302),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_305),
.Y(n_341)
);

INVx2_ASAP7_75t_L g342 ( 
.A(n_310),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_309),
.Y(n_343)
);

BUFx6f_ASAP7_75t_L g344 ( 
.A(n_286),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_306),
.B(n_217),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_311),
.Y(n_346)
);

BUFx6f_ASAP7_75t_L g347 ( 
.A(n_286),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_324),
.B(n_261),
.Y(n_348)
);

AND2x2_ASAP7_75t_L g349 ( 
.A(n_292),
.B(n_227),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_313),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_287),
.Y(n_351)
);

BUFx2_ASAP7_75t_L g352 ( 
.A(n_284),
.Y(n_352)
);

HB1xp67_ASAP7_75t_L g353 ( 
.A(n_284),
.Y(n_353)
);

AND2x4_ASAP7_75t_L g354 ( 
.A(n_298),
.B(n_278),
.Y(n_354)
);

AND2x4_ASAP7_75t_L g355 ( 
.A(n_304),
.B(n_278),
.Y(n_355)
);

NOR2x1_ASAP7_75t_L g356 ( 
.A(n_315),
.B(n_317),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_318),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_320),
.Y(n_358)
);

BUFx6f_ASAP7_75t_L g359 ( 
.A(n_286),
.Y(n_359)
);

INVx2_ASAP7_75t_L g360 ( 
.A(n_295),
.Y(n_360)
);

NOR2x1_ASAP7_75t_L g361 ( 
.A(n_325),
.B(n_239),
.Y(n_361)
);

INVx2_ASAP7_75t_L g362 ( 
.A(n_295),
.Y(n_362)
);

INVx4_ASAP7_75t_L g363 ( 
.A(n_295),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_300),
.Y(n_364)
);

INVx5_ASAP7_75t_L g365 ( 
.A(n_295),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_288),
.Y(n_366)
);

INVx3_ASAP7_75t_L g367 ( 
.A(n_308),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_312),
.Y(n_368)
);

INVx2_ASAP7_75t_L g369 ( 
.A(n_308),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_312),
.Y(n_370)
);

AND2x4_ASAP7_75t_L g371 ( 
.A(n_307),
.B(n_213),
.Y(n_371)
);

BUFx6f_ASAP7_75t_L g372 ( 
.A(n_290),
.Y(n_372)
);

INVx6_ASAP7_75t_L g373 ( 
.A(n_303),
.Y(n_373)
);

AND2x4_ASAP7_75t_L g374 ( 
.A(n_323),
.B(n_252),
.Y(n_374)
);

OAI22xp5_ASAP7_75t_SL g375 ( 
.A1(n_316),
.A2(n_282),
.B1(n_243),
.B2(n_259),
.Y(n_375)
);

BUFx6f_ASAP7_75t_L g376 ( 
.A(n_293),
.Y(n_376)
);

INVx2_ASAP7_75t_L g377 ( 
.A(n_329),
.Y(n_377)
);

AND2x6_ASAP7_75t_L g378 ( 
.A(n_321),
.B(n_252),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_332),
.Y(n_379)
);

INVx2_ASAP7_75t_L g380 ( 
.A(n_326),
.Y(n_380)
);

INVx2_ASAP7_75t_L g381 ( 
.A(n_285),
.Y(n_381)
);

OAI22xp5_ASAP7_75t_L g382 ( 
.A1(n_331),
.A2(n_281),
.B1(n_280),
.B2(n_277),
.Y(n_382)
);

INVx2_ASAP7_75t_L g383 ( 
.A(n_285),
.Y(n_383)
);

BUFx2_ASAP7_75t_L g384 ( 
.A(n_289),
.Y(n_384)
);

BUFx6f_ASAP7_75t_L g385 ( 
.A(n_289),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_314),
.B(n_327),
.Y(n_386)
);

BUFx6f_ASAP7_75t_L g387 ( 
.A(n_291),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_357),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_358),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_333),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_351),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_SL g392 ( 
.A(n_385),
.B(n_314),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_SL g393 ( 
.A(n_385),
.B(n_327),
.Y(n_393)
);

BUFx6f_ASAP7_75t_L g394 ( 
.A(n_335),
.Y(n_394)
);

OR2x6_ASAP7_75t_L g395 ( 
.A(n_380),
.B(n_216),
.Y(n_395)
);

AND2x2_ASAP7_75t_L g396 ( 
.A(n_354),
.B(n_291),
.Y(n_396)
);

INVx2_ASAP7_75t_SL g397 ( 
.A(n_349),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_333),
.Y(n_398)
);

NOR2x1p5_ASAP7_75t_L g399 ( 
.A(n_386),
.B(n_316),
.Y(n_399)
);

INVxp33_ASAP7_75t_L g400 ( 
.A(n_334),
.Y(n_400)
);

INVx2_ASAP7_75t_L g401 ( 
.A(n_342),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_342),
.Y(n_402)
);

HB1xp67_ASAP7_75t_L g403 ( 
.A(n_349),
.Y(n_403)
);

INVx2_ASAP7_75t_L g404 ( 
.A(n_369),
.Y(n_404)
);

INVx2_ASAP7_75t_L g405 ( 
.A(n_369),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_372),
.Y(n_406)
);

AND2x2_ASAP7_75t_L g407 ( 
.A(n_354),
.B(n_355),
.Y(n_407)
);

OR2x2_ASAP7_75t_L g408 ( 
.A(n_377),
.B(n_328),
.Y(n_408)
);

AND3x2_ASAP7_75t_L g409 ( 
.A(n_338),
.B(n_227),
.C(n_301),
.Y(n_409)
);

BUFx6f_ASAP7_75t_L g410 ( 
.A(n_335),
.Y(n_410)
);

HB1xp67_ASAP7_75t_L g411 ( 
.A(n_377),
.Y(n_411)
);

INVx3_ASAP7_75t_L g412 ( 
.A(n_335),
.Y(n_412)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_360),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_SL g414 ( 
.A(n_385),
.B(n_330),
.Y(n_414)
);

NOR2x1p5_ASAP7_75t_L g415 ( 
.A(n_380),
.B(n_319),
.Y(n_415)
);

INVx5_ASAP7_75t_L g416 ( 
.A(n_335),
.Y(n_416)
);

INVx3_ASAP7_75t_L g417 ( 
.A(n_344),
.Y(n_417)
);

INVx8_ASAP7_75t_L g418 ( 
.A(n_378),
.Y(n_418)
);

AND2x2_ASAP7_75t_L g419 ( 
.A(n_354),
.B(n_224),
.Y(n_419)
);

NOR2xp33_ASAP7_75t_L g420 ( 
.A(n_345),
.B(n_330),
.Y(n_420)
);

INVxp33_ASAP7_75t_L g421 ( 
.A(n_353),
.Y(n_421)
);

OR2x2_ASAP7_75t_L g422 ( 
.A(n_379),
.B(n_319),
.Y(n_422)
);

OAI22xp33_ASAP7_75t_L g423 ( 
.A1(n_381),
.A2(n_251),
.B1(n_274),
.B2(n_271),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_SL g424 ( 
.A(n_385),
.B(n_225),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_374),
.B(n_231),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_372),
.Y(n_426)
);

INVxp67_ASAP7_75t_SL g427 ( 
.A(n_344),
.Y(n_427)
);

INVx3_ASAP7_75t_L g428 ( 
.A(n_344),
.Y(n_428)
);

OR2x2_ASAP7_75t_L g429 ( 
.A(n_371),
.B(n_232),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_374),
.B(n_233),
.Y(n_430)
);

INVx2_ASAP7_75t_SL g431 ( 
.A(n_373),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_372),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_336),
.Y(n_433)
);

INVxp67_ASAP7_75t_SL g434 ( 
.A(n_344),
.Y(n_434)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_360),
.Y(n_435)
);

NOR2xp33_ASAP7_75t_L g436 ( 
.A(n_348),
.B(n_322),
.Y(n_436)
);

INVx2_ASAP7_75t_L g437 ( 
.A(n_362),
.Y(n_437)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_362),
.Y(n_438)
);

INVx2_ASAP7_75t_L g439 ( 
.A(n_347),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_337),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_339),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_340),
.Y(n_442)
);

INVx1_ASAP7_75t_SL g443 ( 
.A(n_352),
.Y(n_443)
);

INVx2_ASAP7_75t_L g444 ( 
.A(n_347),
.Y(n_444)
);

INVxp33_ASAP7_75t_SL g445 ( 
.A(n_375),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_341),
.Y(n_446)
);

INVx2_ASAP7_75t_L g447 ( 
.A(n_347),
.Y(n_447)
);

AND2x2_ASAP7_75t_L g448 ( 
.A(n_355),
.B(n_237),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_374),
.B(n_241),
.Y(n_449)
);

INVx1_ASAP7_75t_SL g450 ( 
.A(n_352),
.Y(n_450)
);

OR2x6_ASAP7_75t_L g451 ( 
.A(n_381),
.B(n_383),
.Y(n_451)
);

AND2x2_ASAP7_75t_L g452 ( 
.A(n_355),
.B(n_242),
.Y(n_452)
);

INVx2_ASAP7_75t_L g453 ( 
.A(n_347),
.Y(n_453)
);

NAND2xp33_ASAP7_75t_L g454 ( 
.A(n_378),
.B(n_252),
.Y(n_454)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_359),
.Y(n_455)
);

INVx2_ASAP7_75t_L g456 ( 
.A(n_359),
.Y(n_456)
);

INVx3_ASAP7_75t_L g457 ( 
.A(n_359),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_371),
.B(n_244),
.Y(n_458)
);

INVx2_ASAP7_75t_L g459 ( 
.A(n_359),
.Y(n_459)
);

INVx2_ASAP7_75t_L g460 ( 
.A(n_367),
.Y(n_460)
);

BUFx10_ASAP7_75t_L g461 ( 
.A(n_373),
.Y(n_461)
);

HB1xp67_ASAP7_75t_L g462 ( 
.A(n_382),
.Y(n_462)
);

INVx2_ASAP7_75t_SL g463 ( 
.A(n_373),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_411),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_388),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_388),
.Y(n_466)
);

INVxp67_ASAP7_75t_L g467 ( 
.A(n_408),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_389),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_389),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_391),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_433),
.Y(n_471)
);

BUFx6f_ASAP7_75t_L g472 ( 
.A(n_394),
.Y(n_472)
);

INVx2_ASAP7_75t_SL g473 ( 
.A(n_408),
.Y(n_473)
);

AND2x2_ASAP7_75t_L g474 ( 
.A(n_397),
.B(n_387),
.Y(n_474)
);

NOR2xp33_ASAP7_75t_L g475 ( 
.A(n_420),
.B(n_383),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_440),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_441),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_442),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_446),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_407),
.Y(n_480)
);

NOR2xp33_ASAP7_75t_L g481 ( 
.A(n_400),
.B(n_387),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_407),
.Y(n_482)
);

BUFx6f_ASAP7_75t_L g483 ( 
.A(n_394),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_404),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_404),
.Y(n_485)
);

BUFx6f_ASAP7_75t_L g486 ( 
.A(n_394),
.Y(n_486)
);

CKINVDCx16_ASAP7_75t_R g487 ( 
.A(n_461),
.Y(n_487)
);

NAND2xp33_ASAP7_75t_R g488 ( 
.A(n_445),
.B(n_384),
.Y(n_488)
);

AND2x4_ASAP7_75t_L g489 ( 
.A(n_451),
.B(n_366),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_405),
.Y(n_490)
);

NOR2xp33_ASAP7_75t_L g491 ( 
.A(n_397),
.B(n_387),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_413),
.Y(n_492)
);

NOR2xp67_ASAP7_75t_L g493 ( 
.A(n_406),
.B(n_363),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_413),
.Y(n_494)
);

INVx2_ASAP7_75t_SL g495 ( 
.A(n_396),
.Y(n_495)
);

NOR2xp33_ASAP7_75t_L g496 ( 
.A(n_392),
.B(n_387),
.Y(n_496)
);

CKINVDCx5p33_ASAP7_75t_R g497 ( 
.A(n_461),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_435),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_403),
.B(n_371),
.Y(n_499)
);

NOR2xp33_ASAP7_75t_L g500 ( 
.A(n_422),
.B(n_364),
.Y(n_500)
);

AND2x2_ASAP7_75t_L g501 ( 
.A(n_396),
.B(n_361),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_435),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_419),
.B(n_378),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_437),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_437),
.Y(n_505)
);

NAND2x1p5_ASAP7_75t_L g506 ( 
.A(n_431),
.B(n_252),
.Y(n_506)
);

AND2x2_ASAP7_75t_L g507 ( 
.A(n_443),
.B(n_364),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_438),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_438),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_460),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_460),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_390),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_390),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_398),
.Y(n_514)
);

NOR2xp33_ASAP7_75t_SL g515 ( 
.A(n_445),
.B(n_368),
.Y(n_515)
);

INVx2_ASAP7_75t_SL g516 ( 
.A(n_429),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_398),
.Y(n_517)
);

XOR2x2_ASAP7_75t_L g518 ( 
.A(n_436),
.B(n_322),
.Y(n_518)
);

AND2x2_ASAP7_75t_L g519 ( 
.A(n_450),
.B(n_368),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_419),
.B(n_378),
.Y(n_520)
);

NAND2x1p5_ASAP7_75t_L g521 ( 
.A(n_431),
.B(n_343),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_402),
.Y(n_522)
);

OR2x2_ASAP7_75t_L g523 ( 
.A(n_422),
.B(n_370),
.Y(n_523)
);

CKINVDCx5p33_ASAP7_75t_R g524 ( 
.A(n_461),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_402),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_401),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_401),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_451),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_451),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_448),
.B(n_378),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_451),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_448),
.Y(n_532)
);

NOR2xp33_ASAP7_75t_L g533 ( 
.A(n_462),
.B(n_370),
.Y(n_533)
);

INVxp67_ASAP7_75t_L g534 ( 
.A(n_395),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_452),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_452),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_429),
.Y(n_537)
);

CKINVDCx16_ASAP7_75t_R g538 ( 
.A(n_395),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_406),
.Y(n_539)
);

INVx2_ASAP7_75t_L g540 ( 
.A(n_412),
.Y(n_540)
);

AND2x2_ASAP7_75t_SL g541 ( 
.A(n_454),
.B(n_346),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_426),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_426),
.Y(n_543)
);

CKINVDCx5p33_ASAP7_75t_R g544 ( 
.A(n_463),
.Y(n_544)
);

NOR2xp33_ASAP7_75t_L g545 ( 
.A(n_421),
.B(n_350),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_432),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_432),
.Y(n_547)
);

CKINVDCx16_ASAP7_75t_R g548 ( 
.A(n_395),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_L g549 ( 
.A(n_475),
.B(n_458),
.Y(n_549)
);

INVx2_ASAP7_75t_SL g550 ( 
.A(n_473),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_480),
.B(n_425),
.Y(n_551)
);

INVx2_ASAP7_75t_L g552 ( 
.A(n_484),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_L g553 ( 
.A(n_482),
.B(n_430),
.Y(n_553)
);

INVx2_ASAP7_75t_SL g554 ( 
.A(n_507),
.Y(n_554)
);

O2A1O1Ixp33_ASAP7_75t_L g555 ( 
.A1(n_499),
.A2(n_423),
.B(n_414),
.C(n_393),
.Y(n_555)
);

NOR2x1p5_ASAP7_75t_L g556 ( 
.A(n_497),
.B(n_395),
.Y(n_556)
);

AOI22xp33_ASAP7_75t_L g557 ( 
.A1(n_532),
.A2(n_378),
.B1(n_449),
.B2(n_399),
.Y(n_557)
);

O2A1O1Ixp33_ASAP7_75t_L g558 ( 
.A1(n_499),
.A2(n_424),
.B(n_454),
.C(n_415),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_512),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_L g560 ( 
.A(n_491),
.B(n_412),
.Y(n_560)
);

BUFx3_ASAP7_75t_L g561 ( 
.A(n_544),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_L g562 ( 
.A(n_465),
.B(n_466),
.Y(n_562)
);

OR2x6_ASAP7_75t_L g563 ( 
.A(n_534),
.B(n_463),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_L g564 ( 
.A(n_468),
.B(n_412),
.Y(n_564)
);

BUFx6f_ASAP7_75t_L g565 ( 
.A(n_472),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_L g566 ( 
.A(n_469),
.B(n_474),
.Y(n_566)
);

INVx2_ASAP7_75t_SL g567 ( 
.A(n_519),
.Y(n_567)
);

INVx2_ASAP7_75t_L g568 ( 
.A(n_485),
.Y(n_568)
);

AOI22xp33_ASAP7_75t_L g569 ( 
.A1(n_535),
.A2(n_418),
.B1(n_376),
.B2(n_372),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_SL g570 ( 
.A(n_481),
.B(n_496),
.Y(n_570)
);

NOR2xp33_ASAP7_75t_L g571 ( 
.A(n_500),
.B(n_409),
.Y(n_571)
);

INVx3_ASAP7_75t_L g572 ( 
.A(n_472),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_SL g573 ( 
.A(n_495),
.B(n_418),
.Y(n_573)
);

INVxp67_ASAP7_75t_L g574 ( 
.A(n_545),
.Y(n_574)
);

AOI22xp5_ASAP7_75t_L g575 ( 
.A1(n_501),
.A2(n_418),
.B1(n_427),
.B2(n_434),
.Y(n_575)
);

NOR2x2_ASAP7_75t_L g576 ( 
.A(n_518),
.B(n_439),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_L g577 ( 
.A(n_536),
.B(n_459),
.Y(n_577)
);

CKINVDCx5p33_ASAP7_75t_R g578 ( 
.A(n_487),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_L g579 ( 
.A(n_537),
.B(n_417),
.Y(n_579)
);

INVx2_ASAP7_75t_SL g580 ( 
.A(n_464),
.Y(n_580)
);

BUFx8_ASAP7_75t_L g581 ( 
.A(n_523),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_L g582 ( 
.A(n_470),
.B(n_417),
.Y(n_582)
);

INVxp67_ASAP7_75t_L g583 ( 
.A(n_467),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_513),
.Y(n_584)
);

BUFx5_ASAP7_75t_L g585 ( 
.A(n_510),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_L g586 ( 
.A(n_471),
.B(n_417),
.Y(n_586)
);

NOR2xp33_ASAP7_75t_L g587 ( 
.A(n_533),
.B(n_376),
.Y(n_587)
);

INVx3_ASAP7_75t_L g588 ( 
.A(n_472),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_L g589 ( 
.A(n_476),
.B(n_428),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_L g590 ( 
.A(n_477),
.B(n_428),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_L g591 ( 
.A(n_478),
.B(n_428),
.Y(n_591)
);

AOI22xp5_ASAP7_75t_L g592 ( 
.A1(n_516),
.A2(n_418),
.B1(n_459),
.B2(n_456),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_L g593 ( 
.A(n_479),
.B(n_457),
.Y(n_593)
);

AOI22xp33_ASAP7_75t_L g594 ( 
.A1(n_503),
.A2(n_376),
.B1(n_456),
.B2(n_455),
.Y(n_594)
);

INVx2_ASAP7_75t_SL g595 ( 
.A(n_489),
.Y(n_595)
);

AOI22xp33_ASAP7_75t_L g596 ( 
.A1(n_503),
.A2(n_376),
.B1(n_455),
.B2(n_453),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_SL g597 ( 
.A(n_489),
.B(n_394),
.Y(n_597)
);

NOR2xp33_ASAP7_75t_L g598 ( 
.A(n_528),
.B(n_457),
.Y(n_598)
);

INVxp67_ASAP7_75t_SL g599 ( 
.A(n_483),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_L g600 ( 
.A(n_514),
.B(n_439),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_517),
.Y(n_601)
);

AOI22xp33_ASAP7_75t_L g602 ( 
.A1(n_520),
.A2(n_453),
.B1(n_447),
.B2(n_444),
.Y(n_602)
);

INVx2_ASAP7_75t_L g603 ( 
.A(n_490),
.Y(n_603)
);

AOI22xp33_ASAP7_75t_L g604 ( 
.A1(n_520),
.A2(n_447),
.B1(n_444),
.B2(n_457),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_L g605 ( 
.A(n_522),
.B(n_394),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_SL g606 ( 
.A(n_529),
.B(n_410),
.Y(n_606)
);

NAND2x1_ASAP7_75t_L g607 ( 
.A(n_483),
.B(n_410),
.Y(n_607)
);

INVx2_ASAP7_75t_L g608 ( 
.A(n_526),
.Y(n_608)
);

CKINVDCx20_ASAP7_75t_R g609 ( 
.A(n_524),
.Y(n_609)
);

AOI21x1_ASAP7_75t_L g610 ( 
.A1(n_493),
.A2(n_356),
.B(n_410),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_L g611 ( 
.A(n_525),
.B(n_410),
.Y(n_611)
);

AO22x1_ASAP7_75t_L g612 ( 
.A1(n_531),
.A2(n_246),
.B1(n_248),
.B2(n_250),
.Y(n_612)
);

NAND2xp33_ASAP7_75t_L g613 ( 
.A(n_530),
.B(n_410),
.Y(n_613)
);

BUFx3_ASAP7_75t_L g614 ( 
.A(n_521),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_L g615 ( 
.A(n_530),
.B(n_367),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_SL g616 ( 
.A(n_521),
.B(n_253),
.Y(n_616)
);

AOI22xp33_ASAP7_75t_L g617 ( 
.A1(n_527),
.A2(n_511),
.B1(n_547),
.B2(n_546),
.Y(n_617)
);

OR2x2_ASAP7_75t_L g618 ( 
.A(n_574),
.B(n_538),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_L g619 ( 
.A(n_549),
.B(n_539),
.Y(n_619)
);

INVx2_ASAP7_75t_L g620 ( 
.A(n_552),
.Y(n_620)
);

BUFx4f_ASAP7_75t_L g621 ( 
.A(n_563),
.Y(n_621)
);

NOR2xp33_ASAP7_75t_L g622 ( 
.A(n_583),
.B(n_515),
.Y(n_622)
);

INVx3_ASAP7_75t_L g623 ( 
.A(n_565),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_L g624 ( 
.A(n_549),
.B(n_542),
.Y(n_624)
);

AND2x4_ASAP7_75t_L g625 ( 
.A(n_595),
.B(n_543),
.Y(n_625)
);

BUFx12f_ASAP7_75t_L g626 ( 
.A(n_578),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_559),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_L g628 ( 
.A(n_566),
.B(n_492),
.Y(n_628)
);

INVx4_ASAP7_75t_L g629 ( 
.A(n_565),
.Y(n_629)
);

BUFx4_ASAP7_75t_SL g630 ( 
.A(n_609),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_584),
.Y(n_631)
);

AOI21xp5_ASAP7_75t_L g632 ( 
.A1(n_613),
.A2(n_486),
.B(n_483),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_L g633 ( 
.A(n_551),
.B(n_494),
.Y(n_633)
);

AND2x2_ASAP7_75t_L g634 ( 
.A(n_554),
.B(n_515),
.Y(n_634)
);

HB1xp67_ASAP7_75t_L g635 ( 
.A(n_550),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_601),
.Y(n_636)
);

AND2x4_ASAP7_75t_L g637 ( 
.A(n_614),
.B(n_540),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_L g638 ( 
.A(n_570),
.B(n_541),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_600),
.Y(n_639)
);

BUFx3_ASAP7_75t_L g640 ( 
.A(n_561),
.Y(n_640)
);

BUFx6f_ASAP7_75t_L g641 ( 
.A(n_565),
.Y(n_641)
);

NAND2x1_ASAP7_75t_L g642 ( 
.A(n_572),
.B(n_486),
.Y(n_642)
);

OR2x6_ASAP7_75t_L g643 ( 
.A(n_567),
.B(n_506),
.Y(n_643)
);

INVx2_ASAP7_75t_L g644 ( 
.A(n_568),
.Y(n_644)
);

INVx3_ASAP7_75t_L g645 ( 
.A(n_572),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_L g646 ( 
.A(n_551),
.B(n_498),
.Y(n_646)
);

INVx3_ASAP7_75t_L g647 ( 
.A(n_588),
.Y(n_647)
);

INVxp33_ASAP7_75t_L g648 ( 
.A(n_571),
.Y(n_648)
);

BUFx2_ASAP7_75t_L g649 ( 
.A(n_576),
.Y(n_649)
);

OR2x2_ASAP7_75t_SL g650 ( 
.A(n_553),
.B(n_548),
.Y(n_650)
);

INVx2_ASAP7_75t_L g651 ( 
.A(n_603),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_553),
.B(n_502),
.Y(n_652)
);

HB1xp67_ASAP7_75t_L g653 ( 
.A(n_580),
.Y(n_653)
);

INVx4_ASAP7_75t_L g654 ( 
.A(n_588),
.Y(n_654)
);

INVx2_ASAP7_75t_L g655 ( 
.A(n_608),
.Y(n_655)
);

INVx4_ASAP7_75t_L g656 ( 
.A(n_563),
.Y(n_656)
);

BUFx6f_ASAP7_75t_L g657 ( 
.A(n_563),
.Y(n_657)
);

HB1xp67_ASAP7_75t_L g658 ( 
.A(n_579),
.Y(n_658)
);

O2A1O1Ixp33_ASAP7_75t_L g659 ( 
.A1(n_555),
.A2(n_506),
.B(n_508),
.C(n_509),
.Y(n_659)
);

BUFx2_ASAP7_75t_L g660 ( 
.A(n_581),
.Y(n_660)
);

INVxp67_ASAP7_75t_L g661 ( 
.A(n_581),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_600),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_L g663 ( 
.A(n_562),
.B(n_504),
.Y(n_663)
);

AOI211xp5_ASAP7_75t_L g664 ( 
.A1(n_612),
.A2(n_488),
.B(n_255),
.C(n_268),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_L g665 ( 
.A(n_587),
.B(n_505),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_L g666 ( 
.A(n_577),
.B(n_493),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_577),
.Y(n_667)
);

BUFx2_ASAP7_75t_L g668 ( 
.A(n_556),
.Y(n_668)
);

AND2x2_ASAP7_75t_L g669 ( 
.A(n_557),
.B(n_367),
.Y(n_669)
);

NOR3xp33_ASAP7_75t_SL g670 ( 
.A(n_616),
.B(n_262),
.C(n_257),
.Y(n_670)
);

CKINVDCx20_ASAP7_75t_R g671 ( 
.A(n_597),
.Y(n_671)
);

INVx5_ASAP7_75t_L g672 ( 
.A(n_599),
.Y(n_672)
);

AND2x4_ASAP7_75t_L g673 ( 
.A(n_582),
.B(n_486),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_564),
.Y(n_674)
);

NOR3xp33_ASAP7_75t_SL g675 ( 
.A(n_606),
.B(n_264),
.C(n_263),
.Y(n_675)
);

AOI22xp5_ASAP7_75t_L g676 ( 
.A1(n_586),
.A2(n_270),
.B1(n_363),
.B2(n_416),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_589),
.Y(n_677)
);

BUFx2_ASAP7_75t_L g678 ( 
.A(n_590),
.Y(n_678)
);

HB1xp67_ASAP7_75t_L g679 ( 
.A(n_591),
.Y(n_679)
);

AND2x4_ASAP7_75t_L g680 ( 
.A(n_593),
.B(n_32),
.Y(n_680)
);

BUFx6f_ASAP7_75t_L g681 ( 
.A(n_607),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_L g682 ( 
.A(n_615),
.B(n_363),
.Y(n_682)
);

INVx5_ASAP7_75t_L g683 ( 
.A(n_585),
.Y(n_683)
);

BUFx3_ASAP7_75t_L g684 ( 
.A(n_598),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_627),
.Y(n_685)
);

AND2x2_ASAP7_75t_L g686 ( 
.A(n_634),
.B(n_622),
.Y(n_686)
);

OAI21x1_ASAP7_75t_L g687 ( 
.A1(n_632),
.A2(n_615),
.B(n_602),
.Y(n_687)
);

NAND2x1_ASAP7_75t_L g688 ( 
.A(n_654),
.B(n_629),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_SL g689 ( 
.A(n_618),
.B(n_558),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_667),
.B(n_560),
.Y(n_690)
);

OA22x2_ASAP7_75t_L g691 ( 
.A1(n_649),
.A2(n_575),
.B1(n_592),
.B2(n_605),
.Y(n_691)
);

NAND2x1p5_ASAP7_75t_L g692 ( 
.A(n_683),
.B(n_573),
.Y(n_692)
);

INVx3_ASAP7_75t_L g693 ( 
.A(n_654),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_631),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_619),
.B(n_585),
.Y(n_695)
);

OAI21x1_ASAP7_75t_L g696 ( 
.A1(n_682),
.A2(n_604),
.B(n_605),
.Y(n_696)
);

AOI22xp5_ASAP7_75t_L g697 ( 
.A1(n_648),
.A2(n_569),
.B1(n_585),
.B2(n_617),
.Y(n_697)
);

OAI22xp5_ASAP7_75t_L g698 ( 
.A1(n_619),
.A2(n_611),
.B1(n_596),
.B2(n_594),
.Y(n_698)
);

BUFx3_ASAP7_75t_L g699 ( 
.A(n_640),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_L g700 ( 
.A(n_624),
.B(n_585),
.Y(n_700)
);

OAI21x1_ASAP7_75t_L g701 ( 
.A1(n_682),
.A2(n_611),
.B(n_610),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_L g702 ( 
.A(n_624),
.B(n_585),
.Y(n_702)
);

INVx2_ASAP7_75t_SL g703 ( 
.A(n_635),
.Y(n_703)
);

INVx2_ASAP7_75t_L g704 ( 
.A(n_636),
.Y(n_704)
);

OAI21x1_ASAP7_75t_SL g705 ( 
.A1(n_638),
.A2(n_585),
.B(n_34),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_L g706 ( 
.A(n_639),
.B(n_0),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_662),
.B(n_1),
.Y(n_707)
);

INVx2_ASAP7_75t_L g708 ( 
.A(n_620),
.Y(n_708)
);

AOI21xp5_ASAP7_75t_L g709 ( 
.A1(n_683),
.A2(n_666),
.B(n_665),
.Y(n_709)
);

NOR2xp67_ASAP7_75t_SL g710 ( 
.A(n_683),
.B(n_416),
.Y(n_710)
);

OAI21x1_ASAP7_75t_L g711 ( 
.A1(n_659),
.A2(n_416),
.B(n_35),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_L g712 ( 
.A(n_633),
.B(n_2),
.Y(n_712)
);

AOI21x1_ASAP7_75t_L g713 ( 
.A1(n_665),
.A2(n_416),
.B(n_365),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_L g714 ( 
.A(n_633),
.B(n_2),
.Y(n_714)
);

AOI22xp33_ASAP7_75t_SL g715 ( 
.A1(n_684),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_646),
.B(n_3),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_L g717 ( 
.A(n_646),
.B(n_652),
.Y(n_717)
);

AOI21xp5_ASAP7_75t_L g718 ( 
.A1(n_666),
.A2(n_416),
.B(n_365),
.Y(n_718)
);

OAI21xp5_ASAP7_75t_L g719 ( 
.A1(n_669),
.A2(n_365),
.B(n_36),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_644),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_652),
.B(n_4),
.Y(n_721)
);

OAI21xp5_ASAP7_75t_L g722 ( 
.A1(n_674),
.A2(n_365),
.B(n_37),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_L g723 ( 
.A(n_663),
.B(n_5),
.Y(n_723)
);

AND2x2_ASAP7_75t_L g724 ( 
.A(n_658),
.B(n_6),
.Y(n_724)
);

AOI21xp5_ASAP7_75t_L g725 ( 
.A1(n_663),
.A2(n_365),
.B(n_40),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_L g726 ( 
.A(n_628),
.B(n_677),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_L g727 ( 
.A(n_679),
.B(n_6),
.Y(n_727)
);

AND2x6_ASAP7_75t_L g728 ( 
.A(n_680),
.B(n_33),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_L g729 ( 
.A(n_678),
.B(n_7),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_628),
.B(n_651),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_SL g731 ( 
.A(n_664),
.B(n_7),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_655),
.B(n_8),
.Y(n_732)
);

HB1xp67_ASAP7_75t_L g733 ( 
.A(n_653),
.Y(n_733)
);

OAI21xp5_ASAP7_75t_L g734 ( 
.A1(n_676),
.A2(n_43),
.B(n_41),
.Y(n_734)
);

OAI21x1_ASAP7_75t_L g735 ( 
.A1(n_642),
.A2(n_45),
.B(n_44),
.Y(n_735)
);

OAI21x1_ASAP7_75t_L g736 ( 
.A1(n_645),
.A2(n_48),
.B(n_47),
.Y(n_736)
);

AND2x2_ASAP7_75t_L g737 ( 
.A(n_625),
.B(n_8),
.Y(n_737)
);

NOR2x1_ASAP7_75t_SL g738 ( 
.A(n_643),
.B(n_49),
.Y(n_738)
);

AOI21xp5_ASAP7_75t_L g739 ( 
.A1(n_673),
.A2(n_52),
.B(n_51),
.Y(n_739)
);

BUFx10_ASAP7_75t_L g740 ( 
.A(n_657),
.Y(n_740)
);

OAI22x1_ASAP7_75t_L g741 ( 
.A1(n_656),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_741)
);

OAI21x1_ASAP7_75t_L g742 ( 
.A1(n_645),
.A2(n_54),
.B(n_53),
.Y(n_742)
);

OAI21x1_ASAP7_75t_L g743 ( 
.A1(n_647),
.A2(n_117),
.B(n_210),
.Y(n_743)
);

AND2x2_ASAP7_75t_L g744 ( 
.A(n_625),
.B(n_10),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_704),
.Y(n_745)
);

INVx2_ASAP7_75t_SL g746 ( 
.A(n_699),
.Y(n_746)
);

OAI21x1_ASAP7_75t_L g747 ( 
.A1(n_701),
.A2(n_647),
.B(n_676),
.Y(n_747)
);

O2A1O1Ixp5_ASAP7_75t_L g748 ( 
.A1(n_734),
.A2(n_621),
.B(n_656),
.C(n_680),
.Y(n_748)
);

BUFx2_ASAP7_75t_L g749 ( 
.A(n_733),
.Y(n_749)
);

INVx2_ASAP7_75t_L g750 ( 
.A(n_708),
.Y(n_750)
);

AO31x2_ASAP7_75t_L g751 ( 
.A1(n_709),
.A2(n_629),
.A3(n_675),
.B(n_670),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_L g752 ( 
.A(n_726),
.B(n_671),
.Y(n_752)
);

CKINVDCx5p33_ASAP7_75t_R g753 ( 
.A(n_703),
.Y(n_753)
);

A2O1A1Ixp33_ASAP7_75t_L g754 ( 
.A1(n_734),
.A2(n_664),
.B(n_621),
.C(n_673),
.Y(n_754)
);

BUFx6f_ASAP7_75t_L g755 ( 
.A(n_740),
.Y(n_755)
);

AO31x2_ASAP7_75t_L g756 ( 
.A1(n_698),
.A2(n_668),
.A3(n_650),
.B(n_643),
.Y(n_756)
);

NOR2xp33_ASAP7_75t_L g757 ( 
.A(n_686),
.B(n_626),
.Y(n_757)
);

AO31x2_ASAP7_75t_L g758 ( 
.A1(n_698),
.A2(n_643),
.A3(n_660),
.B(n_672),
.Y(n_758)
);

INVx2_ASAP7_75t_L g759 ( 
.A(n_685),
.Y(n_759)
);

AOI21xp5_ASAP7_75t_L g760 ( 
.A1(n_717),
.A2(n_672),
.B(n_637),
.Y(n_760)
);

AOI21xp5_ASAP7_75t_L g761 ( 
.A1(n_695),
.A2(n_672),
.B(n_637),
.Y(n_761)
);

INVx2_ASAP7_75t_L g762 ( 
.A(n_694),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_SL g763 ( 
.A(n_726),
.B(n_657),
.Y(n_763)
);

INVx3_ASAP7_75t_L g764 ( 
.A(n_740),
.Y(n_764)
);

AOI21xp5_ASAP7_75t_L g765 ( 
.A1(n_695),
.A2(n_702),
.B(n_700),
.Y(n_765)
);

OAI21x1_ASAP7_75t_L g766 ( 
.A1(n_687),
.A2(n_623),
.B(n_681),
.Y(n_766)
);

OAI21x1_ASAP7_75t_L g767 ( 
.A1(n_711),
.A2(n_623),
.B(n_681),
.Y(n_767)
);

O2A1O1Ixp33_ASAP7_75t_L g768 ( 
.A1(n_731),
.A2(n_689),
.B(n_729),
.C(n_727),
.Y(n_768)
);

NOR2x1_ASAP7_75t_SL g769 ( 
.A(n_690),
.B(n_641),
.Y(n_769)
);

A2O1A1Ixp33_ASAP7_75t_L g770 ( 
.A1(n_719),
.A2(n_657),
.B(n_681),
.C(n_641),
.Y(n_770)
);

OAI21x1_ASAP7_75t_L g771 ( 
.A1(n_696),
.A2(n_641),
.B(n_121),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_L g772 ( 
.A(n_730),
.B(n_661),
.Y(n_772)
);

INVx2_ASAP7_75t_SL g773 ( 
.A(n_737),
.Y(n_773)
);

AND2x4_ASAP7_75t_L g774 ( 
.A(n_720),
.B(n_55),
.Y(n_774)
);

AOI21xp5_ASAP7_75t_L g775 ( 
.A1(n_690),
.A2(n_119),
.B(n_211),
.Y(n_775)
);

AOI22xp33_ASAP7_75t_L g776 ( 
.A1(n_691),
.A2(n_630),
.B1(n_13),
.B2(n_14),
.Y(n_776)
);

OAI21x1_ASAP7_75t_L g777 ( 
.A1(n_713),
.A2(n_116),
.B(n_207),
.Y(n_777)
);

O2A1O1Ixp33_ASAP7_75t_L g778 ( 
.A1(n_712),
.A2(n_12),
.B(n_13),
.C(n_15),
.Y(n_778)
);

AND2x2_ASAP7_75t_L g779 ( 
.A(n_724),
.B(n_15),
.Y(n_779)
);

AO31x2_ASAP7_75t_L g780 ( 
.A1(n_725),
.A2(n_16),
.A3(n_17),
.B(n_18),
.Y(n_780)
);

AOI21xp5_ASAP7_75t_L g781 ( 
.A1(n_719),
.A2(n_722),
.B(n_730),
.Y(n_781)
);

OAI22xp5_ASAP7_75t_L g782 ( 
.A1(n_697),
.A2(n_16),
.B1(n_17),
.B2(n_18),
.Y(n_782)
);

O2A1O1Ixp33_ASAP7_75t_SL g783 ( 
.A1(n_707),
.A2(n_19),
.B(n_20),
.C(n_21),
.Y(n_783)
);

AO31x2_ASAP7_75t_L g784 ( 
.A1(n_718),
.A2(n_19),
.A3(n_20),
.B(n_21),
.Y(n_784)
);

NOR2xp67_ASAP7_75t_L g785 ( 
.A(n_714),
.B(n_56),
.Y(n_785)
);

INVx1_ASAP7_75t_SL g786 ( 
.A(n_744),
.Y(n_786)
);

AOI21xp5_ASAP7_75t_L g787 ( 
.A1(n_722),
.A2(n_208),
.B(n_129),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_L g788 ( 
.A(n_723),
.B(n_22),
.Y(n_788)
);

OAI21xp5_ASAP7_75t_L g789 ( 
.A1(n_691),
.A2(n_22),
.B(n_23),
.Y(n_789)
);

OAI21x1_ASAP7_75t_L g790 ( 
.A1(n_736),
.A2(n_130),
.B(n_202),
.Y(n_790)
);

NOR2xp33_ASAP7_75t_L g791 ( 
.A(n_716),
.B(n_57),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_723),
.B(n_721),
.Y(n_792)
);

NOR2xp33_ASAP7_75t_SL g793 ( 
.A(n_728),
.B(n_58),
.Y(n_793)
);

INVx2_ASAP7_75t_L g794 ( 
.A(n_693),
.Y(n_794)
);

AO32x2_ASAP7_75t_L g795 ( 
.A1(n_741),
.A2(n_23),
.A3(n_24),
.B1(n_25),
.B2(n_26),
.Y(n_795)
);

NOR2xp33_ASAP7_75t_L g796 ( 
.A(n_706),
.B(n_59),
.Y(n_796)
);

OR2x6_ASAP7_75t_L g797 ( 
.A(n_688),
.B(n_739),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_728),
.B(n_25),
.Y(n_798)
);

INVx2_ASAP7_75t_SL g799 ( 
.A(n_693),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_L g800 ( 
.A(n_728),
.B(n_26),
.Y(n_800)
);

O2A1O1Ixp33_ASAP7_75t_L g801 ( 
.A1(n_732),
.A2(n_27),
.B(n_28),
.C(n_29),
.Y(n_801)
);

OAI21x1_ASAP7_75t_L g802 ( 
.A1(n_742),
.A2(n_743),
.B(n_735),
.Y(n_802)
);

INVx4_ASAP7_75t_L g803 ( 
.A(n_728),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_738),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_L g805 ( 
.A(n_715),
.B(n_27),
.Y(n_805)
);

NOR2xp67_ASAP7_75t_L g806 ( 
.A(n_705),
.B(n_60),
.Y(n_806)
);

INVx2_ASAP7_75t_SL g807 ( 
.A(n_692),
.Y(n_807)
);

AOI21xp5_ASAP7_75t_L g808 ( 
.A1(n_692),
.A2(n_206),
.B(n_135),
.Y(n_808)
);

AO31x2_ASAP7_75t_L g809 ( 
.A1(n_710),
.A2(n_28),
.A3(n_29),
.B(n_30),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_726),
.B(n_30),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_704),
.Y(n_811)
);

BUFx2_ASAP7_75t_SL g812 ( 
.A(n_699),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_L g813 ( 
.A(n_726),
.B(n_31),
.Y(n_813)
);

AND2x2_ASAP7_75t_L g814 ( 
.A(n_752),
.B(n_61),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_759),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_762),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_745),
.Y(n_817)
);

INVx6_ASAP7_75t_L g818 ( 
.A(n_755),
.Y(n_818)
);

INVx3_ASAP7_75t_L g819 ( 
.A(n_774),
.Y(n_819)
);

AOI22xp33_ASAP7_75t_L g820 ( 
.A1(n_776),
.A2(n_31),
.B1(n_63),
.B2(n_64),
.Y(n_820)
);

INVx2_ASAP7_75t_L g821 ( 
.A(n_750),
.Y(n_821)
);

INVx6_ASAP7_75t_L g822 ( 
.A(n_755),
.Y(n_822)
);

AOI22xp33_ASAP7_75t_L g823 ( 
.A1(n_789),
.A2(n_65),
.B1(n_66),
.B2(n_67),
.Y(n_823)
);

BUFx2_ASAP7_75t_L g824 ( 
.A(n_749),
.Y(n_824)
);

CKINVDCx5p33_ASAP7_75t_R g825 ( 
.A(n_753),
.Y(n_825)
);

INVx2_ASAP7_75t_L g826 ( 
.A(n_811),
.Y(n_826)
);

AOI22xp33_ASAP7_75t_L g827 ( 
.A1(n_782),
.A2(n_68),
.B1(n_70),
.B2(n_71),
.Y(n_827)
);

BUFx2_ASAP7_75t_L g828 ( 
.A(n_773),
.Y(n_828)
);

AOI22xp33_ASAP7_75t_L g829 ( 
.A1(n_791),
.A2(n_73),
.B1(n_74),
.B2(n_77),
.Y(n_829)
);

AOI22xp33_ASAP7_75t_L g830 ( 
.A1(n_796),
.A2(n_79),
.B1(n_80),
.B2(n_82),
.Y(n_830)
);

AOI22xp33_ASAP7_75t_L g831 ( 
.A1(n_798),
.A2(n_85),
.B1(n_86),
.B2(n_89),
.Y(n_831)
);

BUFx12f_ASAP7_75t_L g832 ( 
.A(n_746),
.Y(n_832)
);

AND2x2_ASAP7_75t_L g833 ( 
.A(n_786),
.B(n_94),
.Y(n_833)
);

INVxp67_ASAP7_75t_L g834 ( 
.A(n_763),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_L g835 ( 
.A(n_792),
.B(n_95),
.Y(n_835)
);

INVx2_ASAP7_75t_SL g836 ( 
.A(n_755),
.Y(n_836)
);

OAI22xp33_ASAP7_75t_L g837 ( 
.A1(n_793),
.A2(n_96),
.B1(n_97),
.B2(n_100),
.Y(n_837)
);

BUFx3_ASAP7_75t_L g838 ( 
.A(n_764),
.Y(n_838)
);

INVx1_ASAP7_75t_SL g839 ( 
.A(n_812),
.Y(n_839)
);

OAI22xp5_ASAP7_75t_L g840 ( 
.A1(n_805),
.A2(n_101),
.B1(n_104),
.B2(n_106),
.Y(n_840)
);

BUFx2_ASAP7_75t_L g841 ( 
.A(n_799),
.Y(n_841)
);

INVx2_ASAP7_75t_L g842 ( 
.A(n_794),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_765),
.B(n_756),
.Y(n_843)
);

INVxp67_ASAP7_75t_SL g844 ( 
.A(n_747),
.Y(n_844)
);

AOI22xp5_ASAP7_75t_L g845 ( 
.A1(n_757),
.A2(n_107),
.B1(n_108),
.B2(n_109),
.Y(n_845)
);

BUFx3_ASAP7_75t_L g846 ( 
.A(n_772),
.Y(n_846)
);

BUFx3_ASAP7_75t_L g847 ( 
.A(n_774),
.Y(n_847)
);

AOI22xp33_ASAP7_75t_L g848 ( 
.A1(n_800),
.A2(n_110),
.B1(n_111),
.B2(n_112),
.Y(n_848)
);

BUFx6f_ASAP7_75t_L g849 ( 
.A(n_803),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_784),
.Y(n_850)
);

AOI22xp33_ASAP7_75t_SL g851 ( 
.A1(n_781),
.A2(n_113),
.B1(n_114),
.B2(n_115),
.Y(n_851)
);

AOI22xp33_ASAP7_75t_L g852 ( 
.A1(n_787),
.A2(n_122),
.B1(n_123),
.B2(n_124),
.Y(n_852)
);

AOI22xp5_ASAP7_75t_L g853 ( 
.A1(n_785),
.A2(n_125),
.B1(n_132),
.B2(n_133),
.Y(n_853)
);

NAND2x1p5_ASAP7_75t_L g854 ( 
.A(n_804),
.B(n_134),
.Y(n_854)
);

AOI22xp33_ASAP7_75t_SL g855 ( 
.A1(n_788),
.A2(n_137),
.B1(n_138),
.B2(n_139),
.Y(n_855)
);

BUFx2_ASAP7_75t_SL g856 ( 
.A(n_779),
.Y(n_856)
);

BUFx2_ASAP7_75t_L g857 ( 
.A(n_807),
.Y(n_857)
);

AOI22xp5_ASAP7_75t_SL g858 ( 
.A1(n_810),
.A2(n_140),
.B1(n_142),
.B2(n_143),
.Y(n_858)
);

INVx4_ASAP7_75t_L g859 ( 
.A(n_797),
.Y(n_859)
);

NOR2xp33_ASAP7_75t_L g860 ( 
.A(n_768),
.B(n_145),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_758),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_756),
.B(n_146),
.Y(n_862)
);

INVx6_ASAP7_75t_L g863 ( 
.A(n_797),
.Y(n_863)
);

AOI22xp33_ASAP7_75t_L g864 ( 
.A1(n_813),
.A2(n_148),
.B1(n_151),
.B2(n_152),
.Y(n_864)
);

AOI22xp33_ASAP7_75t_L g865 ( 
.A1(n_775),
.A2(n_153),
.B1(n_154),
.B2(n_156),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_758),
.Y(n_866)
);

OAI21xp5_ASAP7_75t_L g867 ( 
.A1(n_760),
.A2(n_162),
.B(n_163),
.Y(n_867)
);

AOI22xp33_ASAP7_75t_SL g868 ( 
.A1(n_795),
.A2(n_769),
.B1(n_783),
.B2(n_778),
.Y(n_868)
);

INVx2_ASAP7_75t_SL g869 ( 
.A(n_756),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_758),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_809),
.Y(n_871)
);

AND2x4_ASAP7_75t_L g872 ( 
.A(n_859),
.B(n_771),
.Y(n_872)
);

OAI21x1_ASAP7_75t_L g873 ( 
.A1(n_844),
.A2(n_802),
.B(n_777),
.Y(n_873)
);

AOI21x1_ASAP7_75t_L g874 ( 
.A1(n_871),
.A2(n_806),
.B(n_761),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_850),
.Y(n_875)
);

INVx2_ASAP7_75t_SL g876 ( 
.A(n_863),
.Y(n_876)
);

AOI22xp33_ASAP7_75t_L g877 ( 
.A1(n_860),
.A2(n_808),
.B1(n_790),
.B2(n_766),
.Y(n_877)
);

OAI22xp33_ASAP7_75t_L g878 ( 
.A1(n_846),
.A2(n_795),
.B1(n_801),
.B2(n_770),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_861),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_866),
.Y(n_880)
);

INVx4_ASAP7_75t_L g881 ( 
.A(n_863),
.Y(n_881)
);

HB1xp67_ASAP7_75t_L g882 ( 
.A(n_870),
.Y(n_882)
);

INVx2_ASAP7_75t_L g883 ( 
.A(n_817),
.Y(n_883)
);

OAI21xp5_ASAP7_75t_L g884 ( 
.A1(n_867),
.A2(n_748),
.B(n_754),
.Y(n_884)
);

INVx2_ASAP7_75t_L g885 ( 
.A(n_826),
.Y(n_885)
);

INVx4_ASAP7_75t_L g886 ( 
.A(n_863),
.Y(n_886)
);

AND2x2_ASAP7_75t_L g887 ( 
.A(n_844),
.B(n_780),
.Y(n_887)
);

INVx2_ASAP7_75t_L g888 ( 
.A(n_815),
.Y(n_888)
);

AND2x4_ASAP7_75t_L g889 ( 
.A(n_859),
.B(n_767),
.Y(n_889)
);

AND2x2_ASAP7_75t_L g890 ( 
.A(n_843),
.B(n_809),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_843),
.Y(n_891)
);

BUFx4f_ASAP7_75t_SL g892 ( 
.A(n_832),
.Y(n_892)
);

OAI21x1_ASAP7_75t_L g893 ( 
.A1(n_862),
.A2(n_780),
.B(n_809),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_816),
.Y(n_894)
);

HB1xp67_ASAP7_75t_L g895 ( 
.A(n_869),
.Y(n_895)
);

BUFx2_ASAP7_75t_L g896 ( 
.A(n_824),
.Y(n_896)
);

BUFx3_ASAP7_75t_L g897 ( 
.A(n_849),
.Y(n_897)
);

HB1xp67_ASAP7_75t_L g898 ( 
.A(n_834),
.Y(n_898)
);

BUFx3_ASAP7_75t_L g899 ( 
.A(n_849),
.Y(n_899)
);

AND2x2_ASAP7_75t_L g900 ( 
.A(n_862),
.B(n_821),
.Y(n_900)
);

AND2x2_ASAP7_75t_L g901 ( 
.A(n_834),
.B(n_780),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_842),
.Y(n_902)
);

AND2x2_ASAP7_75t_L g903 ( 
.A(n_868),
.B(n_795),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_857),
.Y(n_904)
);

BUFx2_ASAP7_75t_L g905 ( 
.A(n_841),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_835),
.Y(n_906)
);

INVx3_ASAP7_75t_L g907 ( 
.A(n_849),
.Y(n_907)
);

AND2x2_ASAP7_75t_L g908 ( 
.A(n_868),
.B(n_851),
.Y(n_908)
);

BUFx3_ASAP7_75t_L g909 ( 
.A(n_818),
.Y(n_909)
);

CKINVDCx20_ASAP7_75t_R g910 ( 
.A(n_825),
.Y(n_910)
);

AND2x4_ASAP7_75t_L g911 ( 
.A(n_819),
.B(n_751),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_835),
.B(n_751),
.Y(n_912)
);

BUFx3_ASAP7_75t_L g913 ( 
.A(n_818),
.Y(n_913)
);

INVxp67_ASAP7_75t_L g914 ( 
.A(n_896),
.Y(n_914)
);

OR2x2_ASAP7_75t_L g915 ( 
.A(n_891),
.B(n_856),
.Y(n_915)
);

OAI21x1_ASAP7_75t_L g916 ( 
.A1(n_873),
.A2(n_867),
.B(n_854),
.Y(n_916)
);

BUFx4f_ASAP7_75t_SL g917 ( 
.A(n_910),
.Y(n_917)
);

OA21x2_ASAP7_75t_L g918 ( 
.A1(n_893),
.A2(n_823),
.B(n_865),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_883),
.Y(n_919)
);

OAI21xp5_ASAP7_75t_L g920 ( 
.A1(n_884),
.A2(n_851),
.B(n_837),
.Y(n_920)
);

AND2x4_ASAP7_75t_L g921 ( 
.A(n_911),
.B(n_839),
.Y(n_921)
);

OR2x6_ASAP7_75t_L g922 ( 
.A(n_884),
.B(n_854),
.Y(n_922)
);

INVxp33_ASAP7_75t_L g923 ( 
.A(n_896),
.Y(n_923)
);

INVx2_ASAP7_75t_L g924 ( 
.A(n_885),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_L g925 ( 
.A(n_891),
.B(n_828),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_883),
.Y(n_926)
);

NOR2xp67_ASAP7_75t_R g927 ( 
.A(n_881),
.B(n_847),
.Y(n_927)
);

INVx2_ASAP7_75t_L g928 ( 
.A(n_885),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_883),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_885),
.Y(n_930)
);

INVx8_ASAP7_75t_L g931 ( 
.A(n_907),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_888),
.Y(n_932)
);

AOI222xp33_ASAP7_75t_L g933 ( 
.A1(n_908),
.A2(n_820),
.B1(n_840),
.B2(n_837),
.C1(n_827),
.C2(n_852),
.Y(n_933)
);

AO21x2_ASAP7_75t_L g934 ( 
.A1(n_912),
.A2(n_840),
.B(n_853),
.Y(n_934)
);

AOI21xp5_ASAP7_75t_L g935 ( 
.A1(n_878),
.A2(n_858),
.B(n_819),
.Y(n_935)
);

HB1xp67_ASAP7_75t_L g936 ( 
.A(n_898),
.Y(n_936)
);

NOR2xp33_ASAP7_75t_L g937 ( 
.A(n_892),
.B(n_838),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_888),
.Y(n_938)
);

INVxp67_ASAP7_75t_L g939 ( 
.A(n_905),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_888),
.Y(n_940)
);

NOR2x1_ASAP7_75t_L g941 ( 
.A(n_909),
.B(n_833),
.Y(n_941)
);

AO21x2_ASAP7_75t_L g942 ( 
.A1(n_912),
.A2(n_845),
.B(n_814),
.Y(n_942)
);

AND2x4_ASAP7_75t_L g943 ( 
.A(n_911),
.B(n_836),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_L g944 ( 
.A(n_900),
.B(n_751),
.Y(n_944)
);

HB1xp67_ASAP7_75t_L g945 ( 
.A(n_898),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_919),
.Y(n_946)
);

AND2x2_ASAP7_75t_L g947 ( 
.A(n_923),
.B(n_890),
.Y(n_947)
);

AND2x2_ASAP7_75t_L g948 ( 
.A(n_914),
.B(n_890),
.Y(n_948)
);

INVxp67_ASAP7_75t_SL g949 ( 
.A(n_936),
.Y(n_949)
);

AND2x2_ASAP7_75t_L g950 ( 
.A(n_939),
.B(n_901),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_926),
.Y(n_951)
);

AOI211xp5_ASAP7_75t_L g952 ( 
.A1(n_920),
.A2(n_878),
.B(n_908),
.C(n_903),
.Y(n_952)
);

AND2x2_ASAP7_75t_L g953 ( 
.A(n_945),
.B(n_901),
.Y(n_953)
);

INVx2_ASAP7_75t_L g954 ( 
.A(n_929),
.Y(n_954)
);

INVx1_ASAP7_75t_L g955 ( 
.A(n_932),
.Y(n_955)
);

CKINVDCx5p33_ASAP7_75t_R g956 ( 
.A(n_917),
.Y(n_956)
);

AOI22xp33_ASAP7_75t_L g957 ( 
.A1(n_920),
.A2(n_908),
.B1(n_903),
.B2(n_855),
.Y(n_957)
);

HB1xp67_ASAP7_75t_L g958 ( 
.A(n_944),
.Y(n_958)
);

BUFx2_ASAP7_75t_L g959 ( 
.A(n_921),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_L g960 ( 
.A(n_944),
.B(n_901),
.Y(n_960)
);

OR2x2_ASAP7_75t_L g961 ( 
.A(n_925),
.B(n_887),
.Y(n_961)
);

AND2x2_ASAP7_75t_L g962 ( 
.A(n_921),
.B(n_924),
.Y(n_962)
);

AND2x2_ASAP7_75t_L g963 ( 
.A(n_928),
.B(n_887),
.Y(n_963)
);

BUFx2_ASAP7_75t_L g964 ( 
.A(n_943),
.Y(n_964)
);

INVx1_ASAP7_75t_L g965 ( 
.A(n_938),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_940),
.Y(n_966)
);

BUFx3_ASAP7_75t_L g967 ( 
.A(n_931),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_946),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_946),
.Y(n_969)
);

OR2x2_ASAP7_75t_L g970 ( 
.A(n_961),
.B(n_925),
.Y(n_970)
);

AND2x2_ASAP7_75t_L g971 ( 
.A(n_964),
.B(n_943),
.Y(n_971)
);

AND2x2_ASAP7_75t_L g972 ( 
.A(n_964),
.B(n_915),
.Y(n_972)
);

AND2x4_ASAP7_75t_L g973 ( 
.A(n_967),
.B(n_911),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_951),
.Y(n_974)
);

AND2x2_ASAP7_75t_L g975 ( 
.A(n_958),
.B(n_930),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_L g976 ( 
.A(n_947),
.B(n_904),
.Y(n_976)
);

INVx2_ASAP7_75t_L g977 ( 
.A(n_954),
.Y(n_977)
);

AND2x2_ASAP7_75t_L g978 ( 
.A(n_959),
.B(n_905),
.Y(n_978)
);

AND2x2_ASAP7_75t_L g979 ( 
.A(n_959),
.B(n_911),
.Y(n_979)
);

INVx1_ASAP7_75t_L g980 ( 
.A(n_951),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_L g981 ( 
.A(n_947),
.B(n_904),
.Y(n_981)
);

AND2x2_ASAP7_75t_L g982 ( 
.A(n_953),
.B(n_889),
.Y(n_982)
);

OR2x2_ASAP7_75t_L g983 ( 
.A(n_961),
.B(n_960),
.Y(n_983)
);

AND2x2_ASAP7_75t_L g984 ( 
.A(n_953),
.B(n_950),
.Y(n_984)
);

INVx2_ASAP7_75t_L g985 ( 
.A(n_977),
.Y(n_985)
);

INVx3_ASAP7_75t_L g986 ( 
.A(n_973),
.Y(n_986)
);

AND2x2_ASAP7_75t_L g987 ( 
.A(n_972),
.B(n_950),
.Y(n_987)
);

OR2x2_ASAP7_75t_L g988 ( 
.A(n_976),
.B(n_960),
.Y(n_988)
);

INVx1_ASAP7_75t_L g989 ( 
.A(n_968),
.Y(n_989)
);

OR2x2_ASAP7_75t_L g990 ( 
.A(n_981),
.B(n_948),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_L g991 ( 
.A(n_969),
.B(n_952),
.Y(n_991)
);

OR2x2_ASAP7_75t_L g992 ( 
.A(n_970),
.B(n_948),
.Y(n_992)
);

AND2x2_ASAP7_75t_L g993 ( 
.A(n_972),
.B(n_962),
.Y(n_993)
);

INVx1_ASAP7_75t_L g994 ( 
.A(n_974),
.Y(n_994)
);

INVx1_ASAP7_75t_SL g995 ( 
.A(n_978),
.Y(n_995)
);

AND2x2_ASAP7_75t_L g996 ( 
.A(n_971),
.B(n_978),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_L g997 ( 
.A(n_980),
.B(n_952),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_L g998 ( 
.A(n_975),
.B(n_949),
.Y(n_998)
);

INVx1_ASAP7_75t_L g999 ( 
.A(n_989),
.Y(n_999)
);

OR2x2_ASAP7_75t_L g1000 ( 
.A(n_991),
.B(n_983),
.Y(n_1000)
);

INVxp67_ASAP7_75t_SL g1001 ( 
.A(n_991),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_L g1002 ( 
.A(n_997),
.B(n_975),
.Y(n_1002)
);

INVx1_ASAP7_75t_L g1003 ( 
.A(n_994),
.Y(n_1003)
);

INVx2_ASAP7_75t_L g1004 ( 
.A(n_986),
.Y(n_1004)
);

OR2x2_ASAP7_75t_L g1005 ( 
.A(n_997),
.B(n_984),
.Y(n_1005)
);

OR2x2_ASAP7_75t_L g1006 ( 
.A(n_990),
.B(n_992),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_985),
.Y(n_1007)
);

INVx1_ASAP7_75t_L g1008 ( 
.A(n_999),
.Y(n_1008)
);

AOI22xp5_ASAP7_75t_L g1009 ( 
.A1(n_1001),
.A2(n_957),
.B1(n_995),
.B2(n_903),
.Y(n_1009)
);

OAI22xp33_ASAP7_75t_L g1010 ( 
.A1(n_1005),
.A2(n_922),
.B1(n_935),
.B2(n_986),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_L g1011 ( 
.A(n_1002),
.B(n_996),
.Y(n_1011)
);

OR2x2_ASAP7_75t_L g1012 ( 
.A(n_1000),
.B(n_998),
.Y(n_1012)
);

NAND2x1_ASAP7_75t_L g1013 ( 
.A(n_1004),
.B(n_987),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_L g1014 ( 
.A(n_1002),
.B(n_993),
.Y(n_1014)
);

INVx1_ASAP7_75t_SL g1015 ( 
.A(n_1012),
.Y(n_1015)
);

AOI21xp5_ASAP7_75t_SL g1016 ( 
.A1(n_1009),
.A2(n_1008),
.B(n_1010),
.Y(n_1016)
);

NAND2x1p5_ASAP7_75t_L g1017 ( 
.A(n_1013),
.B(n_941),
.Y(n_1017)
);

INVx1_ASAP7_75t_L g1018 ( 
.A(n_1014),
.Y(n_1018)
);

NAND4xp25_ASAP7_75t_L g1019 ( 
.A(n_1011),
.B(n_933),
.C(n_1003),
.D(n_1007),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_L g1020 ( 
.A(n_1011),
.B(n_1006),
.Y(n_1020)
);

INVx1_ASAP7_75t_L g1021 ( 
.A(n_1008),
.Y(n_1021)
);

INVx2_ASAP7_75t_L g1022 ( 
.A(n_1013),
.Y(n_1022)
);

INVx1_ASAP7_75t_L g1023 ( 
.A(n_1008),
.Y(n_1023)
);

INVx1_ASAP7_75t_L g1024 ( 
.A(n_1008),
.Y(n_1024)
);

OAI22xp33_ASAP7_75t_L g1025 ( 
.A1(n_1017),
.A2(n_998),
.B1(n_922),
.B2(n_988),
.Y(n_1025)
);

INVxp67_ASAP7_75t_SL g1026 ( 
.A(n_1022),
.Y(n_1026)
);

NOR2xp67_ASAP7_75t_L g1027 ( 
.A(n_1019),
.B(n_956),
.Y(n_1027)
);

AND2x2_ASAP7_75t_L g1028 ( 
.A(n_1015),
.B(n_971),
.Y(n_1028)
);

INVx1_ASAP7_75t_SL g1029 ( 
.A(n_1020),
.Y(n_1029)
);

NOR2xp33_ASAP7_75t_L g1030 ( 
.A(n_1018),
.B(n_937),
.Y(n_1030)
);

NAND2xp5_ASAP7_75t_SL g1031 ( 
.A(n_1021),
.B(n_973),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_L g1032 ( 
.A(n_1023),
.B(n_984),
.Y(n_1032)
);

NAND2xp5_ASAP7_75t_L g1033 ( 
.A(n_1024),
.B(n_982),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_L g1034 ( 
.A(n_1026),
.B(n_1019),
.Y(n_1034)
);

AOI22xp5_ASAP7_75t_L g1035 ( 
.A1(n_1027),
.A2(n_1016),
.B1(n_922),
.B2(n_942),
.Y(n_1035)
);

NAND2x1_ASAP7_75t_SL g1036 ( 
.A(n_1028),
.B(n_985),
.Y(n_1036)
);

INVx1_ASAP7_75t_SL g1037 ( 
.A(n_1029),
.Y(n_1037)
);

OR2x2_ASAP7_75t_L g1038 ( 
.A(n_1032),
.B(n_949),
.Y(n_1038)
);

NOR2xp67_ASAP7_75t_L g1039 ( 
.A(n_1030),
.B(n_977),
.Y(n_1039)
);

INVxp67_ASAP7_75t_L g1040 ( 
.A(n_1031),
.Y(n_1040)
);

BUFx2_ASAP7_75t_L g1041 ( 
.A(n_1033),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_1025),
.Y(n_1042)
);

INVx1_ASAP7_75t_SL g1043 ( 
.A(n_1036),
.Y(n_1043)
);

OAI211xp5_ASAP7_75t_L g1044 ( 
.A1(n_1035),
.A2(n_855),
.B(n_933),
.C(n_830),
.Y(n_1044)
);

AOI22xp5_ASAP7_75t_L g1045 ( 
.A1(n_1040),
.A2(n_1037),
.B1(n_1042),
.B2(n_1034),
.Y(n_1045)
);

A2O1A1Ixp33_ASAP7_75t_L g1046 ( 
.A1(n_1039),
.A2(n_967),
.B(n_916),
.C(n_973),
.Y(n_1046)
);

INVxp67_ASAP7_75t_L g1047 ( 
.A(n_1041),
.Y(n_1047)
);

OAI21xp33_ASAP7_75t_SL g1048 ( 
.A1(n_1038),
.A2(n_979),
.B(n_982),
.Y(n_1048)
);

INVxp67_ASAP7_75t_L g1049 ( 
.A(n_1034),
.Y(n_1049)
);

INVx1_ASAP7_75t_L g1050 ( 
.A(n_1036),
.Y(n_1050)
);

INVx2_ASAP7_75t_L g1051 ( 
.A(n_1050),
.Y(n_1051)
);

INVxp67_ASAP7_75t_L g1052 ( 
.A(n_1043),
.Y(n_1052)
);

INVx1_ASAP7_75t_L g1053 ( 
.A(n_1045),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_1047),
.Y(n_1054)
);

CKINVDCx5p33_ASAP7_75t_R g1055 ( 
.A(n_1049),
.Y(n_1055)
);

INVx3_ASAP7_75t_L g1056 ( 
.A(n_1048),
.Y(n_1056)
);

INVx2_ASAP7_75t_L g1057 ( 
.A(n_1046),
.Y(n_1057)
);

INVx1_ASAP7_75t_L g1058 ( 
.A(n_1044),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_1045),
.Y(n_1059)
);

INVxp33_ASAP7_75t_SL g1060 ( 
.A(n_1045),
.Y(n_1060)
);

INVx1_ASAP7_75t_L g1061 ( 
.A(n_1045),
.Y(n_1061)
);

NOR2x1_ASAP7_75t_L g1062 ( 
.A(n_1053),
.B(n_967),
.Y(n_1062)
);

AOI22xp5_ASAP7_75t_L g1063 ( 
.A1(n_1060),
.A2(n_1061),
.B1(n_1059),
.B2(n_1054),
.Y(n_1063)
);

NAND4xp25_ASAP7_75t_L g1064 ( 
.A(n_1058),
.B(n_829),
.C(n_831),
.D(n_848),
.Y(n_1064)
);

INVx1_ASAP7_75t_L g1065 ( 
.A(n_1056),
.Y(n_1065)
);

XNOR2xp5_ASAP7_75t_L g1066 ( 
.A(n_1055),
.B(n_897),
.Y(n_1066)
);

NOR2xp33_ASAP7_75t_SL g1067 ( 
.A(n_1052),
.B(n_818),
.Y(n_1067)
);

XOR2x2_ASAP7_75t_L g1068 ( 
.A(n_1052),
.B(n_942),
.Y(n_1068)
);

OAI211xp5_ASAP7_75t_L g1069 ( 
.A1(n_1051),
.A2(n_864),
.B(n_899),
.C(n_897),
.Y(n_1069)
);

INVx1_ASAP7_75t_L g1070 ( 
.A(n_1056),
.Y(n_1070)
);

NAND4xp75_ASAP7_75t_L g1071 ( 
.A(n_1057),
.B(n_979),
.C(n_906),
.D(n_876),
.Y(n_1071)
);

AOI21xp5_ASAP7_75t_L g1072 ( 
.A1(n_1060),
.A2(n_934),
.B(n_927),
.Y(n_1072)
);

NOR2xp67_ASAP7_75t_L g1073 ( 
.A(n_1065),
.B(n_164),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_L g1074 ( 
.A(n_1070),
.B(n_1063),
.Y(n_1074)
);

NAND2xp5_ASAP7_75t_SL g1075 ( 
.A(n_1062),
.B(n_1067),
.Y(n_1075)
);

NOR2xp33_ASAP7_75t_L g1076 ( 
.A(n_1066),
.B(n_822),
.Y(n_1076)
);

NAND4xp75_ASAP7_75t_L g1077 ( 
.A(n_1072),
.B(n_906),
.C(n_876),
.D(n_918),
.Y(n_1077)
);

NAND4xp75_ASAP7_75t_L g1078 ( 
.A(n_1068),
.B(n_876),
.C(n_918),
.D(n_822),
.Y(n_1078)
);

NOR2x1_ASAP7_75t_L g1079 ( 
.A(n_1071),
.B(n_897),
.Y(n_1079)
);

OAI21xp33_ASAP7_75t_L g1080 ( 
.A1(n_1069),
.A2(n_899),
.B(n_909),
.Y(n_1080)
);

OAI21xp5_ASAP7_75t_SL g1081 ( 
.A1(n_1074),
.A2(n_1064),
.B(n_907),
.Y(n_1081)
);

NAND4xp25_ASAP7_75t_L g1082 ( 
.A(n_1076),
.B(n_899),
.C(n_907),
.D(n_877),
.Y(n_1082)
);

OAI221xp5_ASAP7_75t_L g1083 ( 
.A1(n_1080),
.A2(n_822),
.B1(n_907),
.B2(n_886),
.C(n_881),
.Y(n_1083)
);

INVx1_ASAP7_75t_L g1084 ( 
.A(n_1073),
.Y(n_1084)
);

NAND2xp5_ASAP7_75t_SL g1085 ( 
.A(n_1079),
.B(n_913),
.Y(n_1085)
);

AOI311xp33_ASAP7_75t_L g1086 ( 
.A1(n_1075),
.A2(n_966),
.A3(n_965),
.B(n_955),
.C(n_894),
.Y(n_1086)
);

NAND3xp33_ASAP7_75t_SL g1087 ( 
.A(n_1078),
.B(n_881),
.C(n_886),
.Y(n_1087)
);

NAND4xp75_ASAP7_75t_L g1088 ( 
.A(n_1077),
.B(n_962),
.C(n_965),
.D(n_966),
.Y(n_1088)
);

AND2x4_ASAP7_75t_L g1089 ( 
.A(n_1073),
.B(n_913),
.Y(n_1089)
);

NOR2x1p5_ASAP7_75t_L g1090 ( 
.A(n_1084),
.B(n_1089),
.Y(n_1090)
);

INVx1_ASAP7_75t_L g1091 ( 
.A(n_1089),
.Y(n_1091)
);

NOR3xp33_ASAP7_75t_L g1092 ( 
.A(n_1081),
.B(n_881),
.C(n_886),
.Y(n_1092)
);

INVx1_ASAP7_75t_L g1093 ( 
.A(n_1085),
.Y(n_1093)
);

INVx1_ASAP7_75t_L g1094 ( 
.A(n_1088),
.Y(n_1094)
);

NOR3xp33_ASAP7_75t_L g1095 ( 
.A(n_1087),
.B(n_886),
.C(n_893),
.Y(n_1095)
);

NOR3xp33_ASAP7_75t_L g1096 ( 
.A(n_1083),
.B(n_893),
.C(n_900),
.Y(n_1096)
);

NOR2x1_ASAP7_75t_L g1097 ( 
.A(n_1082),
.B(n_913),
.Y(n_1097)
);

NOR2x1_ASAP7_75t_L g1098 ( 
.A(n_1086),
.B(n_909),
.Y(n_1098)
);

OR2x2_ASAP7_75t_L g1099 ( 
.A(n_1084),
.B(n_955),
.Y(n_1099)
);

INVx1_ASAP7_75t_L g1100 ( 
.A(n_1091),
.Y(n_1100)
);

AND2x4_ASAP7_75t_L g1101 ( 
.A(n_1090),
.B(n_954),
.Y(n_1101)
);

NOR2xp67_ASAP7_75t_L g1102 ( 
.A(n_1093),
.B(n_168),
.Y(n_1102)
);

NOR2x1_ASAP7_75t_L g1103 ( 
.A(n_1094),
.B(n_934),
.Y(n_1103)
);

NOR2xp33_ASAP7_75t_L g1104 ( 
.A(n_1099),
.B(n_170),
.Y(n_1104)
);

INVx5_ASAP7_75t_L g1105 ( 
.A(n_1092),
.Y(n_1105)
);

OR2x2_ASAP7_75t_L g1106 ( 
.A(n_1095),
.B(n_1096),
.Y(n_1106)
);

BUFx2_ASAP7_75t_L g1107 ( 
.A(n_1098),
.Y(n_1107)
);

AND3x1_ASAP7_75t_L g1108 ( 
.A(n_1097),
.B(n_954),
.C(n_927),
.Y(n_1108)
);

AND2x2_ASAP7_75t_L g1109 ( 
.A(n_1091),
.B(n_963),
.Y(n_1109)
);

OR2x6_ASAP7_75t_L g1110 ( 
.A(n_1090),
.B(n_931),
.Y(n_1110)
);

INVx2_ASAP7_75t_L g1111 ( 
.A(n_1090),
.Y(n_1111)
);

AND2x2_ASAP7_75t_L g1112 ( 
.A(n_1091),
.B(n_963),
.Y(n_1112)
);

NOR3xp33_ASAP7_75t_L g1113 ( 
.A(n_1100),
.B(n_172),
.C(n_174),
.Y(n_1113)
);

XNOR2xp5_ASAP7_75t_L g1114 ( 
.A(n_1111),
.B(n_175),
.Y(n_1114)
);

INVx1_ASAP7_75t_L g1115 ( 
.A(n_1101),
.Y(n_1115)
);

NOR2xp67_ASAP7_75t_L g1116 ( 
.A(n_1102),
.B(n_176),
.Y(n_1116)
);

OAI22xp5_ASAP7_75t_L g1117 ( 
.A1(n_1110),
.A2(n_931),
.B1(n_872),
.B2(n_894),
.Y(n_1117)
);

OAI22xp5_ASAP7_75t_L g1118 ( 
.A1(n_1108),
.A2(n_872),
.B1(n_902),
.B2(n_889),
.Y(n_1118)
);

INVx1_ASAP7_75t_L g1119 ( 
.A(n_1107),
.Y(n_1119)
);

CKINVDCx20_ASAP7_75t_R g1120 ( 
.A(n_1105),
.Y(n_1120)
);

INVx1_ASAP7_75t_L g1121 ( 
.A(n_1109),
.Y(n_1121)
);

OAI211xp5_ASAP7_75t_L g1122 ( 
.A1(n_1119),
.A2(n_1105),
.B(n_1104),
.C(n_1106),
.Y(n_1122)
);

OAI22xp33_ASAP7_75t_L g1123 ( 
.A1(n_1120),
.A2(n_1103),
.B1(n_1112),
.B2(n_895),
.Y(n_1123)
);

AOI22xp33_ASAP7_75t_L g1124 ( 
.A1(n_1121),
.A2(n_872),
.B1(n_889),
.B2(n_900),
.Y(n_1124)
);

OAI22x1_ASAP7_75t_L g1125 ( 
.A1(n_1115),
.A2(n_872),
.B1(n_889),
.B2(n_874),
.Y(n_1125)
);

INVx2_ASAP7_75t_SL g1126 ( 
.A(n_1114),
.Y(n_1126)
);

HB1xp67_ASAP7_75t_L g1127 ( 
.A(n_1116),
.Y(n_1127)
);

OAI22xp5_ASAP7_75t_SL g1128 ( 
.A1(n_1117),
.A2(n_895),
.B1(n_902),
.B2(n_882),
.Y(n_1128)
);

AOI22xp5_ASAP7_75t_L g1129 ( 
.A1(n_1122),
.A2(n_1113),
.B1(n_1118),
.B2(n_887),
.Y(n_1129)
);

OAI21xp5_ASAP7_75t_L g1130 ( 
.A1(n_1127),
.A2(n_874),
.B(n_873),
.Y(n_1130)
);

INVx2_ASAP7_75t_L g1131 ( 
.A(n_1126),
.Y(n_1131)
);

NAND2xp5_ASAP7_75t_L g1132 ( 
.A(n_1129),
.B(n_1123),
.Y(n_1132)
);

HB1xp67_ASAP7_75t_L g1133 ( 
.A(n_1132),
.Y(n_1133)
);

INVx2_ASAP7_75t_L g1134 ( 
.A(n_1133),
.Y(n_1134)
);

AOI22xp5_ASAP7_75t_L g1135 ( 
.A1(n_1134),
.A2(n_1131),
.B1(n_1128),
.B2(n_1124),
.Y(n_1135)
);

OAI22xp33_ASAP7_75t_L g1136 ( 
.A1(n_1134),
.A2(n_1130),
.B1(n_1125),
.B2(n_882),
.Y(n_1136)
);

AOI22xp5_ASAP7_75t_L g1137 ( 
.A1(n_1134),
.A2(n_880),
.B1(n_879),
.B2(n_875),
.Y(n_1137)
);

XOR2xp5_ASAP7_75t_L g1138 ( 
.A(n_1135),
.B(n_177),
.Y(n_1138)
);

AOI21xp33_ASAP7_75t_SL g1139 ( 
.A1(n_1136),
.A2(n_178),
.B(n_180),
.Y(n_1139)
);

OAI21xp5_ASAP7_75t_L g1140 ( 
.A1(n_1137),
.A2(n_182),
.B(n_183),
.Y(n_1140)
);

INVx1_ASAP7_75t_L g1141 ( 
.A(n_1138),
.Y(n_1141)
);

OA21x2_ASAP7_75t_L g1142 ( 
.A1(n_1140),
.A2(n_185),
.B(n_187),
.Y(n_1142)
);

AOI221xp5_ASAP7_75t_L g1143 ( 
.A1(n_1141),
.A2(n_1139),
.B1(n_1142),
.B2(n_192),
.C(n_194),
.Y(n_1143)
);

AOI211xp5_ASAP7_75t_L g1144 ( 
.A1(n_1143),
.A2(n_190),
.B(n_191),
.C(n_195),
.Y(n_1144)
);


endmodule