module real_jpeg_7044_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_356;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_323;
wire n_215;
wire n_166;
wire n_176;
wire n_286;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_330;
wire n_298;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

INVx8_ASAP7_75t_L g79 ( 
.A(n_0),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_1),
.Y(n_109)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_1),
.Y(n_112)
);

BUFx3_ASAP7_75t_L g185 ( 
.A(n_1),
.Y(n_185)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_2),
.A2(n_116),
.B1(n_118),
.B2(n_122),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_2),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_L g195 ( 
.A1(n_2),
.A2(n_122),
.B1(n_196),
.B2(n_198),
.Y(n_195)
);

AOI22xp33_ASAP7_75t_SL g167 ( 
.A1(n_3),
.A2(n_168),
.B1(n_171),
.B2(n_174),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_3),
.Y(n_174)
);

OAI22xp33_ASAP7_75t_SL g211 ( 
.A1(n_3),
.A2(n_174),
.B1(n_212),
.B2(n_215),
.Y(n_211)
);

OAI22xp33_ASAP7_75t_SL g218 ( 
.A1(n_4),
.A2(n_219),
.B1(n_220),
.B2(n_221),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_4),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_5),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g252 ( 
.A1(n_5),
.A2(n_46),
.B1(n_120),
.B2(n_253),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_5),
.B(n_114),
.C(n_172),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g281 ( 
.A(n_5),
.B(n_75),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_5),
.B(n_270),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_5),
.B(n_103),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_5),
.B(n_330),
.Y(n_329)
);

AOI22xp33_ASAP7_75t_L g96 ( 
.A1(n_6),
.A2(n_90),
.B1(n_97),
.B2(n_100),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_6),
.Y(n_100)
);

OAI22xp33_ASAP7_75t_SL g265 ( 
.A1(n_6),
.A2(n_100),
.B1(n_219),
.B2(n_266),
.Y(n_265)
);

AOI22xp33_ASAP7_75t_SL g320 ( 
.A1(n_6),
.A2(n_100),
.B1(n_321),
.B2(n_323),
.Y(n_320)
);

AOI22xp33_ASAP7_75t_L g180 ( 
.A1(n_7),
.A2(n_168),
.B1(n_181),
.B2(n_182),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_7),
.Y(n_181)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_8),
.Y(n_66)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_9),
.Y(n_161)
);

INVx8_ASAP7_75t_L g178 ( 
.A(n_9),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g202 ( 
.A(n_9),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g226 ( 
.A(n_9),
.Y(n_226)
);

BUFx6f_ASAP7_75t_L g270 ( 
.A(n_9),
.Y(n_270)
);

BUFx5_ASAP7_75t_L g334 ( 
.A(n_9),
.Y(n_334)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_10),
.A2(n_87),
.B1(n_90),
.B2(n_94),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_10),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_10),
.A2(n_44),
.B1(n_94),
.B2(n_236),
.Y(n_235)
);

AOI22xp33_ASAP7_75t_L g278 ( 
.A1(n_10),
.A2(n_94),
.B1(n_215),
.B2(n_279),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_L g293 ( 
.A1(n_10),
.A2(n_94),
.B1(n_294),
.B2(n_297),
.Y(n_293)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_11),
.Y(n_42)
);

BUFx5_ASAP7_75t_L g151 ( 
.A(n_11),
.Y(n_151)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_12),
.Y(n_37)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_13),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_13),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_13),
.Y(n_55)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_13),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g237 ( 
.A(n_13),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_14),
.A2(n_54),
.B1(n_55),
.B2(n_56),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_14),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_14),
.A2(n_54),
.B1(n_119),
.B2(n_125),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_14),
.A2(n_54),
.B1(n_191),
.B2(n_192),
.Y(n_190)
);

AOI22xp33_ASAP7_75t_L g271 ( 
.A1(n_14),
.A2(n_54),
.B1(n_272),
.B2(n_274),
.Y(n_271)
);

BUFx3_ASAP7_75t_L g106 ( 
.A(n_15),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_15),
.Y(n_114)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_15),
.Y(n_134)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_15),
.Y(n_136)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

OAI22xp5_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_244),
.B1(n_245),
.B2(n_363),
.Y(n_17)
);

CKINVDCx16_ASAP7_75t_R g363 ( 
.A(n_18),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_243),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_205),
.Y(n_19)
);

OR2x2_ASAP7_75t_L g243 ( 
.A(n_20),
.B(n_205),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_139),
.C(n_186),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_L g359 ( 
.A(n_21),
.B(n_360),
.Y(n_359)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_23),
.B1(n_59),
.B2(n_138),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_22),
.B(n_60),
.C(n_101),
.Y(n_227)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

AOI21xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_43),
.B(n_51),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_24),
.B(n_53),
.Y(n_238)
);

AND2x2_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_34),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_28),
.B1(n_30),
.B2(n_31),
.Y(n_25)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

AOI22xp5_ASAP7_75t_L g34 ( 
.A1(n_32),
.A2(n_35),
.B1(n_38),
.B2(n_41),
.Y(n_34)
);

INVx6_ASAP7_75t_L g153 ( 
.A(n_32),
.Y(n_153)
);

INVx5_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_34),
.Y(n_58)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_37),
.Y(n_40)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_37),
.Y(n_70)
);

BUFx5_ASAP7_75t_L g93 ( 
.A(n_37),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_37),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g330 ( 
.A(n_37),
.Y(n_330)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx4_ASAP7_75t_L g191 ( 
.A(n_40),
.Y(n_191)
);

HB1xp67_ASAP7_75t_L g192 ( 
.A(n_40),
.Y(n_192)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

OAI21xp33_ASAP7_75t_SL g43 ( 
.A1(n_44),
.A2(n_46),
.B(n_47),
.Y(n_43)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_46),
.B(n_48),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_46),
.B(n_204),
.Y(n_203)
);

AOI21xp5_ASAP7_75t_L g290 ( 
.A1(n_46),
.A2(n_158),
.B(n_268),
.Y(n_290)
);

OAI21xp33_ASAP7_75t_SL g326 ( 
.A1(n_46),
.A2(n_327),
.B(n_328),
.Y(n_326)
);

OAI32xp33_ASAP7_75t_L g142 ( 
.A1(n_47),
.A2(n_143),
.A3(n_146),
.B1(n_149),
.B2(n_152),
.Y(n_142)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_53),
.B(n_58),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_55),
.Y(n_57)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx1_ASAP7_75t_SL g204 ( 
.A(n_58),
.Y(n_204)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_59),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_SL g59 ( 
.A(n_60),
.B(n_101),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_61),
.A2(n_86),
.B1(n_95),
.B2(n_96),
.Y(n_60)
);

INVx3_ASAP7_75t_SL g193 ( 
.A(n_61),
.Y(n_193)
);

OR2x2_ASAP7_75t_L g61 ( 
.A(n_62),
.B(n_75),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_L g62 ( 
.A1(n_63),
.A2(n_67),
.B1(n_71),
.B2(n_73),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_64),
.Y(n_76)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_65),
.Y(n_72)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_66),
.Y(n_85)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx5_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_69),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_70),
.Y(n_89)
);

BUFx5_ASAP7_75t_L g336 ( 
.A(n_70),
.Y(n_336)
);

NAND2xp33_ASAP7_75t_SL g343 ( 
.A(n_71),
.B(n_344),
.Y(n_343)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx1_ASAP7_75t_SL g95 ( 
.A(n_75),
.Y(n_95)
);

AO22x2_ASAP7_75t_L g75 ( 
.A1(n_76),
.A2(n_77),
.B1(n_80),
.B2(n_83),
.Y(n_75)
);

INVx4_ASAP7_75t_SL g279 ( 
.A(n_77),
.Y(n_279)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_79),
.Y(n_82)
);

INVx11_ASAP7_75t_L g121 ( 
.A(n_79),
.Y(n_121)
);

BUFx3_ASAP7_75t_L g131 ( 
.A(n_79),
.Y(n_131)
);

BUFx5_ASAP7_75t_L g261 ( 
.A(n_79),
.Y(n_261)
);

INVx3_ASAP7_75t_L g344 ( 
.A(n_79),
.Y(n_344)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_81),
.Y(n_117)
);

INVx4_ASAP7_75t_L g137 ( 
.A(n_81),
.Y(n_137)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx5_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx4_ASAP7_75t_L g342 ( 
.A(n_85),
.Y(n_342)
);

OAI21xp5_ASAP7_75t_SL g187 ( 
.A1(n_86),
.A2(n_95),
.B(n_188),
.Y(n_187)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

BUFx12f_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx5_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_95),
.B(n_190),
.Y(n_242)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_96),
.Y(n_241)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_99),
.Y(n_145)
);

INVx3_ASAP7_75t_L g155 ( 
.A(n_99),
.Y(n_155)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_99),
.Y(n_327)
);

OAI21xp5_ASAP7_75t_SL g101 ( 
.A1(n_102),
.A2(n_115),
.B(n_123),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_102),
.A2(n_115),
.B1(n_209),
.B2(n_210),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g319 ( 
.A1(n_102),
.A2(n_209),
.B1(n_278),
.B2(n_320),
.Y(n_319)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g257 ( 
.A(n_103),
.B(n_124),
.Y(n_257)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g127 ( 
.A(n_104),
.B(n_128),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_SL g277 ( 
.A1(n_104),
.A2(n_123),
.B(n_278),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_105),
.A2(n_107),
.B1(n_110),
.B2(n_113),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx3_ASAP7_75t_L g274 ( 
.A(n_107),
.Y(n_274)
);

INVx5_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx3_ASAP7_75t_L g170 ( 
.A(n_109),
.Y(n_170)
);

BUFx5_ASAP7_75t_L g219 ( 
.A(n_109),
.Y(n_219)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx8_ASAP7_75t_L g298 ( 
.A(n_111),
.Y(n_298)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_112),
.Y(n_165)
);

BUFx3_ASAP7_75t_L g173 ( 
.A(n_112),
.Y(n_173)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx11_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx5_ASAP7_75t_L g126 ( 
.A(n_121),
.Y(n_126)
);

INVx6_ASAP7_75t_L g256 ( 
.A(n_121),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_127),
.Y(n_123)
);

INVx4_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx5_ASAP7_75t_L g322 ( 
.A(n_126),
.Y(n_322)
);

INVx2_ASAP7_75t_SL g209 ( 
.A(n_127),
.Y(n_209)
);

OAI22xp33_ASAP7_75t_L g128 ( 
.A1(n_129),
.A2(n_132),
.B1(n_135),
.B2(n_137),
.Y(n_128)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx3_ASAP7_75t_L g214 ( 
.A(n_131),
.Y(n_214)
);

INVx4_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVx5_ASAP7_75t_SL g215 ( 
.A(n_137),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g360 ( 
.A1(n_139),
.A2(n_140),
.B1(n_186),
.B2(n_361),
.Y(n_360)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_141),
.A2(n_142),
.B1(n_156),
.B2(n_157),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_142),
.B(n_156),
.Y(n_231)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_154),
.Y(n_152)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_158),
.A2(n_166),
.B1(n_175),
.B2(n_179),
.Y(n_157)
);

AOI21xp5_ASAP7_75t_L g264 ( 
.A1(n_158),
.A2(n_265),
.B(n_268),
.Y(n_264)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_159),
.A2(n_167),
.B1(n_195),
.B2(n_201),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_159),
.A2(n_180),
.B1(n_217),
.B2(n_224),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_159),
.B(n_271),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_SL g305 ( 
.A1(n_159),
.A2(n_306),
.B1(n_307),
.B2(n_308),
.Y(n_305)
);

OR2x2_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_162),
.Y(n_159)
);

INVx3_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

INVx3_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

INVx5_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_165),
.Y(n_200)
);

BUFx6f_ASAP7_75t_L g223 ( 
.A(n_165),
.Y(n_223)
);

INVxp67_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

INVx3_ASAP7_75t_L g273 ( 
.A(n_170),
.Y(n_273)
);

BUFx3_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_173),
.Y(n_296)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

INVx4_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_178),
.Y(n_309)
);

INVxp67_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

INVx8_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

BUFx2_ASAP7_75t_L g197 ( 
.A(n_184),
.Y(n_197)
);

BUFx8_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

BUFx5_ASAP7_75t_L g288 ( 
.A(n_185),
.Y(n_288)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_186),
.Y(n_361)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_194),
.C(n_203),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_SL g353 ( 
.A(n_187),
.B(n_354),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_193),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

AOI21xp5_ASAP7_75t_L g240 ( 
.A1(n_193),
.A2(n_241),
.B(n_242),
.Y(n_240)
);

AOI21xp5_ASAP7_75t_L g325 ( 
.A1(n_193),
.A2(n_242),
.B(n_326),
.Y(n_325)
);

XOR2xp5_ASAP7_75t_L g354 ( 
.A(n_194),
.B(n_203),
.Y(n_354)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_195),
.Y(n_333)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

INVx4_ASAP7_75t_SL g267 ( 
.A(n_199),
.Y(n_267)
);

INVx4_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVx3_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_L g234 ( 
.A1(n_204),
.A2(n_235),
.B(n_238),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_230),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_207),
.A2(n_227),
.B1(n_228),
.B2(n_229),
.Y(n_206)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_207),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_216),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_SL g251 ( 
.A1(n_209),
.A2(n_252),
.B(n_257),
.Y(n_251)
);

OAI21xp5_ASAP7_75t_SL g351 ( 
.A1(n_209),
.A2(n_257),
.B(n_320),
.Y(n_351)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

INVx3_ASAP7_75t_L g323 ( 
.A(n_215),
.Y(n_323)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

INVx6_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

BUFx6f_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

INVx4_ASAP7_75t_L g300 ( 
.A(n_226),
.Y(n_300)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_227),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_232),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_233),
.A2(n_234),
.B1(n_239),
.B2(n_240),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

INVx4_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

AOI21x1_ASAP7_75t_L g245 ( 
.A1(n_246),
.A2(n_357),
.B(n_362),
.Y(n_245)
);

AO21x1_ASAP7_75t_SL g246 ( 
.A1(n_247),
.A2(n_346),
.B(n_356),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_SL g247 ( 
.A1(n_248),
.A2(n_314),
.B(n_345),
.Y(n_247)
);

AOI21xp5_ASAP7_75t_L g248 ( 
.A1(n_249),
.A2(n_282),
.B(n_313),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_263),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_250),
.B(n_263),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_251),
.B(n_258),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g310 ( 
.A1(n_251),
.A2(n_258),
.B1(n_259),
.B2(n_311),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_251),
.Y(n_311)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

HB1xp67_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

INVx2_ASAP7_75t_L g339 ( 
.A(n_256),
.Y(n_339)
);

CKINVDCx16_ASAP7_75t_R g258 ( 
.A(n_259),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_262),
.Y(n_259)
);

INVx3_ASAP7_75t_SL g260 ( 
.A(n_261),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_264),
.B(n_275),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_264),
.B(n_276),
.C(n_281),
.Y(n_315)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_265),
.Y(n_307)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_271),
.Y(n_268)
);

INVx3_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_276),
.A2(n_277),
.B1(n_280),
.B2(n_281),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_L g282 ( 
.A1(n_283),
.A2(n_304),
.B(n_312),
.Y(n_282)
);

AOI21xp5_ASAP7_75t_L g283 ( 
.A1(n_284),
.A2(n_291),
.B(n_303),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_285),
.B(n_290),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_286),
.B(n_289),
.Y(n_285)
);

INVx1_ASAP7_75t_SL g286 ( 
.A(n_287),
.Y(n_286)
);

INVx3_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g291 ( 
.A(n_292),
.B(n_302),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_292),
.B(n_302),
.Y(n_303)
);

AOI21xp5_ASAP7_75t_L g292 ( 
.A1(n_293),
.A2(n_299),
.B(n_301),
.Y(n_292)
);

INVxp67_ASAP7_75t_L g306 ( 
.A(n_293),
.Y(n_306)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

INVx4_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

INVx3_ASAP7_75t_SL g299 ( 
.A(n_300),
.Y(n_299)
);

AOI21xp5_ASAP7_75t_L g332 ( 
.A1(n_301),
.A2(n_333),
.B(n_334),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_305),
.B(n_310),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_305),
.B(n_310),
.Y(n_312)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_315),
.B(n_316),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_315),
.B(n_316),
.Y(n_345)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_317),
.B(n_331),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_318),
.A2(n_319),
.B1(n_324),
.B2(n_325),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_319),
.B(n_324),
.C(n_331),
.Y(n_347)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);

INVxp33_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

AOI32xp33_ASAP7_75t_L g335 ( 
.A1(n_329),
.A2(n_336),
.A3(n_337),
.B1(n_340),
.B2(n_343),
.Y(n_335)
);

XOR2xp5_ASAP7_75t_L g331 ( 
.A(n_332),
.B(n_335),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g352 ( 
.A(n_332),
.B(n_335),
.Y(n_352)
);

BUFx2_ASAP7_75t_L g337 ( 
.A(n_338),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_339),
.Y(n_338)
);

INVx4_ASAP7_75t_L g340 ( 
.A(n_341),
.Y(n_340)
);

INVx8_ASAP7_75t_L g341 ( 
.A(n_342),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_347),
.B(n_348),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_SL g356 ( 
.A(n_347),
.B(n_348),
.Y(n_356)
);

AOI22xp5_ASAP7_75t_L g348 ( 
.A1(n_349),
.A2(n_350),
.B1(n_353),
.B2(n_355),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_350),
.Y(n_349)
);

XNOR2xp5_ASAP7_75t_SL g350 ( 
.A(n_351),
.B(n_352),
.Y(n_350)
);

MAJIxp5_ASAP7_75t_L g358 ( 
.A(n_351),
.B(n_352),
.C(n_355),
.Y(n_358)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_353),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_358),
.B(n_359),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_SL g362 ( 
.A(n_358),
.B(n_359),
.Y(n_362)
);


endmodule