module fake_netlist_1_525_n_32 (n_1, n_2, n_6, n_4, n_3, n_5, n_7, n_8, n_0, n_32);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_5;
input n_7;
input n_8;
input n_0;
output n_32;
wire n_20;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_30;
wire n_13;
wire n_26;
wire n_18;
wire n_12;
wire n_9;
wire n_17;
wire n_14;
wire n_10;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_27;
INVx2_ASAP7_75t_L g9 ( .A(n_2), .Y(n_9) );
INVx2_ASAP7_75t_L g10 ( .A(n_4), .Y(n_10) );
BUFx6f_ASAP7_75t_L g11 ( .A(n_1), .Y(n_11) );
INVx2_ASAP7_75t_L g12 ( .A(n_6), .Y(n_12) );
INVx1_ASAP7_75t_L g13 ( .A(n_9), .Y(n_13) );
INVx1_ASAP7_75t_L g14 ( .A(n_10), .Y(n_14) );
BUFx8_ASAP7_75t_SL g15 ( .A(n_11), .Y(n_15) );
AOI21xp5_ASAP7_75t_L g16 ( .A1(n_12), .A2(n_8), .B(n_7), .Y(n_16) );
INVx1_ASAP7_75t_L g17 ( .A(n_13), .Y(n_17) );
BUFx3_ASAP7_75t_L g18 ( .A(n_13), .Y(n_18) );
AND2x2_ASAP7_75t_SL g19 ( .A(n_14), .B(n_5), .Y(n_19) );
AOI221xp5_ASAP7_75t_L g20 ( .A1(n_17), .A2(n_14), .B1(n_16), .B2(n_15), .C(n_3), .Y(n_20) );
BUFx3_ASAP7_75t_L g21 ( .A(n_18), .Y(n_21) );
INVx1_ASAP7_75t_L g22 ( .A(n_18), .Y(n_22) );
AND2x2_ASAP7_75t_L g23 ( .A(n_21), .B(n_19), .Y(n_23) );
INVx2_ASAP7_75t_L g24 ( .A(n_21), .Y(n_24) );
INVx1_ASAP7_75t_L g25 ( .A(n_24), .Y(n_25) );
INVx1_ASAP7_75t_SL g26 ( .A(n_23), .Y(n_26) );
NAND3xp33_ASAP7_75t_L g27 ( .A(n_25), .B(n_20), .C(n_19), .Y(n_27) );
NAND4xp75_ASAP7_75t_L g28 ( .A(n_25), .B(n_19), .C(n_17), .D(n_22), .Y(n_28) );
INVx2_ASAP7_75t_L g29 ( .A(n_28), .Y(n_29) );
BUFx2_ASAP7_75t_L g30 ( .A(n_27), .Y(n_30) );
INVx1_ASAP7_75t_L g31 ( .A(n_30), .Y(n_31) );
AOI322xp5_ASAP7_75t_L g32 ( .A1(n_31), .A2(n_29), .A3(n_26), .B1(n_3), .B2(n_4), .C1(n_2), .C2(n_0), .Y(n_32) );
endmodule