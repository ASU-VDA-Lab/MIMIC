module real_jpeg_5044_n_4 (n_3, n_1, n_0, n_2, n_4);

input n_3;
input n_1;
input n_0;
input n_2;

output n_4;

wire n_5;
wire n_8;
wire n_12;
wire n_11;
wire n_14;
wire n_13;
wire n_6;
wire n_7;
wire n_10;
wire n_9;

A2O1A1Ixp33_ASAP7_75t_L g4 ( 
.A1(n_0),
.A2(n_5),
.B(n_8),
.C(n_14),
.Y(n_4)
);

INVx1_ASAP7_75t_L g9 ( 
.A(n_0),
.Y(n_9)
);

INVx1_ASAP7_75t_L g10 ( 
.A(n_1),
.Y(n_10)
);

INVx13_ASAP7_75t_L g14 ( 
.A(n_2),
.Y(n_14)
);

INVx3_ASAP7_75t_L g7 ( 
.A(n_3),
.Y(n_7)
);

INVx3_ASAP7_75t_L g5 ( 
.A(n_6),
.Y(n_5)
);

INVx5_ASAP7_75t_L g6 ( 
.A(n_7),
.Y(n_6)
);

INVx8_ASAP7_75t_L g13 ( 
.A(n_7),
.Y(n_13)
);

AOI211xp5_ASAP7_75t_L g8 ( 
.A1(n_9),
.A2(n_10),
.B(n_11),
.C(n_12),
.Y(n_8)
);

NOR2xp33_ASAP7_75t_L g11 ( 
.A(n_9),
.B(n_10),
.Y(n_11)
);

INVx5_ASAP7_75t_L g12 ( 
.A(n_13),
.Y(n_12)
);


endmodule