module fake_netlist_6_3254_n_4109 (n_52, n_435, n_1, n_91, n_326, n_256, n_209, n_367, n_63, n_223, n_278, n_341, n_362, n_148, n_226, n_161, n_22, n_208, n_68, n_316, n_419, n_28, n_304, n_212, n_50, n_7, n_144, n_365, n_125, n_168, n_384, n_297, n_342, n_77, n_106, n_358, n_160, n_131, n_188, n_310, n_186, n_245, n_0, n_368, n_396, n_350, n_78, n_84, n_392, n_142, n_143, n_382, n_180, n_62, n_349, n_233, n_255, n_284, n_400, n_140, n_337, n_214, n_67, n_15, n_246, n_38, n_289, n_421, n_424, n_59, n_181, n_182, n_238, n_202, n_320, n_108, n_327, n_369, n_280, n_287, n_353, n_389, n_415, n_65, n_230, n_141, n_383, n_200, n_176, n_114, n_86, n_198, n_104, n_222, n_179, n_248, n_300, n_71, n_74, n_229, n_305, n_72, n_173, n_250, n_372, n_111, n_314, n_378, n_413, n_377, n_35, n_183, n_79, n_375, n_338, n_56, n_360, n_119, n_235, n_147, n_191, n_340, n_387, n_39, n_344, n_73, n_428, n_432, n_101, n_167, n_174, n_127, n_153, n_156, n_145, n_42, n_133, n_96, n_8, n_371, n_189, n_405, n_213, n_294, n_302, n_380, n_129, n_197, n_11, n_137, n_17, n_343, n_20, n_397, n_155, n_109, n_425, n_122, n_45, n_34, n_218, n_70, n_234, n_37, n_381, n_82, n_27, n_236, n_112, n_172, n_270, n_239, n_126, n_414, n_97, n_58, n_290, n_220, n_118, n_224, n_48, n_25, n_93, n_80, n_196, n_402, n_352, n_9, n_107, n_6, n_417, n_14, n_89, n_374, n_366, n_407, n_103, n_272, n_185, n_348, n_69, n_376, n_390, n_293, n_31, n_334, n_53, n_370, n_44, n_232, n_16, n_163, n_46, n_330, n_298, n_18, n_281, n_258, n_154, n_98, n_260, n_265, n_313, n_279, n_252, n_228, n_356, n_166, n_184, n_216, n_83, n_363, n_395, n_323, n_393, n_411, n_152, n_92, n_321, n_331, n_105, n_227, n_132, n_406, n_102, n_204, n_261, n_420, n_312, n_394, n_32, n_66, n_130, n_164, n_292, n_100, n_121, n_307, n_433, n_23, n_2, n_291, n_219, n_357, n_150, n_264, n_263, n_325, n_329, n_33, n_408, n_61, n_237, n_244, n_399, n_76, n_243, n_124, n_94, n_282, n_436, n_116, n_211, n_117, n_175, n_322, n_345, n_409, n_231, n_354, n_40, n_240, n_139, n_319, n_41, n_134, n_273, n_95, n_311, n_10, n_403, n_253, n_123, n_136, n_249, n_201, n_386, n_159, n_157, n_162, n_115, n_128, n_241, n_30, n_275, n_43, n_276, n_221, n_423, n_146, n_318, n_303, n_306, n_21, n_193, n_269, n_359, n_346, n_88, n_3, n_416, n_277, n_418, n_113, n_4, n_199, n_138, n_266, n_296, n_268, n_271, n_404, n_439, n_158, n_217, n_49, n_210, n_299, n_206, n_5, n_333, n_215, n_178, n_247, n_225, n_308, n_309, n_355, n_426, n_317, n_149, n_431, n_90, n_347, n_24, n_54, n_328, n_429, n_373, n_87, n_195, n_285, n_85, n_99, n_257, n_13, n_203, n_286, n_254, n_207, n_242, n_19, n_47, n_29, n_75, n_401, n_324, n_335, n_430, n_205, n_120, n_251, n_301, n_274, n_110, n_151, n_412, n_81, n_36, n_26, n_55, n_267, n_438, n_339, n_315, n_434, n_64, n_288, n_427, n_422, n_135, n_165, n_351, n_437, n_259, n_177, n_391, n_364, n_295, n_385, n_388, n_190, n_262, n_187, n_60, n_361, n_379, n_170, n_332, n_336, n_12, n_398, n_410, n_194, n_171, n_192, n_57, n_169, n_51, n_283, n_4109);

input n_52;
input n_435;
input n_1;
input n_91;
input n_326;
input n_256;
input n_209;
input n_367;
input n_63;
input n_223;
input n_278;
input n_341;
input n_362;
input n_148;
input n_226;
input n_161;
input n_22;
input n_208;
input n_68;
input n_316;
input n_419;
input n_28;
input n_304;
input n_212;
input n_50;
input n_7;
input n_144;
input n_365;
input n_125;
input n_168;
input n_384;
input n_297;
input n_342;
input n_77;
input n_106;
input n_358;
input n_160;
input n_131;
input n_188;
input n_310;
input n_186;
input n_245;
input n_0;
input n_368;
input n_396;
input n_350;
input n_78;
input n_84;
input n_392;
input n_142;
input n_143;
input n_382;
input n_180;
input n_62;
input n_349;
input n_233;
input n_255;
input n_284;
input n_400;
input n_140;
input n_337;
input n_214;
input n_67;
input n_15;
input n_246;
input n_38;
input n_289;
input n_421;
input n_424;
input n_59;
input n_181;
input n_182;
input n_238;
input n_202;
input n_320;
input n_108;
input n_327;
input n_369;
input n_280;
input n_287;
input n_353;
input n_389;
input n_415;
input n_65;
input n_230;
input n_141;
input n_383;
input n_200;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_179;
input n_248;
input n_300;
input n_71;
input n_74;
input n_229;
input n_305;
input n_72;
input n_173;
input n_250;
input n_372;
input n_111;
input n_314;
input n_378;
input n_413;
input n_377;
input n_35;
input n_183;
input n_79;
input n_375;
input n_338;
input n_56;
input n_360;
input n_119;
input n_235;
input n_147;
input n_191;
input n_340;
input n_387;
input n_39;
input n_344;
input n_73;
input n_428;
input n_432;
input n_101;
input n_167;
input n_174;
input n_127;
input n_153;
input n_156;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_371;
input n_189;
input n_405;
input n_213;
input n_294;
input n_302;
input n_380;
input n_129;
input n_197;
input n_11;
input n_137;
input n_17;
input n_343;
input n_20;
input n_397;
input n_155;
input n_109;
input n_425;
input n_122;
input n_45;
input n_34;
input n_218;
input n_70;
input n_234;
input n_37;
input n_381;
input n_82;
input n_27;
input n_236;
input n_112;
input n_172;
input n_270;
input n_239;
input n_126;
input n_414;
input n_97;
input n_58;
input n_290;
input n_220;
input n_118;
input n_224;
input n_48;
input n_25;
input n_93;
input n_80;
input n_196;
input n_402;
input n_352;
input n_9;
input n_107;
input n_6;
input n_417;
input n_14;
input n_89;
input n_374;
input n_366;
input n_407;
input n_103;
input n_272;
input n_185;
input n_348;
input n_69;
input n_376;
input n_390;
input n_293;
input n_31;
input n_334;
input n_53;
input n_370;
input n_44;
input n_232;
input n_16;
input n_163;
input n_46;
input n_330;
input n_298;
input n_18;
input n_281;
input n_258;
input n_154;
input n_98;
input n_260;
input n_265;
input n_313;
input n_279;
input n_252;
input n_228;
input n_356;
input n_166;
input n_184;
input n_216;
input n_83;
input n_363;
input n_395;
input n_323;
input n_393;
input n_411;
input n_152;
input n_92;
input n_321;
input n_331;
input n_105;
input n_227;
input n_132;
input n_406;
input n_102;
input n_204;
input n_261;
input n_420;
input n_312;
input n_394;
input n_32;
input n_66;
input n_130;
input n_164;
input n_292;
input n_100;
input n_121;
input n_307;
input n_433;
input n_23;
input n_2;
input n_291;
input n_219;
input n_357;
input n_150;
input n_264;
input n_263;
input n_325;
input n_329;
input n_33;
input n_408;
input n_61;
input n_237;
input n_244;
input n_399;
input n_76;
input n_243;
input n_124;
input n_94;
input n_282;
input n_436;
input n_116;
input n_211;
input n_117;
input n_175;
input n_322;
input n_345;
input n_409;
input n_231;
input n_354;
input n_40;
input n_240;
input n_139;
input n_319;
input n_41;
input n_134;
input n_273;
input n_95;
input n_311;
input n_10;
input n_403;
input n_253;
input n_123;
input n_136;
input n_249;
input n_201;
input n_386;
input n_159;
input n_157;
input n_162;
input n_115;
input n_128;
input n_241;
input n_30;
input n_275;
input n_43;
input n_276;
input n_221;
input n_423;
input n_146;
input n_318;
input n_303;
input n_306;
input n_21;
input n_193;
input n_269;
input n_359;
input n_346;
input n_88;
input n_3;
input n_416;
input n_277;
input n_418;
input n_113;
input n_4;
input n_199;
input n_138;
input n_266;
input n_296;
input n_268;
input n_271;
input n_404;
input n_439;
input n_158;
input n_217;
input n_49;
input n_210;
input n_299;
input n_206;
input n_5;
input n_333;
input n_215;
input n_178;
input n_247;
input n_225;
input n_308;
input n_309;
input n_355;
input n_426;
input n_317;
input n_149;
input n_431;
input n_90;
input n_347;
input n_24;
input n_54;
input n_328;
input n_429;
input n_373;
input n_87;
input n_195;
input n_285;
input n_85;
input n_99;
input n_257;
input n_13;
input n_203;
input n_286;
input n_254;
input n_207;
input n_242;
input n_19;
input n_47;
input n_29;
input n_75;
input n_401;
input n_324;
input n_335;
input n_430;
input n_205;
input n_120;
input n_251;
input n_301;
input n_274;
input n_110;
input n_151;
input n_412;
input n_81;
input n_36;
input n_26;
input n_55;
input n_267;
input n_438;
input n_339;
input n_315;
input n_434;
input n_64;
input n_288;
input n_427;
input n_422;
input n_135;
input n_165;
input n_351;
input n_437;
input n_259;
input n_177;
input n_391;
input n_364;
input n_295;
input n_385;
input n_388;
input n_190;
input n_262;
input n_187;
input n_60;
input n_361;
input n_379;
input n_170;
input n_332;
input n_336;
input n_12;
input n_398;
input n_410;
input n_194;
input n_171;
input n_192;
input n_57;
input n_169;
input n_51;
input n_283;

output n_4109;

wire n_992;
wire n_2542;
wire n_1671;
wire n_2817;
wire n_3660;
wire n_3813;
wire n_801;
wire n_3766;
wire n_1613;
wire n_1234;
wire n_2576;
wire n_1458;
wire n_3254;
wire n_3684;
wire n_1199;
wire n_1674;
wire n_3392;
wire n_741;
wire n_1027;
wire n_1351;
wire n_3266;
wire n_3574;
wire n_625;
wire n_1189;
wire n_3152;
wire n_3579;
wire n_1212;
wire n_726;
wire n_2157;
wire n_3335;
wire n_2332;
wire n_3773;
wire n_700;
wire n_3783;
wire n_1307;
wire n_3178;
wire n_2003;
wire n_3849;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_3844;
wire n_1237;
wire n_1061;
wire n_2534;
wire n_2353;
wire n_3089;
wire n_3301;
wire n_4099;
wire n_1357;
wire n_1853;
wire n_3741;
wire n_783;
wire n_2451;
wire n_1738;
wire n_2243;
wire n_798;
wire n_1575;
wire n_1854;
wire n_2324;
wire n_3088;
wire n_3443;
wire n_1923;
wire n_3257;
wire n_509;
wire n_1342;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_2260;
wire n_3222;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_2977;
wire n_3952;
wire n_1739;
wire n_2051;
wire n_2317;
wire n_1380;
wire n_3911;
wire n_2359;
wire n_442;
wire n_480;
wire n_2847;
wire n_1402;
wire n_2557;
wire n_1691;
wire n_1688;
wire n_3332;
wire n_3465;
wire n_1975;
wire n_1009;
wire n_1930;
wire n_1743;
wire n_2405;
wire n_3706;
wire n_4050;
wire n_1160;
wire n_883;
wire n_2647;
wire n_1238;
wire n_1991;
wire n_2570;
wire n_2179;
wire n_2386;
wire n_2997;
wire n_4092;
wire n_1724;
wire n_1032;
wire n_3708;
wire n_2336;
wire n_1247;
wire n_3668;
wire n_4078;
wire n_1547;
wire n_2521;
wire n_3376;
wire n_3046;
wire n_2956;
wire n_1553;
wire n_893;
wire n_1099;
wire n_2491;
wire n_3801;
wire n_1264;
wire n_1192;
wire n_471;
wire n_3564;
wire n_1844;
wire n_3619;
wire n_4087;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_2211;
wire n_1370;
wire n_1786;
wire n_3487;
wire n_2382;
wire n_3754;
wire n_2672;
wire n_3030;
wire n_2291;
wire n_830;
wire n_2299;
wire n_3340;
wire n_461;
wire n_873;
wire n_1371;
wire n_1285;
wire n_2886;
wire n_2974;
wire n_3946;
wire n_1985;
wire n_2989;
wire n_447;
wire n_2838;
wire n_2184;
wire n_3395;
wire n_2982;
wire n_1803;
wire n_3427;
wire n_1172;
wire n_852;
wire n_2509;
wire n_4065;
wire n_4026;
wire n_2513;
wire n_3282;
wire n_1590;
wire n_2645;
wire n_1532;
wire n_2628;
wire n_2313;
wire n_3071;
wire n_3626;
wire n_3757;
wire n_3904;
wire n_1393;
wire n_1517;
wire n_1867;
wire n_2926;
wire n_1704;
wire n_1078;
wire n_544;
wire n_1711;
wire n_2247;
wire n_3106;
wire n_1140;
wire n_2630;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_2344;
wire n_1579;
wire n_3275;
wire n_2365;
wire n_2470;
wire n_2321;
wire n_1263;
wire n_2019;
wire n_3031;
wire n_4029;
wire n_836;
wire n_3345;
wire n_2074;
wire n_2447;
wire n_522;
wire n_2919;
wire n_3678;
wire n_3440;
wire n_2129;
wire n_2340;
wire n_1261;
wire n_945;
wire n_3879;
wire n_4010;
wire n_2286;
wire n_1649;
wire n_2018;
wire n_2094;
wire n_3080;
wire n_1903;
wire n_1511;
wire n_1143;
wire n_2356;
wire n_2399;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_3979;
wire n_616;
wire n_658;
wire n_1874;
wire n_3165;
wire n_1119;
wire n_2865;
wire n_2825;
wire n_3463;
wire n_2013;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_2044;
wire n_1954;
wire n_1735;
wire n_2510;
wire n_2739;
wire n_1300;
wire n_641;
wire n_2480;
wire n_1541;
wire n_3023;
wire n_822;
wire n_3232;
wire n_693;
wire n_1313;
wire n_2791;
wire n_3607;
wire n_3750;
wire n_3251;
wire n_1056;
wire n_3877;
wire n_3316;
wire n_2212;
wire n_3929;
wire n_758;
wire n_516;
wire n_3494;
wire n_3048;
wire n_1455;
wire n_2418;
wire n_2864;
wire n_1163;
wire n_2729;
wire n_3063;
wire n_1180;
wire n_2256;
wire n_2582;
wire n_943;
wire n_1798;
wire n_4060;
wire n_1550;
wire n_2703;
wire n_491;
wire n_3998;
wire n_2786;
wire n_3371;
wire n_1591;
wire n_772;
wire n_3632;
wire n_3122;
wire n_2806;
wire n_1344;
wire n_3261;
wire n_2730;
wire n_2495;
wire n_666;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_1971;
wire n_2058;
wire n_2603;
wire n_2090;
wire n_2660;
wire n_538;
wire n_3028;
wire n_3829;
wire n_3662;
wire n_2981;
wire n_3076;
wire n_2173;
wire n_2004;
wire n_1106;
wire n_886;
wire n_1471;
wire n_953;
wire n_1094;
wire n_3624;
wire n_3077;
wire n_3737;
wire n_1345;
wire n_1820;
wire n_2873;
wire n_3452;
wire n_3655;
wire n_494;
wire n_539;
wire n_493;
wire n_3107;
wire n_3825;
wire n_2880;
wire n_3225;
wire n_2394;
wire n_2108;
wire n_3532;
wire n_454;
wire n_3948;
wire n_1421;
wire n_2836;
wire n_3664;
wire n_1936;
wire n_638;
wire n_1404;
wire n_1211;
wire n_2124;
wire n_2378;
wire n_887;
wire n_1660;
wire n_1961;
wire n_3047;
wire n_1280;
wire n_3765;
wire n_713;
wire n_2655;
wire n_1400;
wire n_2625;
wire n_3296;
wire n_2843;
wire n_1467;
wire n_3297;
wire n_976;
wire n_3760;
wire n_3067;
wire n_2155;
wire n_3906;
wire n_2686;
wire n_1445;
wire n_2364;
wire n_2551;
wire n_1560;
wire n_1526;
wire n_734;
wire n_1088;
wire n_1894;
wire n_2996;
wire n_1231;
wire n_2599;
wire n_2985;
wire n_1978;
wire n_3803;
wire n_2085;
wire n_3963;
wire n_3368;
wire n_917;
wire n_574;
wire n_3639;
wire n_3347;
wire n_2370;
wire n_2612;
wire n_3792;
wire n_907;
wire n_1446;
wire n_3938;
wire n_2591;
wire n_3507;
wire n_659;
wire n_1815;
wire n_2214;
wire n_3351;
wire n_913;
wire n_1658;
wire n_2593;
wire n_808;
wire n_867;
wire n_4071;
wire n_3506;
wire n_3568;
wire n_3269;
wire n_4047;
wire n_3531;
wire n_1230;
wire n_3413;
wire n_3850;
wire n_473;
wire n_1193;
wire n_1967;
wire n_3999;
wire n_1054;
wire n_3928;
wire n_559;
wire n_3412;
wire n_2613;
wire n_3535;
wire n_1333;
wire n_2496;
wire n_2708;
wire n_3313;
wire n_1648;
wire n_3189;
wire n_1911;
wire n_1956;
wire n_1644;
wire n_3791;
wire n_2011;
wire n_2725;
wire n_2277;
wire n_3164;
wire n_1558;
wire n_1732;
wire n_551;
wire n_699;
wire n_1986;
wire n_2300;
wire n_3943;
wire n_564;
wire n_2397;
wire n_3931;
wire n_3884;
wire n_451;
wire n_824;
wire n_686;
wire n_4102;
wire n_757;
wire n_594;
wire n_1641;
wire n_2113;
wire n_1918;
wire n_2190;
wire n_3603;
wire n_3871;
wire n_2907;
wire n_577;
wire n_3438;
wire n_2735;
wire n_1843;
wire n_619;
wire n_3959;
wire n_2268;
wire n_1367;
wire n_1336;
wire n_521;
wire n_2778;
wire n_2850;
wire n_572;
wire n_813;
wire n_1909;
wire n_2080;
wire n_1481;
wire n_3822;
wire n_606;
wire n_1441;
wire n_818;
wire n_3373;
wire n_1123;
wire n_1309;
wire n_2104;
wire n_513;
wire n_645;
wire n_1381;
wire n_2961;
wire n_3812;
wire n_1699;
wire n_3910;
wire n_916;
wire n_3934;
wire n_2093;
wire n_4033;
wire n_4009;
wire n_2633;
wire n_483;
wire n_3883;
wire n_2207;
wire n_1970;
wire n_2770;
wire n_608;
wire n_2101;
wire n_2696;
wire n_3482;
wire n_4080;
wire n_630;
wire n_2059;
wire n_2198;
wire n_3319;
wire n_541;
wire n_512;
wire n_2669;
wire n_2925;
wire n_3728;
wire n_4094;
wire n_2073;
wire n_2273;
wire n_3484;
wire n_3748;
wire n_2546;
wire n_3272;
wire n_3193;
wire n_792;
wire n_2522;
wire n_476;
wire n_3949;
wire n_2792;
wire n_1328;
wire n_3396;
wire n_1957;
wire n_2917;
wire n_2616;
wire n_3912;
wire n_3118;
wire n_3315;
wire n_3720;
wire n_1907;
wire n_3923;
wire n_2529;
wire n_3900;
wire n_1162;
wire n_860;
wire n_1530;
wire n_3798;
wire n_788;
wire n_939;
wire n_3488;
wire n_2811;
wire n_821;
wire n_1543;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_3732;
wire n_982;
wire n_2674;
wire n_2832;
wire n_549;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_3980;
wire n_932;
wire n_2831;
wire n_2998;
wire n_3446;
wire n_3317;
wire n_3857;
wire n_3978;
wire n_1876;
wire n_4107;
wire n_1895;
wire n_2123;
wire n_1697;
wire n_2143;
wire n_979;
wire n_4074;
wire n_3716;
wire n_1873;
wire n_905;
wire n_3630;
wire n_3518;
wire n_3824;
wire n_3859;
wire n_1866;
wire n_4013;
wire n_1680;
wire n_2692;
wire n_993;
wire n_3842;
wire n_689;
wire n_3248;
wire n_2031;
wire n_2130;
wire n_1413;
wire n_1330;
wire n_1605;
wire n_3914;
wire n_3514;
wire n_2228;
wire n_3714;
wire n_3397;
wire n_1988;
wire n_2941;
wire n_1278;
wire n_547;
wire n_3575;
wire n_2455;
wire n_2876;
wire n_558;
wire n_2654;
wire n_3036;
wire n_2469;
wire n_4032;
wire n_1064;
wire n_3099;
wire n_1396;
wire n_634;
wire n_2355;
wire n_3927;
wire n_966;
wire n_3888;
wire n_2908;
wire n_3168;
wire n_764;
wire n_2751;
wire n_2764;
wire n_3357;
wire n_1663;
wire n_2895;
wire n_2009;
wire n_692;
wire n_3403;
wire n_733;
wire n_1793;
wire n_2922;
wire n_3601;
wire n_3882;
wire n_1233;
wire n_1289;
wire n_2714;
wire n_2245;
wire n_487;
wire n_3092;
wire n_3055;
wire n_3492;
wire n_3895;
wire n_3966;
wire n_2068;
wire n_1107;
wire n_2866;
wire n_2457;
wire n_3294;
wire n_1014;
wire n_3734;
wire n_3686;
wire n_1290;
wire n_1703;
wire n_2580;
wire n_3455;
wire n_882;
wire n_2176;
wire n_2072;
wire n_3649;
wire n_1354;
wire n_2821;
wire n_586;
wire n_1865;
wire n_1875;
wire n_1701;
wire n_2459;
wire n_3746;
wire n_1111;
wire n_1713;
wire n_2971;
wire n_715;
wire n_3599;
wire n_2678;
wire n_1251;
wire n_3384;
wire n_3935;
wire n_1265;
wire n_2711;
wire n_3490;
wire n_1726;
wire n_1950;
wire n_530;
wire n_1563;
wire n_1912;
wire n_2434;
wire n_3369;
wire n_3419;
wire n_1982;
wire n_3872;
wire n_2878;
wire n_618;
wire n_3012;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_3875;
wire n_3772;
wire n_1167;
wire n_1359;
wire n_2818;
wire n_2428;
wire n_3581;
wire n_3794;
wire n_674;
wire n_3247;
wire n_871;
wire n_3069;
wire n_3921;
wire n_922;
wire n_1335;
wire n_1760;
wire n_1927;
wire n_2028;
wire n_3715;
wire n_1069;
wire n_2664;
wire n_1722;
wire n_1664;
wire n_612;
wire n_2641;
wire n_3022;
wire n_3052;
wire n_3725;
wire n_1165;
wire n_3933;
wire n_702;
wire n_2008;
wire n_2749;
wire n_3298;
wire n_2192;
wire n_3281;
wire n_2254;
wire n_2345;
wire n_3346;
wire n_1926;
wire n_1175;
wire n_3273;
wire n_1386;
wire n_2311;
wire n_1896;
wire n_2965;
wire n_1747;
wire n_3058;
wire n_1012;
wire n_3691;
wire n_780;
wire n_3861;
wire n_675;
wire n_2624;
wire n_4066;
wire n_903;
wire n_1540;
wire n_1977;
wire n_1802;
wire n_1504;
wire n_3549;
wire n_2350;
wire n_2804;
wire n_2453;
wire n_3891;
wire n_2193;
wire n_3961;
wire n_2676;
wire n_1655;
wire n_3940;
wire n_4072;
wire n_835;
wire n_928;
wire n_1214;
wire n_1801;
wire n_690;
wire n_850;
wire n_1886;
wire n_2347;
wire n_2092;
wire n_3917;
wire n_1654;
wire n_816;
wire n_1157;
wire n_3453;
wire n_1750;
wire n_2994;
wire n_1462;
wire n_3410;
wire n_3153;
wire n_3428;
wire n_1188;
wire n_3689;
wire n_1752;
wire n_877;
wire n_1813;
wire n_2514;
wire n_3768;
wire n_2206;
wire n_604;
wire n_4004;
wire n_2810;
wire n_2967;
wire n_2519;
wire n_2319;
wire n_4043;
wire n_825;
wire n_728;
wire n_2916;
wire n_3415;
wire n_1063;
wire n_1588;
wire n_3785;
wire n_3942;
wire n_3997;
wire n_2963;
wire n_4041;
wire n_2947;
wire n_3918;
wire n_2467;
wire n_2602;
wire n_2468;
wire n_3145;
wire n_1124;
wire n_1624;
wire n_3873;
wire n_3983;
wire n_515;
wire n_2096;
wire n_2980;
wire n_3968;
wire n_1965;
wire n_3538;
wire n_2476;
wire n_3280;
wire n_598;
wire n_3434;
wire n_696;
wire n_1515;
wire n_961;
wire n_3510;
wire n_1317;
wire n_1082;
wire n_3227;
wire n_2733;
wire n_2824;
wire n_3289;
wire n_593;
wire n_514;
wire n_4055;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_2377;
wire n_701;
wire n_2178;
wire n_3271;
wire n_950;
wire n_2812;
wire n_484;
wire n_2644;
wire n_2036;
wire n_3326;
wire n_2976;
wire n_2152;
wire n_1709;
wire n_3009;
wire n_2652;
wire n_3460;
wire n_2411;
wire n_3719;
wire n_2525;
wire n_1825;
wire n_2393;
wire n_1757;
wire n_1796;
wire n_2657;
wire n_1792;
wire n_3827;
wire n_891;
wire n_2067;
wire n_2136;
wire n_2921;
wire n_2409;
wire n_2082;
wire n_3519;
wire n_2252;
wire n_1412;
wire n_2497;
wire n_3889;
wire n_2687;
wire n_3237;
wire n_949;
wire n_1630;
wire n_678;
wire n_2887;
wire n_3809;
wire n_3500;
wire n_3834;
wire n_3526;
wire n_3707;
wire n_2075;
wire n_4045;
wire n_2194;
wire n_2972;
wire n_2619;
wire n_3139;
wire n_3542;
wire n_2763;
wire n_2762;
wire n_4070;
wire n_1987;
wire n_3545;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_3578;
wire n_3885;
wire n_881;
wire n_2271;
wire n_1008;
wire n_3192;
wire n_760;
wire n_3993;
wire n_1546;
wire n_2583;
wire n_590;
wire n_2606;
wire n_4031;
wire n_2279;
wire n_1033;
wire n_462;
wire n_1052;
wire n_2794;
wire n_1296;
wire n_2663;
wire n_1990;
wire n_3352;
wire n_2391;
wire n_3805;
wire n_2431;
wire n_3073;
wire n_4018;
wire n_2987;
wire n_694;
wire n_2938;
wire n_2150;
wire n_1294;
wire n_2943;
wire n_1420;
wire n_3696;
wire n_3780;
wire n_4082;
wire n_2078;
wire n_1634;
wire n_3252;
wire n_2932;
wire n_595;
wire n_627;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_3253;
wire n_3337;
wire n_3450;
wire n_3209;
wire n_4002;
wire n_2622;
wire n_1858;
wire n_1044;
wire n_2658;
wire n_2665;
wire n_2165;
wire n_2133;
wire n_1712;
wire n_3021;
wire n_1391;
wire n_449;
wire n_1523;
wire n_2558;
wire n_2750;
wire n_2775;
wire n_1208;
wire n_2893;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_2954;
wire n_3477;
wire n_2728;
wire n_2349;
wire n_3128;
wire n_3763;
wire n_2684;
wire n_2712;
wire n_1072;
wire n_3146;
wire n_1527;
wire n_1495;
wire n_3733;
wire n_1438;
wire n_495;
wire n_815;
wire n_3953;
wire n_1100;
wire n_585;
wire n_1487;
wire n_2691;
wire n_3421;
wire n_840;
wire n_2913;
wire n_3614;
wire n_874;
wire n_1756;
wire n_3183;
wire n_1128;
wire n_2493;
wire n_673;
wire n_2230;
wire n_2705;
wire n_1969;
wire n_4019;
wire n_2690;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_2145;
wire n_3405;
wire n_1968;
wire n_898;
wire n_1952;
wire n_865;
wire n_3616;
wire n_2573;
wire n_3423;
wire n_2646;
wire n_4044;
wire n_3436;
wire n_925;
wire n_1932;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_2535;
wire n_3442;
wire n_3366;
wire n_2631;
wire n_1364;
wire n_3078;
wire n_3644;
wire n_2436;
wire n_3937;
wire n_615;
wire n_2870;
wire n_1249;
wire n_2706;
wire n_3838;
wire n_1293;
wire n_2693;
wire n_1127;
wire n_1512;
wire n_2151;
wire n_3159;
wire n_1451;
wire n_3941;
wire n_639;
wire n_963;
wire n_794;
wire n_2767;
wire n_3793;
wire n_727;
wire n_894;
wire n_1839;
wire n_2341;
wire n_685;
wire n_1765;
wire n_3727;
wire n_2707;
wire n_3240;
wire n_3576;
wire n_3789;
wire n_605;
wire n_1514;
wire n_1863;
wire n_826;
wire n_3385;
wire n_3747;
wire n_3037;
wire n_1646;
wire n_3293;
wire n_872;
wire n_1139;
wire n_1714;
wire n_3922;
wire n_3179;
wire n_718;
wire n_1018;
wire n_3400;
wire n_3729;
wire n_1521;
wire n_1366;
wire n_4000;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_2537;
wire n_2897;
wire n_3970;
wire n_2554;
wire n_996;
wire n_532;
wire n_1308;
wire n_2089;
wire n_1376;
wire n_3522;
wire n_1513;
wire n_2747;
wire n_3924;
wire n_3171;
wire n_791;
wire n_1913;
wire n_3608;
wire n_510;
wire n_837;
wire n_2097;
wire n_2170;
wire n_3459;
wire n_3491;
wire n_1488;
wire n_2853;
wire n_1808;
wire n_3053;
wire n_948;
wire n_3358;
wire n_2517;
wire n_2713;
wire n_3499;
wire n_704;
wire n_2148;
wire n_977;
wire n_2339;
wire n_1005;
wire n_1947;
wire n_2765;
wire n_2861;
wire n_536;
wire n_3158;
wire n_1788;
wire n_3426;
wire n_1999;
wire n_2731;
wire n_622;
wire n_2643;
wire n_2590;
wire n_3150;
wire n_3018;
wire n_3353;
wire n_3782;
wire n_3975;
wire n_1469;
wire n_2060;
wire n_2608;
wire n_1838;
wire n_2638;
wire n_4011;
wire n_1835;
wire n_3470;
wire n_1766;
wire n_1776;
wire n_1959;
wire n_3133;
wire n_2002;
wire n_581;
wire n_2650;
wire n_2138;
wire n_4098;
wire n_4021;
wire n_765;
wire n_987;
wire n_1492;
wire n_3700;
wire n_2414;
wire n_1340;
wire n_3014;
wire n_3166;
wire n_1771;
wire n_2316;
wire n_4058;
wire n_4103;
wire n_3104;
wire n_631;
wire n_720;
wire n_3435;
wire n_842;
wire n_3148;
wire n_2262;
wire n_3229;
wire n_3348;
wire n_4022;
wire n_1707;
wire n_2239;
wire n_3082;
wire n_3611;
wire n_1432;
wire n_2208;
wire n_843;
wire n_656;
wire n_989;
wire n_2604;
wire n_2407;
wire n_1277;
wire n_2816;
wire n_797;
wire n_2689;
wire n_2933;
wire n_1473;
wire n_2191;
wire n_1723;
wire n_2717;
wire n_1246;
wire n_3799;
wire n_1878;
wire n_2574;
wire n_899;
wire n_738;
wire n_2012;
wire n_3497;
wire n_1304;
wire n_1035;
wire n_2842;
wire n_499;
wire n_2675;
wire n_1426;
wire n_3418;
wire n_705;
wire n_3580;
wire n_3775;
wire n_3537;
wire n_1004;
wire n_1176;
wire n_2134;
wire n_1529;
wire n_2335;
wire n_2473;
wire n_3887;
wire n_1022;
wire n_614;
wire n_529;
wire n_2069;
wire n_2307;
wire n_3704;
wire n_2362;
wire n_684;
wire n_2539;
wire n_2698;
wire n_2667;
wire n_4096;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_3312;
wire n_1571;
wire n_3835;
wire n_1809;
wire n_3119;
wire n_2958;
wire n_1577;
wire n_2948;
wire n_3735;
wire n_2297;
wire n_1181;
wire n_2119;
wire n_3731;
wire n_1822;
wire n_486;
wire n_947;
wire n_2936;
wire n_3224;
wire n_1117;
wire n_2489;
wire n_1087;
wire n_1448;
wire n_3173;
wire n_1992;
wire n_3677;
wire n_3631;
wire n_648;
wire n_657;
wire n_1049;
wire n_3223;
wire n_3996;
wire n_2771;
wire n_2445;
wire n_3020;
wire n_2057;
wire n_2103;
wire n_3140;
wire n_3185;
wire n_3770;
wire n_2605;
wire n_4097;
wire n_1666;
wire n_2772;
wire n_1505;
wire n_803;
wire n_1717;
wire n_926;
wire n_1817;
wire n_2449;
wire n_927;
wire n_3557;
wire n_2610;
wire n_3654;
wire n_3129;
wire n_3880;
wire n_1849;
wire n_2848;
wire n_919;
wire n_3685;
wire n_2868;
wire n_3620;
wire n_1698;
wire n_478;
wire n_4100;
wire n_2231;
wire n_3609;
wire n_929;
wire n_3832;
wire n_2520;
wire n_1228;
wire n_2857;
wire n_446;
wire n_3693;
wire n_3788;
wire n_1568;
wire n_1490;
wire n_2372;
wire n_777;
wire n_1299;
wire n_2896;
wire n_526;
wire n_3837;
wire n_2718;
wire n_3019;
wire n_2639;
wire n_3471;
wire n_1183;
wire n_1436;
wire n_2898;
wire n_2251;
wire n_1384;
wire n_3674;
wire n_2494;
wire n_2959;
wire n_4079;
wire n_2501;
wire n_3203;
wire n_3325;
wire n_2238;
wire n_4085;
wire n_2368;
wire n_458;
wire n_1070;
wire n_2403;
wire n_3342;
wire n_2837;
wire n_998;
wire n_717;
wire n_3200;
wire n_1665;
wire n_3600;
wire n_3259;
wire n_2524;
wire n_3167;
wire n_1383;
wire n_2460;
wire n_3390;
wire n_3656;
wire n_1178;
wire n_2127;
wire n_2338;
wire n_1424;
wire n_3324;
wire n_3593;
wire n_3341;
wire n_3867;
wire n_1073;
wire n_1000;
wire n_796;
wire n_1195;
wire n_3559;
wire n_3025;
wire n_2137;
wire n_1626;
wire n_3191;
wire n_4005;
wire n_2482;
wire n_1507;
wire n_552;
wire n_3810;
wire n_3546;
wire n_2532;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_3661;
wire n_3006;
wire n_2481;
wire n_3561;
wire n_912;
wire n_1857;
wire n_3987;
wire n_1519;
wire n_2144;
wire n_3056;
wire n_745;
wire n_1284;
wire n_2296;
wire n_2424;
wire n_1604;
wire n_3201;
wire n_3633;
wire n_3447;
wire n_3971;
wire n_1142;
wire n_2849;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_2354;
wire n_2682;
wire n_3032;
wire n_3103;
wire n_3638;
wire n_2589;
wire n_1395;
wire n_2110;
wire n_2199;
wire n_2661;
wire n_731;
wire n_2877;
wire n_1502;
wire n_1659;
wire n_1955;
wire n_755;
wire n_931;
wire n_1021;
wire n_3393;
wire n_474;
wire n_683;
wire n_527;
wire n_811;
wire n_1207;
wire n_2442;
wire n_3627;
wire n_1791;
wire n_1368;
wire n_3451;
wire n_3480;
wire n_1418;
wire n_958;
wire n_1250;
wire n_3331;
wire n_1137;
wire n_3615;
wire n_1897;
wire n_2064;
wire n_880;
wire n_3087;
wire n_3072;
wire n_2053;
wire n_3612;
wire n_3505;
wire n_2259;
wire n_2121;
wire n_2773;
wire n_2545;
wire n_3540;
wire n_3577;
wire n_889;
wire n_3509;
wire n_2432;
wire n_2710;
wire n_1478;
wire n_589;
wire n_3606;
wire n_1310;
wire n_3142;
wire n_3598;
wire n_819;
wire n_2966;
wire n_2294;
wire n_1363;
wire n_2581;
wire n_1334;
wire n_1942;
wire n_1966;
wire n_3591;
wire n_767;
wire n_3777;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_1837;
wire n_2788;
wire n_2218;
wire n_477;
wire n_3196;
wire n_3590;
wire n_2435;
wire n_954;
wire n_864;
wire n_2504;
wire n_2797;
wire n_2623;
wire n_1110;
wire n_2213;
wire n_1410;
wire n_2389;
wire n_1440;
wire n_2132;
wire n_2892;
wire n_2063;
wire n_1382;
wire n_1534;
wire n_3892;
wire n_1564;
wire n_1736;
wire n_4069;
wire n_2748;
wire n_4053;
wire n_1483;
wire n_3848;
wire n_1834;
wire n_2331;
wire n_1372;
wire n_2292;
wire n_2860;
wire n_3327;
wire n_2330;
wire n_3441;
wire n_1457;
wire n_505;
wire n_1719;
wire n_3534;
wire n_3718;
wire n_1339;
wire n_1787;
wire n_2701;
wire n_2475;
wire n_537;
wire n_2511;
wire n_3964;
wire n_1993;
wire n_2281;
wire n_1427;
wire n_2416;
wire n_2745;
wire n_2617;
wire n_2776;
wire n_1466;
wire n_1919;
wire n_1080;
wire n_723;
wire n_1877;
wire n_3144;
wire n_3705;
wire n_3211;
wire n_3244;
wire n_596;
wire n_3909;
wire n_3944;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_1939;
wire n_2030;
wire n_1769;
wire n_1220;
wire n_2323;
wire n_1893;
wire n_556;
wire n_2784;
wire n_2209;
wire n_2301;
wire n_3582;
wire n_3605;
wire n_3287;
wire n_2387;
wire n_3322;
wire n_1755;
wire n_1602;
wire n_2421;
wire n_1136;
wire n_3270;
wire n_2618;
wire n_2025;
wire n_2357;
wire n_2846;
wire n_2464;
wire n_3265;
wire n_1125;
wire n_3755;
wire n_4042;
wire n_970;
wire n_3306;
wire n_2488;
wire n_3640;
wire n_2224;
wire n_1980;
wire n_642;
wire n_995;
wire n_1159;
wire n_2329;
wire n_1092;
wire n_3481;
wire n_2237;
wire n_3026;
wire n_441;
wire n_1060;
wire n_1951;
wire n_2250;
wire n_3090;
wire n_444;
wire n_3033;
wire n_3724;
wire n_1252;
wire n_1784;
wire n_3311;
wire n_3571;
wire n_1223;
wire n_3913;
wire n_511;
wire n_2990;
wire n_3847;
wire n_1286;
wire n_1773;
wire n_1775;
wire n_2115;
wire n_2410;
wire n_2552;
wire n_1053;
wire n_3302;
wire n_2374;
wire n_1681;
wire n_520;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_2929;
wire n_2780;
wire n_3226;
wire n_3364;
wire n_3323;
wire n_4020;
wire n_2596;
wire n_2274;
wire n_3163;
wire n_775;
wire n_651;
wire n_1153;
wire n_1618;
wire n_3407;
wire n_518;
wire n_1531;
wire n_2828;
wire n_1185;
wire n_3856;
wire n_453;
wire n_3425;
wire n_2384;
wire n_3894;
wire n_1745;
wire n_914;
wire n_759;
wire n_3479;
wire n_3127;
wire n_2724;
wire n_1831;
wire n_2585;
wire n_2621;
wire n_3623;
wire n_1653;
wire n_2352;
wire n_1679;
wire n_4063;
wire n_1625;
wire n_3986;
wire n_2601;
wire n_2160;
wire n_3454;
wire n_1453;
wire n_2146;
wire n_4006;
wire n_2502;
wire n_2131;
wire n_488;
wire n_2226;
wire n_2801;
wire n_3646;
wire n_497;
wire n_2920;
wire n_4015;
wire n_773;
wire n_3547;
wire n_1901;
wire n_3869;
wire n_920;
wire n_1374;
wire n_2556;
wire n_2648;
wire n_3212;
wire n_1315;
wire n_1647;
wire n_2575;
wire n_2754;
wire n_1224;
wire n_2783;
wire n_3753;
wire n_2306;
wire n_1892;
wire n_1459;
wire n_1614;
wire n_3188;
wire n_3742;
wire n_1933;
wire n_2462;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_2889;
wire n_3243;
wire n_3683;
wire n_4034;
wire n_1617;
wire n_4056;
wire n_3260;
wire n_3370;
wire n_3386;
wire n_3816;
wire n_3960;
wire n_1470;
wire n_2550;
wire n_463;
wire n_3093;
wire n_3175;
wire n_3214;
wire n_1243;
wire n_3736;
wire n_848;
wire n_2732;
wire n_2928;
wire n_1096;
wire n_2249;
wire n_1091;
wire n_1917;
wire n_2000;
wire n_3862;
wire n_1580;
wire n_2227;
wire n_2270;
wire n_2822;
wire n_1425;
wire n_3169;
wire n_3205;
wire n_1881;
wire n_1267;
wire n_1281;
wire n_1806;
wire n_3284;
wire n_983;
wire n_3109;
wire n_2023;
wire n_3354;
wire n_2572;
wire n_2204;
wire n_1520;
wire n_496;
wire n_2720;
wire n_3126;
wire n_2159;
wire n_906;
wire n_1390;
wire n_688;
wire n_2315;
wire n_1077;
wire n_1733;
wire n_2289;
wire n_1419;
wire n_2863;
wire n_3299;
wire n_3663;
wire n_2955;
wire n_2995;
wire n_1731;
wire n_2158;
wire n_2087;
wire n_1855;
wire n_1636;
wire n_3051;
wire n_1437;
wire n_3360;
wire n_2135;
wire n_3956;
wire n_3367;
wire n_1832;
wire n_1645;
wire n_4001;
wire n_1687;
wire n_1439;
wire n_2328;
wire n_1323;
wire n_2859;
wire n_2202;
wire n_858;
wire n_2049;
wire n_1331;
wire n_613;
wire n_736;
wire n_2627;
wire n_501;
wire n_956;
wire n_960;
wire n_2276;
wire n_3234;
wire n_663;
wire n_856;
wire n_2803;
wire n_2100;
wire n_3314;
wire n_3525;
wire n_3016;
wire n_778;
wire n_1668;
wire n_2777;
wire n_1134;
wire n_2993;
wire n_3566;
wire n_3688;
wire n_3004;
wire n_3202;
wire n_2830;
wire n_2781;
wire n_3220;
wire n_4003;
wire n_1129;
wire n_3870;
wire n_554;
wire n_602;
wire n_1696;
wire n_2829;
wire n_1995;
wire n_1594;
wire n_2181;
wire n_3751;
wire n_664;
wire n_1869;
wire n_2911;
wire n_3625;
wire n_3804;
wire n_1764;
wire n_1429;
wire n_2826;
wire n_1610;
wire n_3084;
wire n_3429;
wire n_1889;
wire n_2379;
wire n_2016;
wire n_1905;
wire n_2343;
wire n_793;
wire n_587;
wire n_3466;
wire n_3554;
wire n_1593;
wire n_580;
wire n_762;
wire n_1202;
wire n_1030;
wire n_3901;
wire n_1937;
wire n_465;
wire n_1790;
wire n_1778;
wire n_3749;
wire n_1635;
wire n_2942;
wire n_4014;
wire n_1079;
wire n_2515;
wire n_1744;
wire n_828;
wire n_2139;
wire n_2142;
wire n_4067;
wire n_607;
wire n_1551;
wire n_4028;
wire n_4054;
wire n_2448;
wire n_1103;
wire n_2875;
wire n_3907;
wire n_2555;
wire n_4048;
wire n_3338;
wire n_3586;
wire n_3462;
wire n_3756;
wire n_2219;
wire n_1203;
wire n_3653;
wire n_3636;
wire n_2851;
wire n_3406;
wire n_820;
wire n_2327;
wire n_951;
wire n_2201;
wire n_725;
wire n_952;
wire n_3919;
wire n_999;
wire n_1254;
wire n_2841;
wire n_3349;
wire n_2420;
wire n_3722;
wire n_2984;
wire n_575;
wire n_994;
wire n_2263;
wire n_3539;
wire n_3291;
wire n_2304;
wire n_4024;
wire n_1508;
wire n_2487;
wire n_732;
wire n_974;
wire n_2983;
wire n_2240;
wire n_2278;
wire n_2656;
wire n_2538;
wire n_724;
wire n_2597;
wire n_2375;
wire n_3113;
wire n_3194;
wire n_3250;
wire n_1934;
wire n_3276;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_3981;
wire n_1728;
wire n_3973;
wire n_557;
wire n_2756;
wire n_3572;
wire n_1871;
wire n_3448;
wire n_617;
wire n_3886;
wire n_845;
wire n_807;
wire n_2924;
wire n_1036;
wire n_3595;
wire n_1138;
wire n_3414;
wire n_1661;
wire n_1275;
wire n_2884;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_3637;
wire n_3120;
wire n_1468;
wire n_3991;
wire n_2855;
wire n_3651;
wire n_1859;
wire n_2102;
wire n_3516;
wire n_2563;
wire n_3926;
wire n_3797;
wire n_1095;
wire n_2024;
wire n_1595;
wire n_2156;
wire n_3449;
wire n_1718;
wire n_1749;
wire n_3474;
wire n_1683;
wire n_1916;
wire n_2598;
wire n_597;
wire n_1270;
wire n_2549;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_4101;
wire n_3548;
wire n_3767;
wire n_1024;
wire n_3864;
wire n_4036;
wire n_1768;
wire n_2153;
wire n_2544;
wire n_2381;
wire n_3670;
wire n_3550;
wire n_3974;
wire n_1847;
wire n_2052;
wire n_3634;
wire n_2302;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_3230;
wire n_4016;
wire n_621;
wire n_1037;
wire n_1397;
wire n_3268;
wire n_3236;
wire n_1279;
wire n_750;
wire n_1115;
wire n_901;
wire n_1499;
wire n_3592;
wire n_468;
wire n_2755;
wire n_3141;
wire n_923;
wire n_504;
wire n_1409;
wire n_1841;
wire n_3839;
wire n_2637;
wire n_2823;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_3967;
wire n_1503;
wire n_3112;
wire n_2819;
wire n_3195;
wire n_466;
wire n_2526;
wire n_3041;
wire n_2423;
wire n_1057;
wire n_3277;
wire n_3108;
wire n_2548;
wire n_603;
wire n_991;
wire n_2785;
wire n_1657;
wire n_1126;
wire n_2412;
wire n_1997;
wire n_3817;
wire n_3417;
wire n_2636;
wire n_3131;
wire n_710;
wire n_1108;
wire n_1818;
wire n_2439;
wire n_2404;
wire n_1182;
wire n_3730;
wire n_1298;
wire n_3659;
wire n_2559;
wire n_2177;
wire n_2595;
wire n_3399;
wire n_2088;
wire n_3635;
wire n_1611;
wire n_785;
wire n_2740;
wire n_746;
wire n_609;
wire n_1601;
wire n_3011;
wire n_1960;
wire n_2694;
wire n_2061;
wire n_3416;
wire n_3648;
wire n_1686;
wire n_3498;
wire n_2757;
wire n_2401;
wire n_2337;
wire n_3042;
wire n_1356;
wire n_1589;
wire n_3213;
wire n_3820;
wire n_2309;
wire n_2900;
wire n_2957;
wire n_2607;
wire n_1740;
wire n_2737;
wire n_3994;
wire n_1497;
wire n_2890;
wire n_1168;
wire n_1216;
wire n_1943;
wire n_3228;
wire n_1320;
wire n_2716;
wire n_3249;
wire n_3081;
wire n_3657;
wire n_2452;
wire n_1430;
wire n_3650;
wire n_1316;
wire n_1287;
wire n_2722;
wire n_1452;
wire n_2854;
wire n_3672;
wire n_3010;
wire n_2499;
wire n_3533;
wire n_3043;
wire n_1622;
wire n_1586;
wire n_2543;
wire n_2264;
wire n_3464;
wire n_1694;
wire n_1535;
wire n_3137;
wire n_3382;
wire n_2486;
wire n_3132;
wire n_3560;
wire n_3723;
wire n_2571;
wire n_3138;
wire n_1596;
wire n_3177;
wire n_1190;
wire n_1734;
wire n_3172;
wire n_2902;
wire n_3217;
wire n_1983;
wire n_1938;
wire n_2498;
wire n_2220;
wire n_2577;
wire n_1262;
wire n_2472;
wire n_1891;
wire n_2171;
wire n_1213;
wire n_3238;
wire n_2235;
wire n_3529;
wire n_3570;
wire n_3394;
wire n_2988;
wire n_3136;
wire n_1350;
wire n_1673;
wire n_3828;
wire n_2232;
wire n_1715;
wire n_3536;
wire n_1443;
wire n_1272;
wire n_2392;
wire n_2894;
wire n_3424;
wire n_3957;
wire n_4038;
wire n_2790;
wire n_2037;
wire n_2808;
wire n_3710;
wire n_3784;
wire n_2298;
wire n_782;
wire n_2326;
wire n_1539;
wire n_490;
wire n_3594;
wire n_809;
wire n_1043;
wire n_3819;
wire n_4090;
wire n_3040;
wire n_1797;
wire n_3279;
wire n_1608;
wire n_986;
wire n_2305;
wire n_2120;
wire n_1472;
wire n_2050;
wire n_2373;
wire n_2164;
wire n_2402;
wire n_2225;
wire n_1081;
wire n_3628;
wire n_1870;
wire n_2964;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_2169;
wire n_3485;
wire n_4077;
wire n_2371;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_2006;
wire n_3402;
wire n_1491;
wire n_2187;
wire n_3501;
wire n_662;
wire n_3475;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_3905;
wire n_450;
wire n_3262;
wire n_3544;
wire n_2904;
wire n_4008;
wire n_2244;
wire n_3013;
wire n_3356;
wire n_2586;
wire n_1684;
wire n_921;
wire n_2446;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_2789;
wire n_3105;
wire n_3210;
wire n_2872;
wire n_937;
wire n_2257;
wire n_3692;
wire n_3845;
wire n_1682;
wire n_2017;
wire n_1695;
wire n_1828;
wire n_2046;
wire n_2272;
wire n_2699;
wire n_2200;
wire n_3029;
wire n_650;
wire n_3597;
wire n_1046;
wire n_2560;
wire n_1940;
wire n_1979;
wire n_2760;
wire n_2704;
wire n_3329;
wire n_1145;
wire n_1121;
wire n_1102;
wire n_1963;
wire n_2738;
wire n_972;
wire n_1405;
wire n_2376;
wire n_3826;
wire n_1406;
wire n_456;
wire n_3790;
wire n_3878;
wire n_2766;
wire n_1332;
wire n_2670;
wire n_2700;
wire n_624;
wire n_962;
wire n_1041;
wire n_2346;
wire n_565;
wire n_3134;
wire n_3647;
wire n_1569;
wire n_3681;
wire n_936;
wire n_3045;
wire n_3115;
wire n_1883;
wire n_3821;
wire n_1288;
wire n_3318;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_3278;
wire n_2342;
wire n_2167;
wire n_2084;
wire n_2970;
wire n_3676;
wire n_2882;
wire n_3666;
wire n_3675;
wire n_4017;
wire n_3320;
wire n_2541;
wire n_654;
wire n_2940;
wire n_2518;
wire n_2458;
wire n_1222;
wire n_599;
wire n_776;
wire n_1823;
wire n_2479;
wire n_3050;
wire n_3350;
wire n_2782;
wire n_3977;
wire n_1974;
wire n_3988;
wire n_2673;
wire n_2456;
wire n_1720;
wire n_3476;
wire n_2527;
wire n_482;
wire n_934;
wire n_2635;
wire n_1637;
wire n_3307;
wire n_3439;
wire n_1407;
wire n_1795;
wire n_2768;
wire n_3588;
wire n_2871;
wire n_2688;
wire n_1341;
wire n_1456;
wire n_1845;
wire n_3858;
wire n_1489;
wire n_2314;
wire n_3502;
wire n_942;
wire n_3003;
wire n_2798;
wire n_2852;
wire n_1524;
wire n_543;
wire n_2229;
wire n_1964;
wire n_2288;
wire n_1920;
wire n_2753;
wire n_2099;
wire n_1496;
wire n_1271;
wire n_3292;
wire n_1545;
wire n_2007;
wire n_3121;
wire n_2039;
wire n_3388;
wire n_1946;
wire n_1355;
wire n_1225;
wire n_3184;
wire n_1544;
wire n_2258;
wire n_1485;
wire n_1640;
wire n_4040;
wire n_804;
wire n_464;
wire n_1846;
wire n_3437;
wire n_3245;
wire n_3075;
wire n_2406;
wire n_533;
wire n_2390;
wire n_4007;
wire n_806;
wire n_3712;
wire n_879;
wire n_959;
wire n_2310;
wire n_2506;
wire n_584;
wire n_2141;
wire n_2562;
wire n_2642;
wire n_1343;
wire n_1522;
wire n_2734;
wire n_548;
wire n_1782;
wire n_2383;
wire n_2626;
wire n_1676;
wire n_833;
wire n_1830;
wire n_2351;
wire n_1567;
wire n_4037;
wire n_523;
wire n_1319;
wire n_707;
wire n_2986;
wire n_1900;
wire n_3930;
wire n_3246;
wire n_799;
wire n_1548;
wire n_3381;
wire n_3044;
wire n_3562;
wire n_2973;
wire n_1155;
wire n_2536;
wire n_3915;
wire n_2196;
wire n_2629;
wire n_3665;
wire n_1633;
wire n_2195;
wire n_3208;
wire n_2809;
wire n_3007;
wire n_787;
wire n_2172;
wire n_3528;
wire n_3489;
wire n_2835;
wire n_1416;
wire n_1528;
wire n_2820;
wire n_2293;
wire n_1146;
wire n_3698;
wire n_2021;
wire n_3355;
wire n_2454;
wire n_2114;
wire n_3074;
wire n_3174;
wire n_1086;
wire n_1066;
wire n_3102;
wire n_1948;
wire n_2125;
wire n_2026;
wire n_1282;
wire n_2561;
wire n_550;
wire n_3321;
wire n_2567;
wire n_2322;
wire n_652;
wire n_2154;
wire n_2727;
wire n_2962;
wire n_3377;
wire n_2939;
wire n_560;
wire n_1906;
wire n_1484;
wire n_2992;
wire n_3305;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_2533;
wire n_3157;
wire n_3530;
wire n_1758;
wire n_3221;
wire n_3267;
wire n_3752;
wire n_2283;
wire n_2869;
wire n_2422;
wire n_1925;
wire n_737;
wire n_1318;
wire n_1914;
wire n_1235;
wire n_3457;
wire n_1229;
wire n_2759;
wire n_3517;
wire n_2945;
wire n_3061;
wire n_3893;
wire n_2361;
wire n_1373;
wire n_1292;
wire n_3762;
wire n_3469;
wire n_3932;
wire n_2266;
wire n_2960;
wire n_3958;
wire n_3005;
wire n_3985;
wire n_2427;
wire n_3151;
wire n_3411;
wire n_1029;
wire n_3779;
wire n_1447;
wire n_2388;
wire n_3984;
wire n_2056;
wire n_790;
wire n_2611;
wire n_2901;
wire n_3258;
wire n_1706;
wire n_3389;
wire n_1498;
wire n_3143;
wire n_2653;
wire n_2417;
wire n_3000;
wire n_1210;
wire n_1248;
wire n_1556;
wire n_902;
wire n_2189;
wire n_2680;
wire n_4052;
wire n_2246;
wire n_1047;
wire n_3149;
wire n_3375;
wire n_3899;
wire n_4084;
wire n_3558;
wire n_1984;
wire n_3365;
wire n_2236;
wire n_1385;
wire n_3713;
wire n_3379;
wire n_3156;
wire n_459;
wire n_1269;
wire n_1931;
wire n_2083;
wire n_2834;
wire n_3207;
wire n_502;
wire n_2668;
wire n_672;
wire n_2441;
wire n_1257;
wire n_3008;
wire n_1751;
wire n_3401;
wire n_2840;
wire n_3197;
wire n_3242;
wire n_3939;
wire n_1375;
wire n_1941;
wire n_3483;
wire n_3613;
wire n_3972;
wire n_2128;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1962;
wire n_1236;
wire n_1794;
wire n_2398;
wire n_1725;
wire n_1928;
wire n_1559;
wire n_3855;
wire n_3743;
wire n_1872;
wire n_3091;
wire n_834;
wire n_2695;
wire n_4035;
wire n_3818;
wire n_743;
wire n_766;
wire n_3124;
wire n_1746;
wire n_1741;
wire n_1325;
wire n_1002;
wire n_4088;
wire n_1949;
wire n_3398;
wire n_3761;
wire n_3759;
wire n_545;
wire n_3524;
wire n_2671;
wire n_489;
wire n_2761;
wire n_2885;
wire n_2793;
wire n_2715;
wire n_2923;
wire n_1804;
wire n_2888;
wire n_3711;
wire n_3776;
wire n_1727;
wire n_2508;
wire n_1019;
wire n_636;
wire n_3511;
wire n_2054;
wire n_729;
wire n_876;
wire n_774;
wire n_3744;
wire n_3642;
wire n_2845;
wire n_1337;
wire n_3097;
wire n_660;
wire n_2062;
wire n_2041;
wire n_2975;
wire n_1477;
wire n_1360;
wire n_2839;
wire n_1860;
wire n_2856;
wire n_1904;
wire n_2874;
wire n_1200;
wire n_2070;
wire n_2588;
wire n_479;
wire n_3814;
wire n_1607;
wire n_3781;
wire n_1353;
wire n_1777;
wire n_1908;
wire n_1454;
wire n_2484;
wire n_2348;
wire n_2944;
wire n_2614;
wire n_2126;
wire n_3831;
wire n_869;
wire n_1154;
wire n_3308;
wire n_1113;
wire n_1600;
wire n_2833;
wire n_2253;
wire n_2758;
wire n_3843;
wire n_2366;
wire n_646;
wire n_528;
wire n_1098;
wire n_3694;
wire n_2937;
wire n_1329;
wire n_2045;
wire n_817;
wire n_2261;
wire n_3687;
wire n_2216;
wire n_3589;
wire n_2210;
wire n_3602;
wire n_897;
wire n_846;
wire n_3300;
wire n_2978;
wire n_2066;
wire n_3543;
wire n_841;
wire n_1476;
wire n_3621;
wire n_2516;
wire n_3391;
wire n_1001;
wire n_508;
wire n_1800;
wire n_2241;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_2903;
wire n_2827;
wire n_1177;
wire n_3216;
wire n_3458;
wire n_3515;
wire n_1150;
wire n_3808;
wire n_1742;
wire n_3190;
wire n_1562;
wire n_1690;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1882;
wire n_2951;
wire n_1076;
wire n_1118;
wire n_2949;
wire n_3726;
wire n_1007;
wire n_1929;
wire n_1807;
wire n_1378;
wire n_2369;
wire n_1592;
wire n_855;
wire n_1759;
wire n_2719;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_3758;
wire n_1879;
wire n_853;
wire n_440;
wire n_695;
wire n_3806;
wire n_4081;
wire n_1542;
wire n_2587;
wire n_3199;
wire n_2931;
wire n_875;
wire n_680;
wire n_3339;
wire n_1678;
wire n_2569;
wire n_661;
wire n_2400;
wire n_1716;
wire n_3866;
wire n_3787;
wire n_1256;
wire n_3585;
wire n_671;
wire n_3565;
wire n_1953;
wire n_933;
wire n_740;
wire n_703;
wire n_3343;
wire n_3303;
wire n_978;
wire n_2752;
wire n_3135;
wire n_1976;
wire n_2905;
wire n_1291;
wire n_1217;
wire n_3990;
wire n_751;
wire n_749;
wire n_3865;
wire n_1824;
wire n_3954;
wire n_1628;
wire n_4073;
wire n_1324;
wire n_3890;
wire n_1399;
wire n_2122;
wire n_2109;
wire n_3629;
wire n_1435;
wire n_3920;
wire n_969;
wire n_988;
wire n_2140;
wire n_3503;
wire n_3160;
wire n_1065;
wire n_2796;
wire n_3255;
wire n_2507;
wire n_1401;
wire n_2358;
wire n_1255;
wire n_568;
wire n_3658;
wire n_1516;
wire n_1536;
wire n_3846;
wire n_2186;
wire n_2163;
wire n_3512;
wire n_2029;
wire n_2815;
wire n_1204;
wire n_3951;
wire n_3034;
wire n_823;
wire n_1132;
wire n_643;
wire n_1074;
wire n_698;
wire n_1394;
wire n_3569;
wire n_1327;
wire n_1326;
wire n_955;
wire n_739;
wire n_3874;
wire n_1379;
wire n_2528;
wire n_2814;
wire n_2787;
wire n_1338;
wire n_1097;
wire n_2969;
wire n_2395;
wire n_935;
wire n_3027;
wire n_781;
wire n_789;
wire n_1554;
wire n_3231;
wire n_4083;
wire n_1130;
wire n_3083;
wire n_2979;
wire n_1810;
wire n_2953;
wire n_573;
wire n_769;
wire n_2380;
wire n_676;
wire n_1120;
wire n_832;
wire n_1583;
wire n_3049;
wire n_1730;
wire n_2295;
wire n_555;
wire n_814;
wire n_2746;
wire n_2946;
wire n_1643;
wire n_2020;
wire n_2500;
wire n_3430;
wire n_2269;
wire n_1729;
wire n_669;
wire n_2290;
wire n_2048;
wire n_3652;
wire n_3830;
wire n_3679;
wire n_2005;
wire n_747;
wire n_3541;
wire n_2565;
wire n_4023;
wire n_1389;
wire n_1105;
wire n_3117;
wire n_721;
wire n_1461;
wire n_742;
wire n_3432;
wire n_535;
wire n_691;
wire n_3617;
wire n_2076;
wire n_2736;
wire n_2883;
wire n_3583;
wire n_3860;
wire n_1408;
wire n_3851;
wire n_3567;
wire n_1196;
wire n_1598;
wire n_3493;
wire n_2935;
wire n_4046;
wire n_3807;
wire n_863;
wire n_3015;
wire n_2175;
wire n_601;
wire n_2182;
wire n_3774;
wire n_2910;
wire n_1283;
wire n_2385;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1785;
wire n_1147;
wire n_763;
wire n_1848;
wire n_1754;
wire n_2149;
wire n_3057;
wire n_3154;
wire n_3701;
wire n_2396;
wire n_1506;
wire n_2584;
wire n_1652;
wire n_1812;
wire n_957;
wire n_1994;
wire n_3473;
wire n_895;
wire n_866;
wire n_1227;
wire n_2485;
wire n_2450;
wire n_3739;
wire n_2284;
wire n_3898;
wire n_3520;
wire n_2566;
wire n_2287;
wire n_452;
wire n_744;
wire n_971;
wire n_2702;
wire n_3241;
wire n_946;
wire n_2906;
wire n_761;
wire n_1303;
wire n_2769;
wire n_3622;
wire n_1205;
wire n_2492;
wire n_1258;
wire n_3778;
wire n_4095;
wire n_2438;
wire n_2914;
wire n_1392;
wire n_1173;
wire n_1924;
wire n_525;
wire n_2463;
wire n_3363;
wire n_2881;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_3551;
wire n_3064;
wire n_1780;
wire n_3100;
wire n_3897;
wire n_3721;
wire n_1689;
wire n_2180;
wire n_3372;
wire n_2858;
wire n_3062;
wire n_2679;
wire n_1174;
wire n_3573;
wire n_1944;
wire n_1016;
wire n_1347;
wire n_4106;
wire n_795;
wire n_1501;
wire n_3604;
wire n_1221;
wire n_3334;
wire n_4027;
wire n_1245;
wire n_838;
wire n_3215;
wire n_3969;
wire n_3336;
wire n_647;
wire n_844;
wire n_448;
wire n_2952;
wire n_1017;
wire n_3068;
wire n_3853;
wire n_2117;
wire n_2234;
wire n_2779;
wire n_2685;
wire n_3823;
wire n_1083;
wire n_445;
wire n_3553;
wire n_1561;
wire n_2741;
wire n_3114;
wire n_930;
wire n_888;
wire n_2275;
wire n_1112;
wire n_2465;
wire n_2620;
wire n_2081;
wire n_2168;
wire n_2568;
wire n_2022;
wire n_1945;
wire n_2203;
wire n_910;
wire n_3811;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_2255;
wire n_2112;
wire n_1464;
wire n_653;
wire n_1737;
wire n_2430;
wire n_1414;
wire n_3486;
wire n_4086;
wire n_752;
wire n_908;
wire n_2649;
wire n_2721;
wire n_944;
wire n_3556;
wire n_2034;
wire n_576;
wire n_1028;
wire n_3836;
wire n_2106;
wire n_472;
wire n_2862;
wire n_2265;
wire n_2615;
wire n_2683;
wire n_1922;
wire n_563;
wire n_4068;
wire n_2032;
wire n_2744;
wire n_1011;
wire n_2474;
wire n_3703;
wire n_1566;
wire n_1215;
wire n_2444;
wire n_2437;
wire n_839;
wire n_2743;
wire n_3962;
wire n_708;
wire n_1973;
wire n_3181;
wire n_2267;
wire n_3456;
wire n_3035;
wire n_668;
wire n_626;
wire n_990;
wire n_1821;
wire n_779;
wire n_1537;
wire n_1500;
wire n_2205;
wire n_3699;
wire n_3204;
wire n_1104;
wire n_854;
wire n_1058;
wire n_3378;
wire n_4025;
wire n_2312;
wire n_498;
wire n_3404;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_2242;
wire n_3362;
wire n_3745;
wire n_4059;
wire n_1509;
wire n_3328;
wire n_1693;
wire n_3641;
wire n_2934;
wire n_3667;
wire n_3290;
wire n_1109;
wire n_3523;
wire n_2222;
wire n_712;
wire n_3256;
wire n_1276;
wire n_3802;
wire n_3868;
wire n_3176;
wire n_3309;
wire n_3671;
wire n_2015;
wire n_2118;
wire n_2466;
wire n_2111;
wire n_3982;
wire n_2915;
wire n_2530;
wire n_1148;
wire n_2505;
wire n_2188;
wire n_1989;
wire n_1161;
wire n_2609;
wire n_1085;
wire n_2802;
wire n_3796;
wire n_2999;
wire n_3840;
wire n_2014;
wire n_2042;
wire n_1239;
wire n_3643;
wire n_3697;
wire n_771;
wire n_1584;
wire n_2425;
wire n_470;
wire n_475;
wire n_924;
wire n_3408;
wire n_3461;
wire n_1582;
wire n_492;
wire n_3680;
wire n_2318;
wire n_3286;
wire n_4012;
wire n_2408;
wire n_1149;
wire n_3170;
wire n_3513;
wire n_3468;
wire n_3690;
wire n_1184;
wire n_3645;
wire n_2483;
wire n_2950;
wire n_719;
wire n_1972;
wire n_3060;
wire n_3304;
wire n_3682;
wire n_2592;
wire n_3771;
wire n_1525;
wire n_3098;
wire n_3995;
wire n_4076;
wire n_2594;
wire n_455;
wire n_2666;
wire n_4105;
wire n_1585;
wire n_1851;
wire n_1799;
wire n_1090;
wire n_2147;
wire n_2564;
wire n_592;
wire n_1816;
wire n_4064;
wire n_2503;
wire n_2433;
wire n_1518;
wire n_4049;
wire n_829;
wire n_1362;
wire n_1156;
wire n_3123;
wire n_984;
wire n_2600;
wire n_3380;
wire n_1829;
wire n_503;
wire n_2035;
wire n_3508;
wire n_3024;
wire n_1450;
wire n_1638;
wire n_3422;
wire n_868;
wire n_3038;
wire n_570;
wire n_859;
wire n_2033;
wire n_3086;
wire n_735;
wire n_4104;
wire n_1789;
wire n_2531;
wire n_1770;
wire n_878;
wire n_620;
wire n_3285;
wire n_519;
wire n_2523;
wire n_469;
wire n_1218;
wire n_2413;
wire n_500;
wire n_3769;
wire n_1482;
wire n_3361;
wire n_981;
wire n_3596;
wire n_714;
wire n_3478;
wire n_3936;
wire n_1349;
wire n_4089;
wire n_1144;
wire n_2071;
wire n_3669;
wire n_3863;
wire n_3219;
wire n_2429;
wire n_3130;
wire n_3702;
wire n_985;
wire n_2233;
wire n_2440;
wire n_2723;
wire n_481;
wire n_3521;
wire n_3233;
wire n_997;
wire n_1710;
wire n_2800;
wire n_2161;
wire n_3496;
wire n_1301;
wire n_2805;
wire n_802;
wire n_561;
wire n_3310;
wire n_980;
wire n_2681;
wire n_1306;
wire n_3264;
wire n_2010;
wire n_2282;
wire n_1651;
wire n_1198;
wire n_3096;
wire n_2360;
wire n_3764;
wire n_2047;
wire n_4061;
wire n_2651;
wire n_2095;
wire n_3239;
wire n_1609;
wire n_2174;
wire n_3161;
wire n_2799;
wire n_4075;
wire n_3344;
wire n_2334;
wire n_3902;
wire n_4062;
wire n_3881;
wire n_3295;
wire n_3947;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1998;
wire n_3066;
wire n_3101;
wire n_2426;
wire n_2490;
wire n_2844;
wire n_1574;
wire n_3989;
wire n_756;
wire n_2478;
wire n_1619;
wire n_2303;
wire n_1981;
wire n_2285;
wire n_1606;
wire n_810;
wire n_4108;
wire n_1133;
wire n_635;
wire n_1194;
wire n_3374;
wire n_3786;
wire n_3841;
wire n_2742;
wire n_2640;
wire n_3695;
wire n_4051;
wire n_1051;
wire n_3976;
wire n_1552;
wire n_2918;
wire n_583;
wire n_3288;
wire n_1996;
wire n_3563;
wire n_3992;
wire n_2367;
wire n_3876;
wire n_2867;
wire n_3198;
wire n_1039;
wire n_1442;
wire n_3495;
wire n_2726;
wire n_1034;
wire n_2043;
wire n_1480;
wire n_3125;
wire n_1158;
wire n_2909;
wire n_2248;
wire n_754;
wire n_941;
wire n_3552;
wire n_975;
wire n_3206;
wire n_1031;
wire n_1305;
wire n_2363;
wire n_2578;
wire n_553;
wire n_849;
wire n_2662;
wire n_3116;
wire n_3147;
wire n_3383;
wire n_3709;
wire n_753;
wire n_3925;
wire n_4091;
wire n_1753;
wire n_3095;
wire n_3180;
wire n_3738;
wire n_3359;
wire n_2795;
wire n_3472;
wire n_2471;
wire n_467;
wire n_3187;
wire n_2540;
wire n_973;
wire n_2807;
wire n_1921;
wire n_3218;
wire n_3610;
wire n_3618;
wire n_3330;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_2217;
wire n_2197;
wire n_582;
wire n_2065;
wire n_2879;
wire n_861;
wire n_3717;
wire n_857;
wire n_967;
wire n_571;
wire n_2215;
wire n_2461;
wire n_2001;
wire n_2107;
wire n_1884;
wire n_2040;
wire n_679;
wire n_4057;
wire n_2968;
wire n_633;
wire n_1170;
wire n_665;
wire n_2221;
wire n_1629;
wire n_588;
wire n_1260;
wire n_1819;
wire n_2055;
wire n_3555;
wire n_1010;
wire n_3444;
wire n_2553;
wire n_1040;
wire n_915;
wire n_632;
wire n_3059;
wire n_1166;
wire n_2038;
wire n_812;
wire n_2891;
wire n_1131;
wire n_2634;
wire n_1761;
wire n_2709;
wire n_3155;
wire n_3445;
wire n_534;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_3110;
wire n_1890;
wire n_1632;
wire n_3017;
wire n_3955;
wire n_1805;
wire n_2477;
wire n_1557;
wire n_1888;
wire n_2280;
wire n_1833;
wire n_3903;
wire n_730;
wire n_1311;
wire n_3945;
wire n_1494;
wire n_2325;
wire n_670;
wire n_1850;
wire n_1898;
wire n_2443;
wire n_2697;
wire n_3235;
wire n_3854;
wire n_2308;
wire n_2162;
wire n_3908;
wire n_1868;
wire n_2333;
wire n_2079;
wire n_3467;
wire n_3001;
wire n_3587;
wire n_1089;
wire n_1887;
wire n_1587;
wire n_3916;
wire n_3527;
wire n_3795;
wire n_2512;
wire n_3950;
wire n_3433;
wire n_3852;
wire n_1365;
wire n_1417;
wire n_1242;
wire n_2086;
wire n_2185;
wire n_2927;
wire n_3673;
wire n_1836;
wire n_3833;
wire n_3896;
wire n_2774;
wire n_3815;
wire n_3039;
wire n_681;
wire n_1226;
wire n_3740;
wire n_3162;
wire n_1274;
wire n_1486;
wire n_2166;
wire n_3094;
wire n_2899;
wire n_3333;
wire n_3274;
wire n_3186;
wire n_640;
wire n_1322;
wire n_965;
wire n_1899;
wire n_1428;
wire n_4093;
wire n_1616;
wire n_1576;
wire n_1862;
wire n_1856;
wire n_1958;
wire n_2077;
wire n_784;
wire n_1059;
wire n_1197;
wire n_3065;
wire n_3965;
wire n_2632;
wire n_2579;
wire n_722;
wire n_862;
wire n_2105;
wire n_3079;
wire n_2098;
wire n_3085;
wire n_540;
wire n_1423;
wire n_2813;
wire n_1935;
wire n_3584;
wire n_4039;
wire n_3387;
wire n_2027;
wire n_457;
wire n_3070;
wire n_3800;
wire n_2223;
wire n_2091;
wire n_3263;
wire n_3431;
wire n_3420;
wire n_2991;
wire n_1915;
wire n_629;
wire n_1621;
wire n_1748;
wire n_2547;
wire n_2415;
wire n_900;
wire n_3504;
wire n_1449;
wire n_531;
wire n_827;
wire n_2912;
wire n_2659;
wire n_2930;
wire n_1025;
wire n_3409;
wire n_2419;
wire n_3111;
wire n_2116;
wire n_2320;
wire n_1885;
wire n_2677;
wire n_1013;
wire n_3182;
wire n_1259;
wire n_3054;
wire n_3283;
wire n_2183;
wire n_3002;
wire n_1538;
wire n_649;
wire n_4030;
wire n_1612;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_87),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_384),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_121),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_277),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_438),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_38),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_218),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_108),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_399),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_58),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_7),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_134),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_266),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_145),
.Y(n_453)
);

CKINVDCx20_ASAP7_75t_R g454 ( 
.A(n_368),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_373),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_46),
.Y(n_456)
);

INVxp67_ASAP7_75t_L g457 ( 
.A(n_57),
.Y(n_457)
);

INVx2_ASAP7_75t_L g458 ( 
.A(n_136),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_64),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_184),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_97),
.Y(n_461)
);

BUFx3_ASAP7_75t_L g462 ( 
.A(n_253),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_89),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_309),
.Y(n_464)
);

CKINVDCx5p33_ASAP7_75t_R g465 ( 
.A(n_100),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_287),
.Y(n_466)
);

CKINVDCx5p33_ASAP7_75t_R g467 ( 
.A(n_37),
.Y(n_467)
);

CKINVDCx20_ASAP7_75t_R g468 ( 
.A(n_281),
.Y(n_468)
);

CKINVDCx5p33_ASAP7_75t_R g469 ( 
.A(n_415),
.Y(n_469)
);

CKINVDCx5p33_ASAP7_75t_R g470 ( 
.A(n_285),
.Y(n_470)
);

CKINVDCx5p33_ASAP7_75t_R g471 ( 
.A(n_70),
.Y(n_471)
);

INVx2_ASAP7_75t_L g472 ( 
.A(n_197),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_225),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_419),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_244),
.Y(n_475)
);

CKINVDCx5p33_ASAP7_75t_R g476 ( 
.A(n_82),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_333),
.Y(n_477)
);

INVx2_ASAP7_75t_L g478 ( 
.A(n_349),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_248),
.Y(n_479)
);

INVx1_ASAP7_75t_SL g480 ( 
.A(n_79),
.Y(n_480)
);

CKINVDCx5p33_ASAP7_75t_R g481 ( 
.A(n_356),
.Y(n_481)
);

INVx2_ASAP7_75t_L g482 ( 
.A(n_351),
.Y(n_482)
);

CKINVDCx5p33_ASAP7_75t_R g483 ( 
.A(n_345),
.Y(n_483)
);

CKINVDCx20_ASAP7_75t_R g484 ( 
.A(n_37),
.Y(n_484)
);

CKINVDCx5p33_ASAP7_75t_R g485 ( 
.A(n_208),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_305),
.Y(n_486)
);

INVx2_ASAP7_75t_L g487 ( 
.A(n_210),
.Y(n_487)
);

CKINVDCx5p33_ASAP7_75t_R g488 ( 
.A(n_63),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_420),
.Y(n_489)
);

HB1xp67_ASAP7_75t_L g490 ( 
.A(n_97),
.Y(n_490)
);

CKINVDCx5p33_ASAP7_75t_R g491 ( 
.A(n_234),
.Y(n_491)
);

CKINVDCx5p33_ASAP7_75t_R g492 ( 
.A(n_126),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_203),
.Y(n_493)
);

CKINVDCx5p33_ASAP7_75t_R g494 ( 
.A(n_217),
.Y(n_494)
);

INVxp67_ASAP7_75t_L g495 ( 
.A(n_204),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_240),
.Y(n_496)
);

CKINVDCx5p33_ASAP7_75t_R g497 ( 
.A(n_171),
.Y(n_497)
);

BUFx2_ASAP7_75t_SL g498 ( 
.A(n_385),
.Y(n_498)
);

INVx2_ASAP7_75t_L g499 ( 
.A(n_65),
.Y(n_499)
);

CKINVDCx5p33_ASAP7_75t_R g500 ( 
.A(n_343),
.Y(n_500)
);

CKINVDCx5p33_ASAP7_75t_R g501 ( 
.A(n_134),
.Y(n_501)
);

CKINVDCx20_ASAP7_75t_R g502 ( 
.A(n_20),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_426),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_50),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_138),
.Y(n_505)
);

CKINVDCx5p33_ASAP7_75t_R g506 ( 
.A(n_353),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_405),
.Y(n_507)
);

CKINVDCx5p33_ASAP7_75t_R g508 ( 
.A(n_1),
.Y(n_508)
);

CKINVDCx5p33_ASAP7_75t_R g509 ( 
.A(n_228),
.Y(n_509)
);

CKINVDCx5p33_ASAP7_75t_R g510 ( 
.A(n_403),
.Y(n_510)
);

CKINVDCx5p33_ASAP7_75t_R g511 ( 
.A(n_212),
.Y(n_511)
);

INVx1_ASAP7_75t_SL g512 ( 
.A(n_47),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_360),
.Y(n_513)
);

CKINVDCx5p33_ASAP7_75t_R g514 ( 
.A(n_131),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_409),
.Y(n_515)
);

CKINVDCx5p33_ASAP7_75t_R g516 ( 
.A(n_269),
.Y(n_516)
);

CKINVDCx5p33_ASAP7_75t_R g517 ( 
.A(n_33),
.Y(n_517)
);

CKINVDCx5p33_ASAP7_75t_R g518 ( 
.A(n_40),
.Y(n_518)
);

CKINVDCx5p33_ASAP7_75t_R g519 ( 
.A(n_9),
.Y(n_519)
);

BUFx3_ASAP7_75t_L g520 ( 
.A(n_142),
.Y(n_520)
);

CKINVDCx20_ASAP7_75t_R g521 ( 
.A(n_0),
.Y(n_521)
);

CKINVDCx5p33_ASAP7_75t_R g522 ( 
.A(n_339),
.Y(n_522)
);

BUFx8_ASAP7_75t_SL g523 ( 
.A(n_85),
.Y(n_523)
);

BUFx2_ASAP7_75t_L g524 ( 
.A(n_227),
.Y(n_524)
);

CKINVDCx5p33_ASAP7_75t_R g525 ( 
.A(n_393),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_74),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_65),
.Y(n_527)
);

CKINVDCx5p33_ASAP7_75t_R g528 ( 
.A(n_253),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_231),
.Y(n_529)
);

HB1xp67_ASAP7_75t_L g530 ( 
.A(n_143),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_81),
.Y(n_531)
);

CKINVDCx5p33_ASAP7_75t_R g532 ( 
.A(n_281),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_113),
.Y(n_533)
);

CKINVDCx20_ASAP7_75t_R g534 ( 
.A(n_363),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_124),
.Y(n_535)
);

INVx1_ASAP7_75t_SL g536 ( 
.A(n_32),
.Y(n_536)
);

CKINVDCx5p33_ASAP7_75t_R g537 ( 
.A(n_433),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_303),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_35),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_357),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_20),
.Y(n_541)
);

INVx2_ASAP7_75t_SL g542 ( 
.A(n_254),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_151),
.Y(n_543)
);

BUFx6f_ASAP7_75t_L g544 ( 
.A(n_408),
.Y(n_544)
);

CKINVDCx5p33_ASAP7_75t_R g545 ( 
.A(n_247),
.Y(n_545)
);

CKINVDCx5p33_ASAP7_75t_R g546 ( 
.A(n_352),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_323),
.Y(n_547)
);

CKINVDCx5p33_ASAP7_75t_R g548 ( 
.A(n_181),
.Y(n_548)
);

CKINVDCx5p33_ASAP7_75t_R g549 ( 
.A(n_3),
.Y(n_549)
);

CKINVDCx5p33_ASAP7_75t_R g550 ( 
.A(n_298),
.Y(n_550)
);

BUFx5_ASAP7_75t_L g551 ( 
.A(n_230),
.Y(n_551)
);

CKINVDCx5p33_ASAP7_75t_R g552 ( 
.A(n_246),
.Y(n_552)
);

CKINVDCx5p33_ASAP7_75t_R g553 ( 
.A(n_96),
.Y(n_553)
);

CKINVDCx16_ASAP7_75t_R g554 ( 
.A(n_354),
.Y(n_554)
);

INVx2_ASAP7_75t_L g555 ( 
.A(n_189),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_27),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_249),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_66),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_33),
.Y(n_559)
);

CKINVDCx5p33_ASAP7_75t_R g560 ( 
.A(n_250),
.Y(n_560)
);

CKINVDCx5p33_ASAP7_75t_R g561 ( 
.A(n_152),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_387),
.Y(n_562)
);

BUFx10_ASAP7_75t_L g563 ( 
.A(n_194),
.Y(n_563)
);

INVxp33_ASAP7_75t_L g564 ( 
.A(n_225),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_133),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_177),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_51),
.Y(n_567)
);

CKINVDCx5p33_ASAP7_75t_R g568 ( 
.A(n_36),
.Y(n_568)
);

CKINVDCx5p33_ASAP7_75t_R g569 ( 
.A(n_198),
.Y(n_569)
);

CKINVDCx5p33_ASAP7_75t_R g570 ( 
.A(n_95),
.Y(n_570)
);

CKINVDCx5p33_ASAP7_75t_R g571 ( 
.A(n_258),
.Y(n_571)
);

CKINVDCx5p33_ASAP7_75t_R g572 ( 
.A(n_210),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_308),
.Y(n_573)
);

CKINVDCx5p33_ASAP7_75t_R g574 ( 
.A(n_80),
.Y(n_574)
);

CKINVDCx20_ASAP7_75t_R g575 ( 
.A(n_248),
.Y(n_575)
);

CKINVDCx5p33_ASAP7_75t_R g576 ( 
.A(n_4),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_230),
.Y(n_577)
);

BUFx6f_ASAP7_75t_L g578 ( 
.A(n_427),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_310),
.Y(n_579)
);

CKINVDCx5p33_ASAP7_75t_R g580 ( 
.A(n_171),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_263),
.Y(n_581)
);

INVx1_ASAP7_75t_SL g582 ( 
.A(n_289),
.Y(n_582)
);

CKINVDCx5p33_ASAP7_75t_R g583 ( 
.A(n_377),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_355),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_197),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_383),
.Y(n_586)
);

CKINVDCx5p33_ASAP7_75t_R g587 ( 
.A(n_199),
.Y(n_587)
);

CKINVDCx5p33_ASAP7_75t_R g588 ( 
.A(n_300),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_257),
.Y(n_589)
);

CKINVDCx5p33_ASAP7_75t_R g590 ( 
.A(n_47),
.Y(n_590)
);

CKINVDCx20_ASAP7_75t_R g591 ( 
.A(n_250),
.Y(n_591)
);

BUFx2_ASAP7_75t_L g592 ( 
.A(n_51),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_259),
.Y(n_593)
);

HB1xp67_ASAP7_75t_L g594 ( 
.A(n_185),
.Y(n_594)
);

CKINVDCx5p33_ASAP7_75t_R g595 ( 
.A(n_193),
.Y(n_595)
);

CKINVDCx5p33_ASAP7_75t_R g596 ( 
.A(n_74),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_71),
.Y(n_597)
);

CKINVDCx5p33_ASAP7_75t_R g598 ( 
.A(n_154),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_201),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_264),
.Y(n_600)
);

CKINVDCx5p33_ASAP7_75t_R g601 ( 
.A(n_336),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_156),
.Y(n_602)
);

CKINVDCx5p33_ASAP7_75t_R g603 ( 
.A(n_71),
.Y(n_603)
);

CKINVDCx5p33_ASAP7_75t_R g604 ( 
.A(n_390),
.Y(n_604)
);

BUFx6f_ASAP7_75t_L g605 ( 
.A(n_169),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_311),
.Y(n_606)
);

CKINVDCx5p33_ASAP7_75t_R g607 ( 
.A(n_114),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_338),
.Y(n_608)
);

CKINVDCx5p33_ASAP7_75t_R g609 ( 
.A(n_79),
.Y(n_609)
);

INVx2_ASAP7_75t_L g610 ( 
.A(n_263),
.Y(n_610)
);

CKINVDCx5p33_ASAP7_75t_R g611 ( 
.A(n_278),
.Y(n_611)
);

CKINVDCx5p33_ASAP7_75t_R g612 ( 
.A(n_138),
.Y(n_612)
);

CKINVDCx5p33_ASAP7_75t_R g613 ( 
.A(n_364),
.Y(n_613)
);

CKINVDCx5p33_ASAP7_75t_R g614 ( 
.A(n_100),
.Y(n_614)
);

INVx2_ASAP7_75t_L g615 ( 
.A(n_229),
.Y(n_615)
);

CKINVDCx14_ASAP7_75t_R g616 ( 
.A(n_60),
.Y(n_616)
);

CKINVDCx20_ASAP7_75t_R g617 ( 
.A(n_176),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_365),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_192),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_324),
.Y(n_620)
);

CKINVDCx5p33_ASAP7_75t_R g621 ( 
.A(n_425),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_41),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_147),
.Y(n_623)
);

CKINVDCx5p33_ASAP7_75t_R g624 ( 
.A(n_181),
.Y(n_624)
);

CKINVDCx5p33_ASAP7_75t_R g625 ( 
.A(n_340),
.Y(n_625)
);

CKINVDCx5p33_ASAP7_75t_R g626 ( 
.A(n_193),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_44),
.Y(n_627)
);

INVx1_ASAP7_75t_SL g628 ( 
.A(n_54),
.Y(n_628)
);

INVx1_ASAP7_75t_SL g629 ( 
.A(n_423),
.Y(n_629)
);

CKINVDCx5p33_ASAP7_75t_R g630 ( 
.A(n_379),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_227),
.Y(n_631)
);

CKINVDCx20_ASAP7_75t_R g632 ( 
.A(n_412),
.Y(n_632)
);

CKINVDCx5p33_ASAP7_75t_R g633 ( 
.A(n_158),
.Y(n_633)
);

BUFx10_ASAP7_75t_L g634 ( 
.A(n_388),
.Y(n_634)
);

CKINVDCx5p33_ASAP7_75t_R g635 ( 
.A(n_198),
.Y(n_635)
);

CKINVDCx5p33_ASAP7_75t_R g636 ( 
.A(n_107),
.Y(n_636)
);

CKINVDCx5p33_ASAP7_75t_R g637 ( 
.A(n_366),
.Y(n_637)
);

CKINVDCx5p33_ASAP7_75t_R g638 ( 
.A(n_327),
.Y(n_638)
);

CKINVDCx5p33_ASAP7_75t_R g639 ( 
.A(n_177),
.Y(n_639)
);

CKINVDCx16_ASAP7_75t_R g640 ( 
.A(n_367),
.Y(n_640)
);

CKINVDCx5p33_ASAP7_75t_R g641 ( 
.A(n_188),
.Y(n_641)
);

CKINVDCx5p33_ASAP7_75t_R g642 ( 
.A(n_191),
.Y(n_642)
);

CKINVDCx5p33_ASAP7_75t_R g643 ( 
.A(n_294),
.Y(n_643)
);

CKINVDCx5p33_ASAP7_75t_R g644 ( 
.A(n_150),
.Y(n_644)
);

CKINVDCx16_ASAP7_75t_R g645 ( 
.A(n_28),
.Y(n_645)
);

CKINVDCx20_ASAP7_75t_R g646 ( 
.A(n_124),
.Y(n_646)
);

CKINVDCx5p33_ASAP7_75t_R g647 ( 
.A(n_38),
.Y(n_647)
);

CKINVDCx5p33_ASAP7_75t_R g648 ( 
.A(n_371),
.Y(n_648)
);

CKINVDCx5p33_ASAP7_75t_R g649 ( 
.A(n_61),
.Y(n_649)
);

CKINVDCx5p33_ASAP7_75t_R g650 ( 
.A(n_218),
.Y(n_650)
);

CKINVDCx5p33_ASAP7_75t_R g651 ( 
.A(n_267),
.Y(n_651)
);

CKINVDCx5p33_ASAP7_75t_R g652 ( 
.A(n_199),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_429),
.Y(n_653)
);

INVx2_ASAP7_75t_SL g654 ( 
.A(n_278),
.Y(n_654)
);

CKINVDCx5p33_ASAP7_75t_R g655 ( 
.A(n_165),
.Y(n_655)
);

CKINVDCx5p33_ASAP7_75t_R g656 ( 
.A(n_350),
.Y(n_656)
);

CKINVDCx5p33_ASAP7_75t_R g657 ( 
.A(n_139),
.Y(n_657)
);

CKINVDCx5p33_ASAP7_75t_R g658 ( 
.A(n_369),
.Y(n_658)
);

INVx2_ASAP7_75t_L g659 ( 
.A(n_292),
.Y(n_659)
);

INVxp67_ASAP7_75t_L g660 ( 
.A(n_361),
.Y(n_660)
);

CKINVDCx5p33_ASAP7_75t_R g661 ( 
.A(n_208),
.Y(n_661)
);

CKINVDCx5p33_ASAP7_75t_R g662 ( 
.A(n_191),
.Y(n_662)
);

CKINVDCx20_ASAP7_75t_R g663 ( 
.A(n_277),
.Y(n_663)
);

CKINVDCx20_ASAP7_75t_R g664 ( 
.A(n_7),
.Y(n_664)
);

CKINVDCx5p33_ASAP7_75t_R g665 ( 
.A(n_179),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_154),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_116),
.Y(n_667)
);

BUFx6f_ASAP7_75t_L g668 ( 
.A(n_243),
.Y(n_668)
);

CKINVDCx5p33_ASAP7_75t_R g669 ( 
.A(n_348),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_62),
.Y(n_670)
);

BUFx3_ASAP7_75t_L g671 ( 
.A(n_56),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_83),
.Y(n_672)
);

HB1xp67_ASAP7_75t_L g673 ( 
.A(n_54),
.Y(n_673)
);

CKINVDCx5p33_ASAP7_75t_R g674 ( 
.A(n_70),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_260),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_258),
.Y(n_676)
);

CKINVDCx5p33_ASAP7_75t_R g677 ( 
.A(n_81),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_5),
.Y(n_678)
);

INVx1_ASAP7_75t_SL g679 ( 
.A(n_109),
.Y(n_679)
);

INVx1_ASAP7_75t_SL g680 ( 
.A(n_422),
.Y(n_680)
);

CKINVDCx5p33_ASAP7_75t_R g681 ( 
.A(n_184),
.Y(n_681)
);

CKINVDCx5p33_ASAP7_75t_R g682 ( 
.A(n_46),
.Y(n_682)
);

INVx2_ASAP7_75t_SL g683 ( 
.A(n_320),
.Y(n_683)
);

CKINVDCx5p33_ASAP7_75t_R g684 ( 
.A(n_26),
.Y(n_684)
);

INVxp67_ASAP7_75t_L g685 ( 
.A(n_418),
.Y(n_685)
);

CKINVDCx5p33_ASAP7_75t_R g686 ( 
.A(n_386),
.Y(n_686)
);

CKINVDCx5p33_ASAP7_75t_R g687 ( 
.A(n_275),
.Y(n_687)
);

INVx2_ASAP7_75t_L g688 ( 
.A(n_404),
.Y(n_688)
);

CKINVDCx5p33_ASAP7_75t_R g689 ( 
.A(n_347),
.Y(n_689)
);

INVx2_ASAP7_75t_L g690 ( 
.A(n_407),
.Y(n_690)
);

INVx2_ASAP7_75t_SL g691 ( 
.A(n_216),
.Y(n_691)
);

CKINVDCx20_ASAP7_75t_R g692 ( 
.A(n_173),
.Y(n_692)
);

CKINVDCx5p33_ASAP7_75t_R g693 ( 
.A(n_9),
.Y(n_693)
);

CKINVDCx5p33_ASAP7_75t_R g694 ( 
.A(n_35),
.Y(n_694)
);

CKINVDCx5p33_ASAP7_75t_R g695 ( 
.A(n_205),
.Y(n_695)
);

CKINVDCx5p33_ASAP7_75t_R g696 ( 
.A(n_18),
.Y(n_696)
);

CKINVDCx5p33_ASAP7_75t_R g697 ( 
.A(n_40),
.Y(n_697)
);

CKINVDCx5p33_ASAP7_75t_R g698 ( 
.A(n_304),
.Y(n_698)
);

INVx2_ASAP7_75t_L g699 ( 
.A(n_16),
.Y(n_699)
);

CKINVDCx5p33_ASAP7_75t_R g700 ( 
.A(n_96),
.Y(n_700)
);

BUFx3_ASAP7_75t_L g701 ( 
.A(n_172),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_19),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_273),
.Y(n_703)
);

CKINVDCx5p33_ASAP7_75t_R g704 ( 
.A(n_243),
.Y(n_704)
);

HB1xp67_ASAP7_75t_L g705 ( 
.A(n_163),
.Y(n_705)
);

CKINVDCx5p33_ASAP7_75t_R g706 ( 
.A(n_328),
.Y(n_706)
);

CKINVDCx5p33_ASAP7_75t_R g707 ( 
.A(n_274),
.Y(n_707)
);

CKINVDCx5p33_ASAP7_75t_R g708 ( 
.A(n_389),
.Y(n_708)
);

CKINVDCx20_ASAP7_75t_R g709 ( 
.A(n_155),
.Y(n_709)
);

CKINVDCx5p33_ASAP7_75t_R g710 ( 
.A(n_380),
.Y(n_710)
);

CKINVDCx5p33_ASAP7_75t_R g711 ( 
.A(n_52),
.Y(n_711)
);

CKINVDCx20_ASAP7_75t_R g712 ( 
.A(n_92),
.Y(n_712)
);

INVxp67_ASAP7_75t_L g713 ( 
.A(n_395),
.Y(n_713)
);

CKINVDCx5p33_ASAP7_75t_R g714 ( 
.A(n_187),
.Y(n_714)
);

CKINVDCx5p33_ASAP7_75t_R g715 ( 
.A(n_411),
.Y(n_715)
);

CKINVDCx20_ASAP7_75t_R g716 ( 
.A(n_270),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_101),
.Y(n_717)
);

BUFx6f_ASAP7_75t_L g718 ( 
.A(n_106),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_89),
.Y(n_719)
);

CKINVDCx20_ASAP7_75t_R g720 ( 
.A(n_431),
.Y(n_720)
);

BUFx3_ASAP7_75t_L g721 ( 
.A(n_127),
.Y(n_721)
);

CKINVDCx20_ASAP7_75t_R g722 ( 
.A(n_42),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_301),
.Y(n_723)
);

CKINVDCx5p33_ASAP7_75t_R g724 ( 
.A(n_148),
.Y(n_724)
);

BUFx2_ASAP7_75t_L g725 ( 
.A(n_13),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_432),
.Y(n_726)
);

INVx1_ASAP7_75t_SL g727 ( 
.A(n_101),
.Y(n_727)
);

CKINVDCx5p33_ASAP7_75t_R g728 ( 
.A(n_378),
.Y(n_728)
);

CKINVDCx5p33_ASAP7_75t_R g729 ( 
.A(n_288),
.Y(n_729)
);

INVx2_ASAP7_75t_L g730 ( 
.A(n_108),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_43),
.Y(n_731)
);

CKINVDCx5p33_ASAP7_75t_R g732 ( 
.A(n_73),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_247),
.Y(n_733)
);

CKINVDCx5p33_ASAP7_75t_R g734 ( 
.A(n_117),
.Y(n_734)
);

CKINVDCx5p33_ASAP7_75t_R g735 ( 
.A(n_143),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_205),
.Y(n_736)
);

CKINVDCx5p33_ASAP7_75t_R g737 ( 
.A(n_115),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_185),
.Y(n_738)
);

CKINVDCx5p33_ASAP7_75t_R g739 ( 
.A(n_83),
.Y(n_739)
);

INVx2_ASAP7_75t_L g740 ( 
.A(n_358),
.Y(n_740)
);

CKINVDCx20_ASAP7_75t_R g741 ( 
.A(n_90),
.Y(n_741)
);

BUFx6f_ASAP7_75t_L g742 ( 
.A(n_254),
.Y(n_742)
);

CKINVDCx5p33_ASAP7_75t_R g743 ( 
.A(n_148),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_249),
.Y(n_744)
);

BUFx10_ASAP7_75t_L g745 ( 
.A(n_77),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_113),
.Y(n_746)
);

CKINVDCx5p33_ASAP7_75t_R g747 ( 
.A(n_240),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_14),
.Y(n_748)
);

CKINVDCx5p33_ASAP7_75t_R g749 ( 
.A(n_117),
.Y(n_749)
);

CKINVDCx5p33_ASAP7_75t_R g750 ( 
.A(n_82),
.Y(n_750)
);

CKINVDCx5p33_ASAP7_75t_R g751 ( 
.A(n_213),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_400),
.Y(n_752)
);

CKINVDCx5p33_ASAP7_75t_R g753 ( 
.A(n_76),
.Y(n_753)
);

CKINVDCx5p33_ASAP7_75t_R g754 ( 
.A(n_13),
.Y(n_754)
);

INVx2_ASAP7_75t_SL g755 ( 
.A(n_192),
.Y(n_755)
);

CKINVDCx5p33_ASAP7_75t_R g756 ( 
.A(n_428),
.Y(n_756)
);

BUFx6f_ASAP7_75t_L g757 ( 
.A(n_222),
.Y(n_757)
);

CKINVDCx20_ASAP7_75t_R g758 ( 
.A(n_286),
.Y(n_758)
);

CKINVDCx5p33_ASAP7_75t_R g759 ( 
.A(n_325),
.Y(n_759)
);

CKINVDCx20_ASAP7_75t_R g760 ( 
.A(n_44),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_392),
.Y(n_761)
);

INVx1_ASAP7_75t_SL g762 ( 
.A(n_374),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_58),
.Y(n_763)
);

INVxp67_ASAP7_75t_L g764 ( 
.A(n_295),
.Y(n_764)
);

CKINVDCx5p33_ASAP7_75t_R g765 ( 
.A(n_159),
.Y(n_765)
);

CKINVDCx5p33_ASAP7_75t_R g766 ( 
.A(n_75),
.Y(n_766)
);

CKINVDCx5p33_ASAP7_75t_R g767 ( 
.A(n_187),
.Y(n_767)
);

CKINVDCx5p33_ASAP7_75t_R g768 ( 
.A(n_92),
.Y(n_768)
);

INVx1_ASAP7_75t_SL g769 ( 
.A(n_342),
.Y(n_769)
);

CKINVDCx5p33_ASAP7_75t_R g770 ( 
.A(n_282),
.Y(n_770)
);

CKINVDCx20_ASAP7_75t_R g771 ( 
.A(n_454),
.Y(n_771)
);

CKINVDCx14_ASAP7_75t_R g772 ( 
.A(n_616),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_551),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_551),
.Y(n_774)
);

BUFx2_ASAP7_75t_L g775 ( 
.A(n_524),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_551),
.Y(n_776)
);

CKINVDCx5p33_ASAP7_75t_R g777 ( 
.A(n_523),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_551),
.Y(n_778)
);

CKINVDCx5p33_ASAP7_75t_R g779 ( 
.A(n_645),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_551),
.Y(n_780)
);

INVxp67_ASAP7_75t_SL g781 ( 
.A(n_605),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_551),
.Y(n_782)
);

INVx1_ASAP7_75t_SL g783 ( 
.A(n_524),
.Y(n_783)
);

BUFx6f_ASAP7_75t_L g784 ( 
.A(n_544),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_551),
.Y(n_785)
);

CKINVDCx5p33_ASAP7_75t_R g786 ( 
.A(n_645),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_551),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_551),
.Y(n_788)
);

BUFx3_ASAP7_75t_L g789 ( 
.A(n_634),
.Y(n_789)
);

CKINVDCx5p33_ASAP7_75t_R g790 ( 
.A(n_440),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_464),
.Y(n_791)
);

CKINVDCx5p33_ASAP7_75t_R g792 ( 
.A(n_442),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_464),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_466),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_466),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_474),
.Y(n_796)
);

INVx2_ASAP7_75t_SL g797 ( 
.A(n_462),
.Y(n_797)
);

BUFx8_ASAP7_75t_SL g798 ( 
.A(n_592),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_474),
.Y(n_799)
);

INVx2_ASAP7_75t_L g800 ( 
.A(n_605),
.Y(n_800)
);

CKINVDCx20_ASAP7_75t_R g801 ( 
.A(n_534),
.Y(n_801)
);

INVx2_ASAP7_75t_L g802 ( 
.A(n_605),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_477),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_477),
.Y(n_804)
);

CKINVDCx5p33_ASAP7_75t_R g805 ( 
.A(n_443),
.Y(n_805)
);

CKINVDCx5p33_ASAP7_75t_R g806 ( 
.A(n_445),
.Y(n_806)
);

CKINVDCx5p33_ASAP7_75t_R g807 ( 
.A(n_446),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_486),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_486),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_489),
.Y(n_810)
);

BUFx2_ASAP7_75t_SL g811 ( 
.A(n_683),
.Y(n_811)
);

INVxp33_ASAP7_75t_L g812 ( 
.A(n_490),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_489),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_503),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_503),
.Y(n_815)
);

CKINVDCx16_ASAP7_75t_R g816 ( 
.A(n_554),
.Y(n_816)
);

OR2x2_ASAP7_75t_L g817 ( 
.A(n_450),
.B(n_453),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_507),
.Y(n_818)
);

CKINVDCx5p33_ASAP7_75t_R g819 ( 
.A(n_447),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_507),
.Y(n_820)
);

NOR2xp33_ASAP7_75t_L g821 ( 
.A(n_683),
.B(n_0),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_513),
.Y(n_822)
);

CKINVDCx14_ASAP7_75t_R g823 ( 
.A(n_592),
.Y(n_823)
);

BUFx2_ASAP7_75t_L g824 ( 
.A(n_725),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_513),
.Y(n_825)
);

INVx2_ASAP7_75t_L g826 ( 
.A(n_605),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_515),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_515),
.Y(n_828)
);

INVx1_ASAP7_75t_SL g829 ( 
.A(n_725),
.Y(n_829)
);

INVx1_ASAP7_75t_SL g830 ( 
.A(n_468),
.Y(n_830)
);

CKINVDCx20_ASAP7_75t_R g831 ( 
.A(n_632),
.Y(n_831)
);

CKINVDCx20_ASAP7_75t_R g832 ( 
.A(n_720),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_538),
.Y(n_833)
);

BUFx6f_ASAP7_75t_L g834 ( 
.A(n_544),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_538),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_540),
.Y(n_836)
);

CKINVDCx5p33_ASAP7_75t_R g837 ( 
.A(n_449),
.Y(n_837)
);

INVx2_ASAP7_75t_SL g838 ( 
.A(n_462),
.Y(n_838)
);

INVx2_ASAP7_75t_L g839 ( 
.A(n_605),
.Y(n_839)
);

CKINVDCx5p33_ASAP7_75t_R g840 ( 
.A(n_451),
.Y(n_840)
);

CKINVDCx5p33_ASAP7_75t_R g841 ( 
.A(n_452),
.Y(n_841)
);

CKINVDCx5p33_ASAP7_75t_R g842 ( 
.A(n_456),
.Y(n_842)
);

CKINVDCx20_ASAP7_75t_R g843 ( 
.A(n_554),
.Y(n_843)
);

INVx2_ASAP7_75t_L g844 ( 
.A(n_605),
.Y(n_844)
);

CKINVDCx5p33_ASAP7_75t_R g845 ( 
.A(n_459),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_540),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_547),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_547),
.Y(n_848)
);

CKINVDCx14_ASAP7_75t_R g849 ( 
.A(n_563),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_573),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_573),
.Y(n_851)
);

CKINVDCx5p33_ASAP7_75t_R g852 ( 
.A(n_461),
.Y(n_852)
);

CKINVDCx20_ASAP7_75t_R g853 ( 
.A(n_640),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_579),
.Y(n_854)
);

CKINVDCx16_ASAP7_75t_R g855 ( 
.A(n_640),
.Y(n_855)
);

INVxp67_ASAP7_75t_L g856 ( 
.A(n_530),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_579),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_584),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_584),
.Y(n_859)
);

BUFx10_ASAP7_75t_L g860 ( 
.A(n_668),
.Y(n_860)
);

CKINVDCx20_ASAP7_75t_R g861 ( 
.A(n_441),
.Y(n_861)
);

CKINVDCx5p33_ASAP7_75t_R g862 ( 
.A(n_463),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_586),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_586),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_606),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_606),
.Y(n_866)
);

CKINVDCx20_ASAP7_75t_R g867 ( 
.A(n_444),
.Y(n_867)
);

CKINVDCx5p33_ASAP7_75t_R g868 ( 
.A(n_465),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_608),
.Y(n_869)
);

CKINVDCx16_ASAP7_75t_R g870 ( 
.A(n_563),
.Y(n_870)
);

CKINVDCx16_ASAP7_75t_R g871 ( 
.A(n_563),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_608),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_668),
.Y(n_873)
);

INVxp67_ASAP7_75t_L g874 ( 
.A(n_594),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_668),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_668),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_668),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_668),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_718),
.Y(n_879)
);

CKINVDCx5p33_ASAP7_75t_R g880 ( 
.A(n_467),
.Y(n_880)
);

CKINVDCx20_ASAP7_75t_R g881 ( 
.A(n_448),
.Y(n_881)
);

INVx2_ASAP7_75t_L g882 ( 
.A(n_718),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_618),
.Y(n_883)
);

INVx1_ASAP7_75t_SL g884 ( 
.A(n_484),
.Y(n_884)
);

CKINVDCx5p33_ASAP7_75t_R g885 ( 
.A(n_470),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_618),
.Y(n_886)
);

CKINVDCx5p33_ASAP7_75t_R g887 ( 
.A(n_471),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_620),
.Y(n_888)
);

CKINVDCx20_ASAP7_75t_R g889 ( 
.A(n_455),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_620),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_653),
.Y(n_891)
);

CKINVDCx5p33_ASAP7_75t_R g892 ( 
.A(n_476),
.Y(n_892)
);

CKINVDCx5p33_ASAP7_75t_R g893 ( 
.A(n_485),
.Y(n_893)
);

CKINVDCx5p33_ASAP7_75t_R g894 ( 
.A(n_488),
.Y(n_894)
);

CKINVDCx16_ASAP7_75t_R g895 ( 
.A(n_563),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_653),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_723),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_723),
.Y(n_898)
);

CKINVDCx5p33_ASAP7_75t_R g899 ( 
.A(n_491),
.Y(n_899)
);

INVx2_ASAP7_75t_L g900 ( 
.A(n_718),
.Y(n_900)
);

INVx1_ASAP7_75t_SL g901 ( 
.A(n_502),
.Y(n_901)
);

CKINVDCx20_ASAP7_75t_R g902 ( 
.A(n_469),
.Y(n_902)
);

CKINVDCx5p33_ASAP7_75t_R g903 ( 
.A(n_492),
.Y(n_903)
);

BUFx5_ASAP7_75t_L g904 ( 
.A(n_726),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_726),
.Y(n_905)
);

CKINVDCx5p33_ASAP7_75t_R g906 ( 
.A(n_494),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_752),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_752),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_761),
.Y(n_909)
);

CKINVDCx16_ASAP7_75t_R g910 ( 
.A(n_745),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_761),
.Y(n_911)
);

INVx2_ASAP7_75t_L g912 ( 
.A(n_718),
.Y(n_912)
);

CKINVDCx5p33_ASAP7_75t_R g913 ( 
.A(n_497),
.Y(n_913)
);

INVx2_ASAP7_75t_L g914 ( 
.A(n_718),
.Y(n_914)
);

CKINVDCx20_ASAP7_75t_R g915 ( 
.A(n_481),
.Y(n_915)
);

CKINVDCx5p33_ASAP7_75t_R g916 ( 
.A(n_501),
.Y(n_916)
);

CKINVDCx5p33_ASAP7_75t_R g917 ( 
.A(n_508),
.Y(n_917)
);

CKINVDCx5p33_ASAP7_75t_R g918 ( 
.A(n_509),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_462),
.Y(n_919)
);

BUFx6f_ASAP7_75t_L g920 ( 
.A(n_544),
.Y(n_920)
);

CKINVDCx5p33_ASAP7_75t_R g921 ( 
.A(n_511),
.Y(n_921)
);

INVx2_ASAP7_75t_SL g922 ( 
.A(n_520),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_520),
.Y(n_923)
);

CKINVDCx5p33_ASAP7_75t_R g924 ( 
.A(n_514),
.Y(n_924)
);

CKINVDCx20_ASAP7_75t_R g925 ( 
.A(n_483),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_520),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_671),
.Y(n_927)
);

CKINVDCx5p33_ASAP7_75t_R g928 ( 
.A(n_516),
.Y(n_928)
);

CKINVDCx16_ASAP7_75t_R g929 ( 
.A(n_745),
.Y(n_929)
);

CKINVDCx16_ASAP7_75t_R g930 ( 
.A(n_745),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_671),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_671),
.Y(n_932)
);

INVx1_ASAP7_75t_L g933 ( 
.A(n_701),
.Y(n_933)
);

CKINVDCx5p33_ASAP7_75t_R g934 ( 
.A(n_517),
.Y(n_934)
);

CKINVDCx20_ASAP7_75t_R g935 ( 
.A(n_500),
.Y(n_935)
);

CKINVDCx20_ASAP7_75t_R g936 ( 
.A(n_506),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_701),
.Y(n_937)
);

HB1xp67_ASAP7_75t_L g938 ( 
.A(n_673),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_701),
.Y(n_939)
);

CKINVDCx20_ASAP7_75t_R g940 ( 
.A(n_510),
.Y(n_940)
);

CKINVDCx5p33_ASAP7_75t_R g941 ( 
.A(n_518),
.Y(n_941)
);

INVx1_ASAP7_75t_L g942 ( 
.A(n_721),
.Y(n_942)
);

CKINVDCx5p33_ASAP7_75t_R g943 ( 
.A(n_519),
.Y(n_943)
);

NOR2xp67_ASAP7_75t_L g944 ( 
.A(n_457),
.B(n_1),
.Y(n_944)
);

CKINVDCx5p33_ASAP7_75t_R g945 ( 
.A(n_528),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_721),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_721),
.Y(n_947)
);

INVx1_ASAP7_75t_L g948 ( 
.A(n_478),
.Y(n_948)
);

INVx2_ASAP7_75t_L g949 ( 
.A(n_718),
.Y(n_949)
);

CKINVDCx5p33_ASAP7_75t_R g950 ( 
.A(n_532),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_478),
.Y(n_951)
);

CKINVDCx5p33_ASAP7_75t_R g952 ( 
.A(n_545),
.Y(n_952)
);

INVx1_ASAP7_75t_L g953 ( 
.A(n_742),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_478),
.Y(n_954)
);

INVxp67_ASAP7_75t_L g955 ( 
.A(n_705),
.Y(n_955)
);

INVxp33_ASAP7_75t_L g956 ( 
.A(n_450),
.Y(n_956)
);

CKINVDCx5p33_ASAP7_75t_R g957 ( 
.A(n_548),
.Y(n_957)
);

INVx1_ASAP7_75t_L g958 ( 
.A(n_482),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_482),
.Y(n_959)
);

CKINVDCx5p33_ASAP7_75t_R g960 ( 
.A(n_549),
.Y(n_960)
);

CKINVDCx20_ASAP7_75t_R g961 ( 
.A(n_522),
.Y(n_961)
);

CKINVDCx5p33_ASAP7_75t_R g962 ( 
.A(n_552),
.Y(n_962)
);

BUFx3_ASAP7_75t_L g963 ( 
.A(n_634),
.Y(n_963)
);

CKINVDCx5p33_ASAP7_75t_R g964 ( 
.A(n_553),
.Y(n_964)
);

INVxp67_ASAP7_75t_L g965 ( 
.A(n_453),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_482),
.Y(n_966)
);

INVx2_ASAP7_75t_L g967 ( 
.A(n_742),
.Y(n_967)
);

CKINVDCx5p33_ASAP7_75t_R g968 ( 
.A(n_560),
.Y(n_968)
);

CKINVDCx5p33_ASAP7_75t_R g969 ( 
.A(n_561),
.Y(n_969)
);

HB1xp67_ASAP7_75t_L g970 ( 
.A(n_568),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_562),
.Y(n_971)
);

INVx1_ASAP7_75t_L g972 ( 
.A(n_562),
.Y(n_972)
);

CKINVDCx20_ASAP7_75t_R g973 ( 
.A(n_525),
.Y(n_973)
);

CKINVDCx20_ASAP7_75t_R g974 ( 
.A(n_537),
.Y(n_974)
);

BUFx6f_ASAP7_75t_L g975 ( 
.A(n_544),
.Y(n_975)
);

CKINVDCx5p33_ASAP7_75t_R g976 ( 
.A(n_569),
.Y(n_976)
);

INVx2_ASAP7_75t_SL g977 ( 
.A(n_745),
.Y(n_977)
);

CKINVDCx5p33_ASAP7_75t_R g978 ( 
.A(n_570),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_562),
.Y(n_979)
);

INVx1_ASAP7_75t_L g980 ( 
.A(n_659),
.Y(n_980)
);

INVx1_ASAP7_75t_L g981 ( 
.A(n_659),
.Y(n_981)
);

INVx1_ASAP7_75t_L g982 ( 
.A(n_659),
.Y(n_982)
);

INVxp67_ASAP7_75t_SL g983 ( 
.A(n_742),
.Y(n_983)
);

BUFx6f_ASAP7_75t_L g984 ( 
.A(n_544),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_688),
.Y(n_985)
);

INVx1_ASAP7_75t_L g986 ( 
.A(n_688),
.Y(n_986)
);

CKINVDCx5p33_ASAP7_75t_R g987 ( 
.A(n_571),
.Y(n_987)
);

CKINVDCx5p33_ASAP7_75t_R g988 ( 
.A(n_572),
.Y(n_988)
);

INVxp33_ASAP7_75t_L g989 ( 
.A(n_460),
.Y(n_989)
);

BUFx3_ASAP7_75t_L g990 ( 
.A(n_634),
.Y(n_990)
);

CKINVDCx5p33_ASAP7_75t_R g991 ( 
.A(n_574),
.Y(n_991)
);

CKINVDCx5p33_ASAP7_75t_R g992 ( 
.A(n_576),
.Y(n_992)
);

BUFx6f_ASAP7_75t_L g993 ( 
.A(n_544),
.Y(n_993)
);

CKINVDCx5p33_ASAP7_75t_R g994 ( 
.A(n_580),
.Y(n_994)
);

CKINVDCx20_ASAP7_75t_R g995 ( 
.A(n_546),
.Y(n_995)
);

CKINVDCx5p33_ASAP7_75t_R g996 ( 
.A(n_587),
.Y(n_996)
);

CKINVDCx5p33_ASAP7_75t_R g997 ( 
.A(n_590),
.Y(n_997)
);

CKINVDCx5p33_ASAP7_75t_R g998 ( 
.A(n_595),
.Y(n_998)
);

CKINVDCx5p33_ASAP7_75t_R g999 ( 
.A(n_596),
.Y(n_999)
);

CKINVDCx5p33_ASAP7_75t_R g1000 ( 
.A(n_598),
.Y(n_1000)
);

CKINVDCx5p33_ASAP7_75t_R g1001 ( 
.A(n_603),
.Y(n_1001)
);

CKINVDCx5p33_ASAP7_75t_R g1002 ( 
.A(n_607),
.Y(n_1002)
);

INVx1_ASAP7_75t_L g1003 ( 
.A(n_688),
.Y(n_1003)
);

INVx2_ASAP7_75t_L g1004 ( 
.A(n_742),
.Y(n_1004)
);

INVx1_ASAP7_75t_L g1005 ( 
.A(n_690),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_690),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_690),
.Y(n_1007)
);

INVx1_ASAP7_75t_L g1008 ( 
.A(n_740),
.Y(n_1008)
);

CKINVDCx20_ASAP7_75t_R g1009 ( 
.A(n_550),
.Y(n_1009)
);

CKINVDCx5p33_ASAP7_75t_R g1010 ( 
.A(n_609),
.Y(n_1010)
);

CKINVDCx5p33_ASAP7_75t_R g1011 ( 
.A(n_611),
.Y(n_1011)
);

CKINVDCx16_ASAP7_75t_R g1012 ( 
.A(n_634),
.Y(n_1012)
);

CKINVDCx20_ASAP7_75t_R g1013 ( 
.A(n_583),
.Y(n_1013)
);

CKINVDCx5p33_ASAP7_75t_R g1014 ( 
.A(n_612),
.Y(n_1014)
);

CKINVDCx20_ASAP7_75t_R g1015 ( 
.A(n_588),
.Y(n_1015)
);

CKINVDCx16_ASAP7_75t_R g1016 ( 
.A(n_521),
.Y(n_1016)
);

CKINVDCx5p33_ASAP7_75t_R g1017 ( 
.A(n_614),
.Y(n_1017)
);

BUFx3_ASAP7_75t_L g1018 ( 
.A(n_601),
.Y(n_1018)
);

CKINVDCx20_ASAP7_75t_R g1019 ( 
.A(n_604),
.Y(n_1019)
);

INVx1_ASAP7_75t_L g1020 ( 
.A(n_740),
.Y(n_1020)
);

INVx1_ASAP7_75t_L g1021 ( 
.A(n_740),
.Y(n_1021)
);

INVxp67_ASAP7_75t_L g1022 ( 
.A(n_460),
.Y(n_1022)
);

CKINVDCx5p33_ASAP7_75t_R g1023 ( 
.A(n_624),
.Y(n_1023)
);

INVx1_ASAP7_75t_L g1024 ( 
.A(n_742),
.Y(n_1024)
);

INVxp67_ASAP7_75t_SL g1025 ( 
.A(n_742),
.Y(n_1025)
);

INVx1_ASAP7_75t_L g1026 ( 
.A(n_757),
.Y(n_1026)
);

CKINVDCx20_ASAP7_75t_R g1027 ( 
.A(n_613),
.Y(n_1027)
);

INVx1_ASAP7_75t_L g1028 ( 
.A(n_757),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_757),
.Y(n_1029)
);

BUFx6f_ASAP7_75t_L g1030 ( 
.A(n_578),
.Y(n_1030)
);

INVx1_ASAP7_75t_L g1031 ( 
.A(n_757),
.Y(n_1031)
);

INVxp67_ASAP7_75t_L g1032 ( 
.A(n_473),
.Y(n_1032)
);

INVx1_ASAP7_75t_L g1033 ( 
.A(n_757),
.Y(n_1033)
);

CKINVDCx5p33_ASAP7_75t_R g1034 ( 
.A(n_626),
.Y(n_1034)
);

INVx1_ASAP7_75t_L g1035 ( 
.A(n_757),
.Y(n_1035)
);

XOR2xp5_ASAP7_75t_L g1036 ( 
.A(n_575),
.B(n_2),
.Y(n_1036)
);

AND2x4_ASAP7_75t_L g1037 ( 
.A(n_578),
.B(n_290),
.Y(n_1037)
);

INVx1_ASAP7_75t_L g1038 ( 
.A(n_473),
.Y(n_1038)
);

CKINVDCx20_ASAP7_75t_R g1039 ( 
.A(n_621),
.Y(n_1039)
);

CKINVDCx5p33_ASAP7_75t_R g1040 ( 
.A(n_633),
.Y(n_1040)
);

CKINVDCx20_ASAP7_75t_R g1041 ( 
.A(n_625),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_475),
.Y(n_1042)
);

CKINVDCx5p33_ASAP7_75t_R g1043 ( 
.A(n_635),
.Y(n_1043)
);

INVx1_ASAP7_75t_L g1044 ( 
.A(n_475),
.Y(n_1044)
);

INVx2_ASAP7_75t_SL g1045 ( 
.A(n_458),
.Y(n_1045)
);

CKINVDCx5p33_ASAP7_75t_R g1046 ( 
.A(n_636),
.Y(n_1046)
);

INVx2_ASAP7_75t_L g1047 ( 
.A(n_458),
.Y(n_1047)
);

CKINVDCx5p33_ASAP7_75t_R g1048 ( 
.A(n_639),
.Y(n_1048)
);

INVx1_ASAP7_75t_L g1049 ( 
.A(n_479),
.Y(n_1049)
);

INVx1_ASAP7_75t_L g1050 ( 
.A(n_479),
.Y(n_1050)
);

INVx1_ASAP7_75t_L g1051 ( 
.A(n_493),
.Y(n_1051)
);

CKINVDCx5p33_ASAP7_75t_R g1052 ( 
.A(n_641),
.Y(n_1052)
);

CKINVDCx5p33_ASAP7_75t_R g1053 ( 
.A(n_642),
.Y(n_1053)
);

INVx1_ASAP7_75t_SL g1054 ( 
.A(n_591),
.Y(n_1054)
);

HB1xp67_ASAP7_75t_L g1055 ( 
.A(n_644),
.Y(n_1055)
);

INVx1_ASAP7_75t_L g1056 ( 
.A(n_493),
.Y(n_1056)
);

BUFx10_ASAP7_75t_L g1057 ( 
.A(n_542),
.Y(n_1057)
);

INVx2_ASAP7_75t_SL g1058 ( 
.A(n_458),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_496),
.Y(n_1059)
);

INVx1_ASAP7_75t_L g1060 ( 
.A(n_496),
.Y(n_1060)
);

INVxp67_ASAP7_75t_L g1061 ( 
.A(n_504),
.Y(n_1061)
);

CKINVDCx5p33_ASAP7_75t_R g1062 ( 
.A(n_647),
.Y(n_1062)
);

CKINVDCx5p33_ASAP7_75t_R g1063 ( 
.A(n_649),
.Y(n_1063)
);

CKINVDCx5p33_ASAP7_75t_R g1064 ( 
.A(n_650),
.Y(n_1064)
);

INVx1_ASAP7_75t_L g1065 ( 
.A(n_504),
.Y(n_1065)
);

CKINVDCx5p33_ASAP7_75t_R g1066 ( 
.A(n_651),
.Y(n_1066)
);

BUFx6f_ASAP7_75t_L g1067 ( 
.A(n_578),
.Y(n_1067)
);

INVx1_ASAP7_75t_L g1068 ( 
.A(n_505),
.Y(n_1068)
);

OR2x2_ASAP7_75t_L g1069 ( 
.A(n_505),
.B(n_2),
.Y(n_1069)
);

INVx1_ASAP7_75t_L g1070 ( 
.A(n_526),
.Y(n_1070)
);

CKINVDCx5p33_ASAP7_75t_R g1071 ( 
.A(n_652),
.Y(n_1071)
);

INVx1_ASAP7_75t_L g1072 ( 
.A(n_526),
.Y(n_1072)
);

CKINVDCx5p33_ASAP7_75t_R g1073 ( 
.A(n_655),
.Y(n_1073)
);

INVx1_ASAP7_75t_L g1074 ( 
.A(n_527),
.Y(n_1074)
);

INVx1_ASAP7_75t_L g1075 ( 
.A(n_527),
.Y(n_1075)
);

BUFx2_ASAP7_75t_SL g1076 ( 
.A(n_542),
.Y(n_1076)
);

CKINVDCx5p33_ASAP7_75t_R g1077 ( 
.A(n_657),
.Y(n_1077)
);

CKINVDCx20_ASAP7_75t_R g1078 ( 
.A(n_630),
.Y(n_1078)
);

INVx3_ASAP7_75t_L g1079 ( 
.A(n_472),
.Y(n_1079)
);

INVx1_ASAP7_75t_L g1080 ( 
.A(n_529),
.Y(n_1080)
);

INVx1_ASAP7_75t_L g1081 ( 
.A(n_529),
.Y(n_1081)
);

INVx1_ASAP7_75t_L g1082 ( 
.A(n_531),
.Y(n_1082)
);

INVx1_ASAP7_75t_L g1083 ( 
.A(n_531),
.Y(n_1083)
);

INVx1_ASAP7_75t_L g1084 ( 
.A(n_533),
.Y(n_1084)
);

CKINVDCx5p33_ASAP7_75t_R g1085 ( 
.A(n_661),
.Y(n_1085)
);

BUFx3_ASAP7_75t_L g1086 ( 
.A(n_637),
.Y(n_1086)
);

INVxp67_ASAP7_75t_SL g1087 ( 
.A(n_660),
.Y(n_1087)
);

BUFx2_ASAP7_75t_L g1088 ( 
.A(n_662),
.Y(n_1088)
);

CKINVDCx5p33_ASAP7_75t_R g1089 ( 
.A(n_665),
.Y(n_1089)
);

CKINVDCx20_ASAP7_75t_R g1090 ( 
.A(n_638),
.Y(n_1090)
);

INVx1_ASAP7_75t_L g1091 ( 
.A(n_533),
.Y(n_1091)
);

INVx1_ASAP7_75t_L g1092 ( 
.A(n_535),
.Y(n_1092)
);

HB1xp67_ASAP7_75t_L g1093 ( 
.A(n_674),
.Y(n_1093)
);

CKINVDCx5p33_ASAP7_75t_R g1094 ( 
.A(n_677),
.Y(n_1094)
);

CKINVDCx5p33_ASAP7_75t_R g1095 ( 
.A(n_681),
.Y(n_1095)
);

CKINVDCx5p33_ASAP7_75t_R g1096 ( 
.A(n_682),
.Y(n_1096)
);

NOR2xp67_ASAP7_75t_L g1097 ( 
.A(n_495),
.B(n_3),
.Y(n_1097)
);

BUFx6f_ASAP7_75t_L g1098 ( 
.A(n_578),
.Y(n_1098)
);

INVx1_ASAP7_75t_L g1099 ( 
.A(n_535),
.Y(n_1099)
);

INVx1_ASAP7_75t_L g1100 ( 
.A(n_539),
.Y(n_1100)
);

INVx1_ASAP7_75t_L g1101 ( 
.A(n_539),
.Y(n_1101)
);

CKINVDCx5p33_ASAP7_75t_R g1102 ( 
.A(n_684),
.Y(n_1102)
);

INVx1_ASAP7_75t_L g1103 ( 
.A(n_541),
.Y(n_1103)
);

CKINVDCx5p33_ASAP7_75t_R g1104 ( 
.A(n_687),
.Y(n_1104)
);

CKINVDCx20_ASAP7_75t_R g1105 ( 
.A(n_643),
.Y(n_1105)
);

CKINVDCx5p33_ASAP7_75t_R g1106 ( 
.A(n_693),
.Y(n_1106)
);

CKINVDCx20_ASAP7_75t_R g1107 ( 
.A(n_648),
.Y(n_1107)
);

INVx1_ASAP7_75t_L g1108 ( 
.A(n_541),
.Y(n_1108)
);

CKINVDCx5p33_ASAP7_75t_R g1109 ( 
.A(n_694),
.Y(n_1109)
);

CKINVDCx5p33_ASAP7_75t_R g1110 ( 
.A(n_695),
.Y(n_1110)
);

CKINVDCx20_ASAP7_75t_R g1111 ( 
.A(n_656),
.Y(n_1111)
);

BUFx6f_ASAP7_75t_L g1112 ( 
.A(n_578),
.Y(n_1112)
);

BUFx3_ASAP7_75t_L g1113 ( 
.A(n_658),
.Y(n_1113)
);

CKINVDCx5p33_ASAP7_75t_R g1114 ( 
.A(n_696),
.Y(n_1114)
);

INVx1_ASAP7_75t_L g1115 ( 
.A(n_543),
.Y(n_1115)
);

BUFx2_ASAP7_75t_L g1116 ( 
.A(n_697),
.Y(n_1116)
);

CKINVDCx5p33_ASAP7_75t_R g1117 ( 
.A(n_700),
.Y(n_1117)
);

INVx1_ASAP7_75t_L g1118 ( 
.A(n_543),
.Y(n_1118)
);

INVx1_ASAP7_75t_L g1119 ( 
.A(n_556),
.Y(n_1119)
);

INVx2_ASAP7_75t_SL g1120 ( 
.A(n_472),
.Y(n_1120)
);

INVx1_ASAP7_75t_L g1121 ( 
.A(n_556),
.Y(n_1121)
);

CKINVDCx16_ASAP7_75t_R g1122 ( 
.A(n_617),
.Y(n_1122)
);

CKINVDCx16_ASAP7_75t_R g1123 ( 
.A(n_646),
.Y(n_1123)
);

INVx1_ASAP7_75t_L g1124 ( 
.A(n_557),
.Y(n_1124)
);

CKINVDCx5p33_ASAP7_75t_R g1125 ( 
.A(n_704),
.Y(n_1125)
);

BUFx6f_ASAP7_75t_L g1126 ( 
.A(n_578),
.Y(n_1126)
);

CKINVDCx5p33_ASAP7_75t_R g1127 ( 
.A(n_707),
.Y(n_1127)
);

INVx1_ASAP7_75t_L g1128 ( 
.A(n_557),
.Y(n_1128)
);

CKINVDCx5p33_ASAP7_75t_R g1129 ( 
.A(n_711),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_558),
.Y(n_1130)
);

INVx1_ASAP7_75t_L g1131 ( 
.A(n_558),
.Y(n_1131)
);

INVx1_ASAP7_75t_L g1132 ( 
.A(n_559),
.Y(n_1132)
);

INVxp67_ASAP7_75t_SL g1133 ( 
.A(n_685),
.Y(n_1133)
);

CKINVDCx5p33_ASAP7_75t_R g1134 ( 
.A(n_714),
.Y(n_1134)
);

INVxp67_ASAP7_75t_SL g1135 ( 
.A(n_781),
.Y(n_1135)
);

NOR2xp33_ASAP7_75t_L g1136 ( 
.A(n_811),
.B(n_564),
.Y(n_1136)
);

HB1xp67_ASAP7_75t_L g1137 ( 
.A(n_779),
.Y(n_1137)
);

CKINVDCx20_ASAP7_75t_R g1138 ( 
.A(n_771),
.Y(n_1138)
);

CKINVDCx5p33_ASAP7_75t_R g1139 ( 
.A(n_861),
.Y(n_1139)
);

INVxp67_ASAP7_75t_L g1140 ( 
.A(n_970),
.Y(n_1140)
);

INVx1_ASAP7_75t_L g1141 ( 
.A(n_983),
.Y(n_1141)
);

CKINVDCx16_ASAP7_75t_R g1142 ( 
.A(n_816),
.Y(n_1142)
);

INVx1_ASAP7_75t_L g1143 ( 
.A(n_1025),
.Y(n_1143)
);

NOR2xp33_ASAP7_75t_L g1144 ( 
.A(n_811),
.B(n_582),
.Y(n_1144)
);

CKINVDCx14_ASAP7_75t_R g1145 ( 
.A(n_849),
.Y(n_1145)
);

CKINVDCx20_ASAP7_75t_R g1146 ( 
.A(n_801),
.Y(n_1146)
);

INVx1_ASAP7_75t_L g1147 ( 
.A(n_1024),
.Y(n_1147)
);

CKINVDCx5p33_ASAP7_75t_R g1148 ( 
.A(n_867),
.Y(n_1148)
);

INVx1_ASAP7_75t_L g1149 ( 
.A(n_1026),
.Y(n_1149)
);

HB1xp67_ASAP7_75t_L g1150 ( 
.A(n_779),
.Y(n_1150)
);

INVx1_ASAP7_75t_L g1151 ( 
.A(n_1028),
.Y(n_1151)
);

INVx1_ASAP7_75t_L g1152 ( 
.A(n_1029),
.Y(n_1152)
);

INVx1_ASAP7_75t_L g1153 ( 
.A(n_1031),
.Y(n_1153)
);

NOR2xp33_ASAP7_75t_L g1154 ( 
.A(n_1018),
.B(n_629),
.Y(n_1154)
);

CKINVDCx5p33_ASAP7_75t_R g1155 ( 
.A(n_881),
.Y(n_1155)
);

CKINVDCx5p33_ASAP7_75t_R g1156 ( 
.A(n_889),
.Y(n_1156)
);

INVx1_ASAP7_75t_L g1157 ( 
.A(n_1033),
.Y(n_1157)
);

INVx1_ASAP7_75t_L g1158 ( 
.A(n_1035),
.Y(n_1158)
);

CKINVDCx5p33_ASAP7_75t_R g1159 ( 
.A(n_902),
.Y(n_1159)
);

CKINVDCx5p33_ASAP7_75t_R g1160 ( 
.A(n_915),
.Y(n_1160)
);

CKINVDCx5p33_ASAP7_75t_R g1161 ( 
.A(n_925),
.Y(n_1161)
);

CKINVDCx20_ASAP7_75t_R g1162 ( 
.A(n_831),
.Y(n_1162)
);

INVxp67_ASAP7_75t_SL g1163 ( 
.A(n_1018),
.Y(n_1163)
);

INVxp67_ASAP7_75t_SL g1164 ( 
.A(n_1086),
.Y(n_1164)
);

NOR2xp33_ASAP7_75t_L g1165 ( 
.A(n_1086),
.B(n_680),
.Y(n_1165)
);

INVxp67_ASAP7_75t_L g1166 ( 
.A(n_1055),
.Y(n_1166)
);

CKINVDCx5p33_ASAP7_75t_R g1167 ( 
.A(n_935),
.Y(n_1167)
);

CKINVDCx5p33_ASAP7_75t_R g1168 ( 
.A(n_936),
.Y(n_1168)
);

CKINVDCx20_ASAP7_75t_R g1169 ( 
.A(n_832),
.Y(n_1169)
);

INVxp33_ASAP7_75t_SL g1170 ( 
.A(n_777),
.Y(n_1170)
);

INVxp67_ASAP7_75t_SL g1171 ( 
.A(n_1113),
.Y(n_1171)
);

CKINVDCx20_ASAP7_75t_R g1172 ( 
.A(n_940),
.Y(n_1172)
);

INVx1_ASAP7_75t_L g1173 ( 
.A(n_873),
.Y(n_1173)
);

CKINVDCx5p33_ASAP7_75t_R g1174 ( 
.A(n_961),
.Y(n_1174)
);

INVx1_ASAP7_75t_L g1175 ( 
.A(n_873),
.Y(n_1175)
);

INVx1_ASAP7_75t_L g1176 ( 
.A(n_875),
.Y(n_1176)
);

CKINVDCx20_ASAP7_75t_R g1177 ( 
.A(n_973),
.Y(n_1177)
);

CKINVDCx5p33_ASAP7_75t_R g1178 ( 
.A(n_974),
.Y(n_1178)
);

CKINVDCx5p33_ASAP7_75t_R g1179 ( 
.A(n_995),
.Y(n_1179)
);

INVx1_ASAP7_75t_L g1180 ( 
.A(n_875),
.Y(n_1180)
);

INVx1_ASAP7_75t_L g1181 ( 
.A(n_876),
.Y(n_1181)
);

INVx1_ASAP7_75t_L g1182 ( 
.A(n_876),
.Y(n_1182)
);

CKINVDCx5p33_ASAP7_75t_R g1183 ( 
.A(n_1009),
.Y(n_1183)
);

CKINVDCx20_ASAP7_75t_R g1184 ( 
.A(n_1013),
.Y(n_1184)
);

CKINVDCx5p33_ASAP7_75t_R g1185 ( 
.A(n_1015),
.Y(n_1185)
);

INVx1_ASAP7_75t_L g1186 ( 
.A(n_877),
.Y(n_1186)
);

INVx1_ASAP7_75t_L g1187 ( 
.A(n_877),
.Y(n_1187)
);

INVx1_ASAP7_75t_L g1188 ( 
.A(n_878),
.Y(n_1188)
);

INVx1_ASAP7_75t_L g1189 ( 
.A(n_878),
.Y(n_1189)
);

CKINVDCx20_ASAP7_75t_R g1190 ( 
.A(n_1019),
.Y(n_1190)
);

INVx1_ASAP7_75t_L g1191 ( 
.A(n_879),
.Y(n_1191)
);

INVx1_ASAP7_75t_L g1192 ( 
.A(n_879),
.Y(n_1192)
);

CKINVDCx5p33_ASAP7_75t_R g1193 ( 
.A(n_1027),
.Y(n_1193)
);

CKINVDCx20_ASAP7_75t_R g1194 ( 
.A(n_1039),
.Y(n_1194)
);

INVx1_ASAP7_75t_L g1195 ( 
.A(n_953),
.Y(n_1195)
);

CKINVDCx5p33_ASAP7_75t_R g1196 ( 
.A(n_1041),
.Y(n_1196)
);

INVxp67_ASAP7_75t_SL g1197 ( 
.A(n_1113),
.Y(n_1197)
);

CKINVDCx5p33_ASAP7_75t_R g1198 ( 
.A(n_1078),
.Y(n_1198)
);

INVx1_ASAP7_75t_L g1199 ( 
.A(n_953),
.Y(n_1199)
);

CKINVDCx20_ASAP7_75t_R g1200 ( 
.A(n_1090),
.Y(n_1200)
);

INVx1_ASAP7_75t_L g1201 ( 
.A(n_919),
.Y(n_1201)
);

INVx1_ASAP7_75t_L g1202 ( 
.A(n_800),
.Y(n_1202)
);

INVx1_ASAP7_75t_L g1203 ( 
.A(n_800),
.Y(n_1203)
);

INVx3_ASAP7_75t_L g1204 ( 
.A(n_784),
.Y(n_1204)
);

CKINVDCx16_ASAP7_75t_R g1205 ( 
.A(n_855),
.Y(n_1205)
);

CKINVDCx5p33_ASAP7_75t_R g1206 ( 
.A(n_1105),
.Y(n_1206)
);

INVx1_ASAP7_75t_L g1207 ( 
.A(n_802),
.Y(n_1207)
);

INVxp67_ASAP7_75t_L g1208 ( 
.A(n_1093),
.Y(n_1208)
);

CKINVDCx5p33_ASAP7_75t_R g1209 ( 
.A(n_1107),
.Y(n_1209)
);

INVxp33_ASAP7_75t_SL g1210 ( 
.A(n_777),
.Y(n_1210)
);

CKINVDCx5p33_ASAP7_75t_R g1211 ( 
.A(n_1111),
.Y(n_1211)
);

INVx2_ASAP7_75t_L g1212 ( 
.A(n_802),
.Y(n_1212)
);

INVx1_ASAP7_75t_L g1213 ( 
.A(n_826),
.Y(n_1213)
);

CKINVDCx5p33_ASAP7_75t_R g1214 ( 
.A(n_772),
.Y(n_1214)
);

INVx1_ASAP7_75t_L g1215 ( 
.A(n_826),
.Y(n_1215)
);

INVx1_ASAP7_75t_L g1216 ( 
.A(n_839),
.Y(n_1216)
);

NAND2xp5_ASAP7_75t_L g1217 ( 
.A(n_1087),
.B(n_669),
.Y(n_1217)
);

INVx1_ASAP7_75t_L g1218 ( 
.A(n_839),
.Y(n_1218)
);

NAND2xp5_ASAP7_75t_L g1219 ( 
.A(n_1133),
.B(n_686),
.Y(n_1219)
);

INVx1_ASAP7_75t_L g1220 ( 
.A(n_844),
.Y(n_1220)
);

CKINVDCx20_ASAP7_75t_R g1221 ( 
.A(n_843),
.Y(n_1221)
);

INVx1_ASAP7_75t_L g1222 ( 
.A(n_923),
.Y(n_1222)
);

INVx1_ASAP7_75t_L g1223 ( 
.A(n_926),
.Y(n_1223)
);

CKINVDCx5p33_ASAP7_75t_R g1224 ( 
.A(n_853),
.Y(n_1224)
);

INVx1_ASAP7_75t_L g1225 ( 
.A(n_927),
.Y(n_1225)
);

INVxp33_ASAP7_75t_SL g1226 ( 
.A(n_786),
.Y(n_1226)
);

CKINVDCx5p33_ASAP7_75t_R g1227 ( 
.A(n_790),
.Y(n_1227)
);

INVx1_ASAP7_75t_L g1228 ( 
.A(n_931),
.Y(n_1228)
);

CKINVDCx5p33_ASAP7_75t_R g1229 ( 
.A(n_790),
.Y(n_1229)
);

INVxp67_ASAP7_75t_SL g1230 ( 
.A(n_797),
.Y(n_1230)
);

CKINVDCx20_ASAP7_75t_R g1231 ( 
.A(n_1016),
.Y(n_1231)
);

CKINVDCx5p33_ASAP7_75t_R g1232 ( 
.A(n_792),
.Y(n_1232)
);

INVx1_ASAP7_75t_L g1233 ( 
.A(n_844),
.Y(n_1233)
);

INVx1_ASAP7_75t_L g1234 ( 
.A(n_932),
.Y(n_1234)
);

INVx1_ASAP7_75t_L g1235 ( 
.A(n_933),
.Y(n_1235)
);

INVx1_ASAP7_75t_L g1236 ( 
.A(n_937),
.Y(n_1236)
);

INVx1_ASAP7_75t_L g1237 ( 
.A(n_939),
.Y(n_1237)
);

CKINVDCx5p33_ASAP7_75t_R g1238 ( 
.A(n_792),
.Y(n_1238)
);

INVxp67_ASAP7_75t_SL g1239 ( 
.A(n_797),
.Y(n_1239)
);

CKINVDCx20_ASAP7_75t_R g1240 ( 
.A(n_1122),
.Y(n_1240)
);

INVx1_ASAP7_75t_L g1241 ( 
.A(n_942),
.Y(n_1241)
);

NOR2xp33_ASAP7_75t_L g1242 ( 
.A(n_789),
.B(n_963),
.Y(n_1242)
);

INVx1_ASAP7_75t_L g1243 ( 
.A(n_946),
.Y(n_1243)
);

INVx1_ASAP7_75t_SL g1244 ( 
.A(n_830),
.Y(n_1244)
);

CKINVDCx20_ASAP7_75t_R g1245 ( 
.A(n_1123),
.Y(n_1245)
);

CKINVDCx20_ASAP7_75t_R g1246 ( 
.A(n_884),
.Y(n_1246)
);

CKINVDCx20_ASAP7_75t_R g1247 ( 
.A(n_901),
.Y(n_1247)
);

CKINVDCx5p33_ASAP7_75t_R g1248 ( 
.A(n_805),
.Y(n_1248)
);

INVxp67_ASAP7_75t_SL g1249 ( 
.A(n_838),
.Y(n_1249)
);

NOR2xp33_ASAP7_75t_L g1250 ( 
.A(n_789),
.B(n_762),
.Y(n_1250)
);

INVx1_ASAP7_75t_L g1251 ( 
.A(n_947),
.Y(n_1251)
);

CKINVDCx20_ASAP7_75t_R g1252 ( 
.A(n_1054),
.Y(n_1252)
);

CKINVDCx5p33_ASAP7_75t_R g1253 ( 
.A(n_805),
.Y(n_1253)
);

INVx1_ASAP7_75t_L g1254 ( 
.A(n_791),
.Y(n_1254)
);

INVx1_ASAP7_75t_L g1255 ( 
.A(n_793),
.Y(n_1255)
);

NAND2xp5_ASAP7_75t_L g1256 ( 
.A(n_963),
.B(n_990),
.Y(n_1256)
);

CKINVDCx5p33_ASAP7_75t_R g1257 ( 
.A(n_806),
.Y(n_1257)
);

CKINVDCx5p33_ASAP7_75t_R g1258 ( 
.A(n_806),
.Y(n_1258)
);

CKINVDCx14_ASAP7_75t_R g1259 ( 
.A(n_823),
.Y(n_1259)
);

INVx1_ASAP7_75t_L g1260 ( 
.A(n_794),
.Y(n_1260)
);

CKINVDCx20_ASAP7_75t_R g1261 ( 
.A(n_786),
.Y(n_1261)
);

CKINVDCx5p33_ASAP7_75t_R g1262 ( 
.A(n_807),
.Y(n_1262)
);

INVx1_ASAP7_75t_L g1263 ( 
.A(n_795),
.Y(n_1263)
);

CKINVDCx20_ASAP7_75t_R g1264 ( 
.A(n_1012),
.Y(n_1264)
);

CKINVDCx5p33_ASAP7_75t_R g1265 ( 
.A(n_807),
.Y(n_1265)
);

INVx1_ASAP7_75t_L g1266 ( 
.A(n_796),
.Y(n_1266)
);

NOR2xp33_ASAP7_75t_L g1267 ( 
.A(n_990),
.B(n_769),
.Y(n_1267)
);

CKINVDCx20_ASAP7_75t_R g1268 ( 
.A(n_798),
.Y(n_1268)
);

CKINVDCx20_ASAP7_75t_R g1269 ( 
.A(n_870),
.Y(n_1269)
);

CKINVDCx20_ASAP7_75t_R g1270 ( 
.A(n_871),
.Y(n_1270)
);

CKINVDCx5p33_ASAP7_75t_R g1271 ( 
.A(n_819),
.Y(n_1271)
);

INVx1_ASAP7_75t_L g1272 ( 
.A(n_799),
.Y(n_1272)
);

CKINVDCx5p33_ASAP7_75t_R g1273 ( 
.A(n_819),
.Y(n_1273)
);

NAND2xp5_ASAP7_75t_L g1274 ( 
.A(n_838),
.B(n_689),
.Y(n_1274)
);

CKINVDCx5p33_ASAP7_75t_R g1275 ( 
.A(n_837),
.Y(n_1275)
);

INVxp67_ASAP7_75t_L g1276 ( 
.A(n_1088),
.Y(n_1276)
);

INVx1_ASAP7_75t_L g1277 ( 
.A(n_803),
.Y(n_1277)
);

CKINVDCx5p33_ASAP7_75t_R g1278 ( 
.A(n_837),
.Y(n_1278)
);

CKINVDCx5p33_ASAP7_75t_R g1279 ( 
.A(n_840),
.Y(n_1279)
);

INVx2_ASAP7_75t_L g1280 ( 
.A(n_882),
.Y(n_1280)
);

CKINVDCx20_ASAP7_75t_R g1281 ( 
.A(n_895),
.Y(n_1281)
);

INVx1_ASAP7_75t_L g1282 ( 
.A(n_804),
.Y(n_1282)
);

CKINVDCx20_ASAP7_75t_R g1283 ( 
.A(n_910),
.Y(n_1283)
);

NOR2xp67_ASAP7_75t_L g1284 ( 
.A(n_840),
.B(n_713),
.Y(n_1284)
);

CKINVDCx5p33_ASAP7_75t_R g1285 ( 
.A(n_841),
.Y(n_1285)
);

CKINVDCx20_ASAP7_75t_R g1286 ( 
.A(n_929),
.Y(n_1286)
);

CKINVDCx16_ASAP7_75t_R g1287 ( 
.A(n_930),
.Y(n_1287)
);

HB1xp67_ASAP7_75t_L g1288 ( 
.A(n_841),
.Y(n_1288)
);

INVxp67_ASAP7_75t_L g1289 ( 
.A(n_1088),
.Y(n_1289)
);

CKINVDCx5p33_ASAP7_75t_R g1290 ( 
.A(n_842),
.Y(n_1290)
);

INVxp67_ASAP7_75t_L g1291 ( 
.A(n_1116),
.Y(n_1291)
);

CKINVDCx20_ASAP7_75t_R g1292 ( 
.A(n_842),
.Y(n_1292)
);

INVx1_ASAP7_75t_L g1293 ( 
.A(n_808),
.Y(n_1293)
);

INVx1_ASAP7_75t_L g1294 ( 
.A(n_809),
.Y(n_1294)
);

OR2x2_ASAP7_75t_L g1295 ( 
.A(n_783),
.B(n_654),
.Y(n_1295)
);

CKINVDCx20_ASAP7_75t_R g1296 ( 
.A(n_845),
.Y(n_1296)
);

CKINVDCx16_ASAP7_75t_R g1297 ( 
.A(n_829),
.Y(n_1297)
);

INVx1_ASAP7_75t_L g1298 ( 
.A(n_810),
.Y(n_1298)
);

INVx1_ASAP7_75t_L g1299 ( 
.A(n_813),
.Y(n_1299)
);

INVx1_ASAP7_75t_L g1300 ( 
.A(n_814),
.Y(n_1300)
);

INVx1_ASAP7_75t_L g1301 ( 
.A(n_815),
.Y(n_1301)
);

INVx1_ASAP7_75t_L g1302 ( 
.A(n_818),
.Y(n_1302)
);

INVx1_ASAP7_75t_L g1303 ( 
.A(n_820),
.Y(n_1303)
);

INVx2_ASAP7_75t_L g1304 ( 
.A(n_882),
.Y(n_1304)
);

CKINVDCx5p33_ASAP7_75t_R g1305 ( 
.A(n_845),
.Y(n_1305)
);

CKINVDCx20_ASAP7_75t_R g1306 ( 
.A(n_852),
.Y(n_1306)
);

CKINVDCx5p33_ASAP7_75t_R g1307 ( 
.A(n_852),
.Y(n_1307)
);

NAND2xp5_ASAP7_75t_L g1308 ( 
.A(n_922),
.B(n_698),
.Y(n_1308)
);

NOR2xp33_ASAP7_75t_L g1309 ( 
.A(n_821),
.B(n_764),
.Y(n_1309)
);

NOR2xp33_ASAP7_75t_L g1310 ( 
.A(n_862),
.B(n_868),
.Y(n_1310)
);

CKINVDCx5p33_ASAP7_75t_R g1311 ( 
.A(n_862),
.Y(n_1311)
);

CKINVDCx5p33_ASAP7_75t_R g1312 ( 
.A(n_868),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_822),
.Y(n_1313)
);

NOR2xp33_ASAP7_75t_L g1314 ( 
.A(n_880),
.B(n_885),
.Y(n_1314)
);

INVx1_ASAP7_75t_L g1315 ( 
.A(n_825),
.Y(n_1315)
);

INVx1_ASAP7_75t_L g1316 ( 
.A(n_827),
.Y(n_1316)
);

INVx1_ASAP7_75t_L g1317 ( 
.A(n_828),
.Y(n_1317)
);

CKINVDCx5p33_ASAP7_75t_R g1318 ( 
.A(n_880),
.Y(n_1318)
);

INVxp67_ASAP7_75t_L g1319 ( 
.A(n_1116),
.Y(n_1319)
);

INVxp67_ASAP7_75t_L g1320 ( 
.A(n_977),
.Y(n_1320)
);

OR2x2_ASAP7_75t_L g1321 ( 
.A(n_922),
.B(n_654),
.Y(n_1321)
);

INVx1_ASAP7_75t_L g1322 ( 
.A(n_833),
.Y(n_1322)
);

INVx1_ASAP7_75t_L g1323 ( 
.A(n_900),
.Y(n_1323)
);

INVxp67_ASAP7_75t_L g1324 ( 
.A(n_977),
.Y(n_1324)
);

CKINVDCx16_ASAP7_75t_R g1325 ( 
.A(n_775),
.Y(n_1325)
);

INVxp33_ASAP7_75t_SL g1326 ( 
.A(n_885),
.Y(n_1326)
);

INVx1_ASAP7_75t_L g1327 ( 
.A(n_900),
.Y(n_1327)
);

OR2x2_ASAP7_75t_L g1328 ( 
.A(n_1076),
.B(n_691),
.Y(n_1328)
);

INVx1_ASAP7_75t_L g1329 ( 
.A(n_912),
.Y(n_1329)
);

HB1xp67_ASAP7_75t_L g1330 ( 
.A(n_887),
.Y(n_1330)
);

CKINVDCx20_ASAP7_75t_R g1331 ( 
.A(n_887),
.Y(n_1331)
);

BUFx2_ASAP7_75t_SL g1332 ( 
.A(n_1037),
.Y(n_1332)
);

INVxp67_ASAP7_75t_L g1333 ( 
.A(n_938),
.Y(n_1333)
);

CKINVDCx5p33_ASAP7_75t_R g1334 ( 
.A(n_892),
.Y(n_1334)
);

CKINVDCx16_ASAP7_75t_R g1335 ( 
.A(n_775),
.Y(n_1335)
);

INVxp67_ASAP7_75t_SL g1336 ( 
.A(n_784),
.Y(n_1336)
);

CKINVDCx20_ASAP7_75t_R g1337 ( 
.A(n_892),
.Y(n_1337)
);

NAND2xp5_ASAP7_75t_L g1338 ( 
.A(n_1037),
.B(n_706),
.Y(n_1338)
);

INVx1_ASAP7_75t_L g1339 ( 
.A(n_835),
.Y(n_1339)
);

CKINVDCx16_ASAP7_75t_R g1340 ( 
.A(n_824),
.Y(n_1340)
);

CKINVDCx20_ASAP7_75t_R g1341 ( 
.A(n_893),
.Y(n_1341)
);

INVx1_ASAP7_75t_L g1342 ( 
.A(n_836),
.Y(n_1342)
);

BUFx3_ASAP7_75t_L g1343 ( 
.A(n_860),
.Y(n_1343)
);

INVx2_ASAP7_75t_L g1344 ( 
.A(n_912),
.Y(n_1344)
);

CKINVDCx20_ASAP7_75t_R g1345 ( 
.A(n_893),
.Y(n_1345)
);

INVxp67_ASAP7_75t_L g1346 ( 
.A(n_824),
.Y(n_1346)
);

HB1xp67_ASAP7_75t_L g1347 ( 
.A(n_894),
.Y(n_1347)
);

INVx2_ASAP7_75t_L g1348 ( 
.A(n_914),
.Y(n_1348)
);

INVx2_ASAP7_75t_L g1349 ( 
.A(n_914),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_949),
.Y(n_1350)
);

HB1xp67_ASAP7_75t_L g1351 ( 
.A(n_894),
.Y(n_1351)
);

CKINVDCx5p33_ASAP7_75t_R g1352 ( 
.A(n_899),
.Y(n_1352)
);

INVx1_ASAP7_75t_L g1353 ( 
.A(n_846),
.Y(n_1353)
);

INVx1_ASAP7_75t_L g1354 ( 
.A(n_847),
.Y(n_1354)
);

INVx1_ASAP7_75t_L g1355 ( 
.A(n_848),
.Y(n_1355)
);

INVx1_ASAP7_75t_L g1356 ( 
.A(n_949),
.Y(n_1356)
);

CKINVDCx5p33_ASAP7_75t_R g1357 ( 
.A(n_899),
.Y(n_1357)
);

INVx1_ASAP7_75t_L g1358 ( 
.A(n_850),
.Y(n_1358)
);

NOR2xp67_ASAP7_75t_L g1359 ( 
.A(n_903),
.B(n_708),
.Y(n_1359)
);

CKINVDCx5p33_ASAP7_75t_R g1360 ( 
.A(n_903),
.Y(n_1360)
);

INVxp67_ASAP7_75t_L g1361 ( 
.A(n_906),
.Y(n_1361)
);

INVx2_ASAP7_75t_L g1362 ( 
.A(n_967),
.Y(n_1362)
);

CKINVDCx20_ASAP7_75t_R g1363 ( 
.A(n_906),
.Y(n_1363)
);

INVxp33_ASAP7_75t_SL g1364 ( 
.A(n_913),
.Y(n_1364)
);

CKINVDCx20_ASAP7_75t_R g1365 ( 
.A(n_913),
.Y(n_1365)
);

CKINVDCx5p33_ASAP7_75t_R g1366 ( 
.A(n_916),
.Y(n_1366)
);

CKINVDCx20_ASAP7_75t_R g1367 ( 
.A(n_916),
.Y(n_1367)
);

INVx1_ASAP7_75t_L g1368 ( 
.A(n_851),
.Y(n_1368)
);

CKINVDCx5p33_ASAP7_75t_R g1369 ( 
.A(n_917),
.Y(n_1369)
);

NAND2xp5_ASAP7_75t_L g1370 ( 
.A(n_1037),
.B(n_904),
.Y(n_1370)
);

NOR2xp33_ASAP7_75t_L g1371 ( 
.A(n_917),
.B(n_710),
.Y(n_1371)
);

INVxp33_ASAP7_75t_SL g1372 ( 
.A(n_918),
.Y(n_1372)
);

INVxp67_ASAP7_75t_L g1373 ( 
.A(n_918),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_854),
.Y(n_1374)
);

BUFx3_ASAP7_75t_L g1375 ( 
.A(n_860),
.Y(n_1375)
);

CKINVDCx20_ASAP7_75t_R g1376 ( 
.A(n_921),
.Y(n_1376)
);

INVxp67_ASAP7_75t_SL g1377 ( 
.A(n_784),
.Y(n_1377)
);

INVx1_ASAP7_75t_L g1378 ( 
.A(n_857),
.Y(n_1378)
);

INVx1_ASAP7_75t_L g1379 ( 
.A(n_858),
.Y(n_1379)
);

CKINVDCx5p33_ASAP7_75t_R g1380 ( 
.A(n_921),
.Y(n_1380)
);

CKINVDCx20_ASAP7_75t_R g1381 ( 
.A(n_924),
.Y(n_1381)
);

CKINVDCx20_ASAP7_75t_R g1382 ( 
.A(n_924),
.Y(n_1382)
);

INVx1_ASAP7_75t_L g1383 ( 
.A(n_859),
.Y(n_1383)
);

CKINVDCx20_ASAP7_75t_R g1384 ( 
.A(n_928),
.Y(n_1384)
);

NOR2xp33_ASAP7_75t_L g1385 ( 
.A(n_928),
.B(n_715),
.Y(n_1385)
);

INVxp67_ASAP7_75t_SL g1386 ( 
.A(n_784),
.Y(n_1386)
);

NAND2xp5_ASAP7_75t_L g1387 ( 
.A(n_904),
.B(n_728),
.Y(n_1387)
);

INVx1_ASAP7_75t_L g1388 ( 
.A(n_863),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_864),
.Y(n_1389)
);

NAND2xp5_ASAP7_75t_L g1390 ( 
.A(n_904),
.B(n_729),
.Y(n_1390)
);

CKINVDCx5p33_ASAP7_75t_R g1391 ( 
.A(n_934),
.Y(n_1391)
);

INVx1_ASAP7_75t_L g1392 ( 
.A(n_865),
.Y(n_1392)
);

INVx1_ASAP7_75t_L g1393 ( 
.A(n_866),
.Y(n_1393)
);

CKINVDCx20_ASAP7_75t_R g1394 ( 
.A(n_934),
.Y(n_1394)
);

INVx1_ASAP7_75t_L g1395 ( 
.A(n_869),
.Y(n_1395)
);

CKINVDCx20_ASAP7_75t_R g1396 ( 
.A(n_941),
.Y(n_1396)
);

NOR2xp33_ASAP7_75t_L g1397 ( 
.A(n_941),
.B(n_756),
.Y(n_1397)
);

NAND2xp5_ASAP7_75t_L g1398 ( 
.A(n_904),
.B(n_759),
.Y(n_1398)
);

CKINVDCx20_ASAP7_75t_R g1399 ( 
.A(n_943),
.Y(n_1399)
);

INVx1_ASAP7_75t_L g1400 ( 
.A(n_872),
.Y(n_1400)
);

CKINVDCx5p33_ASAP7_75t_R g1401 ( 
.A(n_943),
.Y(n_1401)
);

CKINVDCx5p33_ASAP7_75t_R g1402 ( 
.A(n_945),
.Y(n_1402)
);

CKINVDCx5p33_ASAP7_75t_R g1403 ( 
.A(n_945),
.Y(n_1403)
);

CKINVDCx5p33_ASAP7_75t_R g1404 ( 
.A(n_950),
.Y(n_1404)
);

CKINVDCx5p33_ASAP7_75t_R g1405 ( 
.A(n_950),
.Y(n_1405)
);

CKINVDCx5p33_ASAP7_75t_R g1406 ( 
.A(n_952),
.Y(n_1406)
);

NAND2xp5_ASAP7_75t_L g1407 ( 
.A(n_904),
.B(n_498),
.Y(n_1407)
);

CKINVDCx5p33_ASAP7_75t_R g1408 ( 
.A(n_952),
.Y(n_1408)
);

INVxp67_ASAP7_75t_SL g1409 ( 
.A(n_784),
.Y(n_1409)
);

CKINVDCx5p33_ASAP7_75t_R g1410 ( 
.A(n_957),
.Y(n_1410)
);

INVxp67_ASAP7_75t_SL g1411 ( 
.A(n_834),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_883),
.Y(n_1412)
);

INVx1_ASAP7_75t_L g1413 ( 
.A(n_886),
.Y(n_1413)
);

CKINVDCx20_ASAP7_75t_R g1414 ( 
.A(n_957),
.Y(n_1414)
);

CKINVDCx5p33_ASAP7_75t_R g1415 ( 
.A(n_960),
.Y(n_1415)
);

CKINVDCx5p33_ASAP7_75t_R g1416 ( 
.A(n_960),
.Y(n_1416)
);

INVx1_ASAP7_75t_L g1417 ( 
.A(n_888),
.Y(n_1417)
);

INVx1_ASAP7_75t_L g1418 ( 
.A(n_890),
.Y(n_1418)
);

INVx1_ASAP7_75t_L g1419 ( 
.A(n_891),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_896),
.Y(n_1420)
);

INVx1_ASAP7_75t_L g1421 ( 
.A(n_897),
.Y(n_1421)
);

INVx1_ASAP7_75t_L g1422 ( 
.A(n_898),
.Y(n_1422)
);

INVx1_ASAP7_75t_L g1423 ( 
.A(n_905),
.Y(n_1423)
);

NOR2xp33_ASAP7_75t_L g1424 ( 
.A(n_962),
.B(n_691),
.Y(n_1424)
);

INVx1_ASAP7_75t_L g1425 ( 
.A(n_907),
.Y(n_1425)
);

INVxp67_ASAP7_75t_SL g1426 ( 
.A(n_834),
.Y(n_1426)
);

CKINVDCx5p33_ASAP7_75t_R g1427 ( 
.A(n_962),
.Y(n_1427)
);

CKINVDCx16_ASAP7_75t_R g1428 ( 
.A(n_1057),
.Y(n_1428)
);

INVx1_ASAP7_75t_L g1429 ( 
.A(n_908),
.Y(n_1429)
);

INVxp67_ASAP7_75t_SL g1430 ( 
.A(n_834),
.Y(n_1430)
);

NOR2xp67_ASAP7_75t_L g1431 ( 
.A(n_964),
.B(n_291),
.Y(n_1431)
);

NOR2xp33_ASAP7_75t_R g1432 ( 
.A(n_964),
.B(n_968),
.Y(n_1432)
);

NOR2xp33_ASAP7_75t_L g1433 ( 
.A(n_968),
.B(n_755),
.Y(n_1433)
);

CKINVDCx20_ASAP7_75t_R g1434 ( 
.A(n_969),
.Y(n_1434)
);

CKINVDCx20_ASAP7_75t_R g1435 ( 
.A(n_969),
.Y(n_1435)
);

CKINVDCx20_ASAP7_75t_R g1436 ( 
.A(n_976),
.Y(n_1436)
);

CKINVDCx16_ASAP7_75t_R g1437 ( 
.A(n_1076),
.Y(n_1437)
);

NAND2xp5_ASAP7_75t_L g1438 ( 
.A(n_904),
.B(n_787),
.Y(n_1438)
);

INVx2_ASAP7_75t_L g1439 ( 
.A(n_1212),
.Y(n_1439)
);

NOR2xp33_ASAP7_75t_L g1440 ( 
.A(n_1309),
.B(n_976),
.Y(n_1440)
);

INVx2_ASAP7_75t_L g1441 ( 
.A(n_1212),
.Y(n_1441)
);

INVx2_ASAP7_75t_L g1442 ( 
.A(n_1280),
.Y(n_1442)
);

INVx2_ASAP7_75t_L g1443 ( 
.A(n_1280),
.Y(n_1443)
);

INVx1_ASAP7_75t_L g1444 ( 
.A(n_1173),
.Y(n_1444)
);

BUFx2_ASAP7_75t_L g1445 ( 
.A(n_1246),
.Y(n_1445)
);

NAND2xp5_ASAP7_75t_L g1446 ( 
.A(n_1135),
.B(n_904),
.Y(n_1446)
);

INVx1_ASAP7_75t_L g1447 ( 
.A(n_1175),
.Y(n_1447)
);

INVx2_ASAP7_75t_L g1448 ( 
.A(n_1304),
.Y(n_1448)
);

BUFx6f_ASAP7_75t_L g1449 ( 
.A(n_1204),
.Y(n_1449)
);

BUFx6f_ASAP7_75t_L g1450 ( 
.A(n_1204),
.Y(n_1450)
);

OA21x2_ASAP7_75t_L g1451 ( 
.A1(n_1176),
.A2(n_774),
.B(n_773),
.Y(n_1451)
);

OAI22xp5_ASAP7_75t_SL g1452 ( 
.A1(n_1297),
.A2(n_1036),
.B1(n_664),
.B2(n_692),
.Y(n_1452)
);

BUFx6f_ASAP7_75t_L g1453 ( 
.A(n_1204),
.Y(n_1453)
);

AOI22xp5_ASAP7_75t_SL g1454 ( 
.A1(n_1247),
.A2(n_1036),
.B1(n_760),
.B2(n_709),
.Y(n_1454)
);

INVx3_ASAP7_75t_L g1455 ( 
.A(n_1304),
.Y(n_1455)
);

INVx3_ASAP7_75t_L g1456 ( 
.A(n_1344),
.Y(n_1456)
);

BUFx3_ASAP7_75t_L g1457 ( 
.A(n_1141),
.Y(n_1457)
);

INVx5_ASAP7_75t_L g1458 ( 
.A(n_1344),
.Y(n_1458)
);

BUFx3_ASAP7_75t_L g1459 ( 
.A(n_1143),
.Y(n_1459)
);

NOR2xp33_ASAP7_75t_L g1460 ( 
.A(n_1371),
.B(n_978),
.Y(n_1460)
);

CKINVDCx20_ASAP7_75t_R g1461 ( 
.A(n_1138),
.Y(n_1461)
);

OA21x2_ASAP7_75t_L g1462 ( 
.A1(n_1180),
.A2(n_778),
.B(n_776),
.Y(n_1462)
);

INVx2_ASAP7_75t_L g1463 ( 
.A(n_1348),
.Y(n_1463)
);

OAI22x1_ASAP7_75t_R g1464 ( 
.A1(n_1221),
.A2(n_712),
.B1(n_716),
.B2(n_663),
.Y(n_1464)
);

BUFx6f_ASAP7_75t_L g1465 ( 
.A(n_1348),
.Y(n_1465)
);

INVx1_ASAP7_75t_L g1466 ( 
.A(n_1181),
.Y(n_1466)
);

BUFx8_ASAP7_75t_L g1467 ( 
.A(n_1295),
.Y(n_1467)
);

INVx2_ASAP7_75t_L g1468 ( 
.A(n_1349),
.Y(n_1468)
);

AND2x2_ASAP7_75t_L g1469 ( 
.A(n_1332),
.B(n_909),
.Y(n_1469)
);

CKINVDCx20_ASAP7_75t_R g1470 ( 
.A(n_1146),
.Y(n_1470)
);

OAI22xp5_ASAP7_75t_L g1471 ( 
.A1(n_1332),
.A2(n_1097),
.B1(n_944),
.B2(n_987),
.Y(n_1471)
);

AOI22xp5_ASAP7_75t_L g1472 ( 
.A1(n_1136),
.A2(n_741),
.B1(n_758),
.B2(n_722),
.Y(n_1472)
);

INVx2_ASAP7_75t_L g1473 ( 
.A(n_1349),
.Y(n_1473)
);

OA21x2_ASAP7_75t_L g1474 ( 
.A1(n_1182),
.A2(n_782),
.B(n_780),
.Y(n_1474)
);

INVx2_ASAP7_75t_SL g1475 ( 
.A(n_1328),
.Y(n_1475)
);

AND2x4_ASAP7_75t_L g1476 ( 
.A(n_1201),
.B(n_1047),
.Y(n_1476)
);

INVx1_ASAP7_75t_L g1477 ( 
.A(n_1186),
.Y(n_1477)
);

BUFx6f_ASAP7_75t_L g1478 ( 
.A(n_1362),
.Y(n_1478)
);

INVx2_ASAP7_75t_L g1479 ( 
.A(n_1362),
.Y(n_1479)
);

INVx5_ASAP7_75t_L g1480 ( 
.A(n_1343),
.Y(n_1480)
);

INVx2_ASAP7_75t_L g1481 ( 
.A(n_1202),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_1187),
.Y(n_1482)
);

NOR2xp33_ASAP7_75t_L g1483 ( 
.A(n_1385),
.B(n_978),
.Y(n_1483)
);

NAND2xp5_ASAP7_75t_SL g1484 ( 
.A(n_1437),
.B(n_987),
.Y(n_1484)
);

AND2x4_ASAP7_75t_L g1485 ( 
.A(n_1222),
.B(n_1047),
.Y(n_1485)
);

INVx1_ASAP7_75t_L g1486 ( 
.A(n_1188),
.Y(n_1486)
);

NAND2x1p5_ASAP7_75t_L g1487 ( 
.A(n_1431),
.B(n_911),
.Y(n_1487)
);

INVx1_ASAP7_75t_L g1488 ( 
.A(n_1189),
.Y(n_1488)
);

INVx3_ASAP7_75t_L g1489 ( 
.A(n_1202),
.Y(n_1489)
);

OAI22xp5_ASAP7_75t_L g1490 ( 
.A1(n_1338),
.A2(n_1289),
.B1(n_1291),
.B2(n_1276),
.Y(n_1490)
);

OAI21x1_ASAP7_75t_L g1491 ( 
.A1(n_1370),
.A2(n_788),
.B(n_785),
.Y(n_1491)
);

INVx2_ASAP7_75t_SL g1492 ( 
.A(n_1328),
.Y(n_1492)
);

INVx1_ASAP7_75t_L g1493 ( 
.A(n_1191),
.Y(n_1493)
);

INVx4_ASAP7_75t_L g1494 ( 
.A(n_1343),
.Y(n_1494)
);

INVxp67_ASAP7_75t_L g1495 ( 
.A(n_1244),
.Y(n_1495)
);

INVx1_ASAP7_75t_L g1496 ( 
.A(n_1192),
.Y(n_1496)
);

BUFx6f_ASAP7_75t_L g1497 ( 
.A(n_1195),
.Y(n_1497)
);

NAND2xp5_ASAP7_75t_L g1498 ( 
.A(n_1230),
.B(n_904),
.Y(n_1498)
);

OAI21x1_ASAP7_75t_L g1499 ( 
.A1(n_1387),
.A2(n_1004),
.B(n_967),
.Y(n_1499)
);

INVx1_ASAP7_75t_L g1500 ( 
.A(n_1199),
.Y(n_1500)
);

INVx1_ASAP7_75t_L g1501 ( 
.A(n_1147),
.Y(n_1501)
);

INVx2_ASAP7_75t_L g1502 ( 
.A(n_1203),
.Y(n_1502)
);

AND2x4_ASAP7_75t_L g1503 ( 
.A(n_1223),
.B(n_948),
.Y(n_1503)
);

AND2x2_ASAP7_75t_SL g1504 ( 
.A(n_1407),
.B(n_1069),
.Y(n_1504)
);

NOR2xp33_ASAP7_75t_L g1505 ( 
.A(n_1397),
.B(n_988),
.Y(n_1505)
);

CKINVDCx20_ASAP7_75t_R g1506 ( 
.A(n_1162),
.Y(n_1506)
);

INVx1_ASAP7_75t_L g1507 ( 
.A(n_1149),
.Y(n_1507)
);

INVx1_ASAP7_75t_L g1508 ( 
.A(n_1151),
.Y(n_1508)
);

NAND2xp5_ASAP7_75t_L g1509 ( 
.A(n_1239),
.B(n_1249),
.Y(n_1509)
);

INVx2_ASAP7_75t_L g1510 ( 
.A(n_1203),
.Y(n_1510)
);

INVx3_ASAP7_75t_L g1511 ( 
.A(n_1207),
.Y(n_1511)
);

INVx1_ASAP7_75t_L g1512 ( 
.A(n_1152),
.Y(n_1512)
);

AND2x6_ASAP7_75t_L g1513 ( 
.A(n_1390),
.B(n_472),
.Y(n_1513)
);

INVx3_ASAP7_75t_L g1514 ( 
.A(n_1207),
.Y(n_1514)
);

BUFx6f_ASAP7_75t_L g1515 ( 
.A(n_1153),
.Y(n_1515)
);

CKINVDCx8_ASAP7_75t_R g1516 ( 
.A(n_1142),
.Y(n_1516)
);

AND2x6_ASAP7_75t_L g1517 ( 
.A(n_1398),
.B(n_487),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_1157),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_1158),
.Y(n_1519)
);

NOR2xp33_ASAP7_75t_L g1520 ( 
.A(n_1217),
.B(n_991),
.Y(n_1520)
);

AND2x2_ASAP7_75t_L g1521 ( 
.A(n_1225),
.B(n_1045),
.Y(n_1521)
);

AND2x4_ASAP7_75t_L g1522 ( 
.A(n_1228),
.B(n_951),
.Y(n_1522)
);

INVxp67_ASAP7_75t_L g1523 ( 
.A(n_1295),
.Y(n_1523)
);

INVx1_ASAP7_75t_L g1524 ( 
.A(n_1438),
.Y(n_1524)
);

INVx2_ASAP7_75t_L g1525 ( 
.A(n_1213),
.Y(n_1525)
);

AND2x2_ASAP7_75t_L g1526 ( 
.A(n_1234),
.B(n_1045),
.Y(n_1526)
);

AND2x4_ASAP7_75t_L g1527 ( 
.A(n_1235),
.B(n_1236),
.Y(n_1527)
);

NOR2x1_ASAP7_75t_L g1528 ( 
.A(n_1375),
.B(n_498),
.Y(n_1528)
);

BUFx6f_ASAP7_75t_L g1529 ( 
.A(n_1213),
.Y(n_1529)
);

INVx2_ASAP7_75t_L g1530 ( 
.A(n_1215),
.Y(n_1530)
);

AND2x4_ASAP7_75t_L g1531 ( 
.A(n_1237),
.B(n_954),
.Y(n_1531)
);

INVx1_ASAP7_75t_L g1532 ( 
.A(n_1254),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_1255),
.Y(n_1533)
);

NOR2xp33_ASAP7_75t_L g1534 ( 
.A(n_1219),
.B(n_991),
.Y(n_1534)
);

BUFx6f_ASAP7_75t_L g1535 ( 
.A(n_1215),
.Y(n_1535)
);

INVx2_ASAP7_75t_L g1536 ( 
.A(n_1216),
.Y(n_1536)
);

INVx1_ASAP7_75t_L g1537 ( 
.A(n_1260),
.Y(n_1537)
);

INVx1_ASAP7_75t_L g1538 ( 
.A(n_1263),
.Y(n_1538)
);

INVx1_ASAP7_75t_L g1539 ( 
.A(n_1266),
.Y(n_1539)
);

NAND2xp33_ASAP7_75t_L g1540 ( 
.A(n_1274),
.B(n_992),
.Y(n_1540)
);

INVx2_ASAP7_75t_L g1541 ( 
.A(n_1216),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_1272),
.Y(n_1542)
);

BUFx6f_ASAP7_75t_L g1543 ( 
.A(n_1218),
.Y(n_1543)
);

BUFx2_ASAP7_75t_L g1544 ( 
.A(n_1252),
.Y(n_1544)
);

OAI22xp5_ASAP7_75t_SL g1545 ( 
.A1(n_1325),
.A2(n_512),
.B1(n_536),
.B2(n_480),
.Y(n_1545)
);

BUFx12f_ASAP7_75t_L g1546 ( 
.A(n_1214),
.Y(n_1546)
);

INVx1_ASAP7_75t_L g1547 ( 
.A(n_1277),
.Y(n_1547)
);

NAND2xp5_ASAP7_75t_L g1548 ( 
.A(n_1144),
.B(n_1154),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_1282),
.Y(n_1549)
);

INVx2_ASAP7_75t_L g1550 ( 
.A(n_1218),
.Y(n_1550)
);

BUFx6f_ASAP7_75t_L g1551 ( 
.A(n_1220),
.Y(n_1551)
);

INVx2_ASAP7_75t_L g1552 ( 
.A(n_1220),
.Y(n_1552)
);

INVx1_ASAP7_75t_L g1553 ( 
.A(n_1293),
.Y(n_1553)
);

INVx2_ASAP7_75t_L g1554 ( 
.A(n_1233),
.Y(n_1554)
);

NAND2xp5_ASAP7_75t_L g1555 ( 
.A(n_1165),
.B(n_1004),
.Y(n_1555)
);

INVx1_ASAP7_75t_L g1556 ( 
.A(n_1294),
.Y(n_1556)
);

OAI22xp5_ASAP7_75t_L g1557 ( 
.A1(n_1319),
.A2(n_994),
.B1(n_996),
.B2(n_992),
.Y(n_1557)
);

BUFx2_ASAP7_75t_L g1558 ( 
.A(n_1335),
.Y(n_1558)
);

INVx2_ASAP7_75t_L g1559 ( 
.A(n_1233),
.Y(n_1559)
);

INVx1_ASAP7_75t_L g1560 ( 
.A(n_1298),
.Y(n_1560)
);

INVx1_ASAP7_75t_L g1561 ( 
.A(n_1299),
.Y(n_1561)
);

INVx2_ASAP7_75t_L g1562 ( 
.A(n_1323),
.Y(n_1562)
);

INVx1_ASAP7_75t_L g1563 ( 
.A(n_1300),
.Y(n_1563)
);

NAND2xp5_ASAP7_75t_L g1564 ( 
.A(n_1163),
.B(n_996),
.Y(n_1564)
);

INVx2_ASAP7_75t_L g1565 ( 
.A(n_1323),
.Y(n_1565)
);

AND2x6_ASAP7_75t_L g1566 ( 
.A(n_1424),
.B(n_487),
.Y(n_1566)
);

INVx2_ASAP7_75t_L g1567 ( 
.A(n_1327),
.Y(n_1567)
);

INVx2_ASAP7_75t_L g1568 ( 
.A(n_1327),
.Y(n_1568)
);

OAI22xp5_ASAP7_75t_L g1569 ( 
.A1(n_1140),
.A2(n_998),
.B1(n_999),
.B2(n_997),
.Y(n_1569)
);

NAND2xp5_ASAP7_75t_L g1570 ( 
.A(n_1164),
.B(n_997),
.Y(n_1570)
);

NOR2x1_ASAP7_75t_L g1571 ( 
.A(n_1375),
.B(n_1069),
.Y(n_1571)
);

CKINVDCx20_ASAP7_75t_R g1572 ( 
.A(n_1169),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_1301),
.Y(n_1573)
);

BUFx6f_ASAP7_75t_L g1574 ( 
.A(n_1329),
.Y(n_1574)
);

INVx3_ASAP7_75t_L g1575 ( 
.A(n_1329),
.Y(n_1575)
);

HB1xp67_ASAP7_75t_L g1576 ( 
.A(n_1320),
.Y(n_1576)
);

HB1xp67_ASAP7_75t_L g1577 ( 
.A(n_1324),
.Y(n_1577)
);

AND2x2_ASAP7_75t_L g1578 ( 
.A(n_1241),
.B(n_1058),
.Y(n_1578)
);

OA21x2_ASAP7_75t_L g1579 ( 
.A1(n_1350),
.A2(n_959),
.B(n_958),
.Y(n_1579)
);

OA21x2_ASAP7_75t_L g1580 ( 
.A1(n_1350),
.A2(n_971),
.B(n_966),
.Y(n_1580)
);

BUFx8_ASAP7_75t_L g1581 ( 
.A(n_1321),
.Y(n_1581)
);

INVx2_ASAP7_75t_L g1582 ( 
.A(n_1356),
.Y(n_1582)
);

INVx3_ASAP7_75t_L g1583 ( 
.A(n_1356),
.Y(n_1583)
);

OAI21x1_ASAP7_75t_L g1584 ( 
.A1(n_1308),
.A2(n_979),
.B(n_972),
.Y(n_1584)
);

BUFx2_ASAP7_75t_L g1585 ( 
.A(n_1340),
.Y(n_1585)
);

NOR2x1_ASAP7_75t_L g1586 ( 
.A(n_1256),
.B(n_980),
.Y(n_1586)
);

CKINVDCx5p33_ASAP7_75t_R g1587 ( 
.A(n_1139),
.Y(n_1587)
);

INVx2_ASAP7_75t_L g1588 ( 
.A(n_1302),
.Y(n_1588)
);

HB1xp67_ASAP7_75t_L g1589 ( 
.A(n_1333),
.Y(n_1589)
);

INVx1_ASAP7_75t_L g1590 ( 
.A(n_1303),
.Y(n_1590)
);

CKINVDCx20_ASAP7_75t_R g1591 ( 
.A(n_1172),
.Y(n_1591)
);

BUFx6f_ASAP7_75t_L g1592 ( 
.A(n_1313),
.Y(n_1592)
);

OAI22x1_ASAP7_75t_SL g1593 ( 
.A1(n_1224),
.A2(n_565),
.B1(n_566),
.B2(n_559),
.Y(n_1593)
);

BUFx6f_ASAP7_75t_L g1594 ( 
.A(n_1315),
.Y(n_1594)
);

AND2x4_ASAP7_75t_L g1595 ( 
.A(n_1243),
.B(n_981),
.Y(n_1595)
);

INVx2_ASAP7_75t_L g1596 ( 
.A(n_1316),
.Y(n_1596)
);

INVx2_ASAP7_75t_L g1597 ( 
.A(n_1317),
.Y(n_1597)
);

OA21x2_ASAP7_75t_L g1598 ( 
.A1(n_1322),
.A2(n_985),
.B(n_982),
.Y(n_1598)
);

INVx6_ASAP7_75t_L g1599 ( 
.A(n_1321),
.Y(n_1599)
);

INVxp67_ASAP7_75t_L g1600 ( 
.A(n_1250),
.Y(n_1600)
);

INVx1_ASAP7_75t_L g1601 ( 
.A(n_1339),
.Y(n_1601)
);

INVx2_ASAP7_75t_L g1602 ( 
.A(n_1342),
.Y(n_1602)
);

OAI22xp5_ASAP7_75t_SL g1603 ( 
.A1(n_1231),
.A2(n_679),
.B1(n_727),
.B2(n_628),
.Y(n_1603)
);

AND2x4_ASAP7_75t_L g1604 ( 
.A(n_1251),
.B(n_986),
.Y(n_1604)
);

HB1xp67_ASAP7_75t_L g1605 ( 
.A(n_1346),
.Y(n_1605)
);

INVx1_ASAP7_75t_L g1606 ( 
.A(n_1353),
.Y(n_1606)
);

INVx2_ASAP7_75t_L g1607 ( 
.A(n_1354),
.Y(n_1607)
);

NOR2xp33_ASAP7_75t_SL g1608 ( 
.A(n_1428),
.B(n_998),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_1355),
.Y(n_1609)
);

NAND2xp5_ASAP7_75t_L g1610 ( 
.A(n_1171),
.B(n_999),
.Y(n_1610)
);

BUFx3_ASAP7_75t_L g1611 ( 
.A(n_1358),
.Y(n_1611)
);

INVx1_ASAP7_75t_L g1612 ( 
.A(n_1368),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1374),
.Y(n_1613)
);

INVx1_ASAP7_75t_L g1614 ( 
.A(n_1378),
.Y(n_1614)
);

INVx2_ASAP7_75t_L g1615 ( 
.A(n_1379),
.Y(n_1615)
);

AOI22xp5_ASAP7_75t_L g1616 ( 
.A1(n_1433),
.A2(n_874),
.B1(n_955),
.B2(n_856),
.Y(n_1616)
);

BUFx6f_ASAP7_75t_L g1617 ( 
.A(n_1383),
.Y(n_1617)
);

INVx3_ASAP7_75t_L g1618 ( 
.A(n_1388),
.Y(n_1618)
);

AND2x2_ASAP7_75t_L g1619 ( 
.A(n_1389),
.B(n_1058),
.Y(n_1619)
);

INVx3_ASAP7_75t_L g1620 ( 
.A(n_1392),
.Y(n_1620)
);

AND2x4_ASAP7_75t_L g1621 ( 
.A(n_1197),
.B(n_1003),
.Y(n_1621)
);

OAI21x1_ASAP7_75t_L g1622 ( 
.A1(n_1393),
.A2(n_1006),
.B(n_1005),
.Y(n_1622)
);

CKINVDCx20_ASAP7_75t_R g1623 ( 
.A(n_1177),
.Y(n_1623)
);

INVx2_ASAP7_75t_SL g1624 ( 
.A(n_1137),
.Y(n_1624)
);

INVx1_ASAP7_75t_L g1625 ( 
.A(n_1395),
.Y(n_1625)
);

AND2x4_ASAP7_75t_L g1626 ( 
.A(n_1400),
.B(n_1007),
.Y(n_1626)
);

INVx1_ASAP7_75t_L g1627 ( 
.A(n_1412),
.Y(n_1627)
);

NAND2xp5_ASAP7_75t_L g1628 ( 
.A(n_1267),
.B(n_1000),
.Y(n_1628)
);

INVx2_ASAP7_75t_L g1629 ( 
.A(n_1413),
.Y(n_1629)
);

BUFx3_ASAP7_75t_L g1630 ( 
.A(n_1417),
.Y(n_1630)
);

AND2x4_ASAP7_75t_L g1631 ( 
.A(n_1418),
.B(n_1008),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_1419),
.Y(n_1632)
);

INVx1_ASAP7_75t_SL g1633 ( 
.A(n_1292),
.Y(n_1633)
);

OA21x2_ASAP7_75t_L g1634 ( 
.A1(n_1420),
.A2(n_1021),
.B(n_1020),
.Y(n_1634)
);

INVx2_ASAP7_75t_L g1635 ( 
.A(n_1421),
.Y(n_1635)
);

NAND2xp5_ASAP7_75t_L g1636 ( 
.A(n_1336),
.B(n_1000),
.Y(n_1636)
);

INVx2_ASAP7_75t_L g1637 ( 
.A(n_1422),
.Y(n_1637)
);

INVx1_ASAP7_75t_L g1638 ( 
.A(n_1423),
.Y(n_1638)
);

INVx2_ASAP7_75t_L g1639 ( 
.A(n_1425),
.Y(n_1639)
);

INVx3_ASAP7_75t_L g1640 ( 
.A(n_1429),
.Y(n_1640)
);

INVx2_ASAP7_75t_L g1641 ( 
.A(n_1377),
.Y(n_1641)
);

INVx2_ASAP7_75t_L g1642 ( 
.A(n_1386),
.Y(n_1642)
);

INVx2_ASAP7_75t_SL g1643 ( 
.A(n_1150),
.Y(n_1643)
);

INVx2_ASAP7_75t_L g1644 ( 
.A(n_1409),
.Y(n_1644)
);

INVx4_ASAP7_75t_L g1645 ( 
.A(n_1214),
.Y(n_1645)
);

BUFx6f_ASAP7_75t_L g1646 ( 
.A(n_1242),
.Y(n_1646)
);

INVx1_ASAP7_75t_L g1647 ( 
.A(n_1411),
.Y(n_1647)
);

BUFx3_ASAP7_75t_L g1648 ( 
.A(n_1310),
.Y(n_1648)
);

INVx2_ASAP7_75t_SL g1649 ( 
.A(n_1288),
.Y(n_1649)
);

INVx1_ASAP7_75t_L g1650 ( 
.A(n_1426),
.Y(n_1650)
);

INVx2_ASAP7_75t_L g1651 ( 
.A(n_1430),
.Y(n_1651)
);

AND2x2_ASAP7_75t_L g1652 ( 
.A(n_1284),
.B(n_1120),
.Y(n_1652)
);

NAND2xp5_ASAP7_75t_L g1653 ( 
.A(n_1359),
.B(n_1001),
.Y(n_1653)
);

INVx1_ASAP7_75t_L g1654 ( 
.A(n_1166),
.Y(n_1654)
);

INVx1_ASAP7_75t_L g1655 ( 
.A(n_1208),
.Y(n_1655)
);

AND2x2_ASAP7_75t_L g1656 ( 
.A(n_1145),
.B(n_1120),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1361),
.Y(n_1657)
);

INVx1_ASAP7_75t_L g1658 ( 
.A(n_1373),
.Y(n_1658)
);

INVx2_ASAP7_75t_L g1659 ( 
.A(n_1330),
.Y(n_1659)
);

INVx3_ASAP7_75t_L g1660 ( 
.A(n_1205),
.Y(n_1660)
);

BUFx6f_ASAP7_75t_L g1661 ( 
.A(n_1314),
.Y(n_1661)
);

AND2x2_ASAP7_75t_L g1662 ( 
.A(n_1259),
.B(n_1079),
.Y(n_1662)
);

OAI22xp5_ASAP7_75t_SL g1663 ( 
.A1(n_1240),
.A2(n_812),
.B1(n_566),
.B2(n_567),
.Y(n_1663)
);

INVx1_ASAP7_75t_L g1664 ( 
.A(n_1347),
.Y(n_1664)
);

BUFx2_ASAP7_75t_L g1665 ( 
.A(n_1245),
.Y(n_1665)
);

INVx4_ASAP7_75t_L g1666 ( 
.A(n_1227),
.Y(n_1666)
);

INVx2_ASAP7_75t_L g1667 ( 
.A(n_1351),
.Y(n_1667)
);

OA21x2_ASAP7_75t_L g1668 ( 
.A1(n_1227),
.A2(n_1042),
.B(n_1038),
.Y(n_1668)
);

NAND2xp5_ASAP7_75t_L g1669 ( 
.A(n_1326),
.B(n_1001),
.Y(n_1669)
);

AND2x4_ASAP7_75t_L g1670 ( 
.A(n_1229),
.B(n_1079),
.Y(n_1670)
);

BUFx12f_ASAP7_75t_L g1671 ( 
.A(n_1229),
.Y(n_1671)
);

OAI22xp5_ASAP7_75t_L g1672 ( 
.A1(n_1326),
.A2(n_1010),
.B1(n_1011),
.B2(n_1002),
.Y(n_1672)
);

OA21x2_ASAP7_75t_L g1673 ( 
.A1(n_1232),
.A2(n_1049),
.B(n_1044),
.Y(n_1673)
);

OA21x2_ASAP7_75t_L g1674 ( 
.A1(n_1232),
.A2(n_1051),
.B(n_1050),
.Y(n_1674)
);

INVx2_ASAP7_75t_L g1675 ( 
.A(n_1238),
.Y(n_1675)
);

INVx2_ASAP7_75t_L g1676 ( 
.A(n_1238),
.Y(n_1676)
);

INVx3_ASAP7_75t_L g1677 ( 
.A(n_1248),
.Y(n_1677)
);

AND2x4_ASAP7_75t_L g1678 ( 
.A(n_1248),
.B(n_1079),
.Y(n_1678)
);

INVx1_ASAP7_75t_L g1679 ( 
.A(n_1432),
.Y(n_1679)
);

BUFx6f_ASAP7_75t_L g1680 ( 
.A(n_1253),
.Y(n_1680)
);

BUFx2_ASAP7_75t_L g1681 ( 
.A(n_1261),
.Y(n_1681)
);

AND2x4_ASAP7_75t_L g1682 ( 
.A(n_1253),
.B(n_1056),
.Y(n_1682)
);

AND2x2_ASAP7_75t_L g1683 ( 
.A(n_1257),
.B(n_956),
.Y(n_1683)
);

AND2x6_ASAP7_75t_L g1684 ( 
.A(n_1364),
.B(n_487),
.Y(n_1684)
);

BUFx6f_ASAP7_75t_L g1685 ( 
.A(n_1257),
.Y(n_1685)
);

INVx5_ASAP7_75t_L g1686 ( 
.A(n_1287),
.Y(n_1686)
);

NAND2xp5_ASAP7_75t_SL g1687 ( 
.A(n_1364),
.B(n_1002),
.Y(n_1687)
);

INVx3_ASAP7_75t_L g1688 ( 
.A(n_1258),
.Y(n_1688)
);

NAND2xp5_ASAP7_75t_L g1689 ( 
.A(n_1372),
.B(n_1010),
.Y(n_1689)
);

INVx1_ASAP7_75t_L g1690 ( 
.A(n_1258),
.Y(n_1690)
);

INVx1_ASAP7_75t_L g1691 ( 
.A(n_1262),
.Y(n_1691)
);

INVx1_ASAP7_75t_L g1692 ( 
.A(n_1262),
.Y(n_1692)
);

INVx1_ASAP7_75t_L g1693 ( 
.A(n_1265),
.Y(n_1693)
);

AND2x6_ASAP7_75t_L g1694 ( 
.A(n_1372),
.B(n_499),
.Y(n_1694)
);

INVx2_ASAP7_75t_L g1695 ( 
.A(n_1265),
.Y(n_1695)
);

INVx2_ASAP7_75t_L g1696 ( 
.A(n_1271),
.Y(n_1696)
);

INVx3_ASAP7_75t_L g1697 ( 
.A(n_1271),
.Y(n_1697)
);

BUFx3_ASAP7_75t_L g1698 ( 
.A(n_1273),
.Y(n_1698)
);

INVx2_ASAP7_75t_L g1699 ( 
.A(n_1273),
.Y(n_1699)
);

INVx1_ASAP7_75t_L g1700 ( 
.A(n_1275),
.Y(n_1700)
);

BUFx2_ASAP7_75t_L g1701 ( 
.A(n_1296),
.Y(n_1701)
);

BUFx2_ASAP7_75t_L g1702 ( 
.A(n_1306),
.Y(n_1702)
);

INVx2_ASAP7_75t_L g1703 ( 
.A(n_1275),
.Y(n_1703)
);

HB1xp67_ASAP7_75t_L g1704 ( 
.A(n_1224),
.Y(n_1704)
);

BUFx6f_ASAP7_75t_L g1705 ( 
.A(n_1278),
.Y(n_1705)
);

AND2x4_ASAP7_75t_L g1706 ( 
.A(n_1278),
.B(n_1059),
.Y(n_1706)
);

AND2x6_ASAP7_75t_L g1707 ( 
.A(n_1226),
.B(n_499),
.Y(n_1707)
);

NAND2xp5_ASAP7_75t_L g1708 ( 
.A(n_1279),
.B(n_1011),
.Y(n_1708)
);

INVx2_ASAP7_75t_L g1709 ( 
.A(n_1279),
.Y(n_1709)
);

INVx2_ASAP7_75t_L g1710 ( 
.A(n_1285),
.Y(n_1710)
);

NOR2xp33_ASAP7_75t_SL g1711 ( 
.A(n_1170),
.B(n_1014),
.Y(n_1711)
);

INVx2_ASAP7_75t_L g1712 ( 
.A(n_1285),
.Y(n_1712)
);

OA21x2_ASAP7_75t_L g1713 ( 
.A1(n_1290),
.A2(n_1065),
.B(n_1060),
.Y(n_1713)
);

CKINVDCx5p33_ASAP7_75t_R g1714 ( 
.A(n_1139),
.Y(n_1714)
);

INVx2_ASAP7_75t_L g1715 ( 
.A(n_1290),
.Y(n_1715)
);

CKINVDCx5p33_ASAP7_75t_R g1716 ( 
.A(n_1148),
.Y(n_1716)
);

INVx3_ASAP7_75t_L g1717 ( 
.A(n_1305),
.Y(n_1717)
);

INVx1_ASAP7_75t_L g1718 ( 
.A(n_1305),
.Y(n_1718)
);

INVx3_ASAP7_75t_L g1719 ( 
.A(n_1307),
.Y(n_1719)
);

AND2x2_ASAP7_75t_L g1720 ( 
.A(n_1307),
.B(n_989),
.Y(n_1720)
);

AND2x4_ASAP7_75t_L g1721 ( 
.A(n_1311),
.B(n_1068),
.Y(n_1721)
);

AND2x2_ASAP7_75t_L g1722 ( 
.A(n_1311),
.B(n_1070),
.Y(n_1722)
);

INVx5_ASAP7_75t_L g1723 ( 
.A(n_1226),
.Y(n_1723)
);

AND2x2_ASAP7_75t_L g1724 ( 
.A(n_1495),
.B(n_1683),
.Y(n_1724)
);

AND2x2_ASAP7_75t_L g1725 ( 
.A(n_1683),
.B(n_1312),
.Y(n_1725)
);

INVx4_ASAP7_75t_L g1726 ( 
.A(n_1592),
.Y(n_1726)
);

INVx1_ASAP7_75t_L g1727 ( 
.A(n_1489),
.Y(n_1727)
);

INVx1_ASAP7_75t_L g1728 ( 
.A(n_1489),
.Y(n_1728)
);

NOR2xp33_ASAP7_75t_L g1729 ( 
.A(n_1600),
.B(n_1548),
.Y(n_1729)
);

AOI22xp5_ASAP7_75t_L g1730 ( 
.A1(n_1504),
.A2(n_1318),
.B1(n_1334),
.B2(n_1312),
.Y(n_1730)
);

AND2x2_ASAP7_75t_L g1731 ( 
.A(n_1720),
.B(n_1318),
.Y(n_1731)
);

BUFx6f_ASAP7_75t_L g1732 ( 
.A(n_1611),
.Y(n_1732)
);

AO22x2_ASAP7_75t_L g1733 ( 
.A1(n_1490),
.A2(n_755),
.B1(n_567),
.B2(n_577),
.Y(n_1733)
);

NOR2xp33_ASAP7_75t_L g1734 ( 
.A(n_1440),
.B(n_1334),
.Y(n_1734)
);

INVx2_ASAP7_75t_L g1735 ( 
.A(n_1455),
.Y(n_1735)
);

OR2x6_ASAP7_75t_L g1736 ( 
.A(n_1445),
.B(n_817),
.Y(n_1736)
);

AND2x2_ASAP7_75t_SL g1737 ( 
.A(n_1558),
.B(n_499),
.Y(n_1737)
);

AND2x2_ASAP7_75t_L g1738 ( 
.A(n_1720),
.B(n_1352),
.Y(n_1738)
);

OR2x6_ASAP7_75t_L g1739 ( 
.A(n_1445),
.B(n_817),
.Y(n_1739)
);

INVx2_ASAP7_75t_L g1740 ( 
.A(n_1455),
.Y(n_1740)
);

OAI22xp33_ASAP7_75t_SL g1741 ( 
.A1(n_1599),
.A2(n_1628),
.B1(n_1570),
.B2(n_1610),
.Y(n_1741)
);

AOI22xp5_ASAP7_75t_L g1742 ( 
.A1(n_1504),
.A2(n_1357),
.B1(n_1360),
.B2(n_1352),
.Y(n_1742)
);

AO22x2_ASAP7_75t_L g1743 ( 
.A1(n_1557),
.A2(n_565),
.B1(n_581),
.B2(n_577),
.Y(n_1743)
);

INVx1_ASAP7_75t_L g1744 ( 
.A(n_1489),
.Y(n_1744)
);

AO22x2_ASAP7_75t_L g1745 ( 
.A1(n_1475),
.A2(n_581),
.B1(n_589),
.B2(n_585),
.Y(n_1745)
);

OAI22xp33_ASAP7_75t_R g1746 ( 
.A1(n_1464),
.A2(n_1454),
.B1(n_1452),
.B2(n_1460),
.Y(n_1746)
);

AND2x2_ASAP7_75t_L g1747 ( 
.A(n_1475),
.B(n_1357),
.Y(n_1747)
);

NOR2xp33_ASAP7_75t_L g1748 ( 
.A(n_1483),
.B(n_1360),
.Y(n_1748)
);

AOI22xp5_ASAP7_75t_L g1749 ( 
.A1(n_1504),
.A2(n_1369),
.B1(n_1380),
.B2(n_1366),
.Y(n_1749)
);

OAI22xp33_ASAP7_75t_L g1750 ( 
.A1(n_1492),
.A2(n_1369),
.B1(n_1380),
.B2(n_1366),
.Y(n_1750)
);

AOI22xp5_ASAP7_75t_L g1751 ( 
.A1(n_1566),
.A2(n_1401),
.B1(n_1402),
.B2(n_1391),
.Y(n_1751)
);

AO22x2_ASAP7_75t_L g1752 ( 
.A1(n_1492),
.A2(n_585),
.B1(n_593),
.B2(n_589),
.Y(n_1752)
);

OR2x6_ASAP7_75t_L g1753 ( 
.A(n_1544),
.B(n_965),
.Y(n_1753)
);

AO22x2_ASAP7_75t_L g1754 ( 
.A1(n_1569),
.A2(n_593),
.B1(n_599),
.B2(n_597),
.Y(n_1754)
);

INVx1_ASAP7_75t_L g1755 ( 
.A(n_1489),
.Y(n_1755)
);

OAI22xp5_ASAP7_75t_SL g1756 ( 
.A1(n_1452),
.A2(n_1190),
.B1(n_1194),
.B2(n_1184),
.Y(n_1756)
);

HB1xp67_ASAP7_75t_L g1757 ( 
.A(n_1670),
.Y(n_1757)
);

AND2x2_ASAP7_75t_L g1758 ( 
.A(n_1523),
.B(n_1391),
.Y(n_1758)
);

INVx1_ASAP7_75t_L g1759 ( 
.A(n_1511),
.Y(n_1759)
);

OAI22xp33_ASAP7_75t_L g1760 ( 
.A1(n_1599),
.A2(n_1402),
.B1(n_1403),
.B2(n_1401),
.Y(n_1760)
);

OAI22xp33_ASAP7_75t_R g1761 ( 
.A1(n_1464),
.A2(n_597),
.B1(n_600),
.B2(n_599),
.Y(n_1761)
);

AOI22xp5_ASAP7_75t_L g1762 ( 
.A1(n_1520),
.A2(n_1404),
.B1(n_1405),
.B2(n_1403),
.Y(n_1762)
);

AOI22xp5_ASAP7_75t_L g1763 ( 
.A1(n_1534),
.A2(n_1405),
.B1(n_1406),
.B2(n_1404),
.Y(n_1763)
);

AO22x2_ASAP7_75t_L g1764 ( 
.A1(n_1690),
.A2(n_600),
.B1(n_619),
.B2(n_602),
.Y(n_1764)
);

INVx8_ASAP7_75t_L g1765 ( 
.A(n_1546),
.Y(n_1765)
);

OAI22xp33_ASAP7_75t_L g1766 ( 
.A1(n_1599),
.A2(n_1408),
.B1(n_1410),
.B2(n_1406),
.Y(n_1766)
);

AOI22xp5_ASAP7_75t_L g1767 ( 
.A1(n_1566),
.A2(n_1410),
.B1(n_1415),
.B2(n_1408),
.Y(n_1767)
);

INVx1_ASAP7_75t_L g1768 ( 
.A(n_1511),
.Y(n_1768)
);

AOI22xp5_ASAP7_75t_L g1769 ( 
.A1(n_1566),
.A2(n_1416),
.B1(n_1427),
.B2(n_1415),
.Y(n_1769)
);

OAI22xp33_ASAP7_75t_L g1770 ( 
.A1(n_1661),
.A2(n_1427),
.B1(n_1416),
.B2(n_1023),
.Y(n_1770)
);

OAI22xp5_ASAP7_75t_SL g1771 ( 
.A1(n_1603),
.A2(n_1200),
.B1(n_1337),
.B2(n_1331),
.Y(n_1771)
);

BUFx6f_ASAP7_75t_SL g1772 ( 
.A(n_1698),
.Y(n_1772)
);

OA22x2_ASAP7_75t_L g1773 ( 
.A1(n_1616),
.A2(n_1034),
.B1(n_1040),
.B2(n_1017),
.Y(n_1773)
);

BUFx10_ASAP7_75t_L g1774 ( 
.A(n_1505),
.Y(n_1774)
);

AO22x2_ASAP7_75t_L g1775 ( 
.A1(n_1690),
.A2(n_602),
.B1(n_622),
.B2(n_619),
.Y(n_1775)
);

AOI22xp5_ASAP7_75t_L g1776 ( 
.A1(n_1566),
.A2(n_1040),
.B1(n_1043),
.B2(n_1034),
.Y(n_1776)
);

XNOR2xp5_ASAP7_75t_L g1777 ( 
.A(n_1461),
.B(n_1148),
.Y(n_1777)
);

AOI22xp5_ASAP7_75t_L g1778 ( 
.A1(n_1566),
.A2(n_1046),
.B1(n_1048),
.B2(n_1043),
.Y(n_1778)
);

OAI22xp33_ASAP7_75t_L g1779 ( 
.A1(n_1661),
.A2(n_1053),
.B1(n_1062),
.B2(n_1052),
.Y(n_1779)
);

INVx2_ASAP7_75t_L g1780 ( 
.A(n_1455),
.Y(n_1780)
);

AND2x4_ASAP7_75t_L g1781 ( 
.A(n_1611),
.B(n_1072),
.Y(n_1781)
);

OAI22xp33_ASAP7_75t_L g1782 ( 
.A1(n_1661),
.A2(n_1062),
.B1(n_1063),
.B2(n_1053),
.Y(n_1782)
);

AO22x2_ASAP7_75t_L g1783 ( 
.A1(n_1691),
.A2(n_623),
.B1(n_627),
.B2(n_622),
.Y(n_1783)
);

INVx1_ASAP7_75t_L g1784 ( 
.A(n_1511),
.Y(n_1784)
);

INVx1_ASAP7_75t_L g1785 ( 
.A(n_1511),
.Y(n_1785)
);

INVx1_ASAP7_75t_L g1786 ( 
.A(n_1514),
.Y(n_1786)
);

OAI22xp33_ASAP7_75t_SL g1787 ( 
.A1(n_1564),
.A2(n_1064),
.B1(n_1066),
.B2(n_1063),
.Y(n_1787)
);

AO22x2_ASAP7_75t_L g1788 ( 
.A1(n_1691),
.A2(n_627),
.B1(n_631),
.B2(n_623),
.Y(n_1788)
);

NAND2xp5_ASAP7_75t_L g1789 ( 
.A(n_1469),
.B(n_1064),
.Y(n_1789)
);

OR2x2_ASAP7_75t_L g1790 ( 
.A(n_1654),
.B(n_1066),
.Y(n_1790)
);

INVx2_ASAP7_75t_L g1791 ( 
.A(n_1456),
.Y(n_1791)
);

INVx8_ASAP7_75t_L g1792 ( 
.A(n_1546),
.Y(n_1792)
);

OR2x6_ASAP7_75t_L g1793 ( 
.A(n_1544),
.B(n_1022),
.Y(n_1793)
);

OAI22xp33_ASAP7_75t_SL g1794 ( 
.A1(n_1472),
.A2(n_1073),
.B1(n_1077),
.B2(n_1071),
.Y(n_1794)
);

AND2x2_ASAP7_75t_L g1795 ( 
.A(n_1722),
.B(n_1071),
.Y(n_1795)
);

BUFx10_ASAP7_75t_L g1796 ( 
.A(n_1682),
.Y(n_1796)
);

OAI22xp33_ASAP7_75t_L g1797 ( 
.A1(n_1661),
.A2(n_1077),
.B1(n_1085),
.B2(n_1073),
.Y(n_1797)
);

INVx1_ASAP7_75t_L g1798 ( 
.A(n_1514),
.Y(n_1798)
);

AND2x4_ASAP7_75t_L g1799 ( 
.A(n_1611),
.B(n_1074),
.Y(n_1799)
);

AOI22xp5_ASAP7_75t_L g1800 ( 
.A1(n_1566),
.A2(n_1089),
.B1(n_1094),
.B2(n_1085),
.Y(n_1800)
);

OAI22xp33_ASAP7_75t_R g1801 ( 
.A1(n_1454),
.A2(n_666),
.B1(n_667),
.B2(n_631),
.Y(n_1801)
);

INVx2_ASAP7_75t_L g1802 ( 
.A(n_1456),
.Y(n_1802)
);

AOI22xp5_ASAP7_75t_L g1803 ( 
.A1(n_1684),
.A2(n_1096),
.B1(n_1102),
.B2(n_1095),
.Y(n_1803)
);

NOR2xp33_ASAP7_75t_L g1804 ( 
.A(n_1661),
.B(n_1096),
.Y(n_1804)
);

AOI22xp5_ASAP7_75t_L g1805 ( 
.A1(n_1684),
.A2(n_1104),
.B1(n_1106),
.B2(n_1102),
.Y(n_1805)
);

AOI22xp5_ASAP7_75t_SL g1806 ( 
.A1(n_1587),
.A2(n_1345),
.B1(n_1363),
.B2(n_1341),
.Y(n_1806)
);

INVx2_ASAP7_75t_L g1807 ( 
.A(n_1456),
.Y(n_1807)
);

INVx1_ASAP7_75t_L g1808 ( 
.A(n_1514),
.Y(n_1808)
);

AOI22xp5_ASAP7_75t_L g1809 ( 
.A1(n_1684),
.A2(n_1106),
.B1(n_1109),
.B2(n_1104),
.Y(n_1809)
);

INVx2_ASAP7_75t_L g1810 ( 
.A(n_1439),
.Y(n_1810)
);

AOI22xp5_ASAP7_75t_L g1811 ( 
.A1(n_1684),
.A2(n_1694),
.B1(n_1707),
.B2(n_1668),
.Y(n_1811)
);

INVx2_ASAP7_75t_L g1812 ( 
.A(n_1439),
.Y(n_1812)
);

OAI22xp33_ASAP7_75t_L g1813 ( 
.A1(n_1668),
.A2(n_1674),
.B1(n_1713),
.B2(n_1673),
.Y(n_1813)
);

AOI22x1_ASAP7_75t_SL g1814 ( 
.A1(n_1714),
.A2(n_1268),
.B1(n_1156),
.B2(n_1159),
.Y(n_1814)
);

BUFx10_ASAP7_75t_L g1815 ( 
.A(n_1682),
.Y(n_1815)
);

INVx1_ASAP7_75t_L g1816 ( 
.A(n_1514),
.Y(n_1816)
);

AOI22xp5_ASAP7_75t_L g1817 ( 
.A1(n_1684),
.A2(n_1114),
.B1(n_1117),
.B2(n_1110),
.Y(n_1817)
);

AOI22xp5_ASAP7_75t_L g1818 ( 
.A1(n_1684),
.A2(n_1125),
.B1(n_1127),
.B2(n_1117),
.Y(n_1818)
);

INVx2_ASAP7_75t_L g1819 ( 
.A(n_1441),
.Y(n_1819)
);

AND2x2_ASAP7_75t_L g1820 ( 
.A(n_1722),
.B(n_1125),
.Y(n_1820)
);

OAI22xp33_ASAP7_75t_SL g1821 ( 
.A1(n_1472),
.A2(n_1129),
.B1(n_1134),
.B2(n_1127),
.Y(n_1821)
);

OAI22xp33_ASAP7_75t_L g1822 ( 
.A1(n_1668),
.A2(n_1134),
.B1(n_1129),
.B2(n_610),
.Y(n_1822)
);

INVx2_ASAP7_75t_L g1823 ( 
.A(n_1441),
.Y(n_1823)
);

INVx1_ASAP7_75t_L g1824 ( 
.A(n_1575),
.Y(n_1824)
);

AND2x2_ASAP7_75t_L g1825 ( 
.A(n_1652),
.B(n_1155),
.Y(n_1825)
);

BUFx6f_ASAP7_75t_L g1826 ( 
.A(n_1630),
.Y(n_1826)
);

INVx2_ASAP7_75t_L g1827 ( 
.A(n_1442),
.Y(n_1827)
);

OAI22xp5_ASAP7_75t_SL g1828 ( 
.A1(n_1603),
.A2(n_1367),
.B1(n_1376),
.B2(n_1365),
.Y(n_1828)
);

AOI22xp5_ASAP7_75t_L g1829 ( 
.A1(n_1684),
.A2(n_1436),
.B1(n_1382),
.B2(n_1384),
.Y(n_1829)
);

OR2x2_ASAP7_75t_L g1830 ( 
.A(n_1654),
.B(n_1155),
.Y(n_1830)
);

OAI22xp33_ASAP7_75t_SL g1831 ( 
.A1(n_1655),
.A2(n_667),
.B1(n_670),
.B2(n_666),
.Y(n_1831)
);

AND2x2_ASAP7_75t_L g1832 ( 
.A(n_1652),
.B(n_1156),
.Y(n_1832)
);

OAI22xp5_ASAP7_75t_SL g1833 ( 
.A1(n_1545),
.A2(n_1394),
.B1(n_1396),
.B2(n_1381),
.Y(n_1833)
);

OAI22xp33_ASAP7_75t_SL g1834 ( 
.A1(n_1655),
.A2(n_672),
.B1(n_675),
.B2(n_670),
.Y(n_1834)
);

AND2x2_ASAP7_75t_L g1835 ( 
.A(n_1670),
.B(n_1159),
.Y(n_1835)
);

INVx1_ASAP7_75t_L g1836 ( 
.A(n_1575),
.Y(n_1836)
);

INVx3_ASAP7_75t_L g1837 ( 
.A(n_1626),
.Y(n_1837)
);

AND2x2_ASAP7_75t_L g1838 ( 
.A(n_1670),
.B(n_1160),
.Y(n_1838)
);

AND2x2_ASAP7_75t_L g1839 ( 
.A(n_1670),
.B(n_1160),
.Y(n_1839)
);

OAI22xp33_ASAP7_75t_L g1840 ( 
.A1(n_1673),
.A2(n_1713),
.B1(n_1674),
.B2(n_1459),
.Y(n_1840)
);

AOI22xp5_ASAP7_75t_L g1841 ( 
.A1(n_1694),
.A2(n_1414),
.B1(n_1434),
.B2(n_1399),
.Y(n_1841)
);

INVx2_ASAP7_75t_L g1842 ( 
.A(n_1442),
.Y(n_1842)
);

AO22x2_ASAP7_75t_L g1843 ( 
.A1(n_1692),
.A2(n_675),
.B1(n_676),
.B2(n_672),
.Y(n_1843)
);

INVx2_ASAP7_75t_L g1844 ( 
.A(n_1443),
.Y(n_1844)
);

INVx2_ASAP7_75t_L g1845 ( 
.A(n_1443),
.Y(n_1845)
);

OAI22xp33_ASAP7_75t_SL g1846 ( 
.A1(n_1657),
.A2(n_678),
.B1(n_702),
.B2(n_676),
.Y(n_1846)
);

OAI22xp33_ASAP7_75t_L g1847 ( 
.A1(n_1673),
.A2(n_610),
.B1(n_615),
.B2(n_555),
.Y(n_1847)
);

OR2x6_ASAP7_75t_L g1848 ( 
.A(n_1558),
.B(n_1032),
.Y(n_1848)
);

BUFx6f_ASAP7_75t_SL g1849 ( 
.A(n_1698),
.Y(n_1849)
);

OAI22xp33_ASAP7_75t_SL g1850 ( 
.A1(n_1657),
.A2(n_702),
.B1(n_703),
.B2(n_678),
.Y(n_1850)
);

OAI22xp33_ASAP7_75t_SL g1851 ( 
.A1(n_1658),
.A2(n_717),
.B1(n_719),
.B2(n_703),
.Y(n_1851)
);

OAI22xp5_ASAP7_75t_L g1852 ( 
.A1(n_1646),
.A2(n_732),
.B1(n_734),
.B2(n_724),
.Y(n_1852)
);

INVx2_ASAP7_75t_L g1853 ( 
.A(n_1448),
.Y(n_1853)
);

INVx2_ASAP7_75t_L g1854 ( 
.A(n_1448),
.Y(n_1854)
);

AOI22xp5_ASAP7_75t_L g1855 ( 
.A1(n_1694),
.A2(n_1435),
.B1(n_1210),
.B2(n_1170),
.Y(n_1855)
);

AOI22xp5_ASAP7_75t_L g1856 ( 
.A1(n_1694),
.A2(n_1210),
.B1(n_1264),
.B2(n_1269),
.Y(n_1856)
);

INVx3_ASAP7_75t_L g1857 ( 
.A(n_1626),
.Y(n_1857)
);

AOI22xp5_ASAP7_75t_L g1858 ( 
.A1(n_1694),
.A2(n_1281),
.B1(n_1283),
.B2(n_1270),
.Y(n_1858)
);

INVx2_ASAP7_75t_SL g1859 ( 
.A(n_1662),
.Y(n_1859)
);

OAI22xp33_ASAP7_75t_L g1860 ( 
.A1(n_1674),
.A2(n_615),
.B1(n_699),
.B2(n_555),
.Y(n_1860)
);

INVx1_ASAP7_75t_SL g1861 ( 
.A(n_1585),
.Y(n_1861)
);

INVx1_ASAP7_75t_L g1862 ( 
.A(n_1575),
.Y(n_1862)
);

AO22x2_ASAP7_75t_L g1863 ( 
.A1(n_1692),
.A2(n_717),
.B1(n_731),
.B2(n_719),
.Y(n_1863)
);

OR2x2_ASAP7_75t_L g1864 ( 
.A(n_1605),
.B(n_1161),
.Y(n_1864)
);

AOI22xp5_ASAP7_75t_L g1865 ( 
.A1(n_1694),
.A2(n_730),
.B1(n_699),
.B2(n_735),
.Y(n_1865)
);

OAI22xp33_ASAP7_75t_L g1866 ( 
.A1(n_1674),
.A2(n_730),
.B1(n_699),
.B2(n_731),
.Y(n_1866)
);

AND2x2_ASAP7_75t_L g1867 ( 
.A(n_1678),
.B(n_1161),
.Y(n_1867)
);

AND2x2_ASAP7_75t_L g1868 ( 
.A(n_1678),
.B(n_1167),
.Y(n_1868)
);

AOI22xp5_ASAP7_75t_L g1869 ( 
.A1(n_1694),
.A2(n_730),
.B1(n_739),
.B2(n_737),
.Y(n_1869)
);

OAI22xp33_ASAP7_75t_L g1870 ( 
.A1(n_1713),
.A2(n_736),
.B1(n_738),
.B2(n_733),
.Y(n_1870)
);

NAND2xp5_ASAP7_75t_L g1871 ( 
.A(n_1646),
.B(n_834),
.Y(n_1871)
);

OAI22xp33_ASAP7_75t_R g1872 ( 
.A1(n_1633),
.A2(n_736),
.B1(n_738),
.B2(n_733),
.Y(n_1872)
);

BUFx10_ASAP7_75t_L g1873 ( 
.A(n_1682),
.Y(n_1873)
);

INVx2_ASAP7_75t_L g1874 ( 
.A(n_1463),
.Y(n_1874)
);

OAI22xp33_ASAP7_75t_SL g1875 ( 
.A1(n_1658),
.A2(n_744),
.B1(n_748),
.B2(n_746),
.Y(n_1875)
);

AOI22xp5_ASAP7_75t_L g1876 ( 
.A1(n_1707),
.A2(n_1286),
.B1(n_1168),
.B2(n_1178),
.Y(n_1876)
);

INVx2_ASAP7_75t_L g1877 ( 
.A(n_1468),
.Y(n_1877)
);

OAI22xp33_ASAP7_75t_SL g1878 ( 
.A1(n_1471),
.A2(n_1616),
.B1(n_1555),
.B2(n_1532),
.Y(n_1878)
);

AND2x2_ASAP7_75t_L g1879 ( 
.A(n_1678),
.B(n_1168),
.Y(n_1879)
);

AND2x2_ASAP7_75t_L g1880 ( 
.A(n_1662),
.B(n_1174),
.Y(n_1880)
);

INVx2_ASAP7_75t_L g1881 ( 
.A(n_1468),
.Y(n_1881)
);

OR2x6_ASAP7_75t_L g1882 ( 
.A(n_1585),
.B(n_1660),
.Y(n_1882)
);

INVx1_ASAP7_75t_SL g1883 ( 
.A(n_1701),
.Y(n_1883)
);

OAI22xp33_ASAP7_75t_L g1884 ( 
.A1(n_1713),
.A2(n_744),
.B1(n_748),
.B2(n_746),
.Y(n_1884)
);

AND2x2_ASAP7_75t_L g1885 ( 
.A(n_1649),
.B(n_1174),
.Y(n_1885)
);

NAND3x1_ASAP7_75t_L g1886 ( 
.A(n_1708),
.B(n_763),
.C(n_1075),
.Y(n_1886)
);

INVx2_ASAP7_75t_L g1887 ( 
.A(n_1473),
.Y(n_1887)
);

INVx1_ASAP7_75t_L g1888 ( 
.A(n_1575),
.Y(n_1888)
);

OAI22xp5_ASAP7_75t_SL g1889 ( 
.A1(n_1545),
.A2(n_1179),
.B1(n_1183),
.B2(n_1178),
.Y(n_1889)
);

AND2x2_ASAP7_75t_L g1890 ( 
.A(n_1649),
.B(n_1179),
.Y(n_1890)
);

OAI22xp33_ASAP7_75t_L g1891 ( 
.A1(n_1457),
.A2(n_763),
.B1(n_747),
.B2(n_749),
.Y(n_1891)
);

AOI22xp5_ASAP7_75t_L g1892 ( 
.A1(n_1707),
.A2(n_1183),
.B1(n_1193),
.B2(n_1185),
.Y(n_1892)
);

NAND3x1_ASAP7_75t_L g1893 ( 
.A(n_1660),
.B(n_1081),
.C(n_1080),
.Y(n_1893)
);

AO22x2_ASAP7_75t_L g1894 ( 
.A1(n_1693),
.A2(n_1061),
.B1(n_1083),
.B2(n_1082),
.Y(n_1894)
);

AND2x2_ASAP7_75t_L g1895 ( 
.A(n_1576),
.B(n_1185),
.Y(n_1895)
);

INVx1_ASAP7_75t_L g1896 ( 
.A(n_1583),
.Y(n_1896)
);

OAI22xp33_ASAP7_75t_L g1897 ( 
.A1(n_1457),
.A2(n_750),
.B1(n_751),
.B2(n_743),
.Y(n_1897)
);

AOI22xp5_ASAP7_75t_L g1898 ( 
.A1(n_1707),
.A2(n_1196),
.B1(n_1198),
.B2(n_1193),
.Y(n_1898)
);

AND2x2_ASAP7_75t_L g1899 ( 
.A(n_1577),
.B(n_1196),
.Y(n_1899)
);

OAI22xp33_ASAP7_75t_L g1900 ( 
.A1(n_1457),
.A2(n_754),
.B1(n_765),
.B2(n_753),
.Y(n_1900)
);

INVx2_ASAP7_75t_L g1901 ( 
.A(n_1479),
.Y(n_1901)
);

INVx1_ASAP7_75t_L g1902 ( 
.A(n_1583),
.Y(n_1902)
);

INVx2_ASAP7_75t_L g1903 ( 
.A(n_1583),
.Y(n_1903)
);

AND2x2_ASAP7_75t_L g1904 ( 
.A(n_1656),
.B(n_1198),
.Y(n_1904)
);

BUFx6f_ASAP7_75t_L g1905 ( 
.A(n_1630),
.Y(n_1905)
);

INVx1_ASAP7_75t_L g1906 ( 
.A(n_1583),
.Y(n_1906)
);

AND2x2_ASAP7_75t_L g1907 ( 
.A(n_1656),
.B(n_1206),
.Y(n_1907)
);

OAI22xp5_ASAP7_75t_L g1908 ( 
.A1(n_1646),
.A2(n_767),
.B1(n_768),
.B2(n_766),
.Y(n_1908)
);

OA22x2_ASAP7_75t_L g1909 ( 
.A1(n_1663),
.A2(n_1682),
.B1(n_1721),
.B2(n_1706),
.Y(n_1909)
);

AO22x2_ASAP7_75t_L g1910 ( 
.A1(n_1693),
.A2(n_1091),
.B1(n_1092),
.B2(n_1084),
.Y(n_1910)
);

OAI22xp33_ASAP7_75t_SL g1911 ( 
.A1(n_1532),
.A2(n_1206),
.B1(n_1211),
.B2(n_1209),
.Y(n_1911)
);

AND2x2_ASAP7_75t_L g1912 ( 
.A(n_1706),
.B(n_1209),
.Y(n_1912)
);

OAI22xp33_ASAP7_75t_SL g1913 ( 
.A1(n_1533),
.A2(n_1211),
.B1(n_770),
.B2(n_1100),
.Y(n_1913)
);

NAND2xp5_ASAP7_75t_L g1914 ( 
.A(n_1646),
.B(n_834),
.Y(n_1914)
);

AO22x2_ASAP7_75t_L g1915 ( 
.A1(n_1700),
.A2(n_1101),
.B1(n_1103),
.B2(n_1099),
.Y(n_1915)
);

AOI22xp5_ASAP7_75t_L g1916 ( 
.A1(n_1707),
.A2(n_1108),
.B1(n_1118),
.B2(n_1115),
.Y(n_1916)
);

AO22x2_ASAP7_75t_L g1917 ( 
.A1(n_1700),
.A2(n_1121),
.B1(n_1124),
.B2(n_1119),
.Y(n_1917)
);

OAI22xp33_ASAP7_75t_L g1918 ( 
.A1(n_1459),
.A2(n_1130),
.B1(n_1131),
.B2(n_1128),
.Y(n_1918)
);

INVx2_ASAP7_75t_L g1919 ( 
.A(n_1536),
.Y(n_1919)
);

AOI22xp5_ASAP7_75t_L g1920 ( 
.A1(n_1707),
.A2(n_1132),
.B1(n_860),
.B2(n_975),
.Y(n_1920)
);

AND2x2_ASAP7_75t_L g1921 ( 
.A(n_1706),
.B(n_1126),
.Y(n_1921)
);

AND2x2_ASAP7_75t_L g1922 ( 
.A(n_1706),
.B(n_1126),
.Y(n_1922)
);

AND2x2_ASAP7_75t_L g1923 ( 
.A(n_1721),
.B(n_1126),
.Y(n_1923)
);

AOI22xp5_ASAP7_75t_L g1924 ( 
.A1(n_1707),
.A2(n_1621),
.B1(n_1721),
.B2(n_1571),
.Y(n_1924)
);

INVx2_ASAP7_75t_L g1925 ( 
.A(n_1536),
.Y(n_1925)
);

AND2x2_ASAP7_75t_L g1926 ( 
.A(n_1721),
.B(n_1126),
.Y(n_1926)
);

INVx1_ASAP7_75t_L g1927 ( 
.A(n_1536),
.Y(n_1927)
);

AOI22xp5_ASAP7_75t_L g1928 ( 
.A1(n_1621),
.A2(n_975),
.B1(n_984),
.B2(n_920),
.Y(n_1928)
);

AND2x2_ASAP7_75t_L g1929 ( 
.A(n_1624),
.B(n_920),
.Y(n_1929)
);

INVxp67_ASAP7_75t_SL g1930 ( 
.A(n_1465),
.Y(n_1930)
);

INVx1_ASAP7_75t_L g1931 ( 
.A(n_1568),
.Y(n_1931)
);

BUFx10_ASAP7_75t_L g1932 ( 
.A(n_1679),
.Y(n_1932)
);

BUFx3_ASAP7_75t_L g1933 ( 
.A(n_1470),
.Y(n_1933)
);

OAI22xp33_ASAP7_75t_SL g1934 ( 
.A1(n_1533),
.A2(n_6),
.B1(n_4),
.B2(n_5),
.Y(n_1934)
);

AOI22xp5_ASAP7_75t_L g1935 ( 
.A1(n_1621),
.A2(n_975),
.B1(n_984),
.B2(n_920),
.Y(n_1935)
);

NAND2xp5_ASAP7_75t_L g1936 ( 
.A(n_1646),
.B(n_920),
.Y(n_1936)
);

OAI22xp33_ASAP7_75t_L g1937 ( 
.A1(n_1648),
.A2(n_975),
.B1(n_984),
.B2(n_920),
.Y(n_1937)
);

AND2x2_ASAP7_75t_SL g1938 ( 
.A(n_1680),
.B(n_984),
.Y(n_1938)
);

OAI22xp33_ASAP7_75t_SL g1939 ( 
.A1(n_1537),
.A2(n_10),
.B1(n_6),
.B2(n_8),
.Y(n_1939)
);

NAND3x1_ASAP7_75t_L g1940 ( 
.A(n_1660),
.B(n_1689),
.C(n_1669),
.Y(n_1940)
);

INVx1_ASAP7_75t_L g1941 ( 
.A(n_1568),
.Y(n_1941)
);

INVx1_ASAP7_75t_L g1942 ( 
.A(n_1568),
.Y(n_1942)
);

OAI22xp33_ASAP7_75t_L g1943 ( 
.A1(n_1648),
.A2(n_1030),
.B1(n_1067),
.B2(n_993),
.Y(n_1943)
);

OAI22xp5_ASAP7_75t_SL g1944 ( 
.A1(n_1663),
.A2(n_11),
.B1(n_8),
.B2(n_10),
.Y(n_1944)
);

AOI22xp5_ASAP7_75t_L g1945 ( 
.A1(n_1621),
.A2(n_1030),
.B1(n_1067),
.B2(n_993),
.Y(n_1945)
);

INVx2_ASAP7_75t_L g1946 ( 
.A(n_1529),
.Y(n_1946)
);

INVx2_ASAP7_75t_L g1947 ( 
.A(n_1529),
.Y(n_1947)
);

OR2x6_ASAP7_75t_L g1948 ( 
.A(n_1660),
.B(n_993),
.Y(n_1948)
);

INVx2_ASAP7_75t_L g1949 ( 
.A(n_1529),
.Y(n_1949)
);

OAI22xp33_ASAP7_75t_L g1950 ( 
.A1(n_1537),
.A2(n_1030),
.B1(n_1067),
.B2(n_993),
.Y(n_1950)
);

INVx2_ASAP7_75t_L g1951 ( 
.A(n_1529),
.Y(n_1951)
);

AOI22xp5_ASAP7_75t_L g1952 ( 
.A1(n_1571),
.A2(n_1067),
.B1(n_1098),
.B2(n_1030),
.Y(n_1952)
);

AO22x2_ASAP7_75t_L g1953 ( 
.A1(n_1718),
.A2(n_14),
.B1(n_11),
.B2(n_12),
.Y(n_1953)
);

AOI22xp5_ASAP7_75t_L g1954 ( 
.A1(n_1540),
.A2(n_1112),
.B1(n_1098),
.B2(n_296),
.Y(n_1954)
);

OAI22xp5_ASAP7_75t_SL g1955 ( 
.A1(n_1506),
.A2(n_16),
.B1(n_12),
.B2(n_15),
.Y(n_1955)
);

AO22x2_ASAP7_75t_L g1956 ( 
.A1(n_1718),
.A2(n_18),
.B1(n_15),
.B2(n_17),
.Y(n_1956)
);

AOI22xp5_ASAP7_75t_L g1957 ( 
.A1(n_1524),
.A2(n_1112),
.B1(n_1098),
.B2(n_297),
.Y(n_1957)
);

BUFx6f_ASAP7_75t_L g1958 ( 
.A(n_1630),
.Y(n_1958)
);

OR2x2_ASAP7_75t_L g1959 ( 
.A(n_1589),
.B(n_17),
.Y(n_1959)
);

AO22x2_ASAP7_75t_L g1960 ( 
.A1(n_1672),
.A2(n_22),
.B1(n_19),
.B2(n_21),
.Y(n_1960)
);

INVx2_ASAP7_75t_L g1961 ( 
.A(n_1529),
.Y(n_1961)
);

AND2x2_ASAP7_75t_L g1962 ( 
.A(n_1624),
.B(n_1112),
.Y(n_1962)
);

OAI22xp33_ASAP7_75t_SL g1963 ( 
.A1(n_1538),
.A2(n_23),
.B1(n_21),
.B2(n_22),
.Y(n_1963)
);

INVx1_ASAP7_75t_L g1964 ( 
.A(n_1622),
.Y(n_1964)
);

HB1xp67_ASAP7_75t_L g1965 ( 
.A(n_1659),
.Y(n_1965)
);

AO22x2_ASAP7_75t_L g1966 ( 
.A1(n_1695),
.A2(n_25),
.B1(n_23),
.B2(n_24),
.Y(n_1966)
);

AO22x2_ASAP7_75t_L g1967 ( 
.A1(n_1695),
.A2(n_26),
.B1(n_24),
.B2(n_25),
.Y(n_1967)
);

AOI22xp5_ASAP7_75t_L g1968 ( 
.A1(n_1524),
.A2(n_1112),
.B1(n_1098),
.B2(n_29),
.Y(n_1968)
);

AO22x2_ASAP7_75t_L g1969 ( 
.A1(n_1695),
.A2(n_29),
.B1(n_27),
.B2(n_28),
.Y(n_1969)
);

AOI22xp5_ASAP7_75t_L g1970 ( 
.A1(n_1626),
.A2(n_1112),
.B1(n_1098),
.B2(n_32),
.Y(n_1970)
);

AOI22xp5_ASAP7_75t_L g1971 ( 
.A1(n_1527),
.A2(n_299),
.B1(n_302),
.B2(n_293),
.Y(n_1971)
);

AND2x2_ASAP7_75t_L g1972 ( 
.A(n_1643),
.B(n_30),
.Y(n_1972)
);

AND2x2_ASAP7_75t_L g1973 ( 
.A(n_1643),
.B(n_30),
.Y(n_1973)
);

INVx1_ASAP7_75t_L g1974 ( 
.A(n_1622),
.Y(n_1974)
);

OR2x2_ASAP7_75t_L g1975 ( 
.A(n_1659),
.B(n_31),
.Y(n_1975)
);

OAI22xp5_ASAP7_75t_SL g1976 ( 
.A1(n_1572),
.A2(n_36),
.B1(n_31),
.B2(n_34),
.Y(n_1976)
);

AOI22xp5_ASAP7_75t_L g1977 ( 
.A1(n_1527),
.A2(n_307),
.B1(n_312),
.B2(n_306),
.Y(n_1977)
);

AOI22xp5_ASAP7_75t_L g1978 ( 
.A1(n_1527),
.A2(n_314),
.B1(n_315),
.B2(n_313),
.Y(n_1978)
);

OAI22xp5_ASAP7_75t_L g1979 ( 
.A1(n_1509),
.A2(n_317),
.B1(n_318),
.B2(n_316),
.Y(n_1979)
);

AOI22xp5_ASAP7_75t_L g1980 ( 
.A1(n_1527),
.A2(n_321),
.B1(n_322),
.B2(n_319),
.Y(n_1980)
);

NOR2x1p5_ASAP7_75t_L g1981 ( 
.A(n_1679),
.B(n_34),
.Y(n_1981)
);

INVx2_ASAP7_75t_L g1982 ( 
.A(n_1535),
.Y(n_1982)
);

OAI22xp5_ASAP7_75t_SL g1983 ( 
.A1(n_1591),
.A2(n_42),
.B1(n_39),
.B2(n_41),
.Y(n_1983)
);

INVx2_ASAP7_75t_L g1984 ( 
.A(n_1535),
.Y(n_1984)
);

OAI22xp33_ASAP7_75t_SL g1985 ( 
.A1(n_1538),
.A2(n_45),
.B1(n_39),
.B2(n_43),
.Y(n_1985)
);

AND2x2_ASAP7_75t_L g1986 ( 
.A(n_1696),
.B(n_45),
.Y(n_1986)
);

INVx1_ASAP7_75t_SL g1987 ( 
.A(n_1701),
.Y(n_1987)
);

AO22x2_ASAP7_75t_L g1988 ( 
.A1(n_1696),
.A2(n_50),
.B1(n_48),
.B2(n_49),
.Y(n_1988)
);

NOR2xp33_ASAP7_75t_L g1989 ( 
.A(n_1636),
.B(n_48),
.Y(n_1989)
);

AOI22xp5_ASAP7_75t_L g1990 ( 
.A1(n_1586),
.A2(n_329),
.B1(n_330),
.B2(n_326),
.Y(n_1990)
);

OAI22xp5_ASAP7_75t_L g1991 ( 
.A1(n_1647),
.A2(n_332),
.B1(n_334),
.B2(n_331),
.Y(n_1991)
);

OAI22xp33_ASAP7_75t_L g1992 ( 
.A1(n_1539),
.A2(n_53),
.B1(n_49),
.B2(n_52),
.Y(n_1992)
);

INVx2_ASAP7_75t_L g1993 ( 
.A(n_1535),
.Y(n_1993)
);

OAI22xp33_ASAP7_75t_L g1994 ( 
.A1(n_1539),
.A2(n_56),
.B1(n_53),
.B2(n_55),
.Y(n_1994)
);

INVx1_ASAP7_75t_L g1995 ( 
.A(n_1481),
.Y(n_1995)
);

OAI22xp5_ASAP7_75t_L g1996 ( 
.A1(n_1647),
.A2(n_337),
.B1(n_341),
.B2(n_335),
.Y(n_1996)
);

AO22x2_ASAP7_75t_L g1997 ( 
.A1(n_1696),
.A2(n_59),
.B1(n_55),
.B2(n_57),
.Y(n_1997)
);

AND2x2_ASAP7_75t_L g1998 ( 
.A(n_1699),
.B(n_59),
.Y(n_1998)
);

OAI22xp33_ASAP7_75t_L g1999 ( 
.A1(n_1542),
.A2(n_62),
.B1(n_60),
.B2(n_61),
.Y(n_1999)
);

AOI22xp5_ASAP7_75t_L g2000 ( 
.A1(n_1586),
.A2(n_346),
.B1(n_359),
.B2(n_344),
.Y(n_2000)
);

OAI22xp33_ASAP7_75t_L g2001 ( 
.A1(n_1542),
.A2(n_66),
.B1(n_63),
.B2(n_64),
.Y(n_2001)
);

NOR2xp33_ASAP7_75t_L g2002 ( 
.A(n_1729),
.B(n_1677),
.Y(n_2002)
);

NAND2xp5_ASAP7_75t_L g2003 ( 
.A(n_1804),
.B(n_1618),
.Y(n_2003)
);

INVx1_ASAP7_75t_L g2004 ( 
.A(n_1727),
.Y(n_2004)
);

AND2x2_ASAP7_75t_L g2005 ( 
.A(n_1724),
.B(n_1677),
.Y(n_2005)
);

AND2x2_ASAP7_75t_SL g2006 ( 
.A(n_1865),
.B(n_1680),
.Y(n_2006)
);

BUFx6f_ASAP7_75t_L g2007 ( 
.A(n_1732),
.Y(n_2007)
);

NOR2xp33_ASAP7_75t_L g2008 ( 
.A(n_1734),
.B(n_1677),
.Y(n_2008)
);

NOR2xp33_ASAP7_75t_L g2009 ( 
.A(n_1748),
.B(n_1677),
.Y(n_2009)
);

BUFx3_ASAP7_75t_L g2010 ( 
.A(n_1933),
.Y(n_2010)
);

INVx4_ASAP7_75t_L g2011 ( 
.A(n_1732),
.Y(n_2011)
);

AOI22xp33_ASAP7_75t_L g2012 ( 
.A1(n_1989),
.A2(n_1909),
.B1(n_1865),
.B2(n_1813),
.Y(n_2012)
);

INVx1_ASAP7_75t_SL g2013 ( 
.A(n_1861),
.Y(n_2013)
);

INVx1_ASAP7_75t_L g2014 ( 
.A(n_1927),
.Y(n_2014)
);

INVx1_ASAP7_75t_L g2015 ( 
.A(n_1931),
.Y(n_2015)
);

INVx2_ASAP7_75t_L g2016 ( 
.A(n_1931),
.Y(n_2016)
);

INVx1_ASAP7_75t_L g2017 ( 
.A(n_1941),
.Y(n_2017)
);

BUFx10_ASAP7_75t_L g2018 ( 
.A(n_1772),
.Y(n_2018)
);

INVx2_ASAP7_75t_L g2019 ( 
.A(n_1941),
.Y(n_2019)
);

NAND2xp5_ASAP7_75t_SL g2020 ( 
.A(n_1789),
.B(n_1723),
.Y(n_2020)
);

INVx4_ASAP7_75t_L g2021 ( 
.A(n_1826),
.Y(n_2021)
);

AND3x1_ASAP7_75t_L g2022 ( 
.A(n_1749),
.B(n_1711),
.C(n_1608),
.Y(n_2022)
);

INVx1_ASAP7_75t_L g2023 ( 
.A(n_1727),
.Y(n_2023)
);

INVx2_ASAP7_75t_L g2024 ( 
.A(n_1942),
.Y(n_2024)
);

BUFx3_ASAP7_75t_L g2025 ( 
.A(n_1826),
.Y(n_2025)
);

INVx1_ASAP7_75t_L g2026 ( 
.A(n_1942),
.Y(n_2026)
);

NOR2xp33_ASAP7_75t_L g2027 ( 
.A(n_1779),
.B(n_1688),
.Y(n_2027)
);

INVx3_ASAP7_75t_L g2028 ( 
.A(n_1903),
.Y(n_2028)
);

INVx2_ASAP7_75t_L g2029 ( 
.A(n_1995),
.Y(n_2029)
);

INVx3_ASAP7_75t_L g2030 ( 
.A(n_1837),
.Y(n_2030)
);

NAND2xp5_ASAP7_75t_SL g2031 ( 
.A(n_1751),
.B(n_1723),
.Y(n_2031)
);

INVx4_ASAP7_75t_L g2032 ( 
.A(n_1826),
.Y(n_2032)
);

INVx1_ASAP7_75t_L g2033 ( 
.A(n_1995),
.Y(n_2033)
);

BUFx10_ASAP7_75t_L g2034 ( 
.A(n_1772),
.Y(n_2034)
);

BUFx4f_ASAP7_75t_L g2035 ( 
.A(n_1905),
.Y(n_2035)
);

INVx2_ASAP7_75t_L g2036 ( 
.A(n_1728),
.Y(n_2036)
);

NOR2xp33_ASAP7_75t_L g2037 ( 
.A(n_1782),
.B(n_1688),
.Y(n_2037)
);

BUFx3_ASAP7_75t_L g2038 ( 
.A(n_1905),
.Y(n_2038)
);

INVx2_ASAP7_75t_L g2039 ( 
.A(n_1728),
.Y(n_2039)
);

INVxp67_ASAP7_75t_SL g2040 ( 
.A(n_1905),
.Y(n_2040)
);

NOR2xp33_ASAP7_75t_L g2041 ( 
.A(n_1797),
.B(n_1688),
.Y(n_2041)
);

INVx1_ASAP7_75t_L g2042 ( 
.A(n_1744),
.Y(n_2042)
);

AND2x2_ASAP7_75t_L g2043 ( 
.A(n_1757),
.B(n_1688),
.Y(n_2043)
);

INVx1_ASAP7_75t_L g2044 ( 
.A(n_1744),
.Y(n_2044)
);

NAND2xp5_ASAP7_75t_SL g2045 ( 
.A(n_1751),
.B(n_1723),
.Y(n_2045)
);

AND2x2_ASAP7_75t_L g2046 ( 
.A(n_1795),
.B(n_1697),
.Y(n_2046)
);

OR2x2_ASAP7_75t_L g2047 ( 
.A(n_1736),
.B(n_1702),
.Y(n_2047)
);

AND2x2_ASAP7_75t_L g2048 ( 
.A(n_1820),
.B(n_1697),
.Y(n_2048)
);

NOR2xp33_ASAP7_75t_L g2049 ( 
.A(n_1774),
.B(n_1697),
.Y(n_2049)
);

INVx1_ASAP7_75t_L g2050 ( 
.A(n_1755),
.Y(n_2050)
);

NOR2xp33_ASAP7_75t_L g2051 ( 
.A(n_1774),
.B(n_1697),
.Y(n_2051)
);

NOR2xp33_ASAP7_75t_L g2052 ( 
.A(n_1770),
.B(n_1717),
.Y(n_2052)
);

INVx1_ASAP7_75t_L g2053 ( 
.A(n_1755),
.Y(n_2053)
);

INVx2_ASAP7_75t_L g2054 ( 
.A(n_1759),
.Y(n_2054)
);

NAND2xp5_ASAP7_75t_SL g2055 ( 
.A(n_1859),
.B(n_1723),
.Y(n_2055)
);

INVx1_ASAP7_75t_L g2056 ( 
.A(n_1759),
.Y(n_2056)
);

NAND2xp5_ASAP7_75t_SL g2057 ( 
.A(n_1747),
.B(n_1723),
.Y(n_2057)
);

INVx2_ASAP7_75t_L g2058 ( 
.A(n_1768),
.Y(n_2058)
);

INVx3_ASAP7_75t_L g2059 ( 
.A(n_1837),
.Y(n_2059)
);

OR2x6_ASAP7_75t_L g2060 ( 
.A(n_1765),
.B(n_1680),
.Y(n_2060)
);

NAND2xp5_ASAP7_75t_SL g2061 ( 
.A(n_1803),
.B(n_1723),
.Y(n_2061)
);

INVx1_ASAP7_75t_L g2062 ( 
.A(n_1768),
.Y(n_2062)
);

NOR2xp33_ASAP7_75t_L g2063 ( 
.A(n_1758),
.B(n_1717),
.Y(n_2063)
);

NAND2xp5_ASAP7_75t_SL g2064 ( 
.A(n_1803),
.B(n_1680),
.Y(n_2064)
);

INVx1_ASAP7_75t_SL g2065 ( 
.A(n_1885),
.Y(n_2065)
);

INVx1_ASAP7_75t_L g2066 ( 
.A(n_1784),
.Y(n_2066)
);

INVx2_ASAP7_75t_L g2067 ( 
.A(n_1784),
.Y(n_2067)
);

AOI22xp33_ASAP7_75t_L g2068 ( 
.A1(n_1857),
.A2(n_1517),
.B1(n_1513),
.B2(n_1618),
.Y(n_2068)
);

AND2x2_ASAP7_75t_L g2069 ( 
.A(n_1929),
.B(n_1717),
.Y(n_2069)
);

INVx4_ASAP7_75t_L g2070 ( 
.A(n_1958),
.Y(n_2070)
);

OR2x6_ASAP7_75t_L g2071 ( 
.A(n_1765),
.B(n_1680),
.Y(n_2071)
);

OAI22xp33_ASAP7_75t_L g2072 ( 
.A1(n_1924),
.A2(n_1703),
.B1(n_1709),
.B2(n_1699),
.Y(n_2072)
);

INVx2_ASAP7_75t_L g2073 ( 
.A(n_1785),
.Y(n_2073)
);

AND2x2_ASAP7_75t_L g2074 ( 
.A(n_1962),
.B(n_1717),
.Y(n_2074)
);

NOR3xp33_ASAP7_75t_L g2075 ( 
.A(n_1750),
.B(n_1484),
.C(n_1687),
.Y(n_2075)
);

NAND2xp5_ASAP7_75t_SL g2076 ( 
.A(n_1796),
.B(n_1685),
.Y(n_2076)
);

OR2x6_ASAP7_75t_L g2077 ( 
.A(n_1792),
.B(n_1685),
.Y(n_2077)
);

INVx2_ASAP7_75t_L g2078 ( 
.A(n_1785),
.Y(n_2078)
);

INVx2_ASAP7_75t_L g2079 ( 
.A(n_1786),
.Y(n_2079)
);

AND2x2_ASAP7_75t_SL g2080 ( 
.A(n_1869),
.B(n_1685),
.Y(n_2080)
);

INVx1_ASAP7_75t_L g2081 ( 
.A(n_1786),
.Y(n_2081)
);

BUFx6f_ASAP7_75t_L g2082 ( 
.A(n_1958),
.Y(n_2082)
);

NAND2xp5_ASAP7_75t_L g2083 ( 
.A(n_1921),
.B(n_1922),
.Y(n_2083)
);

BUFx10_ASAP7_75t_L g2084 ( 
.A(n_1849),
.Y(n_2084)
);

NOR2x1p5_ASAP7_75t_L g2085 ( 
.A(n_1830),
.B(n_1719),
.Y(n_2085)
);

NAND2xp33_ASAP7_75t_SL g2086 ( 
.A(n_1986),
.B(n_1685),
.Y(n_2086)
);

INVx2_ASAP7_75t_L g2087 ( 
.A(n_1798),
.Y(n_2087)
);

NAND2xp33_ASAP7_75t_SL g2088 ( 
.A(n_1998),
.B(n_1685),
.Y(n_2088)
);

INVx1_ASAP7_75t_L g2089 ( 
.A(n_1808),
.Y(n_2089)
);

INVx1_ASAP7_75t_L g2090 ( 
.A(n_1808),
.Y(n_2090)
);

NAND2xp5_ASAP7_75t_SL g2091 ( 
.A(n_1815),
.B(n_1705),
.Y(n_2091)
);

AND2x2_ASAP7_75t_L g2092 ( 
.A(n_1965),
.B(n_1719),
.Y(n_2092)
);

AND2x2_ASAP7_75t_L g2093 ( 
.A(n_1972),
.B(n_1719),
.Y(n_2093)
);

INVx1_ASAP7_75t_L g2094 ( 
.A(n_1816),
.Y(n_2094)
);

AOI22xp33_ASAP7_75t_L g2095 ( 
.A1(n_1857),
.A2(n_1517),
.B1(n_1513),
.B2(n_1618),
.Y(n_2095)
);

INVx3_ASAP7_75t_L g2096 ( 
.A(n_1816),
.Y(n_2096)
);

INVx3_ASAP7_75t_L g2097 ( 
.A(n_1824),
.Y(n_2097)
);

INVx5_ASAP7_75t_L g2098 ( 
.A(n_1726),
.Y(n_2098)
);

INVxp33_ASAP7_75t_L g2099 ( 
.A(n_1890),
.Y(n_2099)
);

OAI22xp33_ASAP7_75t_L g2100 ( 
.A1(n_1869),
.A2(n_1749),
.B1(n_1742),
.B2(n_1730),
.Y(n_2100)
);

INVx4_ASAP7_75t_L g2101 ( 
.A(n_1958),
.Y(n_2101)
);

AND2x2_ASAP7_75t_L g2102 ( 
.A(n_1973),
.B(n_1719),
.Y(n_2102)
);

NOR2xp33_ASAP7_75t_L g2103 ( 
.A(n_1762),
.B(n_1699),
.Y(n_2103)
);

OR2x2_ASAP7_75t_L g2104 ( 
.A(n_1736),
.B(n_1702),
.Y(n_2104)
);

INVx3_ASAP7_75t_L g2105 ( 
.A(n_1824),
.Y(n_2105)
);

INVx1_ASAP7_75t_L g2106 ( 
.A(n_1836),
.Y(n_2106)
);

INVx1_ASAP7_75t_L g2107 ( 
.A(n_1862),
.Y(n_2107)
);

INVx2_ASAP7_75t_L g2108 ( 
.A(n_1862),
.Y(n_2108)
);

BUFx3_ASAP7_75t_L g2109 ( 
.A(n_1792),
.Y(n_2109)
);

BUFx6f_ASAP7_75t_SL g2110 ( 
.A(n_1882),
.Y(n_2110)
);

NAND2xp5_ASAP7_75t_L g2111 ( 
.A(n_1923),
.B(n_1618),
.Y(n_2111)
);

INVx1_ASAP7_75t_L g2112 ( 
.A(n_1888),
.Y(n_2112)
);

AND2x2_ASAP7_75t_L g2113 ( 
.A(n_1737),
.B(n_1703),
.Y(n_2113)
);

NAND2xp5_ASAP7_75t_SL g2114 ( 
.A(n_1873),
.B(n_1705),
.Y(n_2114)
);

AOI22xp33_ASAP7_75t_L g2115 ( 
.A1(n_1840),
.A2(n_1517),
.B1(n_1513),
.B2(n_1620),
.Y(n_2115)
);

NOR2xp33_ASAP7_75t_L g2116 ( 
.A(n_1763),
.B(n_1703),
.Y(n_2116)
);

NAND2xp5_ASAP7_75t_SL g2117 ( 
.A(n_1873),
.B(n_1705),
.Y(n_2117)
);

BUFx6f_ASAP7_75t_L g2118 ( 
.A(n_1938),
.Y(n_2118)
);

INVx2_ASAP7_75t_L g2119 ( 
.A(n_1888),
.Y(n_2119)
);

AND2x2_ASAP7_75t_L g2120 ( 
.A(n_1926),
.B(n_1709),
.Y(n_2120)
);

BUFx4f_ASAP7_75t_L g2121 ( 
.A(n_1882),
.Y(n_2121)
);

INVxp67_ASAP7_75t_SL g2122 ( 
.A(n_1930),
.Y(n_2122)
);

INVx1_ASAP7_75t_L g2123 ( 
.A(n_1896),
.Y(n_2123)
);

INVx3_ASAP7_75t_L g2124 ( 
.A(n_1902),
.Y(n_2124)
);

INVx1_ASAP7_75t_L g2125 ( 
.A(n_1902),
.Y(n_2125)
);

INVx2_ASAP7_75t_L g2126 ( 
.A(n_1906),
.Y(n_2126)
);

AND2x2_ASAP7_75t_L g2127 ( 
.A(n_1781),
.B(n_1667),
.Y(n_2127)
);

INVx2_ASAP7_75t_L g2128 ( 
.A(n_1906),
.Y(n_2128)
);

INVx2_ASAP7_75t_L g2129 ( 
.A(n_1919),
.Y(n_2129)
);

INVx2_ASAP7_75t_L g2130 ( 
.A(n_1925),
.Y(n_2130)
);

INVx2_ASAP7_75t_L g2131 ( 
.A(n_1810),
.Y(n_2131)
);

AND2x6_ASAP7_75t_L g2132 ( 
.A(n_1811),
.B(n_1964),
.Y(n_2132)
);

NAND2xp5_ASAP7_75t_SL g2133 ( 
.A(n_1878),
.B(n_1675),
.Y(n_2133)
);

INVx1_ASAP7_75t_L g2134 ( 
.A(n_1812),
.Y(n_2134)
);

NAND2xp5_ASAP7_75t_L g2135 ( 
.A(n_1781),
.B(n_1620),
.Y(n_2135)
);

INVx3_ASAP7_75t_L g2136 ( 
.A(n_1946),
.Y(n_2136)
);

INVx1_ASAP7_75t_L g2137 ( 
.A(n_1819),
.Y(n_2137)
);

OAI22xp33_ASAP7_75t_L g2138 ( 
.A1(n_1767),
.A2(n_1675),
.B1(n_1710),
.B2(n_1676),
.Y(n_2138)
);

INVx1_ASAP7_75t_L g2139 ( 
.A(n_1823),
.Y(n_2139)
);

NAND2xp5_ASAP7_75t_SL g2140 ( 
.A(n_1769),
.B(n_1676),
.Y(n_2140)
);

AND2x2_ASAP7_75t_L g2141 ( 
.A(n_1799),
.B(n_1710),
.Y(n_2141)
);

AOI22xp5_ASAP7_75t_L g2142 ( 
.A1(n_1741),
.A2(n_1715),
.B1(n_1712),
.B2(n_1620),
.Y(n_2142)
);

INVx2_ASAP7_75t_L g2143 ( 
.A(n_1827),
.Y(n_2143)
);

INVx2_ASAP7_75t_L g2144 ( 
.A(n_1842),
.Y(n_2144)
);

INVx1_ASAP7_75t_L g2145 ( 
.A(n_1844),
.Y(n_2145)
);

INVxp67_ASAP7_75t_SL g2146 ( 
.A(n_1871),
.Y(n_2146)
);

AND2x2_ASAP7_75t_SL g2147 ( 
.A(n_1971),
.B(n_1666),
.Y(n_2147)
);

AND2x2_ASAP7_75t_L g2148 ( 
.A(n_1799),
.B(n_1712),
.Y(n_2148)
);

INVx1_ASAP7_75t_L g2149 ( 
.A(n_1845),
.Y(n_2149)
);

INVx1_ASAP7_75t_L g2150 ( 
.A(n_1853),
.Y(n_2150)
);

INVx2_ASAP7_75t_SL g2151 ( 
.A(n_1948),
.Y(n_2151)
);

NAND2xp5_ASAP7_75t_L g2152 ( 
.A(n_1822),
.B(n_1620),
.Y(n_2152)
);

INVx1_ASAP7_75t_L g2153 ( 
.A(n_1854),
.Y(n_2153)
);

NAND2xp5_ASAP7_75t_L g2154 ( 
.A(n_1726),
.B(n_1640),
.Y(n_2154)
);

INVx1_ASAP7_75t_SL g2155 ( 
.A(n_1883),
.Y(n_2155)
);

NAND2xp5_ASAP7_75t_SL g2156 ( 
.A(n_1760),
.B(n_1715),
.Y(n_2156)
);

INVx1_ASAP7_75t_L g2157 ( 
.A(n_1874),
.Y(n_2157)
);

NAND2xp5_ASAP7_75t_SL g2158 ( 
.A(n_1766),
.B(n_1666),
.Y(n_2158)
);

AOI22xp33_ASAP7_75t_L g2159 ( 
.A1(n_1746),
.A2(n_1517),
.B1(n_1513),
.B2(n_1640),
.Y(n_2159)
);

INVx1_ASAP7_75t_L g2160 ( 
.A(n_1877),
.Y(n_2160)
);

BUFx10_ASAP7_75t_L g2161 ( 
.A(n_1849),
.Y(n_2161)
);

INVx3_ASAP7_75t_L g2162 ( 
.A(n_1947),
.Y(n_2162)
);

INVx2_ASAP7_75t_L g2163 ( 
.A(n_1881),
.Y(n_2163)
);

NAND2xp5_ASAP7_75t_L g2164 ( 
.A(n_1866),
.B(n_1640),
.Y(n_2164)
);

INVx3_ASAP7_75t_L g2165 ( 
.A(n_1949),
.Y(n_2165)
);

AOI22xp5_ASAP7_75t_L g2166 ( 
.A1(n_1940),
.A2(n_1653),
.B1(n_1664),
.B2(n_1528),
.Y(n_2166)
);

NOR2xp33_ASAP7_75t_L g2167 ( 
.A(n_1725),
.B(n_1666),
.Y(n_2167)
);

INVx1_ASAP7_75t_SL g2168 ( 
.A(n_1987),
.Y(n_2168)
);

INVx3_ASAP7_75t_L g2169 ( 
.A(n_1951),
.Y(n_2169)
);

INVx3_ASAP7_75t_L g2170 ( 
.A(n_1961),
.Y(n_2170)
);

NAND2xp5_ASAP7_75t_SL g2171 ( 
.A(n_1776),
.B(n_1666),
.Y(n_2171)
);

NAND2xp33_ASAP7_75t_L g2172 ( 
.A(n_1916),
.B(n_1513),
.Y(n_2172)
);

HB1xp67_ASAP7_75t_L g2173 ( 
.A(n_1739),
.Y(n_2173)
);

NOR2xp33_ASAP7_75t_SL g2174 ( 
.A(n_1895),
.B(n_1671),
.Y(n_2174)
);

INVx1_ASAP7_75t_L g2175 ( 
.A(n_1887),
.Y(n_2175)
);

NAND3xp33_ASAP7_75t_L g2176 ( 
.A(n_1790),
.B(n_1467),
.C(n_1581),
.Y(n_2176)
);

NAND2xp5_ASAP7_75t_SL g2177 ( 
.A(n_1778),
.B(n_1686),
.Y(n_2177)
);

INVx2_ASAP7_75t_L g2178 ( 
.A(n_1901),
.Y(n_2178)
);

AND2x6_ASAP7_75t_L g2179 ( 
.A(n_1964),
.B(n_1528),
.Y(n_2179)
);

NOR2xp33_ASAP7_75t_L g2180 ( 
.A(n_1731),
.B(n_1698),
.Y(n_2180)
);

INVx1_ASAP7_75t_L g2181 ( 
.A(n_1735),
.Y(n_2181)
);

INVx3_ASAP7_75t_L g2182 ( 
.A(n_1982),
.Y(n_2182)
);

BUFx2_ASAP7_75t_L g2183 ( 
.A(n_1739),
.Y(n_2183)
);

NAND2xp5_ASAP7_75t_L g2184 ( 
.A(n_1847),
.B(n_1650),
.Y(n_2184)
);

INVx3_ASAP7_75t_L g2185 ( 
.A(n_1984),
.Y(n_2185)
);

INVx1_ASAP7_75t_L g2186 ( 
.A(n_1740),
.Y(n_2186)
);

NAND2xp5_ASAP7_75t_L g2187 ( 
.A(n_1860),
.B(n_1650),
.Y(n_2187)
);

NAND2xp5_ASAP7_75t_L g2188 ( 
.A(n_1870),
.B(n_1446),
.Y(n_2188)
);

BUFx2_ASAP7_75t_L g2189 ( 
.A(n_1848),
.Y(n_2189)
);

AOI22xp5_ASAP7_75t_L g2190 ( 
.A1(n_1738),
.A2(n_1592),
.B1(n_1617),
.B2(n_1594),
.Y(n_2190)
);

NAND2xp5_ASAP7_75t_L g2191 ( 
.A(n_1884),
.B(n_1444),
.Y(n_2191)
);

INVx1_ASAP7_75t_L g2192 ( 
.A(n_1780),
.Y(n_2192)
);

INVx3_ASAP7_75t_L g2193 ( 
.A(n_1993),
.Y(n_2193)
);

OA22x2_ASAP7_75t_L g2194 ( 
.A1(n_1944),
.A2(n_1549),
.B1(n_1553),
.B2(n_1547),
.Y(n_2194)
);

CKINVDCx5p33_ASAP7_75t_R g2195 ( 
.A(n_1777),
.Y(n_2195)
);

INVxp33_ASAP7_75t_L g2196 ( 
.A(n_1899),
.Y(n_2196)
);

INVx1_ASAP7_75t_L g2197 ( 
.A(n_1791),
.Y(n_2197)
);

INVx1_ASAP7_75t_L g2198 ( 
.A(n_1802),
.Y(n_2198)
);

NOR2x1p5_ASAP7_75t_L g2199 ( 
.A(n_1864),
.B(n_1671),
.Y(n_2199)
);

AND2x2_ASAP7_75t_L g2200 ( 
.A(n_1745),
.B(n_1619),
.Y(n_2200)
);

INVx2_ASAP7_75t_L g2201 ( 
.A(n_1807),
.Y(n_2201)
);

OR2x2_ASAP7_75t_L g2202 ( 
.A(n_1848),
.B(n_1681),
.Y(n_2202)
);

INVx1_ASAP7_75t_L g2203 ( 
.A(n_1974),
.Y(n_2203)
);

NAND2xp5_ASAP7_75t_SL g2204 ( 
.A(n_1800),
.B(n_1805),
.Y(n_2204)
);

OAI22xp5_ASAP7_75t_L g2205 ( 
.A1(n_1809),
.A2(n_1487),
.B1(n_1494),
.B2(n_1641),
.Y(n_2205)
);

CKINVDCx5p33_ASAP7_75t_R g2206 ( 
.A(n_1814),
.Y(n_2206)
);

INVx1_ASAP7_75t_L g2207 ( 
.A(n_1975),
.Y(n_2207)
);

INVx1_ASAP7_75t_L g2208 ( 
.A(n_1948),
.Y(n_2208)
);

AND2x2_ASAP7_75t_L g2209 ( 
.A(n_1745),
.B(n_1619),
.Y(n_2209)
);

INVx1_ASAP7_75t_L g2210 ( 
.A(n_1974),
.Y(n_2210)
);

AND2x4_ASAP7_75t_L g2211 ( 
.A(n_1835),
.B(n_1547),
.Y(n_2211)
);

NOR2xp33_ASAP7_75t_L g2212 ( 
.A(n_1825),
.B(n_1704),
.Y(n_2212)
);

NOR2xp33_ASAP7_75t_L g2213 ( 
.A(n_1832),
.B(n_1716),
.Y(n_2213)
);

INVx6_ASAP7_75t_L g2214 ( 
.A(n_1932),
.Y(n_2214)
);

OR2x6_ASAP7_75t_L g2215 ( 
.A(n_1838),
.B(n_1645),
.Y(n_2215)
);

INVxp33_ASAP7_75t_SL g2216 ( 
.A(n_1806),
.Y(n_2216)
);

NAND2xp5_ASAP7_75t_L g2217 ( 
.A(n_1914),
.B(n_1444),
.Y(n_2217)
);

AOI22xp33_ASAP7_75t_L g2218 ( 
.A1(n_1910),
.A2(n_1517),
.B1(n_1513),
.B2(n_1549),
.Y(n_2218)
);

NAND2xp5_ASAP7_75t_L g2219 ( 
.A(n_1936),
.B(n_1447),
.Y(n_2219)
);

INVx1_ASAP7_75t_L g2220 ( 
.A(n_1928),
.Y(n_2220)
);

AND2x6_ASAP7_75t_L g2221 ( 
.A(n_1970),
.B(n_1553),
.Y(n_2221)
);

BUFx6f_ASAP7_75t_L g2222 ( 
.A(n_1932),
.Y(n_2222)
);

NAND2xp5_ASAP7_75t_SL g2223 ( 
.A(n_1817),
.B(n_1686),
.Y(n_2223)
);

INVx2_ASAP7_75t_L g2224 ( 
.A(n_1966),
.Y(n_2224)
);

AND2x6_ASAP7_75t_L g2225 ( 
.A(n_1970),
.B(n_1556),
.Y(n_2225)
);

NAND2xp5_ASAP7_75t_SL g2226 ( 
.A(n_1818),
.B(n_1686),
.Y(n_2226)
);

INVx1_ASAP7_75t_L g2227 ( 
.A(n_1935),
.Y(n_2227)
);

INVx2_ASAP7_75t_L g2228 ( 
.A(n_1966),
.Y(n_2228)
);

INVx2_ASAP7_75t_SL g2229 ( 
.A(n_1839),
.Y(n_2229)
);

BUFx10_ASAP7_75t_L g2230 ( 
.A(n_1753),
.Y(n_2230)
);

CKINVDCx20_ASAP7_75t_R g2231 ( 
.A(n_1756),
.Y(n_2231)
);

INVx1_ASAP7_75t_SL g2232 ( 
.A(n_1904),
.Y(n_2232)
);

NAND2x1p5_ASAP7_75t_L g2233 ( 
.A(n_1977),
.B(n_1451),
.Y(n_2233)
);

INVx1_ASAP7_75t_L g2234 ( 
.A(n_1945),
.Y(n_2234)
);

AOI22xp33_ASAP7_75t_L g2235 ( 
.A1(n_1910),
.A2(n_1517),
.B1(n_1560),
.B2(n_1556),
.Y(n_2235)
);

INVx1_ASAP7_75t_L g2236 ( 
.A(n_1967),
.Y(n_2236)
);

OAI22xp33_ASAP7_75t_L g2237 ( 
.A1(n_1855),
.A2(n_1686),
.B1(n_1561),
.B2(n_1563),
.Y(n_2237)
);

INVxp67_ASAP7_75t_SL g2238 ( 
.A(n_1937),
.Y(n_2238)
);

INVx1_ASAP7_75t_L g2239 ( 
.A(n_1967),
.Y(n_2239)
);

BUFx2_ASAP7_75t_L g2240 ( 
.A(n_1793),
.Y(n_2240)
);

NOR2xp33_ASAP7_75t_L g2241 ( 
.A(n_1880),
.B(n_1665),
.Y(n_2241)
);

CKINVDCx5p33_ASAP7_75t_R g2242 ( 
.A(n_1814),
.Y(n_2242)
);

INVx1_ASAP7_75t_L g2243 ( 
.A(n_1969),
.Y(n_2243)
);

INVx4_ASAP7_75t_L g2244 ( 
.A(n_1969),
.Y(n_2244)
);

INVx1_ASAP7_75t_L g2245 ( 
.A(n_1915),
.Y(n_2245)
);

BUFx4f_ASAP7_75t_L g2246 ( 
.A(n_1867),
.Y(n_2246)
);

OAI22xp33_ASAP7_75t_L g2247 ( 
.A1(n_1892),
.A2(n_1898),
.B1(n_1856),
.B2(n_1876),
.Y(n_2247)
);

NAND2xp5_ASAP7_75t_L g2248 ( 
.A(n_1852),
.B(n_1447),
.Y(n_2248)
);

BUFx6f_ASAP7_75t_L g2249 ( 
.A(n_1868),
.Y(n_2249)
);

NOR2xp33_ASAP7_75t_L g2250 ( 
.A(n_1794),
.B(n_1665),
.Y(n_2250)
);

AND2x2_ASAP7_75t_L g2251 ( 
.A(n_1752),
.B(n_1521),
.Y(n_2251)
);

INVx1_ASAP7_75t_L g2252 ( 
.A(n_1988),
.Y(n_2252)
);

INVx1_ASAP7_75t_L g2253 ( 
.A(n_1915),
.Y(n_2253)
);

INVx1_ASAP7_75t_L g2254 ( 
.A(n_1917),
.Y(n_2254)
);

AND2x4_ASAP7_75t_L g2255 ( 
.A(n_1879),
.B(n_1560),
.Y(n_2255)
);

NAND2xp5_ASAP7_75t_SL g2256 ( 
.A(n_1912),
.B(n_1686),
.Y(n_2256)
);

AND2x4_ASAP7_75t_L g2257 ( 
.A(n_1981),
.B(n_1561),
.Y(n_2257)
);

BUFx8_ASAP7_75t_SL g2258 ( 
.A(n_1793),
.Y(n_2258)
);

NAND2xp5_ASAP7_75t_SL g2259 ( 
.A(n_1821),
.B(n_1494),
.Y(n_2259)
);

INVx3_ASAP7_75t_L g2260 ( 
.A(n_1893),
.Y(n_2260)
);

INVx2_ASAP7_75t_L g2261 ( 
.A(n_1988),
.Y(n_2261)
);

OA22x2_ASAP7_75t_L g2262 ( 
.A1(n_1955),
.A2(n_1573),
.B1(n_1590),
.B2(n_1563),
.Y(n_2262)
);

NAND2xp5_ASAP7_75t_L g2263 ( 
.A(n_1908),
.B(n_1466),
.Y(n_2263)
);

INVx1_ASAP7_75t_L g2264 ( 
.A(n_1997),
.Y(n_2264)
);

INVx3_ASAP7_75t_L g2265 ( 
.A(n_1886),
.Y(n_2265)
);

NAND2xp5_ASAP7_75t_SL g2266 ( 
.A(n_1907),
.B(n_1494),
.Y(n_2266)
);

INVx3_ASAP7_75t_L g2267 ( 
.A(n_1997),
.Y(n_2267)
);

OAI22xp5_ASAP7_75t_SL g2268 ( 
.A1(n_1828),
.A2(n_1623),
.B1(n_1681),
.B2(n_1516),
.Y(n_2268)
);

BUFx3_ASAP7_75t_L g2269 ( 
.A(n_1959),
.Y(n_2269)
);

INVx2_ASAP7_75t_L g2270 ( 
.A(n_1752),
.Y(n_2270)
);

INVx2_ASAP7_75t_L g2271 ( 
.A(n_1917),
.Y(n_2271)
);

INVx2_ASAP7_75t_L g2272 ( 
.A(n_1733),
.Y(n_2272)
);

AND2x2_ASAP7_75t_L g2273 ( 
.A(n_1733),
.B(n_1521),
.Y(n_2273)
);

INVx3_ASAP7_75t_L g2274 ( 
.A(n_1953),
.Y(n_2274)
);

NOR2xp33_ASAP7_75t_L g2275 ( 
.A(n_1773),
.B(n_1645),
.Y(n_2275)
);

INVx4_ASAP7_75t_SL g2276 ( 
.A(n_2221),
.Y(n_2276)
);

AND2x4_ASAP7_75t_L g2277 ( 
.A(n_2229),
.B(n_1573),
.Y(n_2277)
);

BUFx4f_ASAP7_75t_L g2278 ( 
.A(n_2060),
.Y(n_2278)
);

INVx1_ASAP7_75t_L g2279 ( 
.A(n_2036),
.Y(n_2279)
);

BUFx6f_ASAP7_75t_L g2280 ( 
.A(n_2007),
.Y(n_2280)
);

AND2x4_ASAP7_75t_L g2281 ( 
.A(n_2229),
.B(n_1590),
.Y(n_2281)
);

BUFx6f_ASAP7_75t_L g2282 ( 
.A(n_2007),
.Y(n_2282)
);

BUFx2_ASAP7_75t_L g2283 ( 
.A(n_2013),
.Y(n_2283)
);

CKINVDCx5p33_ASAP7_75t_R g2284 ( 
.A(n_2010),
.Y(n_2284)
);

BUFx2_ASAP7_75t_L g2285 ( 
.A(n_2155),
.Y(n_2285)
);

INVx1_ASAP7_75t_L g2286 ( 
.A(n_2039),
.Y(n_2286)
);

BUFx3_ASAP7_75t_L g2287 ( 
.A(n_2010),
.Y(n_2287)
);

INVx1_ASAP7_75t_L g2288 ( 
.A(n_2039),
.Y(n_2288)
);

CKINVDCx5p33_ASAP7_75t_R g2289 ( 
.A(n_2258),
.Y(n_2289)
);

INVx1_ASAP7_75t_L g2290 ( 
.A(n_2054),
.Y(n_2290)
);

NAND2xp5_ASAP7_75t_SL g2291 ( 
.A(n_2006),
.B(n_1920),
.Y(n_2291)
);

AND2x4_ASAP7_75t_L g2292 ( 
.A(n_2211),
.B(n_1601),
.Y(n_2292)
);

BUFx6f_ASAP7_75t_L g2293 ( 
.A(n_2007),
.Y(n_2293)
);

INVx2_ASAP7_75t_SL g2294 ( 
.A(n_2168),
.Y(n_2294)
);

AND2x4_ASAP7_75t_L g2295 ( 
.A(n_2211),
.B(n_1601),
.Y(n_2295)
);

AND2x6_ASAP7_75t_L g2296 ( 
.A(n_2118),
.B(n_1978),
.Y(n_2296)
);

NAND2xp5_ASAP7_75t_L g2297 ( 
.A(n_2002),
.B(n_1498),
.Y(n_2297)
);

INVx1_ASAP7_75t_L g2298 ( 
.A(n_2054),
.Y(n_2298)
);

NAND2xp5_ASAP7_75t_SL g2299 ( 
.A(n_2006),
.B(n_1787),
.Y(n_2299)
);

NAND3xp33_ASAP7_75t_L g2300 ( 
.A(n_2212),
.B(n_2241),
.C(n_2075),
.Y(n_2300)
);

NAND2x1p5_ASAP7_75t_L g2301 ( 
.A(n_2098),
.B(n_1494),
.Y(n_2301)
);

INVxp67_ASAP7_75t_L g2302 ( 
.A(n_2046),
.Y(n_2302)
);

INVx1_ASAP7_75t_L g2303 ( 
.A(n_2058),
.Y(n_2303)
);

HB1xp67_ASAP7_75t_L g2304 ( 
.A(n_2127),
.Y(n_2304)
);

INVx1_ASAP7_75t_L g2305 ( 
.A(n_2058),
.Y(n_2305)
);

AND2x4_ASAP7_75t_L g2306 ( 
.A(n_2255),
.B(n_1606),
.Y(n_2306)
);

AND2x6_ASAP7_75t_L g2307 ( 
.A(n_2118),
.B(n_1980),
.Y(n_2307)
);

BUFx2_ASAP7_75t_L g2308 ( 
.A(n_2047),
.Y(n_2308)
);

AND2x2_ASAP7_75t_L g2309 ( 
.A(n_2005),
.B(n_1894),
.Y(n_2309)
);

INVxp67_ASAP7_75t_SL g2310 ( 
.A(n_2007),
.Y(n_2310)
);

BUFx6f_ASAP7_75t_L g2311 ( 
.A(n_2007),
.Y(n_2311)
);

CKINVDCx16_ASAP7_75t_R g2312 ( 
.A(n_2268),
.Y(n_2312)
);

INVx1_ASAP7_75t_L g2313 ( 
.A(n_2067),
.Y(n_2313)
);

INVx1_ASAP7_75t_L g2314 ( 
.A(n_2073),
.Y(n_2314)
);

OAI22xp33_ASAP7_75t_SL g2315 ( 
.A1(n_2156),
.A2(n_1761),
.B1(n_1841),
.B2(n_1829),
.Y(n_2315)
);

NAND2xp5_ASAP7_75t_L g2316 ( 
.A(n_2008),
.B(n_2009),
.Y(n_2316)
);

AND2x2_ASAP7_75t_SL g2317 ( 
.A(n_2080),
.B(n_1968),
.Y(n_2317)
);

INVx1_ASAP7_75t_L g2318 ( 
.A(n_2078),
.Y(n_2318)
);

INVx1_ASAP7_75t_L g2319 ( 
.A(n_2078),
.Y(n_2319)
);

CKINVDCx5p33_ASAP7_75t_R g2320 ( 
.A(n_2258),
.Y(n_2320)
);

AOI22xp33_ASAP7_75t_L g2321 ( 
.A1(n_2080),
.A2(n_1801),
.B1(n_1956),
.B2(n_1953),
.Y(n_2321)
);

INVx4_ASAP7_75t_L g2322 ( 
.A(n_2035),
.Y(n_2322)
);

AND2x2_ASAP7_75t_L g2323 ( 
.A(n_2005),
.B(n_1894),
.Y(n_2323)
);

NOR2xp33_ASAP7_75t_L g2324 ( 
.A(n_2099),
.B(n_1858),
.Y(n_2324)
);

BUFx2_ASAP7_75t_L g2325 ( 
.A(n_2047),
.Y(n_2325)
);

BUFx6f_ASAP7_75t_L g2326 ( 
.A(n_2082),
.Y(n_2326)
);

INVx2_ASAP7_75t_L g2327 ( 
.A(n_2016),
.Y(n_2327)
);

AOI22xp5_ASAP7_75t_L g2328 ( 
.A1(n_2103),
.A2(n_1889),
.B1(n_1612),
.B2(n_1613),
.Y(n_2328)
);

BUFx6f_ASAP7_75t_L g2329 ( 
.A(n_2082),
.Y(n_2329)
);

INVx1_ASAP7_75t_L g2330 ( 
.A(n_2079),
.Y(n_2330)
);

INVx1_ASAP7_75t_L g2331 ( 
.A(n_2087),
.Y(n_2331)
);

AND2x4_ASAP7_75t_L g2332 ( 
.A(n_2255),
.B(n_1609),
.Y(n_2332)
);

BUFx12f_ASAP7_75t_L g2333 ( 
.A(n_2018),
.Y(n_2333)
);

BUFx2_ASAP7_75t_L g2334 ( 
.A(n_2104),
.Y(n_2334)
);

AND2x2_ASAP7_75t_L g2335 ( 
.A(n_2046),
.B(n_1764),
.Y(n_2335)
);

AND2x4_ASAP7_75t_L g2336 ( 
.A(n_2255),
.B(n_1609),
.Y(n_2336)
);

AO22x2_ASAP7_75t_L g2337 ( 
.A1(n_2244),
.A2(n_1956),
.B1(n_1960),
.B2(n_1976),
.Y(n_2337)
);

AND2x4_ASAP7_75t_L g2338 ( 
.A(n_2249),
.B(n_2141),
.Y(n_2338)
);

NOR2xp33_ASAP7_75t_L g2339 ( 
.A(n_2232),
.B(n_1911),
.Y(n_2339)
);

INVx2_ASAP7_75t_SL g2340 ( 
.A(n_2104),
.Y(n_2340)
);

AND2x4_ASAP7_75t_L g2341 ( 
.A(n_2249),
.B(n_1612),
.Y(n_2341)
);

AND2x2_ASAP7_75t_L g2342 ( 
.A(n_2048),
.B(n_2065),
.Y(n_2342)
);

NAND2xp5_ASAP7_75t_L g2343 ( 
.A(n_2120),
.B(n_1466),
.Y(n_2343)
);

INVx1_ASAP7_75t_L g2344 ( 
.A(n_2108),
.Y(n_2344)
);

NAND2xp5_ASAP7_75t_L g2345 ( 
.A(n_2120),
.B(n_1477),
.Y(n_2345)
);

NAND3xp33_ASAP7_75t_SL g2346 ( 
.A(n_2027),
.B(n_2041),
.C(n_2037),
.Y(n_2346)
);

INVx1_ASAP7_75t_L g2347 ( 
.A(n_2108),
.Y(n_2347)
);

AND2x6_ASAP7_75t_L g2348 ( 
.A(n_2118),
.B(n_1968),
.Y(n_2348)
);

BUFx3_ASAP7_75t_L g2349 ( 
.A(n_2109),
.Y(n_2349)
);

INVx1_ASAP7_75t_L g2350 ( 
.A(n_2119),
.Y(n_2350)
);

NAND2xp5_ASAP7_75t_SL g2351 ( 
.A(n_2118),
.B(n_1487),
.Y(n_2351)
);

NAND2xp5_ASAP7_75t_SL g2352 ( 
.A(n_2118),
.B(n_1487),
.Y(n_2352)
);

AO21x2_ASAP7_75t_L g2353 ( 
.A1(n_2133),
.A2(n_1499),
.B(n_1491),
.Y(n_2353)
);

OAI22xp5_ASAP7_75t_L g2354 ( 
.A1(n_2012),
.A2(n_1957),
.B1(n_1952),
.B2(n_1954),
.Y(n_2354)
);

INVx3_ASAP7_75t_L g2355 ( 
.A(n_2082),
.Y(n_2355)
);

INVx5_ASAP7_75t_L g2356 ( 
.A(n_2132),
.Y(n_2356)
);

HB1xp67_ASAP7_75t_L g2357 ( 
.A(n_2127),
.Y(n_2357)
);

BUFx3_ASAP7_75t_L g2358 ( 
.A(n_2109),
.Y(n_2358)
);

AO22x2_ASAP7_75t_L g2359 ( 
.A1(n_2244),
.A2(n_1960),
.B1(n_1983),
.B2(n_1872),
.Y(n_2359)
);

NAND2xp5_ASAP7_75t_L g2360 ( 
.A(n_2093),
.B(n_1477),
.Y(n_2360)
);

NOR2xp33_ASAP7_75t_L g2361 ( 
.A(n_2196),
.B(n_1516),
.Y(n_2361)
);

INVxp67_ASAP7_75t_L g2362 ( 
.A(n_2048),
.Y(n_2362)
);

BUFx3_ASAP7_75t_L g2363 ( 
.A(n_2249),
.Y(n_2363)
);

INVx4_ASAP7_75t_L g2364 ( 
.A(n_2035),
.Y(n_2364)
);

AND2x2_ASAP7_75t_L g2365 ( 
.A(n_2180),
.B(n_1764),
.Y(n_2365)
);

CKINVDCx16_ASAP7_75t_R g2366 ( 
.A(n_2174),
.Y(n_2366)
);

INVx2_ASAP7_75t_L g2367 ( 
.A(n_2019),
.Y(n_2367)
);

INVx1_ASAP7_75t_L g2368 ( 
.A(n_2126),
.Y(n_2368)
);

NOR2xp33_ASAP7_75t_L g2369 ( 
.A(n_2116),
.B(n_1897),
.Y(n_2369)
);

NAND3x1_ASAP7_75t_L g2370 ( 
.A(n_2274),
.B(n_1833),
.C(n_1771),
.Y(n_2370)
);

INVx2_ASAP7_75t_L g2371 ( 
.A(n_2019),
.Y(n_2371)
);

INVx1_ASAP7_75t_L g2372 ( 
.A(n_2126),
.Y(n_2372)
);

INVx2_ASAP7_75t_L g2373 ( 
.A(n_2024),
.Y(n_2373)
);

NAND2xp5_ASAP7_75t_L g2374 ( 
.A(n_2093),
.B(n_1482),
.Y(n_2374)
);

INVx1_ASAP7_75t_L g2375 ( 
.A(n_2128),
.Y(n_2375)
);

INVx2_ASAP7_75t_L g2376 ( 
.A(n_2024),
.Y(n_2376)
);

INVx4_ASAP7_75t_L g2377 ( 
.A(n_2035),
.Y(n_2377)
);

INVx1_ASAP7_75t_SL g2378 ( 
.A(n_2202),
.Y(n_2378)
);

INVx1_ASAP7_75t_L g2379 ( 
.A(n_2128),
.Y(n_2379)
);

INVx1_ASAP7_75t_L g2380 ( 
.A(n_2014),
.Y(n_2380)
);

INVx2_ASAP7_75t_L g2381 ( 
.A(n_2029),
.Y(n_2381)
);

OAI22xp33_ASAP7_75t_L g2382 ( 
.A1(n_2194),
.A2(n_1994),
.B1(n_1999),
.B2(n_1992),
.Y(n_2382)
);

INVx2_ASAP7_75t_L g2383 ( 
.A(n_2029),
.Y(n_2383)
);

AO22x2_ASAP7_75t_L g2384 ( 
.A1(n_2244),
.A2(n_1991),
.B1(n_1996),
.B2(n_1743),
.Y(n_2384)
);

INVxp67_ASAP7_75t_L g2385 ( 
.A(n_2092),
.Y(n_2385)
);

INVx2_ASAP7_75t_L g2386 ( 
.A(n_2014),
.Y(n_2386)
);

BUFx2_ASAP7_75t_L g2387 ( 
.A(n_2202),
.Y(n_2387)
);

NOR2xp33_ASAP7_75t_L g2388 ( 
.A(n_2063),
.B(n_1900),
.Y(n_2388)
);

AND2x4_ASAP7_75t_L g2389 ( 
.A(n_2249),
.B(n_2141),
.Y(n_2389)
);

INVx4_ASAP7_75t_L g2390 ( 
.A(n_2082),
.Y(n_2390)
);

INVx2_ASAP7_75t_L g2391 ( 
.A(n_2015),
.Y(n_2391)
);

NOR2xp33_ASAP7_75t_L g2392 ( 
.A(n_2113),
.B(n_1891),
.Y(n_2392)
);

AND2x2_ASAP7_75t_L g2393 ( 
.A(n_2113),
.B(n_1775),
.Y(n_2393)
);

AND2x4_ASAP7_75t_L g2394 ( 
.A(n_2249),
.B(n_1613),
.Y(n_2394)
);

INVxp67_ASAP7_75t_SL g2395 ( 
.A(n_2203),
.Y(n_2395)
);

INVx2_ASAP7_75t_L g2396 ( 
.A(n_2033),
.Y(n_2396)
);

INVx1_ASAP7_75t_L g2397 ( 
.A(n_2015),
.Y(n_2397)
);

NOR2xp33_ASAP7_75t_L g2398 ( 
.A(n_2167),
.B(n_1913),
.Y(n_2398)
);

INVx1_ASAP7_75t_SL g2399 ( 
.A(n_2183),
.Y(n_2399)
);

AO22x2_ASAP7_75t_L g2400 ( 
.A1(n_2236),
.A2(n_1743),
.B1(n_1754),
.B2(n_1775),
.Y(n_2400)
);

AND2x2_ASAP7_75t_L g2401 ( 
.A(n_2092),
.B(n_1783),
.Y(n_2401)
);

INVx1_ASAP7_75t_L g2402 ( 
.A(n_2017),
.Y(n_2402)
);

NOR2xp33_ASAP7_75t_L g2403 ( 
.A(n_2213),
.B(n_1467),
.Y(n_2403)
);

OAI22xp5_ASAP7_75t_SL g2404 ( 
.A1(n_2231),
.A2(n_1645),
.B1(n_1467),
.B2(n_1990),
.Y(n_2404)
);

INVx2_ASAP7_75t_L g2405 ( 
.A(n_2129),
.Y(n_2405)
);

AND2x6_ASAP7_75t_L g2406 ( 
.A(n_2267),
.B(n_2000),
.Y(n_2406)
);

INVx1_ASAP7_75t_L g2407 ( 
.A(n_2017),
.Y(n_2407)
);

AND2x2_ASAP7_75t_L g2408 ( 
.A(n_2148),
.B(n_2207),
.Y(n_2408)
);

OR2x6_ASAP7_75t_L g2409 ( 
.A(n_2060),
.B(n_1645),
.Y(n_2409)
);

AND2x4_ASAP7_75t_L g2410 ( 
.A(n_2148),
.B(n_1614),
.Y(n_2410)
);

AND2x4_ASAP7_75t_L g2411 ( 
.A(n_2257),
.B(n_1614),
.Y(n_2411)
);

INVx4_ASAP7_75t_SL g2412 ( 
.A(n_2221),
.Y(n_2412)
);

NAND2xp5_ASAP7_75t_L g2413 ( 
.A(n_2102),
.B(n_1482),
.Y(n_2413)
);

INVx2_ASAP7_75t_L g2414 ( 
.A(n_2129),
.Y(n_2414)
);

INVx2_ASAP7_75t_L g2415 ( 
.A(n_2130),
.Y(n_2415)
);

CKINVDCx16_ASAP7_75t_R g2416 ( 
.A(n_2018),
.Y(n_2416)
);

INVx2_ASAP7_75t_SL g2417 ( 
.A(n_2269),
.Y(n_2417)
);

CKINVDCx5p33_ASAP7_75t_R g2418 ( 
.A(n_2195),
.Y(n_2418)
);

HB1xp67_ASAP7_75t_L g2419 ( 
.A(n_2043),
.Y(n_2419)
);

NOR2xp33_ASAP7_75t_R g2420 ( 
.A(n_2086),
.B(n_1581),
.Y(n_2420)
);

BUFx6f_ASAP7_75t_L g2421 ( 
.A(n_2025),
.Y(n_2421)
);

AND2x4_ASAP7_75t_L g2422 ( 
.A(n_2257),
.B(n_1625),
.Y(n_2422)
);

NAND2x1p5_ASAP7_75t_L g2423 ( 
.A(n_2098),
.B(n_1480),
.Y(n_2423)
);

INVx1_ASAP7_75t_L g2424 ( 
.A(n_2026),
.Y(n_2424)
);

INVxp67_ASAP7_75t_L g2425 ( 
.A(n_2102),
.Y(n_2425)
);

NAND3xp33_ASAP7_75t_L g2426 ( 
.A(n_2052),
.B(n_1581),
.C(n_1627),
.Y(n_2426)
);

INVx5_ASAP7_75t_L g2427 ( 
.A(n_2132),
.Y(n_2427)
);

INVxp67_ASAP7_75t_L g2428 ( 
.A(n_2273),
.Y(n_2428)
);

OR2x2_ASAP7_75t_L g2429 ( 
.A(n_2183),
.B(n_1627),
.Y(n_2429)
);

BUFx6f_ASAP7_75t_L g2430 ( 
.A(n_2025),
.Y(n_2430)
);

INVx1_ASAP7_75t_L g2431 ( 
.A(n_2042),
.Y(n_2431)
);

INVx1_ASAP7_75t_L g2432 ( 
.A(n_2044),
.Y(n_2432)
);

AND2x4_ASAP7_75t_L g2433 ( 
.A(n_2257),
.B(n_1632),
.Y(n_2433)
);

INVx2_ASAP7_75t_L g2434 ( 
.A(n_2044),
.Y(n_2434)
);

INVx1_ASAP7_75t_L g2435 ( 
.A(n_2050),
.Y(n_2435)
);

INVx3_ASAP7_75t_L g2436 ( 
.A(n_2011),
.Y(n_2436)
);

INVx2_ASAP7_75t_L g2437 ( 
.A(n_2050),
.Y(n_2437)
);

INVx2_ASAP7_75t_L g2438 ( 
.A(n_2053),
.Y(n_2438)
);

NAND2xp5_ASAP7_75t_SL g2439 ( 
.A(n_2098),
.B(n_1592),
.Y(n_2439)
);

BUFx3_ASAP7_75t_L g2440 ( 
.A(n_2121),
.Y(n_2440)
);

AND2x4_ASAP7_75t_L g2441 ( 
.A(n_2085),
.B(n_1638),
.Y(n_2441)
);

INVx2_ASAP7_75t_L g2442 ( 
.A(n_2056),
.Y(n_2442)
);

NAND2x1p5_ASAP7_75t_L g2443 ( 
.A(n_2098),
.B(n_1480),
.Y(n_2443)
);

BUFx3_ASAP7_75t_L g2444 ( 
.A(n_2121),
.Y(n_2444)
);

AND2x4_ASAP7_75t_L g2445 ( 
.A(n_2038),
.B(n_2043),
.Y(n_2445)
);

INVx1_ASAP7_75t_L g2446 ( 
.A(n_2056),
.Y(n_2446)
);

AND2x4_ASAP7_75t_L g2447 ( 
.A(n_2038),
.B(n_1638),
.Y(n_2447)
);

INVx1_ASAP7_75t_L g2448 ( 
.A(n_2062),
.Y(n_2448)
);

AND2x6_ASAP7_75t_L g2449 ( 
.A(n_2267),
.B(n_1588),
.Y(n_2449)
);

INVx2_ASAP7_75t_L g2450 ( 
.A(n_2130),
.Y(n_2450)
);

AND2x2_ASAP7_75t_L g2451 ( 
.A(n_2200),
.B(n_1788),
.Y(n_2451)
);

NOR2xp33_ASAP7_75t_L g2452 ( 
.A(n_2100),
.B(n_1918),
.Y(n_2452)
);

OR2x2_ASAP7_75t_SL g2453 ( 
.A(n_2176),
.B(n_1588),
.Y(n_2453)
);

BUFx2_ASAP7_75t_L g2454 ( 
.A(n_2189),
.Y(n_2454)
);

BUFx3_ASAP7_75t_L g2455 ( 
.A(n_2121),
.Y(n_2455)
);

AND2x2_ASAP7_75t_SL g2456 ( 
.A(n_2147),
.B(n_1596),
.Y(n_2456)
);

HB1xp67_ASAP7_75t_L g2457 ( 
.A(n_2267),
.Y(n_2457)
);

INVx1_ASAP7_75t_L g2458 ( 
.A(n_2066),
.Y(n_2458)
);

INVx2_ASAP7_75t_SL g2459 ( 
.A(n_2173),
.Y(n_2459)
);

INVx1_ASAP7_75t_L g2460 ( 
.A(n_2066),
.Y(n_2460)
);

INVxp67_ASAP7_75t_L g2461 ( 
.A(n_2273),
.Y(n_2461)
);

INVx2_ASAP7_75t_L g2462 ( 
.A(n_2131),
.Y(n_2462)
);

INVx1_ASAP7_75t_L g2463 ( 
.A(n_2081),
.Y(n_2463)
);

BUFx12f_ASAP7_75t_L g2464 ( 
.A(n_2018),
.Y(n_2464)
);

INVx1_ASAP7_75t_L g2465 ( 
.A(n_2106),
.Y(n_2465)
);

INVx1_ASAP7_75t_L g2466 ( 
.A(n_2106),
.Y(n_2466)
);

BUFx6f_ASAP7_75t_L g2467 ( 
.A(n_2021),
.Y(n_2467)
);

INVx2_ASAP7_75t_L g2468 ( 
.A(n_2143),
.Y(n_2468)
);

INVx1_ASAP7_75t_L g2469 ( 
.A(n_2107),
.Y(n_2469)
);

BUFx2_ASAP7_75t_L g2470 ( 
.A(n_2189),
.Y(n_2470)
);

NOR2xp33_ASAP7_75t_L g2471 ( 
.A(n_2049),
.B(n_1846),
.Y(n_2471)
);

INVx1_ASAP7_75t_L g2472 ( 
.A(n_2123),
.Y(n_2472)
);

INVx1_ASAP7_75t_L g2473 ( 
.A(n_2123),
.Y(n_2473)
);

INVx2_ASAP7_75t_L g2474 ( 
.A(n_2143),
.Y(n_2474)
);

CKINVDCx5p33_ASAP7_75t_R g2475 ( 
.A(n_2110),
.Y(n_2475)
);

INVx2_ASAP7_75t_L g2476 ( 
.A(n_2125),
.Y(n_2476)
);

NAND2x1_ASAP7_75t_L g2477 ( 
.A(n_2021),
.B(n_1451),
.Y(n_2477)
);

INVx1_ASAP7_75t_L g2478 ( 
.A(n_2004),
.Y(n_2478)
);

BUFx6f_ASAP7_75t_L g2479 ( 
.A(n_2021),
.Y(n_2479)
);

INVx2_ASAP7_75t_L g2480 ( 
.A(n_2096),
.Y(n_2480)
);

INVx1_ASAP7_75t_L g2481 ( 
.A(n_2023),
.Y(n_2481)
);

NAND2xp5_ASAP7_75t_SL g2482 ( 
.A(n_2098),
.B(n_1592),
.Y(n_2482)
);

INVx4_ASAP7_75t_L g2483 ( 
.A(n_2032),
.Y(n_2483)
);

INVx2_ASAP7_75t_L g2484 ( 
.A(n_2381),
.Y(n_2484)
);

NAND2x1p5_ASAP7_75t_L g2485 ( 
.A(n_2322),
.B(n_2032),
.Y(n_2485)
);

BUFx3_ASAP7_75t_L g2486 ( 
.A(n_2287),
.Y(n_2486)
);

NOR2xp33_ASAP7_75t_L g2487 ( 
.A(n_2300),
.B(n_2051),
.Y(n_2487)
);

INVx2_ASAP7_75t_L g2488 ( 
.A(n_2381),
.Y(n_2488)
);

BUFx6f_ASAP7_75t_L g2489 ( 
.A(n_2287),
.Y(n_2489)
);

INVx1_ASAP7_75t_L g2490 ( 
.A(n_2457),
.Y(n_2490)
);

NAND2xp5_ASAP7_75t_L g2491 ( 
.A(n_2316),
.B(n_2069),
.Y(n_2491)
);

AOI22xp33_ASAP7_75t_L g2492 ( 
.A1(n_2369),
.A2(n_2247),
.B1(n_2262),
.B2(n_2204),
.Y(n_2492)
);

NAND2xp5_ASAP7_75t_L g2493 ( 
.A(n_2316),
.B(n_2069),
.Y(n_2493)
);

NAND2xp5_ASAP7_75t_L g2494 ( 
.A(n_2302),
.B(n_2074),
.Y(n_2494)
);

NAND2xp5_ASAP7_75t_SL g2495 ( 
.A(n_2338),
.B(n_2246),
.Y(n_2495)
);

BUFx6f_ASAP7_75t_L g2496 ( 
.A(n_2421),
.Y(n_2496)
);

INVx2_ASAP7_75t_L g2497 ( 
.A(n_2383),
.Y(n_2497)
);

NAND2xp5_ASAP7_75t_L g2498 ( 
.A(n_2302),
.B(n_2074),
.Y(n_2498)
);

NAND2xp5_ASAP7_75t_L g2499 ( 
.A(n_2362),
.B(n_2270),
.Y(n_2499)
);

NAND2xp5_ASAP7_75t_SL g2500 ( 
.A(n_2338),
.B(n_2389),
.Y(n_2500)
);

INVx2_ASAP7_75t_L g2501 ( 
.A(n_2383),
.Y(n_2501)
);

AND2x4_ASAP7_75t_L g2502 ( 
.A(n_2440),
.B(n_2215),
.Y(n_2502)
);

NAND2xp5_ASAP7_75t_SL g2503 ( 
.A(n_2389),
.B(n_2246),
.Y(n_2503)
);

INVx2_ASAP7_75t_SL g2504 ( 
.A(n_2284),
.Y(n_2504)
);

INVx1_ASAP7_75t_L g2505 ( 
.A(n_2457),
.Y(n_2505)
);

NAND2xp5_ASAP7_75t_SL g2506 ( 
.A(n_2294),
.B(n_2315),
.Y(n_2506)
);

NAND2xp5_ASAP7_75t_SL g2507 ( 
.A(n_2403),
.B(n_2222),
.Y(n_2507)
);

NAND2xp5_ASAP7_75t_L g2508 ( 
.A(n_2342),
.B(n_2209),
.Y(n_2508)
);

NOR2xp33_ASAP7_75t_L g2509 ( 
.A(n_2324),
.B(n_2216),
.Y(n_2509)
);

NAND3xp33_ASAP7_75t_L g2510 ( 
.A(n_2398),
.B(n_2022),
.C(n_2250),
.Y(n_2510)
);

INVx1_ASAP7_75t_L g2511 ( 
.A(n_2395),
.Y(n_2511)
);

NAND2xp5_ASAP7_75t_L g2512 ( 
.A(n_2304),
.B(n_2357),
.Y(n_2512)
);

CKINVDCx5p33_ASAP7_75t_R g2513 ( 
.A(n_2418),
.Y(n_2513)
);

NAND2xp5_ASAP7_75t_L g2514 ( 
.A(n_2357),
.B(n_2251),
.Y(n_2514)
);

NAND2xp5_ASAP7_75t_L g2515 ( 
.A(n_2392),
.B(n_2271),
.Y(n_2515)
);

NAND3xp33_ASAP7_75t_L g2516 ( 
.A(n_2398),
.B(n_2275),
.C(n_2166),
.Y(n_2516)
);

INVx1_ASAP7_75t_L g2517 ( 
.A(n_2478),
.Y(n_2517)
);

INVx1_ASAP7_75t_L g2518 ( 
.A(n_2481),
.Y(n_2518)
);

NAND2xp5_ASAP7_75t_L g2519 ( 
.A(n_2385),
.B(n_2271),
.Y(n_2519)
);

NAND2xp5_ASAP7_75t_L g2520 ( 
.A(n_2408),
.B(n_2138),
.Y(n_2520)
);

NAND2xp5_ASAP7_75t_L g2521 ( 
.A(n_2419),
.B(n_2245),
.Y(n_2521)
);

NAND2xp5_ASAP7_75t_SL g2522 ( 
.A(n_2366),
.B(n_2222),
.Y(n_2522)
);

NAND2xp5_ASAP7_75t_L g2523 ( 
.A(n_2419),
.B(n_2362),
.Y(n_2523)
);

NAND2xp5_ASAP7_75t_L g2524 ( 
.A(n_2393),
.B(n_2253),
.Y(n_2524)
);

NAND2xp5_ASAP7_75t_L g2525 ( 
.A(n_2388),
.B(n_2254),
.Y(n_2525)
);

NAND2xp5_ASAP7_75t_L g2526 ( 
.A(n_2388),
.B(n_2072),
.Y(n_2526)
);

NAND2xp5_ASAP7_75t_SL g2527 ( 
.A(n_2410),
.B(n_2222),
.Y(n_2527)
);

INVx2_ASAP7_75t_SL g2528 ( 
.A(n_2349),
.Y(n_2528)
);

NAND2xp5_ASAP7_75t_L g2529 ( 
.A(n_2471),
.B(n_2272),
.Y(n_2529)
);

HB1xp67_ASAP7_75t_L g2530 ( 
.A(n_2283),
.Y(n_2530)
);

NAND2xp5_ASAP7_75t_L g2531 ( 
.A(n_2471),
.B(n_2272),
.Y(n_2531)
);

NAND3xp33_ASAP7_75t_L g2532 ( 
.A(n_2452),
.B(n_2140),
.C(n_2142),
.Y(n_2532)
);

INVx2_ASAP7_75t_L g2533 ( 
.A(n_2327),
.Y(n_2533)
);

INVx2_ASAP7_75t_SL g2534 ( 
.A(n_2349),
.Y(n_2534)
);

NAND2xp5_ASAP7_75t_L g2535 ( 
.A(n_2425),
.B(n_2270),
.Y(n_2535)
);

AOI22xp33_ASAP7_75t_SL g2536 ( 
.A1(n_2359),
.A2(n_2216),
.B1(n_2262),
.B2(n_2231),
.Y(n_2536)
);

NAND2xp5_ASAP7_75t_L g2537 ( 
.A(n_2425),
.B(n_2274),
.Y(n_2537)
);

INVxp33_ASAP7_75t_SL g2538 ( 
.A(n_2289),
.Y(n_2538)
);

AOI22xp33_ASAP7_75t_L g2539 ( 
.A1(n_2346),
.A2(n_2262),
.B1(n_2194),
.B2(n_2147),
.Y(n_2539)
);

BUFx6f_ASAP7_75t_L g2540 ( 
.A(n_2421),
.Y(n_2540)
);

INVxp67_ASAP7_75t_L g2541 ( 
.A(n_2285),
.Y(n_2541)
);

BUFx6f_ASAP7_75t_L g2542 ( 
.A(n_2421),
.Y(n_2542)
);

NAND2xp5_ASAP7_75t_L g2543 ( 
.A(n_2401),
.B(n_2274),
.Y(n_2543)
);

INVx1_ASAP7_75t_L g2544 ( 
.A(n_2431),
.Y(n_2544)
);

OR2x2_ASAP7_75t_L g2545 ( 
.A(n_2378),
.B(n_2240),
.Y(n_2545)
);

INVxp67_ASAP7_75t_SL g2546 ( 
.A(n_2310),
.Y(n_2546)
);

AOI22xp33_ASAP7_75t_L g2547 ( 
.A1(n_2346),
.A2(n_2194),
.B1(n_2265),
.B2(n_2064),
.Y(n_2547)
);

NAND2xp5_ASAP7_75t_L g2548 ( 
.A(n_2343),
.B(n_2221),
.Y(n_2548)
);

NAND2xp5_ASAP7_75t_SL g2549 ( 
.A(n_2410),
.B(n_2222),
.Y(n_2549)
);

AOI21xp5_ASAP7_75t_L g2550 ( 
.A1(n_2291),
.A2(n_2003),
.B(n_2086),
.Y(n_2550)
);

INVx2_ASAP7_75t_L g2551 ( 
.A(n_2327),
.Y(n_2551)
);

AOI22xp5_ASAP7_75t_L g2552 ( 
.A1(n_2361),
.A2(n_2158),
.B1(n_2266),
.B2(n_2240),
.Y(n_2552)
);

AOI21xp5_ASAP7_75t_L g2553 ( 
.A1(n_2291),
.A2(n_2088),
.B(n_2083),
.Y(n_2553)
);

INVx2_ASAP7_75t_L g2554 ( 
.A(n_2367),
.Y(n_2554)
);

INVx1_ASAP7_75t_L g2555 ( 
.A(n_2432),
.Y(n_2555)
);

OAI221xp5_ASAP7_75t_L g2556 ( 
.A1(n_2339),
.A2(n_2321),
.B1(n_2328),
.B2(n_2361),
.C(n_2299),
.Y(n_2556)
);

AND2x2_ASAP7_75t_L g2557 ( 
.A(n_2365),
.B(n_1981),
.Y(n_2557)
);

INVx1_ASAP7_75t_L g2558 ( 
.A(n_2435),
.Y(n_2558)
);

NAND2x1p5_ASAP7_75t_L g2559 ( 
.A(n_2322),
.B(n_2070),
.Y(n_2559)
);

AND2x6_ASAP7_75t_SL g2560 ( 
.A(n_2339),
.B(n_2060),
.Y(n_2560)
);

NAND2xp5_ASAP7_75t_L g2561 ( 
.A(n_2343),
.B(n_2236),
.Y(n_2561)
);

NOR2xp33_ASAP7_75t_L g2562 ( 
.A(n_2428),
.B(n_2222),
.Y(n_2562)
);

AOI22xp33_ASAP7_75t_L g2563 ( 
.A1(n_2317),
.A2(n_2265),
.B1(n_2225),
.B2(n_2221),
.Y(n_2563)
);

NAND2xp5_ASAP7_75t_SL g2564 ( 
.A(n_2292),
.B(n_2230),
.Y(n_2564)
);

NAND2xp5_ASAP7_75t_L g2565 ( 
.A(n_2345),
.B(n_2239),
.Y(n_2565)
);

AND2x2_ASAP7_75t_L g2566 ( 
.A(n_2309),
.B(n_1754),
.Y(n_2566)
);

INVx2_ASAP7_75t_SL g2567 ( 
.A(n_2358),
.Y(n_2567)
);

INVx2_ASAP7_75t_SL g2568 ( 
.A(n_2358),
.Y(n_2568)
);

NOR2xp33_ASAP7_75t_L g2569 ( 
.A(n_2428),
.B(n_2214),
.Y(n_2569)
);

NAND2xp5_ASAP7_75t_L g2570 ( 
.A(n_2345),
.B(n_2239),
.Y(n_2570)
);

NAND2xp5_ASAP7_75t_L g2571 ( 
.A(n_2360),
.B(n_2243),
.Y(n_2571)
);

AND2x2_ASAP7_75t_L g2572 ( 
.A(n_2323),
.B(n_1843),
.Y(n_2572)
);

NAND2x1p5_ASAP7_75t_L g2573 ( 
.A(n_2364),
.B(n_2070),
.Y(n_2573)
);

NAND2xp5_ASAP7_75t_L g2574 ( 
.A(n_2360),
.B(n_2243),
.Y(n_2574)
);

BUFx6f_ASAP7_75t_L g2575 ( 
.A(n_2421),
.Y(n_2575)
);

NOR2xp33_ASAP7_75t_L g2576 ( 
.A(n_2461),
.B(n_2214),
.Y(n_2576)
);

INVx2_ASAP7_75t_L g2577 ( 
.A(n_2367),
.Y(n_2577)
);

NAND2xp5_ASAP7_75t_L g2578 ( 
.A(n_2374),
.B(n_2252),
.Y(n_2578)
);

INVx2_ASAP7_75t_SL g2579 ( 
.A(n_2387),
.Y(n_2579)
);

A2O1A1Ixp33_ASAP7_75t_L g2580 ( 
.A1(n_2299),
.A2(n_2088),
.B(n_2263),
.C(n_2248),
.Y(n_2580)
);

NAND2xp5_ASAP7_75t_L g2581 ( 
.A(n_2374),
.B(n_2413),
.Y(n_2581)
);

NAND2xp5_ASAP7_75t_SL g2582 ( 
.A(n_2292),
.B(n_2230),
.Y(n_2582)
);

NAND2xp5_ASAP7_75t_SL g2583 ( 
.A(n_2295),
.B(n_2230),
.Y(n_2583)
);

AOI21xp5_ASAP7_75t_L g2584 ( 
.A1(n_2297),
.A2(n_2061),
.B(n_2020),
.Y(n_2584)
);

INVx2_ASAP7_75t_L g2585 ( 
.A(n_2371),
.Y(n_2585)
);

A2O1A1Ixp33_ASAP7_75t_L g2586 ( 
.A1(n_2456),
.A2(n_2171),
.B(n_2259),
.C(n_2265),
.Y(n_2586)
);

NAND2xp5_ASAP7_75t_L g2587 ( 
.A(n_2413),
.B(n_2252),
.Y(n_2587)
);

AND2x2_ASAP7_75t_L g2588 ( 
.A(n_2451),
.B(n_1863),
.Y(n_2588)
);

INVx1_ASAP7_75t_L g2589 ( 
.A(n_2446),
.Y(n_2589)
);

NOR2xp33_ASAP7_75t_L g2590 ( 
.A(n_2461),
.B(n_2214),
.Y(n_2590)
);

OR2x6_ASAP7_75t_L g2591 ( 
.A(n_2364),
.B(n_2071),
.Y(n_2591)
);

NOR2xp33_ASAP7_75t_L g2592 ( 
.A(n_2308),
.B(n_2214),
.Y(n_2592)
);

OR2x6_ASAP7_75t_L g2593 ( 
.A(n_2377),
.B(n_2071),
.Y(n_2593)
);

NAND2xp5_ASAP7_75t_L g2594 ( 
.A(n_2386),
.B(n_2391),
.Y(n_2594)
);

NAND2xp5_ASAP7_75t_L g2595 ( 
.A(n_2335),
.B(n_2221),
.Y(n_2595)
);

INVx1_ASAP7_75t_L g2596 ( 
.A(n_2448),
.Y(n_2596)
);

INVx1_ASAP7_75t_L g2597 ( 
.A(n_2458),
.Y(n_2597)
);

NAND2xp5_ASAP7_75t_L g2598 ( 
.A(n_2386),
.B(n_2264),
.Y(n_2598)
);

NAND2xp5_ASAP7_75t_L g2599 ( 
.A(n_2445),
.B(n_2221),
.Y(n_2599)
);

BUFx6f_ASAP7_75t_L g2600 ( 
.A(n_2430),
.Y(n_2600)
);

NAND2xp5_ASAP7_75t_L g2601 ( 
.A(n_2445),
.B(n_2225),
.Y(n_2601)
);

BUFx6f_ASAP7_75t_L g2602 ( 
.A(n_2430),
.Y(n_2602)
);

INVx1_ASAP7_75t_L g2603 ( 
.A(n_2460),
.Y(n_2603)
);

NOR2xp33_ASAP7_75t_L g2604 ( 
.A(n_2325),
.B(n_2334),
.Y(n_2604)
);

NAND2xp33_ASAP7_75t_L g2605 ( 
.A(n_2467),
.B(n_2225),
.Y(n_2605)
);

NAND2xp5_ASAP7_75t_L g2606 ( 
.A(n_2391),
.B(n_2264),
.Y(n_2606)
);

AND2x4_ASAP7_75t_L g2607 ( 
.A(n_2440),
.B(n_2215),
.Y(n_2607)
);

INVx2_ASAP7_75t_SL g2608 ( 
.A(n_2340),
.Y(n_2608)
);

INVx8_ASAP7_75t_L g2609 ( 
.A(n_2449),
.Y(n_2609)
);

NAND2xp5_ASAP7_75t_L g2610 ( 
.A(n_2297),
.B(n_2225),
.Y(n_2610)
);

O2A1O1Ixp33_ASAP7_75t_L g2611 ( 
.A1(n_2382),
.A2(n_2001),
.B(n_2237),
.C(n_1851),
.Y(n_2611)
);

NAND2xp5_ASAP7_75t_L g2612 ( 
.A(n_2380),
.B(n_2224),
.Y(n_2612)
);

NAND2xp5_ASAP7_75t_L g2613 ( 
.A(n_2397),
.B(n_2224),
.Y(n_2613)
);

INVx4_ASAP7_75t_L g2614 ( 
.A(n_2467),
.Y(n_2614)
);

NAND2xp5_ASAP7_75t_SL g2615 ( 
.A(n_2295),
.B(n_2034),
.Y(n_2615)
);

AND2x6_ASAP7_75t_L g2616 ( 
.A(n_2480),
.B(n_2228),
.Y(n_2616)
);

INVx1_ASAP7_75t_L g2617 ( 
.A(n_2463),
.Y(n_2617)
);

NAND2xp5_ASAP7_75t_L g2618 ( 
.A(n_2402),
.B(n_2228),
.Y(n_2618)
);

O2A1O1Ixp33_ASAP7_75t_L g2619 ( 
.A1(n_2382),
.A2(n_1875),
.B(n_1850),
.C(n_2260),
.Y(n_2619)
);

NOR2xp33_ASAP7_75t_L g2620 ( 
.A(n_2399),
.B(n_2260),
.Y(n_2620)
);

NAND2xp5_ASAP7_75t_L g2621 ( 
.A(n_2407),
.B(n_2261),
.Y(n_2621)
);

AOI22xp5_ASAP7_75t_L g2622 ( 
.A1(n_2404),
.A2(n_2260),
.B1(n_2215),
.B2(n_2256),
.Y(n_2622)
);

HB1xp67_ASAP7_75t_L g2623 ( 
.A(n_2454),
.Y(n_2623)
);

AND2x2_ASAP7_75t_L g2624 ( 
.A(n_2306),
.B(n_2071),
.Y(n_2624)
);

NOR2xp33_ASAP7_75t_L g2625 ( 
.A(n_2429),
.B(n_2208),
.Y(n_2625)
);

NAND2xp5_ASAP7_75t_L g2626 ( 
.A(n_2306),
.B(n_2261),
.Y(n_2626)
);

NAND3xp33_ASAP7_75t_L g2627 ( 
.A(n_2426),
.B(n_2159),
.C(n_2235),
.Y(n_2627)
);

INVx1_ASAP7_75t_L g2628 ( 
.A(n_2465),
.Y(n_2628)
);

NAND2xp5_ASAP7_75t_L g2629 ( 
.A(n_2332),
.B(n_2217),
.Y(n_2629)
);

AOI22xp5_ASAP7_75t_L g2630 ( 
.A1(n_2456),
.A2(n_2199),
.B1(n_2110),
.B2(n_2076),
.Y(n_2630)
);

NAND2xp5_ASAP7_75t_SL g2631 ( 
.A(n_2332),
.B(n_2034),
.Y(n_2631)
);

OR2x2_ASAP7_75t_L g2632 ( 
.A(n_2470),
.B(n_2175),
.Y(n_2632)
);

NAND2xp5_ASAP7_75t_L g2633 ( 
.A(n_2336),
.B(n_2219),
.Y(n_2633)
);

CKINVDCx5p33_ASAP7_75t_R g2634 ( 
.A(n_2320),
.Y(n_2634)
);

NAND2xp5_ASAP7_75t_L g2635 ( 
.A(n_2336),
.B(n_2122),
.Y(n_2635)
);

NAND2xp5_ASAP7_75t_L g2636 ( 
.A(n_2277),
.B(n_2191),
.Y(n_2636)
);

AND2x2_ASAP7_75t_L g2637 ( 
.A(n_2359),
.B(n_2071),
.Y(n_2637)
);

INVx3_ASAP7_75t_L g2638 ( 
.A(n_2467),
.Y(n_2638)
);

INVx1_ASAP7_75t_L g2639 ( 
.A(n_2466),
.Y(n_2639)
);

AOI22xp5_ASAP7_75t_L g2640 ( 
.A1(n_2441),
.A2(n_2091),
.B1(n_2117),
.B2(n_2114),
.Y(n_2640)
);

NAND2xp33_ASAP7_75t_L g2641 ( 
.A(n_2467),
.B(n_2179),
.Y(n_2641)
);

NAND2xp5_ASAP7_75t_SL g2642 ( 
.A(n_2411),
.B(n_2034),
.Y(n_2642)
);

OR2x2_ASAP7_75t_L g2643 ( 
.A(n_2459),
.B(n_2077),
.Y(n_2643)
);

XNOR2xp5_ASAP7_75t_L g2644 ( 
.A(n_2370),
.B(n_2206),
.Y(n_2644)
);

NAND2x1p5_ASAP7_75t_L g2645 ( 
.A(n_2377),
.B(n_2101),
.Y(n_2645)
);

AOI221x1_ASAP7_75t_L g2646 ( 
.A1(n_2384),
.A2(n_2152),
.B1(n_2205),
.B2(n_2164),
.C(n_1934),
.Y(n_2646)
);

NAND2xp5_ASAP7_75t_L g2647 ( 
.A(n_2281),
.B(n_2341),
.Y(n_2647)
);

BUFx6f_ASAP7_75t_L g2648 ( 
.A(n_2430),
.Y(n_2648)
);

O2A1O1Ixp5_ASAP7_75t_L g2649 ( 
.A1(n_2354),
.A2(n_2031),
.B(n_2045),
.C(n_2177),
.Y(n_2649)
);

NOR2xp33_ASAP7_75t_L g2650 ( 
.A(n_2417),
.B(n_2077),
.Y(n_2650)
);

NAND2xp5_ASAP7_75t_L g2651 ( 
.A(n_2341),
.B(n_2394),
.Y(n_2651)
);

AOI22xp33_ASAP7_75t_L g2652 ( 
.A1(n_2317),
.A2(n_2132),
.B1(n_2059),
.B2(n_2030),
.Y(n_2652)
);

NOR2xp33_ASAP7_75t_L g2653 ( 
.A(n_2411),
.B(n_2077),
.Y(n_2653)
);

INVxp67_ASAP7_75t_L g2654 ( 
.A(n_2422),
.Y(n_2654)
);

INVx1_ASAP7_75t_L g2655 ( 
.A(n_2469),
.Y(n_2655)
);

AND2x2_ASAP7_75t_SL g2656 ( 
.A(n_2563),
.B(n_2278),
.Y(n_2656)
);

INVx2_ASAP7_75t_L g2657 ( 
.A(n_2484),
.Y(n_2657)
);

INVx1_ASAP7_75t_SL g2658 ( 
.A(n_2545),
.Y(n_2658)
);

NAND2xp5_ASAP7_75t_SL g2659 ( 
.A(n_2487),
.B(n_2356),
.Y(n_2659)
);

INVx1_ASAP7_75t_L g2660 ( 
.A(n_2517),
.Y(n_2660)
);

INVx1_ASAP7_75t_L g2661 ( 
.A(n_2518),
.Y(n_2661)
);

INVx5_ASAP7_75t_L g2662 ( 
.A(n_2591),
.Y(n_2662)
);

AOI22xp33_ASAP7_75t_L g2663 ( 
.A1(n_2492),
.A2(n_2359),
.B1(n_2337),
.B2(n_2406),
.Y(n_2663)
);

INVx4_ASAP7_75t_L g2664 ( 
.A(n_2489),
.Y(n_2664)
);

AND2x4_ASAP7_75t_L g2665 ( 
.A(n_2591),
.B(n_2444),
.Y(n_2665)
);

NAND2xp5_ASAP7_75t_L g2666 ( 
.A(n_2525),
.B(n_2422),
.Y(n_2666)
);

OR2x6_ASAP7_75t_L g2667 ( 
.A(n_2609),
.B(n_2409),
.Y(n_2667)
);

AO22x1_ASAP7_75t_L g2668 ( 
.A1(n_2509),
.A2(n_2475),
.B1(n_2242),
.B2(n_2206),
.Y(n_2668)
);

INVx2_ASAP7_75t_SL g2669 ( 
.A(n_2489),
.Y(n_2669)
);

AO22x1_ASAP7_75t_L g2670 ( 
.A1(n_2620),
.A2(n_2242),
.B1(n_2455),
.B2(n_2444),
.Y(n_2670)
);

AOI22xp33_ASAP7_75t_SL g2671 ( 
.A1(n_2556),
.A2(n_2337),
.B1(n_2348),
.B2(n_2356),
.Y(n_2671)
);

INVx4_ASAP7_75t_L g2672 ( 
.A(n_2489),
.Y(n_2672)
);

INVx2_ASAP7_75t_L g2673 ( 
.A(n_2488),
.Y(n_2673)
);

INVx1_ASAP7_75t_L g2674 ( 
.A(n_2544),
.Y(n_2674)
);

INVx2_ASAP7_75t_L g2675 ( 
.A(n_2497),
.Y(n_2675)
);

INVx2_ASAP7_75t_L g2676 ( 
.A(n_2501),
.Y(n_2676)
);

NAND2xp5_ASAP7_75t_L g2677 ( 
.A(n_2515),
.B(n_2433),
.Y(n_2677)
);

INVx1_ASAP7_75t_L g2678 ( 
.A(n_2555),
.Y(n_2678)
);

INVx1_ASAP7_75t_L g2679 ( 
.A(n_2558),
.Y(n_2679)
);

INVx2_ASAP7_75t_SL g2680 ( 
.A(n_2486),
.Y(n_2680)
);

NAND2xp5_ASAP7_75t_L g2681 ( 
.A(n_2636),
.B(n_2433),
.Y(n_2681)
);

INVx1_ASAP7_75t_SL g2682 ( 
.A(n_2530),
.Y(n_2682)
);

AOI22xp33_ASAP7_75t_L g2683 ( 
.A1(n_2526),
.A2(n_2337),
.B1(n_2406),
.B2(n_2348),
.Y(n_2683)
);

AOI22xp5_ASAP7_75t_L g2684 ( 
.A1(n_2510),
.A2(n_2296),
.B1(n_2307),
.B2(n_2312),
.Y(n_2684)
);

NAND2xp5_ASAP7_75t_L g2685 ( 
.A(n_2529),
.B(n_2394),
.Y(n_2685)
);

OR2x2_ASAP7_75t_SL g2686 ( 
.A(n_2516),
.B(n_2416),
.Y(n_2686)
);

AND2x2_ASAP7_75t_L g2687 ( 
.A(n_2588),
.B(n_2400),
.Y(n_2687)
);

INVx1_ASAP7_75t_L g2688 ( 
.A(n_2589),
.Y(n_2688)
);

INVx2_ASAP7_75t_L g2689 ( 
.A(n_2533),
.Y(n_2689)
);

INVx2_ASAP7_75t_L g2690 ( 
.A(n_2551),
.Y(n_2690)
);

BUFx3_ASAP7_75t_L g2691 ( 
.A(n_2496),
.Y(n_2691)
);

NAND2xp5_ASAP7_75t_L g2692 ( 
.A(n_2531),
.B(n_2400),
.Y(n_2692)
);

OAI22xp5_ASAP7_75t_L g2693 ( 
.A1(n_2552),
.A2(n_2427),
.B1(n_2356),
.B2(n_2278),
.Y(n_2693)
);

INVx2_ASAP7_75t_L g2694 ( 
.A(n_2554),
.Y(n_2694)
);

AND2x2_ASAP7_75t_SL g2695 ( 
.A(n_2605),
.B(n_2276),
.Y(n_2695)
);

INVx2_ASAP7_75t_L g2696 ( 
.A(n_2577),
.Y(n_2696)
);

OR2x6_ASAP7_75t_L g2697 ( 
.A(n_2609),
.B(n_2409),
.Y(n_2697)
);

NAND2xp5_ASAP7_75t_L g2698 ( 
.A(n_2629),
.B(n_2400),
.Y(n_2698)
);

OR2x6_ASAP7_75t_L g2699 ( 
.A(n_2609),
.B(n_2409),
.Y(n_2699)
);

NAND2xp5_ASAP7_75t_L g2700 ( 
.A(n_2633),
.B(n_2447),
.Y(n_2700)
);

BUFx2_ASAP7_75t_L g2701 ( 
.A(n_2623),
.Y(n_2701)
);

AND2x4_ASAP7_75t_SL g2702 ( 
.A(n_2591),
.B(n_2084),
.Y(n_2702)
);

INVx2_ASAP7_75t_L g2703 ( 
.A(n_2585),
.Y(n_2703)
);

BUFx3_ASAP7_75t_L g2704 ( 
.A(n_2496),
.Y(n_2704)
);

NOR2xp33_ASAP7_75t_L g2705 ( 
.A(n_2506),
.B(n_2356),
.Y(n_2705)
);

INVx2_ASAP7_75t_L g2706 ( 
.A(n_2596),
.Y(n_2706)
);

INVx1_ASAP7_75t_L g2707 ( 
.A(n_2597),
.Y(n_2707)
);

INVx4_ASAP7_75t_L g2708 ( 
.A(n_2496),
.Y(n_2708)
);

INVx1_ASAP7_75t_L g2709 ( 
.A(n_2603),
.Y(n_2709)
);

BUFx8_ASAP7_75t_L g2710 ( 
.A(n_2504),
.Y(n_2710)
);

OR2x6_ASAP7_75t_L g2711 ( 
.A(n_2593),
.B(n_2077),
.Y(n_2711)
);

CKINVDCx6p67_ASAP7_75t_R g2712 ( 
.A(n_2540),
.Y(n_2712)
);

AND2x4_ASAP7_75t_L g2713 ( 
.A(n_2593),
.B(n_2455),
.Y(n_2713)
);

AND2x6_ASAP7_75t_L g2714 ( 
.A(n_2622),
.B(n_2434),
.Y(n_2714)
);

NAND2xp5_ASAP7_75t_L g2715 ( 
.A(n_2508),
.B(n_2447),
.Y(n_2715)
);

AOI22xp5_ASAP7_75t_SL g2716 ( 
.A1(n_2644),
.A2(n_1963),
.B1(n_1985),
.B2(n_1939),
.Y(n_2716)
);

INVx2_ASAP7_75t_L g2717 ( 
.A(n_2617),
.Y(n_2717)
);

NAND2xp5_ASAP7_75t_SL g2718 ( 
.A(n_2507),
.B(n_2491),
.Y(n_2718)
);

INVx3_ASAP7_75t_L g2719 ( 
.A(n_2614),
.Y(n_2719)
);

NAND2xp5_ASAP7_75t_SL g2720 ( 
.A(n_2491),
.B(n_2427),
.Y(n_2720)
);

NAND2xp5_ASAP7_75t_SL g2721 ( 
.A(n_2493),
.B(n_2427),
.Y(n_2721)
);

OR2x2_ASAP7_75t_L g2722 ( 
.A(n_2524),
.B(n_2396),
.Y(n_2722)
);

BUFx6f_ASAP7_75t_L g2723 ( 
.A(n_2540),
.Y(n_2723)
);

BUFx6f_ASAP7_75t_L g2724 ( 
.A(n_2540),
.Y(n_2724)
);

AND2x6_ASAP7_75t_SL g2725 ( 
.A(n_2604),
.B(n_1593),
.Y(n_2725)
);

OAI22xp5_ASAP7_75t_L g2726 ( 
.A1(n_2539),
.A2(n_2427),
.B1(n_2190),
.B2(n_2384),
.Y(n_2726)
);

NAND2x1p5_ASAP7_75t_L g2727 ( 
.A(n_2511),
.B(n_2479),
.Y(n_2727)
);

AND2x4_ASAP7_75t_L g2728 ( 
.A(n_2502),
.B(n_2276),
.Y(n_2728)
);

BUFx6f_ASAP7_75t_L g2729 ( 
.A(n_2542),
.Y(n_2729)
);

INVx3_ASAP7_75t_L g2730 ( 
.A(n_2614),
.Y(n_2730)
);

INVx2_ASAP7_75t_L g2731 ( 
.A(n_2594),
.Y(n_2731)
);

CKINVDCx5p33_ASAP7_75t_R g2732 ( 
.A(n_2513),
.Y(n_2732)
);

AOI22xp33_ASAP7_75t_L g2733 ( 
.A1(n_2536),
.A2(n_2406),
.B1(n_2348),
.B2(n_2296),
.Y(n_2733)
);

INVxp67_ASAP7_75t_L g2734 ( 
.A(n_2625),
.Y(n_2734)
);

INVx5_ASAP7_75t_L g2735 ( 
.A(n_2542),
.Y(n_2735)
);

OAI22xp5_ASAP7_75t_L g2736 ( 
.A1(n_2630),
.A2(n_2384),
.B1(n_2453),
.B2(n_2151),
.Y(n_2736)
);

INVx1_ASAP7_75t_L g2737 ( 
.A(n_2628),
.Y(n_2737)
);

INVx1_ASAP7_75t_L g2738 ( 
.A(n_2639),
.Y(n_2738)
);

INVx2_ASAP7_75t_L g2739 ( 
.A(n_2655),
.Y(n_2739)
);

AND2x4_ASAP7_75t_L g2740 ( 
.A(n_2502),
.B(n_2276),
.Y(n_2740)
);

AOI22xp33_ASAP7_75t_L g2741 ( 
.A1(n_2532),
.A2(n_2406),
.B1(n_2348),
.B2(n_2307),
.Y(n_2741)
);

NAND2xp5_ASAP7_75t_L g2742 ( 
.A(n_2647),
.B(n_2424),
.Y(n_2742)
);

INVx2_ASAP7_75t_L g2743 ( 
.A(n_2598),
.Y(n_2743)
);

BUFx6f_ASAP7_75t_L g2744 ( 
.A(n_2542),
.Y(n_2744)
);

OR2x2_ASAP7_75t_L g2745 ( 
.A(n_2514),
.B(n_2363),
.Y(n_2745)
);

NAND2xp5_ASAP7_75t_L g2746 ( 
.A(n_2512),
.B(n_2472),
.Y(n_2746)
);

AOI22xp33_ASAP7_75t_L g2747 ( 
.A1(n_2572),
.A2(n_2406),
.B1(n_2348),
.B2(n_2307),
.Y(n_2747)
);

BUFx2_ASAP7_75t_L g2748 ( 
.A(n_2541),
.Y(n_2748)
);

BUFx8_ASAP7_75t_L g2749 ( 
.A(n_2579),
.Y(n_2749)
);

NAND2xp5_ASAP7_75t_L g2750 ( 
.A(n_2635),
.B(n_2520),
.Y(n_2750)
);

BUFx2_ASAP7_75t_L g2751 ( 
.A(n_2608),
.Y(n_2751)
);

AND2x4_ASAP7_75t_L g2752 ( 
.A(n_2607),
.B(n_2412),
.Y(n_2752)
);

BUFx4f_ASAP7_75t_L g2753 ( 
.A(n_2575),
.Y(n_2753)
);

BUFx12f_ASAP7_75t_L g2754 ( 
.A(n_2634),
.Y(n_2754)
);

AOI22xp33_ASAP7_75t_L g2755 ( 
.A1(n_2547),
.A2(n_2307),
.B1(n_2296),
.B2(n_2412),
.Y(n_2755)
);

CKINVDCx5p33_ASAP7_75t_R g2756 ( 
.A(n_2538),
.Y(n_2756)
);

AOI22xp33_ASAP7_75t_SL g2757 ( 
.A1(n_2637),
.A2(n_2296),
.B1(n_2307),
.B2(n_2420),
.Y(n_2757)
);

INVxp33_ASAP7_75t_SL g2758 ( 
.A(n_2592),
.Y(n_2758)
);

INVx2_ASAP7_75t_L g2759 ( 
.A(n_2606),
.Y(n_2759)
);

NOR2xp33_ASAP7_75t_L g2760 ( 
.A(n_2595),
.B(n_2351),
.Y(n_2760)
);

INVx1_ASAP7_75t_L g2761 ( 
.A(n_2490),
.Y(n_2761)
);

BUFx3_ASAP7_75t_L g2762 ( 
.A(n_2575),
.Y(n_2762)
);

INVx2_ASAP7_75t_L g2763 ( 
.A(n_2505),
.Y(n_2763)
);

INVx2_ASAP7_75t_L g2764 ( 
.A(n_2537),
.Y(n_2764)
);

INVx4_ASAP7_75t_L g2765 ( 
.A(n_2575),
.Y(n_2765)
);

INVx1_ASAP7_75t_L g2766 ( 
.A(n_2521),
.Y(n_2766)
);

INVx2_ASAP7_75t_SL g2767 ( 
.A(n_2528),
.Y(n_2767)
);

INVx1_ASAP7_75t_L g2768 ( 
.A(n_2523),
.Y(n_2768)
);

INVx1_ASAP7_75t_L g2769 ( 
.A(n_2519),
.Y(n_2769)
);

INVx1_ASAP7_75t_L g2770 ( 
.A(n_2612),
.Y(n_2770)
);

INVx1_ASAP7_75t_L g2771 ( 
.A(n_2612),
.Y(n_2771)
);

HB1xp67_ASAP7_75t_L g2772 ( 
.A(n_2546),
.Y(n_2772)
);

INVx1_ASAP7_75t_L g2773 ( 
.A(n_2613),
.Y(n_2773)
);

INVx2_ASAP7_75t_L g2774 ( 
.A(n_2613),
.Y(n_2774)
);

AND2x4_ASAP7_75t_L g2775 ( 
.A(n_2607),
.B(n_2412),
.Y(n_2775)
);

INVx2_ASAP7_75t_SL g2776 ( 
.A(n_2534),
.Y(n_2776)
);

INVx1_ASAP7_75t_L g2777 ( 
.A(n_2618),
.Y(n_2777)
);

CKINVDCx5p33_ASAP7_75t_R g2778 ( 
.A(n_2560),
.Y(n_2778)
);

INVx1_ASAP7_75t_L g2779 ( 
.A(n_2618),
.Y(n_2779)
);

BUFx2_ASAP7_75t_L g2780 ( 
.A(n_2654),
.Y(n_2780)
);

BUFx6f_ASAP7_75t_L g2781 ( 
.A(n_2600),
.Y(n_2781)
);

INVxp67_ASAP7_75t_L g2782 ( 
.A(n_2632),
.Y(n_2782)
);

NAND2xp5_ASAP7_75t_SL g2783 ( 
.A(n_2610),
.B(n_2420),
.Y(n_2783)
);

INVx1_ASAP7_75t_L g2784 ( 
.A(n_2621),
.Y(n_2784)
);

NAND2xp5_ASAP7_75t_SL g2785 ( 
.A(n_2581),
.B(n_2352),
.Y(n_2785)
);

INVx1_ASAP7_75t_L g2786 ( 
.A(n_2621),
.Y(n_2786)
);

INVx5_ASAP7_75t_L g2787 ( 
.A(n_2600),
.Y(n_2787)
);

NAND2xp5_ASAP7_75t_L g2788 ( 
.A(n_2581),
.B(n_2473),
.Y(n_2788)
);

INVx1_ASAP7_75t_L g2789 ( 
.A(n_2626),
.Y(n_2789)
);

INVx2_ASAP7_75t_L g2790 ( 
.A(n_2494),
.Y(n_2790)
);

INVx3_ASAP7_75t_L g2791 ( 
.A(n_2638),
.Y(n_2791)
);

BUFx4f_ASAP7_75t_L g2792 ( 
.A(n_2600),
.Y(n_2792)
);

AOI22xp33_ASAP7_75t_L g2793 ( 
.A1(n_2557),
.A2(n_1834),
.B1(n_1831),
.B2(n_1979),
.Y(n_2793)
);

INVx1_ASAP7_75t_L g2794 ( 
.A(n_2499),
.Y(n_2794)
);

NAND2xp5_ASAP7_75t_SL g2795 ( 
.A(n_2580),
.B(n_2586),
.Y(n_2795)
);

INVx1_ASAP7_75t_L g2796 ( 
.A(n_2535),
.Y(n_2796)
);

INVx4_ASAP7_75t_L g2797 ( 
.A(n_2602),
.Y(n_2797)
);

BUFx3_ASAP7_75t_L g2798 ( 
.A(n_2602),
.Y(n_2798)
);

NAND2xp5_ASAP7_75t_L g2799 ( 
.A(n_2561),
.B(n_2434),
.Y(n_2799)
);

INVxp67_ASAP7_75t_L g2800 ( 
.A(n_2543),
.Y(n_2800)
);

INVx5_ASAP7_75t_L g2801 ( 
.A(n_2602),
.Y(n_2801)
);

AOI22xp33_ASAP7_75t_L g2802 ( 
.A1(n_2566),
.A2(n_2188),
.B1(n_2449),
.B2(n_2438),
.Y(n_2802)
);

INVx1_ASAP7_75t_L g2803 ( 
.A(n_2616),
.Y(n_2803)
);

INVxp67_ASAP7_75t_L g2804 ( 
.A(n_2567),
.Y(n_2804)
);

BUFx6f_ASAP7_75t_SL g2805 ( 
.A(n_2568),
.Y(n_2805)
);

AOI22xp5_ASAP7_75t_L g2806 ( 
.A1(n_2495),
.A2(n_2057),
.B1(n_2226),
.B2(n_2223),
.Y(n_2806)
);

BUFx3_ASAP7_75t_L g2807 ( 
.A(n_2648),
.Y(n_2807)
);

INVx1_ASAP7_75t_L g2808 ( 
.A(n_2616),
.Y(n_2808)
);

HB1xp67_ASAP7_75t_L g2809 ( 
.A(n_2548),
.Y(n_2809)
);

HB1xp67_ASAP7_75t_L g2810 ( 
.A(n_2494),
.Y(n_2810)
);

NAND2x1p5_ASAP7_75t_L g2811 ( 
.A(n_2503),
.B(n_2479),
.Y(n_2811)
);

AND2x2_ASAP7_75t_SL g2812 ( 
.A(n_2641),
.B(n_2172),
.Y(n_2812)
);

INVx2_ASAP7_75t_L g2813 ( 
.A(n_2498),
.Y(n_2813)
);

BUFx4f_ASAP7_75t_SL g2814 ( 
.A(n_2522),
.Y(n_2814)
);

INVx2_ASAP7_75t_L g2815 ( 
.A(n_2571),
.Y(n_2815)
);

NAND2xp5_ASAP7_75t_L g2816 ( 
.A(n_2565),
.B(n_2437),
.Y(n_2816)
);

BUFx4f_ASAP7_75t_L g2817 ( 
.A(n_2648),
.Y(n_2817)
);

INVx3_ASAP7_75t_L g2818 ( 
.A(n_2638),
.Y(n_2818)
);

INVxp67_ASAP7_75t_L g2819 ( 
.A(n_2648),
.Y(n_2819)
);

INVx1_ASAP7_75t_L g2820 ( 
.A(n_2565),
.Y(n_2820)
);

OR2x6_ASAP7_75t_SL g2821 ( 
.A(n_2643),
.B(n_1596),
.Y(n_2821)
);

AOI21xp5_ASAP7_75t_L g2822 ( 
.A1(n_2795),
.A2(n_2584),
.B(n_2550),
.Y(n_2822)
);

O2A1O1Ixp33_ASAP7_75t_L g2823 ( 
.A1(n_2795),
.A2(n_2611),
.B(n_2619),
.C(n_2615),
.Y(n_2823)
);

AOI21xp5_ASAP7_75t_L g2824 ( 
.A1(n_2741),
.A2(n_2649),
.B(n_2553),
.Y(n_2824)
);

BUFx6f_ASAP7_75t_L g2825 ( 
.A(n_2753),
.Y(n_2825)
);

NOR2x1p5_ASAP7_75t_SL g2826 ( 
.A(n_2803),
.B(n_2373),
.Y(n_2826)
);

OAI21xp5_ASAP7_75t_L g2827 ( 
.A1(n_2734),
.A2(n_2627),
.B(n_2646),
.Y(n_2827)
);

OAI22x1_ASAP7_75t_L g2828 ( 
.A1(n_2684),
.A2(n_2631),
.B1(n_2642),
.B2(n_2640),
.Y(n_2828)
);

INVx8_ASAP7_75t_L g2829 ( 
.A(n_2735),
.Y(n_2829)
);

NAND2xp5_ASAP7_75t_SL g2830 ( 
.A(n_2734),
.B(n_2562),
.Y(n_2830)
);

O2A1O1Ixp33_ASAP7_75t_SL g2831 ( 
.A1(n_2788),
.A2(n_2549),
.B(n_2527),
.C(n_2571),
.Y(n_2831)
);

AOI21xp5_ASAP7_75t_L g2832 ( 
.A1(n_2741),
.A2(n_2482),
.B(n_2439),
.Y(n_2832)
);

INVx5_ASAP7_75t_L g2833 ( 
.A(n_2711),
.Y(n_2833)
);

OAI22xp5_ASAP7_75t_L g2834 ( 
.A1(n_2733),
.A2(n_2576),
.B1(n_2590),
.B2(n_2569),
.Y(n_2834)
);

O2A1O1Ixp33_ASAP7_75t_L g2835 ( 
.A1(n_2736),
.A2(n_2582),
.B(n_2583),
.C(n_2564),
.Y(n_2835)
);

INVx5_ASAP7_75t_L g2836 ( 
.A(n_2711),
.Y(n_2836)
);

AOI21xp5_ASAP7_75t_L g2837 ( 
.A1(n_2812),
.A2(n_2482),
.B(n_2439),
.Y(n_2837)
);

NAND2xp5_ASAP7_75t_L g2838 ( 
.A(n_2750),
.B(n_2570),
.Y(n_2838)
);

BUFx12f_ASAP7_75t_L g2839 ( 
.A(n_2732),
.Y(n_2839)
);

BUFx2_ASAP7_75t_L g2840 ( 
.A(n_2701),
.Y(n_2840)
);

NAND2xp5_ASAP7_75t_SL g2841 ( 
.A(n_2778),
.B(n_2814),
.Y(n_2841)
);

AOI21xp5_ASAP7_75t_L g2842 ( 
.A1(n_2812),
.A2(n_2301),
.B(n_2172),
.Y(n_2842)
);

NAND2xp5_ASAP7_75t_L g2843 ( 
.A(n_2658),
.B(n_2570),
.Y(n_2843)
);

OAI22xp5_ASAP7_75t_L g2844 ( 
.A1(n_2733),
.A2(n_2652),
.B1(n_2653),
.B2(n_2601),
.Y(n_2844)
);

NAND2xp5_ASAP7_75t_L g2845 ( 
.A(n_2789),
.B(n_2574),
.Y(n_2845)
);

BUFx6f_ASAP7_75t_L g2846 ( 
.A(n_2753),
.Y(n_2846)
);

AOI21xp5_ASAP7_75t_L g2847 ( 
.A1(n_2695),
.A2(n_2301),
.B(n_2310),
.Y(n_2847)
);

AOI21xp5_ASAP7_75t_L g2848 ( 
.A1(n_2695),
.A2(n_2055),
.B(n_2115),
.Y(n_2848)
);

AOI21xp5_ASAP7_75t_L g2849 ( 
.A1(n_2785),
.A2(n_2146),
.B(n_2423),
.Y(n_2849)
);

OR2x2_ASAP7_75t_L g2850 ( 
.A(n_2809),
.B(n_2599),
.Y(n_2850)
);

NAND2xp5_ASAP7_75t_L g2851 ( 
.A(n_2666),
.B(n_2574),
.Y(n_2851)
);

NAND2xp5_ASAP7_75t_L g2852 ( 
.A(n_2677),
.B(n_2578),
.Y(n_2852)
);

NAND2xp5_ASAP7_75t_L g2853 ( 
.A(n_2800),
.B(n_2578),
.Y(n_2853)
);

NAND2xp5_ASAP7_75t_SL g2854 ( 
.A(n_2814),
.B(n_2651),
.Y(n_2854)
);

AOI22xp5_ASAP7_75t_L g2855 ( 
.A1(n_2671),
.A2(n_2500),
.B1(n_2624),
.B2(n_2587),
.Y(n_2855)
);

O2A1O1Ixp33_ASAP7_75t_L g2856 ( 
.A1(n_2726),
.A2(n_2705),
.B(n_2800),
.C(n_2782),
.Y(n_2856)
);

AOI21x1_ASAP7_75t_L g2857 ( 
.A1(n_2783),
.A2(n_2587),
.B(n_2210),
.Y(n_2857)
);

BUFx4f_ASAP7_75t_L g2858 ( 
.A(n_2754),
.Y(n_2858)
);

AO32x1_ASAP7_75t_L g2859 ( 
.A1(n_2693),
.A2(n_2820),
.A3(n_2771),
.B1(n_2777),
.B2(n_2773),
.Y(n_2859)
);

BUFx3_ASAP7_75t_L g2860 ( 
.A(n_2710),
.Y(n_2860)
);

AO32x1_ASAP7_75t_L g2861 ( 
.A1(n_2770),
.A2(n_2210),
.A3(n_2203),
.B1(n_2438),
.B2(n_2437),
.Y(n_2861)
);

NAND2xp5_ASAP7_75t_L g2862 ( 
.A(n_2685),
.B(n_2650),
.Y(n_2862)
);

INVx2_ASAP7_75t_L g2863 ( 
.A(n_2739),
.Y(n_2863)
);

NOR2xp67_ASAP7_75t_L g2864 ( 
.A(n_2662),
.B(n_2279),
.Y(n_2864)
);

OR2x6_ASAP7_75t_L g2865 ( 
.A(n_2711),
.B(n_2485),
.Y(n_2865)
);

NOR2xp33_ASAP7_75t_L g2866 ( 
.A(n_2758),
.B(n_1593),
.Y(n_2866)
);

INVx2_ASAP7_75t_L g2867 ( 
.A(n_2739),
.Y(n_2867)
);

NAND2xp5_ASAP7_75t_L g2868 ( 
.A(n_2769),
.B(n_2796),
.Y(n_2868)
);

INVx2_ASAP7_75t_L g2869 ( 
.A(n_2706),
.Y(n_2869)
);

NAND2xp5_ASAP7_75t_SL g2870 ( 
.A(n_2705),
.B(n_2084),
.Y(n_2870)
);

OAI21xp5_ASAP7_75t_L g2871 ( 
.A1(n_2793),
.A2(n_2135),
.B(n_2218),
.Y(n_2871)
);

NAND2xp5_ASAP7_75t_L g2872 ( 
.A(n_2768),
.B(n_2442),
.Y(n_2872)
);

NAND2xp5_ASAP7_75t_L g2873 ( 
.A(n_2681),
.B(n_2442),
.Y(n_2873)
);

OAI22xp5_ASAP7_75t_L g2874 ( 
.A1(n_2663),
.A2(n_2485),
.B1(n_2573),
.B2(n_2559),
.Y(n_2874)
);

NOR2xp33_ASAP7_75t_L g2875 ( 
.A(n_2682),
.B(n_2084),
.Y(n_2875)
);

BUFx8_ASAP7_75t_L g2876 ( 
.A(n_2805),
.Y(n_2876)
);

OAI22x1_ASAP7_75t_L g2877 ( 
.A1(n_2659),
.A2(n_2559),
.B1(n_2645),
.B2(n_2573),
.Y(n_2877)
);

OAI22xp5_ASAP7_75t_L g2878 ( 
.A1(n_2663),
.A2(n_2645),
.B1(n_2238),
.B2(n_2040),
.Y(n_2878)
);

INVx3_ASAP7_75t_L g2879 ( 
.A(n_2728),
.Y(n_2879)
);

AOI21xp5_ASAP7_75t_L g2880 ( 
.A1(n_2785),
.A2(n_2443),
.B(n_2423),
.Y(n_2880)
);

NAND2xp5_ASAP7_75t_L g2881 ( 
.A(n_2766),
.B(n_2476),
.Y(n_2881)
);

INVx4_ASAP7_75t_L g2882 ( 
.A(n_2735),
.Y(n_2882)
);

OR2x2_ASAP7_75t_L g2883 ( 
.A(n_2809),
.B(n_2698),
.Y(n_2883)
);

AND2x2_ASAP7_75t_L g2884 ( 
.A(n_2687),
.B(n_2745),
.Y(n_2884)
);

AOI22x1_ASAP7_75t_L g2885 ( 
.A1(n_2716),
.A2(n_2811),
.B1(n_2751),
.B2(n_2764),
.Y(n_2885)
);

NAND2xp5_ASAP7_75t_L g2886 ( 
.A(n_2742),
.B(n_2700),
.Y(n_2886)
);

NAND2xp5_ASAP7_75t_L g2887 ( 
.A(n_2790),
.B(n_2476),
.Y(n_2887)
);

NAND3xp33_ASAP7_75t_L g2888 ( 
.A(n_2683),
.B(n_1602),
.C(n_1597),
.Y(n_2888)
);

NAND2xp5_ASAP7_75t_L g2889 ( 
.A(n_2790),
.B(n_2286),
.Y(n_2889)
);

A2O1A1Ixp33_ASAP7_75t_L g2890 ( 
.A1(n_2671),
.A2(n_2187),
.B(n_2184),
.C(n_1607),
.Y(n_2890)
);

NAND2xp5_ASAP7_75t_L g2891 ( 
.A(n_2813),
.B(n_2288),
.Y(n_2891)
);

INVx3_ASAP7_75t_L g2892 ( 
.A(n_2740),
.Y(n_2892)
);

INVx1_ASAP7_75t_L g2893 ( 
.A(n_2761),
.Y(n_2893)
);

AOI21xp5_ASAP7_75t_L g2894 ( 
.A1(n_2720),
.A2(n_2233),
.B(n_2154),
.Y(n_2894)
);

AOI21xp5_ASAP7_75t_L g2895 ( 
.A1(n_2721),
.A2(n_2233),
.B(n_2111),
.Y(n_2895)
);

AOI21xp5_ASAP7_75t_L g2896 ( 
.A1(n_2721),
.A2(n_2755),
.B(n_2799),
.Y(n_2896)
);

INVx4_ASAP7_75t_L g2897 ( 
.A(n_2735),
.Y(n_2897)
);

NOR2xp33_ASAP7_75t_L g2898 ( 
.A(n_2748),
.B(n_2161),
.Y(n_2898)
);

O2A1O1Ixp33_ASAP7_75t_L g2899 ( 
.A1(n_2718),
.A2(n_1615),
.B(n_1629),
.C(n_1597),
.Y(n_2899)
);

OA21x2_ASAP7_75t_L g2900 ( 
.A1(n_2718),
.A2(n_1584),
.B(n_1491),
.Y(n_2900)
);

NOR2xp67_ASAP7_75t_L g2901 ( 
.A(n_2662),
.B(n_2290),
.Y(n_2901)
);

AOI21xp5_ASAP7_75t_L g2902 ( 
.A1(n_2816),
.A2(n_2477),
.B(n_2436),
.Y(n_2902)
);

OAI22xp5_ASAP7_75t_L g2903 ( 
.A1(n_2683),
.A2(n_2464),
.B1(n_2333),
.B2(n_2095),
.Y(n_2903)
);

O2A1O1Ixp33_ASAP7_75t_L g2904 ( 
.A1(n_2715),
.A2(n_1629),
.B(n_1635),
.C(n_1615),
.Y(n_2904)
);

BUFx6f_ASAP7_75t_L g2905 ( 
.A(n_2792),
.Y(n_2905)
);

NAND2xp5_ASAP7_75t_SL g2906 ( 
.A(n_2656),
.B(n_2161),
.Y(n_2906)
);

NAND2xp5_ASAP7_75t_L g2907 ( 
.A(n_2813),
.B(n_2298),
.Y(n_2907)
);

AND2x4_ASAP7_75t_L g2908 ( 
.A(n_2665),
.B(n_2355),
.Y(n_2908)
);

OAI22xp5_ASAP7_75t_L g2909 ( 
.A1(n_2686),
.A2(n_2068),
.B1(n_2305),
.B2(n_2303),
.Y(n_2909)
);

INVx2_ASAP7_75t_L g2910 ( 
.A(n_2717),
.Y(n_2910)
);

NAND2x1p5_ASAP7_75t_L g2911 ( 
.A(n_2787),
.B(n_2479),
.Y(n_2911)
);

AOI21xp5_ASAP7_75t_L g2912 ( 
.A1(n_2656),
.A2(n_2436),
.B(n_2101),
.Y(n_2912)
);

NAND3xp33_ASAP7_75t_L g2913 ( 
.A(n_2760),
.B(n_1637),
.C(n_1635),
.Y(n_2913)
);

AOI21xp5_ASAP7_75t_L g2914 ( 
.A1(n_2667),
.A2(n_2479),
.B(n_2353),
.Y(n_2914)
);

AOI21xp5_ASAP7_75t_L g2915 ( 
.A1(n_2667),
.A2(n_2353),
.B(n_1943),
.Y(n_2915)
);

INVx2_ASAP7_75t_L g2916 ( 
.A(n_2675),
.Y(n_2916)
);

NAND2x1p5_ASAP7_75t_L g2917 ( 
.A(n_2787),
.B(n_2483),
.Y(n_2917)
);

INVx1_ASAP7_75t_L g2918 ( 
.A(n_2674),
.Y(n_2918)
);

A2O1A1Ixp33_ASAP7_75t_L g2919 ( 
.A1(n_2747),
.A2(n_1639),
.B(n_1637),
.C(n_2220),
.Y(n_2919)
);

NAND2xp5_ASAP7_75t_L g2920 ( 
.A(n_2815),
.B(n_2313),
.Y(n_2920)
);

AOI21xp5_ASAP7_75t_L g2921 ( 
.A1(n_2697),
.A2(n_2282),
.B(n_2280),
.Y(n_2921)
);

AOI22xp5_ASAP7_75t_L g2922 ( 
.A1(n_2665),
.A2(n_1631),
.B1(n_1522),
.B2(n_1531),
.Y(n_2922)
);

INVx1_ASAP7_75t_L g2923 ( 
.A(n_2678),
.Y(n_2923)
);

NAND2x1p5_ASAP7_75t_L g2924 ( 
.A(n_2787),
.B(n_2390),
.Y(n_2924)
);

BUFx6f_ASAP7_75t_L g2925 ( 
.A(n_2792),
.Y(n_2925)
);

AND2x2_ASAP7_75t_L g2926 ( 
.A(n_2740),
.B(n_2462),
.Y(n_2926)
);

INVx2_ASAP7_75t_L g2927 ( 
.A(n_2676),
.Y(n_2927)
);

INVx3_ASAP7_75t_L g2928 ( 
.A(n_2752),
.Y(n_2928)
);

NOR2xp33_ASAP7_75t_L g2929 ( 
.A(n_2756),
.B(n_2161),
.Y(n_2929)
);

INVx1_ASAP7_75t_L g2930 ( 
.A(n_2679),
.Y(n_2930)
);

NAND2xp5_ASAP7_75t_L g2931 ( 
.A(n_2815),
.B(n_2314),
.Y(n_2931)
);

OAI21xp33_ASAP7_75t_L g2932 ( 
.A1(n_2760),
.A2(n_1578),
.B(n_1526),
.Y(n_2932)
);

AOI21xp5_ASAP7_75t_L g2933 ( 
.A1(n_2697),
.A2(n_2282),
.B(n_2280),
.Y(n_2933)
);

A2O1A1Ixp33_ASAP7_75t_L g2934 ( 
.A1(n_2747),
.A2(n_1639),
.B(n_2227),
.C(n_2220),
.Y(n_2934)
);

NAND2xp5_ASAP7_75t_L g2935 ( 
.A(n_2794),
.B(n_2318),
.Y(n_2935)
);

OAI22xp5_ASAP7_75t_L g2936 ( 
.A1(n_2821),
.A2(n_2330),
.B1(n_2331),
.B2(n_2319),
.Y(n_2936)
);

INVx3_ASAP7_75t_L g2937 ( 
.A(n_2752),
.Y(n_2937)
);

AOI21xp5_ASAP7_75t_L g2938 ( 
.A1(n_2699),
.A2(n_2282),
.B(n_2280),
.Y(n_2938)
);

O2A1O1Ixp33_ASAP7_75t_L g2939 ( 
.A1(n_2804),
.A2(n_1507),
.B(n_1508),
.C(n_1501),
.Y(n_2939)
);

AND2x2_ASAP7_75t_L g2940 ( 
.A(n_2775),
.B(n_2468),
.Y(n_2940)
);

NOR2xp33_ASAP7_75t_L g2941 ( 
.A(n_2725),
.B(n_1526),
.Y(n_2941)
);

OAI22xp5_ASAP7_75t_L g2942 ( 
.A1(n_2692),
.A2(n_2347),
.B1(n_2350),
.B2(n_2344),
.Y(n_2942)
);

OR2x6_ASAP7_75t_SL g2943 ( 
.A(n_2722),
.B(n_2474),
.Y(n_2943)
);

BUFx3_ASAP7_75t_L g2944 ( 
.A(n_2749),
.Y(n_2944)
);

INVx2_ASAP7_75t_L g2945 ( 
.A(n_2689),
.Y(n_2945)
);

NAND2xp5_ASAP7_75t_L g2946 ( 
.A(n_2810),
.B(n_2368),
.Y(n_2946)
);

OAI22xp5_ASAP7_75t_L g2947 ( 
.A1(n_2802),
.A2(n_2375),
.B1(n_2379),
.B2(n_2372),
.Y(n_2947)
);

INVxp67_ASAP7_75t_L g2948 ( 
.A(n_2780),
.Y(n_2948)
);

INVx2_ASAP7_75t_L g2949 ( 
.A(n_2690),
.Y(n_2949)
);

INVx2_ASAP7_75t_L g2950 ( 
.A(n_2657),
.Y(n_2950)
);

HB1xp67_ASAP7_75t_L g2951 ( 
.A(n_2772),
.Y(n_2951)
);

AOI21xp5_ASAP7_75t_L g2952 ( 
.A1(n_2699),
.A2(n_2311),
.B(n_2293),
.Y(n_2952)
);

NAND2xp5_ASAP7_75t_SL g2953 ( 
.A(n_2713),
.B(n_2376),
.Y(n_2953)
);

INVx1_ASAP7_75t_L g2954 ( 
.A(n_2688),
.Y(n_2954)
);

NAND2xp5_ASAP7_75t_L g2955 ( 
.A(n_2810),
.B(n_2376),
.Y(n_2955)
);

NAND2xp5_ASAP7_75t_L g2956 ( 
.A(n_2743),
.B(n_2405),
.Y(n_2956)
);

NOR2x1_ASAP7_75t_L g2957 ( 
.A(n_2774),
.B(n_2390),
.Y(n_2957)
);

OAI22x1_ASAP7_75t_L g2958 ( 
.A1(n_2660),
.A2(n_2414),
.B1(n_2450),
.B2(n_2415),
.Y(n_2958)
);

AND2x2_ASAP7_75t_L g2959 ( 
.A(n_2775),
.B(n_2355),
.Y(n_2959)
);

O2A1O1Ixp5_ASAP7_75t_L g2960 ( 
.A1(n_2670),
.A2(n_2234),
.B(n_2480),
.C(n_2030),
.Y(n_2960)
);

NOR2xp33_ASAP7_75t_L g2961 ( 
.A(n_2668),
.B(n_1578),
.Y(n_2961)
);

AO32x1_ASAP7_75t_L g2962 ( 
.A1(n_2779),
.A2(n_2786),
.A3(n_2784),
.B1(n_2808),
.B2(n_2759),
.Y(n_2962)
);

NAND2xp5_ASAP7_75t_SL g2963 ( 
.A(n_2713),
.B(n_2757),
.Y(n_2963)
);

INVx3_ASAP7_75t_L g2964 ( 
.A(n_2723),
.Y(n_2964)
);

NAND2xp5_ASAP7_75t_SL g2965 ( 
.A(n_2757),
.B(n_2293),
.Y(n_2965)
);

O2A1O1Ixp33_ASAP7_75t_L g2966 ( 
.A1(n_2746),
.A2(n_2661),
.B(n_2776),
.C(n_2767),
.Y(n_2966)
);

OAI22xp5_ASAP7_75t_L g2967 ( 
.A1(n_2802),
.A2(n_2030),
.B1(n_2059),
.B2(n_2134),
.Y(n_2967)
);

NOR2xp33_ASAP7_75t_L g2968 ( 
.A(n_2680),
.B(n_1512),
.Y(n_2968)
);

OAI22xp5_ASAP7_75t_L g2969 ( 
.A1(n_2806),
.A2(n_2059),
.B1(n_2137),
.B2(n_2134),
.Y(n_2969)
);

HB1xp67_ASAP7_75t_L g2970 ( 
.A(n_2763),
.Y(n_2970)
);

INVx4_ASAP7_75t_L g2971 ( 
.A(n_2801),
.Y(n_2971)
);

AND2x2_ASAP7_75t_L g2972 ( 
.A(n_2819),
.B(n_2181),
.Y(n_2972)
);

A2O1A1Ixp33_ASAP7_75t_SL g2973 ( 
.A1(n_2719),
.A2(n_1518),
.B(n_1519),
.C(n_1512),
.Y(n_2973)
);

CKINVDCx5p33_ASAP7_75t_R g2974 ( 
.A(n_2749),
.Y(n_2974)
);

NAND2xp5_ASAP7_75t_L g2975 ( 
.A(n_2731),
.B(n_1503),
.Y(n_2975)
);

NAND2xp5_ASAP7_75t_SL g2976 ( 
.A(n_2664),
.B(n_2311),
.Y(n_2976)
);

INVx1_ASAP7_75t_L g2977 ( 
.A(n_2707),
.Y(n_2977)
);

OAI22xp5_ASAP7_75t_L g2978 ( 
.A1(n_2702),
.A2(n_2139),
.B1(n_2145),
.B2(n_2137),
.Y(n_2978)
);

BUFx8_ASAP7_75t_L g2979 ( 
.A(n_2805),
.Y(n_2979)
);

O2A1O1Ixp33_ASAP7_75t_L g2980 ( 
.A1(n_2709),
.A2(n_1488),
.B(n_1493),
.C(n_1486),
.Y(n_2980)
);

AO32x1_ASAP7_75t_L g2981 ( 
.A1(n_2737),
.A2(n_2145),
.A3(n_2150),
.B1(n_2149),
.B2(n_2139),
.Y(n_2981)
);

AO21x1_ASAP7_75t_L g2982 ( 
.A1(n_2966),
.A2(n_2727),
.B(n_2738),
.Y(n_2982)
);

AO31x2_ASAP7_75t_L g2983 ( 
.A1(n_2877),
.A2(n_2673),
.A3(n_2694),
.B(n_2657),
.Y(n_2983)
);

OAI22xp5_ASAP7_75t_L g2984 ( 
.A1(n_2855),
.A2(n_2819),
.B1(n_2694),
.B2(n_2696),
.Y(n_2984)
);

BUFx6f_ASAP7_75t_L g2985 ( 
.A(n_2825),
.Y(n_2985)
);

AOI221x1_ASAP7_75t_L g2986 ( 
.A1(n_2827),
.A2(n_2818),
.B1(n_2791),
.B2(n_2729),
.C(n_2744),
.Y(n_2986)
);

AND2x2_ASAP7_75t_L g2987 ( 
.A(n_2884),
.B(n_2669),
.Y(n_2987)
);

OR2x2_ASAP7_75t_L g2988 ( 
.A(n_2883),
.B(n_2703),
.Y(n_2988)
);

NAND2xp5_ASAP7_75t_L g2989 ( 
.A(n_2886),
.B(n_2714),
.Y(n_2989)
);

NOR2xp33_ASAP7_75t_L g2990 ( 
.A(n_2866),
.B(n_2664),
.Y(n_2990)
);

OAI21x1_ASAP7_75t_L g2991 ( 
.A1(n_2894),
.A2(n_2895),
.B(n_2824),
.Y(n_2991)
);

CKINVDCx8_ASAP7_75t_R g2992 ( 
.A(n_2974),
.Y(n_2992)
);

INVx2_ASAP7_75t_L g2993 ( 
.A(n_2869),
.Y(n_2993)
);

INVx1_ASAP7_75t_L g2994 ( 
.A(n_2918),
.Y(n_2994)
);

INVx2_ASAP7_75t_SL g2995 ( 
.A(n_2876),
.Y(n_2995)
);

NAND2xp5_ASAP7_75t_L g2996 ( 
.A(n_2853),
.B(n_2714),
.Y(n_2996)
);

AOI21xp5_ASAP7_75t_L g2997 ( 
.A1(n_2831),
.A2(n_2817),
.B(n_2730),
.Y(n_2997)
);

OAI21x1_ASAP7_75t_L g2998 ( 
.A1(n_2914),
.A2(n_2818),
.B(n_2791),
.Y(n_2998)
);

OAI21x1_ASAP7_75t_L g2999 ( 
.A1(n_2915),
.A2(n_2162),
.B(n_2136),
.Y(n_2999)
);

NOR2xp33_ASAP7_75t_L g3000 ( 
.A(n_2862),
.B(n_2672),
.Y(n_3000)
);

NAND2xp5_ASAP7_75t_SL g3001 ( 
.A(n_2885),
.B(n_2723),
.Y(n_3001)
);

NAND2xp5_ASAP7_75t_L g3002 ( 
.A(n_2838),
.B(n_2714),
.Y(n_3002)
);

OAI21x1_ASAP7_75t_L g3003 ( 
.A1(n_2880),
.A2(n_2162),
.B(n_2136),
.Y(n_3003)
);

AO21x2_ASAP7_75t_L g3004 ( 
.A1(n_2864),
.A2(n_1950),
.B(n_2198),
.Y(n_3004)
);

OAI21x1_ASAP7_75t_L g3005 ( 
.A1(n_2902),
.A2(n_2849),
.B(n_2842),
.Y(n_3005)
);

OAI21x1_ASAP7_75t_L g3006 ( 
.A1(n_2857),
.A2(n_2162),
.B(n_2136),
.Y(n_3006)
);

AOI22xp5_ASAP7_75t_L g3007 ( 
.A1(n_2906),
.A2(n_2714),
.B1(n_2449),
.B2(n_2132),
.Y(n_3007)
);

INVx5_ASAP7_75t_L g3008 ( 
.A(n_2829),
.Y(n_3008)
);

INVx1_ASAP7_75t_SL g3009 ( 
.A(n_2840),
.Y(n_3009)
);

AOI21xp5_ASAP7_75t_L g3010 ( 
.A1(n_2847),
.A2(n_2329),
.B(n_2326),
.Y(n_3010)
);

OAI21xp5_ASAP7_75t_L g3011 ( 
.A1(n_2823),
.A2(n_2913),
.B(n_2960),
.Y(n_3011)
);

AO31x2_ASAP7_75t_L g3012 ( 
.A1(n_2958),
.A2(n_2765),
.A3(n_2797),
.B(n_2708),
.Y(n_3012)
);

NAND2xp5_ASAP7_75t_L g3013 ( 
.A(n_2851),
.B(n_2852),
.Y(n_3013)
);

OAI21xp5_ASAP7_75t_L g3014 ( 
.A1(n_2890),
.A2(n_2132),
.B(n_2179),
.Y(n_3014)
);

CKINVDCx11_ASAP7_75t_R g3015 ( 
.A(n_2839),
.Y(n_3015)
);

NAND2xp33_ASAP7_75t_L g3016 ( 
.A(n_2828),
.B(n_2932),
.Y(n_3016)
);

NAND2xp5_ASAP7_75t_L g3017 ( 
.A(n_2970),
.B(n_2723),
.Y(n_3017)
);

OAI21x1_ASAP7_75t_L g3018 ( 
.A1(n_2832),
.A2(n_2169),
.B(n_2165),
.Y(n_3018)
);

INVx1_ASAP7_75t_L g3019 ( 
.A(n_2923),
.Y(n_3019)
);

OAI21x1_ASAP7_75t_L g3020 ( 
.A1(n_2837),
.A2(n_2182),
.B(n_2170),
.Y(n_3020)
);

OAI21xp5_ASAP7_75t_L g3021 ( 
.A1(n_2904),
.A2(n_2888),
.B(n_2871),
.Y(n_3021)
);

OAI21xp5_ASAP7_75t_L g3022 ( 
.A1(n_2896),
.A2(n_2934),
.B(n_2848),
.Y(n_3022)
);

OAI21x1_ASAP7_75t_L g3023 ( 
.A1(n_2912),
.A2(n_2182),
.B(n_2170),
.Y(n_3023)
);

BUFx3_ASAP7_75t_L g3024 ( 
.A(n_2876),
.Y(n_3024)
);

AO31x2_ASAP7_75t_L g3025 ( 
.A1(n_2942),
.A2(n_2797),
.A3(n_2090),
.B(n_2094),
.Y(n_3025)
);

INVx4_ASAP7_75t_L g3026 ( 
.A(n_2829),
.Y(n_3026)
);

NAND2xp5_ASAP7_75t_L g3027 ( 
.A(n_2843),
.B(n_2724),
.Y(n_3027)
);

NAND2xp5_ASAP7_75t_L g3028 ( 
.A(n_2868),
.B(n_2724),
.Y(n_3028)
);

A2O1A1Ixp33_ASAP7_75t_L g3029 ( 
.A1(n_2961),
.A2(n_2704),
.B(n_2762),
.C(n_2691),
.Y(n_3029)
);

INVx2_ASAP7_75t_L g3030 ( 
.A(n_2910),
.Y(n_3030)
);

INVx2_ASAP7_75t_L g3031 ( 
.A(n_2863),
.Y(n_3031)
);

INVx4_ASAP7_75t_L g3032 ( 
.A(n_2882),
.Y(n_3032)
);

OAI21x1_ASAP7_75t_L g3033 ( 
.A1(n_2921),
.A2(n_2193),
.B(n_2185),
.Y(n_3033)
);

AND2x2_ASAP7_75t_L g3034 ( 
.A(n_2943),
.B(n_2850),
.Y(n_3034)
);

OAI22xp5_ASAP7_75t_L g3035 ( 
.A1(n_2855),
.A2(n_2712),
.B1(n_2704),
.B2(n_2691),
.Y(n_3035)
);

OAI21x1_ASAP7_75t_L g3036 ( 
.A1(n_2933),
.A2(n_2193),
.B(n_2185),
.Y(n_3036)
);

OAI21x1_ASAP7_75t_L g3037 ( 
.A1(n_2938),
.A2(n_2097),
.B(n_2096),
.Y(n_3037)
);

A2O1A1Ixp33_ASAP7_75t_L g3038 ( 
.A1(n_2835),
.A2(n_2798),
.B(n_2807),
.C(n_2762),
.Y(n_3038)
);

NAND2xp5_ASAP7_75t_L g3039 ( 
.A(n_2845),
.B(n_2724),
.Y(n_3039)
);

INVx2_ASAP7_75t_L g3040 ( 
.A(n_2867),
.Y(n_3040)
);

AND2x4_ASAP7_75t_L g3041 ( 
.A(n_2833),
.B(n_2798),
.Y(n_3041)
);

NAND2xp5_ASAP7_75t_SL g3042 ( 
.A(n_2856),
.B(n_2834),
.Y(n_3042)
);

INVx1_ASAP7_75t_L g3043 ( 
.A(n_2930),
.Y(n_3043)
);

OAI21x1_ASAP7_75t_L g3044 ( 
.A1(n_2952),
.A2(n_2105),
.B(n_2097),
.Y(n_3044)
);

A2O1A1Ixp33_ASAP7_75t_L g3045 ( 
.A1(n_2939),
.A2(n_2807),
.B(n_2729),
.C(n_2744),
.Y(n_3045)
);

AO31x2_ASAP7_75t_L g3046 ( 
.A1(n_2947),
.A2(n_2874),
.A3(n_2969),
.B(n_2919),
.Y(n_3046)
);

NAND2x1p5_ASAP7_75t_L g3047 ( 
.A(n_2836),
.B(n_2724),
.Y(n_3047)
);

AOI211x1_ASAP7_75t_L g3048 ( 
.A1(n_2830),
.A2(n_69),
.B(n_67),
.C(n_68),
.Y(n_3048)
);

INVx1_ASAP7_75t_L g3049 ( 
.A(n_2954),
.Y(n_3049)
);

OAI21xp5_ASAP7_75t_SL g3050 ( 
.A1(n_2941),
.A2(n_2744),
.B(n_2729),
.Y(n_3050)
);

OAI21xp5_ASAP7_75t_L g3051 ( 
.A1(n_2909),
.A2(n_2936),
.B(n_2878),
.Y(n_3051)
);

A2O1A1Ixp33_ASAP7_75t_L g3052 ( 
.A1(n_2968),
.A2(n_2744),
.B(n_2781),
.C(n_2729),
.Y(n_3052)
);

AOI21xp33_ASAP7_75t_L g3053 ( 
.A1(n_2844),
.A2(n_2873),
.B(n_2973),
.Y(n_3053)
);

AO31x2_ASAP7_75t_L g3054 ( 
.A1(n_2967),
.A2(n_2112),
.A3(n_2089),
.B(n_2186),
.Y(n_3054)
);

OAI21xp5_ASAP7_75t_L g3055 ( 
.A1(n_2899),
.A2(n_2179),
.B(n_2449),
.Y(n_3055)
);

AO31x2_ASAP7_75t_L g3056 ( 
.A1(n_2977),
.A2(n_2192),
.A3(n_2197),
.B(n_2186),
.Y(n_3056)
);

OAI22xp5_ASAP7_75t_L g3057 ( 
.A1(n_2948),
.A2(n_2781),
.B1(n_2105),
.B2(n_2124),
.Y(n_3057)
);

A2O1A1Ixp33_ASAP7_75t_L g3058 ( 
.A1(n_2903),
.A2(n_2781),
.B(n_1522),
.C(n_1531),
.Y(n_3058)
);

INVx4_ASAP7_75t_L g3059 ( 
.A(n_2882),
.Y(n_3059)
);

OAI21x1_ASAP7_75t_L g3060 ( 
.A1(n_2957),
.A2(n_2124),
.B(n_2028),
.Y(n_3060)
);

AO31x2_ASAP7_75t_L g3061 ( 
.A1(n_2978),
.A2(n_2197),
.A3(n_2192),
.B(n_2150),
.Y(n_3061)
);

NAND2xp5_ASAP7_75t_L g3062 ( 
.A(n_2893),
.B(n_2946),
.Y(n_3062)
);

OAI21xp5_ASAP7_75t_L g3063 ( 
.A1(n_2854),
.A2(n_2179),
.B(n_2153),
.Y(n_3063)
);

NAND2xp5_ASAP7_75t_SL g3064 ( 
.A(n_2875),
.B(n_1594),
.Y(n_3064)
);

NAND2xp5_ASAP7_75t_L g3065 ( 
.A(n_2955),
.B(n_2950),
.Y(n_3065)
);

OAI21xp5_ASAP7_75t_L g3066 ( 
.A1(n_2870),
.A2(n_2179),
.B(n_2157),
.Y(n_3066)
);

AOI21x1_ASAP7_75t_L g3067 ( 
.A1(n_2901),
.A2(n_1500),
.B(n_1496),
.Y(n_3067)
);

OAI22xp5_ASAP7_75t_L g3068 ( 
.A1(n_2965),
.A2(n_2160),
.B1(n_2163),
.B2(n_2144),
.Y(n_3068)
);

NAND2xp5_ASAP7_75t_SL g3069 ( 
.A(n_2836),
.B(n_1594),
.Y(n_3069)
);

INVx1_ASAP7_75t_L g3070 ( 
.A(n_2916),
.Y(n_3070)
);

NAND2xp5_ASAP7_75t_SL g3071 ( 
.A(n_2836),
.B(n_2898),
.Y(n_3071)
);

OAI21xp5_ASAP7_75t_L g3072 ( 
.A1(n_2980),
.A2(n_1500),
.B(n_2201),
.Y(n_3072)
);

NAND2xp5_ASAP7_75t_L g3073 ( 
.A(n_2927),
.B(n_1503),
.Y(n_3073)
);

NAND2xp5_ASAP7_75t_L g3074 ( 
.A(n_2945),
.B(n_1522),
.Y(n_3074)
);

OAI21x1_ASAP7_75t_L g3075 ( 
.A1(n_2900),
.A2(n_2163),
.B(n_2144),
.Y(n_3075)
);

INVx1_ASAP7_75t_L g3076 ( 
.A(n_2949),
.Y(n_3076)
);

OAI21xp5_ASAP7_75t_L g3077 ( 
.A1(n_2975),
.A2(n_2953),
.B(n_2872),
.Y(n_3077)
);

INVx1_ASAP7_75t_L g3078 ( 
.A(n_2962),
.Y(n_3078)
);

OAI21xp5_ASAP7_75t_L g3079 ( 
.A1(n_2881),
.A2(n_2935),
.B(n_2891),
.Y(n_3079)
);

OAI21xp5_ASAP7_75t_L g3080 ( 
.A1(n_2889),
.A2(n_2178),
.B(n_1595),
.Y(n_3080)
);

INVx1_ASAP7_75t_L g3081 ( 
.A(n_2962),
.Y(n_3081)
);

OA21x2_ASAP7_75t_L g3082 ( 
.A1(n_2963),
.A2(n_2178),
.B(n_1502),
.Y(n_3082)
);

INVx1_ASAP7_75t_L g3083 ( 
.A(n_2962),
.Y(n_3083)
);

AO21x1_ASAP7_75t_L g3084 ( 
.A1(n_2976),
.A2(n_1595),
.B(n_1531),
.Y(n_3084)
);

OAI21x1_ASAP7_75t_L g3085 ( 
.A1(n_2907),
.A2(n_2931),
.B(n_2920),
.Y(n_3085)
);

OAI21xp33_ASAP7_75t_L g3086 ( 
.A1(n_2826),
.A2(n_1595),
.B(n_1531),
.Y(n_3086)
);

INVx2_ASAP7_75t_SL g3087 ( 
.A(n_2979),
.Y(n_3087)
);

OAI21x1_ASAP7_75t_L g3088 ( 
.A1(n_2887),
.A2(n_1502),
.B(n_1481),
.Y(n_3088)
);

BUFx6f_ASAP7_75t_L g3089 ( 
.A(n_2825),
.Y(n_3089)
);

AO31x2_ASAP7_75t_L g3090 ( 
.A1(n_2897),
.A2(n_1525),
.A3(n_1530),
.B(n_1510),
.Y(n_3090)
);

OAI21x1_ASAP7_75t_L g3091 ( 
.A1(n_2956),
.A2(n_1525),
.B(n_1510),
.Y(n_3091)
);

BUFx6f_ASAP7_75t_SL g3092 ( 
.A(n_2860),
.Y(n_3092)
);

BUFx6f_ASAP7_75t_L g3093 ( 
.A(n_2825),
.Y(n_3093)
);

AOI22xp5_ASAP7_75t_L g3094 ( 
.A1(n_2841),
.A2(n_1604),
.B1(n_1485),
.B2(n_1476),
.Y(n_3094)
);

NAND2xp5_ASAP7_75t_L g3095 ( 
.A(n_2972),
.B(n_1604),
.Y(n_3095)
);

AOI21xp5_ASAP7_75t_L g3096 ( 
.A1(n_2859),
.A2(n_1617),
.B(n_1594),
.Y(n_3096)
);

NAND2xp5_ASAP7_75t_SL g3097 ( 
.A(n_2908),
.B(n_1617),
.Y(n_3097)
);

AOI22xp5_ASAP7_75t_L g3098 ( 
.A1(n_2922),
.A2(n_1604),
.B1(n_1485),
.B2(n_1476),
.Y(n_3098)
);

AOI21xp5_ASAP7_75t_L g3099 ( 
.A1(n_2859),
.A2(n_1617),
.B(n_1541),
.Y(n_3099)
);

BUFx6f_ASAP7_75t_L g3100 ( 
.A(n_2846),
.Y(n_3100)
);

AOI221xp5_ASAP7_75t_SL g3101 ( 
.A1(n_2926),
.A2(n_67),
.B1(n_68),
.B2(n_69),
.C(n_72),
.Y(n_3101)
);

NAND2xp5_ASAP7_75t_L g3102 ( 
.A(n_2940),
.B(n_72),
.Y(n_3102)
);

BUFx6f_ASAP7_75t_L g3103 ( 
.A(n_2846),
.Y(n_3103)
);

HB1xp67_ASAP7_75t_L g3104 ( 
.A(n_2865),
.Y(n_3104)
);

A2O1A1Ixp33_ASAP7_75t_L g3105 ( 
.A1(n_2858),
.A2(n_1485),
.B(n_1476),
.C(n_1550),
.Y(n_3105)
);

AOI21xp5_ASAP7_75t_L g3106 ( 
.A1(n_2859),
.A2(n_1552),
.B(n_1550),
.Y(n_3106)
);

AOI21xp5_ASAP7_75t_L g3107 ( 
.A1(n_2981),
.A2(n_1554),
.B(n_1552),
.Y(n_3107)
);

NAND2xp5_ASAP7_75t_L g3108 ( 
.A(n_2908),
.B(n_2879),
.Y(n_3108)
);

OAI21x1_ASAP7_75t_SL g3109 ( 
.A1(n_2897),
.A2(n_1634),
.B(n_1598),
.Y(n_3109)
);

NAND2xp5_ASAP7_75t_L g3110 ( 
.A(n_2879),
.B(n_2892),
.Y(n_3110)
);

AOI21xp5_ASAP7_75t_L g3111 ( 
.A1(n_2981),
.A2(n_1559),
.B(n_1554),
.Y(n_3111)
);

OAI21xp33_ASAP7_75t_L g3112 ( 
.A1(n_2929),
.A2(n_1562),
.B(n_1559),
.Y(n_3112)
);

AOI21xp5_ASAP7_75t_L g3113 ( 
.A1(n_2981),
.A2(n_1565),
.B(n_1562),
.Y(n_3113)
);

HB1xp67_ASAP7_75t_L g3114 ( 
.A(n_2964),
.Y(n_3114)
);

NOR2xp67_ASAP7_75t_L g3115 ( 
.A(n_2892),
.B(n_76),
.Y(n_3115)
);

INVx2_ASAP7_75t_L g3116 ( 
.A(n_2928),
.Y(n_3116)
);

OAI21x1_ASAP7_75t_L g3117 ( 
.A1(n_2911),
.A2(n_1567),
.B(n_1565),
.Y(n_3117)
);

OAI21x1_ASAP7_75t_L g3118 ( 
.A1(n_2917),
.A2(n_1582),
.B(n_1567),
.Y(n_3118)
);

AO21x2_ASAP7_75t_L g3119 ( 
.A1(n_2861),
.A2(n_1582),
.B(n_1641),
.Y(n_3119)
);

OAI21x1_ASAP7_75t_L g3120 ( 
.A1(n_2924),
.A2(n_1634),
.B(n_1598),
.Y(n_3120)
);

OAI21x1_ASAP7_75t_L g3121 ( 
.A1(n_2937),
.A2(n_2959),
.B(n_2861),
.Y(n_3121)
);

A2O1A1Ixp33_ASAP7_75t_L g3122 ( 
.A1(n_2858),
.A2(n_84),
.B(n_78),
.C(n_80),
.Y(n_3122)
);

OAI21x1_ASAP7_75t_L g3123 ( 
.A1(n_2971),
.A2(n_1580),
.B(n_1579),
.Y(n_3123)
);

NAND2xp5_ASAP7_75t_L g3124 ( 
.A(n_2846),
.B(n_78),
.Y(n_3124)
);

AO31x2_ASAP7_75t_L g3125 ( 
.A1(n_2905),
.A2(n_1644),
.A3(n_1651),
.B(n_1642),
.Y(n_3125)
);

OAI21xp5_ASAP7_75t_L g3126 ( 
.A1(n_2944),
.A2(n_1580),
.B(n_1579),
.Y(n_3126)
);

INVx1_ASAP7_75t_L g3127 ( 
.A(n_2979),
.Y(n_3127)
);

AO31x2_ASAP7_75t_L g3128 ( 
.A1(n_2905),
.A2(n_1651),
.A3(n_1580),
.B(n_1579),
.Y(n_3128)
);

NAND2xp5_ASAP7_75t_L g3129 ( 
.A(n_2905),
.B(n_1580),
.Y(n_3129)
);

AND2x4_ASAP7_75t_L g3130 ( 
.A(n_2925),
.B(n_362),
.Y(n_3130)
);

NAND3xp33_ASAP7_75t_SL g3131 ( 
.A(n_2925),
.B(n_84),
.C(n_85),
.Y(n_3131)
);

INVx2_ASAP7_75t_L g3132 ( 
.A(n_2925),
.Y(n_3132)
);

INVx6_ASAP7_75t_L g3133 ( 
.A(n_2876),
.Y(n_3133)
);

OAI21x1_ASAP7_75t_L g3134 ( 
.A1(n_2822),
.A2(n_1579),
.B(n_1462),
.Y(n_3134)
);

AND2x2_ASAP7_75t_L g3135 ( 
.A(n_2884),
.B(n_86),
.Y(n_3135)
);

INVx1_ASAP7_75t_L g3136 ( 
.A(n_2951),
.Y(n_3136)
);

OAI21x1_ASAP7_75t_L g3137 ( 
.A1(n_2822),
.A2(n_1462),
.B(n_1451),
.Y(n_3137)
);

NAND3xp33_ASAP7_75t_SL g3138 ( 
.A(n_2966),
.B(n_86),
.C(n_87),
.Y(n_3138)
);

AOI221x1_ASAP7_75t_L g3139 ( 
.A1(n_2827),
.A2(n_88),
.B1(n_90),
.B2(n_91),
.C(n_93),
.Y(n_3139)
);

OAI21xp5_ASAP7_75t_L g3140 ( 
.A1(n_2822),
.A2(n_1462),
.B(n_1451),
.Y(n_3140)
);

O2A1O1Ixp33_ASAP7_75t_L g3141 ( 
.A1(n_3122),
.A2(n_93),
.B(n_88),
.C(n_91),
.Y(n_3141)
);

AOI21x1_ASAP7_75t_L g3142 ( 
.A1(n_3001),
.A2(n_1474),
.B(n_94),
.Y(n_3142)
);

INVx4_ASAP7_75t_L g3143 ( 
.A(n_3008),
.Y(n_3143)
);

OAI21xp5_ASAP7_75t_L g3144 ( 
.A1(n_3042),
.A2(n_98),
.B(n_99),
.Y(n_3144)
);

INVx1_ASAP7_75t_L g3145 ( 
.A(n_2994),
.Y(n_3145)
);

AND2x4_ASAP7_75t_L g3146 ( 
.A(n_3104),
.B(n_98),
.Y(n_3146)
);

OAI21x1_ASAP7_75t_SL g3147 ( 
.A1(n_2982),
.A2(n_99),
.B(n_102),
.Y(n_3147)
);

INVx3_ASAP7_75t_L g3148 ( 
.A(n_3041),
.Y(n_3148)
);

INVx1_ASAP7_75t_L g3149 ( 
.A(n_3019),
.Y(n_3149)
);

OAI21x1_ASAP7_75t_L g3150 ( 
.A1(n_3005),
.A2(n_2999),
.B(n_2991),
.Y(n_3150)
);

NAND2xp5_ASAP7_75t_L g3151 ( 
.A(n_3013),
.B(n_102),
.Y(n_3151)
);

OAI22xp33_ASAP7_75t_L g3152 ( 
.A1(n_3139),
.A2(n_1515),
.B1(n_1497),
.B2(n_1535),
.Y(n_3152)
);

NAND3xp33_ASAP7_75t_SL g3153 ( 
.A(n_3058),
.B(n_103),
.C(n_104),
.Y(n_3153)
);

INVx1_ASAP7_75t_L g3154 ( 
.A(n_3043),
.Y(n_3154)
);

OAI21xp5_ASAP7_75t_L g3155 ( 
.A1(n_3016),
.A2(n_103),
.B(n_104),
.Y(n_3155)
);

O2A1O1Ixp33_ASAP7_75t_L g3156 ( 
.A1(n_3138),
.A2(n_107),
.B(n_105),
.C(n_106),
.Y(n_3156)
);

NAND3x1_ASAP7_75t_L g3157 ( 
.A(n_3127),
.B(n_105),
.C(n_109),
.Y(n_3157)
);

NAND2xp5_ASAP7_75t_L g3158 ( 
.A(n_3034),
.B(n_110),
.Y(n_3158)
);

AND2x6_ASAP7_75t_SL g3159 ( 
.A(n_2990),
.B(n_110),
.Y(n_3159)
);

AOI221x1_ASAP7_75t_L g3160 ( 
.A1(n_3038),
.A2(n_111),
.B1(n_112),
.B2(n_114),
.C(n_115),
.Y(n_3160)
);

NAND2xp5_ASAP7_75t_SL g3161 ( 
.A(n_3029),
.B(n_1515),
.Y(n_3161)
);

O2A1O1Ixp5_ASAP7_75t_L g3162 ( 
.A1(n_3022),
.A2(n_111),
.B(n_112),
.C(n_116),
.Y(n_3162)
);

OA21x2_ASAP7_75t_L g3163 ( 
.A1(n_3078),
.A2(n_118),
.B(n_119),
.Y(n_3163)
);

OAI21xp5_ASAP7_75t_SL g3164 ( 
.A1(n_3131),
.A2(n_3051),
.B(n_3050),
.Y(n_3164)
);

AO221x2_ASAP7_75t_L g3165 ( 
.A1(n_3050),
.A2(n_118),
.B1(n_119),
.B2(n_120),
.C(n_121),
.Y(n_3165)
);

AOI21xp5_ASAP7_75t_L g3166 ( 
.A1(n_3014),
.A2(n_1515),
.B(n_1497),
.Y(n_3166)
);

INVx2_ASAP7_75t_L g3167 ( 
.A(n_3049),
.Y(n_3167)
);

AOI21xp5_ASAP7_75t_L g3168 ( 
.A1(n_3014),
.A2(n_1515),
.B(n_1497),
.Y(n_3168)
);

NAND2xp5_ASAP7_75t_L g3169 ( 
.A(n_3002),
.B(n_122),
.Y(n_3169)
);

BUFx6f_ASAP7_75t_L g3170 ( 
.A(n_3015),
.Y(n_3170)
);

AOI21xp5_ASAP7_75t_L g3171 ( 
.A1(n_3021),
.A2(n_1497),
.B(n_1535),
.Y(n_3171)
);

CKINVDCx20_ASAP7_75t_R g3172 ( 
.A(n_2992),
.Y(n_3172)
);

BUFx3_ASAP7_75t_L g3173 ( 
.A(n_3133),
.Y(n_3173)
);

OAI21xp5_ASAP7_75t_L g3174 ( 
.A1(n_3101),
.A2(n_3011),
.B(n_3045),
.Y(n_3174)
);

NAND2xp5_ASAP7_75t_L g3175 ( 
.A(n_2996),
.B(n_122),
.Y(n_3175)
);

O2A1O1Ixp33_ASAP7_75t_SL g3176 ( 
.A1(n_3052),
.A2(n_123),
.B(n_125),
.C(n_126),
.Y(n_3176)
);

CKINVDCx6p67_ASAP7_75t_R g3177 ( 
.A(n_3092),
.Y(n_3177)
);

NAND3xp33_ASAP7_75t_SL g3178 ( 
.A(n_3064),
.B(n_123),
.C(n_125),
.Y(n_3178)
);

INVx3_ASAP7_75t_L g3179 ( 
.A(n_3041),
.Y(n_3179)
);

INVx5_ASAP7_75t_L g3180 ( 
.A(n_3133),
.Y(n_3180)
);

AOI21x1_ASAP7_75t_L g3181 ( 
.A1(n_2997),
.A2(n_127),
.B(n_128),
.Y(n_3181)
);

AND2x2_ASAP7_75t_L g3182 ( 
.A(n_3009),
.B(n_128),
.Y(n_3182)
);

BUFx3_ASAP7_75t_L g3183 ( 
.A(n_3024),
.Y(n_3183)
);

O2A1O1Ixp33_ASAP7_75t_L g3184 ( 
.A1(n_3053),
.A2(n_129),
.B(n_130),
.C(n_131),
.Y(n_3184)
);

OA21x2_ASAP7_75t_L g3185 ( 
.A1(n_3081),
.A2(n_129),
.B(n_130),
.Y(n_3185)
);

OR2x6_ASAP7_75t_L g3186 ( 
.A(n_3010),
.B(n_3121),
.Y(n_3186)
);

OAI21xp5_ASAP7_75t_L g3187 ( 
.A1(n_3053),
.A2(n_132),
.B(n_133),
.Y(n_3187)
);

NOR2xp33_ASAP7_75t_SL g3188 ( 
.A(n_3026),
.B(n_3008),
.Y(n_3188)
);

NAND2xp5_ASAP7_75t_L g3189 ( 
.A(n_2989),
.B(n_135),
.Y(n_3189)
);

AOI21xp5_ASAP7_75t_L g3190 ( 
.A1(n_3055),
.A2(n_1551),
.B(n_1543),
.Y(n_3190)
);

AO31x2_ASAP7_75t_L g3191 ( 
.A1(n_2986),
.A2(n_135),
.A3(n_136),
.B(n_137),
.Y(n_3191)
);

A2O1A1Ixp33_ASAP7_75t_L g3192 ( 
.A1(n_3007),
.A2(n_137),
.B(n_139),
.C(n_140),
.Y(n_3192)
);

NAND2xp5_ASAP7_75t_L g3193 ( 
.A(n_3136),
.B(n_140),
.Y(n_3193)
);

AO31x2_ASAP7_75t_L g3194 ( 
.A1(n_3096),
.A2(n_141),
.A3(n_142),
.B(n_144),
.Y(n_3194)
);

AOI21xp5_ASAP7_75t_L g3195 ( 
.A1(n_3055),
.A2(n_1551),
.B(n_1543),
.Y(n_3195)
);

INVxp67_ASAP7_75t_L g3196 ( 
.A(n_3114),
.Y(n_3196)
);

INVx1_ASAP7_75t_L g3197 ( 
.A(n_3062),
.Y(n_3197)
);

AOI221xp5_ASAP7_75t_L g3198 ( 
.A1(n_3048),
.A2(n_141),
.B1(n_144),
.B2(n_145),
.C(n_146),
.Y(n_3198)
);

OA21x2_ASAP7_75t_L g3199 ( 
.A1(n_3083),
.A2(n_146),
.B(n_147),
.Y(n_3199)
);

NAND2xp5_ASAP7_75t_L g3200 ( 
.A(n_3062),
.B(n_3065),
.Y(n_3200)
);

O2A1O1Ixp33_ASAP7_75t_SL g3201 ( 
.A1(n_2995),
.A2(n_149),
.B(n_150),
.C(n_151),
.Y(n_3201)
);

AOI22x1_ASAP7_75t_L g3202 ( 
.A1(n_3130),
.A2(n_149),
.B1(n_152),
.B2(n_153),
.Y(n_3202)
);

AOI22xp5_ASAP7_75t_L g3203 ( 
.A1(n_3035),
.A2(n_153),
.B1(n_155),
.B2(n_156),
.Y(n_3203)
);

INVx1_ASAP7_75t_L g3204 ( 
.A(n_3031),
.Y(n_3204)
);

AOI21xp5_ASAP7_75t_L g3205 ( 
.A1(n_3069),
.A2(n_1574),
.B(n_1478),
.Y(n_3205)
);

CKINVDCx8_ASAP7_75t_R g3206 ( 
.A(n_2985),
.Y(n_3206)
);

OAI21x1_ASAP7_75t_L g3207 ( 
.A1(n_3006),
.A2(n_372),
.B(n_370),
.Y(n_3207)
);

O2A1O1Ixp33_ASAP7_75t_L g3208 ( 
.A1(n_3035),
.A2(n_157),
.B(n_158),
.C(n_159),
.Y(n_3208)
);

OAI21x1_ASAP7_75t_L g3209 ( 
.A1(n_3075),
.A2(n_376),
.B(n_375),
.Y(n_3209)
);

AOI21xp5_ASAP7_75t_L g3210 ( 
.A1(n_3080),
.A2(n_1574),
.B(n_1478),
.Y(n_3210)
);

AOI21xp5_ASAP7_75t_L g3211 ( 
.A1(n_3080),
.A2(n_1574),
.B(n_1478),
.Y(n_3211)
);

BUFx6f_ASAP7_75t_L g3212 ( 
.A(n_2985),
.Y(n_3212)
);

INVx3_ASAP7_75t_L g3213 ( 
.A(n_3032),
.Y(n_3213)
);

AOI21xp5_ASAP7_75t_L g3214 ( 
.A1(n_3140),
.A2(n_1478),
.B(n_1465),
.Y(n_3214)
);

BUFx3_ASAP7_75t_L g3215 ( 
.A(n_3087),
.Y(n_3215)
);

NOR2xp33_ASAP7_75t_SL g3216 ( 
.A(n_3026),
.B(n_160),
.Y(n_3216)
);

INVx2_ASAP7_75t_L g3217 ( 
.A(n_3040),
.Y(n_3217)
);

OAI21x1_ASAP7_75t_L g3218 ( 
.A1(n_3018),
.A2(n_382),
.B(n_381),
.Y(n_3218)
);

INVx1_ASAP7_75t_SL g3219 ( 
.A(n_3017),
.Y(n_3219)
);

AO21x2_ASAP7_75t_L g3220 ( 
.A1(n_3099),
.A2(n_3106),
.B(n_3119),
.Y(n_3220)
);

BUFx12f_ASAP7_75t_L g3221 ( 
.A(n_2985),
.Y(n_3221)
);

INVx2_ASAP7_75t_L g3222 ( 
.A(n_2993),
.Y(n_3222)
);

OAI21xp33_ASAP7_75t_L g3223 ( 
.A1(n_3102),
.A2(n_161),
.B(n_162),
.Y(n_3223)
);

AOI21xp5_ASAP7_75t_L g3224 ( 
.A1(n_3140),
.A2(n_1465),
.B(n_1458),
.Y(n_3224)
);

NOR2xp33_ASAP7_75t_L g3225 ( 
.A(n_3000),
.B(n_161),
.Y(n_3225)
);

AOI221xp5_ASAP7_75t_SL g3226 ( 
.A1(n_2984),
.A2(n_3124),
.B1(n_3071),
.B2(n_3079),
.C(n_3077),
.Y(n_3226)
);

AO31x2_ASAP7_75t_L g3227 ( 
.A1(n_3084),
.A2(n_3111),
.A3(n_3113),
.B(n_3107),
.Y(n_3227)
);

AOI21x1_ASAP7_75t_L g3228 ( 
.A1(n_3067),
.A2(n_162),
.B(n_163),
.Y(n_3228)
);

OR2x6_ASAP7_75t_L g3229 ( 
.A(n_2998),
.B(n_1465),
.Y(n_3229)
);

OAI21x1_ASAP7_75t_L g3230 ( 
.A1(n_3091),
.A2(n_439),
.B(n_437),
.Y(n_3230)
);

O2A1O1Ixp5_ASAP7_75t_SL g3231 ( 
.A1(n_3070),
.A2(n_164),
.B(n_165),
.C(n_166),
.Y(n_3231)
);

INVx1_ASAP7_75t_L g3232 ( 
.A(n_3076),
.Y(n_3232)
);

NAND2xp5_ASAP7_75t_L g3233 ( 
.A(n_2988),
.B(n_164),
.Y(n_3233)
);

AOI221x1_ASAP7_75t_L g3234 ( 
.A1(n_3112),
.A2(n_166),
.B1(n_167),
.B2(n_168),
.C(n_169),
.Y(n_3234)
);

OAI21x1_ASAP7_75t_L g3235 ( 
.A1(n_3088),
.A2(n_436),
.B(n_435),
.Y(n_3235)
);

OAI21x1_ASAP7_75t_L g3236 ( 
.A1(n_3020),
.A2(n_434),
.B(n_430),
.Y(n_3236)
);

OAI21x1_ASAP7_75t_L g3237 ( 
.A1(n_3003),
.A2(n_424),
.B(n_421),
.Y(n_3237)
);

AOI22xp33_ASAP7_75t_L g3238 ( 
.A1(n_3007),
.A2(n_1453),
.B1(n_1450),
.B2(n_1449),
.Y(n_3238)
);

OAI22xp33_ASAP7_75t_L g3239 ( 
.A1(n_3115),
.A2(n_167),
.B1(n_168),
.B2(n_170),
.Y(n_3239)
);

NAND2xp5_ASAP7_75t_L g3240 ( 
.A(n_3027),
.B(n_170),
.Y(n_3240)
);

NOR2xp33_ASAP7_75t_L g3241 ( 
.A(n_3108),
.B(n_172),
.Y(n_3241)
);

AOI21xp5_ASAP7_75t_L g3242 ( 
.A1(n_3066),
.A2(n_1458),
.B(n_1453),
.Y(n_3242)
);

NOR3xp33_ASAP7_75t_L g3243 ( 
.A(n_3095),
.B(n_173),
.C(n_174),
.Y(n_3243)
);

AND2x2_ASAP7_75t_L g3244 ( 
.A(n_2987),
.B(n_174),
.Y(n_3244)
);

INVx1_ASAP7_75t_L g3245 ( 
.A(n_3030),
.Y(n_3245)
);

BUFx6f_ASAP7_75t_L g3246 ( 
.A(n_3089),
.Y(n_3246)
);

OAI21x1_ASAP7_75t_L g3247 ( 
.A1(n_3060),
.A2(n_417),
.B(n_416),
.Y(n_3247)
);

AOI21xp5_ASAP7_75t_L g3248 ( 
.A1(n_3066),
.A2(n_1458),
.B(n_1453),
.Y(n_3248)
);

INVx2_ASAP7_75t_L g3249 ( 
.A(n_2983),
.Y(n_3249)
);

INVx2_ASAP7_75t_SL g3250 ( 
.A(n_3089),
.Y(n_3250)
);

OAI21x1_ASAP7_75t_SL g3251 ( 
.A1(n_3077),
.A2(n_3063),
.B(n_2984),
.Y(n_3251)
);

NAND2x1p5_ASAP7_75t_L g3252 ( 
.A(n_3008),
.B(n_1449),
.Y(n_3252)
);

NOR2xp33_ASAP7_75t_L g3253 ( 
.A(n_3092),
.B(n_175),
.Y(n_3253)
);

OR2x2_ASAP7_75t_L g3254 ( 
.A(n_3039),
.B(n_3028),
.Y(n_3254)
);

AOI22xp5_ASAP7_75t_L g3255 ( 
.A1(n_3135),
.A2(n_3098),
.B1(n_3068),
.B2(n_3063),
.Y(n_3255)
);

AO31x2_ASAP7_75t_L g3256 ( 
.A1(n_3059),
.A2(n_175),
.A3(n_176),
.B(n_178),
.Y(n_3256)
);

AND2x4_ASAP7_75t_L g3257 ( 
.A(n_3116),
.B(n_178),
.Y(n_3257)
);

OAI21x1_ASAP7_75t_L g3258 ( 
.A1(n_3023),
.A2(n_414),
.B(n_413),
.Y(n_3258)
);

INVx4_ASAP7_75t_L g3259 ( 
.A(n_3059),
.Y(n_3259)
);

BUFx2_ASAP7_75t_R g3260 ( 
.A(n_3110),
.Y(n_3260)
);

INVx1_ASAP7_75t_L g3261 ( 
.A(n_2983),
.Y(n_3261)
);

OAI22xp5_ASAP7_75t_L g3262 ( 
.A1(n_3132),
.A2(n_180),
.B1(n_182),
.B2(n_183),
.Y(n_3262)
);

OAI21xp5_ASAP7_75t_L g3263 ( 
.A1(n_3105),
.A2(n_186),
.B(n_188),
.Y(n_3263)
);

NAND2xp5_ASAP7_75t_L g3264 ( 
.A(n_3085),
.B(n_189),
.Y(n_3264)
);

AO32x2_ASAP7_75t_L g3265 ( 
.A1(n_3057),
.A2(n_190),
.A3(n_194),
.B1(n_195),
.B2(n_196),
.Y(n_3265)
);

OAI21x1_ASAP7_75t_L g3266 ( 
.A1(n_3150),
.A2(n_3249),
.B(n_3261),
.Y(n_3266)
);

BUFx12f_ASAP7_75t_L g3267 ( 
.A(n_3170),
.Y(n_3267)
);

INVx4_ASAP7_75t_L g3268 ( 
.A(n_3180),
.Y(n_3268)
);

AND2x4_ASAP7_75t_L g3269 ( 
.A(n_3148),
.B(n_3179),
.Y(n_3269)
);

CKINVDCx5p33_ASAP7_75t_R g3270 ( 
.A(n_3172),
.Y(n_3270)
);

AOI221xp5_ASAP7_75t_L g3271 ( 
.A1(n_3155),
.A2(n_3068),
.B1(n_3057),
.B2(n_3073),
.C(n_3074),
.Y(n_3271)
);

OR2x6_ASAP7_75t_L g3272 ( 
.A(n_3251),
.B(n_3047),
.Y(n_3272)
);

OAI21x1_ASAP7_75t_L g3273 ( 
.A1(n_3171),
.A2(n_3047),
.B(n_3036),
.Y(n_3273)
);

BUFx3_ASAP7_75t_L g3274 ( 
.A(n_3170),
.Y(n_3274)
);

INVx2_ASAP7_75t_L g3275 ( 
.A(n_3167),
.Y(n_3275)
);

OAI22xp5_ASAP7_75t_L g3276 ( 
.A1(n_3203),
.A2(n_3164),
.B1(n_3192),
.B2(n_3263),
.Y(n_3276)
);

BUFx2_ASAP7_75t_L g3277 ( 
.A(n_3148),
.Y(n_3277)
);

OA21x2_ASAP7_75t_L g3278 ( 
.A1(n_3226),
.A2(n_3126),
.B(n_3033),
.Y(n_3278)
);

INVx1_ASAP7_75t_SL g3279 ( 
.A(n_3177),
.Y(n_3279)
);

AO21x1_ASAP7_75t_L g3280 ( 
.A1(n_3164),
.A2(n_3097),
.B(n_3126),
.Y(n_3280)
);

OA21x2_ASAP7_75t_L g3281 ( 
.A1(n_3226),
.A2(n_3174),
.B(n_3264),
.Y(n_3281)
);

OAI21x1_ASAP7_75t_L g3282 ( 
.A1(n_3224),
.A2(n_3044),
.B(n_3037),
.Y(n_3282)
);

NOR2xp67_ASAP7_75t_SL g3283 ( 
.A(n_3180),
.B(n_3089),
.Y(n_3283)
);

AND2x4_ASAP7_75t_L g3284 ( 
.A(n_3179),
.B(n_3025),
.Y(n_3284)
);

INVx2_ASAP7_75t_L g3285 ( 
.A(n_3145),
.Y(n_3285)
);

NAND2x1p5_ASAP7_75t_L g3286 ( 
.A(n_3143),
.B(n_3082),
.Y(n_3286)
);

OAI21xp5_ASAP7_75t_L g3287 ( 
.A1(n_3162),
.A2(n_3098),
.B(n_3086),
.Y(n_3287)
);

O2A1O1Ixp33_ASAP7_75t_L g3288 ( 
.A1(n_3141),
.A2(n_3086),
.B(n_3109),
.C(n_3129),
.Y(n_3288)
);

NAND2xp33_ASAP7_75t_L g3289 ( 
.A(n_3243),
.B(n_3093),
.Y(n_3289)
);

NOR2xp33_ASAP7_75t_L g3290 ( 
.A(n_3159),
.B(n_3093),
.Y(n_3290)
);

O2A1O1Ixp33_ASAP7_75t_L g3291 ( 
.A1(n_3208),
.A2(n_3129),
.B(n_3072),
.C(n_3082),
.Y(n_3291)
);

AOI22xp33_ASAP7_75t_L g3292 ( 
.A1(n_3153),
.A2(n_3072),
.B1(n_3094),
.B2(n_3004),
.Y(n_3292)
);

INVx2_ASAP7_75t_L g3293 ( 
.A(n_3149),
.Y(n_3293)
);

AO21x2_ASAP7_75t_L g3294 ( 
.A1(n_3214),
.A2(n_3119),
.B(n_3004),
.Y(n_3294)
);

INVx2_ASAP7_75t_L g3295 ( 
.A(n_3154),
.Y(n_3295)
);

OAI22xp5_ASAP7_75t_L g3296 ( 
.A1(n_3203),
.A2(n_3093),
.B1(n_3100),
.B2(n_3103),
.Y(n_3296)
);

OAI21x1_ASAP7_75t_L g3297 ( 
.A1(n_3242),
.A2(n_3117),
.B(n_3118),
.Y(n_3297)
);

INVx3_ASAP7_75t_L g3298 ( 
.A(n_3259),
.Y(n_3298)
);

CKINVDCx6p67_ASAP7_75t_R g3299 ( 
.A(n_3180),
.Y(n_3299)
);

OAI21x1_ASAP7_75t_L g3300 ( 
.A1(n_3248),
.A2(n_3120),
.B(n_3123),
.Y(n_3300)
);

CKINVDCx5p33_ASAP7_75t_R g3301 ( 
.A(n_3159),
.Y(n_3301)
);

AOI221xp5_ASAP7_75t_L g3302 ( 
.A1(n_3223),
.A2(n_3103),
.B1(n_3100),
.B2(n_3094),
.C(n_201),
.Y(n_3302)
);

AO21x2_ASAP7_75t_L g3303 ( 
.A1(n_3147),
.A2(n_3134),
.B(n_3137),
.Y(n_3303)
);

AND2x4_ASAP7_75t_L g3304 ( 
.A(n_3213),
.B(n_3025),
.Y(n_3304)
);

AOI22xp33_ASAP7_75t_L g3305 ( 
.A1(n_3165),
.A2(n_3103),
.B1(n_3100),
.B2(n_3046),
.Y(n_3305)
);

BUFx8_ASAP7_75t_L g3306 ( 
.A(n_3182),
.Y(n_3306)
);

INVx2_ASAP7_75t_L g3307 ( 
.A(n_3232),
.Y(n_3307)
);

NAND2xp5_ASAP7_75t_L g3308 ( 
.A(n_3219),
.B(n_3046),
.Y(n_3308)
);

NOR2xp33_ASAP7_75t_SL g3309 ( 
.A(n_3260),
.B(n_3012),
.Y(n_3309)
);

OAI21x1_ASAP7_75t_L g3310 ( 
.A1(n_3228),
.A2(n_3090),
.B(n_3025),
.Y(n_3310)
);

NOR2xp33_ASAP7_75t_L g3311 ( 
.A(n_3151),
.B(n_195),
.Y(n_3311)
);

INVx1_ASAP7_75t_SL g3312 ( 
.A(n_3219),
.Y(n_3312)
);

AOI21xp5_ASAP7_75t_L g3313 ( 
.A1(n_3152),
.A2(n_3061),
.B(n_3054),
.Y(n_3313)
);

INVx1_ASAP7_75t_L g3314 ( 
.A(n_3204),
.Y(n_3314)
);

BUFx3_ASAP7_75t_L g3315 ( 
.A(n_3173),
.Y(n_3315)
);

BUFx4f_ASAP7_75t_L g3316 ( 
.A(n_3146),
.Y(n_3316)
);

INVxp67_ASAP7_75t_SL g3317 ( 
.A(n_3163),
.Y(n_3317)
);

BUFx3_ASAP7_75t_L g3318 ( 
.A(n_3183),
.Y(n_3318)
);

NAND2x1p5_ASAP7_75t_L g3319 ( 
.A(n_3143),
.B(n_3061),
.Y(n_3319)
);

INVx2_ASAP7_75t_L g3320 ( 
.A(n_3217),
.Y(n_3320)
);

AOI22xp33_ASAP7_75t_L g3321 ( 
.A1(n_3165),
.A2(n_196),
.B1(n_200),
.B2(n_202),
.Y(n_3321)
);

AOI22xp33_ASAP7_75t_SL g3322 ( 
.A1(n_3216),
.A2(n_3012),
.B1(n_3125),
.B2(n_3054),
.Y(n_3322)
);

AOI21xp5_ASAP7_75t_L g3323 ( 
.A1(n_3156),
.A2(n_3125),
.B(n_3056),
.Y(n_3323)
);

OA21x2_ASAP7_75t_L g3324 ( 
.A1(n_3160),
.A2(n_3128),
.B(n_202),
.Y(n_3324)
);

OA21x2_ASAP7_75t_L g3325 ( 
.A1(n_3166),
.A2(n_3128),
.B(n_203),
.Y(n_3325)
);

OAI22xp33_ASAP7_75t_L g3326 ( 
.A1(n_3216),
.A2(n_200),
.B1(n_204),
.B2(n_206),
.Y(n_3326)
);

OAI22xp5_ASAP7_75t_L g3327 ( 
.A1(n_3255),
.A2(n_206),
.B1(n_207),
.B2(n_209),
.Y(n_3327)
);

INVx2_ASAP7_75t_L g3328 ( 
.A(n_3222),
.Y(n_3328)
);

INVx1_ASAP7_75t_L g3329 ( 
.A(n_3245),
.Y(n_3329)
);

OR2x6_ASAP7_75t_L g3330 ( 
.A(n_3186),
.B(n_1450),
.Y(n_3330)
);

OAI21x1_ASAP7_75t_L g3331 ( 
.A1(n_3168),
.A2(n_207),
.B(n_209),
.Y(n_3331)
);

INVx3_ASAP7_75t_L g3332 ( 
.A(n_3259),
.Y(n_3332)
);

OA21x2_ASAP7_75t_L g3333 ( 
.A1(n_3190),
.A2(n_211),
.B(n_213),
.Y(n_3333)
);

OA21x2_ASAP7_75t_L g3334 ( 
.A1(n_3195),
.A2(n_214),
.B(n_215),
.Y(n_3334)
);

OAI222xp33_ASAP7_75t_L g3335 ( 
.A1(n_3255),
.A2(n_214),
.B1(n_215),
.B2(n_216),
.C1(n_217),
.C2(n_219),
.Y(n_3335)
);

OAI21xp5_ASAP7_75t_L g3336 ( 
.A1(n_3187),
.A2(n_219),
.B(n_220),
.Y(n_3336)
);

AO21x2_ASAP7_75t_L g3337 ( 
.A1(n_3175),
.A2(n_220),
.B(n_221),
.Y(n_3337)
);

HB1xp67_ASAP7_75t_L g3338 ( 
.A(n_3185),
.Y(n_3338)
);

HB1xp67_ASAP7_75t_L g3339 ( 
.A(n_3199),
.Y(n_3339)
);

INVx2_ASAP7_75t_L g3340 ( 
.A(n_3197),
.Y(n_3340)
);

NAND2xp5_ASAP7_75t_L g3341 ( 
.A(n_3200),
.B(n_223),
.Y(n_3341)
);

AOI22xp5_ASAP7_75t_L g3342 ( 
.A1(n_3161),
.A2(n_223),
.B1(n_224),
.B2(n_226),
.Y(n_3342)
);

INVx1_ASAP7_75t_L g3343 ( 
.A(n_3196),
.Y(n_3343)
);

NAND3xp33_ASAP7_75t_L g3344 ( 
.A(n_3184),
.B(n_224),
.C(n_226),
.Y(n_3344)
);

OAI21xp5_ASAP7_75t_L g3345 ( 
.A1(n_3157),
.A2(n_228),
.B(n_229),
.Y(n_3345)
);

INVx2_ASAP7_75t_SL g3346 ( 
.A(n_3215),
.Y(n_3346)
);

OAI22xp5_ASAP7_75t_L g3347 ( 
.A1(n_3198),
.A2(n_231),
.B1(n_232),
.B2(n_233),
.Y(n_3347)
);

OAI21xp5_ASAP7_75t_L g3348 ( 
.A1(n_3144),
.A2(n_232),
.B(n_233),
.Y(n_3348)
);

OAI21x1_ASAP7_75t_L g3349 ( 
.A1(n_3209),
.A2(n_234),
.B(n_235),
.Y(n_3349)
);

OA21x2_ASAP7_75t_L g3350 ( 
.A1(n_3169),
.A2(n_235),
.B(n_236),
.Y(n_3350)
);

NAND2xp5_ASAP7_75t_L g3351 ( 
.A(n_3254),
.B(n_237),
.Y(n_3351)
);

AOI22xp33_ASAP7_75t_L g3352 ( 
.A1(n_3223),
.A2(n_238),
.B1(n_239),
.B2(n_241),
.Y(n_3352)
);

OAI22xp5_ASAP7_75t_L g3353 ( 
.A1(n_3202),
.A2(n_239),
.B1(n_241),
.B2(n_242),
.Y(n_3353)
);

INVx2_ASAP7_75t_L g3354 ( 
.A(n_3199),
.Y(n_3354)
);

HB1xp67_ASAP7_75t_L g3355 ( 
.A(n_3186),
.Y(n_3355)
);

CKINVDCx5p33_ASAP7_75t_R g3356 ( 
.A(n_3221),
.Y(n_3356)
);

AOI21xp5_ASAP7_75t_L g3357 ( 
.A1(n_3210),
.A2(n_410),
.B(n_406),
.Y(n_3357)
);

OR2x2_ASAP7_75t_L g3358 ( 
.A(n_3158),
.B(n_245),
.Y(n_3358)
);

OAI21x1_ASAP7_75t_SL g3359 ( 
.A1(n_3181),
.A2(n_245),
.B(n_246),
.Y(n_3359)
);

OAI21x1_ASAP7_75t_L g3360 ( 
.A1(n_3211),
.A2(n_251),
.B(n_252),
.Y(n_3360)
);

AO21x2_ASAP7_75t_L g3361 ( 
.A1(n_3189),
.A2(n_255),
.B(n_256),
.Y(n_3361)
);

INVx1_ASAP7_75t_L g3362 ( 
.A(n_3193),
.Y(n_3362)
);

OAI22xp5_ASAP7_75t_L g3363 ( 
.A1(n_3206),
.A2(n_255),
.B1(n_256),
.B2(n_257),
.Y(n_3363)
);

NAND3xp33_ASAP7_75t_L g3364 ( 
.A(n_3241),
.B(n_3225),
.C(n_3234),
.Y(n_3364)
);

AOI21xp5_ASAP7_75t_R g3365 ( 
.A1(n_3262),
.A2(n_259),
.B(n_260),
.Y(n_3365)
);

BUFx6f_ASAP7_75t_L g3366 ( 
.A(n_3212),
.Y(n_3366)
);

INVx1_ASAP7_75t_L g3367 ( 
.A(n_3194),
.Y(n_3367)
);

AO31x2_ASAP7_75t_L g3368 ( 
.A1(n_3354),
.A2(n_3233),
.A3(n_3240),
.B(n_3253),
.Y(n_3368)
);

AOI21xp33_ASAP7_75t_SL g3369 ( 
.A1(n_3301),
.A2(n_3239),
.B(n_3146),
.Y(n_3369)
);

OA21x2_ASAP7_75t_L g3370 ( 
.A1(n_3317),
.A2(n_3237),
.B(n_3247),
.Y(n_3370)
);

AOI21xp5_ASAP7_75t_L g3371 ( 
.A1(n_3289),
.A2(n_3178),
.B(n_3176),
.Y(n_3371)
);

BUFx2_ASAP7_75t_L g3372 ( 
.A(n_3268),
.Y(n_3372)
);

AOI21xp5_ASAP7_75t_L g3373 ( 
.A1(n_3289),
.A2(n_3201),
.B(n_3188),
.Y(n_3373)
);

AO21x2_ASAP7_75t_L g3374 ( 
.A1(n_3317),
.A2(n_3142),
.B(n_3205),
.Y(n_3374)
);

BUFx10_ASAP7_75t_L g3375 ( 
.A(n_3290),
.Y(n_3375)
);

BUFx2_ASAP7_75t_R g3376 ( 
.A(n_3301),
.Y(n_3376)
);

OR2x6_ASAP7_75t_L g3377 ( 
.A(n_3268),
.B(n_3229),
.Y(n_3377)
);

BUFx2_ASAP7_75t_L g3378 ( 
.A(n_3299),
.Y(n_3378)
);

OAI21x1_ASAP7_75t_L g3379 ( 
.A1(n_3266),
.A2(n_3236),
.B(n_3218),
.Y(n_3379)
);

AOI21xp5_ASAP7_75t_L g3380 ( 
.A1(n_3324),
.A2(n_3220),
.B(n_3229),
.Y(n_3380)
);

OAI21xp5_ASAP7_75t_L g3381 ( 
.A1(n_3364),
.A2(n_3231),
.B(n_3257),
.Y(n_3381)
);

INVxp67_ASAP7_75t_SL g3382 ( 
.A(n_3338),
.Y(n_3382)
);

AND2x2_ASAP7_75t_L g3383 ( 
.A(n_3269),
.B(n_3250),
.Y(n_3383)
);

AO21x2_ASAP7_75t_L g3384 ( 
.A1(n_3338),
.A2(n_3207),
.B(n_3258),
.Y(n_3384)
);

NAND2xp5_ASAP7_75t_L g3385 ( 
.A(n_3312),
.B(n_3244),
.Y(n_3385)
);

AOI21x1_ASAP7_75t_L g3386 ( 
.A1(n_3339),
.A2(n_3229),
.B(n_3230),
.Y(n_3386)
);

HB1xp67_ASAP7_75t_L g3387 ( 
.A(n_3339),
.Y(n_3387)
);

NAND2xp5_ASAP7_75t_L g3388 ( 
.A(n_3362),
.B(n_3194),
.Y(n_3388)
);

INVx1_ASAP7_75t_SL g3389 ( 
.A(n_3270),
.Y(n_3389)
);

NAND2xp5_ASAP7_75t_L g3390 ( 
.A(n_3281),
.B(n_3343),
.Y(n_3390)
);

INVx1_ASAP7_75t_L g3391 ( 
.A(n_3285),
.Y(n_3391)
);

AND2x4_ASAP7_75t_L g3392 ( 
.A(n_3298),
.B(n_3246),
.Y(n_3392)
);

OR2x6_ASAP7_75t_L g3393 ( 
.A(n_3272),
.B(n_3252),
.Y(n_3393)
);

INVx1_ASAP7_75t_L g3394 ( 
.A(n_3293),
.Y(n_3394)
);

OAI21x1_ASAP7_75t_L g3395 ( 
.A1(n_3319),
.A2(n_3235),
.B(n_3238),
.Y(n_3395)
);

INVx1_ASAP7_75t_L g3396 ( 
.A(n_3295),
.Y(n_3396)
);

BUFx6f_ASAP7_75t_L g3397 ( 
.A(n_3267),
.Y(n_3397)
);

OR2x2_ASAP7_75t_L g3398 ( 
.A(n_3308),
.B(n_3194),
.Y(n_3398)
);

INVx1_ASAP7_75t_L g3399 ( 
.A(n_3295),
.Y(n_3399)
);

OA21x2_ASAP7_75t_L g3400 ( 
.A1(n_3354),
.A2(n_3265),
.B(n_3256),
.Y(n_3400)
);

INVxp67_ASAP7_75t_L g3401 ( 
.A(n_3350),
.Y(n_3401)
);

OAI21xp5_ASAP7_75t_L g3402 ( 
.A1(n_3344),
.A2(n_3336),
.B(n_3348),
.Y(n_3402)
);

INVx2_ASAP7_75t_L g3403 ( 
.A(n_3307),
.Y(n_3403)
);

OR2x6_ASAP7_75t_L g3404 ( 
.A(n_3272),
.B(n_3246),
.Y(n_3404)
);

INVx3_ASAP7_75t_L g3405 ( 
.A(n_3269),
.Y(n_3405)
);

BUFx2_ASAP7_75t_L g3406 ( 
.A(n_3272),
.Y(n_3406)
);

OA21x2_ASAP7_75t_L g3407 ( 
.A1(n_3355),
.A2(n_3256),
.B(n_3191),
.Y(n_3407)
);

OAI221xp5_ASAP7_75t_SL g3408 ( 
.A1(n_3321),
.A2(n_3191),
.B1(n_262),
.B2(n_264),
.C(n_265),
.Y(n_3408)
);

BUFx8_ASAP7_75t_L g3409 ( 
.A(n_3267),
.Y(n_3409)
);

AOI21xp5_ASAP7_75t_L g3410 ( 
.A1(n_3324),
.A2(n_3246),
.B(n_3227),
.Y(n_3410)
);

AOI21xp5_ASAP7_75t_L g3411 ( 
.A1(n_3313),
.A2(n_3227),
.B(n_262),
.Y(n_3411)
);

INVx2_ASAP7_75t_L g3412 ( 
.A(n_3340),
.Y(n_3412)
);

OAI21xp5_ASAP7_75t_L g3413 ( 
.A1(n_3311),
.A2(n_3227),
.B(n_265),
.Y(n_3413)
);

OA21x2_ASAP7_75t_L g3414 ( 
.A1(n_3355),
.A2(n_261),
.B(n_266),
.Y(n_3414)
);

OAI21x1_ASAP7_75t_L g3415 ( 
.A1(n_3310),
.A2(n_261),
.B(n_267),
.Y(n_3415)
);

NAND2xp5_ASAP7_75t_L g3416 ( 
.A(n_3314),
.B(n_268),
.Y(n_3416)
);

AOI21xp5_ASAP7_75t_L g3417 ( 
.A1(n_3357),
.A2(n_268),
.B(n_269),
.Y(n_3417)
);

NAND2xp5_ASAP7_75t_L g3418 ( 
.A(n_3329),
.B(n_270),
.Y(n_3418)
);

NOR2xp33_ASAP7_75t_L g3419 ( 
.A(n_3290),
.B(n_271),
.Y(n_3419)
);

INVx5_ASAP7_75t_L g3420 ( 
.A(n_3330),
.Y(n_3420)
);

INVx2_ASAP7_75t_L g3421 ( 
.A(n_3275),
.Y(n_3421)
);

OAI21x1_ASAP7_75t_L g3422 ( 
.A1(n_3273),
.A2(n_271),
.B(n_272),
.Y(n_3422)
);

BUFx12f_ASAP7_75t_L g3423 ( 
.A(n_3270),
.Y(n_3423)
);

INVx3_ASAP7_75t_L g3424 ( 
.A(n_3269),
.Y(n_3424)
);

INVx2_ASAP7_75t_L g3425 ( 
.A(n_3275),
.Y(n_3425)
);

A2O1A1Ixp33_ASAP7_75t_L g3426 ( 
.A1(n_3345),
.A2(n_272),
.B(n_273),
.C(n_274),
.Y(n_3426)
);

OAI21x1_ASAP7_75t_L g3427 ( 
.A1(n_3286),
.A2(n_275),
.B(n_276),
.Y(n_3427)
);

AND2x2_ASAP7_75t_L g3428 ( 
.A(n_3277),
.B(n_276),
.Y(n_3428)
);

INVx2_ASAP7_75t_L g3429 ( 
.A(n_3284),
.Y(n_3429)
);

AO31x2_ASAP7_75t_L g3430 ( 
.A1(n_3280),
.A2(n_279),
.A3(n_280),
.B(n_282),
.Y(n_3430)
);

AND2x2_ASAP7_75t_L g3431 ( 
.A(n_3298),
.B(n_279),
.Y(n_3431)
);

AND2x4_ASAP7_75t_L g3432 ( 
.A(n_3332),
.B(n_280),
.Y(n_3432)
);

AOI21x1_ASAP7_75t_L g3433 ( 
.A1(n_3283),
.A2(n_283),
.B(n_284),
.Y(n_3433)
);

INVx2_ASAP7_75t_L g3434 ( 
.A(n_3284),
.Y(n_3434)
);

NAND2xp5_ASAP7_75t_L g3435 ( 
.A(n_3320),
.B(n_283),
.Y(n_3435)
);

OAI22xp5_ASAP7_75t_L g3436 ( 
.A1(n_3321),
.A2(n_284),
.B1(n_285),
.B2(n_286),
.Y(n_3436)
);

OAI21x1_ASAP7_75t_L g3437 ( 
.A1(n_3286),
.A2(n_391),
.B(n_394),
.Y(n_3437)
);

AO21x2_ASAP7_75t_L g3438 ( 
.A1(n_3367),
.A2(n_396),
.B(n_397),
.Y(n_3438)
);

OA21x2_ASAP7_75t_L g3439 ( 
.A1(n_3284),
.A2(n_402),
.B(n_398),
.Y(n_3439)
);

HB1xp67_ASAP7_75t_L g3440 ( 
.A(n_3350),
.Y(n_3440)
);

CKINVDCx5p33_ASAP7_75t_R g3441 ( 
.A(n_3356),
.Y(n_3441)
);

OAI22xp33_ASAP7_75t_L g3442 ( 
.A1(n_3302),
.A2(n_3309),
.B1(n_3342),
.B2(n_3326),
.Y(n_3442)
);

INVx1_ASAP7_75t_L g3443 ( 
.A(n_3328),
.Y(n_3443)
);

AOI21xp5_ASAP7_75t_L g3444 ( 
.A1(n_3333),
.A2(n_401),
.B(n_3334),
.Y(n_3444)
);

INVx2_ASAP7_75t_L g3445 ( 
.A(n_3328),
.Y(n_3445)
);

INVx3_ASAP7_75t_L g3446 ( 
.A(n_3332),
.Y(n_3446)
);

INVx2_ASAP7_75t_L g3447 ( 
.A(n_3304),
.Y(n_3447)
);

NOR2xp33_ASAP7_75t_L g3448 ( 
.A(n_3341),
.B(n_3351),
.Y(n_3448)
);

NAND2xp5_ASAP7_75t_L g3449 ( 
.A(n_3337),
.B(n_3361),
.Y(n_3449)
);

INVx3_ASAP7_75t_SL g3450 ( 
.A(n_3356),
.Y(n_3450)
);

NAND2x1p5_ASAP7_75t_L g3451 ( 
.A(n_3304),
.B(n_3325),
.Y(n_3451)
);

BUFx2_ASAP7_75t_L g3452 ( 
.A(n_3318),
.Y(n_3452)
);

AND2x2_ASAP7_75t_L g3453 ( 
.A(n_3346),
.B(n_3279),
.Y(n_3453)
);

INVx1_ASAP7_75t_L g3454 ( 
.A(n_3304),
.Y(n_3454)
);

NOR2xp33_ASAP7_75t_L g3455 ( 
.A(n_3358),
.B(n_3274),
.Y(n_3455)
);

AOI21xp5_ASAP7_75t_L g3456 ( 
.A1(n_3333),
.A2(n_3334),
.B(n_3287),
.Y(n_3456)
);

OAI21xp5_ASAP7_75t_L g3457 ( 
.A1(n_3456),
.A2(n_3327),
.B(n_3352),
.Y(n_3457)
);

AOI22xp33_ASAP7_75t_L g3458 ( 
.A1(n_3402),
.A2(n_3347),
.B1(n_3352),
.B2(n_3353),
.Y(n_3458)
);

OAI22xp5_ASAP7_75t_L g3459 ( 
.A1(n_3408),
.A2(n_3365),
.B1(n_3305),
.B2(n_3292),
.Y(n_3459)
);

BUFx6f_ASAP7_75t_SL g3460 ( 
.A(n_3397),
.Y(n_3460)
);

AOI222xp33_ASAP7_75t_L g3461 ( 
.A1(n_3442),
.A2(n_3335),
.B1(n_3326),
.B2(n_3363),
.C1(n_3296),
.C2(n_3359),
.Y(n_3461)
);

BUFx2_ASAP7_75t_L g3462 ( 
.A(n_3378),
.Y(n_3462)
);

OAI21xp33_ASAP7_75t_L g3463 ( 
.A1(n_3413),
.A2(n_3305),
.B(n_3292),
.Y(n_3463)
);

AOI22xp33_ASAP7_75t_L g3464 ( 
.A1(n_3442),
.A2(n_3333),
.B1(n_3334),
.B2(n_3271),
.Y(n_3464)
);

AOI22xp33_ASAP7_75t_L g3465 ( 
.A1(n_3436),
.A2(n_3419),
.B1(n_3371),
.B2(n_3448),
.Y(n_3465)
);

INVxp67_ASAP7_75t_L g3466 ( 
.A(n_3376),
.Y(n_3466)
);

NAND2xp5_ASAP7_75t_L g3467 ( 
.A(n_3368),
.B(n_3322),
.Y(n_3467)
);

AOI22xp33_ASAP7_75t_L g3468 ( 
.A1(n_3419),
.A2(n_3325),
.B1(n_3360),
.B2(n_3278),
.Y(n_3468)
);

BUFx3_ASAP7_75t_L g3469 ( 
.A(n_3409),
.Y(n_3469)
);

AND2x2_ASAP7_75t_L g3470 ( 
.A(n_3383),
.B(n_3315),
.Y(n_3470)
);

AND2x2_ASAP7_75t_L g3471 ( 
.A(n_3406),
.B(n_3318),
.Y(n_3471)
);

NOR2x1_ASAP7_75t_L g3472 ( 
.A(n_3372),
.B(n_3330),
.Y(n_3472)
);

AND2x2_ASAP7_75t_L g3473 ( 
.A(n_3375),
.B(n_3316),
.Y(n_3473)
);

BUFx3_ASAP7_75t_L g3474 ( 
.A(n_3409),
.Y(n_3474)
);

OAI21xp33_ASAP7_75t_L g3475 ( 
.A1(n_3426),
.A2(n_3323),
.B(n_3331),
.Y(n_3475)
);

BUFx6f_ASAP7_75t_SL g3476 ( 
.A(n_3397),
.Y(n_3476)
);

OAI21xp5_ASAP7_75t_SL g3477 ( 
.A1(n_3426),
.A2(n_3288),
.B(n_3291),
.Y(n_3477)
);

CKINVDCx5p33_ASAP7_75t_R g3478 ( 
.A(n_3423),
.Y(n_3478)
);

CKINVDCx5p33_ASAP7_75t_R g3479 ( 
.A(n_3441),
.Y(n_3479)
);

CKINVDCx20_ASAP7_75t_R g3480 ( 
.A(n_3450),
.Y(n_3480)
);

NAND2xp5_ASAP7_75t_SL g3481 ( 
.A(n_3375),
.B(n_3306),
.Y(n_3481)
);

HB1xp67_ASAP7_75t_L g3482 ( 
.A(n_3387),
.Y(n_3482)
);

AOI22xp33_ASAP7_75t_L g3483 ( 
.A1(n_3448),
.A2(n_3303),
.B1(n_3294),
.B2(n_3349),
.Y(n_3483)
);

BUFx12f_ASAP7_75t_L g3484 ( 
.A(n_3397),
.Y(n_3484)
);

NOR2x1_ASAP7_75t_R g3485 ( 
.A(n_3397),
.B(n_3366),
.Y(n_3485)
);

OAI22xp5_ASAP7_75t_L g3486 ( 
.A1(n_3373),
.A2(n_3300),
.B1(n_3297),
.B2(n_3282),
.Y(n_3486)
);

AND2x2_ASAP7_75t_L g3487 ( 
.A(n_3452),
.B(n_3405),
.Y(n_3487)
);

AOI22xp33_ASAP7_75t_L g3488 ( 
.A1(n_3417),
.A2(n_3381),
.B1(n_3449),
.B2(n_3455),
.Y(n_3488)
);

OAI21xp5_ASAP7_75t_SL g3489 ( 
.A1(n_3369),
.A2(n_3417),
.B(n_3444),
.Y(n_3489)
);

AOI22xp33_ASAP7_75t_SL g3490 ( 
.A1(n_3440),
.A2(n_3414),
.B1(n_3400),
.B2(n_3382),
.Y(n_3490)
);

AOI222xp33_ASAP7_75t_L g3491 ( 
.A1(n_3401),
.A2(n_3390),
.B1(n_3382),
.B2(n_3418),
.C1(n_3416),
.C2(n_3388),
.Y(n_3491)
);

AOI22xp5_ASAP7_75t_L g3492 ( 
.A1(n_3453),
.A2(n_3404),
.B1(n_3393),
.B2(n_3389),
.Y(n_3492)
);

AOI22xp33_ASAP7_75t_L g3493 ( 
.A1(n_3411),
.A2(n_3400),
.B1(n_3444),
.B2(n_3407),
.Y(n_3493)
);

OAI211xp5_ASAP7_75t_L g3494 ( 
.A1(n_3380),
.A2(n_3387),
.B(n_3400),
.C(n_3410),
.Y(n_3494)
);

OAI21xp5_ASAP7_75t_SL g3495 ( 
.A1(n_3380),
.A2(n_3433),
.B(n_3410),
.Y(n_3495)
);

AND2x2_ASAP7_75t_L g3496 ( 
.A(n_3405),
.B(n_3424),
.Y(n_3496)
);

AOI22xp33_ASAP7_75t_SL g3497 ( 
.A1(n_3438),
.A2(n_3439),
.B1(n_3407),
.B2(n_3384),
.Y(n_3497)
);

BUFx4f_ASAP7_75t_SL g3498 ( 
.A(n_3450),
.Y(n_3498)
);

OAI21xp33_ASAP7_75t_L g3499 ( 
.A1(n_3398),
.A2(n_3435),
.B(n_3451),
.Y(n_3499)
);

INVx2_ASAP7_75t_SL g3500 ( 
.A(n_3392),
.Y(n_3500)
);

AOI22xp33_ASAP7_75t_L g3501 ( 
.A1(n_3407),
.A2(n_3438),
.B1(n_3374),
.B2(n_3384),
.Y(n_3501)
);

AOI22xp33_ASAP7_75t_SL g3502 ( 
.A1(n_3439),
.A2(n_3370),
.B1(n_3432),
.B2(n_3374),
.Y(n_3502)
);

CKINVDCx5p33_ASAP7_75t_R g3503 ( 
.A(n_3432),
.Y(n_3503)
);

INVx1_ASAP7_75t_L g3504 ( 
.A(n_3391),
.Y(n_3504)
);

AOI22xp5_ASAP7_75t_L g3505 ( 
.A1(n_3404),
.A2(n_3393),
.B1(n_3377),
.B2(n_3424),
.Y(n_3505)
);

AOI22xp33_ASAP7_75t_L g3506 ( 
.A1(n_3385),
.A2(n_3370),
.B1(n_3439),
.B2(n_3415),
.Y(n_3506)
);

OAI21xp5_ASAP7_75t_SL g3507 ( 
.A1(n_3451),
.A2(n_3428),
.B(n_3386),
.Y(n_3507)
);

BUFx4f_ASAP7_75t_SL g3508 ( 
.A(n_3431),
.Y(n_3508)
);

AOI22xp33_ASAP7_75t_L g3509 ( 
.A1(n_3370),
.A2(n_3422),
.B1(n_3427),
.B2(n_3395),
.Y(n_3509)
);

CKINVDCx5p33_ASAP7_75t_R g3510 ( 
.A(n_3446),
.Y(n_3510)
);

OAI21xp33_ASAP7_75t_L g3511 ( 
.A1(n_3454),
.A2(n_3429),
.B(n_3434),
.Y(n_3511)
);

OAI22xp33_ASAP7_75t_L g3512 ( 
.A1(n_3420),
.A2(n_3377),
.B1(n_3430),
.B2(n_3434),
.Y(n_3512)
);

OAI222xp33_ASAP7_75t_L g3513 ( 
.A1(n_3420),
.A2(n_3429),
.B1(n_3447),
.B2(n_3430),
.C1(n_3443),
.C2(n_3394),
.Y(n_3513)
);

CKINVDCx5p33_ASAP7_75t_R g3514 ( 
.A(n_3420),
.Y(n_3514)
);

CKINVDCx20_ASAP7_75t_R g3515 ( 
.A(n_3396),
.Y(n_3515)
);

AOI22xp33_ASAP7_75t_L g3516 ( 
.A1(n_3437),
.A2(n_3445),
.B1(n_3421),
.B2(n_3425),
.Y(n_3516)
);

OAI22xp33_ASAP7_75t_L g3517 ( 
.A1(n_3430),
.A2(n_3399),
.B1(n_3412),
.B2(n_3403),
.Y(n_3517)
);

HB1xp67_ASAP7_75t_L g3518 ( 
.A(n_3403),
.Y(n_3518)
);

AOI22xp33_ASAP7_75t_L g3519 ( 
.A1(n_3379),
.A2(n_3276),
.B1(n_3402),
.B2(n_3442),
.Y(n_3519)
);

OAI22xp5_ASAP7_75t_L g3520 ( 
.A1(n_3408),
.A2(n_3301),
.B1(n_3321),
.B2(n_3276),
.Y(n_3520)
);

OAI22xp5_ASAP7_75t_L g3521 ( 
.A1(n_3408),
.A2(n_3301),
.B1(n_3321),
.B2(n_3276),
.Y(n_3521)
);

AOI22xp33_ASAP7_75t_L g3522 ( 
.A1(n_3402),
.A2(n_3276),
.B1(n_3442),
.B2(n_3301),
.Y(n_3522)
);

HB1xp67_ASAP7_75t_L g3523 ( 
.A(n_3387),
.Y(n_3523)
);

AOI22xp5_ASAP7_75t_L g3524 ( 
.A1(n_3442),
.A2(n_3276),
.B1(n_3301),
.B2(n_3289),
.Y(n_3524)
);

AOI22xp33_ASAP7_75t_L g3525 ( 
.A1(n_3402),
.A2(n_3276),
.B1(n_3442),
.B2(n_3301),
.Y(n_3525)
);

AOI22xp33_ASAP7_75t_L g3526 ( 
.A1(n_3402),
.A2(n_3276),
.B1(n_3442),
.B2(n_3301),
.Y(n_3526)
);

AOI22xp5_ASAP7_75t_L g3527 ( 
.A1(n_3442),
.A2(n_3276),
.B1(n_3301),
.B2(n_3289),
.Y(n_3527)
);

OAI21xp5_ASAP7_75t_SL g3528 ( 
.A1(n_3402),
.A2(n_3276),
.B(n_3442),
.Y(n_3528)
);

OAI22xp5_ASAP7_75t_L g3529 ( 
.A1(n_3408),
.A2(n_3301),
.B1(n_3321),
.B2(n_3276),
.Y(n_3529)
);

OAI22xp5_ASAP7_75t_L g3530 ( 
.A1(n_3408),
.A2(n_3301),
.B1(n_3321),
.B2(n_3276),
.Y(n_3530)
);

AOI22xp5_ASAP7_75t_L g3531 ( 
.A1(n_3442),
.A2(n_3276),
.B1(n_3301),
.B2(n_3289),
.Y(n_3531)
);

AND2x2_ASAP7_75t_L g3532 ( 
.A(n_3383),
.B(n_3378),
.Y(n_3532)
);

OAI22xp5_ASAP7_75t_L g3533 ( 
.A1(n_3408),
.A2(n_3301),
.B1(n_3321),
.B2(n_3276),
.Y(n_3533)
);

OAI22xp5_ASAP7_75t_L g3534 ( 
.A1(n_3408),
.A2(n_3301),
.B1(n_3321),
.B2(n_3276),
.Y(n_3534)
);

AND2x4_ASAP7_75t_L g3535 ( 
.A(n_3472),
.B(n_3482),
.Y(n_3535)
);

AOI21x1_ASAP7_75t_L g3536 ( 
.A1(n_3481),
.A2(n_3462),
.B(n_3523),
.Y(n_3536)
);

HB1xp67_ASAP7_75t_L g3537 ( 
.A(n_3482),
.Y(n_3537)
);

INVx3_ASAP7_75t_L g3538 ( 
.A(n_3484),
.Y(n_3538)
);

AND2x2_ASAP7_75t_L g3539 ( 
.A(n_3487),
.B(n_3496),
.Y(n_3539)
);

NAND2xp5_ASAP7_75t_L g3540 ( 
.A(n_3519),
.B(n_3488),
.Y(n_3540)
);

AND2x4_ASAP7_75t_L g3541 ( 
.A(n_3523),
.B(n_3505),
.Y(n_3541)
);

INVx2_ASAP7_75t_L g3542 ( 
.A(n_3518),
.Y(n_3542)
);

BUFx3_ASAP7_75t_L g3543 ( 
.A(n_3498),
.Y(n_3543)
);

AO21x2_ASAP7_75t_L g3544 ( 
.A1(n_3494),
.A2(n_3517),
.B(n_3513),
.Y(n_3544)
);

AO21x2_ASAP7_75t_L g3545 ( 
.A1(n_3517),
.A2(n_3512),
.B(n_3495),
.Y(n_3545)
);

AND2x2_ASAP7_75t_L g3546 ( 
.A(n_3500),
.B(n_3532),
.Y(n_3546)
);

INVx3_ASAP7_75t_L g3547 ( 
.A(n_3460),
.Y(n_3547)
);

AND2x2_ASAP7_75t_L g3548 ( 
.A(n_3473),
.B(n_3471),
.Y(n_3548)
);

NAND2xp5_ASAP7_75t_L g3549 ( 
.A(n_3519),
.B(n_3522),
.Y(n_3549)
);

HB1xp67_ASAP7_75t_L g3550 ( 
.A(n_3504),
.Y(n_3550)
);

AND2x2_ASAP7_75t_L g3551 ( 
.A(n_3492),
.B(n_3514),
.Y(n_3551)
);

BUFx3_ASAP7_75t_L g3552 ( 
.A(n_3498),
.Y(n_3552)
);

INVx1_ASAP7_75t_SL g3553 ( 
.A(n_3480),
.Y(n_3553)
);

AO21x2_ASAP7_75t_L g3554 ( 
.A1(n_3507),
.A2(n_3467),
.B(n_3457),
.Y(n_3554)
);

AO21x2_ASAP7_75t_L g3555 ( 
.A1(n_3486),
.A2(n_3489),
.B(n_3477),
.Y(n_3555)
);

BUFx2_ASAP7_75t_SL g3556 ( 
.A(n_3460),
.Y(n_3556)
);

AND2x4_ASAP7_75t_L g3557 ( 
.A(n_3501),
.B(n_3493),
.Y(n_3557)
);

INVx2_ASAP7_75t_L g3558 ( 
.A(n_3515),
.Y(n_3558)
);

INVx2_ASAP7_75t_L g3559 ( 
.A(n_3476),
.Y(n_3559)
);

AO21x2_ASAP7_75t_L g3560 ( 
.A1(n_3524),
.A2(n_3531),
.B(n_3527),
.Y(n_3560)
);

INVx1_ASAP7_75t_L g3561 ( 
.A(n_3490),
.Y(n_3561)
);

NOR2xp33_ASAP7_75t_L g3562 ( 
.A(n_3466),
.B(n_3474),
.Y(n_3562)
);

AND2x2_ASAP7_75t_L g3563 ( 
.A(n_3502),
.B(n_3506),
.Y(n_3563)
);

AND2x2_ASAP7_75t_L g3564 ( 
.A(n_3506),
.B(n_3470),
.Y(n_3564)
);

INVx2_ASAP7_75t_L g3565 ( 
.A(n_3476),
.Y(n_3565)
);

INVx2_ASAP7_75t_L g3566 ( 
.A(n_3485),
.Y(n_3566)
);

INVx1_ASAP7_75t_L g3567 ( 
.A(n_3511),
.Y(n_3567)
);

HB1xp67_ASAP7_75t_L g3568 ( 
.A(n_3534),
.Y(n_3568)
);

AND2x2_ASAP7_75t_L g3569 ( 
.A(n_3509),
.B(n_3510),
.Y(n_3569)
);

OR2x2_ASAP7_75t_L g3570 ( 
.A(n_3464),
.B(n_3468),
.Y(n_3570)
);

INVx2_ASAP7_75t_SL g3571 ( 
.A(n_3469),
.Y(n_3571)
);

OR2x6_ASAP7_75t_L g3572 ( 
.A(n_3475),
.B(n_3459),
.Y(n_3572)
);

INVx2_ASAP7_75t_L g3573 ( 
.A(n_3508),
.Y(n_3573)
);

INVx2_ASAP7_75t_L g3574 ( 
.A(n_3508),
.Y(n_3574)
);

AND2x2_ASAP7_75t_L g3575 ( 
.A(n_3499),
.B(n_3491),
.Y(n_3575)
);

INVx2_ASAP7_75t_L g3576 ( 
.A(n_3503),
.Y(n_3576)
);

NAND2xp5_ASAP7_75t_L g3577 ( 
.A(n_3522),
.B(n_3526),
.Y(n_3577)
);

INVx1_ASAP7_75t_L g3578 ( 
.A(n_3520),
.Y(n_3578)
);

HB1xp67_ASAP7_75t_L g3579 ( 
.A(n_3521),
.Y(n_3579)
);

OR2x2_ASAP7_75t_L g3580 ( 
.A(n_3483),
.B(n_3516),
.Y(n_3580)
);

OA21x2_ASAP7_75t_L g3581 ( 
.A1(n_3463),
.A2(n_3526),
.B(n_3525),
.Y(n_3581)
);

HB1xp67_ASAP7_75t_L g3582 ( 
.A(n_3529),
.Y(n_3582)
);

AND2x2_ASAP7_75t_L g3583 ( 
.A(n_3497),
.B(n_3516),
.Y(n_3583)
);

INVx1_ASAP7_75t_L g3584 ( 
.A(n_3530),
.Y(n_3584)
);

AND2x2_ASAP7_75t_L g3585 ( 
.A(n_3525),
.B(n_3465),
.Y(n_3585)
);

INVx2_ASAP7_75t_L g3586 ( 
.A(n_3533),
.Y(n_3586)
);

BUFx2_ASAP7_75t_SL g3587 ( 
.A(n_3478),
.Y(n_3587)
);

BUFx2_ASAP7_75t_L g3588 ( 
.A(n_3479),
.Y(n_3588)
);

INVx2_ASAP7_75t_L g3589 ( 
.A(n_3465),
.Y(n_3589)
);

INVx1_ASAP7_75t_L g3590 ( 
.A(n_3458),
.Y(n_3590)
);

AND2x2_ASAP7_75t_L g3591 ( 
.A(n_3461),
.B(n_3458),
.Y(n_3591)
);

INVx1_ASAP7_75t_L g3592 ( 
.A(n_3482),
.Y(n_3592)
);

AND2x2_ASAP7_75t_L g3593 ( 
.A(n_3462),
.B(n_3487),
.Y(n_3593)
);

NOR2xp33_ASAP7_75t_L g3594 ( 
.A(n_3498),
.B(n_3466),
.Y(n_3594)
);

OA21x2_ASAP7_75t_L g3595 ( 
.A1(n_3501),
.A2(n_3493),
.B(n_3495),
.Y(n_3595)
);

INVx1_ASAP7_75t_L g3596 ( 
.A(n_3482),
.Y(n_3596)
);

AND2x4_ASAP7_75t_L g3597 ( 
.A(n_3472),
.B(n_3482),
.Y(n_3597)
);

INVx1_ASAP7_75t_L g3598 ( 
.A(n_3482),
.Y(n_3598)
);

OAI21xp5_ASAP7_75t_L g3599 ( 
.A1(n_3528),
.A2(n_3525),
.B(n_3522),
.Y(n_3599)
);

INVx1_ASAP7_75t_L g3600 ( 
.A(n_3482),
.Y(n_3600)
);

INVx2_ASAP7_75t_L g3601 ( 
.A(n_3482),
.Y(n_3601)
);

AOI21xp5_ASAP7_75t_L g3602 ( 
.A1(n_3528),
.A2(n_3525),
.B(n_3522),
.Y(n_3602)
);

AO21x2_ASAP7_75t_L g3603 ( 
.A1(n_3494),
.A2(n_3517),
.B(n_3513),
.Y(n_3603)
);

INVxp67_ASAP7_75t_L g3604 ( 
.A(n_3462),
.Y(n_3604)
);

NAND2xp5_ASAP7_75t_L g3605 ( 
.A(n_3519),
.B(n_3401),
.Y(n_3605)
);

INVx1_ASAP7_75t_L g3606 ( 
.A(n_3482),
.Y(n_3606)
);

INVx1_ASAP7_75t_L g3607 ( 
.A(n_3482),
.Y(n_3607)
);

AO21x2_ASAP7_75t_L g3608 ( 
.A1(n_3494),
.A2(n_3517),
.B(n_3513),
.Y(n_3608)
);

AO21x2_ASAP7_75t_L g3609 ( 
.A1(n_3494),
.A2(n_3517),
.B(n_3513),
.Y(n_3609)
);

AO21x2_ASAP7_75t_L g3610 ( 
.A1(n_3494),
.A2(n_3517),
.B(n_3513),
.Y(n_3610)
);

INVx2_ASAP7_75t_L g3611 ( 
.A(n_3482),
.Y(n_3611)
);

INVx1_ASAP7_75t_L g3612 ( 
.A(n_3482),
.Y(n_3612)
);

AO21x2_ASAP7_75t_L g3613 ( 
.A1(n_3494),
.A2(n_3517),
.B(n_3513),
.Y(n_3613)
);

INVx3_ASAP7_75t_L g3614 ( 
.A(n_3613),
.Y(n_3614)
);

INVx1_ASAP7_75t_L g3615 ( 
.A(n_3537),
.Y(n_3615)
);

INVx1_ASAP7_75t_L g3616 ( 
.A(n_3601),
.Y(n_3616)
);

INVx1_ASAP7_75t_L g3617 ( 
.A(n_3601),
.Y(n_3617)
);

INVx1_ASAP7_75t_L g3618 ( 
.A(n_3601),
.Y(n_3618)
);

INVx1_ASAP7_75t_SL g3619 ( 
.A(n_3587),
.Y(n_3619)
);

AOI22xp33_ASAP7_75t_SL g3620 ( 
.A1(n_3591),
.A2(n_3575),
.B1(n_3585),
.B2(n_3563),
.Y(n_3620)
);

INVx2_ASAP7_75t_L g3621 ( 
.A(n_3544),
.Y(n_3621)
);

INVx1_ASAP7_75t_L g3622 ( 
.A(n_3611),
.Y(n_3622)
);

AND2x2_ASAP7_75t_L g3623 ( 
.A(n_3593),
.B(n_3548),
.Y(n_3623)
);

OR2x2_ASAP7_75t_L g3624 ( 
.A(n_3604),
.B(n_3592),
.Y(n_3624)
);

INVx1_ASAP7_75t_L g3625 ( 
.A(n_3542),
.Y(n_3625)
);

INVx2_ASAP7_75t_L g3626 ( 
.A(n_3544),
.Y(n_3626)
);

HB1xp67_ASAP7_75t_L g3627 ( 
.A(n_3604),
.Y(n_3627)
);

INVx2_ASAP7_75t_L g3628 ( 
.A(n_3544),
.Y(n_3628)
);

AND2x2_ASAP7_75t_L g3629 ( 
.A(n_3593),
.B(n_3548),
.Y(n_3629)
);

INVx1_ASAP7_75t_L g3630 ( 
.A(n_3542),
.Y(n_3630)
);

NAND3xp33_ASAP7_75t_L g3631 ( 
.A(n_3599),
.B(n_3602),
.C(n_3540),
.Y(n_3631)
);

OA222x2_ASAP7_75t_L g3632 ( 
.A1(n_3580),
.A2(n_3561),
.B1(n_3572),
.B2(n_3605),
.C1(n_3570),
.C2(n_3540),
.Y(n_3632)
);

AO31x2_ASAP7_75t_L g3633 ( 
.A1(n_3561),
.A2(n_3605),
.A3(n_3549),
.B(n_3577),
.Y(n_3633)
);

AND2x2_ASAP7_75t_L g3634 ( 
.A(n_3539),
.B(n_3546),
.Y(n_3634)
);

INVx2_ASAP7_75t_SL g3635 ( 
.A(n_3547),
.Y(n_3635)
);

AND2x2_ASAP7_75t_L g3636 ( 
.A(n_3539),
.B(n_3546),
.Y(n_3636)
);

INVx1_ASAP7_75t_L g3637 ( 
.A(n_3542),
.Y(n_3637)
);

NOR2x1_ASAP7_75t_L g3638 ( 
.A(n_3544),
.B(n_3603),
.Y(n_3638)
);

AND2x2_ASAP7_75t_L g3639 ( 
.A(n_3551),
.B(n_3566),
.Y(n_3639)
);

AND2x2_ASAP7_75t_L g3640 ( 
.A(n_3551),
.B(n_3566),
.Y(n_3640)
);

INVx1_ASAP7_75t_L g3641 ( 
.A(n_3592),
.Y(n_3641)
);

AND2x2_ASAP7_75t_L g3642 ( 
.A(n_3566),
.B(n_3564),
.Y(n_3642)
);

BUFx2_ASAP7_75t_L g3643 ( 
.A(n_3547),
.Y(n_3643)
);

INVx2_ASAP7_75t_L g3644 ( 
.A(n_3603),
.Y(n_3644)
);

NAND2xp5_ASAP7_75t_L g3645 ( 
.A(n_3591),
.B(n_3585),
.Y(n_3645)
);

HB1xp67_ASAP7_75t_L g3646 ( 
.A(n_3535),
.Y(n_3646)
);

AND2x4_ASAP7_75t_L g3647 ( 
.A(n_3535),
.B(n_3597),
.Y(n_3647)
);

AND2x2_ASAP7_75t_L g3648 ( 
.A(n_3564),
.B(n_3573),
.Y(n_3648)
);

OR2x2_ASAP7_75t_L g3649 ( 
.A(n_3596),
.B(n_3598),
.Y(n_3649)
);

AND2x2_ASAP7_75t_L g3650 ( 
.A(n_3573),
.B(n_3574),
.Y(n_3650)
);

INVx2_ASAP7_75t_L g3651 ( 
.A(n_3603),
.Y(n_3651)
);

INVx3_ASAP7_75t_L g3652 ( 
.A(n_3613),
.Y(n_3652)
);

BUFx4f_ASAP7_75t_L g3653 ( 
.A(n_3538),
.Y(n_3653)
);

INVx2_ASAP7_75t_L g3654 ( 
.A(n_3603),
.Y(n_3654)
);

AND2x2_ASAP7_75t_L g3655 ( 
.A(n_3573),
.B(n_3574),
.Y(n_3655)
);

OR2x2_ASAP7_75t_L g3656 ( 
.A(n_3600),
.B(n_3606),
.Y(n_3656)
);

NAND2xp5_ASAP7_75t_L g3657 ( 
.A(n_3602),
.B(n_3568),
.Y(n_3657)
);

INVx2_ASAP7_75t_SL g3658 ( 
.A(n_3547),
.Y(n_3658)
);

OAI33xp33_ASAP7_75t_L g3659 ( 
.A1(n_3549),
.A2(n_3577),
.A3(n_3584),
.B1(n_3578),
.B2(n_3570),
.B3(n_3590),
.Y(n_3659)
);

AND2x4_ASAP7_75t_L g3660 ( 
.A(n_3535),
.B(n_3597),
.Y(n_3660)
);

INVx2_ASAP7_75t_L g3661 ( 
.A(n_3608),
.Y(n_3661)
);

NAND2xp5_ASAP7_75t_L g3662 ( 
.A(n_3568),
.B(n_3579),
.Y(n_3662)
);

INVx2_ASAP7_75t_L g3663 ( 
.A(n_3608),
.Y(n_3663)
);

INVx2_ASAP7_75t_L g3664 ( 
.A(n_3608),
.Y(n_3664)
);

INVxp33_ASAP7_75t_L g3665 ( 
.A(n_3562),
.Y(n_3665)
);

AND2x2_ASAP7_75t_L g3666 ( 
.A(n_3574),
.B(n_3569),
.Y(n_3666)
);

AND2x4_ASAP7_75t_SL g3667 ( 
.A(n_3547),
.B(n_3576),
.Y(n_3667)
);

INVx1_ASAP7_75t_SL g3668 ( 
.A(n_3587),
.Y(n_3668)
);

HB1xp67_ASAP7_75t_L g3669 ( 
.A(n_3535),
.Y(n_3669)
);

AND2x2_ASAP7_75t_L g3670 ( 
.A(n_3569),
.B(n_3541),
.Y(n_3670)
);

AND2x2_ASAP7_75t_L g3671 ( 
.A(n_3541),
.B(n_3576),
.Y(n_3671)
);

AND2x2_ASAP7_75t_L g3672 ( 
.A(n_3541),
.B(n_3576),
.Y(n_3672)
);

HB1xp67_ASAP7_75t_L g3673 ( 
.A(n_3597),
.Y(n_3673)
);

BUFx6f_ASAP7_75t_L g3674 ( 
.A(n_3543),
.Y(n_3674)
);

AND2x4_ASAP7_75t_L g3675 ( 
.A(n_3597),
.B(n_3559),
.Y(n_3675)
);

INVx2_ASAP7_75t_L g3676 ( 
.A(n_3608),
.Y(n_3676)
);

AO21x2_ASAP7_75t_L g3677 ( 
.A1(n_3613),
.A2(n_3610),
.B(n_3609),
.Y(n_3677)
);

OAI221xp5_ASAP7_75t_L g3678 ( 
.A1(n_3599),
.A2(n_3572),
.B1(n_3581),
.B2(n_3582),
.C(n_3590),
.Y(n_3678)
);

AND2x2_ASAP7_75t_L g3679 ( 
.A(n_3541),
.B(n_3536),
.Y(n_3679)
);

OR2x2_ASAP7_75t_L g3680 ( 
.A(n_3607),
.B(n_3612),
.Y(n_3680)
);

INVx2_ASAP7_75t_L g3681 ( 
.A(n_3609),
.Y(n_3681)
);

INVx2_ASAP7_75t_L g3682 ( 
.A(n_3609),
.Y(n_3682)
);

BUFx2_ASAP7_75t_L g3683 ( 
.A(n_3609),
.Y(n_3683)
);

OAI211xp5_ASAP7_75t_SL g3684 ( 
.A1(n_3578),
.A2(n_3584),
.B(n_3586),
.C(n_3589),
.Y(n_3684)
);

AOI22xp33_ASAP7_75t_L g3685 ( 
.A1(n_3581),
.A2(n_3572),
.B1(n_3560),
.B2(n_3589),
.Y(n_3685)
);

INVx2_ASAP7_75t_L g3686 ( 
.A(n_3610),
.Y(n_3686)
);

INVx2_ASAP7_75t_L g3687 ( 
.A(n_3610),
.Y(n_3687)
);

INVx2_ASAP7_75t_L g3688 ( 
.A(n_3610),
.Y(n_3688)
);

INVx1_ASAP7_75t_L g3689 ( 
.A(n_3550),
.Y(n_3689)
);

INVx1_ASAP7_75t_L g3690 ( 
.A(n_3550),
.Y(n_3690)
);

OR2x6_ASAP7_75t_L g3691 ( 
.A(n_3556),
.B(n_3543),
.Y(n_3691)
);

HB1xp67_ASAP7_75t_L g3692 ( 
.A(n_3558),
.Y(n_3692)
);

AND2x2_ASAP7_75t_L g3693 ( 
.A(n_3536),
.B(n_3558),
.Y(n_3693)
);

AND2x2_ASAP7_75t_L g3694 ( 
.A(n_3623),
.B(n_3629),
.Y(n_3694)
);

INVx4_ASAP7_75t_L g3695 ( 
.A(n_3674),
.Y(n_3695)
);

AND2x2_ASAP7_75t_L g3696 ( 
.A(n_3623),
.B(n_3559),
.Y(n_3696)
);

INVx1_ASAP7_75t_L g3697 ( 
.A(n_3683),
.Y(n_3697)
);

INVx2_ASAP7_75t_L g3698 ( 
.A(n_3677),
.Y(n_3698)
);

INVx1_ASAP7_75t_L g3699 ( 
.A(n_3683),
.Y(n_3699)
);

OR2x2_ASAP7_75t_L g3700 ( 
.A(n_3677),
.B(n_3589),
.Y(n_3700)
);

AOI22xp33_ASAP7_75t_L g3701 ( 
.A1(n_3631),
.A2(n_3572),
.B1(n_3581),
.B2(n_3560),
.Y(n_3701)
);

NAND2xp5_ASAP7_75t_L g3702 ( 
.A(n_3629),
.B(n_3571),
.Y(n_3702)
);

AND2x2_ASAP7_75t_L g3703 ( 
.A(n_3634),
.B(n_3559),
.Y(n_3703)
);

INVx1_ASAP7_75t_L g3704 ( 
.A(n_3638),
.Y(n_3704)
);

NAND2xp5_ASAP7_75t_L g3705 ( 
.A(n_3620),
.B(n_3642),
.Y(n_3705)
);

INVx1_ASAP7_75t_L g3706 ( 
.A(n_3689),
.Y(n_3706)
);

INVx1_ASAP7_75t_L g3707 ( 
.A(n_3689),
.Y(n_3707)
);

INVx1_ASAP7_75t_L g3708 ( 
.A(n_3690),
.Y(n_3708)
);

INVx1_ASAP7_75t_L g3709 ( 
.A(n_3690),
.Y(n_3709)
);

AND2x2_ASAP7_75t_L g3710 ( 
.A(n_3634),
.B(n_3565),
.Y(n_3710)
);

INVx3_ASAP7_75t_L g3711 ( 
.A(n_3677),
.Y(n_3711)
);

INVx1_ASAP7_75t_L g3712 ( 
.A(n_3627),
.Y(n_3712)
);

INVx1_ASAP7_75t_L g3713 ( 
.A(n_3646),
.Y(n_3713)
);

INVx2_ASAP7_75t_L g3714 ( 
.A(n_3647),
.Y(n_3714)
);

OR2x2_ASAP7_75t_L g3715 ( 
.A(n_3624),
.B(n_3692),
.Y(n_3715)
);

HB1xp67_ASAP7_75t_L g3716 ( 
.A(n_3669),
.Y(n_3716)
);

AND2x2_ASAP7_75t_L g3717 ( 
.A(n_3636),
.B(n_3565),
.Y(n_3717)
);

AND2x2_ASAP7_75t_L g3718 ( 
.A(n_3636),
.B(n_3565),
.Y(n_3718)
);

AND2x2_ASAP7_75t_L g3719 ( 
.A(n_3639),
.B(n_3556),
.Y(n_3719)
);

BUFx2_ASAP7_75t_L g3720 ( 
.A(n_3614),
.Y(n_3720)
);

AND2x2_ASAP7_75t_L g3721 ( 
.A(n_3639),
.B(n_3571),
.Y(n_3721)
);

AND2x2_ASAP7_75t_L g3722 ( 
.A(n_3640),
.B(n_3571),
.Y(n_3722)
);

INVx1_ASAP7_75t_L g3723 ( 
.A(n_3673),
.Y(n_3723)
);

INVx2_ASAP7_75t_L g3724 ( 
.A(n_3647),
.Y(n_3724)
);

INVx1_ASAP7_75t_L g3725 ( 
.A(n_3649),
.Y(n_3725)
);

AND2x2_ASAP7_75t_L g3726 ( 
.A(n_3640),
.B(n_3552),
.Y(n_3726)
);

BUFx6f_ASAP7_75t_L g3727 ( 
.A(n_3674),
.Y(n_3727)
);

INVx1_ASAP7_75t_L g3728 ( 
.A(n_3649),
.Y(n_3728)
);

OR2x2_ASAP7_75t_L g3729 ( 
.A(n_3624),
.B(n_3586),
.Y(n_3729)
);

INVx2_ASAP7_75t_L g3730 ( 
.A(n_3647),
.Y(n_3730)
);

OR2x2_ASAP7_75t_L g3731 ( 
.A(n_3614),
.B(n_3586),
.Y(n_3731)
);

AND2x2_ASAP7_75t_L g3732 ( 
.A(n_3667),
.B(n_3552),
.Y(n_3732)
);

NAND2xp5_ASAP7_75t_L g3733 ( 
.A(n_3642),
.B(n_3648),
.Y(n_3733)
);

BUFx3_ASAP7_75t_L g3734 ( 
.A(n_3643),
.Y(n_3734)
);

BUFx3_ASAP7_75t_L g3735 ( 
.A(n_3643),
.Y(n_3735)
);

INVx1_ASAP7_75t_L g3736 ( 
.A(n_3656),
.Y(n_3736)
);

OAI211xp5_ASAP7_75t_L g3737 ( 
.A1(n_3685),
.A2(n_3563),
.B(n_3581),
.C(n_3583),
.Y(n_3737)
);

INVx1_ASAP7_75t_L g3738 ( 
.A(n_3656),
.Y(n_3738)
);

INVx2_ASAP7_75t_L g3739 ( 
.A(n_3614),
.Y(n_3739)
);

BUFx6f_ASAP7_75t_L g3740 ( 
.A(n_3674),
.Y(n_3740)
);

OR2x2_ASAP7_75t_L g3741 ( 
.A(n_3652),
.B(n_3567),
.Y(n_3741)
);

INVx1_ASAP7_75t_L g3742 ( 
.A(n_3680),
.Y(n_3742)
);

INVx1_ASAP7_75t_L g3743 ( 
.A(n_3680),
.Y(n_3743)
);

OR2x2_ASAP7_75t_L g3744 ( 
.A(n_3652),
.B(n_3613),
.Y(n_3744)
);

INVx1_ASAP7_75t_L g3745 ( 
.A(n_3652),
.Y(n_3745)
);

INVx2_ASAP7_75t_L g3746 ( 
.A(n_3621),
.Y(n_3746)
);

NOR2xp33_ASAP7_75t_L g3747 ( 
.A(n_3665),
.B(n_3553),
.Y(n_3747)
);

NAND3xp33_ASAP7_75t_L g3748 ( 
.A(n_3701),
.B(n_3678),
.C(n_3657),
.Y(n_3748)
);

INVx2_ASAP7_75t_L g3749 ( 
.A(n_3711),
.Y(n_3749)
);

INVx2_ASAP7_75t_L g3750 ( 
.A(n_3711),
.Y(n_3750)
);

AND2x4_ASAP7_75t_SL g3751 ( 
.A(n_3727),
.B(n_3691),
.Y(n_3751)
);

BUFx3_ASAP7_75t_L g3752 ( 
.A(n_3720),
.Y(n_3752)
);

AND2x2_ASAP7_75t_L g3753 ( 
.A(n_3719),
.B(n_3632),
.Y(n_3753)
);

AND2x4_ASAP7_75t_L g3754 ( 
.A(n_3734),
.B(n_3660),
.Y(n_3754)
);

INVx2_ASAP7_75t_L g3755 ( 
.A(n_3711),
.Y(n_3755)
);

AND4x1_ASAP7_75t_L g3756 ( 
.A(n_3747),
.B(n_3659),
.C(n_3645),
.D(n_3594),
.Y(n_3756)
);

AND2x2_ASAP7_75t_L g3757 ( 
.A(n_3719),
.B(n_3679),
.Y(n_3757)
);

NAND2xp5_ASAP7_75t_L g3758 ( 
.A(n_3737),
.B(n_3633),
.Y(n_3758)
);

OR2x2_ASAP7_75t_L g3759 ( 
.A(n_3711),
.B(n_3621),
.Y(n_3759)
);

NAND2xp5_ASAP7_75t_L g3760 ( 
.A(n_3734),
.B(n_3633),
.Y(n_3760)
);

AND2x2_ASAP7_75t_L g3761 ( 
.A(n_3721),
.B(n_3722),
.Y(n_3761)
);

AND2x2_ASAP7_75t_L g3762 ( 
.A(n_3721),
.B(n_3679),
.Y(n_3762)
);

INVx1_ASAP7_75t_L g3763 ( 
.A(n_3720),
.Y(n_3763)
);

AND2x2_ASAP7_75t_L g3764 ( 
.A(n_3722),
.B(n_3691),
.Y(n_3764)
);

BUFx3_ASAP7_75t_L g3765 ( 
.A(n_3734),
.Y(n_3765)
);

NAND2xp5_ASAP7_75t_L g3766 ( 
.A(n_3735),
.B(n_3633),
.Y(n_3766)
);

INVx2_ASAP7_75t_L g3767 ( 
.A(n_3698),
.Y(n_3767)
);

AND2x2_ASAP7_75t_L g3768 ( 
.A(n_3726),
.B(n_3691),
.Y(n_3768)
);

NAND2xp5_ASAP7_75t_L g3769 ( 
.A(n_3735),
.B(n_3633),
.Y(n_3769)
);

INVx1_ASAP7_75t_L g3770 ( 
.A(n_3698),
.Y(n_3770)
);

INVx2_ASAP7_75t_L g3771 ( 
.A(n_3698),
.Y(n_3771)
);

INVx1_ASAP7_75t_L g3772 ( 
.A(n_3735),
.Y(n_3772)
);

AND2x4_ASAP7_75t_L g3773 ( 
.A(n_3695),
.B(n_3660),
.Y(n_3773)
);

AND2x4_ASAP7_75t_L g3774 ( 
.A(n_3695),
.B(n_3660),
.Y(n_3774)
);

NOR2xp33_ASAP7_75t_L g3775 ( 
.A(n_3705),
.B(n_3619),
.Y(n_3775)
);

NAND2xp5_ASAP7_75t_L g3776 ( 
.A(n_3716),
.B(n_3633),
.Y(n_3776)
);

BUFx3_ASAP7_75t_L g3777 ( 
.A(n_3704),
.Y(n_3777)
);

AND2x2_ASAP7_75t_L g3778 ( 
.A(n_3726),
.B(n_3694),
.Y(n_3778)
);

NAND2xp5_ASAP7_75t_L g3779 ( 
.A(n_3694),
.B(n_3581),
.Y(n_3779)
);

INVx1_ASAP7_75t_L g3780 ( 
.A(n_3715),
.Y(n_3780)
);

INVx2_ASAP7_75t_SL g3781 ( 
.A(n_3727),
.Y(n_3781)
);

NOR2xp33_ASAP7_75t_L g3782 ( 
.A(n_3733),
.B(n_3668),
.Y(n_3782)
);

INVx1_ASAP7_75t_L g3783 ( 
.A(n_3715),
.Y(n_3783)
);

NAND2xp5_ASAP7_75t_SL g3784 ( 
.A(n_3700),
.B(n_3557),
.Y(n_3784)
);

NAND2xp5_ASAP7_75t_L g3785 ( 
.A(n_3712),
.B(n_3713),
.Y(n_3785)
);

AND2x2_ASAP7_75t_L g3786 ( 
.A(n_3732),
.B(n_3691),
.Y(n_3786)
);

HB1xp67_ASAP7_75t_L g3787 ( 
.A(n_3704),
.Y(n_3787)
);

OA21x2_ASAP7_75t_L g3788 ( 
.A1(n_3744),
.A2(n_3664),
.B(n_3686),
.Y(n_3788)
);

AND2x2_ASAP7_75t_L g3789 ( 
.A(n_3732),
.B(n_3545),
.Y(n_3789)
);

OAI221xp5_ASAP7_75t_SL g3790 ( 
.A1(n_3700),
.A2(n_3572),
.B1(n_3580),
.B2(n_3583),
.C(n_3575),
.Y(n_3790)
);

INVx1_ASAP7_75t_L g3791 ( 
.A(n_3739),
.Y(n_3791)
);

INVx2_ASAP7_75t_L g3792 ( 
.A(n_3744),
.Y(n_3792)
);

INVx2_ASAP7_75t_L g3793 ( 
.A(n_3697),
.Y(n_3793)
);

INVx2_ASAP7_75t_L g3794 ( 
.A(n_3697),
.Y(n_3794)
);

INVx2_ASAP7_75t_L g3795 ( 
.A(n_3699),
.Y(n_3795)
);

INVx2_ASAP7_75t_L g3796 ( 
.A(n_3699),
.Y(n_3796)
);

AND2x2_ASAP7_75t_L g3797 ( 
.A(n_3696),
.B(n_3545),
.Y(n_3797)
);

AND2x2_ASAP7_75t_L g3798 ( 
.A(n_3696),
.B(n_3703),
.Y(n_3798)
);

AND2x4_ASAP7_75t_L g3799 ( 
.A(n_3695),
.B(n_3635),
.Y(n_3799)
);

INVx1_ASAP7_75t_SL g3800 ( 
.A(n_3753),
.Y(n_3800)
);

INVx2_ASAP7_75t_L g3801 ( 
.A(n_3752),
.Y(n_3801)
);

INVx1_ASAP7_75t_L g3802 ( 
.A(n_3752),
.Y(n_3802)
);

HB1xp67_ASAP7_75t_L g3803 ( 
.A(n_3765),
.Y(n_3803)
);

AND2x2_ASAP7_75t_L g3804 ( 
.A(n_3798),
.B(n_3703),
.Y(n_3804)
);

INVx1_ASAP7_75t_L g3805 ( 
.A(n_3752),
.Y(n_3805)
);

OR2x2_ASAP7_75t_L g3806 ( 
.A(n_3758),
.B(n_3626),
.Y(n_3806)
);

NOR2xp33_ASAP7_75t_SL g3807 ( 
.A(n_3790),
.B(n_3543),
.Y(n_3807)
);

INVx1_ASAP7_75t_L g3808 ( 
.A(n_3752),
.Y(n_3808)
);

INVx2_ASAP7_75t_L g3809 ( 
.A(n_3765),
.Y(n_3809)
);

OR2x2_ASAP7_75t_L g3810 ( 
.A(n_3758),
.B(n_3626),
.Y(n_3810)
);

INVx2_ASAP7_75t_L g3811 ( 
.A(n_3765),
.Y(n_3811)
);

OR2x2_ASAP7_75t_L g3812 ( 
.A(n_3784),
.B(n_3628),
.Y(n_3812)
);

AND2x2_ASAP7_75t_L g3813 ( 
.A(n_3798),
.B(n_3710),
.Y(n_3813)
);

HB1xp67_ASAP7_75t_L g3814 ( 
.A(n_3765),
.Y(n_3814)
);

INVx2_ASAP7_75t_L g3815 ( 
.A(n_3788),
.Y(n_3815)
);

AND2x2_ASAP7_75t_L g3816 ( 
.A(n_3798),
.B(n_3710),
.Y(n_3816)
);

AND2x2_ASAP7_75t_L g3817 ( 
.A(n_3778),
.B(n_3717),
.Y(n_3817)
);

NOR2xp33_ASAP7_75t_L g3818 ( 
.A(n_3756),
.B(n_3538),
.Y(n_3818)
);

NOR2x1_ASAP7_75t_L g3819 ( 
.A(n_3760),
.B(n_3695),
.Y(n_3819)
);

INVx1_ASAP7_75t_SL g3820 ( 
.A(n_3753),
.Y(n_3820)
);

INVx1_ASAP7_75t_L g3821 ( 
.A(n_3763),
.Y(n_3821)
);

INVx1_ASAP7_75t_L g3822 ( 
.A(n_3763),
.Y(n_3822)
);

INVx2_ASAP7_75t_L g3823 ( 
.A(n_3788),
.Y(n_3823)
);

NAND2xp5_ASAP7_75t_L g3824 ( 
.A(n_3756),
.B(n_3712),
.Y(n_3824)
);

AND2x2_ASAP7_75t_L g3825 ( 
.A(n_3778),
.B(n_3761),
.Y(n_3825)
);

INVx2_ASAP7_75t_L g3826 ( 
.A(n_3788),
.Y(n_3826)
);

INVx1_ASAP7_75t_L g3827 ( 
.A(n_3759),
.Y(n_3827)
);

INVx4_ASAP7_75t_L g3828 ( 
.A(n_3751),
.Y(n_3828)
);

INVx2_ASAP7_75t_L g3829 ( 
.A(n_3788),
.Y(n_3829)
);

INVx2_ASAP7_75t_L g3830 ( 
.A(n_3788),
.Y(n_3830)
);

NOR2xp33_ASAP7_75t_L g3831 ( 
.A(n_3790),
.B(n_3538),
.Y(n_3831)
);

AND2x2_ASAP7_75t_L g3832 ( 
.A(n_3778),
.B(n_3717),
.Y(n_3832)
);

INVx5_ASAP7_75t_L g3833 ( 
.A(n_3781),
.Y(n_3833)
);

INVx1_ASAP7_75t_L g3834 ( 
.A(n_3759),
.Y(n_3834)
);

INVx1_ASAP7_75t_L g3835 ( 
.A(n_3759),
.Y(n_3835)
);

INVx2_ASAP7_75t_SL g3836 ( 
.A(n_3751),
.Y(n_3836)
);

INVx2_ASAP7_75t_L g3837 ( 
.A(n_3788),
.Y(n_3837)
);

INVx4_ASAP7_75t_L g3838 ( 
.A(n_3751),
.Y(n_3838)
);

AND2x2_ASAP7_75t_L g3839 ( 
.A(n_3825),
.B(n_3761),
.Y(n_3839)
);

INVx1_ASAP7_75t_L g3840 ( 
.A(n_3814),
.Y(n_3840)
);

OR2x2_ASAP7_75t_L g3841 ( 
.A(n_3800),
.B(n_3779),
.Y(n_3841)
);

AND2x2_ASAP7_75t_L g3842 ( 
.A(n_3825),
.B(n_3761),
.Y(n_3842)
);

INVx1_ASAP7_75t_L g3843 ( 
.A(n_3814),
.Y(n_3843)
);

NAND2xp67_ASAP7_75t_L g3844 ( 
.A(n_3809),
.B(n_3751),
.Y(n_3844)
);

NAND2xp5_ASAP7_75t_L g3845 ( 
.A(n_3817),
.B(n_3753),
.Y(n_3845)
);

AND2x2_ASAP7_75t_L g3846 ( 
.A(n_3817),
.B(n_3762),
.Y(n_3846)
);

INVx1_ASAP7_75t_L g3847 ( 
.A(n_3803),
.Y(n_3847)
);

AND2x4_ASAP7_75t_L g3848 ( 
.A(n_3801),
.B(n_3754),
.Y(n_3848)
);

INVx1_ASAP7_75t_L g3849 ( 
.A(n_3801),
.Y(n_3849)
);

INVx1_ASAP7_75t_L g3850 ( 
.A(n_3801),
.Y(n_3850)
);

NAND2xp5_ASAP7_75t_L g3851 ( 
.A(n_3832),
.B(n_3718),
.Y(n_3851)
);

AND2x2_ASAP7_75t_L g3852 ( 
.A(n_3832),
.B(n_3762),
.Y(n_3852)
);

INVx1_ASAP7_75t_L g3853 ( 
.A(n_3804),
.Y(n_3853)
);

OR2x2_ASAP7_75t_L g3854 ( 
.A(n_3800),
.B(n_3820),
.Y(n_3854)
);

INVx1_ASAP7_75t_L g3855 ( 
.A(n_3804),
.Y(n_3855)
);

AND2x2_ASAP7_75t_L g3856 ( 
.A(n_3813),
.B(n_3762),
.Y(n_3856)
);

NAND2xp5_ASAP7_75t_L g3857 ( 
.A(n_3813),
.B(n_3718),
.Y(n_3857)
);

OR2x2_ASAP7_75t_L g3858 ( 
.A(n_3820),
.B(n_3779),
.Y(n_3858)
);

INVx2_ASAP7_75t_L g3859 ( 
.A(n_3833),
.Y(n_3859)
);

AND2x2_ASAP7_75t_L g3860 ( 
.A(n_3816),
.B(n_3757),
.Y(n_3860)
);

INVx1_ASAP7_75t_L g3861 ( 
.A(n_3816),
.Y(n_3861)
);

AND2x4_ASAP7_75t_L g3862 ( 
.A(n_3809),
.B(n_3754),
.Y(n_3862)
);

AND2x4_ASAP7_75t_L g3863 ( 
.A(n_3809),
.B(n_3754),
.Y(n_3863)
);

INVx1_ASAP7_75t_L g3864 ( 
.A(n_3802),
.Y(n_3864)
);

NOR2x1p5_ASAP7_75t_L g3865 ( 
.A(n_3851),
.B(n_3552),
.Y(n_3865)
);

NAND2xp5_ASAP7_75t_L g3866 ( 
.A(n_3839),
.B(n_3764),
.Y(n_3866)
);

INVx2_ASAP7_75t_L g3867 ( 
.A(n_3848),
.Y(n_3867)
);

NAND2xp5_ASAP7_75t_L g3868 ( 
.A(n_3839),
.B(n_3764),
.Y(n_3868)
);

INVx1_ASAP7_75t_L g3869 ( 
.A(n_3842),
.Y(n_3869)
);

NOR2x1_ASAP7_75t_L g3870 ( 
.A(n_3854),
.B(n_3838),
.Y(n_3870)
);

AND2x2_ASAP7_75t_L g3871 ( 
.A(n_3842),
.B(n_3768),
.Y(n_3871)
);

INVx1_ASAP7_75t_L g3872 ( 
.A(n_3860),
.Y(n_3872)
);

INVx2_ASAP7_75t_L g3873 ( 
.A(n_3848),
.Y(n_3873)
);

INVx2_ASAP7_75t_L g3874 ( 
.A(n_3848),
.Y(n_3874)
);

AND2x2_ASAP7_75t_L g3875 ( 
.A(n_3860),
.B(n_3768),
.Y(n_3875)
);

AND2x2_ASAP7_75t_L g3876 ( 
.A(n_3846),
.B(n_3768),
.Y(n_3876)
);

AND2x2_ASAP7_75t_L g3877 ( 
.A(n_3846),
.B(n_3764),
.Y(n_3877)
);

AND2x2_ASAP7_75t_L g3878 ( 
.A(n_3852),
.B(n_3786),
.Y(n_3878)
);

INVx2_ASAP7_75t_L g3879 ( 
.A(n_3862),
.Y(n_3879)
);

INVx2_ASAP7_75t_L g3880 ( 
.A(n_3862),
.Y(n_3880)
);

INVx1_ASAP7_75t_L g3881 ( 
.A(n_3862),
.Y(n_3881)
);

NAND2xp5_ASAP7_75t_L g3882 ( 
.A(n_3852),
.B(n_3757),
.Y(n_3882)
);

INVx1_ASAP7_75t_L g3883 ( 
.A(n_3863),
.Y(n_3883)
);

OR2x2_ASAP7_75t_L g3884 ( 
.A(n_3845),
.B(n_3729),
.Y(n_3884)
);

INVx1_ASAP7_75t_L g3885 ( 
.A(n_3867),
.Y(n_3885)
);

OR2x2_ASAP7_75t_L g3886 ( 
.A(n_3882),
.B(n_3841),
.Y(n_3886)
);

INVxp67_ASAP7_75t_SL g3887 ( 
.A(n_3870),
.Y(n_3887)
);

NOR2xp33_ASAP7_75t_SL g3888 ( 
.A(n_3878),
.B(n_3786),
.Y(n_3888)
);

NAND2x1p5_ASAP7_75t_L g3889 ( 
.A(n_3881),
.B(n_3828),
.Y(n_3889)
);

INVx1_ASAP7_75t_SL g3890 ( 
.A(n_3878),
.Y(n_3890)
);

AND2x2_ASAP7_75t_L g3891 ( 
.A(n_3875),
.B(n_3786),
.Y(n_3891)
);

INVx1_ASAP7_75t_L g3892 ( 
.A(n_3867),
.Y(n_3892)
);

NAND2xp5_ASAP7_75t_L g3893 ( 
.A(n_3871),
.B(n_3856),
.Y(n_3893)
);

INVx2_ASAP7_75t_L g3894 ( 
.A(n_3873),
.Y(n_3894)
);

AND2x2_ASAP7_75t_L g3895 ( 
.A(n_3871),
.B(n_3856),
.Y(n_3895)
);

AND2x2_ASAP7_75t_L g3896 ( 
.A(n_3875),
.B(n_3650),
.Y(n_3896)
);

OAI21xp5_ASAP7_75t_SL g3897 ( 
.A1(n_3876),
.A2(n_3748),
.B(n_3824),
.Y(n_3897)
);

AND2x2_ASAP7_75t_L g3898 ( 
.A(n_3876),
.B(n_3650),
.Y(n_3898)
);

AND2x2_ASAP7_75t_L g3899 ( 
.A(n_3877),
.B(n_3655),
.Y(n_3899)
);

INVx1_ASAP7_75t_L g3900 ( 
.A(n_3873),
.Y(n_3900)
);

HB1xp67_ASAP7_75t_L g3901 ( 
.A(n_3874),
.Y(n_3901)
);

NAND2xp5_ASAP7_75t_L g3902 ( 
.A(n_3895),
.B(n_3877),
.Y(n_3902)
);

NAND2xp5_ASAP7_75t_L g3903 ( 
.A(n_3895),
.B(n_3896),
.Y(n_3903)
);

INVx1_ASAP7_75t_L g3904 ( 
.A(n_3901),
.Y(n_3904)
);

INVx1_ASAP7_75t_L g3905 ( 
.A(n_3901),
.Y(n_3905)
);

AND2x2_ASAP7_75t_L g3906 ( 
.A(n_3891),
.B(n_3674),
.Y(n_3906)
);

AND2x4_ASAP7_75t_L g3907 ( 
.A(n_3896),
.B(n_3836),
.Y(n_3907)
);

NAND2x1_ASAP7_75t_L g3908 ( 
.A(n_3898),
.B(n_3754),
.Y(n_3908)
);

AOI21xp5_ASAP7_75t_L g3909 ( 
.A1(n_3897),
.A2(n_3824),
.B(n_3748),
.Y(n_3909)
);

AND2x2_ASAP7_75t_L g3910 ( 
.A(n_3898),
.B(n_3674),
.Y(n_3910)
);

OR2x2_ASAP7_75t_L g3911 ( 
.A(n_3890),
.B(n_3858),
.Y(n_3911)
);

INVx2_ASAP7_75t_SL g3912 ( 
.A(n_3889),
.Y(n_3912)
);

NAND2xp5_ASAP7_75t_L g3913 ( 
.A(n_3899),
.B(n_3836),
.Y(n_3913)
);

OAI322xp33_ASAP7_75t_L g3914 ( 
.A1(n_3909),
.A2(n_3807),
.A3(n_3831),
.B1(n_3818),
.B2(n_3766),
.C1(n_3760),
.C2(n_3769),
.Y(n_3914)
);

INVx2_ASAP7_75t_L g3915 ( 
.A(n_3908),
.Y(n_3915)
);

AOI21xp5_ASAP7_75t_L g3916 ( 
.A1(n_3902),
.A2(n_3653),
.B(n_3887),
.Y(n_3916)
);

INVx1_ASAP7_75t_L g3917 ( 
.A(n_3907),
.Y(n_3917)
);

INVx1_ASAP7_75t_L g3918 ( 
.A(n_3907),
.Y(n_3918)
);

AOI22xp5_ASAP7_75t_L g3919 ( 
.A1(n_3906),
.A2(n_3807),
.B1(n_3775),
.B2(n_3888),
.Y(n_3919)
);

INVx1_ASAP7_75t_L g3920 ( 
.A(n_3903),
.Y(n_3920)
);

INVx1_ASAP7_75t_L g3921 ( 
.A(n_3913),
.Y(n_3921)
);

NAND2xp5_ASAP7_75t_L g3922 ( 
.A(n_3917),
.B(n_3802),
.Y(n_3922)
);

INVx1_ASAP7_75t_L g3923 ( 
.A(n_3918),
.Y(n_3923)
);

AND2x2_ASAP7_75t_L g3924 ( 
.A(n_3919),
.B(n_3899),
.Y(n_3924)
);

OAI22xp5_ASAP7_75t_L g3925 ( 
.A1(n_3915),
.A2(n_3653),
.B1(n_3784),
.B2(n_3775),
.Y(n_3925)
);

INVx2_ASAP7_75t_L g3926 ( 
.A(n_3920),
.Y(n_3926)
);

OAI211xp5_ASAP7_75t_L g3927 ( 
.A1(n_3916),
.A2(n_3838),
.B(n_3828),
.C(n_3893),
.Y(n_3927)
);

INVx1_ASAP7_75t_L g3928 ( 
.A(n_3921),
.Y(n_3928)
);

AND2x2_ASAP7_75t_L g3929 ( 
.A(n_3914),
.B(n_3853),
.Y(n_3929)
);

INVx2_ASAP7_75t_L g3930 ( 
.A(n_3914),
.Y(n_3930)
);

AND2x2_ASAP7_75t_L g3931 ( 
.A(n_3919),
.B(n_3855),
.Y(n_3931)
);

NAND2xp5_ASAP7_75t_L g3932 ( 
.A(n_3917),
.B(n_3836),
.Y(n_3932)
);

OAI32xp33_ASAP7_75t_L g3933 ( 
.A1(n_3917),
.A2(n_3810),
.A3(n_3806),
.B1(n_3812),
.B2(n_3776),
.Y(n_3933)
);

INVx1_ASAP7_75t_L g3934 ( 
.A(n_3917),
.Y(n_3934)
);

OAI221xp5_ASAP7_75t_L g3935 ( 
.A1(n_3925),
.A2(n_3653),
.B1(n_3912),
.B2(n_3889),
.C(n_3780),
.Y(n_3935)
);

INVx1_ASAP7_75t_L g3936 ( 
.A(n_3922),
.Y(n_3936)
);

INVx1_ASAP7_75t_L g3937 ( 
.A(n_3922),
.Y(n_3937)
);

XNOR2xp5_ASAP7_75t_L g3938 ( 
.A(n_3925),
.B(n_3865),
.Y(n_3938)
);

NAND2xp5_ASAP7_75t_L g3939 ( 
.A(n_3929),
.B(n_3828),
.Y(n_3939)
);

INVx1_ASAP7_75t_L g3940 ( 
.A(n_3932),
.Y(n_3940)
);

INVx2_ASAP7_75t_SL g3941 ( 
.A(n_3923),
.Y(n_3941)
);

INVx1_ASAP7_75t_L g3942 ( 
.A(n_3934),
.Y(n_3942)
);

INVx1_ASAP7_75t_L g3943 ( 
.A(n_3924),
.Y(n_3943)
);

AND2x2_ASAP7_75t_L g3944 ( 
.A(n_3931),
.B(n_3861),
.Y(n_3944)
);

INVx2_ASAP7_75t_L g3945 ( 
.A(n_3926),
.Y(n_3945)
);

INVx1_ASAP7_75t_L g3946 ( 
.A(n_3927),
.Y(n_3946)
);

NAND2xp5_ASAP7_75t_SL g3947 ( 
.A(n_3930),
.B(n_3754),
.Y(n_3947)
);

OR2x2_ASAP7_75t_L g3948 ( 
.A(n_3928),
.B(n_3780),
.Y(n_3948)
);

OAI21xp33_ASAP7_75t_SL g3949 ( 
.A1(n_3933),
.A2(n_3769),
.B(n_3766),
.Y(n_3949)
);

AOI211xp5_ASAP7_75t_L g3950 ( 
.A1(n_3925),
.A2(n_3869),
.B(n_3872),
.C(n_3883),
.Y(n_3950)
);

INVx1_ASAP7_75t_L g3951 ( 
.A(n_3922),
.Y(n_3951)
);

NAND2xp5_ASAP7_75t_L g3952 ( 
.A(n_3925),
.B(n_3828),
.Y(n_3952)
);

NAND2xp33_ASAP7_75t_L g3953 ( 
.A(n_3925),
.B(n_3727),
.Y(n_3953)
);

AOI21xp5_ASAP7_75t_L g3954 ( 
.A1(n_3925),
.A2(n_3868),
.B(n_3866),
.Y(n_3954)
);

INVxp67_ASAP7_75t_SL g3955 ( 
.A(n_3922),
.Y(n_3955)
);

AOI321xp33_ASAP7_75t_L g3956 ( 
.A1(n_3925),
.A2(n_3847),
.A3(n_3910),
.B1(n_3885),
.B2(n_3892),
.C(n_3900),
.Y(n_3956)
);

OAI31xp33_ASAP7_75t_L g3957 ( 
.A1(n_3935),
.A2(n_3772),
.A3(n_3840),
.B(n_3843),
.Y(n_3957)
);

AOI221xp5_ASAP7_75t_L g3958 ( 
.A1(n_3947),
.A2(n_3772),
.B1(n_3838),
.B2(n_3805),
.C(n_3808),
.Y(n_3958)
);

NAND2xp5_ASAP7_75t_L g3959 ( 
.A(n_3950),
.B(n_3838),
.Y(n_3959)
);

OAI21xp5_ASAP7_75t_L g3960 ( 
.A1(n_3954),
.A2(n_3911),
.B(n_3886),
.Y(n_3960)
);

OAI22xp5_ASAP7_75t_L g3961 ( 
.A1(n_3939),
.A2(n_3857),
.B1(n_3635),
.B2(n_3658),
.Y(n_3961)
);

AOI22xp5_ASAP7_75t_L g3962 ( 
.A1(n_3943),
.A2(n_3782),
.B1(n_3655),
.B2(n_3667),
.Y(n_3962)
);

AOI22xp5_ASAP7_75t_L g3963 ( 
.A1(n_3944),
.A2(n_3782),
.B1(n_3658),
.B2(n_3773),
.Y(n_3963)
);

OAI22xp5_ASAP7_75t_L g3964 ( 
.A1(n_3946),
.A2(n_3724),
.B1(n_3714),
.B2(n_3730),
.Y(n_3964)
);

NAND2xp5_ASAP7_75t_L g3965 ( 
.A(n_3941),
.B(n_3874),
.Y(n_3965)
);

INVx1_ASAP7_75t_L g3966 ( 
.A(n_3948),
.Y(n_3966)
);

INVx1_ASAP7_75t_L g3967 ( 
.A(n_3952),
.Y(n_3967)
);

AOI221xp5_ASAP7_75t_L g3968 ( 
.A1(n_3953),
.A2(n_3805),
.B1(n_3808),
.B2(n_3822),
.C(n_3821),
.Y(n_3968)
);

NAND2xp5_ASAP7_75t_L g3969 ( 
.A(n_3955),
.B(n_3879),
.Y(n_3969)
);

OAI211xp5_ASAP7_75t_SL g3970 ( 
.A1(n_3956),
.A2(n_3942),
.B(n_3940),
.C(n_3904),
.Y(n_3970)
);

AOI31xp33_ASAP7_75t_L g3971 ( 
.A1(n_3938),
.A2(n_3905),
.A3(n_3894),
.B(n_3879),
.Y(n_3971)
);

NAND2x1_ASAP7_75t_L g3972 ( 
.A(n_3936),
.B(n_3863),
.Y(n_3972)
);

INVx1_ASAP7_75t_L g3973 ( 
.A(n_3937),
.Y(n_3973)
);

INVx1_ASAP7_75t_L g3974 ( 
.A(n_3951),
.Y(n_3974)
);

OAI21xp5_ASAP7_75t_SL g3975 ( 
.A1(n_3945),
.A2(n_3884),
.B(n_3863),
.Y(n_3975)
);

OAI221xp5_ASAP7_75t_SL g3976 ( 
.A1(n_3949),
.A2(n_3806),
.B1(n_3810),
.B2(n_3812),
.C(n_3785),
.Y(n_3976)
);

NAND2xp5_ASAP7_75t_L g3977 ( 
.A(n_3949),
.B(n_3880),
.Y(n_3977)
);

OAI21xp5_ASAP7_75t_L g3978 ( 
.A1(n_3954),
.A2(n_3880),
.B(n_3894),
.Y(n_3978)
);

AO21x1_ASAP7_75t_L g3979 ( 
.A1(n_3947),
.A2(n_3850),
.B(n_3849),
.Y(n_3979)
);

INVx1_ASAP7_75t_L g3980 ( 
.A(n_3939),
.Y(n_3980)
);

OAI211xp5_ASAP7_75t_L g3981 ( 
.A1(n_3950),
.A2(n_3811),
.B(n_3864),
.C(n_3859),
.Y(n_3981)
);

INVxp67_ASAP7_75t_SL g3982 ( 
.A(n_3948),
.Y(n_3982)
);

NOR3x1_ASAP7_75t_L g3983 ( 
.A(n_3975),
.B(n_3960),
.C(n_3978),
.Y(n_3983)
);

NOR2xp33_ASAP7_75t_L g3984 ( 
.A(n_3962),
.B(n_3844),
.Y(n_3984)
);

NAND4xp25_ASAP7_75t_L g3985 ( 
.A(n_3958),
.B(n_3811),
.C(n_3821),
.D(n_3822),
.Y(n_3985)
);

AOI222xp33_ASAP7_75t_L g3986 ( 
.A1(n_3968),
.A2(n_3776),
.B1(n_3777),
.B2(n_3783),
.C1(n_3787),
.C2(n_3785),
.Y(n_3986)
);

INVx1_ASAP7_75t_L g3987 ( 
.A(n_3963),
.Y(n_3987)
);

AOI221xp5_ASAP7_75t_L g3988 ( 
.A1(n_3971),
.A2(n_3811),
.B1(n_3777),
.B2(n_3740),
.C(n_3727),
.Y(n_3988)
);

AOI21xp5_ASAP7_75t_L g3989 ( 
.A1(n_3972),
.A2(n_3859),
.B(n_3819),
.Y(n_3989)
);

AOI322xp5_ASAP7_75t_L g3990 ( 
.A1(n_3967),
.A2(n_3783),
.A3(n_3787),
.B1(n_3687),
.B2(n_3651),
.C1(n_3628),
.C2(n_3676),
.Y(n_3990)
);

NOR3xp33_ASAP7_75t_L g3991 ( 
.A(n_3970),
.B(n_3819),
.C(n_3553),
.Y(n_3991)
);

NAND4xp25_ASAP7_75t_SL g3992 ( 
.A(n_3959),
.B(n_3835),
.C(n_3834),
.D(n_3827),
.Y(n_3992)
);

NAND2xp5_ASAP7_75t_L g3993 ( 
.A(n_3961),
.B(n_3773),
.Y(n_3993)
);

NAND3xp33_ASAP7_75t_L g3994 ( 
.A(n_3957),
.B(n_3833),
.C(n_3740),
.Y(n_3994)
);

AND2x4_ASAP7_75t_L g3995 ( 
.A(n_3982),
.B(n_3773),
.Y(n_3995)
);

AOI221x1_ASAP7_75t_L g3996 ( 
.A1(n_3977),
.A2(n_3835),
.B1(n_3834),
.B2(n_3827),
.C(n_3794),
.Y(n_3996)
);

AOI32xp33_ASAP7_75t_L g3997 ( 
.A1(n_3964),
.A2(n_3781),
.A3(n_3774),
.B1(n_3773),
.B2(n_3777),
.Y(n_3997)
);

NAND3xp33_ASAP7_75t_L g3998 ( 
.A(n_3981),
.B(n_3833),
.C(n_3740),
.Y(n_3998)
);

NOR3xp33_ASAP7_75t_L g3999 ( 
.A(n_3969),
.B(n_3538),
.C(n_3781),
.Y(n_3999)
);

AOI221xp5_ASAP7_75t_SL g4000 ( 
.A1(n_3965),
.A2(n_3794),
.B1(n_3793),
.B2(n_3795),
.C(n_3796),
.Y(n_4000)
);

NAND2xp5_ASAP7_75t_L g4001 ( 
.A(n_3979),
.B(n_3773),
.Y(n_4001)
);

NOR3xp33_ASAP7_75t_L g4002 ( 
.A(n_3980),
.B(n_3966),
.C(n_3973),
.Y(n_4002)
);

OAI211xp5_ASAP7_75t_SL g4003 ( 
.A1(n_3974),
.A2(n_3794),
.B(n_3793),
.C(n_3795),
.Y(n_4003)
);

OAI211xp5_ASAP7_75t_L g4004 ( 
.A1(n_3976),
.A2(n_3833),
.B(n_3777),
.C(n_3793),
.Y(n_4004)
);

AOI211xp5_ASAP7_75t_L g4005 ( 
.A1(n_3964),
.A2(n_3740),
.B(n_3727),
.C(n_3774),
.Y(n_4005)
);

AOI21xp5_ASAP7_75t_L g4006 ( 
.A1(n_3972),
.A2(n_3833),
.B(n_3796),
.Y(n_4006)
);

NAND4xp25_ASAP7_75t_L g4007 ( 
.A(n_3991),
.B(n_3774),
.C(n_3795),
.D(n_3796),
.Y(n_4007)
);

AOI322xp5_ASAP7_75t_L g4008 ( 
.A1(n_3984),
.A2(n_3774),
.A3(n_3644),
.B1(n_3688),
.B2(n_3651),
.C1(n_3654),
.C2(n_3661),
.Y(n_4008)
);

OAI211xp5_ASAP7_75t_L g4009 ( 
.A1(n_3988),
.A2(n_3833),
.B(n_3740),
.C(n_3727),
.Y(n_4009)
);

OAI21xp33_ASAP7_75t_L g4010 ( 
.A1(n_3987),
.A2(n_3774),
.B(n_3740),
.Y(n_4010)
);

AOI221xp5_ASAP7_75t_L g4011 ( 
.A1(n_3992),
.A2(n_3796),
.B1(n_3795),
.B2(n_3833),
.C(n_3799),
.Y(n_4011)
);

NAND4xp75_ASAP7_75t_L g4012 ( 
.A(n_3983),
.B(n_3723),
.C(n_3713),
.D(n_3757),
.Y(n_4012)
);

AOI21xp5_ASAP7_75t_L g4013 ( 
.A1(n_4006),
.A2(n_3771),
.B(n_3767),
.Y(n_4013)
);

OAI21xp33_ASAP7_75t_L g4014 ( 
.A1(n_3993),
.A2(n_3723),
.B(n_3799),
.Y(n_4014)
);

OAI221xp5_ASAP7_75t_L g4015 ( 
.A1(n_3997),
.A2(n_3709),
.B1(n_3706),
.B2(n_3707),
.C(n_3708),
.Y(n_4015)
);

NAND2xp5_ASAP7_75t_SL g4016 ( 
.A(n_3995),
.B(n_3799),
.Y(n_4016)
);

AOI321xp33_ASAP7_75t_L g4017 ( 
.A1(n_3999),
.A2(n_3770),
.A3(n_3767),
.B1(n_3771),
.B2(n_3755),
.C(n_3749),
.Y(n_4017)
);

OAI21xp5_ASAP7_75t_L g4018 ( 
.A1(n_3989),
.A2(n_3799),
.B(n_3770),
.Y(n_4018)
);

O2A1O1Ixp33_ASAP7_75t_SL g4019 ( 
.A1(n_4001),
.A2(n_3791),
.B(n_3792),
.C(n_3745),
.Y(n_4019)
);

XNOR2x1_ASAP7_75t_L g4020 ( 
.A(n_3995),
.B(n_3666),
.Y(n_4020)
);

AOI21xp5_ASAP7_75t_L g4021 ( 
.A1(n_4004),
.A2(n_3767),
.B(n_3771),
.Y(n_4021)
);

INVx1_ASAP7_75t_L g4022 ( 
.A(n_3996),
.Y(n_4022)
);

OAI21xp5_ASAP7_75t_L g4023 ( 
.A1(n_3994),
.A2(n_3799),
.B(n_3791),
.Y(n_4023)
);

NAND3xp33_ASAP7_75t_L g4024 ( 
.A(n_4016),
.B(n_4002),
.C(n_3998),
.Y(n_4024)
);

INVx2_ASAP7_75t_L g4025 ( 
.A(n_4020),
.Y(n_4025)
);

HB1xp67_ASAP7_75t_L g4026 ( 
.A(n_4012),
.Y(n_4026)
);

NOR2x1p5_ASAP7_75t_L g4027 ( 
.A(n_4007),
.B(n_3985),
.Y(n_4027)
);

OAI211xp5_ASAP7_75t_L g4028 ( 
.A1(n_4010),
.A2(n_4005),
.B(n_3986),
.C(n_4003),
.Y(n_4028)
);

A2O1A1Ixp33_ASAP7_75t_L g4029 ( 
.A1(n_4014),
.A2(n_4008),
.B(n_3990),
.C(n_4011),
.Y(n_4029)
);

NOR2xp33_ASAP7_75t_SL g4030 ( 
.A(n_4022),
.B(n_3671),
.Y(n_4030)
);

NAND4xp25_ASAP7_75t_L g4031 ( 
.A(n_4017),
.B(n_4000),
.C(n_3731),
.D(n_3729),
.Y(n_4031)
);

INVx1_ASAP7_75t_L g4032 ( 
.A(n_4019),
.Y(n_4032)
);

NAND3xp33_ASAP7_75t_SL g4033 ( 
.A(n_4009),
.B(n_3731),
.C(n_3741),
.Y(n_4033)
);

NAND4xp25_ASAP7_75t_L g4034 ( 
.A(n_4023),
.B(n_3724),
.C(n_3730),
.D(n_3714),
.Y(n_4034)
);

NOR2x1_ASAP7_75t_L g4035 ( 
.A(n_4018),
.B(n_3792),
.Y(n_4035)
);

OAI22xp5_ASAP7_75t_L g4036 ( 
.A1(n_4015),
.A2(n_3702),
.B1(n_3662),
.B2(n_3709),
.Y(n_4036)
);

INVx1_ASAP7_75t_L g4037 ( 
.A(n_4013),
.Y(n_4037)
);

AOI21xp5_ASAP7_75t_L g4038 ( 
.A1(n_4021),
.A2(n_3755),
.B(n_3750),
.Y(n_4038)
);

NAND2xp5_ASAP7_75t_L g4039 ( 
.A(n_4030),
.B(n_3666),
.Y(n_4039)
);

INVx2_ASAP7_75t_L g4040 ( 
.A(n_4035),
.Y(n_4040)
);

NAND2xp5_ASAP7_75t_SL g4041 ( 
.A(n_4024),
.B(n_3675),
.Y(n_4041)
);

NAND2xp5_ASAP7_75t_L g4042 ( 
.A(n_4036),
.B(n_3706),
.Y(n_4042)
);

NAND4xp25_ASAP7_75t_L g4043 ( 
.A(n_4029),
.B(n_3750),
.C(n_3749),
.D(n_3755),
.Y(n_4043)
);

NAND3xp33_ASAP7_75t_L g4044 ( 
.A(n_4028),
.B(n_3708),
.C(n_3707),
.Y(n_4044)
);

INVx1_ASAP7_75t_L g4045 ( 
.A(n_4034),
.Y(n_4045)
);

NOR2xp33_ASAP7_75t_L g4046 ( 
.A(n_4031),
.B(n_4026),
.Y(n_4046)
);

NAND4xp25_ASAP7_75t_L g4047 ( 
.A(n_4025),
.B(n_3750),
.C(n_3749),
.D(n_3741),
.Y(n_4047)
);

AOI211xp5_ASAP7_75t_L g4048 ( 
.A1(n_4033),
.A2(n_3738),
.B(n_3725),
.C(n_3728),
.Y(n_4048)
);

NAND2xp5_ASAP7_75t_L g4049 ( 
.A(n_4038),
.B(n_3648),
.Y(n_4049)
);

AOI211x1_ASAP7_75t_L g4050 ( 
.A1(n_4032),
.A2(n_3745),
.B(n_3789),
.C(n_3797),
.Y(n_4050)
);

AOI21xp33_ASAP7_75t_SL g4051 ( 
.A1(n_4037),
.A2(n_3837),
.B(n_3830),
.Y(n_4051)
);

OAI211xp5_ASAP7_75t_SL g4052 ( 
.A1(n_4027),
.A2(n_3746),
.B(n_3792),
.C(n_3829),
.Y(n_4052)
);

INVx1_ASAP7_75t_L g4053 ( 
.A(n_4035),
.Y(n_4053)
);

OAI211xp5_ASAP7_75t_SL g4054 ( 
.A1(n_4029),
.A2(n_3746),
.B(n_3830),
.C(n_3829),
.Y(n_4054)
);

NOR4xp75_ASAP7_75t_L g4055 ( 
.A(n_4033),
.B(n_3789),
.C(n_3797),
.D(n_3671),
.Y(n_4055)
);

NOR3xp33_ASAP7_75t_L g4056 ( 
.A(n_4024),
.B(n_3672),
.C(n_3588),
.Y(n_4056)
);

HB1xp67_ASAP7_75t_L g4057 ( 
.A(n_4055),
.Y(n_4057)
);

NOR2x1_ASAP7_75t_L g4058 ( 
.A(n_4053),
.B(n_3815),
.Y(n_4058)
);

INVx1_ASAP7_75t_L g4059 ( 
.A(n_4049),
.Y(n_4059)
);

AO211x2_ASAP7_75t_L g4060 ( 
.A1(n_4043),
.A2(n_3728),
.B(n_3743),
.C(n_3742),
.Y(n_4060)
);

OAI21xp5_ASAP7_75t_SL g4061 ( 
.A1(n_4056),
.A2(n_3789),
.B(n_3670),
.Y(n_4061)
);

INVx1_ASAP7_75t_L g4062 ( 
.A(n_4039),
.Y(n_4062)
);

HB1xp67_ASAP7_75t_L g4063 ( 
.A(n_4050),
.Y(n_4063)
);

AOI22xp33_ASAP7_75t_L g4064 ( 
.A1(n_4054),
.A2(n_3746),
.B1(n_3739),
.B2(n_3829),
.Y(n_4064)
);

NOR2x1_ASAP7_75t_L g4065 ( 
.A(n_4040),
.B(n_3815),
.Y(n_4065)
);

INVxp33_ASAP7_75t_SL g4066 ( 
.A(n_4046),
.Y(n_4066)
);

AOI22xp5_ASAP7_75t_L g4067 ( 
.A1(n_4041),
.A2(n_3675),
.B1(n_3672),
.B2(n_3670),
.Y(n_4067)
);

NOR2x1_ASAP7_75t_L g4068 ( 
.A(n_4052),
.B(n_3815),
.Y(n_4068)
);

AOI22xp5_ASAP7_75t_L g4069 ( 
.A1(n_4045),
.A2(n_3675),
.B1(n_3725),
.B2(n_3736),
.Y(n_4069)
);

INVx1_ASAP7_75t_L g4070 ( 
.A(n_4044),
.Y(n_4070)
);

NAND3xp33_ASAP7_75t_L g4071 ( 
.A(n_4051),
.B(n_3837),
.C(n_3823),
.Y(n_4071)
);

NAND2xp5_ASAP7_75t_SL g4072 ( 
.A(n_4048),
.B(n_3823),
.Y(n_4072)
);

AOI22xp5_ASAP7_75t_L g4073 ( 
.A1(n_4047),
.A2(n_3736),
.B1(n_3743),
.B2(n_3738),
.Y(n_4073)
);

NAND2xp5_ASAP7_75t_L g4074 ( 
.A(n_4067),
.B(n_4061),
.Y(n_4074)
);

OAI211xp5_ASAP7_75t_L g4075 ( 
.A1(n_4057),
.A2(n_4042),
.B(n_3837),
.C(n_3830),
.Y(n_4075)
);

NOR2xp33_ASAP7_75t_L g4076 ( 
.A(n_4066),
.B(n_3588),
.Y(n_4076)
);

NOR3xp33_ASAP7_75t_L g4077 ( 
.A(n_4062),
.B(n_3826),
.C(n_3823),
.Y(n_4077)
);

NAND4xp25_ASAP7_75t_SL g4078 ( 
.A(n_4069),
.B(n_3682),
.C(n_3664),
.D(n_3663),
.Y(n_4078)
);

NOR2x1_ASAP7_75t_L g4079 ( 
.A(n_4058),
.B(n_3826),
.Y(n_4079)
);

OR2x2_ASAP7_75t_L g4080 ( 
.A(n_4073),
.B(n_3742),
.Y(n_4080)
);

NOR2x1_ASAP7_75t_L g4081 ( 
.A(n_4065),
.B(n_3826),
.Y(n_4081)
);

AOI221xp5_ASAP7_75t_L g4082 ( 
.A1(n_4064),
.A2(n_3739),
.B1(n_3687),
.B2(n_3686),
.C(n_3682),
.Y(n_4082)
);

OAI22xp5_ASAP7_75t_L g4083 ( 
.A1(n_4059),
.A2(n_3654),
.B1(n_3644),
.B2(n_3688),
.Y(n_4083)
);

AND2x2_ASAP7_75t_L g4084 ( 
.A(n_4068),
.B(n_3693),
.Y(n_4084)
);

AND2x2_ASAP7_75t_L g4085 ( 
.A(n_4076),
.B(n_4063),
.Y(n_4085)
);

NAND2xp5_ASAP7_75t_L g4086 ( 
.A(n_4084),
.B(n_4060),
.Y(n_4086)
);

NOR2x1_ASAP7_75t_L g4087 ( 
.A(n_4079),
.B(n_4071),
.Y(n_4087)
);

AOI32xp33_ASAP7_75t_L g4088 ( 
.A1(n_4077),
.A2(n_4070),
.A3(n_4072),
.B1(n_3797),
.B2(n_3663),
.Y(n_4088)
);

NAND4xp75_ASAP7_75t_L g4089 ( 
.A(n_4074),
.B(n_3693),
.C(n_3661),
.D(n_3681),
.Y(n_4089)
);

AOI21xp5_ASAP7_75t_L g4090 ( 
.A1(n_4075),
.A2(n_3676),
.B(n_3681),
.Y(n_4090)
);

NOR2x1_ASAP7_75t_L g4091 ( 
.A(n_4087),
.B(n_4081),
.Y(n_4091)
);

OR2x2_ASAP7_75t_L g4092 ( 
.A(n_4089),
.B(n_4080),
.Y(n_4092)
);

NOR3xp33_ASAP7_75t_L g4093 ( 
.A(n_4086),
.B(n_4078),
.C(n_4083),
.Y(n_4093)
);

INVx2_ASAP7_75t_L g4094 ( 
.A(n_4091),
.Y(n_4094)
);

INVx1_ASAP7_75t_L g4095 ( 
.A(n_4092),
.Y(n_4095)
);

XOR2xp5_ASAP7_75t_L g4096 ( 
.A(n_4095),
.B(n_4085),
.Y(n_4096)
);

OAI21xp33_ASAP7_75t_L g4097 ( 
.A1(n_4096),
.A2(n_4088),
.B(n_4094),
.Y(n_4097)
);

NOR2xp33_ASAP7_75t_L g4098 ( 
.A(n_4097),
.B(n_4093),
.Y(n_4098)
);

AOI22xp5_ASAP7_75t_L g4099 ( 
.A1(n_4098),
.A2(n_4090),
.B1(n_4082),
.B2(n_3615),
.Y(n_4099)
);

OAI22xp5_ASAP7_75t_SL g4100 ( 
.A1(n_4099),
.A2(n_3615),
.B1(n_3595),
.B2(n_3617),
.Y(n_4100)
);

INVx1_ASAP7_75t_L g4101 ( 
.A(n_4100),
.Y(n_4101)
);

NAND2xp5_ASAP7_75t_L g4102 ( 
.A(n_4101),
.B(n_3641),
.Y(n_4102)
);

INVx1_ASAP7_75t_L g4103 ( 
.A(n_4102),
.Y(n_4103)
);

NAND3xp33_ASAP7_75t_L g4104 ( 
.A(n_4103),
.B(n_3617),
.C(n_3616),
.Y(n_4104)
);

INVx1_ASAP7_75t_L g4105 ( 
.A(n_4104),
.Y(n_4105)
);

OA21x2_ASAP7_75t_L g4106 ( 
.A1(n_4105),
.A2(n_3616),
.B(n_3618),
.Y(n_4106)
);

OAI221xp5_ASAP7_75t_R g4107 ( 
.A1(n_4106),
.A2(n_3684),
.B1(n_3555),
.B2(n_3622),
.C(n_3554),
.Y(n_4107)
);

AOI21xp33_ASAP7_75t_SL g4108 ( 
.A1(n_4107),
.A2(n_3595),
.B(n_3555),
.Y(n_4108)
);

AOI211xp5_ASAP7_75t_L g4109 ( 
.A1(n_4108),
.A2(n_3630),
.B(n_3637),
.C(n_3625),
.Y(n_4109)
);


endmodule