module fake_jpeg_14401_n_256 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_256);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_256;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_251;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_125;
wire n_80;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_247;
wire n_87;
wire n_46;
wire n_157;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_140;
wire n_128;
wire n_82;
wire n_96;

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_10),
.Y(n_15)
);

INVx3_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_14),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

INVx4_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

INVx2_ASAP7_75t_SL g25 ( 
.A(n_12),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_10),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_5),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_13),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_5),
.Y(n_35)
);

INVxp67_ASAP7_75t_L g36 ( 
.A(n_2),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_5),
.Y(n_37)
);

BUFx10_ASAP7_75t_L g38 ( 
.A(n_6),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_3),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_10),
.Y(n_40)
);

HAxp5_ASAP7_75t_SL g41 ( 
.A(n_38),
.B(n_0),
.CON(n_41),
.SN(n_41)
);

NAND2xp33_ASAP7_75t_SL g118 ( 
.A(n_41),
.B(n_73),
.Y(n_118)
);

INVx4_ASAP7_75t_SL g42 ( 
.A(n_38),
.Y(n_42)
);

AND2x2_ASAP7_75t_L g115 ( 
.A(n_42),
.B(n_46),
.Y(n_115)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_21),
.Y(n_43)
);

BUFx2_ASAP7_75t_L g81 ( 
.A(n_43),
.Y(n_81)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_20),
.Y(n_44)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_44),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g45 ( 
.A(n_30),
.B(n_33),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_45),
.B(n_58),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g46 ( 
.A(n_25),
.B(n_0),
.Y(n_46)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_15),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_47),
.Y(n_79)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_20),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g92 ( 
.A(n_48),
.Y(n_92)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_29),
.Y(n_49)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_49),
.Y(n_102)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_28),
.Y(n_50)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_50),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_15),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_51),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_32),
.B(n_0),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_52),
.B(n_54),
.Y(n_86)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_29),
.Y(n_53)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_53),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_36),
.B(n_1),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_36),
.B(n_1),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_55),
.B(n_57),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

INVx6_ASAP7_75t_L g82 ( 
.A(n_56),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_37),
.B(n_2),
.Y(n_57)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_25),
.B(n_3),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_37),
.B(n_4),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_59),
.B(n_6),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_38),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_60),
.B(n_67),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_39),
.Y(n_61)
);

INVx6_ASAP7_75t_L g87 ( 
.A(n_61),
.Y(n_87)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_21),
.Y(n_62)
);

BUFx2_ASAP7_75t_L g85 ( 
.A(n_62),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_17),
.Y(n_63)
);

INVx6_ASAP7_75t_L g89 ( 
.A(n_63),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_28),
.B(n_6),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_64),
.B(n_78),
.Y(n_91)
);

INVx11_ASAP7_75t_L g65 ( 
.A(n_38),
.Y(n_65)
);

INVx11_ASAP7_75t_L g114 ( 
.A(n_65),
.Y(n_114)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_17),
.Y(n_66)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_66),
.Y(n_107)
);

INVx13_ASAP7_75t_L g67 ( 
.A(n_25),
.Y(n_67)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_17),
.Y(n_68)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_68),
.Y(n_83)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_17),
.Y(n_69)
);

INVx5_ASAP7_75t_L g116 ( 
.A(n_69),
.Y(n_116)
);

BUFx2_ASAP7_75t_L g70 ( 
.A(n_16),
.Y(n_70)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_70),
.Y(n_93)
);

BUFx12f_ASAP7_75t_L g71 ( 
.A(n_23),
.Y(n_71)
);

INVx6_ASAP7_75t_L g110 ( 
.A(n_71),
.Y(n_110)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_19),
.Y(n_72)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_72),
.Y(n_113)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_19),
.Y(n_73)
);

BUFx12f_ASAP7_75t_L g74 ( 
.A(n_23),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_74),
.B(n_77),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_19),
.Y(n_75)
);

INVx8_ASAP7_75t_L g104 ( 
.A(n_75),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_19),
.Y(n_76)
);

INVx8_ASAP7_75t_L g109 ( 
.A(n_76),
.Y(n_109)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_34),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_34),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_88),
.B(n_105),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_L g90 ( 
.A1(n_51),
.A2(n_16),
.B1(n_40),
.B2(n_18),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_90),
.A2(n_97),
.B1(n_99),
.B2(n_111),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_52),
.B(n_40),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_95),
.B(n_96),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_57),
.B(n_35),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_46),
.A2(n_58),
.B1(n_61),
.B2(n_56),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_L g99 ( 
.A1(n_70),
.A2(n_22),
.B1(n_27),
.B2(n_26),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_54),
.B(n_22),
.C(n_27),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_SL g151 ( 
.A1(n_100),
.A2(n_108),
.B(n_118),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_59),
.B(n_18),
.Y(n_105)
);

AOI21xp33_ASAP7_75t_SL g108 ( 
.A1(n_55),
.A2(n_34),
.B(n_24),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_71),
.A2(n_24),
.B1(n_31),
.B2(n_34),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_63),
.B(n_35),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_112),
.B(n_85),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_74),
.A2(n_31),
.B1(n_26),
.B2(n_11),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_117),
.A2(n_78),
.B1(n_76),
.B2(n_75),
.Y(n_121)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_99),
.Y(n_120)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_120),
.Y(n_159)
);

OAI22xp33_ASAP7_75t_L g169 ( 
.A1(n_121),
.A2(n_116),
.B1(n_119),
.B2(n_89),
.Y(n_169)
);

INVx2_ASAP7_75t_SL g122 ( 
.A(n_107),
.Y(n_122)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_122),
.Y(n_161)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_104),
.Y(n_123)
);

BUFx2_ASAP7_75t_L g166 ( 
.A(n_123),
.Y(n_166)
);

BUFx10_ASAP7_75t_L g125 ( 
.A(n_114),
.Y(n_125)
);

BUFx2_ASAP7_75t_L g168 ( 
.A(n_125),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_86),
.B(n_8),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_SL g180 ( 
.A(n_126),
.B(n_128),
.Y(n_180)
);

INVx13_ASAP7_75t_L g127 ( 
.A(n_101),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_127),
.B(n_135),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_98),
.B(n_8),
.Y(n_128)
);

INVx1_ASAP7_75t_SL g129 ( 
.A(n_81),
.Y(n_129)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_129),
.Y(n_163)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_93),
.Y(n_130)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_130),
.Y(n_173)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_104),
.Y(n_131)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_131),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_84),
.B(n_9),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g181 ( 
.A(n_132),
.B(n_136),
.Y(n_181)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_80),
.Y(n_133)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_133),
.Y(n_176)
);

INVx11_ASAP7_75t_L g134 ( 
.A(n_114),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_134),
.Y(n_157)
);

BUFx3_ASAP7_75t_L g135 ( 
.A(n_110),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_91),
.B(n_11),
.Y(n_136)
);

INVx4_ASAP7_75t_L g137 ( 
.A(n_109),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_137),
.B(n_139),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_90),
.A2(n_42),
.B1(n_12),
.B2(n_13),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_138),
.A2(n_140),
.B1(n_92),
.B2(n_85),
.Y(n_162)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_109),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_111),
.A2(n_11),
.B1(n_12),
.B2(n_117),
.Y(n_140)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_83),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_142),
.B(n_143),
.Y(n_174)
);

INVx1_ASAP7_75t_SL g143 ( 
.A(n_81),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_115),
.A2(n_79),
.B1(n_82),
.B2(n_87),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_144),
.A2(n_122),
.B1(n_143),
.B2(n_129),
.Y(n_172)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_113),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_145),
.B(n_146),
.Y(n_175)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_110),
.Y(n_146)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_107),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_147),
.B(n_150),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_115),
.B(n_103),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_149),
.B(n_151),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_89),
.Y(n_150)
);

OAI21xp33_ASAP7_75t_L g164 ( 
.A1(n_152),
.A2(n_106),
.B(n_92),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_94),
.B(n_102),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_153),
.B(n_154),
.Y(n_160)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_82),
.Y(n_154)
);

BUFx2_ASAP7_75t_L g155 ( 
.A(n_116),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_155),
.B(n_122),
.Y(n_182)
);

OA22x2_ASAP7_75t_L g158 ( 
.A1(n_120),
.A2(n_106),
.B1(n_79),
.B2(n_119),
.Y(n_158)
);

OA21x2_ASAP7_75t_L g202 ( 
.A1(n_158),
.A2(n_125),
.B(n_172),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_162),
.A2(n_177),
.B1(n_144),
.B2(n_131),
.Y(n_190)
);

AND2x2_ASAP7_75t_L g199 ( 
.A(n_164),
.B(n_179),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_152),
.B(n_87),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_167),
.B(n_178),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_169),
.A2(n_172),
.B1(n_125),
.B2(n_135),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_124),
.A2(n_138),
.B1(n_140),
.B2(n_151),
.Y(n_177)
);

AO22x2_ASAP7_75t_L g179 ( 
.A1(n_137),
.A2(n_133),
.B1(n_123),
.B2(n_139),
.Y(n_179)
);

CKINVDCx14_ASAP7_75t_R g188 ( 
.A(n_182),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_183),
.B(n_185),
.Y(n_206)
);

BUFx3_ASAP7_75t_L g184 ( 
.A(n_166),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_184),
.B(n_189),
.Y(n_203)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_173),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_165),
.B(n_148),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_SL g204 ( 
.A(n_186),
.B(n_191),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_156),
.B(n_167),
.C(n_177),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_187),
.B(n_195),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_182),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_190),
.A2(n_202),
.B1(n_199),
.B2(n_188),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_181),
.B(n_141),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_160),
.B(n_130),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_192),
.B(n_193),
.Y(n_211)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_173),
.Y(n_193)
);

BUFx2_ASAP7_75t_L g194 ( 
.A(n_161),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_194),
.B(n_197),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_160),
.B(n_127),
.Y(n_195)
);

AOI22xp33_ASAP7_75t_L g196 ( 
.A1(n_159),
.A2(n_154),
.B1(n_146),
.B2(n_147),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_196),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_180),
.B(n_155),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_SL g198 ( 
.A1(n_162),
.A2(n_125),
.B(n_134),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_198),
.B(n_158),
.Y(n_209)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_161),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_200),
.B(n_159),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_201),
.A2(n_169),
.B1(n_158),
.B2(n_171),
.Y(n_216)
);

AND2x2_ASAP7_75t_L g222 ( 
.A(n_209),
.B(n_212),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_191),
.B(n_175),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_210),
.B(n_213),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_183),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_192),
.Y(n_214)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_214),
.Y(n_223)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_215),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_216),
.A2(n_202),
.B1(n_198),
.B2(n_201),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_205),
.B(n_187),
.C(n_195),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_217),
.B(n_219),
.C(n_221),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_205),
.B(n_189),
.C(n_190),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_216),
.A2(n_199),
.B1(n_200),
.B2(n_194),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_220),
.B(n_212),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_206),
.B(n_185),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_206),
.B(n_193),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_224),
.B(n_203),
.C(n_211),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_213),
.A2(n_199),
.B1(n_202),
.B2(n_194),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_225),
.B(n_226),
.Y(n_229)
);

AOI21xp5_ASAP7_75t_L g238 ( 
.A1(n_230),
.A2(n_231),
.B(n_235),
.Y(n_238)
);

AND2x2_ASAP7_75t_L g231 ( 
.A(n_219),
.B(n_208),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_232),
.B(n_233),
.C(n_234),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_217),
.B(n_211),
.C(n_214),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_218),
.B(n_204),
.C(n_170),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_223),
.B(n_204),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_L g236 ( 
.A1(n_229),
.A2(n_227),
.B1(n_225),
.B2(n_215),
.Y(n_236)
);

OR2x2_ASAP7_75t_L g242 ( 
.A(n_236),
.B(n_179),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_228),
.B(n_224),
.C(n_221),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_237),
.B(n_184),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_229),
.A2(n_222),
.B1(n_207),
.B2(n_202),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_L g243 ( 
.A1(n_240),
.A2(n_241),
.B(n_207),
.Y(n_243)
);

AOI21xp5_ASAP7_75t_L g241 ( 
.A1(n_234),
.A2(n_222),
.B(n_174),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_242),
.A2(n_243),
.B1(n_238),
.B2(n_179),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_244),
.B(n_245),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_239),
.B(n_170),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_237),
.B(n_166),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_SL g250 ( 
.A1(n_246),
.A2(n_176),
.B(n_163),
.Y(n_250)
);

INVxp67_ASAP7_75t_L g251 ( 
.A(n_247),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_245),
.A2(n_158),
.B1(n_157),
.B2(n_168),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_249),
.B(n_250),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_252),
.B(n_248),
.C(n_247),
.Y(n_253)
);

AOI22xp33_ASAP7_75t_L g255 ( 
.A1(n_253),
.A2(n_254),
.B1(n_157),
.B2(n_179),
.Y(n_255)
);

OAI21xp5_ASAP7_75t_L g254 ( 
.A1(n_251),
.A2(n_249),
.B(n_168),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_255),
.B(n_163),
.Y(n_256)
);


endmodule