module fake_jpeg_19756_n_35 (n_3, n_2, n_1, n_0, n_4, n_5, n_35);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_35;

wire n_13;
wire n_21;
wire n_33;
wire n_10;
wire n_23;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_34;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_9;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

BUFx12f_ASAP7_75t_L g6 ( 
.A(n_5),
.Y(n_6)
);

CKINVDCx20_ASAP7_75t_R g7 ( 
.A(n_1),
.Y(n_7)
);

INVx5_ASAP7_75t_L g8 ( 
.A(n_0),
.Y(n_8)
);

BUFx6f_ASAP7_75t_L g9 ( 
.A(n_5),
.Y(n_9)
);

INVx2_ASAP7_75t_L g10 ( 
.A(n_3),
.Y(n_10)
);

INVx4_ASAP7_75t_L g11 ( 
.A(n_6),
.Y(n_11)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

INVx8_ASAP7_75t_L g12 ( 
.A(n_6),
.Y(n_12)
);

AOI22xp5_ASAP7_75t_SL g16 ( 
.A1(n_12),
.A2(n_13),
.B1(n_14),
.B2(n_10),
.Y(n_16)
);

AO22x1_ASAP7_75t_SL g13 ( 
.A1(n_8),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_13)
);

INVx3_ASAP7_75t_L g14 ( 
.A(n_10),
.Y(n_14)
);

CKINVDCx12_ASAP7_75t_R g15 ( 
.A(n_12),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_15),
.B(n_12),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_SL g21 ( 
.A1(n_16),
.A2(n_11),
.B1(n_14),
.B2(n_13),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_17),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_SL g23 ( 
.A(n_18),
.B(n_20),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_19),
.B(n_6),
.Y(n_25)
);

AOI22xp5_ASAP7_75t_L g20 ( 
.A1(n_16),
.A2(n_14),
.B1(n_13),
.B2(n_11),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_L g22 ( 
.A(n_21),
.B(n_13),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_SL g26 ( 
.A(n_22),
.B(n_25),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_SL g24 ( 
.A(n_18),
.B(n_7),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_SL g28 ( 
.A(n_24),
.B(n_7),
.Y(n_28)
);

BUFx12f_ASAP7_75t_SL g27 ( 
.A(n_23),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_27),
.B(n_28),
.Y(n_30)
);

HB1xp67_ASAP7_75t_L g29 ( 
.A(n_27),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_29),
.B(n_31),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_L g31 ( 
.A1(n_26),
.A2(n_20),
.B1(n_21),
.B2(n_22),
.Y(n_31)
);

AOI21xp33_ASAP7_75t_L g33 ( 
.A1(n_32),
.A2(n_4),
.B(n_9),
.Y(n_33)
);

OAI321xp33_ASAP7_75t_L g34 ( 
.A1(n_33),
.A2(n_2),
.A3(n_3),
.B1(n_4),
.B2(n_9),
.C(n_30),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_34),
.Y(n_35)
);


endmodule