module real_jpeg_29385_n_7 (n_5, n_4, n_0, n_1, n_2, n_6, n_30, n_28, n_29, n_3, n_7);

input n_5;
input n_4;
input n_0;
input n_1;
input n_2;
input n_6;
input n_30;
input n_28;
input n_29;
input n_3;

output n_7;

wire n_17;
wire n_8;
wire n_21;
wire n_10;
wire n_9;
wire n_12;
wire n_24;
wire n_23;
wire n_11;
wire n_14;
wire n_25;
wire n_22;
wire n_18;
wire n_26;
wire n_20;
wire n_19;
wire n_16;
wire n_15;
wire n_13;

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_0),
.Y(n_12)
);

AOI21xp5_ASAP7_75t_L g25 ( 
.A1(n_1),
.A2(n_3),
.B(n_19),
.Y(n_25)
);

NAND3xp33_ASAP7_75t_L g26 ( 
.A(n_1),
.B(n_3),
.C(n_19),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_2),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_4),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_5),
.Y(n_22)
);

NAND3xp33_ASAP7_75t_L g24 ( 
.A(n_5),
.B(n_19),
.C(n_30),
.Y(n_24)
);

NOR3xp33_ASAP7_75t_L g10 ( 
.A(n_6),
.B(n_11),
.C(n_12),
.Y(n_10)
);

OAI21xp5_ASAP7_75t_L g13 ( 
.A1(n_6),
.A2(n_11),
.B(n_12),
.Y(n_13)
);

INVx4_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

OAI21xp5_ASAP7_75t_L g20 ( 
.A1(n_6),
.A2(n_21),
.B(n_22),
.Y(n_20)
);

XOR2xp5_ASAP7_75t_L g7 ( 
.A(n_8),
.B(n_14),
.Y(n_7)
);

NAND2xp5_ASAP7_75t_L g8 ( 
.A(n_9),
.B(n_13),
.Y(n_8)
);

CKINVDCx20_ASAP7_75t_R g9 ( 
.A(n_10),
.Y(n_9)
);

OAI21xp5_ASAP7_75t_SL g14 ( 
.A1(n_15),
.A2(n_25),
.B(n_26),
.Y(n_14)
);

AOI21xp5_ASAP7_75t_L g15 ( 
.A1(n_16),
.A2(n_20),
.B(n_23),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_18),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_28),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_24),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_29),
.Y(n_21)
);


endmodule