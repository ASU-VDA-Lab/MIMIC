module fake_jpeg_2709_n_473 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_473);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_473;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_2),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_13),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

INVx11_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

INVx6_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_1),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_16),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_1),
.Y(n_35)
);

INVx6_ASAP7_75t_SL g36 ( 
.A(n_15),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_9),
.Y(n_37)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_1),
.Y(n_39)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_2),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_13),
.Y(n_41)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_12),
.Y(n_42)
);

INVx1_ASAP7_75t_SL g43 ( 
.A(n_6),
.Y(n_43)
);

INVx8_ASAP7_75t_SL g44 ( 
.A(n_0),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_7),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_9),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_13),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_7),
.Y(n_48)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_4),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_0),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_15),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_10),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_14),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_10),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_9),
.Y(n_55)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_11),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_19),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_57),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_36),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_58),
.B(n_72),
.Y(n_122)
);

INVx11_ASAP7_75t_L g59 ( 
.A(n_33),
.Y(n_59)
);

INVx4_ASAP7_75t_L g123 ( 
.A(n_59),
.Y(n_123)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_36),
.Y(n_60)
);

INVx4_ASAP7_75t_SL g153 ( 
.A(n_60),
.Y(n_153)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_19),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_61),
.Y(n_151)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_49),
.Y(n_62)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_62),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_19),
.Y(n_63)
);

INVx6_ASAP7_75t_L g141 ( 
.A(n_63),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_51),
.B(n_15),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_64),
.B(n_65),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_51),
.B(n_16),
.Y(n_65)
);

BUFx2_ASAP7_75t_L g66 ( 
.A(n_22),
.Y(n_66)
);

BUFx2_ASAP7_75t_L g120 ( 
.A(n_66),
.Y(n_120)
);

BUFx4f_ASAP7_75t_L g67 ( 
.A(n_29),
.Y(n_67)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_67),
.Y(n_139)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_33),
.Y(n_68)
);

INVx5_ASAP7_75t_L g117 ( 
.A(n_68),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_32),
.Y(n_69)
);

INVx6_ASAP7_75t_L g157 ( 
.A(n_69),
.Y(n_157)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_33),
.Y(n_70)
);

INVx5_ASAP7_75t_L g124 ( 
.A(n_70),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_32),
.Y(n_71)
);

INVx6_ASAP7_75t_L g175 ( 
.A(n_71),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_44),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_44),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_73),
.B(n_82),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_32),
.Y(n_74)
);

INVx8_ASAP7_75t_L g121 ( 
.A(n_74),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_41),
.Y(n_75)
);

INVx8_ASAP7_75t_L g130 ( 
.A(n_75),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_24),
.B(n_3),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_76),
.B(n_93),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_41),
.Y(n_77)
);

BUFx3_ASAP7_75t_L g155 ( 
.A(n_77),
.Y(n_155)
);

INVx2_ASAP7_75t_SL g78 ( 
.A(n_29),
.Y(n_78)
);

INVx4_ASAP7_75t_L g126 ( 
.A(n_78),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_49),
.B(n_14),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g156 ( 
.A(n_79),
.B(n_86),
.Y(n_156)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_24),
.Y(n_80)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_80),
.Y(n_145)
);

BUFx12_ASAP7_75t_L g81 ( 
.A(n_30),
.Y(n_81)
);

BUFx12f_ASAP7_75t_L g181 ( 
.A(n_81),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_21),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_41),
.Y(n_83)
);

INVx5_ASAP7_75t_L g137 ( 
.A(n_83),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_52),
.Y(n_84)
);

INVx5_ASAP7_75t_L g138 ( 
.A(n_84),
.Y(n_138)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_29),
.Y(n_85)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_85),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_55),
.B(n_14),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_52),
.Y(n_87)
);

INVx4_ASAP7_75t_L g134 ( 
.A(n_87),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_21),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_88),
.B(n_97),
.Y(n_129)
);

BUFx12f_ASAP7_75t_L g89 ( 
.A(n_56),
.Y(n_89)
);

INVx4_ASAP7_75t_L g140 ( 
.A(n_89),
.Y(n_140)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_55),
.Y(n_90)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_90),
.Y(n_147)
);

HB1xp67_ASAP7_75t_L g91 ( 
.A(n_22),
.Y(n_91)
);

HB1xp67_ASAP7_75t_L g186 ( 
.A(n_91),
.Y(n_186)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_22),
.Y(n_92)
);

INVx3_ASAP7_75t_L g162 ( 
.A(n_92),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_30),
.B(n_3),
.Y(n_93)
);

INVx11_ASAP7_75t_L g94 ( 
.A(n_33),
.Y(n_94)
);

INVx4_ASAP7_75t_L g149 ( 
.A(n_94),
.Y(n_149)
);

BUFx5_ASAP7_75t_L g95 ( 
.A(n_23),
.Y(n_95)
);

INVx4_ASAP7_75t_L g179 ( 
.A(n_95),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_52),
.Y(n_96)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_96),
.Y(n_148)
);

NOR3xp33_ASAP7_75t_L g97 ( 
.A(n_43),
.B(n_4),
.C(n_5),
.Y(n_97)
);

INVx8_ASAP7_75t_L g98 ( 
.A(n_33),
.Y(n_98)
);

INVx3_ASAP7_75t_L g176 ( 
.A(n_98),
.Y(n_176)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_26),
.Y(n_99)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_99),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_30),
.B(n_4),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g178 ( 
.A(n_100),
.B(n_5),
.Y(n_178)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_26),
.Y(n_101)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_101),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_54),
.Y(n_102)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_102),
.Y(n_171)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_23),
.Y(n_103)
);

INVx3_ASAP7_75t_L g183 ( 
.A(n_103),
.Y(n_183)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_27),
.Y(n_104)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_104),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_54),
.Y(n_105)
);

NAND2x1_ASAP7_75t_SL g163 ( 
.A(n_105),
.B(n_110),
.Y(n_163)
);

INVx6_ASAP7_75t_SL g106 ( 
.A(n_38),
.Y(n_106)
);

INVx13_ASAP7_75t_L g150 ( 
.A(n_106),
.Y(n_150)
);

BUFx4f_ASAP7_75t_L g107 ( 
.A(n_20),
.Y(n_107)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_107),
.Y(n_164)
);

BUFx3_ASAP7_75t_L g108 ( 
.A(n_56),
.Y(n_108)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_108),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_21),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_109),
.B(n_111),
.Y(n_132)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_23),
.Y(n_110)
);

BUFx12f_ASAP7_75t_L g111 ( 
.A(n_56),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_54),
.Y(n_112)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_112),
.Y(n_168)
);

BUFx3_ASAP7_75t_L g113 ( 
.A(n_26),
.Y(n_113)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_113),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_40),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_114),
.B(n_31),
.Y(n_166)
);

INVx8_ASAP7_75t_L g115 ( 
.A(n_30),
.Y(n_115)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_115),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_40),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_116),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_101),
.B(n_37),
.C(n_50),
.Y(n_118)
);

AND2x2_ASAP7_75t_L g221 ( 
.A(n_118),
.B(n_161),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_57),
.A2(n_37),
.B1(n_50),
.B2(n_48),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_119),
.A2(n_133),
.B1(n_159),
.B2(n_160),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_61),
.A2(n_30),
.B1(n_40),
.B2(n_25),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_131),
.A2(n_146),
.B1(n_182),
.B2(n_95),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_63),
.A2(n_53),
.B1(n_25),
.B2(n_18),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_106),
.A2(n_43),
.B1(n_20),
.B2(n_47),
.Y(n_136)
);

OA22x2_ASAP7_75t_L g243 ( 
.A1(n_136),
.A2(n_144),
.B1(n_172),
.B2(n_81),
.Y(n_243)
);

AOI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_78),
.A2(n_43),
.B1(n_20),
.B2(n_47),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_116),
.A2(n_18),
.B1(n_17),
.B2(n_53),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_L g159 ( 
.A1(n_69),
.A2(n_27),
.B1(n_46),
.B2(n_45),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_71),
.A2(n_28),
.B1(n_46),
.B2(n_45),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_92),
.B(n_48),
.C(n_35),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_L g165 ( 
.A1(n_74),
.A2(n_28),
.B1(n_35),
.B2(n_31),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_165),
.A2(n_174),
.B1(n_180),
.B2(n_185),
.Y(n_212)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_166),
.Y(n_189)
);

AOI22xp33_ASAP7_75t_SL g172 ( 
.A1(n_107),
.A2(n_103),
.B1(n_110),
.B2(n_108),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_L g174 ( 
.A1(n_75),
.A2(n_17),
.B1(n_39),
.B2(n_34),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_60),
.B(n_5),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_SL g188 ( 
.A(n_177),
.B(n_67),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_178),
.B(n_60),
.Y(n_203)
);

OAI22xp33_ASAP7_75t_L g180 ( 
.A1(n_77),
.A2(n_39),
.B1(n_42),
.B2(n_34),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_83),
.A2(n_38),
.B1(n_42),
.B2(n_39),
.Y(n_182)
);

AND2x2_ASAP7_75t_SL g184 ( 
.A(n_85),
.B(n_38),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_184),
.Y(n_244)
);

AOI22xp33_ASAP7_75t_L g185 ( 
.A1(n_84),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_185)
);

INVx3_ASAP7_75t_L g187 ( 
.A(n_126),
.Y(n_187)
);

INVx3_ASAP7_75t_L g287 ( 
.A(n_187),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_188),
.B(n_194),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_156),
.B(n_67),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_191),
.B(n_198),
.Y(n_247)
);

OR2x2_ASAP7_75t_L g192 ( 
.A(n_125),
.B(n_66),
.Y(n_192)
);

CKINVDCx14_ASAP7_75t_R g248 ( 
.A(n_192),
.Y(n_248)
);

AOI22xp33_ASAP7_75t_SL g193 ( 
.A1(n_129),
.A2(n_107),
.B1(n_111),
.B2(n_89),
.Y(n_193)
);

INVxp67_ASAP7_75t_L g250 ( 
.A(n_193),
.Y(n_250)
);

OR2x2_ASAP7_75t_L g194 ( 
.A(n_145),
.B(n_113),
.Y(n_194)
);

CKINVDCx16_ASAP7_75t_R g195 ( 
.A(n_122),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_195),
.B(n_203),
.Y(n_284)
);

BUFx2_ASAP7_75t_L g196 ( 
.A(n_120),
.Y(n_196)
);

INVx1_ASAP7_75t_SL g286 ( 
.A(n_196),
.Y(n_286)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_139),
.Y(n_197)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_197),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_156),
.B(n_96),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_152),
.B(n_132),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_199),
.B(n_200),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_135),
.B(n_102),
.Y(n_200)
);

INVx4_ASAP7_75t_L g201 ( 
.A(n_117),
.Y(n_201)
);

HB1xp67_ASAP7_75t_L g249 ( 
.A(n_201),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_147),
.B(n_105),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_202),
.B(n_225),
.Y(n_283)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_148),
.Y(n_204)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_204),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_SL g205 ( 
.A1(n_163),
.A2(n_128),
.B(n_158),
.Y(n_205)
);

AOI21xp5_ASAP7_75t_L g274 ( 
.A1(n_205),
.A2(n_230),
.B(n_238),
.Y(n_274)
);

INVx4_ASAP7_75t_L g206 ( 
.A(n_124),
.Y(n_206)
);

HB1xp67_ASAP7_75t_L g263 ( 
.A(n_206),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_169),
.B(n_115),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_207),
.B(n_209),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_174),
.A2(n_112),
.B1(n_87),
.B2(n_89),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_208),
.A2(n_137),
.B1(n_138),
.B2(n_134),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_153),
.B(n_98),
.Y(n_209)
);

INVx3_ASAP7_75t_L g210 ( 
.A(n_126),
.Y(n_210)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_210),
.Y(n_264)
);

CKINVDCx16_ASAP7_75t_R g211 ( 
.A(n_163),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_211),
.B(n_219),
.Y(n_293)
);

OAI22xp33_ASAP7_75t_SL g256 ( 
.A1(n_213),
.A2(n_216),
.B1(n_241),
.B2(n_245),
.Y(n_256)
);

INVx6_ASAP7_75t_L g214 ( 
.A(n_143),
.Y(n_214)
);

INVx8_ASAP7_75t_L g292 ( 
.A(n_214),
.Y(n_292)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_171),
.Y(n_215)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_215),
.Y(n_265)
);

AOI22xp33_ASAP7_75t_L g216 ( 
.A1(n_180),
.A2(n_142),
.B1(n_168),
.B2(n_165),
.Y(n_216)
);

INVx8_ASAP7_75t_L g217 ( 
.A(n_181),
.Y(n_217)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_217),
.Y(n_270)
);

INVx3_ASAP7_75t_L g218 ( 
.A(n_140),
.Y(n_218)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_218),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_186),
.B(n_111),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_120),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_220),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_SL g222 ( 
.A(n_183),
.B(n_6),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_222),
.B(n_228),
.Y(n_285)
);

BUFx8_ASAP7_75t_L g223 ( 
.A(n_150),
.Y(n_223)
);

BUFx2_ASAP7_75t_SL g288 ( 
.A(n_223),
.Y(n_288)
);

AOI22xp33_ASAP7_75t_SL g224 ( 
.A1(n_179),
.A2(n_94),
.B1(n_59),
.B2(n_68),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_224),
.A2(n_231),
.B1(n_232),
.B2(n_233),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_184),
.B(n_6),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_153),
.B(n_70),
.Y(n_226)
);

CKINVDCx16_ASAP7_75t_R g291 ( 
.A(n_226),
.Y(n_291)
);

BUFx6f_ASAP7_75t_L g227 ( 
.A(n_143),
.Y(n_227)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_227),
.Y(n_289)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_164),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_134),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_229),
.Y(n_278)
);

OAI21xp5_ASAP7_75t_L g230 ( 
.A1(n_144),
.A2(n_159),
.B(n_136),
.Y(n_230)
);

INVx4_ASAP7_75t_L g231 ( 
.A(n_140),
.Y(n_231)
);

NOR3xp33_ASAP7_75t_L g232 ( 
.A(n_150),
.B(n_81),
.C(n_9),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_162),
.B(n_8),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_173),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_234),
.B(n_236),
.C(n_237),
.Y(n_266)
);

BUFx6f_ASAP7_75t_L g235 ( 
.A(n_141),
.Y(n_235)
);

AOI22xp33_ASAP7_75t_L g255 ( 
.A1(n_235),
.A2(n_242),
.B1(n_243),
.B2(n_123),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_154),
.B(n_8),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_167),
.B(n_10),
.Y(n_237)
);

INVx1_ASAP7_75t_SL g238 ( 
.A(n_181),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_185),
.B(n_11),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_239),
.B(n_240),
.C(n_246),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_151),
.B(n_11),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_170),
.B(n_12),
.Y(n_241)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_151),
.Y(n_242)
);

AOI22xp33_ASAP7_75t_SL g245 ( 
.A1(n_179),
.A2(n_12),
.B1(n_14),
.B2(n_176),
.Y(n_245)
);

NAND2x1_ASAP7_75t_SL g246 ( 
.A(n_123),
.B(n_12),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_251),
.A2(n_257),
.B1(n_259),
.B2(n_268),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_212),
.A2(n_121),
.B1(n_130),
.B2(n_155),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_L g324 ( 
.A1(n_253),
.A2(n_254),
.B1(n_258),
.B2(n_261),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_208),
.A2(n_121),
.B1(n_130),
.B2(n_155),
.Y(n_254)
);

INVxp33_ASAP7_75t_L g326 ( 
.A(n_255),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_213),
.A2(n_239),
.B1(n_230),
.B2(n_221),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_190),
.A2(n_127),
.B1(n_149),
.B2(n_172),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_L g259 ( 
.A1(n_221),
.A2(n_141),
.B1(n_157),
.B2(n_175),
.Y(n_259)
);

AOI22xp33_ASAP7_75t_L g261 ( 
.A1(n_198),
.A2(n_127),
.B1(n_149),
.B2(n_157),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_221),
.A2(n_175),
.B1(n_181),
.B2(n_191),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_192),
.A2(n_200),
.B1(n_202),
.B2(n_225),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_271),
.A2(n_281),
.B1(n_246),
.B2(n_201),
.Y(n_294)
);

AOI22xp33_ASAP7_75t_L g272 ( 
.A1(n_237),
.A2(n_240),
.B1(n_229),
.B2(n_228),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_272),
.A2(n_273),
.B1(n_279),
.B2(n_280),
.Y(n_298)
);

AOI22xp33_ASAP7_75t_L g273 ( 
.A1(n_197),
.A2(n_242),
.B1(n_215),
.B2(n_204),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_194),
.A2(n_244),
.B1(n_243),
.B2(n_199),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_244),
.A2(n_243),
.B1(n_189),
.B2(n_235),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_243),
.A2(n_205),
.B1(n_214),
.B2(n_227),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_238),
.B(n_218),
.C(n_210),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_282),
.B(n_274),
.C(n_250),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_SL g341 ( 
.A1(n_294),
.A2(n_267),
.B1(n_270),
.B2(n_292),
.Y(n_341)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_262),
.Y(n_295)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_295),
.Y(n_339)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_262),
.Y(n_296)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_296),
.Y(n_347)
);

OAI21xp5_ASAP7_75t_L g297 ( 
.A1(n_248),
.A2(n_223),
.B(n_217),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_SL g337 ( 
.A1(n_297),
.A2(n_325),
.B(n_267),
.Y(n_337)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_265),
.Y(n_299)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_299),
.Y(n_352)
);

INVx1_ASAP7_75t_SL g300 ( 
.A(n_288),
.Y(n_300)
);

BUFx3_ASAP7_75t_L g345 ( 
.A(n_300),
.Y(n_345)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_289),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_301),
.B(n_302),
.Y(n_344)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_289),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_291),
.B(n_187),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_SL g335 ( 
.A(n_303),
.B(n_307),
.Y(n_335)
);

A2O1A1Ixp33_ASAP7_75t_L g304 ( 
.A1(n_257),
.A2(n_223),
.B(n_206),
.C(n_231),
.Y(n_304)
);

OAI21xp5_ASAP7_75t_L g346 ( 
.A1(n_304),
.A2(n_316),
.B(n_318),
.Y(n_346)
);

INVx3_ASAP7_75t_L g305 ( 
.A(n_288),
.Y(n_305)
);

AOI22xp33_ASAP7_75t_SL g343 ( 
.A1(n_305),
.A2(n_327),
.B1(n_328),
.B2(n_286),
.Y(n_343)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_265),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_306),
.B(n_315),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_291),
.B(n_196),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_252),
.B(n_247),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_308),
.B(n_311),
.Y(n_354)
);

OAI22xp5_ASAP7_75t_SL g309 ( 
.A1(n_280),
.A2(n_279),
.B1(n_253),
.B2(n_258),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_L g333 ( 
.A1(n_309),
.A2(n_314),
.B1(n_275),
.B2(n_278),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_252),
.B(n_247),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_271),
.B(n_283),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_312),
.B(n_313),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_284),
.B(n_290),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_248),
.A2(n_274),
.B1(n_293),
.B2(n_283),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_269),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_284),
.B(n_290),
.Y(n_316)
);

INVxp67_ASAP7_75t_L g317 ( 
.A(n_293),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g330 ( 
.A(n_317),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_285),
.B(n_260),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_249),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_319),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_266),
.B(n_276),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_SL g350 ( 
.A(n_320),
.B(n_323),
.Y(n_350)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_263),
.Y(n_321)
);

AOI22xp33_ASAP7_75t_L g338 ( 
.A1(n_321),
.A2(n_286),
.B1(n_287),
.B2(n_264),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_322),
.B(n_275),
.C(n_282),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_SL g323 ( 
.A(n_266),
.B(n_268),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_285),
.B(n_260),
.Y(n_325)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_269),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_264),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_276),
.B(n_278),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_L g348 ( 
.A(n_329),
.B(n_292),
.Y(n_348)
);

AOI21xp5_ASAP7_75t_L g331 ( 
.A1(n_297),
.A2(n_281),
.B(n_256),
.Y(n_331)
);

AOI21xp5_ASAP7_75t_L g376 ( 
.A1(n_331),
.A2(n_300),
.B(n_305),
.Y(n_376)
);

OAI22xp5_ASAP7_75t_L g332 ( 
.A1(n_310),
.A2(n_254),
.B1(n_259),
.B2(n_251),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_L g370 ( 
.A1(n_332),
.A2(n_333),
.B1(n_338),
.B2(n_295),
.Y(n_370)
);

MAJIxp5_ASAP7_75t_L g361 ( 
.A(n_334),
.B(n_336),
.C(n_356),
.Y(n_361)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_320),
.B(n_277),
.C(n_270),
.Y(n_336)
);

INVxp67_ASAP7_75t_L g366 ( 
.A(n_337),
.Y(n_366)
);

INVxp67_ASAP7_75t_L g375 ( 
.A(n_341),
.Y(n_375)
);

OAI21xp5_ASAP7_75t_SL g342 ( 
.A1(n_294),
.A2(n_277),
.B(n_287),
.Y(n_342)
);

AO21x1_ASAP7_75t_L g360 ( 
.A1(n_342),
.A2(n_351),
.B(n_326),
.Y(n_360)
);

HB1xp67_ASAP7_75t_L g377 ( 
.A(n_343),
.Y(n_377)
);

XNOR2xp5_ASAP7_75t_SL g367 ( 
.A(n_348),
.B(n_355),
.Y(n_367)
);

OAI22xp5_ASAP7_75t_SL g349 ( 
.A1(n_310),
.A2(n_292),
.B1(n_312),
.B2(n_311),
.Y(n_349)
);

AOI22xp5_ASAP7_75t_L g380 ( 
.A1(n_349),
.A2(n_306),
.B1(n_301),
.B2(n_302),
.Y(n_380)
);

AO21x2_ASAP7_75t_SL g351 ( 
.A1(n_309),
.A2(n_324),
.B(n_304),
.Y(n_351)
);

XNOR2xp5_ASAP7_75t_L g355 ( 
.A(n_308),
.B(n_329),
.Y(n_355)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_323),
.B(n_322),
.C(n_314),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_SL g358 ( 
.A(n_330),
.B(n_318),
.Y(n_358)
);

CKINVDCx14_ASAP7_75t_R g390 ( 
.A(n_358),
.Y(n_390)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_353),
.Y(n_359)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_359),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_360),
.B(n_376),
.Y(n_400)
);

XNOR2xp5_ASAP7_75t_L g362 ( 
.A(n_355),
.B(n_316),
.Y(n_362)
);

MAJIxp5_ASAP7_75t_L g386 ( 
.A(n_362),
.B(n_363),
.C(n_381),
.Y(n_386)
);

MAJIxp5_ASAP7_75t_L g363 ( 
.A(n_356),
.B(n_313),
.C(n_304),
.Y(n_363)
);

OAI22xp5_ASAP7_75t_SL g364 ( 
.A1(n_351),
.A2(n_298),
.B1(n_325),
.B2(n_324),
.Y(n_364)
);

AOI22xp5_ASAP7_75t_L g383 ( 
.A1(n_364),
.A2(n_370),
.B1(n_351),
.B2(n_349),
.Y(n_383)
);

OAI21xp5_ASAP7_75t_L g365 ( 
.A1(n_337),
.A2(n_303),
.B(n_307),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_L g384 ( 
.A(n_365),
.B(n_368),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_L g368 ( 
.A(n_330),
.B(n_321),
.Y(n_368)
);

BUFx24_ASAP7_75t_SL g369 ( 
.A(n_357),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_L g387 ( 
.A(n_369),
.B(n_371),
.Y(n_387)
);

XOR2x2_ASAP7_75t_L g371 ( 
.A(n_357),
.B(n_298),
.Y(n_371)
);

OAI22xp5_ASAP7_75t_L g372 ( 
.A1(n_333),
.A2(n_296),
.B1(n_319),
.B2(n_299),
.Y(n_372)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_372),
.Y(n_399)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_353),
.Y(n_373)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_373),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_SL g374 ( 
.A(n_354),
.B(n_328),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_L g395 ( 
.A(n_374),
.B(n_373),
.Y(n_395)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_339),
.Y(n_378)
);

INVx2_ASAP7_75t_L g391 ( 
.A(n_378),
.Y(n_391)
);

OR2x2_ASAP7_75t_L g379 ( 
.A(n_346),
.B(n_335),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_SL g385 ( 
.A(n_379),
.B(n_346),
.Y(n_385)
);

OAI22xp5_ASAP7_75t_SL g392 ( 
.A1(n_380),
.A2(n_339),
.B1(n_347),
.B2(n_378),
.Y(n_392)
);

MAJIxp5_ASAP7_75t_L g381 ( 
.A(n_350),
.B(n_315),
.C(n_327),
.Y(n_381)
);

CKINVDCx20_ASAP7_75t_R g382 ( 
.A(n_379),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_382),
.B(n_397),
.Y(n_408)
);

AOI22xp5_ASAP7_75t_L g411 ( 
.A1(n_383),
.A2(n_389),
.B1(n_392),
.B2(n_396),
.Y(n_411)
);

OR2x2_ASAP7_75t_L g414 ( 
.A(n_385),
.B(n_394),
.Y(n_414)
);

INVx5_ASAP7_75t_L g388 ( 
.A(n_371),
.Y(n_388)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_388),
.Y(n_419)
);

OAI22xp5_ASAP7_75t_L g389 ( 
.A1(n_375),
.A2(n_351),
.B1(n_331),
.B2(n_354),
.Y(n_389)
);

MAJIxp5_ASAP7_75t_L g393 ( 
.A(n_361),
.B(n_334),
.C(n_336),
.Y(n_393)
);

MAJIxp5_ASAP7_75t_L g417 ( 
.A(n_393),
.B(n_363),
.C(n_367),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_SL g394 ( 
.A(n_359),
.B(n_335),
.Y(n_394)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_395),
.Y(n_404)
);

AOI22xp5_ASAP7_75t_L g396 ( 
.A1(n_364),
.A2(n_351),
.B1(n_341),
.B2(n_332),
.Y(n_396)
);

CKINVDCx20_ASAP7_75t_R g397 ( 
.A(n_376),
.Y(n_397)
);

CKINVDCx20_ASAP7_75t_R g401 ( 
.A(n_380),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_401),
.B(n_360),
.Y(n_418)
);

XOR2x2_ASAP7_75t_SL g403 ( 
.A(n_389),
.B(n_350),
.Y(n_403)
);

MAJIxp5_ASAP7_75t_L g424 ( 
.A(n_403),
.B(n_409),
.C(n_416),
.Y(n_424)
);

XNOR2xp5_ASAP7_75t_L g405 ( 
.A(n_393),
.B(n_361),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_L g421 ( 
.A(n_405),
.B(n_410),
.Y(n_421)
);

OAI21xp5_ASAP7_75t_L g406 ( 
.A1(n_400),
.A2(n_366),
.B(n_375),
.Y(n_406)
);

OAI21xp5_ASAP7_75t_SL g426 ( 
.A1(n_406),
.A2(n_400),
.B(n_397),
.Y(n_426)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_395),
.Y(n_407)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_407),
.Y(n_431)
);

XOR2xp5_ASAP7_75t_L g409 ( 
.A(n_386),
.B(n_381),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_398),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_L g412 ( 
.A(n_382),
.B(n_362),
.Y(n_412)
);

CKINVDCx16_ASAP7_75t_R g420 ( 
.A(n_412),
.Y(n_420)
);

INVxp33_ASAP7_75t_L g413 ( 
.A(n_394),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_413),
.B(n_418),
.Y(n_432)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_398),
.Y(n_415)
);

NOR2xp33_ASAP7_75t_L g422 ( 
.A(n_415),
.B(n_340),
.Y(n_422)
);

XOR2x2_ASAP7_75t_SL g416 ( 
.A(n_385),
.B(n_367),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_SL g423 ( 
.A(n_417),
.B(n_386),
.Y(n_423)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_422),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_SL g441 ( 
.A(n_423),
.B(n_348),
.Y(n_441)
);

OAI22xp5_ASAP7_75t_L g425 ( 
.A1(n_414),
.A2(n_390),
.B1(n_387),
.B2(n_383),
.Y(n_425)
);

OAI22xp5_ASAP7_75t_L g439 ( 
.A1(n_425),
.A2(n_429),
.B1(n_399),
.B2(n_402),
.Y(n_439)
);

AOI21xp5_ASAP7_75t_L g438 ( 
.A1(n_426),
.A2(n_428),
.B(n_430),
.Y(n_438)
);

BUFx2_ASAP7_75t_L g427 ( 
.A(n_404),
.Y(n_427)
);

CKINVDCx20_ASAP7_75t_R g443 ( 
.A(n_427),
.Y(n_443)
);

OAI21xp5_ASAP7_75t_SL g428 ( 
.A1(n_419),
.A2(n_388),
.B(n_384),
.Y(n_428)
);

AOI22xp5_ASAP7_75t_L g429 ( 
.A1(n_411),
.A2(n_396),
.B1(n_399),
.B2(n_401),
.Y(n_429)
);

OAI21xp5_ASAP7_75t_SL g430 ( 
.A1(n_419),
.A2(n_384),
.B(n_366),
.Y(n_430)
);

OAI22xp5_ASAP7_75t_SL g433 ( 
.A1(n_411),
.A2(n_414),
.B1(n_413),
.B2(n_408),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_433),
.B(n_408),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_434),
.B(n_435),
.Y(n_446)
);

NOR2xp33_ASAP7_75t_L g435 ( 
.A(n_420),
.B(n_387),
.Y(n_435)
);

MAJIxp5_ASAP7_75t_L g437 ( 
.A(n_421),
.B(n_405),
.C(n_409),
.Y(n_437)
);

NOR2xp33_ASAP7_75t_L g445 ( 
.A(n_437),
.B(n_440),
.Y(n_445)
);

AOI22xp5_ASAP7_75t_L g451 ( 
.A1(n_439),
.A2(n_432),
.B1(n_418),
.B2(n_429),
.Y(n_451)
);

MAJIxp5_ASAP7_75t_L g440 ( 
.A(n_424),
.B(n_417),
.C(n_403),
.Y(n_440)
);

XNOR2xp5_ASAP7_75t_L g452 ( 
.A(n_441),
.B(n_365),
.Y(n_452)
);

MAJIxp5_ASAP7_75t_L g442 ( 
.A(n_424),
.B(n_406),
.C(n_416),
.Y(n_442)
);

NOR2xp33_ASAP7_75t_L g447 ( 
.A(n_442),
.B(n_428),
.Y(n_447)
);

AOI22xp33_ASAP7_75t_SL g444 ( 
.A1(n_436),
.A2(n_433),
.B1(n_431),
.B2(n_427),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_444),
.B(n_447),
.Y(n_457)
);

NOR2xp33_ASAP7_75t_L g448 ( 
.A(n_443),
.B(n_430),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_448),
.B(n_449),
.Y(n_459)
);

CKINVDCx20_ASAP7_75t_R g449 ( 
.A(n_434),
.Y(n_449)
);

NOR2xp33_ASAP7_75t_L g450 ( 
.A(n_437),
.B(n_402),
.Y(n_450)
);

NAND3xp33_ASAP7_75t_L g453 ( 
.A(n_450),
.B(n_438),
.C(n_442),
.Y(n_453)
);

NOR2xp33_ASAP7_75t_L g456 ( 
.A(n_451),
.B(n_432),
.Y(n_456)
);

NOR2xp33_ASAP7_75t_L g454 ( 
.A(n_452),
.B(n_446),
.Y(n_454)
);

AOI21xp5_ASAP7_75t_L g462 ( 
.A1(n_453),
.A2(n_458),
.B(n_438),
.Y(n_462)
);

XNOR2xp5_ASAP7_75t_SL g461 ( 
.A(n_454),
.B(n_452),
.Y(n_461)
);

AND2x2_ASAP7_75t_L g455 ( 
.A(n_445),
.B(n_440),
.Y(n_455)
);

AO21x1_ASAP7_75t_L g463 ( 
.A1(n_455),
.A2(n_426),
.B(n_451),
.Y(n_463)
);

INVxp67_ASAP7_75t_L g460 ( 
.A(n_456),
.Y(n_460)
);

INVx11_ASAP7_75t_L g458 ( 
.A(n_446),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_461),
.B(n_462),
.Y(n_467)
);

AOI22xp5_ASAP7_75t_SL g465 ( 
.A1(n_463),
.A2(n_457),
.B1(n_456),
.B2(n_340),
.Y(n_465)
);

XOR2xp5_ASAP7_75t_L g464 ( 
.A(n_459),
.B(n_377),
.Y(n_464)
);

AO221x1_ASAP7_75t_L g466 ( 
.A1(n_464),
.A2(n_391),
.B1(n_392),
.B2(n_344),
.C(n_360),
.Y(n_466)
);

OAI321xp33_ASAP7_75t_L g469 ( 
.A1(n_465),
.A2(n_347),
.A3(n_352),
.B1(n_344),
.B2(n_391),
.C(n_300),
.Y(n_469)
);

AOI21xp5_ASAP7_75t_L g468 ( 
.A1(n_466),
.A2(n_460),
.B(n_342),
.Y(n_468)
);

MAJIxp5_ASAP7_75t_L g470 ( 
.A(n_468),
.B(n_469),
.C(n_467),
.Y(n_470)
);

AOI21xp5_ASAP7_75t_L g471 ( 
.A1(n_470),
.A2(n_352),
.B(n_305),
.Y(n_471)
);

NAND3xp33_ASAP7_75t_L g472 ( 
.A(n_471),
.B(n_345),
.C(n_453),
.Y(n_472)
);

XOR2xp5_ASAP7_75t_L g473 ( 
.A(n_472),
.B(n_345),
.Y(n_473)
);


endmodule