module fake_jpeg_21648_n_105 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_8, n_15, n_7, n_105);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_8;
input n_15;
input n_7;

output n_105;

wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_44;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

BUFx24_ASAP7_75t_L g32 ( 
.A(n_28),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_27),
.Y(n_33)
);

INVx5_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_18),
.B(n_15),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_12),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_17),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_29),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_16),
.Y(n_39)
);

INVx2_ASAP7_75t_SL g40 ( 
.A(n_2),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_2),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_22),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_11),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_3),
.Y(n_45)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_32),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_46),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_32),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_47),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_39),
.Y(n_48)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_48),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_39),
.Y(n_49)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_49),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_SL g50 ( 
.A(n_40),
.B(n_0),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_50),
.B(n_51),
.Y(n_59)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_41),
.Y(n_51)
);

BUFx5_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_52),
.Y(n_54)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_34),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_53),
.B(n_0),
.Y(n_65)
);

NOR2x1_ASAP7_75t_L g57 ( 
.A(n_50),
.B(n_45),
.Y(n_57)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_57),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_51),
.B(n_44),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_58),
.B(n_60),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g60 ( 
.A(n_51),
.B(n_44),
.C(n_42),
.Y(n_60)
);

OAI22xp33_ASAP7_75t_L g62 ( 
.A1(n_53),
.A2(n_43),
.B1(n_38),
.B2(n_36),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_62),
.A2(n_63),
.B1(n_35),
.B2(n_20),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_46),
.A2(n_33),
.B1(n_21),
.B2(n_30),
.Y(n_63)
);

CKINVDCx16_ASAP7_75t_R g67 ( 
.A(n_65),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_68),
.B(n_70),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_59),
.A2(n_63),
.B1(n_65),
.B2(n_56),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_69),
.A2(n_72),
.B1(n_10),
.B2(n_13),
.Y(n_89)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_61),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_54),
.Y(n_71)
);

OR2x2_ASAP7_75t_L g82 ( 
.A(n_71),
.B(n_4),
.Y(n_82)
);

O2A1O1Ixp33_ASAP7_75t_L g72 ( 
.A1(n_59),
.A2(n_19),
.B(n_26),
.C(n_25),
.Y(n_72)
);

CKINVDCx16_ASAP7_75t_R g74 ( 
.A(n_54),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_74),
.B(n_77),
.Y(n_85)
);

INVx5_ASAP7_75t_L g75 ( 
.A(n_64),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_75),
.Y(n_86)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_55),
.Y(n_76)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_76),
.Y(n_84)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_54),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_58),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_78),
.A2(n_79),
.B1(n_1),
.B2(n_3),
.Y(n_80)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_58),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_80),
.B(n_82),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_L g83 ( 
.A1(n_76),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_83)
);

OR2x2_ASAP7_75t_L g93 ( 
.A(n_83),
.B(n_87),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_L g87 ( 
.A1(n_67),
.A2(n_5),
.B1(n_7),
.B2(n_8),
.Y(n_87)
);

XNOR2xp5_ASAP7_75t_L g88 ( 
.A(n_73),
.B(n_9),
.Y(n_88)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_88),
.Y(n_90)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_89),
.Y(n_91)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_85),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_92),
.B(n_66),
.C(n_81),
.Y(n_95)
);

XOR2xp5_ASAP7_75t_L g97 ( 
.A(n_95),
.B(n_96),
.Y(n_97)
);

A2O1A1O1Ixp25_ASAP7_75t_L g96 ( 
.A1(n_90),
.A2(n_72),
.B(n_87),
.C(n_83),
.D(n_24),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_97),
.B(n_94),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_98),
.B(n_91),
.C(n_93),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_99),
.A2(n_93),
.B1(n_84),
.B2(n_77),
.Y(n_100)
);

BUFx24_ASAP7_75t_SL g101 ( 
.A(n_100),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_L g102 ( 
.A(n_101),
.B(n_14),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_102),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_103),
.B(n_86),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_104),
.B(n_23),
.Y(n_105)
);


endmodule