module fake_netlist_6_1108_n_1919 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_193, n_147, n_154, n_191, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_166, n_28, n_184, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_188, n_102, n_186, n_0, n_87, n_195, n_189, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_104, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_190, n_14, n_123, n_136, n_72, n_187, n_89, n_173, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_194, n_171, n_31, n_192, n_57, n_169, n_53, n_51, n_44, n_56, n_1919);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_193;
input n_147;
input n_154;
input n_191;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_184;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_188;
input n_102;
input n_186;
input n_0;
input n_87;
input n_195;
input n_189;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_104;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_190;
input n_14;
input n_123;
input n_136;
input n_72;
input n_187;
input n_89;
input n_173;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_194;
input n_171;
input n_31;
input n_192;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1919;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_1853;
wire n_783;
wire n_1738;
wire n_798;
wire n_1575;
wire n_1854;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1691;
wire n_1688;
wire n_1009;
wire n_1743;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_1844;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1803;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1867;
wire n_1704;
wire n_1078;
wire n_250;
wire n_544;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1903;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_658;
wire n_616;
wire n_1874;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1560;
wire n_1526;
wire n_734;
wire n_1088;
wire n_1894;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_1815;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1911;
wire n_1644;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_1918;
wire n_577;
wire n_1843;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1909;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_1907;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1876;
wire n_1895;
wire n_1697;
wire n_243;
wire n_979;
wire n_1873;
wire n_905;
wire n_1866;
wire n_1680;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1605;
wire n_1413;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1865;
wire n_1875;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_530;
wire n_1563;
wire n_1912;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_210;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_1896;
wire n_429;
wire n_1747;
wire n_1012;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1802;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_850;
wire n_690;
wire n_1801;
wire n_1886;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_697;
wire n_687;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_484;
wire n_1709;
wire n_1825;
wire n_1757;
wire n_1796;
wire n_1792;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_297;
wire n_627;
wire n_595;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1858;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_1839;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_1863;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_1913;
wire n_510;
wire n_837;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_1788;
wire n_622;
wire n_1469;
wire n_1838;
wire n_1835;
wire n_1776;
wire n_1766;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_1878;
wire n_899;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_1181;
wire n_1822;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_1817;
wire n_927;
wire n_1849;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_552;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_216;
wire n_912;
wire n_1857;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1774;
wire n_884;
wire n_1398;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_1021;
wire n_931;
wire n_474;
wire n_527;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_1897;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_1837;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_211;
wire n_1483;
wire n_1834;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_1877;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1769;
wire n_1220;
wire n_1893;
wire n_556;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_1286;
wire n_1775;
wire n_1773;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_1745;
wire n_914;
wire n_759;
wire n_1831;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_1901;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1892;
wire n_1135;
wire n_1179;
wire n_1169;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1917;
wire n_1580;
wire n_1425;
wire n_1881;
wire n_1267;
wire n_1281;
wire n_1806;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_1855;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_1832;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_1869;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_1889;
wire n_435;
wire n_1905;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_1871;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_1859;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_1916;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_198;
wire n_1847;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1841;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1818;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1262;
wire n_218;
wire n_1891;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_1870;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_1695;
wire n_1828;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1883;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_1823;
wire n_227;
wire n_1720;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_1846;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_1676;
wire n_833;
wire n_1830;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_1900;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1906;
wire n_1484;
wire n_1321;
wire n_1241;
wire n_1672;
wire n_569;
wire n_1758;
wire n_737;
wire n_1318;
wire n_1914;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1794;
wire n_786;
wire n_1650;
wire n_1236;
wire n_1559;
wire n_1725;
wire n_1872;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1741;
wire n_1325;
wire n_1002;
wire n_1746;
wire n_545;
wire n_489;
wire n_1804;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1860;
wire n_1904;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1908;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1800;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1882;
wire n_1076;
wire n_1118;
wire n_1007;
wire n_1807;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_1879;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_1810;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_1729;
wire n_669;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1785;
wire n_763;
wire n_1147;
wire n_1848;
wire n_360;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_1851;
wire n_363;
wire n_1799;
wire n_1090;
wire n_592;
wire n_1816;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_1829;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_404;
wire n_271;
wire n_1884;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1819;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_373;
wire n_1632;
wire n_1890;
wire n_1805;
wire n_257;
wire n_1557;
wire n_1888;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_1850;
wire n_1898;
wire n_1868;
wire n_207;
wire n_1089;
wire n_1887;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_1836;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1899;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1862;
wire n_1856;
wire n_339;
wire n_784;
wire n_434;
wire n_315;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_1915;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1885;
wire n_1013;
wire n_1259;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

INVx2_ASAP7_75t_L g196 ( 
.A(n_112),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_80),
.Y(n_197)
);

BUFx3_ASAP7_75t_L g198 ( 
.A(n_166),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_53),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_70),
.Y(n_200)
);

BUFx10_ASAP7_75t_L g201 ( 
.A(n_131),
.Y(n_201)
);

INVx1_ASAP7_75t_SL g202 ( 
.A(n_81),
.Y(n_202)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_153),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_38),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_184),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_36),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_78),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_3),
.Y(n_208)
);

CKINVDCx11_ASAP7_75t_R g209 ( 
.A(n_36),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_21),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_73),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_187),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_97),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_9),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_139),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_135),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_150),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_47),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_148),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_179),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_158),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_161),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_137),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_114),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_40),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_178),
.Y(n_226)
);

INVxp33_ASAP7_75t_R g227 ( 
.A(n_57),
.Y(n_227)
);

BUFx2_ASAP7_75t_L g228 ( 
.A(n_19),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_188),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_46),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_41),
.Y(n_231)
);

BUFx2_ASAP7_75t_L g232 ( 
.A(n_136),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_121),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_10),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_147),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_88),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_48),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_140),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_102),
.Y(n_239)
);

BUFx2_ASAP7_75t_L g240 ( 
.A(n_82),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_30),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_27),
.Y(n_242)
);

CKINVDCx14_ASAP7_75t_R g243 ( 
.A(n_1),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_165),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_105),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_124),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_8),
.Y(n_247)
);

BUFx6f_ASAP7_75t_L g248 ( 
.A(n_160),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_174),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_94),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_100),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_113),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_86),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_66),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_129),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_28),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_25),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_31),
.Y(n_258)
);

INVx1_ASAP7_75t_SL g259 ( 
.A(n_85),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_1),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_99),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_69),
.Y(n_262)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_190),
.Y(n_263)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_84),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_55),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_91),
.Y(n_266)
);

CKINVDCx16_ASAP7_75t_R g267 ( 
.A(n_96),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_90),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_169),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_108),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_63),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_67),
.Y(n_272)
);

CKINVDCx16_ASAP7_75t_R g273 ( 
.A(n_95),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_117),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_120),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_162),
.Y(n_276)
);

INVxp67_ASAP7_75t_L g277 ( 
.A(n_183),
.Y(n_277)
);

BUFx2_ASAP7_75t_SL g278 ( 
.A(n_171),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_21),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_15),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_173),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_71),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_107),
.Y(n_283)
);

HB1xp67_ASAP7_75t_L g284 ( 
.A(n_43),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_61),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_56),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_29),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_15),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_149),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_144),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_55),
.Y(n_291)
);

INVx1_ASAP7_75t_SL g292 ( 
.A(n_24),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_146),
.Y(n_293)
);

CKINVDCx14_ASAP7_75t_R g294 ( 
.A(n_182),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_68),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_43),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_170),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_185),
.Y(n_298)
);

BUFx6f_ASAP7_75t_L g299 ( 
.A(n_192),
.Y(n_299)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_52),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_56),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_3),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_181),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_128),
.Y(n_304)
);

INVx2_ASAP7_75t_L g305 ( 
.A(n_79),
.Y(n_305)
);

BUFx2_ASAP7_75t_L g306 ( 
.A(n_195),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_83),
.Y(n_307)
);

INVx1_ASAP7_75t_SL g308 ( 
.A(n_14),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_29),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_20),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_13),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_16),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_98),
.Y(n_313)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_157),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_75),
.Y(n_315)
);

CKINVDCx14_ASAP7_75t_R g316 ( 
.A(n_61),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_48),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_125),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_176),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_37),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_172),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_4),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_45),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_133),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_45),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_145),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_52),
.Y(n_327)
);

HB1xp67_ASAP7_75t_L g328 ( 
.A(n_134),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_5),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_5),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_194),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_60),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_40),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_87),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_111),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_35),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_130),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_64),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_23),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_141),
.Y(n_340)
);

INVx1_ASAP7_75t_SL g341 ( 
.A(n_7),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_123),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_167),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_104),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g345 ( 
.A(n_62),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_106),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g347 ( 
.A(n_132),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_116),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_46),
.Y(n_349)
);

INVx2_ASAP7_75t_SL g350 ( 
.A(n_50),
.Y(n_350)
);

BUFx2_ASAP7_75t_L g351 ( 
.A(n_64),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_92),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_2),
.Y(n_353)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_103),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_8),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_127),
.Y(n_356)
);

CKINVDCx20_ASAP7_75t_R g357 ( 
.A(n_62),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_19),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_38),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g360 ( 
.A(n_33),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_13),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_119),
.Y(n_362)
);

CKINVDCx20_ASAP7_75t_R g363 ( 
.A(n_77),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_72),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_28),
.Y(n_365)
);

CKINVDCx16_ASAP7_75t_R g366 ( 
.A(n_175),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_22),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_35),
.Y(n_368)
);

BUFx10_ASAP7_75t_L g369 ( 
.A(n_74),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_189),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_0),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_168),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_186),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_34),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_37),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_138),
.Y(n_376)
);

INVx4_ASAP7_75t_R g377 ( 
.A(n_30),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_154),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_109),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_0),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_118),
.Y(n_381)
);

CKINVDCx16_ASAP7_75t_R g382 ( 
.A(n_152),
.Y(n_382)
);

BUFx8_ASAP7_75t_SL g383 ( 
.A(n_27),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_122),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_159),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_41),
.Y(n_386)
);

BUFx2_ASAP7_75t_L g387 ( 
.A(n_17),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_180),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_177),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_23),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_54),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_65),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_51),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_155),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_89),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_7),
.Y(n_396)
);

CKINVDCx20_ASAP7_75t_R g397 ( 
.A(n_236),
.Y(n_397)
);

INVxp67_ASAP7_75t_L g398 ( 
.A(n_228),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_300),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_243),
.B(n_316),
.Y(n_400)
);

INVxp67_ASAP7_75t_L g401 ( 
.A(n_228),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_300),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_199),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_209),
.Y(n_404)
);

INVxp67_ASAP7_75t_L g405 ( 
.A(n_351),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_383),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_199),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_210),
.Y(n_408)
);

AND2x2_ASAP7_75t_L g409 ( 
.A(n_351),
.B(n_2),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_200),
.Y(n_410)
);

NOR2xp67_ASAP7_75t_L g411 ( 
.A(n_284),
.B(n_4),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_205),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_207),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_212),
.Y(n_414)
);

INVxp33_ASAP7_75t_SL g415 ( 
.A(n_387),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_210),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_231),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_213),
.Y(n_418)
);

CKINVDCx20_ASAP7_75t_R g419 ( 
.A(n_252),
.Y(n_419)
);

INVx2_ASAP7_75t_L g420 ( 
.A(n_211),
.Y(n_420)
);

CKINVDCx20_ASAP7_75t_R g421 ( 
.A(n_269),
.Y(n_421)
);

CKINVDCx20_ASAP7_75t_R g422 ( 
.A(n_272),
.Y(n_422)
);

INVxp67_ASAP7_75t_L g423 ( 
.A(n_387),
.Y(n_423)
);

NOR2xp33_ASAP7_75t_L g424 ( 
.A(n_232),
.B(n_6),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_215),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_216),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_217),
.Y(n_427)
);

INVx2_ASAP7_75t_L g428 ( 
.A(n_211),
.Y(n_428)
);

NOR2xp33_ASAP7_75t_L g429 ( 
.A(n_232),
.B(n_6),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_222),
.Y(n_430)
);

INVxp67_ASAP7_75t_L g431 ( 
.A(n_231),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_247),
.Y(n_432)
);

HB1xp67_ASAP7_75t_L g433 ( 
.A(n_204),
.Y(n_433)
);

INVx3_ASAP7_75t_L g434 ( 
.A(n_198),
.Y(n_434)
);

CKINVDCx20_ASAP7_75t_R g435 ( 
.A(n_293),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_247),
.Y(n_436)
);

INVxp67_ASAP7_75t_L g437 ( 
.A(n_286),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_223),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_224),
.Y(n_439)
);

CKINVDCx20_ASAP7_75t_R g440 ( 
.A(n_347),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_229),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_286),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_287),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_287),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_235),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_238),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_288),
.Y(n_447)
);

CKINVDCx20_ASAP7_75t_R g448 ( 
.A(n_363),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_288),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_249),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_317),
.Y(n_451)
);

NOR2xp33_ASAP7_75t_R g452 ( 
.A(n_294),
.B(n_193),
.Y(n_452)
);

BUFx2_ASAP7_75t_L g453 ( 
.A(n_206),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_317),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_325),
.Y(n_455)
);

CKINVDCx20_ASAP7_75t_R g456 ( 
.A(n_267),
.Y(n_456)
);

CKINVDCx20_ASAP7_75t_R g457 ( 
.A(n_273),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_325),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_250),
.Y(n_459)
);

HB1xp67_ASAP7_75t_L g460 ( 
.A(n_208),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_327),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_327),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_333),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_333),
.Y(n_464)
);

CKINVDCx5p33_ASAP7_75t_R g465 ( 
.A(n_251),
.Y(n_465)
);

NOR2xp33_ASAP7_75t_L g466 ( 
.A(n_240),
.B(n_9),
.Y(n_466)
);

CKINVDCx5p33_ASAP7_75t_R g467 ( 
.A(n_253),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_338),
.Y(n_468)
);

CKINVDCx5p33_ASAP7_75t_R g469 ( 
.A(n_254),
.Y(n_469)
);

INVxp67_ASAP7_75t_L g470 ( 
.A(n_338),
.Y(n_470)
);

CKINVDCx20_ASAP7_75t_R g471 ( 
.A(n_366),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_339),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_339),
.Y(n_473)
);

CKINVDCx5p33_ASAP7_75t_R g474 ( 
.A(n_255),
.Y(n_474)
);

INVxp67_ASAP7_75t_L g475 ( 
.A(n_349),
.Y(n_475)
);

CKINVDCx5p33_ASAP7_75t_R g476 ( 
.A(n_268),
.Y(n_476)
);

CKINVDCx5p33_ASAP7_75t_R g477 ( 
.A(n_270),
.Y(n_477)
);

CKINVDCx20_ASAP7_75t_R g478 ( 
.A(n_382),
.Y(n_478)
);

CKINVDCx5p33_ASAP7_75t_R g479 ( 
.A(n_274),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_349),
.Y(n_480)
);

BUFx3_ASAP7_75t_L g481 ( 
.A(n_198),
.Y(n_481)
);

INVxp67_ASAP7_75t_SL g482 ( 
.A(n_328),
.Y(n_482)
);

CKINVDCx5p33_ASAP7_75t_R g483 ( 
.A(n_275),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_359),
.Y(n_484)
);

INVxp67_ASAP7_75t_SL g485 ( 
.A(n_240),
.Y(n_485)
);

NOR2xp33_ASAP7_75t_L g486 ( 
.A(n_306),
.B(n_10),
.Y(n_486)
);

INVxp67_ASAP7_75t_SL g487 ( 
.A(n_306),
.Y(n_487)
);

CKINVDCx5p33_ASAP7_75t_R g488 ( 
.A(n_276),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_359),
.Y(n_489)
);

INVxp67_ASAP7_75t_SL g490 ( 
.A(n_277),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_367),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_196),
.B(n_11),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_367),
.Y(n_493)
);

INVx2_ASAP7_75t_L g494 ( 
.A(n_219),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_368),
.Y(n_495)
);

CKINVDCx20_ASAP7_75t_R g496 ( 
.A(n_282),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_368),
.Y(n_497)
);

INVxp67_ASAP7_75t_L g498 ( 
.A(n_374),
.Y(n_498)
);

CKINVDCx5p33_ASAP7_75t_R g499 ( 
.A(n_289),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_410),
.B(n_196),
.Y(n_500)
);

CKINVDCx5p33_ASAP7_75t_R g501 ( 
.A(n_496),
.Y(n_501)
);

INVx2_ASAP7_75t_L g502 ( 
.A(n_420),
.Y(n_502)
);

CKINVDCx20_ASAP7_75t_R g503 ( 
.A(n_397),
.Y(n_503)
);

CKINVDCx20_ASAP7_75t_R g504 ( 
.A(n_419),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_420),
.Y(n_505)
);

INVx2_ASAP7_75t_L g506 ( 
.A(n_428),
.Y(n_506)
);

HB1xp67_ASAP7_75t_L g507 ( 
.A(n_433),
.Y(n_507)
);

BUFx6f_ASAP7_75t_L g508 ( 
.A(n_428),
.Y(n_508)
);

HB1xp67_ASAP7_75t_L g509 ( 
.A(n_460),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_SL g510 ( 
.A(n_400),
.B(n_201),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_494),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_494),
.Y(n_512)
);

INVx2_ASAP7_75t_L g513 ( 
.A(n_399),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_481),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_481),
.Y(n_515)
);

CKINVDCx5p33_ASAP7_75t_R g516 ( 
.A(n_412),
.Y(n_516)
);

CKINVDCx8_ASAP7_75t_R g517 ( 
.A(n_406),
.Y(n_517)
);

NOR2xp33_ASAP7_75t_L g518 ( 
.A(n_485),
.B(n_202),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_403),
.Y(n_519)
);

INVxp67_ASAP7_75t_L g520 ( 
.A(n_453),
.Y(n_520)
);

NAND2xp33_ASAP7_75t_SL g521 ( 
.A(n_409),
.B(n_350),
.Y(n_521)
);

NOR2xp67_ASAP7_75t_L g522 ( 
.A(n_499),
.B(n_197),
.Y(n_522)
);

BUFx6f_ASAP7_75t_L g523 ( 
.A(n_399),
.Y(n_523)
);

AND2x4_ASAP7_75t_L g524 ( 
.A(n_434),
.B(n_203),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_403),
.Y(n_525)
);

CKINVDCx5p33_ASAP7_75t_R g526 ( 
.A(n_413),
.Y(n_526)
);

CKINVDCx5p33_ASAP7_75t_R g527 ( 
.A(n_414),
.Y(n_527)
);

CKINVDCx20_ASAP7_75t_R g528 ( 
.A(n_421),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_407),
.Y(n_529)
);

OAI22xp5_ASAP7_75t_SL g530 ( 
.A1(n_415),
.A2(n_230),
.B1(n_242),
.B2(n_280),
.Y(n_530)
);

BUFx10_ASAP7_75t_L g531 ( 
.A(n_418),
.Y(n_531)
);

CKINVDCx5p33_ASAP7_75t_R g532 ( 
.A(n_425),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_407),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_408),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_408),
.Y(n_535)
);

AND2x2_ASAP7_75t_L g536 ( 
.A(n_487),
.B(n_434),
.Y(n_536)
);

OAI21x1_ASAP7_75t_L g537 ( 
.A1(n_492),
.A2(n_263),
.B(n_203),
.Y(n_537)
);

CKINVDCx5p33_ASAP7_75t_R g538 ( 
.A(n_426),
.Y(n_538)
);

INVx3_ASAP7_75t_L g539 ( 
.A(n_402),
.Y(n_539)
);

CKINVDCx5p33_ASAP7_75t_R g540 ( 
.A(n_427),
.Y(n_540)
);

CKINVDCx20_ASAP7_75t_R g541 ( 
.A(n_422),
.Y(n_541)
);

AND2x4_ASAP7_75t_L g542 ( 
.A(n_434),
.B(n_263),
.Y(n_542)
);

AND2x6_ASAP7_75t_L g543 ( 
.A(n_409),
.B(n_248),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_416),
.Y(n_544)
);

BUFx6f_ASAP7_75t_L g545 ( 
.A(n_402),
.Y(n_545)
);

INVx3_ASAP7_75t_L g546 ( 
.A(n_416),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_417),
.Y(n_547)
);

CKINVDCx5p33_ASAP7_75t_R g548 ( 
.A(n_430),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_417),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_432),
.Y(n_550)
);

CKINVDCx5p33_ASAP7_75t_R g551 ( 
.A(n_438),
.Y(n_551)
);

INVx2_ASAP7_75t_L g552 ( 
.A(n_432),
.Y(n_552)
);

AND2x6_ASAP7_75t_L g553 ( 
.A(n_424),
.B(n_248),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_436),
.Y(n_554)
);

CKINVDCx5p33_ASAP7_75t_R g555 ( 
.A(n_439),
.Y(n_555)
);

CKINVDCx5p33_ASAP7_75t_R g556 ( 
.A(n_441),
.Y(n_556)
);

CKINVDCx5p33_ASAP7_75t_R g557 ( 
.A(n_445),
.Y(n_557)
);

BUFx6f_ASAP7_75t_L g558 ( 
.A(n_436),
.Y(n_558)
);

CKINVDCx20_ASAP7_75t_R g559 ( 
.A(n_435),
.Y(n_559)
);

INVx2_ASAP7_75t_L g560 ( 
.A(n_442),
.Y(n_560)
);

CKINVDCx5p33_ASAP7_75t_R g561 ( 
.A(n_446),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_442),
.Y(n_562)
);

INVx3_ASAP7_75t_L g563 ( 
.A(n_443),
.Y(n_563)
);

CKINVDCx5p33_ASAP7_75t_R g564 ( 
.A(n_450),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_L g565 ( 
.A(n_459),
.B(n_264),
.Y(n_565)
);

AOI22xp33_ASAP7_75t_L g566 ( 
.A1(n_429),
.A2(n_350),
.B1(n_392),
.B2(n_386),
.Y(n_566)
);

INVxp67_ASAP7_75t_L g567 ( 
.A(n_453),
.Y(n_567)
);

CKINVDCx5p33_ASAP7_75t_R g568 ( 
.A(n_465),
.Y(n_568)
);

INVx1_ASAP7_75t_SL g569 ( 
.A(n_456),
.Y(n_569)
);

CKINVDCx5p33_ASAP7_75t_R g570 ( 
.A(n_467),
.Y(n_570)
);

BUFx6f_ASAP7_75t_L g571 ( 
.A(n_443),
.Y(n_571)
);

CKINVDCx5p33_ASAP7_75t_R g572 ( 
.A(n_469),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_444),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_444),
.Y(n_574)
);

BUFx6f_ASAP7_75t_L g575 ( 
.A(n_447),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_447),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_449),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_449),
.Y(n_578)
);

CKINVDCx5p33_ASAP7_75t_R g579 ( 
.A(n_474),
.Y(n_579)
);

INVx2_ASAP7_75t_L g580 ( 
.A(n_451),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_451),
.Y(n_581)
);

INVxp33_ASAP7_75t_L g582 ( 
.A(n_518),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_SL g583 ( 
.A(n_536),
.B(n_264),
.Y(n_583)
);

INVx3_ASAP7_75t_L g584 ( 
.A(n_508),
.Y(n_584)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_508),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_525),
.Y(n_586)
);

OAI22xp33_ASAP7_75t_L g587 ( 
.A1(n_520),
.A2(n_482),
.B1(n_411),
.B2(n_466),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_SL g588 ( 
.A(n_536),
.B(n_305),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_L g589 ( 
.A(n_500),
.B(n_476),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_L g590 ( 
.A(n_565),
.B(n_477),
.Y(n_590)
);

AND2x6_ASAP7_75t_L g591 ( 
.A(n_524),
.B(n_305),
.Y(n_591)
);

BUFx3_ASAP7_75t_L g592 ( 
.A(n_514),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_L g593 ( 
.A(n_553),
.B(n_522),
.Y(n_593)
);

AO22x2_ASAP7_75t_L g594 ( 
.A1(n_567),
.A2(n_401),
.B1(n_405),
.B2(n_398),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_508),
.Y(n_595)
);

BUFx8_ASAP7_75t_SL g596 ( 
.A(n_503),
.Y(n_596)
);

AOI22xp33_ASAP7_75t_L g597 ( 
.A1(n_553),
.A2(n_486),
.B1(n_490),
.B2(n_423),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_529),
.Y(n_598)
);

OR2x2_ASAP7_75t_L g599 ( 
.A(n_515),
.B(n_479),
.Y(n_599)
);

INVx2_ASAP7_75t_L g600 ( 
.A(n_508),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_L g601 ( 
.A(n_553),
.B(n_483),
.Y(n_601)
);

AND2x2_ASAP7_75t_L g602 ( 
.A(n_546),
.B(n_454),
.Y(n_602)
);

NOR2xp33_ASAP7_75t_L g603 ( 
.A(n_510),
.B(n_488),
.Y(n_603)
);

AOI22xp33_ASAP7_75t_L g604 ( 
.A1(n_553),
.A2(n_375),
.B1(n_386),
.B2(n_374),
.Y(n_604)
);

INVx3_ASAP7_75t_L g605 ( 
.A(n_558),
.Y(n_605)
);

NOR2xp33_ASAP7_75t_L g606 ( 
.A(n_516),
.B(n_457),
.Y(n_606)
);

NAND3xp33_ASAP7_75t_L g607 ( 
.A(n_566),
.B(n_521),
.C(n_509),
.Y(n_607)
);

AOI22xp5_ASAP7_75t_L g608 ( 
.A1(n_507),
.A2(n_478),
.B1(n_471),
.B2(n_440),
.Y(n_608)
);

BUFx3_ASAP7_75t_L g609 ( 
.A(n_524),
.Y(n_609)
);

INVx2_ASAP7_75t_L g610 ( 
.A(n_523),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_533),
.Y(n_611)
);

BUFx2_ASAP7_75t_L g612 ( 
.A(n_501),
.Y(n_612)
);

OAI22xp33_ASAP7_75t_L g613 ( 
.A1(n_516),
.A2(n_341),
.B1(n_308),
.B2(n_292),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_534),
.Y(n_614)
);

NOR2xp33_ASAP7_75t_L g615 ( 
.A(n_526),
.B(n_404),
.Y(n_615)
);

AND2x2_ASAP7_75t_L g616 ( 
.A(n_546),
.B(n_454),
.Y(n_616)
);

AOI22xp33_ASAP7_75t_L g617 ( 
.A1(n_553),
.A2(n_375),
.B1(n_392),
.B2(n_452),
.Y(n_617)
);

AOI22xp33_ASAP7_75t_L g618 ( 
.A1(n_553),
.A2(n_258),
.B1(n_291),
.B2(n_301),
.Y(n_618)
);

INVxp67_ASAP7_75t_L g619 ( 
.A(n_530),
.Y(n_619)
);

AND2x4_ASAP7_75t_L g620 ( 
.A(n_524),
.B(n_219),
.Y(n_620)
);

INVx3_ASAP7_75t_L g621 ( 
.A(n_558),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_L g622 ( 
.A(n_553),
.B(n_259),
.Y(n_622)
);

NOR2xp33_ASAP7_75t_L g623 ( 
.A(n_526),
.B(n_448),
.Y(n_623)
);

INVxp67_ASAP7_75t_SL g624 ( 
.A(n_558),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_543),
.B(n_290),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_535),
.Y(n_626)
);

OR2x2_ASAP7_75t_L g627 ( 
.A(n_569),
.B(n_431),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_SL g628 ( 
.A(n_542),
.B(n_314),
.Y(n_628)
);

BUFx3_ASAP7_75t_L g629 ( 
.A(n_542),
.Y(n_629)
);

INVx4_ASAP7_75t_L g630 ( 
.A(n_558),
.Y(n_630)
);

OR2x6_ASAP7_75t_L g631 ( 
.A(n_542),
.B(n_278),
.Y(n_631)
);

INVx2_ASAP7_75t_L g632 ( 
.A(n_523),
.Y(n_632)
);

OAI22xp5_ASAP7_75t_L g633 ( 
.A1(n_527),
.A2(n_323),
.B1(n_218),
.B2(n_225),
.Y(n_633)
);

INVx2_ASAP7_75t_L g634 ( 
.A(n_523),
.Y(n_634)
);

INVx2_ASAP7_75t_L g635 ( 
.A(n_523),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_SL g636 ( 
.A(n_527),
.B(n_314),
.Y(n_636)
);

BUFx6f_ASAP7_75t_SL g637 ( 
.A(n_531),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_544),
.Y(n_638)
);

INVx6_ASAP7_75t_L g639 ( 
.A(n_531),
.Y(n_639)
);

OR2x6_ASAP7_75t_L g640 ( 
.A(n_537),
.B(n_278),
.Y(n_640)
);

OR2x2_ASAP7_75t_L g641 ( 
.A(n_546),
.B(n_437),
.Y(n_641)
);

BUFx10_ASAP7_75t_L g642 ( 
.A(n_532),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_L g643 ( 
.A(n_543),
.B(n_295),
.Y(n_643)
);

OAI22xp33_ASAP7_75t_L g644 ( 
.A1(n_532),
.A2(n_279),
.B1(n_271),
.B2(n_265),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_547),
.Y(n_645)
);

AOI22xp33_ASAP7_75t_L g646 ( 
.A1(n_543),
.A2(n_563),
.B1(n_571),
.B2(n_558),
.Y(n_646)
);

AND2x2_ASAP7_75t_SL g647 ( 
.A(n_519),
.B(n_354),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_549),
.Y(n_648)
);

AND2x4_ASAP7_75t_L g649 ( 
.A(n_550),
.B(n_220),
.Y(n_649)
);

INVx4_ASAP7_75t_L g650 ( 
.A(n_571),
.Y(n_650)
);

CKINVDCx20_ASAP7_75t_R g651 ( 
.A(n_504),
.Y(n_651)
);

NOR2xp33_ASAP7_75t_L g652 ( 
.A(n_538),
.B(n_470),
.Y(n_652)
);

BUFx3_ASAP7_75t_L g653 ( 
.A(n_571),
.Y(n_653)
);

OR2x2_ASAP7_75t_L g654 ( 
.A(n_563),
.B(n_475),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_543),
.B(n_304),
.Y(n_655)
);

NAND2xp33_ASAP7_75t_L g656 ( 
.A(n_543),
.B(n_248),
.Y(n_656)
);

INVxp67_ASAP7_75t_SL g657 ( 
.A(n_571),
.Y(n_657)
);

NOR2xp33_ASAP7_75t_L g658 ( 
.A(n_538),
.B(n_498),
.Y(n_658)
);

BUFx2_ASAP7_75t_L g659 ( 
.A(n_501),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_554),
.Y(n_660)
);

INVx5_ASAP7_75t_L g661 ( 
.A(n_543),
.Y(n_661)
);

INVx2_ASAP7_75t_SL g662 ( 
.A(n_531),
.Y(n_662)
);

INVx8_ASAP7_75t_L g663 ( 
.A(n_543),
.Y(n_663)
);

INVx2_ASAP7_75t_L g664 ( 
.A(n_545),
.Y(n_664)
);

INVx2_ASAP7_75t_L g665 ( 
.A(n_545),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_573),
.Y(n_666)
);

INVx3_ASAP7_75t_L g667 ( 
.A(n_575),
.Y(n_667)
);

NOR2xp33_ASAP7_75t_SL g668 ( 
.A(n_540),
.B(n_548),
.Y(n_668)
);

AND2x2_ASAP7_75t_SL g669 ( 
.A(n_519),
.B(n_354),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_576),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_577),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_563),
.B(n_307),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_578),
.Y(n_673)
);

AND2x2_ASAP7_75t_L g674 ( 
.A(n_552),
.B(n_455),
.Y(n_674)
);

NOR2xp33_ASAP7_75t_L g675 ( 
.A(n_540),
.B(n_214),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_SL g676 ( 
.A(n_548),
.B(n_248),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_502),
.B(n_315),
.Y(n_677)
);

INVx3_ASAP7_75t_L g678 ( 
.A(n_575),
.Y(n_678)
);

INVx4_ASAP7_75t_L g679 ( 
.A(n_575),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_502),
.B(n_318),
.Y(n_680)
);

CKINVDCx5p33_ASAP7_75t_R g681 ( 
.A(n_528),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_SL g682 ( 
.A(n_551),
.B(n_299),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_581),
.Y(n_683)
);

INVx2_ASAP7_75t_L g684 ( 
.A(n_545),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_575),
.Y(n_685)
);

INVx4_ASAP7_75t_SL g686 ( 
.A(n_575),
.Y(n_686)
);

NOR2xp33_ASAP7_75t_L g687 ( 
.A(n_551),
.B(n_234),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_L g688 ( 
.A(n_506),
.B(n_321),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_L g689 ( 
.A(n_506),
.B(n_326),
.Y(n_689)
);

INVx4_ASAP7_75t_SL g690 ( 
.A(n_505),
.Y(n_690)
);

INVx3_ASAP7_75t_L g691 ( 
.A(n_539),
.Y(n_691)
);

BUFx6f_ASAP7_75t_L g692 ( 
.A(n_560),
.Y(n_692)
);

INVx4_ASAP7_75t_L g693 ( 
.A(n_539),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_L g694 ( 
.A(n_511),
.B(n_331),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_SL g695 ( 
.A(n_555),
.B(n_299),
.Y(n_695)
);

INVx2_ASAP7_75t_L g696 ( 
.A(n_539),
.Y(n_696)
);

INVx2_ASAP7_75t_L g697 ( 
.A(n_513),
.Y(n_697)
);

BUFx4f_ASAP7_75t_L g698 ( 
.A(n_512),
.Y(n_698)
);

AND2x2_ASAP7_75t_L g699 ( 
.A(n_560),
.B(n_455),
.Y(n_699)
);

INVx2_ASAP7_75t_L g700 ( 
.A(n_513),
.Y(n_700)
);

INVx4_ASAP7_75t_SL g701 ( 
.A(n_537),
.Y(n_701)
);

AOI22xp33_ASAP7_75t_L g702 ( 
.A1(n_562),
.A2(n_580),
.B1(n_574),
.B2(n_309),
.Y(n_702)
);

INVx2_ASAP7_75t_L g703 ( 
.A(n_580),
.Y(n_703)
);

INVx2_ASAP7_75t_L g704 ( 
.A(n_562),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_574),
.Y(n_705)
);

BUFx8_ASAP7_75t_SL g706 ( 
.A(n_541),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_555),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_556),
.Y(n_708)
);

INVx2_ASAP7_75t_L g709 ( 
.A(n_556),
.Y(n_709)
);

INVxp33_ASAP7_75t_SL g710 ( 
.A(n_557),
.Y(n_710)
);

INVxp67_ASAP7_75t_SL g711 ( 
.A(n_559),
.Y(n_711)
);

BUFx10_ASAP7_75t_L g712 ( 
.A(n_561),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_561),
.Y(n_713)
);

NOR2xp33_ASAP7_75t_L g714 ( 
.A(n_564),
.B(n_237),
.Y(n_714)
);

INVx4_ASAP7_75t_L g715 ( 
.A(n_568),
.Y(n_715)
);

OAI22xp33_ASAP7_75t_L g716 ( 
.A1(n_568),
.A2(n_336),
.B1(n_332),
.B2(n_330),
.Y(n_716)
);

INVx2_ASAP7_75t_L g717 ( 
.A(n_570),
.Y(n_717)
);

AOI22xp33_ASAP7_75t_L g718 ( 
.A1(n_570),
.A2(n_297),
.B1(n_395),
.B2(n_394),
.Y(n_718)
);

INVx2_ASAP7_75t_L g719 ( 
.A(n_572),
.Y(n_719)
);

OR2x6_ASAP7_75t_L g720 ( 
.A(n_517),
.B(n_220),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_572),
.Y(n_721)
);

AND2x2_ASAP7_75t_L g722 ( 
.A(n_579),
.B(n_458),
.Y(n_722)
);

INVx2_ASAP7_75t_L g723 ( 
.A(n_579),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_L g724 ( 
.A(n_517),
.B(n_335),
.Y(n_724)
);

INVx2_ASAP7_75t_L g725 ( 
.A(n_508),
.Y(n_725)
);

INVx3_ASAP7_75t_L g726 ( 
.A(n_508),
.Y(n_726)
);

INVx3_ASAP7_75t_L g727 ( 
.A(n_609),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_609),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_629),
.Y(n_729)
);

NOR2xp67_ASAP7_75t_L g730 ( 
.A(n_662),
.B(n_340),
.Y(n_730)
);

BUFx3_ASAP7_75t_L g731 ( 
.A(n_629),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_647),
.B(n_221),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_SL g733 ( 
.A(n_647),
.B(n_299),
.Y(n_733)
);

INVxp67_ASAP7_75t_L g734 ( 
.A(n_652),
.Y(n_734)
);

INVx3_ASAP7_75t_L g735 ( 
.A(n_691),
.Y(n_735)
);

AOI22xp5_ASAP7_75t_L g736 ( 
.A1(n_669),
.A2(n_343),
.B1(n_376),
.B2(n_379),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_674),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_L g738 ( 
.A(n_669),
.B(n_221),
.Y(n_738)
);

INVx2_ASAP7_75t_L g739 ( 
.A(n_703),
.Y(n_739)
);

AOI21xp5_ASAP7_75t_L g740 ( 
.A1(n_624),
.A2(n_262),
.B(n_261),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_L g741 ( 
.A(n_691),
.B(n_226),
.Y(n_741)
);

INVx2_ASAP7_75t_L g742 ( 
.A(n_703),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_L g743 ( 
.A(n_691),
.B(n_226),
.Y(n_743)
);

OAI22xp5_ASAP7_75t_L g744 ( 
.A1(n_582),
.A2(n_297),
.B1(n_281),
.B2(n_395),
.Y(n_744)
);

INVx2_ASAP7_75t_L g745 ( 
.A(n_704),
.Y(n_745)
);

AOI22xp33_ASAP7_75t_L g746 ( 
.A1(n_583),
.A2(n_334),
.B1(n_239),
.B2(n_394),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_589),
.B(n_233),
.Y(n_747)
);

INVx2_ASAP7_75t_L g748 ( 
.A(n_697),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_590),
.B(n_233),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_674),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_699),
.Y(n_751)
);

AND2x2_ASAP7_75t_L g752 ( 
.A(n_722),
.B(n_458),
.Y(n_752)
);

NOR2xp33_ASAP7_75t_L g753 ( 
.A(n_722),
.B(n_241),
.Y(n_753)
);

AOI22xp33_ASAP7_75t_L g754 ( 
.A1(n_583),
.A2(n_337),
.B1(n_245),
.B2(n_246),
.Y(n_754)
);

NOR2xp33_ASAP7_75t_L g755 ( 
.A(n_658),
.B(n_256),
.Y(n_755)
);

INVxp67_ASAP7_75t_L g756 ( 
.A(n_627),
.Y(n_756)
);

INVx2_ASAP7_75t_SL g757 ( 
.A(n_627),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_699),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_586),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_693),
.B(n_244),
.Y(n_760)
);

O2A1O1Ixp5_ASAP7_75t_L g761 ( 
.A1(n_588),
.A2(n_334),
.B(n_389),
.C(n_388),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_598),
.Y(n_762)
);

INVx2_ASAP7_75t_L g763 ( 
.A(n_697),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_L g764 ( 
.A(n_693),
.B(n_244),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_SL g765 ( 
.A(n_661),
.B(n_299),
.Y(n_765)
);

NOR3xp33_ASAP7_75t_L g766 ( 
.A(n_613),
.B(n_257),
.C(n_396),
.Y(n_766)
);

AND2x2_ASAP7_75t_L g767 ( 
.A(n_662),
.B(n_461),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_SL g768 ( 
.A(n_661),
.B(n_693),
.Y(n_768)
);

NOR2xp67_ASAP7_75t_L g769 ( 
.A(n_715),
.B(n_344),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_L g770 ( 
.A(n_588),
.B(n_245),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_611),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_614),
.Y(n_772)
);

BUFx6f_ASAP7_75t_L g773 ( 
.A(n_591),
.Y(n_773)
);

CKINVDCx5p33_ASAP7_75t_R g774 ( 
.A(n_596),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_SL g775 ( 
.A(n_661),
.B(n_299),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_602),
.B(n_616),
.Y(n_776)
);

INVx3_ASAP7_75t_L g777 ( 
.A(n_692),
.Y(n_777)
);

AND2x2_ASAP7_75t_L g778 ( 
.A(n_639),
.B(n_675),
.Y(n_778)
);

AOI22xp33_ASAP7_75t_L g779 ( 
.A1(n_591),
.A2(n_378),
.B1(n_246),
.B2(n_266),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_602),
.B(n_266),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_616),
.B(n_281),
.Y(n_781)
);

NOR2xp33_ASAP7_75t_L g782 ( 
.A(n_636),
.B(n_260),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_626),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_638),
.Y(n_784)
);

OAI22xp33_ASAP7_75t_L g785 ( 
.A1(n_607),
.A2(n_283),
.B1(n_313),
.B2(n_319),
.Y(n_785)
);

INVx2_ASAP7_75t_SL g786 ( 
.A(n_592),
.Y(n_786)
);

AOI22xp5_ASAP7_75t_L g787 ( 
.A1(n_603),
.A2(n_356),
.B1(n_346),
.B2(n_352),
.Y(n_787)
);

AO22x1_ASAP7_75t_L g788 ( 
.A1(n_687),
.A2(n_714),
.B1(n_619),
.B2(n_620),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_645),
.Y(n_789)
);

OAI22xp33_ASAP7_75t_L g790 ( 
.A1(n_720),
.A2(n_283),
.B1(n_313),
.B2(n_319),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_648),
.Y(n_791)
);

INVx2_ASAP7_75t_L g792 ( 
.A(n_700),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_L g793 ( 
.A(n_660),
.B(n_324),
.Y(n_793)
);

AOI22xp5_ASAP7_75t_L g794 ( 
.A1(n_631),
.A2(n_370),
.B1(n_372),
.B2(n_373),
.Y(n_794)
);

NOR2xp33_ASAP7_75t_L g795 ( 
.A(n_636),
.B(n_285),
.Y(n_795)
);

AOI22xp33_ASAP7_75t_L g796 ( 
.A1(n_591),
.A2(n_381),
.B1(n_324),
.B2(n_337),
.Y(n_796)
);

CKINVDCx5p33_ASAP7_75t_R g797 ( 
.A(n_596),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_SL g798 ( 
.A(n_661),
.B(n_298),
.Y(n_798)
);

NOR2xp33_ASAP7_75t_L g799 ( 
.A(n_587),
.B(n_302),
.Y(n_799)
);

OR2x2_ASAP7_75t_L g800 ( 
.A(n_633),
.B(n_461),
.Y(n_800)
);

BUFx6f_ASAP7_75t_SL g801 ( 
.A(n_642),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_SL g802 ( 
.A(n_661),
.B(n_303),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_666),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_L g804 ( 
.A(n_670),
.B(n_342),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_SL g805 ( 
.A(n_593),
.B(n_384),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_L g806 ( 
.A(n_671),
.B(n_342),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_673),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_683),
.Y(n_808)
);

HB1xp67_ASAP7_75t_L g809 ( 
.A(n_599),
.Y(n_809)
);

NOR3xp33_ASAP7_75t_L g810 ( 
.A(n_644),
.B(n_329),
.C(n_320),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_L g811 ( 
.A(n_672),
.B(n_348),
.Y(n_811)
);

INVxp67_ASAP7_75t_L g812 ( 
.A(n_623),
.Y(n_812)
);

INVx4_ASAP7_75t_L g813 ( 
.A(n_692),
.Y(n_813)
);

AND2x2_ASAP7_75t_L g814 ( 
.A(n_639),
.B(n_462),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_SL g815 ( 
.A(n_622),
.B(n_348),
.Y(n_815)
);

INVx2_ASAP7_75t_SL g816 ( 
.A(n_592),
.Y(n_816)
);

INVx2_ASAP7_75t_L g817 ( 
.A(n_700),
.Y(n_817)
);

INVx4_ASAP7_75t_L g818 ( 
.A(n_663),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_L g819 ( 
.A(n_692),
.B(n_362),
.Y(n_819)
);

NOR3xp33_ASAP7_75t_L g820 ( 
.A(n_716),
.B(n_365),
.C(n_310),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_L g821 ( 
.A(n_641),
.B(n_362),
.Y(n_821)
);

BUFx6f_ASAP7_75t_SL g822 ( 
.A(n_642),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_L g823 ( 
.A(n_641),
.B(n_364),
.Y(n_823)
);

INVx2_ASAP7_75t_L g824 ( 
.A(n_696),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_L g825 ( 
.A(n_654),
.B(n_364),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_L g826 ( 
.A(n_654),
.B(n_378),
.Y(n_826)
);

INVx4_ASAP7_75t_L g827 ( 
.A(n_663),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_L g828 ( 
.A(n_677),
.B(n_680),
.Y(n_828)
);

NOR2xp33_ASAP7_75t_L g829 ( 
.A(n_676),
.B(n_311),
.Y(n_829)
);

INVx2_ASAP7_75t_L g830 ( 
.A(n_705),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_SL g831 ( 
.A(n_646),
.B(n_381),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_SL g832 ( 
.A(n_601),
.B(n_385),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_649),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_688),
.B(n_385),
.Y(n_834)
);

A2O1A1Ixp33_ASAP7_75t_L g835 ( 
.A1(n_718),
.A2(n_388),
.B(n_389),
.C(n_493),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_L g836 ( 
.A(n_689),
.B(n_462),
.Y(n_836)
);

NAND2xp33_ASAP7_75t_L g837 ( 
.A(n_617),
.B(n_312),
.Y(n_837)
);

AOI22xp5_ASAP7_75t_L g838 ( 
.A1(n_631),
.A2(n_296),
.B1(n_322),
.B2(n_345),
.Y(n_838)
);

AND2x4_ASAP7_75t_L g839 ( 
.A(n_620),
.B(n_463),
.Y(n_839)
);

INVx4_ASAP7_75t_L g840 ( 
.A(n_663),
.Y(n_840)
);

NOR3x1_ASAP7_75t_L g841 ( 
.A(n_612),
.B(n_227),
.C(n_495),
.Y(n_841)
);

INVx4_ASAP7_75t_L g842 ( 
.A(n_663),
.Y(n_842)
);

NOR2xp33_ASAP7_75t_L g843 ( 
.A(n_676),
.B(n_353),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_L g844 ( 
.A(n_657),
.B(n_463),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_SL g845 ( 
.A(n_698),
.B(n_597),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_L g846 ( 
.A(n_620),
.B(n_464),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_L g847 ( 
.A(n_694),
.B(n_464),
.Y(n_847)
);

NOR2xp67_ASAP7_75t_L g848 ( 
.A(n_715),
.B(n_615),
.Y(n_848)
);

OAI22xp33_ASAP7_75t_L g849 ( 
.A1(n_720),
.A2(n_360),
.B1(n_357),
.B2(n_355),
.Y(n_849)
);

HB1xp67_ASAP7_75t_L g850 ( 
.A(n_681),
.Y(n_850)
);

OAI22xp33_ASAP7_75t_L g851 ( 
.A1(n_720),
.A2(n_393),
.B1(n_358),
.B2(n_361),
.Y(n_851)
);

INVx2_ASAP7_75t_L g852 ( 
.A(n_585),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_649),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_605),
.B(n_621),
.Y(n_854)
);

INVx2_ASAP7_75t_L g855 ( 
.A(n_595),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_SL g856 ( 
.A(n_698),
.B(n_595),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_605),
.B(n_468),
.Y(n_857)
);

INVx2_ASAP7_75t_L g858 ( 
.A(n_600),
.Y(n_858)
);

NAND3xp33_ASAP7_75t_SL g859 ( 
.A(n_608),
.B(n_371),
.C(n_380),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_L g860 ( 
.A(n_605),
.B(n_621),
.Y(n_860)
);

INVx2_ASAP7_75t_L g861 ( 
.A(n_600),
.Y(n_861)
);

OAI221xp5_ASAP7_75t_L g862 ( 
.A1(n_702),
.A2(n_497),
.B1(n_495),
.B2(n_493),
.C(n_491),
.Y(n_862)
);

OAI22xp5_ASAP7_75t_L g863 ( 
.A1(n_631),
.A2(n_390),
.B1(n_391),
.B2(n_489),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_621),
.B(n_497),
.Y(n_864)
);

NOR2xp33_ASAP7_75t_L g865 ( 
.A(n_682),
.B(n_695),
.Y(n_865)
);

OR2x2_ASAP7_75t_L g866 ( 
.A(n_720),
.B(n_491),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_667),
.B(n_489),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_667),
.B(n_484),
.Y(n_868)
);

INVx1_ASAP7_75t_SL g869 ( 
.A(n_659),
.Y(n_869)
);

AND2x4_ASAP7_75t_L g870 ( 
.A(n_649),
.B(n_484),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_L g871 ( 
.A(n_667),
.B(n_678),
.Y(n_871)
);

INVx2_ASAP7_75t_L g872 ( 
.A(n_725),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_SL g873 ( 
.A(n_698),
.B(n_369),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_L g874 ( 
.A(n_678),
.B(n_480),
.Y(n_874)
);

NOR2xp33_ASAP7_75t_SL g875 ( 
.A(n_637),
.B(n_369),
.Y(n_875)
);

BUFx3_ASAP7_75t_L g876 ( 
.A(n_639),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_SL g877 ( 
.A(n_725),
.B(n_369),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_SL g878 ( 
.A(n_610),
.B(n_632),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_678),
.B(n_480),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_628),
.Y(n_880)
);

NOR3xp33_ASAP7_75t_L g881 ( 
.A(n_606),
.B(n_473),
.C(n_472),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_SL g882 ( 
.A(n_610),
.B(n_201),
.Y(n_882)
);

CKINVDCx5p33_ASAP7_75t_R g883 ( 
.A(n_706),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_L g884 ( 
.A(n_653),
.B(n_473),
.Y(n_884)
);

NOR2xp67_ASAP7_75t_L g885 ( 
.A(n_715),
.B(n_156),
.Y(n_885)
);

OR2x2_ASAP7_75t_L g886 ( 
.A(n_682),
.B(n_468),
.Y(n_886)
);

AOI22xp33_ASAP7_75t_L g887 ( 
.A1(n_591),
.A2(n_604),
.B1(n_618),
.B2(n_640),
.Y(n_887)
);

AOI21xp5_ASAP7_75t_L g888 ( 
.A1(n_625),
.A2(n_201),
.B(n_377),
.Y(n_888)
);

INVx8_ASAP7_75t_L g889 ( 
.A(n_631),
.Y(n_889)
);

AO21x1_ASAP7_75t_L g890 ( 
.A1(n_733),
.A2(n_695),
.B(n_643),
.Y(n_890)
);

INVx4_ASAP7_75t_L g891 ( 
.A(n_876),
.Y(n_891)
);

AND2x4_ASAP7_75t_L g892 ( 
.A(n_731),
.B(n_709),
.Y(n_892)
);

AO21x2_ASAP7_75t_L g893 ( 
.A1(n_832),
.A2(n_845),
.B(n_738),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_SL g894 ( 
.A(n_848),
.B(n_709),
.Y(n_894)
);

OAI22xp5_ASAP7_75t_L g895 ( 
.A1(n_887),
.A2(n_719),
.B1(n_723),
.B2(n_717),
.Y(n_895)
);

AOI21xp5_ASAP7_75t_L g896 ( 
.A1(n_818),
.A2(n_679),
.B(n_630),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_L g897 ( 
.A(n_865),
.B(n_717),
.Y(n_897)
);

AOI21xp5_ASAP7_75t_L g898 ( 
.A1(n_818),
.A2(n_679),
.B(n_630),
.Y(n_898)
);

O2A1O1Ixp33_ASAP7_75t_L g899 ( 
.A1(n_744),
.A2(n_656),
.B(n_719),
.C(n_655),
.Y(n_899)
);

BUFx12f_ASAP7_75t_L g900 ( 
.A(n_757),
.Y(n_900)
);

NOR2xp33_ASAP7_75t_SL g901 ( 
.A(n_869),
.B(n_710),
.Y(n_901)
);

INVx5_ASAP7_75t_L g902 ( 
.A(n_773),
.Y(n_902)
);

BUFx3_ASAP7_75t_L g903 ( 
.A(n_876),
.Y(n_903)
);

AOI21xp5_ASAP7_75t_L g904 ( 
.A1(n_818),
.A2(n_679),
.B(n_650),
.Y(n_904)
);

AND2x2_ASAP7_75t_L g905 ( 
.A(n_752),
.B(n_756),
.Y(n_905)
);

BUFx3_ASAP7_75t_L g906 ( 
.A(n_774),
.Y(n_906)
);

OAI21xp5_ASAP7_75t_L g907 ( 
.A1(n_776),
.A2(n_640),
.B(n_591),
.Y(n_907)
);

AOI21xp5_ASAP7_75t_L g908 ( 
.A1(n_827),
.A2(n_842),
.B(n_840),
.Y(n_908)
);

INVx3_ASAP7_75t_L g909 ( 
.A(n_727),
.Y(n_909)
);

NAND3xp33_ASAP7_75t_L g910 ( 
.A(n_755),
.B(n_668),
.C(n_707),
.Y(n_910)
);

O2A1O1Ixp33_ASAP7_75t_SL g911 ( 
.A1(n_733),
.A2(n_724),
.B(n_685),
.C(n_635),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_865),
.B(n_591),
.Y(n_912)
);

O2A1O1Ixp33_ASAP7_75t_L g913 ( 
.A1(n_785),
.A2(n_708),
.B(n_721),
.C(n_713),
.Y(n_913)
);

OAI21xp5_ASAP7_75t_L g914 ( 
.A1(n_845),
.A2(n_640),
.B(n_634),
.Y(n_914)
);

AOI21xp5_ASAP7_75t_L g915 ( 
.A1(n_840),
.A2(n_842),
.B(n_768),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_SL g916 ( 
.A(n_734),
.B(n_778),
.Y(n_916)
);

OAI21x1_ASAP7_75t_L g917 ( 
.A1(n_878),
.A2(n_860),
.B(n_854),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_L g918 ( 
.A(n_755),
.B(n_584),
.Y(n_918)
);

BUFx2_ASAP7_75t_L g919 ( 
.A(n_850),
.Y(n_919)
);

BUFx2_ASAP7_75t_L g920 ( 
.A(n_814),
.Y(n_920)
);

AOI21xp5_ASAP7_75t_L g921 ( 
.A1(n_813),
.A2(n_684),
.B(n_664),
.Y(n_921)
);

INVx2_ASAP7_75t_L g922 ( 
.A(n_824),
.Y(n_922)
);

OAI22xp5_ASAP7_75t_L g923 ( 
.A1(n_746),
.A2(n_710),
.B1(n_594),
.B2(n_637),
.Y(n_923)
);

AOI21xp5_ASAP7_75t_L g924 ( 
.A1(n_813),
.A2(n_664),
.B(n_665),
.Y(n_924)
);

CKINVDCx20_ASAP7_75t_R g925 ( 
.A(n_797),
.Y(n_925)
);

OAI21xp33_ASAP7_75t_L g926 ( 
.A1(n_753),
.A2(n_594),
.B(n_711),
.Y(n_926)
);

AOI21xp5_ASAP7_75t_L g927 ( 
.A1(n_856),
.A2(n_871),
.B(n_878),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_824),
.Y(n_928)
);

OAI21xp5_ASAP7_75t_L g929 ( 
.A1(n_780),
.A2(n_684),
.B(n_584),
.Y(n_929)
);

AO21x1_ASAP7_75t_L g930 ( 
.A1(n_832),
.A2(n_701),
.B(n_594),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_SL g931 ( 
.A(n_767),
.B(n_712),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_SL g932 ( 
.A(n_786),
.B(n_712),
.Y(n_932)
);

BUFx2_ASAP7_75t_L g933 ( 
.A(n_809),
.Y(n_933)
);

AOI21xp5_ASAP7_75t_L g934 ( 
.A1(n_856),
.A2(n_726),
.B(n_584),
.Y(n_934)
);

INVxp67_ASAP7_75t_L g935 ( 
.A(n_753),
.Y(n_935)
);

AOI21xp5_ASAP7_75t_L g936 ( 
.A1(n_805),
.A2(n_726),
.B(n_686),
.Y(n_936)
);

NOR3xp33_ASAP7_75t_L g937 ( 
.A(n_788),
.B(n_681),
.C(n_637),
.Y(n_937)
);

NOR2xp67_ASAP7_75t_L g938 ( 
.A(n_812),
.B(n_726),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_SL g939 ( 
.A(n_816),
.B(n_712),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_L g940 ( 
.A(n_747),
.B(n_701),
.Y(n_940)
);

AND2x4_ASAP7_75t_L g941 ( 
.A(n_731),
.B(n_690),
.Y(n_941)
);

AOI21xp5_ASAP7_75t_L g942 ( 
.A1(n_805),
.A2(n_686),
.B(n_701),
.Y(n_942)
);

AO32x1_ASAP7_75t_L g943 ( 
.A1(n_863),
.A2(n_701),
.A3(n_690),
.B1(n_14),
.B2(n_16),
.Y(n_943)
);

NOR3xp33_ASAP7_75t_L g944 ( 
.A(n_859),
.B(n_642),
.C(n_706),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_L g945 ( 
.A(n_749),
.B(n_686),
.Y(n_945)
);

NOR2xp33_ASAP7_75t_L g946 ( 
.A(n_799),
.B(n_651),
.Y(n_946)
);

A2O1A1Ixp33_ASAP7_75t_L g947 ( 
.A1(n_782),
.A2(n_651),
.B(n_690),
.C(n_17),
.Y(n_947)
);

AOI21xp5_ASAP7_75t_L g948 ( 
.A1(n_844),
.A2(n_764),
.B(n_760),
.Y(n_948)
);

NOR2xp33_ASAP7_75t_L g949 ( 
.A(n_799),
.B(n_11),
.Y(n_949)
);

NOR2xp33_ASAP7_75t_L g950 ( 
.A(n_849),
.B(n_12),
.Y(n_950)
);

AOI21xp5_ASAP7_75t_L g951 ( 
.A1(n_836),
.A2(n_686),
.B(n_690),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_L g952 ( 
.A(n_847),
.B(n_12),
.Y(n_952)
);

NOR2xp33_ASAP7_75t_L g953 ( 
.A(n_838),
.B(n_18),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_L g954 ( 
.A(n_737),
.B(n_18),
.Y(n_954)
);

NAND3xp33_ASAP7_75t_L g955 ( 
.A(n_782),
.B(n_20),
.C(n_22),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_L g956 ( 
.A(n_750),
.B(n_24),
.Y(n_956)
);

AND2x6_ASAP7_75t_L g957 ( 
.A(n_773),
.B(n_191),
.Y(n_957)
);

AND2x2_ASAP7_75t_L g958 ( 
.A(n_751),
.B(n_25),
.Y(n_958)
);

INVx2_ASAP7_75t_L g959 ( 
.A(n_739),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_L g960 ( 
.A(n_758),
.B(n_26),
.Y(n_960)
);

OAI22xp5_ASAP7_75t_L g961 ( 
.A1(n_754),
.A2(n_26),
.B1(n_31),
.B2(n_32),
.Y(n_961)
);

INVx2_ASAP7_75t_L g962 ( 
.A(n_742),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_L g963 ( 
.A(n_833),
.B(n_853),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_L g964 ( 
.A(n_870),
.B(n_32),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_L g965 ( 
.A(n_870),
.B(n_821),
.Y(n_965)
);

AND2x2_ASAP7_75t_L g966 ( 
.A(n_881),
.B(n_33),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_L g967 ( 
.A(n_870),
.B(n_34),
.Y(n_967)
);

O2A1O1Ixp33_ASAP7_75t_L g968 ( 
.A1(n_837),
.A2(n_39),
.B(n_42),
.C(n_44),
.Y(n_968)
);

INVx2_ASAP7_75t_SL g969 ( 
.A(n_866),
.Y(n_969)
);

NOR2xp33_ASAP7_75t_L g970 ( 
.A(n_795),
.B(n_39),
.Y(n_970)
);

OAI21xp5_ASAP7_75t_L g971 ( 
.A1(n_781),
.A2(n_164),
.B(n_163),
.Y(n_971)
);

INVx2_ASAP7_75t_L g972 ( 
.A(n_742),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_L g973 ( 
.A(n_735),
.B(n_115),
.Y(n_973)
);

AOI21xp5_ASAP7_75t_L g974 ( 
.A1(n_735),
.A2(n_151),
.B(n_143),
.Y(n_974)
);

AOI22xp5_ASAP7_75t_L g975 ( 
.A1(n_795),
.A2(n_142),
.B1(n_126),
.B2(n_110),
.Y(n_975)
);

NOR2xp33_ASAP7_75t_L g976 ( 
.A(n_800),
.B(n_42),
.Y(n_976)
);

AOI21xp5_ASAP7_75t_L g977 ( 
.A1(n_777),
.A2(n_101),
.B(n_93),
.Y(n_977)
);

A2O1A1Ixp33_ASAP7_75t_L g978 ( 
.A1(n_829),
.A2(n_44),
.B(n_47),
.C(n_49),
.Y(n_978)
);

NAND2xp5_ASAP7_75t_L g979 ( 
.A(n_823),
.B(n_825),
.Y(n_979)
);

OAI22xp5_ASAP7_75t_L g980 ( 
.A1(n_826),
.A2(n_49),
.B1(n_50),
.B2(n_51),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_L g981 ( 
.A(n_811),
.B(n_76),
.Y(n_981)
);

AOI21xp5_ASAP7_75t_L g982 ( 
.A1(n_777),
.A2(n_53),
.B(n_54),
.Y(n_982)
);

BUFx6f_ASAP7_75t_L g983 ( 
.A(n_773),
.Y(n_983)
);

AND2x2_ASAP7_75t_L g984 ( 
.A(n_839),
.B(n_57),
.Y(n_984)
);

AOI21x1_ASAP7_75t_L g985 ( 
.A1(n_741),
.A2(n_58),
.B(n_59),
.Y(n_985)
);

AOI21xp5_ASAP7_75t_L g986 ( 
.A1(n_846),
.A2(n_58),
.B(n_59),
.Y(n_986)
);

HB1xp67_ASAP7_75t_L g987 ( 
.A(n_839),
.Y(n_987)
);

OAI21xp5_ASAP7_75t_L g988 ( 
.A1(n_770),
.A2(n_815),
.B(n_743),
.Y(n_988)
);

AO32x1_ASAP7_75t_L g989 ( 
.A1(n_852),
.A2(n_872),
.A3(n_861),
.B1(n_858),
.B2(n_855),
.Y(n_989)
);

OR2x6_ASAP7_75t_L g990 ( 
.A(n_889),
.B(n_65),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_L g991 ( 
.A(n_834),
.B(n_60),
.Y(n_991)
);

O2A1O1Ixp33_ASAP7_75t_L g992 ( 
.A1(n_835),
.A2(n_63),
.B(n_815),
.C(n_831),
.Y(n_992)
);

A2O1A1Ixp33_ASAP7_75t_L g993 ( 
.A1(n_829),
.A2(n_843),
.B(n_886),
.C(n_839),
.Y(n_993)
);

AOI22xp5_ASAP7_75t_L g994 ( 
.A1(n_843),
.A2(n_728),
.B1(n_729),
.B2(n_873),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_L g995 ( 
.A(n_759),
.B(n_762),
.Y(n_995)
);

CKINVDCx11_ASAP7_75t_R g996 ( 
.A(n_889),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_830),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_L g998 ( 
.A(n_771),
.B(n_807),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_L g999 ( 
.A(n_772),
.B(n_803),
.Y(n_999)
);

O2A1O1Ixp33_ASAP7_75t_SL g1000 ( 
.A1(n_835),
.A2(n_831),
.B(n_873),
.C(n_775),
.Y(n_1000)
);

INVx1_ASAP7_75t_SL g1001 ( 
.A(n_883),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_L g1002 ( 
.A(n_783),
.B(n_791),
.Y(n_1002)
);

O2A1O1Ixp5_ASAP7_75t_L g1003 ( 
.A1(n_888),
.A2(n_761),
.B(n_830),
.C(n_819),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_L g1004 ( 
.A(n_784),
.B(n_808),
.Y(n_1004)
);

INVx1_ASAP7_75t_SL g1005 ( 
.A(n_877),
.Y(n_1005)
);

NOR2xp33_ASAP7_75t_L g1006 ( 
.A(n_851),
.B(n_789),
.Y(n_1006)
);

OAI22xp5_ASAP7_75t_L g1007 ( 
.A1(n_779),
.A2(n_796),
.B1(n_790),
.B2(n_804),
.Y(n_1007)
);

AND2x2_ASAP7_75t_L g1008 ( 
.A(n_766),
.B(n_810),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_L g1009 ( 
.A(n_884),
.B(n_857),
.Y(n_1009)
);

BUFx8_ASAP7_75t_L g1010 ( 
.A(n_801),
.Y(n_1010)
);

CKINVDCx6p67_ASAP7_75t_R g1011 ( 
.A(n_801),
.Y(n_1011)
);

INVx2_ASAP7_75t_L g1012 ( 
.A(n_745),
.Y(n_1012)
);

AO22x1_ASAP7_75t_L g1013 ( 
.A1(n_820),
.A2(n_841),
.B1(n_793),
.B2(n_806),
.Y(n_1013)
);

AOI21xp5_ASAP7_75t_L g1014 ( 
.A1(n_745),
.A2(n_817),
.B(n_792),
.Y(n_1014)
);

AOI21xp5_ASAP7_75t_L g1015 ( 
.A1(n_748),
.A2(n_817),
.B(n_763),
.Y(n_1015)
);

INVx2_ASAP7_75t_L g1016 ( 
.A(n_864),
.Y(n_1016)
);

INVx2_ASAP7_75t_L g1017 ( 
.A(n_867),
.Y(n_1017)
);

CKINVDCx10_ASAP7_75t_R g1018 ( 
.A(n_822),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_SL g1019 ( 
.A(n_769),
.B(n_730),
.Y(n_1019)
);

INVx2_ASAP7_75t_L g1020 ( 
.A(n_868),
.Y(n_1020)
);

OAI21xp5_ASAP7_75t_L g1021 ( 
.A1(n_874),
.A2(n_879),
.B(n_740),
.Y(n_1021)
);

NAND2xp5_ASAP7_75t_L g1022 ( 
.A(n_885),
.B(n_787),
.Y(n_1022)
);

AO21x1_ASAP7_75t_L g1023 ( 
.A1(n_877),
.A2(n_882),
.B(n_802),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_L g1024 ( 
.A(n_736),
.B(n_882),
.Y(n_1024)
);

NAND2xp5_ASAP7_75t_SL g1025 ( 
.A(n_875),
.B(n_794),
.Y(n_1025)
);

INVx3_ASAP7_75t_L g1026 ( 
.A(n_773),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_862),
.Y(n_1027)
);

AND2x2_ASAP7_75t_L g1028 ( 
.A(n_889),
.B(n_798),
.Y(n_1028)
);

NOR2xp33_ASAP7_75t_L g1029 ( 
.A(n_822),
.B(n_765),
.Y(n_1029)
);

NOR3xp33_ASAP7_75t_L g1030 ( 
.A(n_788),
.B(n_755),
.C(n_859),
.Y(n_1030)
);

NAND2xp5_ASAP7_75t_L g1031 ( 
.A(n_865),
.B(n_647),
.Y(n_1031)
);

AOI21xp5_ASAP7_75t_L g1032 ( 
.A1(n_818),
.A2(n_840),
.B(n_827),
.Y(n_1032)
);

O2A1O1Ixp33_ASAP7_75t_L g1033 ( 
.A1(n_732),
.A2(n_738),
.B(n_744),
.C(n_785),
.Y(n_1033)
);

AOI21xp5_ASAP7_75t_L g1034 ( 
.A1(n_818),
.A2(n_840),
.B(n_827),
.Y(n_1034)
);

NAND2xp5_ASAP7_75t_L g1035 ( 
.A(n_865),
.B(n_647),
.Y(n_1035)
);

AOI22xp33_ASAP7_75t_L g1036 ( 
.A1(n_845),
.A2(n_669),
.B1(n_647),
.B2(n_799),
.Y(n_1036)
);

BUFx6f_ASAP7_75t_L g1037 ( 
.A(n_731),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_L g1038 ( 
.A(n_776),
.B(n_828),
.Y(n_1038)
);

A2O1A1Ixp33_ASAP7_75t_L g1039 ( 
.A1(n_865),
.A2(n_755),
.B(n_795),
.C(n_782),
.Y(n_1039)
);

INVx3_ASAP7_75t_L g1040 ( 
.A(n_727),
.Y(n_1040)
);

NAND2xp5_ASAP7_75t_L g1041 ( 
.A(n_776),
.B(n_828),
.Y(n_1041)
);

INVx6_ASAP7_75t_L g1042 ( 
.A(n_876),
.Y(n_1042)
);

OAI21xp5_ASAP7_75t_L g1043 ( 
.A1(n_776),
.A2(n_845),
.B(n_738),
.Y(n_1043)
);

OAI22xp5_ASAP7_75t_L g1044 ( 
.A1(n_887),
.A2(n_738),
.B1(n_732),
.B2(n_647),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_L g1045 ( 
.A(n_865),
.B(n_647),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_SL g1046 ( 
.A(n_848),
.B(n_662),
.Y(n_1046)
);

OAI22xp5_ASAP7_75t_L g1047 ( 
.A1(n_887),
.A2(n_738),
.B1(n_732),
.B2(n_647),
.Y(n_1047)
);

BUFx3_ASAP7_75t_L g1048 ( 
.A(n_876),
.Y(n_1048)
);

NAND2xp5_ASAP7_75t_L g1049 ( 
.A(n_865),
.B(n_647),
.Y(n_1049)
);

O2A1O1Ixp33_ASAP7_75t_L g1050 ( 
.A1(n_732),
.A2(n_738),
.B(n_744),
.C(n_785),
.Y(n_1050)
);

AOI22xp5_ASAP7_75t_L g1051 ( 
.A1(n_865),
.A2(n_845),
.B1(n_755),
.B2(n_880),
.Y(n_1051)
);

NAND2xp5_ASAP7_75t_SL g1052 ( 
.A(n_848),
.B(n_662),
.Y(n_1052)
);

AOI21xp5_ASAP7_75t_L g1053 ( 
.A1(n_1038),
.A2(n_1041),
.B(n_948),
.Y(n_1053)
);

NAND2xp5_ASAP7_75t_L g1054 ( 
.A(n_1038),
.B(n_1041),
.Y(n_1054)
);

AO21x2_ASAP7_75t_L g1055 ( 
.A1(n_914),
.A2(n_1039),
.B(n_929),
.Y(n_1055)
);

NAND2xp5_ASAP7_75t_L g1056 ( 
.A(n_935),
.B(n_979),
.Y(n_1056)
);

AOI21xp33_ASAP7_75t_L g1057 ( 
.A1(n_970),
.A2(n_949),
.B(n_1033),
.Y(n_1057)
);

AOI221x1_ASAP7_75t_L g1058 ( 
.A1(n_926),
.A2(n_1030),
.B1(n_1044),
.B2(n_1047),
.C(n_947),
.Y(n_1058)
);

AOI21xp5_ASAP7_75t_L g1059 ( 
.A1(n_912),
.A2(n_907),
.B(n_915),
.Y(n_1059)
);

OAI21x1_ASAP7_75t_L g1060 ( 
.A1(n_917),
.A2(n_927),
.B(n_934),
.Y(n_1060)
);

INVx1_ASAP7_75t_L g1061 ( 
.A(n_963),
.Y(n_1061)
);

INVx1_ASAP7_75t_L g1062 ( 
.A(n_928),
.Y(n_1062)
);

BUFx3_ASAP7_75t_L g1063 ( 
.A(n_900),
.Y(n_1063)
);

AOI21x1_ASAP7_75t_L g1064 ( 
.A1(n_940),
.A2(n_918),
.B(n_973),
.Y(n_1064)
);

AOI21xp5_ASAP7_75t_L g1065 ( 
.A1(n_907),
.A2(n_1009),
.B(n_965),
.Y(n_1065)
);

AOI21xp33_ASAP7_75t_L g1066 ( 
.A1(n_1050),
.A2(n_1047),
.B(n_1044),
.Y(n_1066)
);

OAI21x1_ASAP7_75t_L g1067 ( 
.A1(n_896),
.A2(n_904),
.B(n_898),
.Y(n_1067)
);

OR2x6_ASAP7_75t_L g1068 ( 
.A(n_990),
.B(n_919),
.Y(n_1068)
);

OAI21xp5_ASAP7_75t_SL g1069 ( 
.A1(n_953),
.A2(n_1036),
.B(n_950),
.Y(n_1069)
);

NAND2xp5_ASAP7_75t_L g1070 ( 
.A(n_979),
.B(n_1051),
.Y(n_1070)
);

NAND2xp5_ASAP7_75t_L g1071 ( 
.A(n_897),
.B(n_1031),
.Y(n_1071)
);

OAI21xp5_ASAP7_75t_L g1072 ( 
.A1(n_1043),
.A2(n_1045),
.B(n_1035),
.Y(n_1072)
);

OAI21x1_ASAP7_75t_SL g1073 ( 
.A1(n_930),
.A2(n_971),
.B(n_1023),
.Y(n_1073)
);

AOI21xp33_ASAP7_75t_L g1074 ( 
.A1(n_1049),
.A2(n_976),
.B(n_1024),
.Y(n_1074)
);

INVx2_ASAP7_75t_L g1075 ( 
.A(n_922),
.Y(n_1075)
);

AND2x2_ASAP7_75t_L g1076 ( 
.A(n_905),
.B(n_920),
.Y(n_1076)
);

NAND2xp5_ASAP7_75t_L g1077 ( 
.A(n_895),
.B(n_993),
.Y(n_1077)
);

BUFx6f_ASAP7_75t_L g1078 ( 
.A(n_1037),
.Y(n_1078)
);

OR2x2_ASAP7_75t_L g1079 ( 
.A(n_969),
.B(n_933),
.Y(n_1079)
);

AOI21xp5_ASAP7_75t_L g1080 ( 
.A1(n_1022),
.A2(n_1021),
.B(n_1043),
.Y(n_1080)
);

NAND2xp5_ASAP7_75t_L g1081 ( 
.A(n_895),
.B(n_1006),
.Y(n_1081)
);

OAI21xp5_ASAP7_75t_L g1082 ( 
.A1(n_914),
.A2(n_929),
.B(n_1015),
.Y(n_1082)
);

AOI21x1_ASAP7_75t_L g1083 ( 
.A1(n_973),
.A2(n_942),
.B(n_936),
.Y(n_1083)
);

INVx1_ASAP7_75t_SL g1084 ( 
.A(n_892),
.Y(n_1084)
);

AO31x2_ASAP7_75t_L g1085 ( 
.A1(n_890),
.A2(n_978),
.A3(n_981),
.B(n_1007),
.Y(n_1085)
);

OAI21x1_ASAP7_75t_SL g1086 ( 
.A1(n_971),
.A2(n_968),
.B(n_992),
.Y(n_1086)
);

BUFx3_ASAP7_75t_L g1087 ( 
.A(n_903),
.Y(n_1087)
);

AOI21x1_ASAP7_75t_L g1088 ( 
.A1(n_981),
.A2(n_921),
.B(n_924),
.Y(n_1088)
);

BUFx2_ASAP7_75t_L g1089 ( 
.A(n_892),
.Y(n_1089)
);

O2A1O1Ixp5_ASAP7_75t_L g1090 ( 
.A1(n_894),
.A2(n_1019),
.B(n_1003),
.C(n_952),
.Y(n_1090)
);

OAI21xp5_ASAP7_75t_L g1091 ( 
.A1(n_1014),
.A2(n_988),
.B(n_1021),
.Y(n_1091)
);

OAI22xp5_ASAP7_75t_L g1092 ( 
.A1(n_1027),
.A2(n_994),
.B1(n_910),
.B2(n_1007),
.Y(n_1092)
);

AOI21xp5_ASAP7_75t_L g1093 ( 
.A1(n_988),
.A2(n_945),
.B(n_911),
.Y(n_1093)
);

NAND2xp5_ASAP7_75t_L g1094 ( 
.A(n_1016),
.B(n_1017),
.Y(n_1094)
);

BUFx4_ASAP7_75t_SL g1095 ( 
.A(n_925),
.Y(n_1095)
);

INVx1_ASAP7_75t_L g1096 ( 
.A(n_997),
.Y(n_1096)
);

AND2x2_ASAP7_75t_L g1097 ( 
.A(n_987),
.B(n_916),
.Y(n_1097)
);

CKINVDCx5p33_ASAP7_75t_R g1098 ( 
.A(n_1018),
.Y(n_1098)
);

NAND2xp5_ASAP7_75t_L g1099 ( 
.A(n_995),
.B(n_998),
.Y(n_1099)
);

AOI21xp5_ASAP7_75t_L g1100 ( 
.A1(n_902),
.A2(n_893),
.B(n_1020),
.Y(n_1100)
);

AO31x2_ASAP7_75t_L g1101 ( 
.A1(n_991),
.A2(n_980),
.A3(n_954),
.B(n_960),
.Y(n_1101)
);

O2A1O1Ixp5_ASAP7_75t_L g1102 ( 
.A1(n_1013),
.A2(n_991),
.B(n_1025),
.C(n_1052),
.Y(n_1102)
);

NAND2x1p5_ASAP7_75t_L g1103 ( 
.A(n_902),
.B(n_983),
.Y(n_1103)
);

CKINVDCx5p33_ASAP7_75t_R g1104 ( 
.A(n_996),
.Y(n_1104)
);

OAI21xp5_ASAP7_75t_L g1105 ( 
.A1(n_899),
.A2(n_964),
.B(n_967),
.Y(n_1105)
);

NOR2xp33_ASAP7_75t_SL g1106 ( 
.A(n_957),
.B(n_961),
.Y(n_1106)
);

INVx3_ASAP7_75t_SL g1107 ( 
.A(n_1011),
.Y(n_1107)
);

A2O1A1Ixp33_ASAP7_75t_L g1108 ( 
.A1(n_913),
.A2(n_1008),
.B(n_1002),
.C(n_1004),
.Y(n_1108)
);

NAND3xp33_ASAP7_75t_L g1109 ( 
.A(n_946),
.B(n_901),
.C(n_955),
.Y(n_1109)
);

INVx3_ASAP7_75t_L g1110 ( 
.A(n_983),
.Y(n_1110)
);

NAND2xp5_ASAP7_75t_L g1111 ( 
.A(n_999),
.B(n_938),
.Y(n_1111)
);

AOI22xp5_ASAP7_75t_L g1112 ( 
.A1(n_1005),
.A2(n_931),
.B1(n_937),
.B2(n_923),
.Y(n_1112)
);

OAI21xp5_ASAP7_75t_L g1113 ( 
.A1(n_956),
.A2(n_1000),
.B(n_962),
.Y(n_1113)
);

OAI22x1_ASAP7_75t_L g1114 ( 
.A1(n_966),
.A2(n_939),
.B1(n_932),
.B2(n_1029),
.Y(n_1114)
);

AOI21xp5_ASAP7_75t_L g1115 ( 
.A1(n_902),
.A2(n_893),
.B(n_909),
.Y(n_1115)
);

AOI21xp5_ASAP7_75t_L g1116 ( 
.A1(n_909),
.A2(n_1040),
.B(n_1026),
.Y(n_1116)
);

AOI21xp5_ASAP7_75t_L g1117 ( 
.A1(n_1040),
.A2(n_1026),
.B(n_1046),
.Y(n_1117)
);

OAI22xp5_ASAP7_75t_L g1118 ( 
.A1(n_958),
.A2(n_961),
.B1(n_1042),
.B2(n_975),
.Y(n_1118)
);

INVx2_ASAP7_75t_SL g1119 ( 
.A(n_1048),
.Y(n_1119)
);

INVx2_ASAP7_75t_L g1120 ( 
.A(n_959),
.Y(n_1120)
);

OAI21xp5_ASAP7_75t_L g1121 ( 
.A1(n_972),
.A2(n_1012),
.B(n_951),
.Y(n_1121)
);

AOI21xp5_ASAP7_75t_L g1122 ( 
.A1(n_1028),
.A2(n_983),
.B(n_941),
.Y(n_1122)
);

NAND2xp5_ASAP7_75t_L g1123 ( 
.A(n_984),
.B(n_1037),
.Y(n_1123)
);

AND2x2_ASAP7_75t_L g1124 ( 
.A(n_1037),
.B(n_990),
.Y(n_1124)
);

NAND2xp5_ASAP7_75t_L g1125 ( 
.A(n_891),
.B(n_1042),
.Y(n_1125)
);

AOI21x1_ASAP7_75t_L g1126 ( 
.A1(n_974),
.A2(n_977),
.B(n_985),
.Y(n_1126)
);

NAND2xp5_ASAP7_75t_L g1127 ( 
.A(n_891),
.B(n_1042),
.Y(n_1127)
);

INVx2_ASAP7_75t_L g1128 ( 
.A(n_941),
.Y(n_1128)
);

NOR2xp33_ASAP7_75t_L g1129 ( 
.A(n_923),
.B(n_1001),
.Y(n_1129)
);

AO31x2_ASAP7_75t_L g1130 ( 
.A1(n_980),
.A2(n_982),
.A3(n_986),
.B(n_989),
.Y(n_1130)
);

INVx2_ASAP7_75t_L g1131 ( 
.A(n_989),
.Y(n_1131)
);

NAND2xp5_ASAP7_75t_L g1132 ( 
.A(n_957),
.B(n_944),
.Y(n_1132)
);

NAND2x1_ASAP7_75t_L g1133 ( 
.A(n_957),
.B(n_990),
.Y(n_1133)
);

INVx4_ASAP7_75t_L g1134 ( 
.A(n_957),
.Y(n_1134)
);

O2A1O1Ixp33_ASAP7_75t_SL g1135 ( 
.A1(n_943),
.A2(n_989),
.B(n_957),
.C(n_1010),
.Y(n_1135)
);

AOI21x1_ASAP7_75t_L g1136 ( 
.A1(n_943),
.A2(n_1010),
.B(n_906),
.Y(n_1136)
);

NAND2xp5_ASAP7_75t_L g1137 ( 
.A(n_943),
.B(n_1038),
.Y(n_1137)
);

INVx3_ASAP7_75t_L g1138 ( 
.A(n_983),
.Y(n_1138)
);

AOI22xp5_ASAP7_75t_L g1139 ( 
.A1(n_1030),
.A2(n_970),
.B1(n_935),
.B2(n_949),
.Y(n_1139)
);

BUFx6f_ASAP7_75t_L g1140 ( 
.A(n_1037),
.Y(n_1140)
);

BUFx2_ASAP7_75t_L g1141 ( 
.A(n_933),
.Y(n_1141)
);

OAI21x1_ASAP7_75t_L g1142 ( 
.A1(n_908),
.A2(n_1034),
.B(n_1032),
.Y(n_1142)
);

NAND2xp5_ASAP7_75t_SL g1143 ( 
.A(n_935),
.B(n_910),
.Y(n_1143)
);

NAND2xp5_ASAP7_75t_L g1144 ( 
.A(n_1038),
.B(n_1041),
.Y(n_1144)
);

AND2x4_ASAP7_75t_L g1145 ( 
.A(n_892),
.B(n_903),
.Y(n_1145)
);

AND2x2_ASAP7_75t_L g1146 ( 
.A(n_905),
.B(n_722),
.Y(n_1146)
);

OAI22xp5_ASAP7_75t_L g1147 ( 
.A1(n_1036),
.A2(n_1039),
.B1(n_1041),
.B2(n_1038),
.Y(n_1147)
);

OAI21x1_ASAP7_75t_L g1148 ( 
.A1(n_908),
.A2(n_1034),
.B(n_1032),
.Y(n_1148)
);

OR2x6_ASAP7_75t_L g1149 ( 
.A(n_900),
.B(n_889),
.Y(n_1149)
);

NAND2xp5_ASAP7_75t_L g1150 ( 
.A(n_1038),
.B(n_1041),
.Y(n_1150)
);

AND2x2_ASAP7_75t_L g1151 ( 
.A(n_905),
.B(n_722),
.Y(n_1151)
);

AOI21xp5_ASAP7_75t_L g1152 ( 
.A1(n_1038),
.A2(n_827),
.B(n_818),
.Y(n_1152)
);

INVx1_ASAP7_75t_SL g1153 ( 
.A(n_933),
.Y(n_1153)
);

AOI21xp5_ASAP7_75t_L g1154 ( 
.A1(n_1038),
.A2(n_827),
.B(n_818),
.Y(n_1154)
);

AO21x1_ASAP7_75t_L g1155 ( 
.A1(n_970),
.A2(n_949),
.B(n_1044),
.Y(n_1155)
);

INVx3_ASAP7_75t_L g1156 ( 
.A(n_983),
.Y(n_1156)
);

NAND2xp5_ASAP7_75t_L g1157 ( 
.A(n_1038),
.B(n_1041),
.Y(n_1157)
);

NAND3xp33_ASAP7_75t_L g1158 ( 
.A(n_949),
.B(n_755),
.C(n_970),
.Y(n_1158)
);

AOI21x1_ASAP7_75t_L g1159 ( 
.A1(n_940),
.A2(n_918),
.B(n_832),
.Y(n_1159)
);

AO21x2_ASAP7_75t_L g1160 ( 
.A1(n_914),
.A2(n_1039),
.B(n_929),
.Y(n_1160)
);

NAND2xp5_ASAP7_75t_L g1161 ( 
.A(n_1038),
.B(n_1041),
.Y(n_1161)
);

NOR2xp67_ASAP7_75t_L g1162 ( 
.A(n_910),
.B(n_662),
.Y(n_1162)
);

AO21x1_ASAP7_75t_L g1163 ( 
.A1(n_970),
.A2(n_949),
.B(n_1044),
.Y(n_1163)
);

OAI21xp5_ASAP7_75t_L g1164 ( 
.A1(n_1039),
.A2(n_1043),
.B(n_1035),
.Y(n_1164)
);

AOI22xp33_ASAP7_75t_L g1165 ( 
.A1(n_970),
.A2(n_949),
.B1(n_1030),
.B2(n_1036),
.Y(n_1165)
);

OAI21x1_ASAP7_75t_L g1166 ( 
.A1(n_908),
.A2(n_1034),
.B(n_1032),
.Y(n_1166)
);

INVx3_ASAP7_75t_L g1167 ( 
.A(n_983),
.Y(n_1167)
);

NAND2xp5_ASAP7_75t_L g1168 ( 
.A(n_1038),
.B(n_1041),
.Y(n_1168)
);

AO31x2_ASAP7_75t_L g1169 ( 
.A1(n_890),
.A2(n_930),
.A3(n_1039),
.B(n_1044),
.Y(n_1169)
);

NAND2xp5_ASAP7_75t_L g1170 ( 
.A(n_1038),
.B(n_1041),
.Y(n_1170)
);

INVx5_ASAP7_75t_L g1171 ( 
.A(n_957),
.Y(n_1171)
);

AND2x4_ASAP7_75t_L g1172 ( 
.A(n_892),
.B(n_903),
.Y(n_1172)
);

NAND2xp5_ASAP7_75t_L g1173 ( 
.A(n_1038),
.B(n_1041),
.Y(n_1173)
);

OAI21xp5_ASAP7_75t_L g1174 ( 
.A1(n_1039),
.A2(n_1043),
.B(n_1035),
.Y(n_1174)
);

INVx1_ASAP7_75t_L g1175 ( 
.A(n_963),
.Y(n_1175)
);

AND2x6_ASAP7_75t_L g1176 ( 
.A(n_983),
.B(n_1026),
.Y(n_1176)
);

NAND2xp5_ASAP7_75t_L g1177 ( 
.A(n_1038),
.B(n_1041),
.Y(n_1177)
);

NAND2xp5_ASAP7_75t_L g1178 ( 
.A(n_1038),
.B(n_1041),
.Y(n_1178)
);

AND2x4_ASAP7_75t_L g1179 ( 
.A(n_892),
.B(n_903),
.Y(n_1179)
);

AOI21xp33_ASAP7_75t_L g1180 ( 
.A1(n_970),
.A2(n_1039),
.B(n_949),
.Y(n_1180)
);

AOI21xp5_ASAP7_75t_SL g1181 ( 
.A1(n_1039),
.A2(n_827),
.B(n_818),
.Y(n_1181)
);

OAI21x1_ASAP7_75t_L g1182 ( 
.A1(n_908),
.A2(n_1034),
.B(n_1032),
.Y(n_1182)
);

INVx1_ASAP7_75t_SL g1183 ( 
.A(n_933),
.Y(n_1183)
);

A2O1A1Ixp33_ASAP7_75t_L g1184 ( 
.A1(n_1039),
.A2(n_970),
.B(n_949),
.C(n_865),
.Y(n_1184)
);

AND2x4_ASAP7_75t_L g1185 ( 
.A(n_892),
.B(n_903),
.Y(n_1185)
);

NOR2x1_ASAP7_75t_SL g1186 ( 
.A(n_902),
.B(n_983),
.Y(n_1186)
);

A2O1A1Ixp33_ASAP7_75t_L g1187 ( 
.A1(n_1039),
.A2(n_970),
.B(n_949),
.C(n_865),
.Y(n_1187)
);

OAI21x1_ASAP7_75t_SL g1188 ( 
.A1(n_930),
.A2(n_971),
.B(n_1023),
.Y(n_1188)
);

A2O1A1Ixp33_ASAP7_75t_L g1189 ( 
.A1(n_1039),
.A2(n_970),
.B(n_949),
.C(n_865),
.Y(n_1189)
);

NAND2xp5_ASAP7_75t_L g1190 ( 
.A(n_1038),
.B(n_1041),
.Y(n_1190)
);

NAND2xp5_ASAP7_75t_L g1191 ( 
.A(n_1038),
.B(n_1041),
.Y(n_1191)
);

BUFx3_ASAP7_75t_L g1192 ( 
.A(n_1141),
.Y(n_1192)
);

NAND2xp5_ASAP7_75t_SL g1193 ( 
.A(n_1139),
.B(n_1054),
.Y(n_1193)
);

AOI22xp33_ASAP7_75t_L g1194 ( 
.A1(n_1158),
.A2(n_1165),
.B1(n_1180),
.B2(n_1057),
.Y(n_1194)
);

OAI22xp5_ASAP7_75t_L g1195 ( 
.A1(n_1144),
.A2(n_1161),
.B1(n_1168),
.B2(n_1170),
.Y(n_1195)
);

NAND2xp5_ASAP7_75t_L g1196 ( 
.A(n_1173),
.B(n_1177),
.Y(n_1196)
);

OR2x6_ASAP7_75t_SL g1197 ( 
.A(n_1098),
.B(n_1104),
.Y(n_1197)
);

NAND2xp5_ASAP7_75t_L g1198 ( 
.A(n_1178),
.B(n_1150),
.Y(n_1198)
);

AND2x4_ASAP7_75t_L g1199 ( 
.A(n_1145),
.B(n_1172),
.Y(n_1199)
);

INVx3_ASAP7_75t_L g1200 ( 
.A(n_1134),
.Y(n_1200)
);

AOI21xp5_ASAP7_75t_L g1201 ( 
.A1(n_1053),
.A2(n_1157),
.B(n_1150),
.Y(n_1201)
);

AOI21xp5_ASAP7_75t_L g1202 ( 
.A1(n_1157),
.A2(n_1191),
.B(n_1190),
.Y(n_1202)
);

BUFx6f_ASAP7_75t_L g1203 ( 
.A(n_1078),
.Y(n_1203)
);

O2A1O1Ixp5_ASAP7_75t_L g1204 ( 
.A1(n_1180),
.A2(n_1057),
.B(n_1163),
.C(n_1155),
.Y(n_1204)
);

HB1xp67_ASAP7_75t_L g1205 ( 
.A(n_1153),
.Y(n_1205)
);

AOI21xp5_ASAP7_75t_L g1206 ( 
.A1(n_1190),
.A2(n_1191),
.B(n_1065),
.Y(n_1206)
);

BUFx3_ASAP7_75t_L g1207 ( 
.A(n_1087),
.Y(n_1207)
);

AOI21xp5_ASAP7_75t_L g1208 ( 
.A1(n_1059),
.A2(n_1080),
.B(n_1184),
.Y(n_1208)
);

INVx2_ASAP7_75t_L g1209 ( 
.A(n_1075),
.Y(n_1209)
);

NAND2x1p5_ASAP7_75t_L g1210 ( 
.A(n_1171),
.B(n_1134),
.Y(n_1210)
);

AND2x2_ASAP7_75t_L g1211 ( 
.A(n_1146),
.B(n_1151),
.Y(n_1211)
);

INVx1_ASAP7_75t_L g1212 ( 
.A(n_1096),
.Y(n_1212)
);

INVx2_ASAP7_75t_L g1213 ( 
.A(n_1120),
.Y(n_1213)
);

BUFx3_ASAP7_75t_L g1214 ( 
.A(n_1063),
.Y(n_1214)
);

AND2x2_ASAP7_75t_L g1215 ( 
.A(n_1076),
.B(n_1097),
.Y(n_1215)
);

AND2x2_ASAP7_75t_L g1216 ( 
.A(n_1089),
.B(n_1084),
.Y(n_1216)
);

AND2x4_ASAP7_75t_L g1217 ( 
.A(n_1145),
.B(n_1172),
.Y(n_1217)
);

BUFx3_ASAP7_75t_L g1218 ( 
.A(n_1079),
.Y(n_1218)
);

AND2x4_ASAP7_75t_L g1219 ( 
.A(n_1179),
.B(n_1185),
.Y(n_1219)
);

NOR2xp67_ASAP7_75t_SL g1220 ( 
.A(n_1171),
.B(n_1069),
.Y(n_1220)
);

HB1xp67_ASAP7_75t_L g1221 ( 
.A(n_1153),
.Y(n_1221)
);

OAI22xp5_ASAP7_75t_L g1222 ( 
.A1(n_1081),
.A2(n_1189),
.B1(n_1187),
.B2(n_1069),
.Y(n_1222)
);

NAND2xp5_ASAP7_75t_L g1223 ( 
.A(n_1071),
.B(n_1070),
.Y(n_1223)
);

BUFx6f_ASAP7_75t_L g1224 ( 
.A(n_1078),
.Y(n_1224)
);

INVx2_ASAP7_75t_L g1225 ( 
.A(n_1061),
.Y(n_1225)
);

AND2x4_ASAP7_75t_L g1226 ( 
.A(n_1179),
.B(n_1185),
.Y(n_1226)
);

AND2x4_ASAP7_75t_L g1227 ( 
.A(n_1124),
.B(n_1128),
.Y(n_1227)
);

CKINVDCx16_ASAP7_75t_R g1228 ( 
.A(n_1149),
.Y(n_1228)
);

OR2x6_ASAP7_75t_L g1229 ( 
.A(n_1133),
.B(n_1149),
.Y(n_1229)
);

NOR2xp33_ASAP7_75t_SL g1230 ( 
.A(n_1171),
.B(n_1106),
.Y(n_1230)
);

OAI22xp5_ASAP7_75t_L g1231 ( 
.A1(n_1070),
.A2(n_1099),
.B1(n_1147),
.B2(n_1056),
.Y(n_1231)
);

AOI21xp5_ASAP7_75t_L g1232 ( 
.A1(n_1091),
.A2(n_1077),
.B(n_1147),
.Y(n_1232)
);

NAND2xp5_ASAP7_75t_L g1233 ( 
.A(n_1071),
.B(n_1175),
.Y(n_1233)
);

INVx1_ASAP7_75t_L g1234 ( 
.A(n_1094),
.Y(n_1234)
);

NAND2xp5_ASAP7_75t_L g1235 ( 
.A(n_1074),
.B(n_1094),
.Y(n_1235)
);

INVx3_ASAP7_75t_L g1236 ( 
.A(n_1103),
.Y(n_1236)
);

NAND2xp5_ASAP7_75t_L g1237 ( 
.A(n_1074),
.B(n_1072),
.Y(n_1237)
);

NAND2xp5_ASAP7_75t_L g1238 ( 
.A(n_1072),
.B(n_1108),
.Y(n_1238)
);

OAI31xp33_ASAP7_75t_L g1239 ( 
.A1(n_1109),
.A2(n_1129),
.A3(n_1092),
.B(n_1118),
.Y(n_1239)
);

NOR2xp33_ASAP7_75t_SL g1240 ( 
.A(n_1171),
.B(n_1106),
.Y(n_1240)
);

AND2x4_ASAP7_75t_L g1241 ( 
.A(n_1084),
.B(n_1123),
.Y(n_1241)
);

NAND2x1_ASAP7_75t_L g1242 ( 
.A(n_1176),
.B(n_1110),
.Y(n_1242)
);

OR2x6_ASAP7_75t_L g1243 ( 
.A(n_1149),
.B(n_1068),
.Y(n_1243)
);

HB1xp67_ASAP7_75t_L g1244 ( 
.A(n_1183),
.Y(n_1244)
);

AND2x4_ASAP7_75t_L g1245 ( 
.A(n_1140),
.B(n_1119),
.Y(n_1245)
);

INVx1_ASAP7_75t_SL g1246 ( 
.A(n_1183),
.Y(n_1246)
);

INVx1_ASAP7_75t_SL g1247 ( 
.A(n_1095),
.Y(n_1247)
);

BUFx6f_ASAP7_75t_L g1248 ( 
.A(n_1140),
.Y(n_1248)
);

NAND2xp5_ASAP7_75t_L g1249 ( 
.A(n_1092),
.B(n_1164),
.Y(n_1249)
);

NAND2xp5_ASAP7_75t_L g1250 ( 
.A(n_1164),
.B(n_1174),
.Y(n_1250)
);

AND2x4_ASAP7_75t_L g1251 ( 
.A(n_1140),
.B(n_1125),
.Y(n_1251)
);

AOI22xp33_ASAP7_75t_L g1252 ( 
.A1(n_1066),
.A2(n_1118),
.B1(n_1143),
.B2(n_1086),
.Y(n_1252)
);

CKINVDCx16_ASAP7_75t_R g1253 ( 
.A(n_1068),
.Y(n_1253)
);

OAI21xp33_ASAP7_75t_L g1254 ( 
.A1(n_1112),
.A2(n_1066),
.B(n_1111),
.Y(n_1254)
);

INVx2_ASAP7_75t_SL g1255 ( 
.A(n_1068),
.Y(n_1255)
);

INVxp67_ASAP7_75t_SL g1256 ( 
.A(n_1186),
.Y(n_1256)
);

NOR2xp33_ASAP7_75t_L g1257 ( 
.A(n_1132),
.B(n_1162),
.Y(n_1257)
);

NAND2xp33_ASAP7_75t_L g1258 ( 
.A(n_1132),
.B(n_1176),
.Y(n_1258)
);

OR2x2_ASAP7_75t_L g1259 ( 
.A(n_1127),
.B(n_1101),
.Y(n_1259)
);

BUFx2_ASAP7_75t_SL g1260 ( 
.A(n_1138),
.Y(n_1260)
);

NAND2xp5_ASAP7_75t_SL g1261 ( 
.A(n_1102),
.B(n_1114),
.Y(n_1261)
);

BUFx2_ASAP7_75t_L g1262 ( 
.A(n_1156),
.Y(n_1262)
);

BUFx6f_ASAP7_75t_L g1263 ( 
.A(n_1103),
.Y(n_1263)
);

HB1xp67_ASAP7_75t_L g1264 ( 
.A(n_1156),
.Y(n_1264)
);

OR2x2_ASAP7_75t_SL g1265 ( 
.A(n_1107),
.B(n_1137),
.Y(n_1265)
);

NAND2x1_ASAP7_75t_L g1266 ( 
.A(n_1176),
.B(n_1167),
.Y(n_1266)
);

NAND2xp5_ASAP7_75t_L g1267 ( 
.A(n_1174),
.B(n_1058),
.Y(n_1267)
);

INVx3_ASAP7_75t_SL g1268 ( 
.A(n_1176),
.Y(n_1268)
);

AND2x2_ASAP7_75t_L g1269 ( 
.A(n_1122),
.B(n_1105),
.Y(n_1269)
);

BUFx6f_ASAP7_75t_L g1270 ( 
.A(n_1136),
.Y(n_1270)
);

CKINVDCx20_ASAP7_75t_R g1271 ( 
.A(n_1105),
.Y(n_1271)
);

INVx4_ASAP7_75t_L g1272 ( 
.A(n_1055),
.Y(n_1272)
);

INVx5_ASAP7_75t_L g1273 ( 
.A(n_1131),
.Y(n_1273)
);

NAND2xp5_ASAP7_75t_SL g1274 ( 
.A(n_1090),
.B(n_1113),
.Y(n_1274)
);

INVx1_ASAP7_75t_SL g1275 ( 
.A(n_1055),
.Y(n_1275)
);

AND2x2_ASAP7_75t_L g1276 ( 
.A(n_1169),
.B(n_1085),
.Y(n_1276)
);

NOR2xp67_ASAP7_75t_R g1277 ( 
.A(n_1073),
.B(n_1188),
.Y(n_1277)
);

NOR2xp33_ASAP7_75t_R g1278 ( 
.A(n_1126),
.B(n_1159),
.Y(n_1278)
);

AND2x4_ASAP7_75t_L g1279 ( 
.A(n_1117),
.B(n_1116),
.Y(n_1279)
);

INVx2_ASAP7_75t_L g1280 ( 
.A(n_1085),
.Y(n_1280)
);

AND2x4_ASAP7_75t_L g1281 ( 
.A(n_1121),
.B(n_1115),
.Y(n_1281)
);

OR2x2_ASAP7_75t_L g1282 ( 
.A(n_1137),
.B(n_1085),
.Y(n_1282)
);

OR2x6_ASAP7_75t_L g1283 ( 
.A(n_1181),
.B(n_1100),
.Y(n_1283)
);

NAND2xp5_ASAP7_75t_L g1284 ( 
.A(n_1160),
.B(n_1082),
.Y(n_1284)
);

BUFx10_ASAP7_75t_L g1285 ( 
.A(n_1130),
.Y(n_1285)
);

BUFx3_ASAP7_75t_L g1286 ( 
.A(n_1060),
.Y(n_1286)
);

INVx2_ASAP7_75t_SL g1287 ( 
.A(n_1160),
.Y(n_1287)
);

BUFx6f_ASAP7_75t_L g1288 ( 
.A(n_1083),
.Y(n_1288)
);

INVx1_ASAP7_75t_L g1289 ( 
.A(n_1135),
.Y(n_1289)
);

AOI22xp5_ASAP7_75t_L g1290 ( 
.A1(n_1152),
.A2(n_1154),
.B1(n_1067),
.B2(n_1148),
.Y(n_1290)
);

NAND2xp5_ASAP7_75t_L g1291 ( 
.A(n_1064),
.B(n_1088),
.Y(n_1291)
);

AOI21xp33_ASAP7_75t_L g1292 ( 
.A1(n_1142),
.A2(n_1166),
.B(n_1182),
.Y(n_1292)
);

INVx1_ASAP7_75t_L g1293 ( 
.A(n_1062),
.Y(n_1293)
);

AOI21xp5_ASAP7_75t_L g1294 ( 
.A1(n_1053),
.A2(n_1144),
.B(n_1054),
.Y(n_1294)
);

OA21x2_ASAP7_75t_L g1295 ( 
.A1(n_1082),
.A2(n_1091),
.B(n_1093),
.Y(n_1295)
);

NAND2xp5_ASAP7_75t_L g1296 ( 
.A(n_1054),
.B(n_1144),
.Y(n_1296)
);

INVx2_ASAP7_75t_SL g1297 ( 
.A(n_1087),
.Y(n_1297)
);

INVx3_ASAP7_75t_L g1298 ( 
.A(n_1134),
.Y(n_1298)
);

BUFx3_ASAP7_75t_L g1299 ( 
.A(n_1141),
.Y(n_1299)
);

OR2x6_ASAP7_75t_L g1300 ( 
.A(n_1133),
.B(n_1134),
.Y(n_1300)
);

HB1xp67_ASAP7_75t_L g1301 ( 
.A(n_1153),
.Y(n_1301)
);

INVxp67_ASAP7_75t_SL g1302 ( 
.A(n_1054),
.Y(n_1302)
);

CKINVDCx5p33_ASAP7_75t_R g1303 ( 
.A(n_1095),
.Y(n_1303)
);

INVx1_ASAP7_75t_L g1304 ( 
.A(n_1062),
.Y(n_1304)
);

NAND2xp5_ASAP7_75t_L g1305 ( 
.A(n_1054),
.B(n_1144),
.Y(n_1305)
);

NOR2xp33_ASAP7_75t_L g1306 ( 
.A(n_1158),
.B(n_734),
.Y(n_1306)
);

A2O1A1Ixp33_ASAP7_75t_SL g1307 ( 
.A1(n_1180),
.A2(n_970),
.B(n_949),
.C(n_1057),
.Y(n_1307)
);

OAI22xp5_ASAP7_75t_L g1308 ( 
.A1(n_1054),
.A2(n_1161),
.B1(n_1168),
.B2(n_1144),
.Y(n_1308)
);

A2O1A1Ixp33_ASAP7_75t_L g1309 ( 
.A1(n_1158),
.A2(n_1039),
.B(n_1187),
.C(n_1184),
.Y(n_1309)
);

INVx2_ASAP7_75t_L g1310 ( 
.A(n_1075),
.Y(n_1310)
);

BUFx3_ASAP7_75t_L g1311 ( 
.A(n_1141),
.Y(n_1311)
);

O2A1O1Ixp5_ASAP7_75t_L g1312 ( 
.A1(n_1180),
.A2(n_1158),
.B(n_1057),
.C(n_1155),
.Y(n_1312)
);

O2A1O1Ixp33_ASAP7_75t_L g1313 ( 
.A1(n_1180),
.A2(n_1039),
.B(n_1187),
.C(n_1184),
.Y(n_1313)
);

OAI22xp5_ASAP7_75t_L g1314 ( 
.A1(n_1054),
.A2(n_1161),
.B1(n_1168),
.B2(n_1144),
.Y(n_1314)
);

BUFx2_ASAP7_75t_L g1315 ( 
.A(n_1141),
.Y(n_1315)
);

NAND2xp5_ASAP7_75t_L g1316 ( 
.A(n_1054),
.B(n_1144),
.Y(n_1316)
);

BUFx6f_ASAP7_75t_L g1317 ( 
.A(n_1078),
.Y(n_1317)
);

BUFx3_ASAP7_75t_L g1318 ( 
.A(n_1141),
.Y(n_1318)
);

OAI22xp33_ASAP7_75t_L g1319 ( 
.A1(n_1158),
.A2(n_1106),
.B1(n_1069),
.B2(n_1139),
.Y(n_1319)
);

AND2x2_ASAP7_75t_L g1320 ( 
.A(n_1146),
.B(n_1151),
.Y(n_1320)
);

NOR2xp33_ASAP7_75t_R g1321 ( 
.A(n_1104),
.B(n_651),
.Y(n_1321)
);

BUFx3_ASAP7_75t_L g1322 ( 
.A(n_1141),
.Y(n_1322)
);

NOR2xp33_ASAP7_75t_SL g1323 ( 
.A(n_1171),
.B(n_1134),
.Y(n_1323)
);

AND2x2_ASAP7_75t_L g1324 ( 
.A(n_1146),
.B(n_1151),
.Y(n_1324)
);

BUFx2_ASAP7_75t_L g1325 ( 
.A(n_1141),
.Y(n_1325)
);

BUFx6f_ASAP7_75t_L g1326 ( 
.A(n_1078),
.Y(n_1326)
);

CKINVDCx14_ASAP7_75t_R g1327 ( 
.A(n_1321),
.Y(n_1327)
);

NAND2xp5_ASAP7_75t_L g1328 ( 
.A(n_1302),
.B(n_1196),
.Y(n_1328)
);

NAND2x1p5_ASAP7_75t_L g1329 ( 
.A(n_1220),
.B(n_1269),
.Y(n_1329)
);

AOI22xp33_ASAP7_75t_L g1330 ( 
.A1(n_1239),
.A2(n_1319),
.B1(n_1271),
.B2(n_1194),
.Y(n_1330)
);

NAND2x1p5_ASAP7_75t_L g1331 ( 
.A(n_1273),
.B(n_1275),
.Y(n_1331)
);

AOI22xp33_ASAP7_75t_L g1332 ( 
.A1(n_1222),
.A2(n_1193),
.B1(n_1306),
.B2(n_1252),
.Y(n_1332)
);

CKINVDCx20_ASAP7_75t_R g1333 ( 
.A(n_1303),
.Y(n_1333)
);

AOI22xp33_ASAP7_75t_L g1334 ( 
.A1(n_1222),
.A2(n_1254),
.B1(n_1249),
.B2(n_1257),
.Y(n_1334)
);

CKINVDCx11_ASAP7_75t_R g1335 ( 
.A(n_1197),
.Y(n_1335)
);

OR2x2_ASAP7_75t_L g1336 ( 
.A(n_1237),
.B(n_1250),
.Y(n_1336)
);

OA21x2_ASAP7_75t_L g1337 ( 
.A1(n_1204),
.A2(n_1291),
.B(n_1208),
.Y(n_1337)
);

AOI22xp33_ASAP7_75t_SL g1338 ( 
.A1(n_1230),
.A2(n_1240),
.B1(n_1249),
.B2(n_1253),
.Y(n_1338)
);

AND2x4_ASAP7_75t_L g1339 ( 
.A(n_1229),
.B(n_1300),
.Y(n_1339)
);

BUFx4f_ASAP7_75t_SL g1340 ( 
.A(n_1247),
.Y(n_1340)
);

CKINVDCx20_ASAP7_75t_R g1341 ( 
.A(n_1247),
.Y(n_1341)
);

AND2x2_ASAP7_75t_L g1342 ( 
.A(n_1198),
.B(n_1196),
.Y(n_1342)
);

INVx4_ASAP7_75t_L g1343 ( 
.A(n_1268),
.Y(n_1343)
);

BUFx2_ASAP7_75t_L g1344 ( 
.A(n_1205),
.Y(n_1344)
);

INVx1_ASAP7_75t_SL g1345 ( 
.A(n_1246),
.Y(n_1345)
);

OAI22xp5_ASAP7_75t_L g1346 ( 
.A1(n_1296),
.A2(n_1305),
.B1(n_1316),
.B2(n_1198),
.Y(n_1346)
);

HB1xp67_ASAP7_75t_L g1347 ( 
.A(n_1221),
.Y(n_1347)
);

OAI22xp33_ASAP7_75t_L g1348 ( 
.A1(n_1230),
.A2(n_1240),
.B1(n_1296),
.B2(n_1305),
.Y(n_1348)
);

INVx2_ASAP7_75t_L g1349 ( 
.A(n_1212),
.Y(n_1349)
);

INVx2_ASAP7_75t_L g1350 ( 
.A(n_1293),
.Y(n_1350)
);

HB1xp67_ASAP7_75t_L g1351 ( 
.A(n_1244),
.Y(n_1351)
);

INVx2_ASAP7_75t_L g1352 ( 
.A(n_1304),
.Y(n_1352)
);

INVx1_ASAP7_75t_L g1353 ( 
.A(n_1209),
.Y(n_1353)
);

INVx1_ASAP7_75t_L g1354 ( 
.A(n_1213),
.Y(n_1354)
);

HB1xp67_ASAP7_75t_L g1355 ( 
.A(n_1301),
.Y(n_1355)
);

AND2x2_ASAP7_75t_L g1356 ( 
.A(n_1195),
.B(n_1308),
.Y(n_1356)
);

NAND2xp5_ASAP7_75t_L g1357 ( 
.A(n_1233),
.B(n_1314),
.Y(n_1357)
);

AOI22xp33_ASAP7_75t_SL g1358 ( 
.A1(n_1323),
.A2(n_1228),
.B1(n_1238),
.B2(n_1231),
.Y(n_1358)
);

INVx2_ASAP7_75t_L g1359 ( 
.A(n_1234),
.Y(n_1359)
);

BUFx2_ASAP7_75t_L g1360 ( 
.A(n_1241),
.Y(n_1360)
);

AOI22xp5_ASAP7_75t_L g1361 ( 
.A1(n_1211),
.A2(n_1320),
.B1(n_1324),
.B2(n_1255),
.Y(n_1361)
);

AOI22xp33_ASAP7_75t_SL g1362 ( 
.A1(n_1323),
.A2(n_1238),
.B1(n_1231),
.B2(n_1233),
.Y(n_1362)
);

OAI22xp33_ASAP7_75t_L g1363 ( 
.A1(n_1218),
.A2(n_1223),
.B1(n_1243),
.B2(n_1235),
.Y(n_1363)
);

INVx6_ASAP7_75t_L g1364 ( 
.A(n_1199),
.Y(n_1364)
);

NAND2x1_ASAP7_75t_L g1365 ( 
.A(n_1283),
.B(n_1279),
.Y(n_1365)
);

BUFx2_ASAP7_75t_L g1366 ( 
.A(n_1241),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_1310),
.Y(n_1367)
);

BUFx6f_ASAP7_75t_L g1368 ( 
.A(n_1300),
.Y(n_1368)
);

AND2x4_ASAP7_75t_L g1369 ( 
.A(n_1229),
.B(n_1300),
.Y(n_1369)
);

CKINVDCx20_ASAP7_75t_R g1370 ( 
.A(n_1207),
.Y(n_1370)
);

AOI22xp33_ASAP7_75t_SL g1371 ( 
.A1(n_1215),
.A2(n_1267),
.B1(n_1250),
.B2(n_1243),
.Y(n_1371)
);

BUFx2_ASAP7_75t_L g1372 ( 
.A(n_1273),
.Y(n_1372)
);

OA21x2_ASAP7_75t_L g1373 ( 
.A1(n_1208),
.A2(n_1274),
.B(n_1312),
.Y(n_1373)
);

AND2x4_ASAP7_75t_L g1374 ( 
.A(n_1229),
.B(n_1200),
.Y(n_1374)
);

AND2x2_ASAP7_75t_L g1375 ( 
.A(n_1235),
.B(n_1202),
.Y(n_1375)
);

INVx1_ASAP7_75t_L g1376 ( 
.A(n_1264),
.Y(n_1376)
);

INVx3_ASAP7_75t_L g1377 ( 
.A(n_1200),
.Y(n_1377)
);

AOI22xp33_ASAP7_75t_L g1378 ( 
.A1(n_1261),
.A2(n_1237),
.B1(n_1227),
.B2(n_1232),
.Y(n_1378)
);

OR2x6_ASAP7_75t_L g1379 ( 
.A(n_1283),
.B(n_1201),
.Y(n_1379)
);

BUFx2_ASAP7_75t_L g1380 ( 
.A(n_1273),
.Y(n_1380)
);

OAI22xp5_ASAP7_75t_L g1381 ( 
.A1(n_1309),
.A2(n_1315),
.B1(n_1325),
.B2(n_1192),
.Y(n_1381)
);

BUFx2_ASAP7_75t_L g1382 ( 
.A(n_1273),
.Y(n_1382)
);

AOI22xp33_ASAP7_75t_L g1383 ( 
.A1(n_1227),
.A2(n_1232),
.B1(n_1267),
.B2(n_1216),
.Y(n_1383)
);

BUFx6f_ASAP7_75t_L g1384 ( 
.A(n_1263),
.Y(n_1384)
);

BUFx2_ASAP7_75t_L g1385 ( 
.A(n_1289),
.Y(n_1385)
);

OA21x2_ASAP7_75t_L g1386 ( 
.A1(n_1292),
.A2(n_1206),
.B(n_1294),
.Y(n_1386)
);

INVx2_ASAP7_75t_L g1387 ( 
.A(n_1288),
.Y(n_1387)
);

AND2x2_ASAP7_75t_L g1388 ( 
.A(n_1276),
.B(n_1259),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_1262),
.Y(n_1389)
);

HB1xp67_ASAP7_75t_L g1390 ( 
.A(n_1299),
.Y(n_1390)
);

INVx2_ASAP7_75t_L g1391 ( 
.A(n_1288),
.Y(n_1391)
);

INVx1_ASAP7_75t_L g1392 ( 
.A(n_1251),
.Y(n_1392)
);

INVx2_ASAP7_75t_L g1393 ( 
.A(n_1288),
.Y(n_1393)
);

OAI22xp5_ASAP7_75t_L g1394 ( 
.A1(n_1311),
.A2(n_1322),
.B1(n_1318),
.B2(n_1243),
.Y(n_1394)
);

INVx1_ASAP7_75t_L g1395 ( 
.A(n_1251),
.Y(n_1395)
);

CKINVDCx5p33_ASAP7_75t_R g1396 ( 
.A(n_1214),
.Y(n_1396)
);

INVx1_ASAP7_75t_L g1397 ( 
.A(n_1260),
.Y(n_1397)
);

BUFx4f_ASAP7_75t_SL g1398 ( 
.A(n_1297),
.Y(n_1398)
);

INVx6_ASAP7_75t_L g1399 ( 
.A(n_1217),
.Y(n_1399)
);

BUFx6f_ASAP7_75t_L g1400 ( 
.A(n_1263),
.Y(n_1400)
);

OA21x2_ASAP7_75t_L g1401 ( 
.A1(n_1292),
.A2(n_1206),
.B(n_1294),
.Y(n_1401)
);

AND2x2_ASAP7_75t_L g1402 ( 
.A(n_1282),
.B(n_1280),
.Y(n_1402)
);

INVx2_ASAP7_75t_L g1403 ( 
.A(n_1295),
.Y(n_1403)
);

AOI22xp33_ASAP7_75t_L g1404 ( 
.A1(n_1270),
.A2(n_1226),
.B1(n_1217),
.B2(n_1219),
.Y(n_1404)
);

NAND2x1p5_ASAP7_75t_L g1405 ( 
.A(n_1275),
.B(n_1272),
.Y(n_1405)
);

INVx1_ASAP7_75t_SL g1406 ( 
.A(n_1245),
.Y(n_1406)
);

INVx2_ASAP7_75t_L g1407 ( 
.A(n_1287),
.Y(n_1407)
);

INVx2_ASAP7_75t_L g1408 ( 
.A(n_1285),
.Y(n_1408)
);

BUFx3_ASAP7_75t_L g1409 ( 
.A(n_1219),
.Y(n_1409)
);

BUFx3_ASAP7_75t_L g1410 ( 
.A(n_1226),
.Y(n_1410)
);

INVx3_ASAP7_75t_L g1411 ( 
.A(n_1298),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_1284),
.Y(n_1412)
);

CKINVDCx11_ASAP7_75t_R g1413 ( 
.A(n_1203),
.Y(n_1413)
);

OAI21x1_ASAP7_75t_L g1414 ( 
.A1(n_1290),
.A2(n_1313),
.B(n_1298),
.Y(n_1414)
);

INVx2_ASAP7_75t_L g1415 ( 
.A(n_1285),
.Y(n_1415)
);

OAI21x1_ASAP7_75t_L g1416 ( 
.A1(n_1242),
.A2(n_1266),
.B(n_1236),
.Y(n_1416)
);

NAND2x1p5_ASAP7_75t_L g1417 ( 
.A(n_1272),
.B(n_1281),
.Y(n_1417)
);

AOI22xp33_ASAP7_75t_SL g1418 ( 
.A1(n_1270),
.A2(n_1258),
.B1(n_1256),
.B2(n_1307),
.Y(n_1418)
);

HB1xp67_ASAP7_75t_L g1419 ( 
.A(n_1245),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_1224),
.Y(n_1420)
);

AND2x2_ASAP7_75t_L g1421 ( 
.A(n_1236),
.B(n_1281),
.Y(n_1421)
);

HB1xp67_ASAP7_75t_L g1422 ( 
.A(n_1248),
.Y(n_1422)
);

BUFx3_ASAP7_75t_L g1423 ( 
.A(n_1326),
.Y(n_1423)
);

OAI22xp5_ASAP7_75t_L g1424 ( 
.A1(n_1283),
.A2(n_1265),
.B1(n_1279),
.B2(n_1248),
.Y(n_1424)
);

CKINVDCx20_ASAP7_75t_R g1425 ( 
.A(n_1248),
.Y(n_1425)
);

OAI22xp5_ASAP7_75t_L g1426 ( 
.A1(n_1317),
.A2(n_1326),
.B1(n_1286),
.B2(n_1277),
.Y(n_1426)
);

BUFx2_ASAP7_75t_L g1427 ( 
.A(n_1278),
.Y(n_1427)
);

BUFx8_ASAP7_75t_L g1428 ( 
.A(n_1317),
.Y(n_1428)
);

INVx1_ASAP7_75t_L g1429 ( 
.A(n_1225),
.Y(n_1429)
);

AOI22xp33_ASAP7_75t_L g1430 ( 
.A1(n_1239),
.A2(n_1158),
.B1(n_949),
.B2(n_1319),
.Y(n_1430)
);

BUFx3_ASAP7_75t_L g1431 ( 
.A(n_1207),
.Y(n_1431)
);

AND2x2_ASAP7_75t_L g1432 ( 
.A(n_1302),
.B(n_1198),
.Y(n_1432)
);

AOI22xp33_ASAP7_75t_L g1433 ( 
.A1(n_1239),
.A2(n_1158),
.B1(n_949),
.B2(n_1319),
.Y(n_1433)
);

NOR2xp67_ASAP7_75t_L g1434 ( 
.A(n_1225),
.B(n_662),
.Y(n_1434)
);

AOI22xp33_ASAP7_75t_SL g1435 ( 
.A1(n_1230),
.A2(n_946),
.B1(n_1106),
.B2(n_1240),
.Y(n_1435)
);

INVx1_ASAP7_75t_SL g1436 ( 
.A(n_1246),
.Y(n_1436)
);

AOI22xp33_ASAP7_75t_SL g1437 ( 
.A1(n_1230),
.A2(n_946),
.B1(n_1106),
.B2(n_1240),
.Y(n_1437)
);

INVx1_ASAP7_75t_L g1438 ( 
.A(n_1225),
.Y(n_1438)
);

INVx3_ASAP7_75t_L g1439 ( 
.A(n_1210),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_1225),
.Y(n_1440)
);

BUFx4_ASAP7_75t_R g1441 ( 
.A(n_1230),
.Y(n_1441)
);

INVx1_ASAP7_75t_SL g1442 ( 
.A(n_1246),
.Y(n_1442)
);

AND2x4_ASAP7_75t_L g1443 ( 
.A(n_1229),
.B(n_1300),
.Y(n_1443)
);

INVx2_ASAP7_75t_L g1444 ( 
.A(n_1225),
.Y(n_1444)
);

CKINVDCx5p33_ASAP7_75t_R g1445 ( 
.A(n_1303),
.Y(n_1445)
);

NAND2xp5_ASAP7_75t_L g1446 ( 
.A(n_1342),
.B(n_1432),
.Y(n_1446)
);

AND2x2_ASAP7_75t_L g1447 ( 
.A(n_1388),
.B(n_1375),
.Y(n_1447)
);

INVx2_ASAP7_75t_SL g1448 ( 
.A(n_1372),
.Y(n_1448)
);

NAND2xp5_ASAP7_75t_L g1449 ( 
.A(n_1342),
.B(n_1432),
.Y(n_1449)
);

HB1xp67_ASAP7_75t_L g1450 ( 
.A(n_1344),
.Y(n_1450)
);

AND2x2_ASAP7_75t_L g1451 ( 
.A(n_1388),
.B(n_1375),
.Y(n_1451)
);

BUFx2_ASAP7_75t_L g1452 ( 
.A(n_1385),
.Y(n_1452)
);

BUFx12f_ASAP7_75t_L g1453 ( 
.A(n_1445),
.Y(n_1453)
);

INVx1_ASAP7_75t_L g1454 ( 
.A(n_1412),
.Y(n_1454)
);

AND2x2_ASAP7_75t_L g1455 ( 
.A(n_1356),
.B(n_1402),
.Y(n_1455)
);

AND2x2_ASAP7_75t_L g1456 ( 
.A(n_1356),
.B(n_1402),
.Y(n_1456)
);

INVx3_ASAP7_75t_L g1457 ( 
.A(n_1331),
.Y(n_1457)
);

INVx2_ASAP7_75t_L g1458 ( 
.A(n_1403),
.Y(n_1458)
);

AND2x2_ASAP7_75t_L g1459 ( 
.A(n_1336),
.B(n_1421),
.Y(n_1459)
);

BUFx3_ASAP7_75t_L g1460 ( 
.A(n_1331),
.Y(n_1460)
);

AND2x2_ASAP7_75t_L g1461 ( 
.A(n_1336),
.B(n_1421),
.Y(n_1461)
);

HB1xp67_ASAP7_75t_L g1462 ( 
.A(n_1344),
.Y(n_1462)
);

INVxp33_ASAP7_75t_L g1463 ( 
.A(n_1390),
.Y(n_1463)
);

INVx1_ASAP7_75t_L g1464 ( 
.A(n_1405),
.Y(n_1464)
);

INVx1_ASAP7_75t_L g1465 ( 
.A(n_1405),
.Y(n_1465)
);

INVxp67_ASAP7_75t_L g1466 ( 
.A(n_1347),
.Y(n_1466)
);

OAI21xp5_ASAP7_75t_L g1467 ( 
.A1(n_1430),
.A2(n_1433),
.B(n_1332),
.Y(n_1467)
);

BUFx2_ASAP7_75t_SL g1468 ( 
.A(n_1434),
.Y(n_1468)
);

OR2x2_ASAP7_75t_L g1469 ( 
.A(n_1357),
.B(n_1417),
.Y(n_1469)
);

INVx1_ASAP7_75t_L g1470 ( 
.A(n_1405),
.Y(n_1470)
);

INVxp67_ASAP7_75t_SL g1471 ( 
.A(n_1328),
.Y(n_1471)
);

CKINVDCx20_ASAP7_75t_R g1472 ( 
.A(n_1333),
.Y(n_1472)
);

INVx1_ASAP7_75t_L g1473 ( 
.A(n_1407),
.Y(n_1473)
);

AND2x2_ASAP7_75t_L g1474 ( 
.A(n_1334),
.B(n_1373),
.Y(n_1474)
);

HB1xp67_ASAP7_75t_L g1475 ( 
.A(n_1351),
.Y(n_1475)
);

OR2x2_ASAP7_75t_L g1476 ( 
.A(n_1417),
.B(n_1337),
.Y(n_1476)
);

AND2x2_ASAP7_75t_L g1477 ( 
.A(n_1373),
.B(n_1349),
.Y(n_1477)
);

INVx2_ASAP7_75t_L g1478 ( 
.A(n_1337),
.Y(n_1478)
);

AND2x2_ASAP7_75t_L g1479 ( 
.A(n_1373),
.B(n_1349),
.Y(n_1479)
);

INVxp67_ASAP7_75t_L g1480 ( 
.A(n_1355),
.Y(n_1480)
);

INVx1_ASAP7_75t_L g1481 ( 
.A(n_1385),
.Y(n_1481)
);

HB1xp67_ASAP7_75t_L g1482 ( 
.A(n_1360),
.Y(n_1482)
);

INVx1_ASAP7_75t_L g1483 ( 
.A(n_1359),
.Y(n_1483)
);

BUFx4f_ASAP7_75t_SL g1484 ( 
.A(n_1333),
.Y(n_1484)
);

INVx1_ASAP7_75t_L g1485 ( 
.A(n_1359),
.Y(n_1485)
);

OAI21x1_ASAP7_75t_L g1486 ( 
.A1(n_1414),
.A2(n_1365),
.B(n_1386),
.Y(n_1486)
);

AND2x2_ASAP7_75t_L g1487 ( 
.A(n_1350),
.B(n_1352),
.Y(n_1487)
);

HB1xp67_ASAP7_75t_L g1488 ( 
.A(n_1360),
.Y(n_1488)
);

OAI21x1_ASAP7_75t_L g1489 ( 
.A1(n_1365),
.A2(n_1386),
.B(n_1401),
.Y(n_1489)
);

NAND2xp5_ASAP7_75t_SL g1490 ( 
.A(n_1346),
.B(n_1435),
.Y(n_1490)
);

INVx1_ASAP7_75t_L g1491 ( 
.A(n_1408),
.Y(n_1491)
);

BUFx6f_ASAP7_75t_L g1492 ( 
.A(n_1368),
.Y(n_1492)
);

NAND3xp33_ASAP7_75t_L g1493 ( 
.A(n_1330),
.B(n_1437),
.C(n_1358),
.Y(n_1493)
);

BUFx3_ASAP7_75t_L g1494 ( 
.A(n_1339),
.Y(n_1494)
);

INVxp67_ASAP7_75t_L g1495 ( 
.A(n_1345),
.Y(n_1495)
);

OAI21x1_ASAP7_75t_L g1496 ( 
.A1(n_1401),
.A2(n_1424),
.B(n_1415),
.Y(n_1496)
);

INVx1_ASAP7_75t_L g1497 ( 
.A(n_1408),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_1415),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_1379),
.Y(n_1499)
);

BUFx2_ASAP7_75t_L g1500 ( 
.A(n_1379),
.Y(n_1500)
);

INVx1_ASAP7_75t_L g1501 ( 
.A(n_1379),
.Y(n_1501)
);

OAI21xp5_ASAP7_75t_L g1502 ( 
.A1(n_1418),
.A2(n_1362),
.B(n_1378),
.Y(n_1502)
);

CKINVDCx5p33_ASAP7_75t_R g1503 ( 
.A(n_1445),
.Y(n_1503)
);

INVx4_ASAP7_75t_L g1504 ( 
.A(n_1441),
.Y(n_1504)
);

OAI21xp33_ASAP7_75t_SL g1505 ( 
.A1(n_1441),
.A2(n_1379),
.B(n_1383),
.Y(n_1505)
);

OR2x2_ASAP7_75t_L g1506 ( 
.A(n_1366),
.B(n_1329),
.Y(n_1506)
);

NAND2xp5_ASAP7_75t_L g1507 ( 
.A(n_1436),
.B(n_1442),
.Y(n_1507)
);

AO21x2_ASAP7_75t_L g1508 ( 
.A1(n_1363),
.A2(n_1348),
.B(n_1387),
.Y(n_1508)
);

BUFx3_ASAP7_75t_L g1509 ( 
.A(n_1339),
.Y(n_1509)
);

OAI21xp5_ASAP7_75t_L g1510 ( 
.A1(n_1381),
.A2(n_1329),
.B(n_1338),
.Y(n_1510)
);

AO31x2_ASAP7_75t_L g1511 ( 
.A1(n_1391),
.A2(n_1393),
.A3(n_1382),
.B(n_1380),
.Y(n_1511)
);

INVx3_ASAP7_75t_L g1512 ( 
.A(n_1368),
.Y(n_1512)
);

INVx3_ASAP7_75t_L g1513 ( 
.A(n_1368),
.Y(n_1513)
);

HB1xp67_ASAP7_75t_L g1514 ( 
.A(n_1366),
.Y(n_1514)
);

HB1xp67_ASAP7_75t_L g1515 ( 
.A(n_1376),
.Y(n_1515)
);

HB1xp67_ASAP7_75t_L g1516 ( 
.A(n_1389),
.Y(n_1516)
);

AND2x2_ASAP7_75t_L g1517 ( 
.A(n_1444),
.B(n_1329),
.Y(n_1517)
);

AND2x2_ASAP7_75t_L g1518 ( 
.A(n_1444),
.B(n_1429),
.Y(n_1518)
);

INVx3_ASAP7_75t_L g1519 ( 
.A(n_1368),
.Y(n_1519)
);

INVx1_ASAP7_75t_L g1520 ( 
.A(n_1438),
.Y(n_1520)
);

INVx2_ASAP7_75t_L g1521 ( 
.A(n_1440),
.Y(n_1521)
);

INVx1_ASAP7_75t_L g1522 ( 
.A(n_1353),
.Y(n_1522)
);

CKINVDCx5p33_ASAP7_75t_R g1523 ( 
.A(n_1335),
.Y(n_1523)
);

INVx1_ASAP7_75t_SL g1524 ( 
.A(n_1370),
.Y(n_1524)
);

INVx1_ASAP7_75t_L g1525 ( 
.A(n_1354),
.Y(n_1525)
);

INVx2_ASAP7_75t_L g1526 ( 
.A(n_1367),
.Y(n_1526)
);

NOR2xp33_ASAP7_75t_L g1527 ( 
.A(n_1340),
.B(n_1341),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_1339),
.Y(n_1528)
);

BUFx10_ASAP7_75t_L g1529 ( 
.A(n_1374),
.Y(n_1529)
);

INVx2_ASAP7_75t_L g1530 ( 
.A(n_1369),
.Y(n_1530)
);

INVx1_ASAP7_75t_L g1531 ( 
.A(n_1443),
.Y(n_1531)
);

HB1xp67_ASAP7_75t_L g1532 ( 
.A(n_1392),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_1369),
.Y(n_1533)
);

BUFx3_ASAP7_75t_L g1534 ( 
.A(n_1460),
.Y(n_1534)
);

AOI22xp33_ASAP7_75t_SL g1535 ( 
.A1(n_1467),
.A2(n_1443),
.B1(n_1369),
.B2(n_1427),
.Y(n_1535)
);

INVx1_ASAP7_75t_SL g1536 ( 
.A(n_1452),
.Y(n_1536)
);

BUFx2_ASAP7_75t_L g1537 ( 
.A(n_1460),
.Y(n_1537)
);

NAND2xp5_ASAP7_75t_L g1538 ( 
.A(n_1471),
.B(n_1447),
.Y(n_1538)
);

NOR2x1p5_ASAP7_75t_L g1539 ( 
.A(n_1504),
.B(n_1443),
.Y(n_1539)
);

AND2x4_ASAP7_75t_L g1540 ( 
.A(n_1499),
.B(n_1374),
.Y(n_1540)
);

AND2x2_ASAP7_75t_L g1541 ( 
.A(n_1477),
.B(n_1371),
.Y(n_1541)
);

INVxp67_ASAP7_75t_SL g1542 ( 
.A(n_1478),
.Y(n_1542)
);

AND2x2_ASAP7_75t_L g1543 ( 
.A(n_1477),
.B(n_1361),
.Y(n_1543)
);

NAND2xp5_ASAP7_75t_L g1544 ( 
.A(n_1447),
.B(n_1427),
.Y(n_1544)
);

AND2x2_ASAP7_75t_L g1545 ( 
.A(n_1479),
.B(n_1395),
.Y(n_1545)
);

INVx2_ASAP7_75t_SL g1546 ( 
.A(n_1511),
.Y(n_1546)
);

AND2x2_ASAP7_75t_L g1547 ( 
.A(n_1479),
.B(n_1374),
.Y(n_1547)
);

AND2x2_ASAP7_75t_L g1548 ( 
.A(n_1451),
.B(n_1411),
.Y(n_1548)
);

OR2x2_ASAP7_75t_L g1549 ( 
.A(n_1451),
.B(n_1394),
.Y(n_1549)
);

AND2x2_ASAP7_75t_L g1550 ( 
.A(n_1474),
.B(n_1377),
.Y(n_1550)
);

AND2x2_ASAP7_75t_L g1551 ( 
.A(n_1459),
.B(n_1397),
.Y(n_1551)
);

BUFx2_ASAP7_75t_L g1552 ( 
.A(n_1460),
.Y(n_1552)
);

AND2x2_ASAP7_75t_L g1553 ( 
.A(n_1474),
.B(n_1377),
.Y(n_1553)
);

BUFx3_ASAP7_75t_L g1554 ( 
.A(n_1452),
.Y(n_1554)
);

AND2x4_ASAP7_75t_SL g1555 ( 
.A(n_1529),
.B(n_1343),
.Y(n_1555)
);

AND2x2_ASAP7_75t_L g1556 ( 
.A(n_1459),
.B(n_1461),
.Y(n_1556)
);

NAND2xp5_ASAP7_75t_L g1557 ( 
.A(n_1446),
.B(n_1426),
.Y(n_1557)
);

NAND2xp5_ASAP7_75t_L g1558 ( 
.A(n_1449),
.B(n_1454),
.Y(n_1558)
);

AND2x2_ASAP7_75t_L g1559 ( 
.A(n_1461),
.B(n_1411),
.Y(n_1559)
);

INVx1_ASAP7_75t_SL g1560 ( 
.A(n_1450),
.Y(n_1560)
);

AND2x2_ASAP7_75t_L g1561 ( 
.A(n_1455),
.B(n_1411),
.Y(n_1561)
);

AND2x2_ASAP7_75t_L g1562 ( 
.A(n_1455),
.B(n_1377),
.Y(n_1562)
);

NAND2xp5_ASAP7_75t_L g1563 ( 
.A(n_1454),
.B(n_1419),
.Y(n_1563)
);

AND2x4_ASAP7_75t_L g1564 ( 
.A(n_1499),
.B(n_1416),
.Y(n_1564)
);

AND2x2_ASAP7_75t_L g1565 ( 
.A(n_1456),
.B(n_1420),
.Y(n_1565)
);

OAI22xp33_ASAP7_75t_L g1566 ( 
.A1(n_1493),
.A2(n_1409),
.B1(n_1410),
.B2(n_1343),
.Y(n_1566)
);

NAND2xp5_ASAP7_75t_SL g1567 ( 
.A(n_1504),
.B(n_1343),
.Y(n_1567)
);

HB1xp67_ASAP7_75t_L g1568 ( 
.A(n_1481),
.Y(n_1568)
);

AND2x4_ASAP7_75t_L g1569 ( 
.A(n_1501),
.B(n_1416),
.Y(n_1569)
);

AND2x2_ASAP7_75t_L g1570 ( 
.A(n_1530),
.B(n_1469),
.Y(n_1570)
);

AND2x2_ASAP7_75t_L g1571 ( 
.A(n_1530),
.B(n_1439),
.Y(n_1571)
);

INVx2_ASAP7_75t_SL g1572 ( 
.A(n_1511),
.Y(n_1572)
);

HB1xp67_ASAP7_75t_L g1573 ( 
.A(n_1511),
.Y(n_1573)
);

NOR2xp33_ASAP7_75t_L g1574 ( 
.A(n_1524),
.B(n_1341),
.Y(n_1574)
);

AND2x2_ASAP7_75t_L g1575 ( 
.A(n_1469),
.B(n_1439),
.Y(n_1575)
);

BUFx6f_ASAP7_75t_L g1576 ( 
.A(n_1496),
.Y(n_1576)
);

OAI22xp5_ASAP7_75t_L g1577 ( 
.A1(n_1535),
.A2(n_1504),
.B1(n_1490),
.B2(n_1502),
.Y(n_1577)
);

AND2x2_ASAP7_75t_L g1578 ( 
.A(n_1547),
.B(n_1500),
.Y(n_1578)
);

NAND3xp33_ASAP7_75t_L g1579 ( 
.A(n_1535),
.B(n_1510),
.C(n_1517),
.Y(n_1579)
);

NAND3xp33_ASAP7_75t_L g1580 ( 
.A(n_1557),
.B(n_1517),
.C(n_1501),
.Y(n_1580)
);

AND2x2_ASAP7_75t_L g1581 ( 
.A(n_1547),
.B(n_1476),
.Y(n_1581)
);

AND2x2_ASAP7_75t_SL g1582 ( 
.A(n_1537),
.B(n_1504),
.Y(n_1582)
);

NAND2xp5_ASAP7_75t_L g1583 ( 
.A(n_1538),
.B(n_1462),
.Y(n_1583)
);

NAND2xp5_ASAP7_75t_L g1584 ( 
.A(n_1538),
.B(n_1475),
.Y(n_1584)
);

OAI21xp5_ASAP7_75t_L g1585 ( 
.A1(n_1566),
.A2(n_1505),
.B(n_1463),
.Y(n_1585)
);

AND2x2_ASAP7_75t_L g1586 ( 
.A(n_1570),
.B(n_1476),
.Y(n_1586)
);

OAI221xp5_ASAP7_75t_L g1587 ( 
.A1(n_1567),
.A2(n_1505),
.B1(n_1468),
.B2(n_1557),
.C(n_1574),
.Y(n_1587)
);

NOR3xp33_ASAP7_75t_L g1588 ( 
.A(n_1566),
.B(n_1480),
.C(n_1466),
.Y(n_1588)
);

OAI21xp5_ASAP7_75t_SL g1589 ( 
.A1(n_1541),
.A2(n_1327),
.B(n_1527),
.Y(n_1589)
);

OA21x2_ASAP7_75t_L g1590 ( 
.A1(n_1542),
.A2(n_1489),
.B(n_1486),
.Y(n_1590)
);

NAND2xp5_ASAP7_75t_L g1591 ( 
.A(n_1544),
.B(n_1515),
.Y(n_1591)
);

NAND4xp25_ASAP7_75t_L g1592 ( 
.A(n_1560),
.B(n_1507),
.C(n_1495),
.D(n_1520),
.Y(n_1592)
);

NAND2xp5_ASAP7_75t_L g1593 ( 
.A(n_1544),
.B(n_1516),
.Y(n_1593)
);

NAND3xp33_ASAP7_75t_L g1594 ( 
.A(n_1576),
.B(n_1506),
.C(n_1465),
.Y(n_1594)
);

AND2x2_ASAP7_75t_L g1595 ( 
.A(n_1570),
.B(n_1496),
.Y(n_1595)
);

NAND2xp5_ASAP7_75t_L g1596 ( 
.A(n_1560),
.B(n_1482),
.Y(n_1596)
);

AOI21xp5_ASAP7_75t_SL g1597 ( 
.A1(n_1539),
.A2(n_1508),
.B(n_1523),
.Y(n_1597)
);

AND2x2_ASAP7_75t_L g1598 ( 
.A(n_1550),
.B(n_1464),
.Y(n_1598)
);

AND2x2_ASAP7_75t_L g1599 ( 
.A(n_1550),
.B(n_1464),
.Y(n_1599)
);

NAND2xp5_ASAP7_75t_L g1600 ( 
.A(n_1556),
.B(n_1488),
.Y(n_1600)
);

NAND2xp5_ASAP7_75t_L g1601 ( 
.A(n_1556),
.B(n_1514),
.Y(n_1601)
);

OAI221xp5_ASAP7_75t_SL g1602 ( 
.A1(n_1549),
.A2(n_1506),
.B1(n_1404),
.B2(n_1406),
.C(n_1528),
.Y(n_1602)
);

OAI221xp5_ASAP7_75t_SL g1603 ( 
.A1(n_1549),
.A2(n_1533),
.B1(n_1531),
.B2(n_1528),
.C(n_1494),
.Y(n_1603)
);

AOI21xp33_ASAP7_75t_SL g1604 ( 
.A1(n_1551),
.A2(n_1503),
.B(n_1396),
.Y(n_1604)
);

OAI221xp5_ASAP7_75t_L g1605 ( 
.A1(n_1563),
.A2(n_1468),
.B1(n_1533),
.B2(n_1531),
.C(n_1513),
.Y(n_1605)
);

OAI22xp5_ASAP7_75t_L g1606 ( 
.A1(n_1539),
.A2(n_1494),
.B1(n_1509),
.B2(n_1425),
.Y(n_1606)
);

OAI221xp5_ASAP7_75t_SL g1607 ( 
.A1(n_1541),
.A2(n_1536),
.B1(n_1543),
.B2(n_1558),
.C(n_1563),
.Y(n_1607)
);

OAI21xp5_ASAP7_75t_SL g1608 ( 
.A1(n_1541),
.A2(n_1335),
.B(n_1519),
.Y(n_1608)
);

NAND2xp5_ASAP7_75t_L g1609 ( 
.A(n_1558),
.B(n_1491),
.Y(n_1609)
);

AND2x2_ASAP7_75t_L g1610 ( 
.A(n_1553),
.B(n_1470),
.Y(n_1610)
);

AOI22xp5_ASAP7_75t_L g1611 ( 
.A1(n_1540),
.A2(n_1508),
.B1(n_1509),
.B2(n_1494),
.Y(n_1611)
);

NAND2xp5_ASAP7_75t_L g1612 ( 
.A(n_1543),
.B(n_1491),
.Y(n_1612)
);

AND2x2_ASAP7_75t_SL g1613 ( 
.A(n_1537),
.B(n_1492),
.Y(n_1613)
);

NAND3xp33_ASAP7_75t_L g1614 ( 
.A(n_1576),
.B(n_1470),
.C(n_1497),
.Y(n_1614)
);

OAI21xp33_ASAP7_75t_L g1615 ( 
.A1(n_1543),
.A2(n_1551),
.B(n_1575),
.Y(n_1615)
);

OAI21xp5_ASAP7_75t_L g1616 ( 
.A1(n_1564),
.A2(n_1486),
.B(n_1532),
.Y(n_1616)
);

AOI221xp5_ASAP7_75t_L g1617 ( 
.A1(n_1536),
.A2(n_1520),
.B1(n_1522),
.B2(n_1525),
.C(n_1497),
.Y(n_1617)
);

NAND2xp5_ASAP7_75t_L g1618 ( 
.A(n_1548),
.B(n_1498),
.Y(n_1618)
);

NAND2xp5_ASAP7_75t_L g1619 ( 
.A(n_1548),
.B(n_1498),
.Y(n_1619)
);

NOR2xp33_ASAP7_75t_L g1620 ( 
.A(n_1540),
.B(n_1575),
.Y(n_1620)
);

NAND2xp5_ASAP7_75t_L g1621 ( 
.A(n_1548),
.B(n_1487),
.Y(n_1621)
);

AND2x2_ASAP7_75t_L g1622 ( 
.A(n_1553),
.B(n_1458),
.Y(n_1622)
);

NAND2xp5_ASAP7_75t_SL g1623 ( 
.A(n_1540),
.B(n_1457),
.Y(n_1623)
);

NAND2xp5_ASAP7_75t_L g1624 ( 
.A(n_1559),
.B(n_1487),
.Y(n_1624)
);

NAND2xp5_ASAP7_75t_L g1625 ( 
.A(n_1559),
.B(n_1521),
.Y(n_1625)
);

NAND2xp5_ASAP7_75t_L g1626 ( 
.A(n_1545),
.B(n_1521),
.Y(n_1626)
);

NAND3xp33_ASAP7_75t_L g1627 ( 
.A(n_1576),
.B(n_1522),
.C(n_1525),
.Y(n_1627)
);

OAI21xp5_ASAP7_75t_SL g1628 ( 
.A1(n_1555),
.A2(n_1513),
.B(n_1512),
.Y(n_1628)
);

NAND2xp5_ASAP7_75t_L g1629 ( 
.A(n_1545),
.B(n_1561),
.Y(n_1629)
);

NAND2xp5_ASAP7_75t_L g1630 ( 
.A(n_1545),
.B(n_1521),
.Y(n_1630)
);

AOI22xp33_ASAP7_75t_L g1631 ( 
.A1(n_1565),
.A2(n_1508),
.B1(n_1399),
.B2(n_1364),
.Y(n_1631)
);

NAND2xp5_ASAP7_75t_L g1632 ( 
.A(n_1561),
.B(n_1473),
.Y(n_1632)
);

NAND3xp33_ASAP7_75t_L g1633 ( 
.A(n_1576),
.B(n_1483),
.C(n_1485),
.Y(n_1633)
);

OAI22xp5_ASAP7_75t_L g1634 ( 
.A1(n_1540),
.A2(n_1509),
.B1(n_1425),
.B2(n_1364),
.Y(n_1634)
);

OAI21xp5_ASAP7_75t_SL g1635 ( 
.A1(n_1555),
.A2(n_1513),
.B(n_1512),
.Y(n_1635)
);

OAI221xp5_ASAP7_75t_L g1636 ( 
.A1(n_1552),
.A2(n_1519),
.B1(n_1513),
.B2(n_1512),
.C(n_1409),
.Y(n_1636)
);

NAND2xp5_ASAP7_75t_L g1637 ( 
.A(n_1562),
.B(n_1473),
.Y(n_1637)
);

NAND2xp5_ASAP7_75t_L g1638 ( 
.A(n_1562),
.B(n_1571),
.Y(n_1638)
);

NAND2xp5_ASAP7_75t_L g1639 ( 
.A(n_1612),
.B(n_1568),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_1622),
.Y(n_1640)
);

INVxp33_ASAP7_75t_L g1641 ( 
.A(n_1600),
.Y(n_1641)
);

AND2x2_ASAP7_75t_L g1642 ( 
.A(n_1581),
.B(n_1586),
.Y(n_1642)
);

NOR2xp33_ASAP7_75t_L g1643 ( 
.A(n_1589),
.B(n_1484),
.Y(n_1643)
);

NAND3xp33_ASAP7_75t_L g1644 ( 
.A(n_1588),
.B(n_1518),
.C(n_1526),
.Y(n_1644)
);

NAND2x1_ASAP7_75t_SL g1645 ( 
.A(n_1611),
.B(n_1573),
.Y(n_1645)
);

BUFx2_ASAP7_75t_L g1646 ( 
.A(n_1613),
.Y(n_1646)
);

INVx1_ASAP7_75t_L g1647 ( 
.A(n_1622),
.Y(n_1647)
);

OR2x2_ASAP7_75t_L g1648 ( 
.A(n_1583),
.B(n_1554),
.Y(n_1648)
);

OR2x2_ASAP7_75t_L g1649 ( 
.A(n_1584),
.B(n_1554),
.Y(n_1649)
);

INVx2_ASAP7_75t_L g1650 ( 
.A(n_1590),
.Y(n_1650)
);

INVx2_ASAP7_75t_L g1651 ( 
.A(n_1590),
.Y(n_1651)
);

INVx2_ASAP7_75t_L g1652 ( 
.A(n_1595),
.Y(n_1652)
);

AND2x4_ASAP7_75t_L g1653 ( 
.A(n_1616),
.B(n_1564),
.Y(n_1653)
);

INVx1_ASAP7_75t_L g1654 ( 
.A(n_1626),
.Y(n_1654)
);

INVxp67_ASAP7_75t_L g1655 ( 
.A(n_1580),
.Y(n_1655)
);

AND2x4_ASAP7_75t_L g1656 ( 
.A(n_1623),
.B(n_1564),
.Y(n_1656)
);

AND2x2_ASAP7_75t_L g1657 ( 
.A(n_1595),
.B(n_1564),
.Y(n_1657)
);

AND2x2_ASAP7_75t_L g1658 ( 
.A(n_1620),
.B(n_1578),
.Y(n_1658)
);

INVx1_ASAP7_75t_L g1659 ( 
.A(n_1630),
.Y(n_1659)
);

AND2x4_ASAP7_75t_L g1660 ( 
.A(n_1623),
.B(n_1569),
.Y(n_1660)
);

INVx2_ASAP7_75t_L g1661 ( 
.A(n_1598),
.Y(n_1661)
);

NAND2xp5_ASAP7_75t_L g1662 ( 
.A(n_1591),
.B(n_1609),
.Y(n_1662)
);

OR2x2_ASAP7_75t_L g1663 ( 
.A(n_1593),
.B(n_1629),
.Y(n_1663)
);

INVx2_ASAP7_75t_L g1664 ( 
.A(n_1598),
.Y(n_1664)
);

HB1xp67_ASAP7_75t_L g1665 ( 
.A(n_1627),
.Y(n_1665)
);

INVx2_ASAP7_75t_L g1666 ( 
.A(n_1599),
.Y(n_1666)
);

OR2x6_ASAP7_75t_L g1667 ( 
.A(n_1597),
.B(n_1628),
.Y(n_1667)
);

AND2x4_ASAP7_75t_L g1668 ( 
.A(n_1594),
.B(n_1546),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_1625),
.Y(n_1669)
);

INVxp67_ASAP7_75t_L g1670 ( 
.A(n_1614),
.Y(n_1670)
);

INVx4_ASAP7_75t_L g1671 ( 
.A(n_1582),
.Y(n_1671)
);

BUFx2_ASAP7_75t_L g1672 ( 
.A(n_1613),
.Y(n_1672)
);

HB1xp67_ASAP7_75t_L g1673 ( 
.A(n_1633),
.Y(n_1673)
);

NAND2x1_ASAP7_75t_L g1674 ( 
.A(n_1610),
.B(n_1546),
.Y(n_1674)
);

OR2x2_ASAP7_75t_L g1675 ( 
.A(n_1618),
.B(n_1572),
.Y(n_1675)
);

BUFx6f_ASAP7_75t_L g1676 ( 
.A(n_1582),
.Y(n_1676)
);

INVxp67_ASAP7_75t_R g1677 ( 
.A(n_1585),
.Y(n_1677)
);

HB1xp67_ASAP7_75t_L g1678 ( 
.A(n_1596),
.Y(n_1678)
);

INVx2_ASAP7_75t_SL g1679 ( 
.A(n_1619),
.Y(n_1679)
);

INVx2_ASAP7_75t_L g1680 ( 
.A(n_1652),
.Y(n_1680)
);

INVx2_ASAP7_75t_L g1681 ( 
.A(n_1652),
.Y(n_1681)
);

INVx1_ASAP7_75t_L g1682 ( 
.A(n_1640),
.Y(n_1682)
);

AND2x2_ASAP7_75t_L g1683 ( 
.A(n_1657),
.B(n_1638),
.Y(n_1683)
);

INVx1_ASAP7_75t_L g1684 ( 
.A(n_1640),
.Y(n_1684)
);

OR2x2_ASAP7_75t_L g1685 ( 
.A(n_1655),
.B(n_1601),
.Y(n_1685)
);

NAND2xp5_ASAP7_75t_L g1686 ( 
.A(n_1678),
.B(n_1615),
.Y(n_1686)
);

AOI22xp5_ASAP7_75t_L g1687 ( 
.A1(n_1677),
.A2(n_1577),
.B1(n_1579),
.B2(n_1587),
.Y(n_1687)
);

NAND2xp5_ASAP7_75t_L g1688 ( 
.A(n_1678),
.B(n_1632),
.Y(n_1688)
);

NAND2xp5_ASAP7_75t_L g1689 ( 
.A(n_1655),
.B(n_1662),
.Y(n_1689)
);

AND2x2_ASAP7_75t_L g1690 ( 
.A(n_1657),
.B(n_1621),
.Y(n_1690)
);

NAND2xp5_ASAP7_75t_L g1691 ( 
.A(n_1662),
.B(n_1637),
.Y(n_1691)
);

AND2x2_ASAP7_75t_L g1692 ( 
.A(n_1646),
.B(n_1672),
.Y(n_1692)
);

AND2x2_ASAP7_75t_L g1693 ( 
.A(n_1646),
.B(n_1635),
.Y(n_1693)
);

AND2x2_ASAP7_75t_L g1694 ( 
.A(n_1672),
.B(n_1534),
.Y(n_1694)
);

NAND2xp5_ASAP7_75t_L g1695 ( 
.A(n_1669),
.B(n_1624),
.Y(n_1695)
);

NAND2xp5_ASAP7_75t_SL g1696 ( 
.A(n_1676),
.B(n_1604),
.Y(n_1696)
);

INVx1_ASAP7_75t_L g1697 ( 
.A(n_1647),
.Y(n_1697)
);

AND2x4_ASAP7_75t_SL g1698 ( 
.A(n_1676),
.B(n_1529),
.Y(n_1698)
);

INVx1_ASAP7_75t_L g1699 ( 
.A(n_1647),
.Y(n_1699)
);

NAND2xp5_ASAP7_75t_L g1700 ( 
.A(n_1669),
.B(n_1592),
.Y(n_1700)
);

INVx2_ASAP7_75t_L g1701 ( 
.A(n_1652),
.Y(n_1701)
);

INVx1_ASAP7_75t_L g1702 ( 
.A(n_1661),
.Y(n_1702)
);

INVx2_ASAP7_75t_L g1703 ( 
.A(n_1661),
.Y(n_1703)
);

INVx1_ASAP7_75t_L g1704 ( 
.A(n_1661),
.Y(n_1704)
);

NOR2x1p5_ASAP7_75t_L g1705 ( 
.A(n_1671),
.B(n_1453),
.Y(n_1705)
);

AND2x2_ASAP7_75t_L g1706 ( 
.A(n_1676),
.B(n_1534),
.Y(n_1706)
);

AND2x2_ASAP7_75t_L g1707 ( 
.A(n_1676),
.B(n_1534),
.Y(n_1707)
);

BUFx3_ASAP7_75t_L g1708 ( 
.A(n_1676),
.Y(n_1708)
);

OR2x2_ASAP7_75t_L g1709 ( 
.A(n_1673),
.B(n_1607),
.Y(n_1709)
);

INVx1_ASAP7_75t_L g1710 ( 
.A(n_1664),
.Y(n_1710)
);

NOR2xp33_ASAP7_75t_L g1711 ( 
.A(n_1643),
.B(n_1453),
.Y(n_1711)
);

AND2x4_ASAP7_75t_SL g1712 ( 
.A(n_1676),
.B(n_1529),
.Y(n_1712)
);

INVx1_ASAP7_75t_L g1713 ( 
.A(n_1664),
.Y(n_1713)
);

NOR2xp33_ASAP7_75t_L g1714 ( 
.A(n_1641),
.B(n_1663),
.Y(n_1714)
);

INVx3_ASAP7_75t_L g1715 ( 
.A(n_1674),
.Y(n_1715)
);

NAND2x1p5_ASAP7_75t_SL g1716 ( 
.A(n_1677),
.B(n_1448),
.Y(n_1716)
);

OR2x2_ASAP7_75t_L g1717 ( 
.A(n_1673),
.B(n_1568),
.Y(n_1717)
);

AND2x4_ASAP7_75t_L g1718 ( 
.A(n_1656),
.B(n_1572),
.Y(n_1718)
);

NAND2xp5_ASAP7_75t_SL g1719 ( 
.A(n_1671),
.B(n_1606),
.Y(n_1719)
);

INVx1_ASAP7_75t_L g1720 ( 
.A(n_1664),
.Y(n_1720)
);

NOR2x1_ASAP7_75t_SL g1721 ( 
.A(n_1667),
.B(n_1608),
.Y(n_1721)
);

INVx1_ASAP7_75t_L g1722 ( 
.A(n_1666),
.Y(n_1722)
);

AND2x2_ASAP7_75t_L g1723 ( 
.A(n_1671),
.B(n_1656),
.Y(n_1723)
);

INVx1_ASAP7_75t_L g1724 ( 
.A(n_1666),
.Y(n_1724)
);

INVx1_ASAP7_75t_L g1725 ( 
.A(n_1717),
.Y(n_1725)
);

INVxp67_ASAP7_75t_L g1726 ( 
.A(n_1700),
.Y(n_1726)
);

INVx1_ASAP7_75t_L g1727 ( 
.A(n_1717),
.Y(n_1727)
);

INVx2_ASAP7_75t_L g1728 ( 
.A(n_1680),
.Y(n_1728)
);

INVx2_ASAP7_75t_L g1729 ( 
.A(n_1680),
.Y(n_1729)
);

OR2x2_ASAP7_75t_L g1730 ( 
.A(n_1685),
.B(n_1663),
.Y(n_1730)
);

AND2x2_ASAP7_75t_L g1731 ( 
.A(n_1692),
.B(n_1667),
.Y(n_1731)
);

OR2x2_ASAP7_75t_L g1732 ( 
.A(n_1709),
.B(n_1665),
.Y(n_1732)
);

INVxp67_ASAP7_75t_L g1733 ( 
.A(n_1689),
.Y(n_1733)
);

NAND2xp5_ASAP7_75t_L g1734 ( 
.A(n_1714),
.B(n_1670),
.Y(n_1734)
);

A2O1A1Ixp33_ASAP7_75t_L g1735 ( 
.A1(n_1687),
.A2(n_1645),
.B(n_1644),
.C(n_1670),
.Y(n_1735)
);

OR2x2_ASAP7_75t_L g1736 ( 
.A(n_1709),
.B(n_1665),
.Y(n_1736)
);

NAND2xp33_ASAP7_75t_L g1737 ( 
.A(n_1687),
.B(n_1644),
.Y(n_1737)
);

OR2x2_ASAP7_75t_L g1738 ( 
.A(n_1685),
.B(n_1675),
.Y(n_1738)
);

AND2x2_ASAP7_75t_L g1739 ( 
.A(n_1692),
.B(n_1723),
.Y(n_1739)
);

INVx2_ASAP7_75t_L g1740 ( 
.A(n_1681),
.Y(n_1740)
);

OR2x2_ASAP7_75t_L g1741 ( 
.A(n_1686),
.B(n_1675),
.Y(n_1741)
);

INVx2_ASAP7_75t_L g1742 ( 
.A(n_1681),
.Y(n_1742)
);

INVx1_ASAP7_75t_L g1743 ( 
.A(n_1682),
.Y(n_1743)
);

INVx1_ASAP7_75t_L g1744 ( 
.A(n_1682),
.Y(n_1744)
);

AND2x2_ASAP7_75t_L g1745 ( 
.A(n_1723),
.B(n_1667),
.Y(n_1745)
);

OR2x2_ASAP7_75t_L g1746 ( 
.A(n_1691),
.B(n_1649),
.Y(n_1746)
);

NAND2xp5_ASAP7_75t_L g1747 ( 
.A(n_1690),
.B(n_1679),
.Y(n_1747)
);

NAND2x2_ASAP7_75t_L g1748 ( 
.A(n_1705),
.B(n_1431),
.Y(n_1748)
);

NAND2xp5_ASAP7_75t_L g1749 ( 
.A(n_1690),
.B(n_1679),
.Y(n_1749)
);

INVx1_ASAP7_75t_L g1750 ( 
.A(n_1684),
.Y(n_1750)
);

INVx1_ASAP7_75t_L g1751 ( 
.A(n_1684),
.Y(n_1751)
);

NAND2xp5_ASAP7_75t_L g1752 ( 
.A(n_1683),
.B(n_1679),
.Y(n_1752)
);

INVx1_ASAP7_75t_SL g1753 ( 
.A(n_1696),
.Y(n_1753)
);

OR2x2_ASAP7_75t_L g1754 ( 
.A(n_1688),
.B(n_1649),
.Y(n_1754)
);

AND2x2_ASAP7_75t_L g1755 ( 
.A(n_1708),
.B(n_1667),
.Y(n_1755)
);

NAND2xp5_ASAP7_75t_L g1756 ( 
.A(n_1683),
.B(n_1695),
.Y(n_1756)
);

INVx1_ASAP7_75t_L g1757 ( 
.A(n_1697),
.Y(n_1757)
);

AND2x2_ASAP7_75t_L g1758 ( 
.A(n_1708),
.B(n_1667),
.Y(n_1758)
);

INVxp67_ASAP7_75t_L g1759 ( 
.A(n_1694),
.Y(n_1759)
);

NAND2xp5_ASAP7_75t_L g1760 ( 
.A(n_1694),
.B(n_1654),
.Y(n_1760)
);

AND2x4_ASAP7_75t_L g1761 ( 
.A(n_1705),
.B(n_1671),
.Y(n_1761)
);

AND2x2_ASAP7_75t_SL g1762 ( 
.A(n_1698),
.B(n_1555),
.Y(n_1762)
);

AND2x2_ASAP7_75t_L g1763 ( 
.A(n_1708),
.B(n_1653),
.Y(n_1763)
);

INVx1_ASAP7_75t_L g1764 ( 
.A(n_1697),
.Y(n_1764)
);

NAND2xp5_ASAP7_75t_L g1765 ( 
.A(n_1706),
.B(n_1654),
.Y(n_1765)
);

INVx1_ASAP7_75t_L g1766 ( 
.A(n_1699),
.Y(n_1766)
);

INVx1_ASAP7_75t_L g1767 ( 
.A(n_1699),
.Y(n_1767)
);

AND2x2_ASAP7_75t_L g1768 ( 
.A(n_1693),
.B(n_1653),
.Y(n_1768)
);

AOI22xp5_ASAP7_75t_L g1769 ( 
.A1(n_1719),
.A2(n_1653),
.B1(n_1660),
.B2(n_1656),
.Y(n_1769)
);

AND2x2_ASAP7_75t_L g1770 ( 
.A(n_1693),
.B(n_1653),
.Y(n_1770)
);

BUFx2_ASAP7_75t_L g1771 ( 
.A(n_1739),
.Y(n_1771)
);

NAND2xp5_ASAP7_75t_L g1772 ( 
.A(n_1726),
.B(n_1706),
.Y(n_1772)
);

INVx1_ASAP7_75t_L g1773 ( 
.A(n_1743),
.Y(n_1773)
);

INVx1_ASAP7_75t_SL g1774 ( 
.A(n_1753),
.Y(n_1774)
);

AOI22xp33_ASAP7_75t_L g1775 ( 
.A1(n_1737),
.A2(n_1707),
.B1(n_1712),
.B2(n_1698),
.Y(n_1775)
);

INVx1_ASAP7_75t_SL g1776 ( 
.A(n_1732),
.Y(n_1776)
);

INVxp67_ASAP7_75t_L g1777 ( 
.A(n_1732),
.Y(n_1777)
);

NOR2x1_ASAP7_75t_L g1778 ( 
.A(n_1737),
.B(n_1711),
.Y(n_1778)
);

NAND2xp5_ASAP7_75t_L g1779 ( 
.A(n_1733),
.B(n_1707),
.Y(n_1779)
);

NOR2xp33_ASAP7_75t_L g1780 ( 
.A(n_1734),
.B(n_1472),
.Y(n_1780)
);

AND2x2_ASAP7_75t_L g1781 ( 
.A(n_1739),
.B(n_1721),
.Y(n_1781)
);

INVx3_ASAP7_75t_SL g1782 ( 
.A(n_1761),
.Y(n_1782)
);

NAND2xp5_ASAP7_75t_L g1783 ( 
.A(n_1759),
.B(n_1658),
.Y(n_1783)
);

INVx1_ASAP7_75t_SL g1784 ( 
.A(n_1736),
.Y(n_1784)
);

INVxp67_ASAP7_75t_L g1785 ( 
.A(n_1736),
.Y(n_1785)
);

NAND2xp5_ASAP7_75t_L g1786 ( 
.A(n_1735),
.B(n_1725),
.Y(n_1786)
);

OR2x2_ASAP7_75t_L g1787 ( 
.A(n_1730),
.B(n_1716),
.Y(n_1787)
);

NAND2xp33_ASAP7_75t_L g1788 ( 
.A(n_1735),
.B(n_1716),
.Y(n_1788)
);

NAND2xp5_ASAP7_75t_L g1789 ( 
.A(n_1727),
.B(n_1658),
.Y(n_1789)
);

INVx2_ASAP7_75t_SL g1790 ( 
.A(n_1763),
.Y(n_1790)
);

NAND2xp5_ASAP7_75t_L g1791 ( 
.A(n_1756),
.B(n_1659),
.Y(n_1791)
);

INVx1_ASAP7_75t_L g1792 ( 
.A(n_1744),
.Y(n_1792)
);

HB1xp67_ASAP7_75t_L g1793 ( 
.A(n_1738),
.Y(n_1793)
);

NOR2x1_ASAP7_75t_L g1794 ( 
.A(n_1755),
.B(n_1715),
.Y(n_1794)
);

HB1xp67_ASAP7_75t_L g1795 ( 
.A(n_1738),
.Y(n_1795)
);

INVx1_ASAP7_75t_SL g1796 ( 
.A(n_1761),
.Y(n_1796)
);

AND2x2_ASAP7_75t_L g1797 ( 
.A(n_1768),
.B(n_1721),
.Y(n_1797)
);

NAND4xp25_ASAP7_75t_L g1798 ( 
.A(n_1755),
.B(n_1602),
.C(n_1631),
.D(n_1605),
.Y(n_1798)
);

NAND2xp5_ASAP7_75t_L g1799 ( 
.A(n_1765),
.B(n_1659),
.Y(n_1799)
);

HB1xp67_ASAP7_75t_L g1800 ( 
.A(n_1750),
.Y(n_1800)
);

OR2x2_ASAP7_75t_L g1801 ( 
.A(n_1741),
.B(n_1716),
.Y(n_1801)
);

AND2x4_ASAP7_75t_SL g1802 ( 
.A(n_1761),
.B(n_1715),
.Y(n_1802)
);

NAND2xp5_ASAP7_75t_L g1803 ( 
.A(n_1760),
.B(n_1642),
.Y(n_1803)
);

CKINVDCx16_ASAP7_75t_R g1804 ( 
.A(n_1758),
.Y(n_1804)
);

INVx3_ASAP7_75t_L g1805 ( 
.A(n_1762),
.Y(n_1805)
);

BUFx3_ASAP7_75t_L g1806 ( 
.A(n_1758),
.Y(n_1806)
);

NOR2x1_ASAP7_75t_L g1807 ( 
.A(n_1731),
.B(n_1715),
.Y(n_1807)
);

INVx1_ASAP7_75t_SL g1808 ( 
.A(n_1731),
.Y(n_1808)
);

INVx2_ASAP7_75t_L g1809 ( 
.A(n_1771),
.Y(n_1809)
);

OR2x2_ASAP7_75t_L g1810 ( 
.A(n_1776),
.B(n_1741),
.Y(n_1810)
);

OAI21xp5_ASAP7_75t_SL g1811 ( 
.A1(n_1778),
.A2(n_1745),
.B(n_1769),
.Y(n_1811)
);

OAI22xp33_ASAP7_75t_L g1812 ( 
.A1(n_1786),
.A2(n_1748),
.B1(n_1752),
.B2(n_1749),
.Y(n_1812)
);

INVx2_ASAP7_75t_L g1813 ( 
.A(n_1771),
.Y(n_1813)
);

INVx1_ASAP7_75t_L g1814 ( 
.A(n_1793),
.Y(n_1814)
);

NOR2x1_ASAP7_75t_L g1815 ( 
.A(n_1788),
.B(n_1763),
.Y(n_1815)
);

INVx1_ASAP7_75t_L g1816 ( 
.A(n_1795),
.Y(n_1816)
);

NAND2xp5_ASAP7_75t_L g1817 ( 
.A(n_1774),
.B(n_1746),
.Y(n_1817)
);

NAND2xp5_ASAP7_75t_L g1818 ( 
.A(n_1784),
.B(n_1768),
.Y(n_1818)
);

OAI21xp5_ASAP7_75t_L g1819 ( 
.A1(n_1788),
.A2(n_1745),
.B(n_1645),
.Y(n_1819)
);

OAI221xp5_ASAP7_75t_L g1820 ( 
.A1(n_1775),
.A2(n_1748),
.B1(n_1770),
.B2(n_1754),
.C(n_1747),
.Y(n_1820)
);

NOR2xp67_ASAP7_75t_L g1821 ( 
.A(n_1805),
.B(n_1770),
.Y(n_1821)
);

AND2x2_ASAP7_75t_L g1822 ( 
.A(n_1804),
.B(n_1782),
.Y(n_1822)
);

INVxp67_ASAP7_75t_L g1823 ( 
.A(n_1806),
.Y(n_1823)
);

A2O1A1Ixp33_ASAP7_75t_L g1824 ( 
.A1(n_1777),
.A2(n_1712),
.B(n_1668),
.C(n_1762),
.Y(n_1824)
);

INVx1_ASAP7_75t_L g1825 ( 
.A(n_1800),
.Y(n_1825)
);

NOR2xp33_ASAP7_75t_L g1826 ( 
.A(n_1804),
.B(n_1396),
.Y(n_1826)
);

OAI21xp5_ASAP7_75t_L g1827 ( 
.A1(n_1807),
.A2(n_1757),
.B(n_1751),
.Y(n_1827)
);

INVx1_ASAP7_75t_L g1828 ( 
.A(n_1773),
.Y(n_1828)
);

AOI221xp5_ASAP7_75t_L g1829 ( 
.A1(n_1785),
.A2(n_1767),
.B1(n_1766),
.B2(n_1764),
.C(n_1742),
.Y(n_1829)
);

OAI22xp5_ASAP7_75t_L g1830 ( 
.A1(n_1782),
.A2(n_1656),
.B1(n_1660),
.B2(n_1631),
.Y(n_1830)
);

INVx1_ASAP7_75t_L g1831 ( 
.A(n_1773),
.Y(n_1831)
);

NAND2xp5_ASAP7_75t_L g1832 ( 
.A(n_1808),
.B(n_1742),
.Y(n_1832)
);

NOR3xp33_ASAP7_75t_L g1833 ( 
.A(n_1772),
.B(n_1413),
.C(n_1431),
.Y(n_1833)
);

INVx1_ASAP7_75t_L g1834 ( 
.A(n_1792),
.Y(n_1834)
);

INVx1_ASAP7_75t_L g1835 ( 
.A(n_1792),
.Y(n_1835)
);

INVx2_ASAP7_75t_L g1836 ( 
.A(n_1806),
.Y(n_1836)
);

NAND2xp5_ASAP7_75t_L g1837 ( 
.A(n_1823),
.B(n_1796),
.Y(n_1837)
);

NOR2xp33_ASAP7_75t_L g1838 ( 
.A(n_1826),
.B(n_1780),
.Y(n_1838)
);

NAND2xp5_ASAP7_75t_L g1839 ( 
.A(n_1836),
.B(n_1790),
.Y(n_1839)
);

INVx1_ASAP7_75t_L g1840 ( 
.A(n_1809),
.Y(n_1840)
);

INVx1_ASAP7_75t_L g1841 ( 
.A(n_1809),
.Y(n_1841)
);

NOR2xp33_ASAP7_75t_L g1842 ( 
.A(n_1826),
.B(n_1779),
.Y(n_1842)
);

NAND2xp5_ASAP7_75t_L g1843 ( 
.A(n_1813),
.B(n_1790),
.Y(n_1843)
);

AOI22xp5_ASAP7_75t_L g1844 ( 
.A1(n_1815),
.A2(n_1805),
.B1(n_1781),
.B2(n_1797),
.Y(n_1844)
);

AND2x2_ASAP7_75t_L g1845 ( 
.A(n_1822),
.B(n_1797),
.Y(n_1845)
);

NOR2xp33_ASAP7_75t_L g1846 ( 
.A(n_1814),
.B(n_1805),
.Y(n_1846)
);

INVx1_ASAP7_75t_L g1847 ( 
.A(n_1813),
.Y(n_1847)
);

INVx1_ASAP7_75t_L g1848 ( 
.A(n_1828),
.Y(n_1848)
);

NAND2xp5_ASAP7_75t_L g1849 ( 
.A(n_1816),
.B(n_1783),
.Y(n_1849)
);

NAND2xp5_ASAP7_75t_L g1850 ( 
.A(n_1825),
.B(n_1789),
.Y(n_1850)
);

NAND2xp5_ASAP7_75t_L g1851 ( 
.A(n_1817),
.B(n_1781),
.Y(n_1851)
);

AND2x2_ASAP7_75t_L g1852 ( 
.A(n_1821),
.B(n_1802),
.Y(n_1852)
);

INVx1_ASAP7_75t_L g1853 ( 
.A(n_1831),
.Y(n_1853)
);

AOI22xp33_ASAP7_75t_L g1854 ( 
.A1(n_1833),
.A2(n_1798),
.B1(n_1801),
.B2(n_1787),
.Y(n_1854)
);

NAND2xp5_ASAP7_75t_L g1855 ( 
.A(n_1818),
.B(n_1803),
.Y(n_1855)
);

INVx1_ASAP7_75t_L g1856 ( 
.A(n_1834),
.Y(n_1856)
);

INVx1_ASAP7_75t_L g1857 ( 
.A(n_1835),
.Y(n_1857)
);

OAI21xp33_ASAP7_75t_SL g1858 ( 
.A1(n_1844),
.A2(n_1827),
.B(n_1819),
.Y(n_1858)
);

AOI22xp5_ASAP7_75t_L g1859 ( 
.A1(n_1845),
.A2(n_1833),
.B1(n_1811),
.B2(n_1812),
.Y(n_1859)
);

NAND2xp5_ASAP7_75t_L g1860 ( 
.A(n_1846),
.B(n_1810),
.Y(n_1860)
);

O2A1O1Ixp33_ASAP7_75t_L g1861 ( 
.A1(n_1854),
.A2(n_1812),
.B(n_1824),
.C(n_1801),
.Y(n_1861)
);

AOI211x1_ASAP7_75t_SL g1862 ( 
.A1(n_1843),
.A2(n_1832),
.B(n_1824),
.C(n_1830),
.Y(n_1862)
);

OA21x2_ASAP7_75t_SL g1863 ( 
.A1(n_1837),
.A2(n_1799),
.B(n_1791),
.Y(n_1863)
);

OAI21xp33_ASAP7_75t_L g1864 ( 
.A1(n_1854),
.A2(n_1820),
.B(n_1829),
.Y(n_1864)
);

INVx1_ASAP7_75t_L g1865 ( 
.A(n_1840),
.Y(n_1865)
);

AOI211x1_ASAP7_75t_L g1866 ( 
.A1(n_1851),
.A2(n_1794),
.B(n_1636),
.C(n_1802),
.Y(n_1866)
);

HB1xp67_ASAP7_75t_L g1867 ( 
.A(n_1841),
.Y(n_1867)
);

OAI21xp5_ASAP7_75t_L g1868 ( 
.A1(n_1838),
.A2(n_1787),
.B(n_1729),
.Y(n_1868)
);

NAND2xp5_ASAP7_75t_L g1869 ( 
.A(n_1846),
.B(n_1728),
.Y(n_1869)
);

AOI222xp33_ASAP7_75t_L g1870 ( 
.A1(n_1842),
.A2(n_1668),
.B1(n_1740),
.B2(n_1729),
.C1(n_1728),
.C2(n_1651),
.Y(n_1870)
);

NAND4xp25_ASAP7_75t_L g1871 ( 
.A(n_1849),
.B(n_1740),
.C(n_1603),
.D(n_1634),
.Y(n_1871)
);

NAND2xp5_ASAP7_75t_L g1872 ( 
.A(n_1862),
.B(n_1847),
.Y(n_1872)
);

NAND3xp33_ASAP7_75t_L g1873 ( 
.A(n_1861),
.B(n_1839),
.C(n_1848),
.Y(n_1873)
);

HB1xp67_ASAP7_75t_L g1874 ( 
.A(n_1867),
.Y(n_1874)
);

NOR2x1_ASAP7_75t_L g1875 ( 
.A(n_1860),
.B(n_1853),
.Y(n_1875)
);

NAND2xp5_ASAP7_75t_L g1876 ( 
.A(n_1864),
.B(n_1838),
.Y(n_1876)
);

AND5x1_ASAP7_75t_L g1877 ( 
.A(n_1859),
.B(n_1863),
.C(n_1858),
.D(n_1866),
.E(n_1870),
.Y(n_1877)
);

NAND3xp33_ASAP7_75t_L g1878 ( 
.A(n_1868),
.B(n_1857),
.C(n_1856),
.Y(n_1878)
);

NAND3xp33_ASAP7_75t_SL g1879 ( 
.A(n_1869),
.B(n_1852),
.C(n_1850),
.Y(n_1879)
);

NOR2xp33_ASAP7_75t_L g1880 ( 
.A(n_1865),
.B(n_1855),
.Y(n_1880)
);

NOR2x1_ASAP7_75t_L g1881 ( 
.A(n_1871),
.B(n_1370),
.Y(n_1881)
);

NAND2xp5_ASAP7_75t_L g1882 ( 
.A(n_1867),
.B(n_1703),
.Y(n_1882)
);

NAND3xp33_ASAP7_75t_L g1883 ( 
.A(n_1861),
.B(n_1413),
.C(n_1428),
.Y(n_1883)
);

NOR2x1_ASAP7_75t_L g1884 ( 
.A(n_1860),
.B(n_1715),
.Y(n_1884)
);

NOR2xp33_ASAP7_75t_L g1885 ( 
.A(n_1876),
.B(n_1398),
.Y(n_1885)
);

NOR3xp33_ASAP7_75t_SL g1886 ( 
.A(n_1873),
.B(n_1639),
.C(n_1702),
.Y(n_1886)
);

OAI211xp5_ASAP7_75t_SL g1887 ( 
.A1(n_1883),
.A2(n_1648),
.B(n_1722),
.C(n_1720),
.Y(n_1887)
);

NOR2xp33_ASAP7_75t_L g1888 ( 
.A(n_1879),
.B(n_1703),
.Y(n_1888)
);

NAND2xp5_ASAP7_75t_L g1889 ( 
.A(n_1875),
.B(n_1702),
.Y(n_1889)
);

NAND3xp33_ASAP7_75t_SL g1890 ( 
.A(n_1872),
.B(n_1674),
.C(n_1617),
.Y(n_1890)
);

NAND2xp5_ASAP7_75t_L g1891 ( 
.A(n_1888),
.B(n_1874),
.Y(n_1891)
);

INVxp67_ASAP7_75t_SL g1892 ( 
.A(n_1885),
.Y(n_1892)
);

INVx1_ASAP7_75t_L g1893 ( 
.A(n_1889),
.Y(n_1893)
);

NAND2xp5_ASAP7_75t_L g1894 ( 
.A(n_1886),
.B(n_1880),
.Y(n_1894)
);

HB1xp67_ASAP7_75t_L g1895 ( 
.A(n_1890),
.Y(n_1895)
);

OAI22xp5_ASAP7_75t_L g1896 ( 
.A1(n_1887),
.A2(n_1878),
.B1(n_1881),
.B2(n_1884),
.Y(n_1896)
);

NOR2x1_ASAP7_75t_L g1897 ( 
.A(n_1885),
.B(n_1882),
.Y(n_1897)
);

OAI211xp5_ASAP7_75t_SL g1898 ( 
.A1(n_1897),
.A2(n_1877),
.B(n_1648),
.C(n_1722),
.Y(n_1898)
);

NAND2xp5_ASAP7_75t_L g1899 ( 
.A(n_1895),
.B(n_1704),
.Y(n_1899)
);

INVx1_ASAP7_75t_SL g1900 ( 
.A(n_1891),
.Y(n_1900)
);

INVx1_ASAP7_75t_SL g1901 ( 
.A(n_1894),
.Y(n_1901)
);

INVx1_ASAP7_75t_L g1902 ( 
.A(n_1893),
.Y(n_1902)
);

NAND2xp5_ASAP7_75t_L g1903 ( 
.A(n_1892),
.B(n_1704),
.Y(n_1903)
);

OAI21xp5_ASAP7_75t_L g1904 ( 
.A1(n_1898),
.A2(n_1896),
.B(n_1713),
.Y(n_1904)
);

XOR2x1_ASAP7_75t_L g1905 ( 
.A(n_1902),
.B(n_1900),
.Y(n_1905)
);

XOR2xp5_ASAP7_75t_L g1906 ( 
.A(n_1901),
.B(n_1422),
.Y(n_1906)
);

AND2x2_ASAP7_75t_L g1907 ( 
.A(n_1899),
.B(n_1642),
.Y(n_1907)
);

INVx1_ASAP7_75t_L g1908 ( 
.A(n_1905),
.Y(n_1908)
);

AOI22xp5_ASAP7_75t_L g1909 ( 
.A1(n_1906),
.A2(n_1903),
.B1(n_1718),
.B2(n_1668),
.Y(n_1909)
);

AND4x2_ASAP7_75t_L g1910 ( 
.A(n_1908),
.B(n_1904),
.C(n_1907),
.D(n_1428),
.Y(n_1910)
);

INVx1_ASAP7_75t_L g1911 ( 
.A(n_1910),
.Y(n_1911)
);

INVx1_ASAP7_75t_L g1912 ( 
.A(n_1910),
.Y(n_1912)
);

AO21x2_ASAP7_75t_L g1913 ( 
.A1(n_1911),
.A2(n_1909),
.B(n_1650),
.Y(n_1913)
);

NAND2xp5_ASAP7_75t_L g1914 ( 
.A(n_1912),
.B(n_1701),
.Y(n_1914)
);

NAND2xp5_ASAP7_75t_L g1915 ( 
.A(n_1913),
.B(n_1701),
.Y(n_1915)
);

AOI21xp5_ASAP7_75t_SL g1916 ( 
.A1(n_1915),
.A2(n_1914),
.B(n_1423),
.Y(n_1916)
);

AOI22xp33_ASAP7_75t_L g1917 ( 
.A1(n_1916),
.A2(n_1428),
.B1(n_1651),
.B2(n_1650),
.Y(n_1917)
);

OAI221xp5_ASAP7_75t_R g1918 ( 
.A1(n_1917),
.A2(n_1724),
.B1(n_1720),
.B2(n_1710),
.C(n_1713),
.Y(n_1918)
);

AOI211xp5_ASAP7_75t_L g1919 ( 
.A1(n_1918),
.A2(n_1423),
.B(n_1400),
.C(n_1384),
.Y(n_1919)
);


endmodule