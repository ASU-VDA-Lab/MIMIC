module fake_jpeg_17513_n_283 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_283);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_283;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_127;
wire n_76;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_272;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_258;
wire n_282;
wire n_96;

INVx1_ASAP7_75t_L g13 ( 
.A(n_10),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_11),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_11),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

BUFx12_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_4),
.Y(n_23)
);

BUFx8_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

INVx2_ASAP7_75t_SL g26 ( 
.A(n_5),
.Y(n_26)
);

INVx11_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_20),
.Y(n_28)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_28),
.Y(n_45)
);

INVx2_ASAP7_75t_SL g29 ( 
.A(n_17),
.Y(n_29)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_29),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_25),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_30),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_25),
.Y(n_31)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_31),
.Y(n_43)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_17),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_32),
.B(n_34),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_25),
.Y(n_33)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_33),
.Y(n_46)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_17),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_20),
.Y(n_35)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_25),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_37),
.Y(n_38)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_37),
.Y(n_39)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_39),
.Y(n_67)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_32),
.Y(n_40)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

CKINVDCx14_ASAP7_75t_R g41 ( 
.A(n_34),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_41),
.B(n_21),
.Y(n_57)
);

AND2x2_ASAP7_75t_L g42 ( 
.A(n_28),
.B(n_16),
.Y(n_42)
);

INVx1_ASAP7_75t_SL g53 ( 
.A(n_42),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_35),
.B(n_20),
.Y(n_44)
);

AND2x2_ASAP7_75t_SL g60 ( 
.A(n_44),
.B(n_16),
.Y(n_60)
);

INVx2_ASAP7_75t_SL g49 ( 
.A(n_29),
.Y(n_49)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_49),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_45),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_54),
.B(n_64),
.Y(n_80)
);

XNOR2xp5_ASAP7_75t_L g56 ( 
.A(n_44),
.B(n_24),
.Y(n_56)
);

XOR2xp5_ASAP7_75t_L g95 ( 
.A(n_56),
.B(n_24),
.Y(n_95)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_57),
.Y(n_90)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_51),
.Y(n_58)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_58),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_40),
.A2(n_26),
.B1(n_27),
.B2(n_18),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_59),
.A2(n_70),
.B1(n_26),
.B2(n_27),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_60),
.B(n_71),
.Y(n_83)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_51),
.Y(n_61)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_61),
.Y(n_85)
);

HB1xp67_ASAP7_75t_L g62 ( 
.A(n_45),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_62),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_52),
.B(n_18),
.Y(n_64)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_47),
.Y(n_65)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_65),
.Y(n_76)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_47),
.Y(n_66)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_66),
.Y(n_79)
);

BUFx2_ASAP7_75t_L g68 ( 
.A(n_47),
.Y(n_68)
);

INVxp67_ASAP7_75t_L g75 ( 
.A(n_68),
.Y(n_75)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_47),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_69),
.Y(n_77)
);

OAI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_42),
.A2(n_27),
.B1(n_23),
.B2(n_31),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_43),
.Y(n_71)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_49),
.Y(n_72)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_72),
.Y(n_94)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_49),
.Y(n_73)
);

BUFx3_ASAP7_75t_L g91 ( 
.A(n_73),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_53),
.A2(n_42),
.B1(n_18),
.B2(n_26),
.Y(n_74)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_74),
.Y(n_101)
);

AOI21xp33_ASAP7_75t_SL g78 ( 
.A1(n_53),
.A2(n_50),
.B(n_52),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_78),
.B(n_87),
.C(n_24),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_82),
.A2(n_88),
.B1(n_89),
.B2(n_92),
.Y(n_99)
);

AOI21xp5_ASAP7_75t_L g84 ( 
.A1(n_60),
.A2(n_17),
.B(n_43),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_84),
.Y(n_111)
);

FAx1_ASAP7_75t_SL g86 ( 
.A(n_56),
.B(n_60),
.CI(n_63),
.CON(n_86),
.SN(n_86)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_86),
.B(n_24),
.Y(n_107)
);

XNOR2xp5_ASAP7_75t_L g87 ( 
.A(n_61),
.B(n_29),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_67),
.A2(n_46),
.B1(n_39),
.B2(n_33),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_58),
.A2(n_46),
.B1(n_31),
.B2(n_33),
.Y(n_89)
);

OAI22xp33_ASAP7_75t_L g92 ( 
.A1(n_67),
.A2(n_48),
.B1(n_36),
.B2(n_30),
.Y(n_92)
);

XNOR2xp5_ASAP7_75t_L g100 ( 
.A(n_95),
.B(n_24),
.Y(n_100)
);

XOR2xp5_ASAP7_75t_SL g136 ( 
.A(n_96),
.B(n_21),
.Y(n_136)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_94),
.Y(n_97)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_97),
.Y(n_119)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_94),
.Y(n_98)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_98),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_100),
.B(n_102),
.C(n_17),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_95),
.B(n_69),
.C(n_17),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_85),
.Y(n_103)
);

HB1xp67_ASAP7_75t_L g121 ( 
.A(n_103),
.Y(n_121)
);

CKINVDCx16_ASAP7_75t_R g104 ( 
.A(n_80),
.Y(n_104)
);

HB1xp67_ASAP7_75t_L g139 ( 
.A(n_104),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_93),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_105),
.B(n_114),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_86),
.B(n_83),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_106),
.B(n_110),
.Y(n_117)
);

OAI21xp33_ASAP7_75t_L g118 ( 
.A1(n_107),
.A2(n_112),
.B(n_113),
.Y(n_118)
);

AND2x2_ASAP7_75t_SL g108 ( 
.A(n_84),
.B(n_73),
.Y(n_108)
);

INVx1_ASAP7_75t_SL g131 ( 
.A(n_108),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_86),
.A2(n_72),
.B1(n_55),
.B2(n_26),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_109),
.A2(n_101),
.B1(n_107),
.B2(n_112),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_87),
.B(n_48),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_74),
.B(n_19),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_90),
.B(n_19),
.Y(n_113)
);

CKINVDCx14_ASAP7_75t_R g114 ( 
.A(n_88),
.Y(n_114)
);

BUFx3_ASAP7_75t_L g115 ( 
.A(n_77),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_115),
.B(n_103),
.Y(n_137)
);

OA21x2_ASAP7_75t_L g116 ( 
.A1(n_92),
.A2(n_55),
.B(n_38),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_116),
.A2(n_85),
.B1(n_75),
.B2(n_81),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_97),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_120),
.B(n_132),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_123),
.A2(n_127),
.B1(n_129),
.B2(n_130),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_SL g153 ( 
.A(n_124),
.B(n_126),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_100),
.B(n_91),
.C(n_89),
.Y(n_125)
);

XOR2xp5_ASAP7_75t_L g146 ( 
.A(n_125),
.B(n_102),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_111),
.A2(n_75),
.B1(n_76),
.B2(n_79),
.Y(n_127)
);

AOI21xp5_ASAP7_75t_L g128 ( 
.A1(n_108),
.A2(n_0),
.B(n_1),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_SL g154 ( 
.A1(n_128),
.A2(n_113),
.B(n_104),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_108),
.A2(n_79),
.B1(n_76),
.B2(n_13),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_114),
.A2(n_13),
.B1(n_23),
.B2(n_77),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_98),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_99),
.A2(n_48),
.B1(n_38),
.B2(n_13),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_134),
.A2(n_140),
.B1(n_116),
.B2(n_109),
.Y(n_147)
);

BUFx2_ASAP7_75t_L g135 ( 
.A(n_115),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_135),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_SL g165 ( 
.A1(n_136),
.A2(n_21),
.B(n_22),
.Y(n_165)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_137),
.Y(n_142)
);

OAI22x1_ASAP7_75t_SL g138 ( 
.A1(n_108),
.A2(n_15),
.B1(n_14),
.B2(n_68),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_138),
.A2(n_116),
.B1(n_105),
.B2(n_110),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_99),
.A2(n_15),
.B1(n_14),
.B2(n_91),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g141 ( 
.A(n_127),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_141),
.B(n_145),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_SL g187 ( 
.A1(n_143),
.A2(n_154),
.B(n_160),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_119),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_146),
.B(n_153),
.C(n_164),
.Y(n_172)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_147),
.Y(n_189)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_119),
.Y(n_148)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_148),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_L g149 ( 
.A1(n_128),
.A2(n_96),
.B(n_106),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_L g181 ( 
.A1(n_149),
.A2(n_163),
.B(n_7),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_L g151 ( 
.A1(n_138),
.A2(n_133),
.B1(n_131),
.B2(n_116),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_151),
.A2(n_22),
.B1(n_1),
.B2(n_3),
.Y(n_183)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_122),
.Y(n_152)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_152),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_117),
.B(n_15),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_155),
.B(n_157),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_122),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_SL g185 ( 
.A(n_156),
.B(n_22),
.Y(n_185)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_129),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_123),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_158),
.B(n_159),
.Y(n_173)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_135),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_SL g160 ( 
.A1(n_131),
.A2(n_115),
.B(n_22),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_117),
.B(n_14),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_162),
.B(n_164),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_SL g163 ( 
.A1(n_136),
.A2(n_126),
.B(n_125),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_124),
.B(n_15),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_165),
.B(n_134),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_144),
.B(n_139),
.Y(n_166)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_166),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_150),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_169),
.B(n_171),
.Y(n_199)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_161),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_170),
.B(n_180),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_148),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_172),
.B(n_162),
.C(n_155),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_174),
.B(n_146),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_158),
.A2(n_140),
.B1(n_118),
.B2(n_121),
.Y(n_175)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_175),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_152),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_176),
.B(n_177),
.Y(n_204)
);

HB1xp67_ASAP7_75t_L g177 ( 
.A(n_142),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_141),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_180)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_181),
.B(n_165),
.Y(n_196)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_183),
.Y(n_193)
);

AOI21xp5_ASAP7_75t_L g184 ( 
.A1(n_160),
.A2(n_0),
.B(n_3),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_SL g202 ( 
.A1(n_184),
.A2(n_188),
.B(n_154),
.Y(n_202)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_185),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_157),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_186)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_186),
.Y(n_197)
);

XNOR2x1_ASAP7_75t_SL g188 ( 
.A(n_153),
.B(n_22),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_SL g210 ( 
.A(n_190),
.B(n_202),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_168),
.Y(n_192)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_192),
.Y(n_226)
);

OR2x2_ASAP7_75t_L g194 ( 
.A(n_173),
.B(n_143),
.Y(n_194)
);

OR2x2_ASAP7_75t_L g218 ( 
.A(n_194),
.B(n_178),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_196),
.B(n_201),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_168),
.Y(n_200)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_200),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_172),
.B(n_188),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_SL g203 ( 
.A1(n_173),
.A2(n_163),
.B(n_142),
.Y(n_203)
);

INVxp67_ASAP7_75t_L g213 ( 
.A(n_203),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_187),
.B(n_149),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_205),
.B(n_206),
.C(n_209),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_187),
.B(n_181),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_179),
.Y(n_207)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_207),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_198),
.A2(n_170),
.B1(n_189),
.B2(n_179),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_212),
.A2(n_224),
.B1(n_225),
.B2(n_197),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_199),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_214),
.B(n_215),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_204),
.Y(n_215)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_191),
.Y(n_217)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_217),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_L g228 ( 
.A1(n_218),
.A2(n_167),
.B(n_184),
.Y(n_228)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_203),
.Y(n_219)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_219),
.Y(n_234)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_195),
.Y(n_221)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_221),
.Y(n_235)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_208),
.Y(n_223)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_223),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_208),
.A2(n_189),
.B1(n_193),
.B2(n_198),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_194),
.A2(n_167),
.B1(n_182),
.B2(n_174),
.Y(n_225)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_228),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_220),
.B(n_190),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_229),
.B(n_233),
.C(n_147),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_218),
.B(n_182),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_231),
.B(n_237),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_232),
.B(n_212),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_220),
.B(n_205),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_222),
.B(n_209),
.C(n_201),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_236),
.B(n_240),
.C(n_183),
.Y(n_250)
);

FAx1_ASAP7_75t_L g237 ( 
.A(n_225),
.B(n_206),
.CI(n_175),
.CON(n_237),
.SN(n_237)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_211),
.B(n_159),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_239),
.B(n_3),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_222),
.B(n_196),
.C(n_202),
.Y(n_240)
);

INVxp67_ASAP7_75t_SL g241 ( 
.A(n_228),
.Y(n_241)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_241),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_242),
.B(n_244),
.Y(n_256)
);

OAI21xp5_ASAP7_75t_L g243 ( 
.A1(n_234),
.A2(n_213),
.B(n_226),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_243),
.B(n_249),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_229),
.B(n_210),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_235),
.A2(n_213),
.B1(n_216),
.B2(n_210),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_245),
.A2(n_237),
.B1(n_238),
.B2(n_230),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_246),
.B(n_236),
.C(n_240),
.Y(n_258)
);

BUFx24_ASAP7_75t_SL g249 ( 
.A(n_227),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_250),
.B(n_237),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_233),
.B(n_186),
.C(n_180),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_251),
.B(n_252),
.Y(n_253)
);

AND2x2_ASAP7_75t_L g270 ( 
.A(n_254),
.B(n_261),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_SL g268 ( 
.A(n_255),
.B(n_6),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_258),
.B(n_262),
.C(n_6),
.Y(n_267)
);

OAI21xp5_ASAP7_75t_L g259 ( 
.A1(n_250),
.A2(n_8),
.B(n_10),
.Y(n_259)
);

AOI21xp5_ASAP7_75t_L g263 ( 
.A1(n_259),
.A2(n_241),
.B(n_7),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_247),
.B(n_4),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_248),
.B(n_4),
.C(n_5),
.Y(n_262)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_263),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_257),
.B(n_253),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_264),
.B(n_265),
.Y(n_272)
);

INVxp67_ASAP7_75t_L g265 ( 
.A(n_256),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_261),
.B(n_6),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_266),
.B(n_267),
.Y(n_275)
);

INVxp67_ASAP7_75t_L g274 ( 
.A(n_268),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_254),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_L g271 ( 
.A1(n_269),
.A2(n_262),
.B(n_260),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_271),
.B(n_270),
.Y(n_276)
);

AOI21xp5_ASAP7_75t_L g279 ( 
.A1(n_276),
.A2(n_273),
.B(n_275),
.Y(n_279)
);

AOI21xp5_ASAP7_75t_L g277 ( 
.A1(n_272),
.A2(n_264),
.B(n_258),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_277),
.B(n_274),
.Y(n_278)
);

OAI21x1_ASAP7_75t_SL g280 ( 
.A1(n_278),
.A2(n_279),
.B(n_9),
.Y(n_280)
);

INVxp67_ASAP7_75t_L g281 ( 
.A(n_280),
.Y(n_281)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_281),
.B(n_12),
.Y(n_282)
);

AOI21xp5_ASAP7_75t_L g283 ( 
.A1(n_282),
.A2(n_12),
.B(n_270),
.Y(n_283)
);


endmodule