module fake_jpeg_1177_n_137 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_137);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_137;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_13),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_13),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_7),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_5),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_0),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_2),
.B(n_8),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

BUFx8_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_17),
.Y(n_30)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_30),
.Y(n_50)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_28),
.Y(n_31)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_31),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_17),
.Y(n_32)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_32),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_28),
.Y(n_33)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_33),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_26),
.B(n_21),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_34),
.B(n_3),
.Y(n_60)
);

INVx11_ASAP7_75t_L g35 ( 
.A(n_28),
.Y(n_35)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_35),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_14),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_36),
.B(n_19),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g37 ( 
.A(n_23),
.B(n_1),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_37),
.B(n_41),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_14),
.Y(n_38)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

INVx13_ASAP7_75t_L g39 ( 
.A(n_22),
.Y(n_39)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_39),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_22),
.Y(n_40)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g41 ( 
.A(n_23),
.B(n_2),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_38),
.Y(n_42)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_42),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g45 ( 
.A1(n_37),
.A2(n_24),
.B1(n_27),
.B2(n_29),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_45),
.A2(n_46),
.B1(n_56),
.B2(n_58),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g46 ( 
.A1(n_41),
.A2(n_24),
.B1(n_27),
.B2(n_29),
.Y(n_46)
);

AND2x2_ASAP7_75t_L g48 ( 
.A(n_33),
.B(n_25),
.Y(n_48)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_48),
.B(n_33),
.Y(n_63)
);

INVxp67_ASAP7_75t_L g75 ( 
.A(n_51),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_34),
.B(n_25),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_53),
.B(n_59),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_L g56 ( 
.A1(n_36),
.A2(n_18),
.B1(n_20),
.B2(n_16),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g58 ( 
.A1(n_38),
.A2(n_20),
.B1(n_16),
.B2(n_18),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_33),
.B(n_15),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_60),
.B(n_3),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_61),
.B(n_66),
.Y(n_86)
);

CKINVDCx16_ASAP7_75t_R g89 ( 
.A(n_63),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g64 ( 
.A1(n_46),
.A2(n_30),
.B1(n_32),
.B2(n_40),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_64),
.A2(n_71),
.B1(n_54),
.B2(n_50),
.Y(n_87)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_52),
.Y(n_65)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_65),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_57),
.B(n_31),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_57),
.B(n_4),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_67),
.B(n_75),
.Y(n_88)
);

HB1xp67_ASAP7_75t_L g69 ( 
.A(n_44),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_69),
.Y(n_80)
);

OAI22x1_ASAP7_75t_L g70 ( 
.A1(n_58),
.A2(n_40),
.B1(n_39),
.B2(n_35),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_70),
.A2(n_54),
.B1(n_50),
.B2(n_47),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_44),
.A2(n_31),
.B1(n_32),
.B2(n_30),
.Y(n_71)
);

A2O1A1Ixp33_ASAP7_75t_L g73 ( 
.A1(n_48),
.A2(n_39),
.B(n_5),
.C(n_6),
.Y(n_73)
);

XOR2x1_ASAP7_75t_L g82 ( 
.A(n_73),
.B(n_4),
.Y(n_82)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_55),
.Y(n_74)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_74),
.Y(n_84)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_52),
.Y(n_76)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_76),
.Y(n_85)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_55),
.Y(n_77)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_77),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_48),
.B(n_47),
.C(n_49),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_78),
.B(n_63),
.C(n_72),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_79),
.A2(n_87),
.B1(n_89),
.B2(n_80),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_82),
.B(n_90),
.Y(n_103)
);

XOR2xp5_ASAP7_75t_L g83 ( 
.A(n_66),
.B(n_49),
.Y(n_83)
);

XOR2xp5_ASAP7_75t_L g96 ( 
.A(n_83),
.B(n_93),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_88),
.B(n_73),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_78),
.B(n_9),
.Y(n_90)
);

INVx13_ASAP7_75t_L g92 ( 
.A(n_65),
.Y(n_92)
);

INVx13_ASAP7_75t_L g102 ( 
.A(n_92),
.Y(n_102)
);

XNOR2xp5_ASAP7_75t_SL g94 ( 
.A(n_93),
.B(n_62),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_94),
.B(n_90),
.C(n_83),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_86),
.B(n_75),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_95),
.B(n_98),
.Y(n_108)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_84),
.Y(n_97)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_97),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_88),
.B(n_68),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_79),
.A2(n_64),
.B1(n_71),
.B2(n_70),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_99),
.B(n_101),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_100),
.B(n_105),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_L g104 ( 
.A1(n_80),
.A2(n_76),
.B(n_43),
.Y(n_104)
);

AOI21xp5_ASAP7_75t_L g109 ( 
.A1(n_104),
.A2(n_85),
.B(n_81),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_92),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_107),
.B(n_114),
.C(n_94),
.Y(n_118)
);

INVx1_ASAP7_75t_SL g116 ( 
.A(n_109),
.Y(n_116)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_97),
.Y(n_112)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_112),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_103),
.B(n_85),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_113),
.B(n_91),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_96),
.B(n_84),
.C(n_91),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_111),
.Y(n_115)
);

HB1xp67_ASAP7_75t_L g122 ( 
.A(n_115),
.Y(n_122)
);

OR2x2_ASAP7_75t_L g126 ( 
.A(n_117),
.B(n_120),
.Y(n_126)
);

XOR2xp5_ASAP7_75t_L g125 ( 
.A(n_118),
.B(n_107),
.Y(n_125)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_106),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_110),
.A2(n_103),
.B1(n_99),
.B2(n_82),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_L g123 ( 
.A1(n_121),
.A2(n_108),
.B(n_110),
.Y(n_123)
);

NAND3xp33_ASAP7_75t_L g130 ( 
.A(n_123),
.B(n_104),
.C(n_81),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_115),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_124),
.B(n_119),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_125),
.B(n_116),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_L g132 ( 
.A1(n_127),
.A2(n_130),
.B(n_122),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_126),
.A2(n_116),
.B1(n_114),
.B2(n_96),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_128),
.B(n_129),
.C(n_102),
.Y(n_133)
);

AOI21xp5_ASAP7_75t_L g131 ( 
.A1(n_129),
.A2(n_122),
.B(n_102),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_131),
.B(n_133),
.C(n_43),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_132),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_134),
.B(n_135),
.C(n_10),
.Y(n_136)
);

XOR2xp5_ASAP7_75t_L g137 ( 
.A(n_136),
.B(n_10),
.Y(n_137)
);


endmodule