module fake_jpeg_11355_n_619 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_619);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_619;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_19;
wire n_182;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_582;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_387;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_615;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_384;
wire n_296;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_599;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_613;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx3_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

INVx6_ASAP7_75t_SL g19 ( 
.A(n_1),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_4),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_6),
.Y(n_22)
);

INVx11_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_4),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_17),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_11),
.Y(n_34)
);

HB1xp67_ASAP7_75t_L g35 ( 
.A(n_3),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_4),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_9),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_11),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_6),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_8),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_10),
.Y(n_41)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_1),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_16),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_0),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_10),
.Y(n_45)
);

INVx11_ASAP7_75t_L g46 ( 
.A(n_10),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_8),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_0),
.Y(n_48)
);

INVx11_ASAP7_75t_SL g49 ( 
.A(n_17),
.Y(n_49)
);

INVx11_ASAP7_75t_L g50 ( 
.A(n_16),
.Y(n_50)
);

INVx6_ASAP7_75t_SL g51 ( 
.A(n_12),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_15),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_8),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_4),
.Y(n_54)
);

BUFx5_ASAP7_75t_L g55 ( 
.A(n_7),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_1),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_11),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_5),
.Y(n_58)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_19),
.Y(n_59)
);

BUFx2_ASAP7_75t_L g154 ( 
.A(n_59),
.Y(n_154)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_42),
.Y(n_60)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_60),
.Y(n_134)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_29),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_61),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_26),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_62),
.Y(n_129)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_63),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_26),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_64),
.Y(n_148)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_42),
.Y(n_65)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_65),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_26),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_66),
.Y(n_161)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_19),
.Y(n_67)
);

INVx5_ASAP7_75t_L g140 ( 
.A(n_67),
.Y(n_140)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_27),
.Y(n_68)
);

INVx4_ASAP7_75t_L g151 ( 
.A(n_68),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_22),
.B(n_9),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g178 ( 
.A(n_69),
.B(n_80),
.Y(n_178)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_19),
.Y(n_70)
);

INVx5_ASAP7_75t_L g157 ( 
.A(n_70),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_26),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_71),
.Y(n_163)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_27),
.Y(n_72)
);

INVx4_ASAP7_75t_L g165 ( 
.A(n_72),
.Y(n_165)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_18),
.Y(n_73)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_73),
.Y(n_128)
);

INVx5_ASAP7_75t_L g74 ( 
.A(n_51),
.Y(n_74)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_74),
.Y(n_138)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_30),
.Y(n_75)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_75),
.Y(n_146)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_18),
.Y(n_76)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_76),
.Y(n_130)
);

BUFx4f_ASAP7_75t_SL g77 ( 
.A(n_51),
.Y(n_77)
);

BUFx8_ASAP7_75t_L g143 ( 
.A(n_77),
.Y(n_143)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_18),
.Y(n_78)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_78),
.Y(n_176)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_30),
.Y(n_79)
);

INVx3_ASAP7_75t_L g169 ( 
.A(n_79),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_22),
.B(n_9),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_54),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g170 ( 
.A(n_81),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_54),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g182 ( 
.A(n_82),
.Y(n_182)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_35),
.Y(n_83)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_83),
.Y(n_132)
);

BUFx3_ASAP7_75t_L g84 ( 
.A(n_27),
.Y(n_84)
);

INVx4_ASAP7_75t_L g204 ( 
.A(n_84),
.Y(n_204)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_55),
.Y(n_85)
);

INVx4_ASAP7_75t_L g145 ( 
.A(n_85),
.Y(n_145)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_35),
.Y(n_86)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_86),
.Y(n_137)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_30),
.Y(n_87)
);

INVx3_ASAP7_75t_L g171 ( 
.A(n_87),
.Y(n_171)
);

BUFx2_ASAP7_75t_L g88 ( 
.A(n_51),
.Y(n_88)
);

INVx1_ASAP7_75t_SL g152 ( 
.A(n_88),
.Y(n_152)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_55),
.Y(n_89)
);

INVx3_ASAP7_75t_L g177 ( 
.A(n_89),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_54),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g206 ( 
.A(n_90),
.Y(n_206)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_55),
.Y(n_91)
);

INVx3_ASAP7_75t_L g183 ( 
.A(n_91),
.Y(n_183)
);

BUFx12_ASAP7_75t_L g92 ( 
.A(n_46),
.Y(n_92)
);

BUFx8_ASAP7_75t_L g205 ( 
.A(n_92),
.Y(n_205)
);

BUFx5_ASAP7_75t_L g93 ( 
.A(n_46),
.Y(n_93)
);

INVx2_ASAP7_75t_SL g196 ( 
.A(n_93),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_43),
.B(n_9),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_94),
.B(n_112),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_54),
.Y(n_95)
);

INVx6_ASAP7_75t_L g133 ( 
.A(n_95),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_29),
.Y(n_96)
);

INVx6_ASAP7_75t_L g168 ( 
.A(n_96),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_29),
.Y(n_97)
);

INVx6_ASAP7_75t_L g208 ( 
.A(n_97),
.Y(n_208)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_36),
.Y(n_98)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_98),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_29),
.Y(n_99)
);

INVx4_ASAP7_75t_L g162 ( 
.A(n_99),
.Y(n_162)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_48),
.Y(n_100)
);

INVx3_ASAP7_75t_L g184 ( 
.A(n_100),
.Y(n_184)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_48),
.Y(n_101)
);

INVx3_ASAP7_75t_L g190 ( 
.A(n_101),
.Y(n_190)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_36),
.Y(n_102)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_102),
.Y(n_155)
);

INVx13_ASAP7_75t_L g103 ( 
.A(n_46),
.Y(n_103)
);

INVx4_ASAP7_75t_SL g172 ( 
.A(n_103),
.Y(n_172)
);

BUFx12f_ASAP7_75t_L g104 ( 
.A(n_48),
.Y(n_104)
);

INVx4_ASAP7_75t_L g167 ( 
.A(n_104),
.Y(n_167)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_36),
.Y(n_105)
);

INVx3_ASAP7_75t_L g198 ( 
.A(n_105),
.Y(n_198)
);

BUFx3_ASAP7_75t_L g106 ( 
.A(n_36),
.Y(n_106)
);

HB1xp67_ASAP7_75t_L g127 ( 
.A(n_106),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_32),
.Y(n_107)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_107),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_32),
.Y(n_108)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_108),
.Y(n_173)
);

INVx6_ASAP7_75t_L g109 ( 
.A(n_32),
.Y(n_109)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_109),
.Y(n_193)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_36),
.Y(n_110)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_110),
.Y(n_199)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_32),
.Y(n_111)
);

HB1xp67_ASAP7_75t_L g175 ( 
.A(n_111),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_43),
.B(n_8),
.Y(n_112)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_36),
.Y(n_113)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_113),
.Y(n_180)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_50),
.Y(n_114)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_114),
.Y(n_188)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_33),
.Y(n_115)
);

INVx4_ASAP7_75t_SL g174 ( 
.A(n_115),
.Y(n_174)
);

INVx8_ASAP7_75t_L g116 ( 
.A(n_33),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_116),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_33),
.Y(n_117)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_117),
.Y(n_209)
);

INVx11_ASAP7_75t_L g118 ( 
.A(n_23),
.Y(n_118)
);

INVx11_ASAP7_75t_L g141 ( 
.A(n_118),
.Y(n_141)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_33),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_119),
.B(n_124),
.Y(n_160)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_34),
.Y(n_120)
);

AND2x2_ASAP7_75t_L g192 ( 
.A(n_120),
.B(n_121),
.Y(n_192)
);

INVx8_ASAP7_75t_L g121 ( 
.A(n_50),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_34),
.Y(n_122)
);

NAND2xp33_ASAP7_75t_SL g139 ( 
.A(n_122),
.B(n_123),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_34),
.Y(n_123)
);

OR2x2_ASAP7_75t_L g124 ( 
.A(n_24),
.B(n_10),
.Y(n_124)
);

BUFx3_ASAP7_75t_L g125 ( 
.A(n_34),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_125),
.B(n_77),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_69),
.A2(n_57),
.B1(n_45),
.B2(n_53),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_131),
.A2(n_149),
.B1(n_150),
.B2(n_186),
.Y(n_244)
);

AOI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_88),
.A2(n_50),
.B1(n_53),
.B2(n_38),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_SL g220 ( 
.A1(n_136),
.A2(n_179),
.B1(n_181),
.B2(n_189),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_80),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_SL g217 ( 
.A(n_142),
.B(n_156),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_94),
.B(n_57),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_144),
.B(n_164),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_112),
.A2(n_53),
.B1(n_40),
.B2(n_38),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_124),
.A2(n_45),
.B1(n_53),
.B2(n_40),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_92),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_59),
.B(n_56),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_L g166 ( 
.A1(n_62),
.A2(n_38),
.B1(n_40),
.B2(n_21),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_166),
.A2(n_195),
.B1(n_202),
.B2(n_20),
.Y(n_223)
);

AOI22xp33_ASAP7_75t_SL g179 ( 
.A1(n_67),
.A2(n_70),
.B1(n_40),
.B2(n_38),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_SL g181 ( 
.A1(n_116),
.A2(n_23),
.B1(n_104),
.B2(n_52),
.Y(n_181)
);

OA22x2_ASAP7_75t_L g185 ( 
.A1(n_64),
.A2(n_21),
.B1(n_56),
.B2(n_25),
.Y(n_185)
);

OA22x2_ASAP7_75t_L g218 ( 
.A1(n_185),
.A2(n_39),
.B1(n_37),
.B2(n_41),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_96),
.A2(n_37),
.B1(n_39),
.B2(n_58),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_66),
.B(n_25),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_187),
.B(n_200),
.Y(n_222)
);

AOI22xp33_ASAP7_75t_SL g189 ( 
.A1(n_71),
.A2(n_23),
.B1(n_52),
.B2(n_47),
.Y(n_189)
);

INVxp67_ASAP7_75t_L g281 ( 
.A(n_191),
.Y(n_281)
);

AOI22xp33_ASAP7_75t_L g195 ( 
.A1(n_81),
.A2(n_24),
.B1(n_52),
.B2(n_28),
.Y(n_195)
);

AOI22xp33_ASAP7_75t_SL g197 ( 
.A1(n_82),
.A2(n_24),
.B1(n_28),
.B2(n_47),
.Y(n_197)
);

AOI22xp33_ASAP7_75t_SL g232 ( 
.A1(n_197),
.A2(n_20),
.B1(n_44),
.B2(n_41),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_90),
.B(n_58),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_95),
.B(n_58),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_201),
.B(n_185),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_97),
.A2(n_39),
.B1(n_37),
.B2(n_28),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_103),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_203),
.B(n_207),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_99),
.B(n_47),
.C(n_41),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_175),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_210),
.B(n_212),
.Y(n_303)
);

INVx6_ASAP7_75t_L g211 ( 
.A(n_129),
.Y(n_211)
);

INVx5_ASAP7_75t_L g291 ( 
.A(n_211),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_175),
.Y(n_212)
);

AND2x4_ASAP7_75t_SL g213 ( 
.A(n_132),
.B(n_122),
.Y(n_213)
);

AND2x2_ASAP7_75t_L g300 ( 
.A(n_213),
.B(n_218),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_127),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_214),
.B(n_216),
.Y(n_308)
);

INVx3_ASAP7_75t_L g215 ( 
.A(n_140),
.Y(n_215)
);

BUFx2_ASAP7_75t_L g283 ( 
.A(n_215),
.Y(n_283)
);

CKINVDCx16_ASAP7_75t_R g216 ( 
.A(n_127),
.Y(n_216)
);

BUFx6f_ASAP7_75t_L g221 ( 
.A(n_129),
.Y(n_221)
);

INVx4_ASAP7_75t_L g321 ( 
.A(n_221),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_223),
.A2(n_227),
.B1(n_251),
.B2(n_265),
.Y(n_292)
);

INVx1_ASAP7_75t_SL g224 ( 
.A(n_198),
.Y(n_224)
);

AND2x2_ASAP7_75t_L g335 ( 
.A(n_224),
.B(n_248),
.Y(n_335)
);

HB1xp67_ASAP7_75t_L g225 ( 
.A(n_184),
.Y(n_225)
);

INVxp67_ASAP7_75t_SL g334 ( 
.A(n_225),
.Y(n_334)
);

CKINVDCx14_ASAP7_75t_R g226 ( 
.A(n_143),
.Y(n_226)
);

NAND3xp33_ASAP7_75t_L g285 ( 
.A(n_226),
.B(n_234),
.C(n_262),
.Y(n_285)
);

OAI22xp33_ASAP7_75t_SL g227 ( 
.A1(n_185),
.A2(n_179),
.B1(n_136),
.B2(n_197),
.Y(n_227)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_193),
.Y(n_228)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_228),
.Y(n_296)
);

INVx6_ASAP7_75t_L g230 ( 
.A(n_148),
.Y(n_230)
);

INVx3_ASAP7_75t_L g320 ( 
.A(n_230),
.Y(n_320)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_159),
.Y(n_231)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_231),
.Y(n_301)
);

AOI21xp5_ASAP7_75t_L g295 ( 
.A1(n_232),
.A2(n_274),
.B(n_181),
.Y(n_295)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_173),
.Y(n_233)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_233),
.Y(n_311)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_134),
.Y(n_235)
);

INVx2_ASAP7_75t_SL g314 ( 
.A(n_235),
.Y(n_314)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_147),
.Y(n_236)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_236),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_194),
.B(n_31),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_SL g297 ( 
.A(n_237),
.B(n_245),
.Y(n_297)
);

CKINVDCx6p67_ASAP7_75t_R g238 ( 
.A(n_172),
.Y(n_238)
);

INVx4_ASAP7_75t_SL g318 ( 
.A(n_238),
.Y(n_318)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_155),
.Y(n_239)
);

INVx3_ASAP7_75t_L g330 ( 
.A(n_239),
.Y(n_330)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_199),
.Y(n_240)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_240),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_192),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_241),
.B(n_252),
.Y(n_319)
);

BUFx3_ASAP7_75t_L g242 ( 
.A(n_154),
.Y(n_242)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_242),
.Y(n_312)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_153),
.Y(n_243)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_243),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_160),
.B(n_31),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_158),
.Y(n_246)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_246),
.Y(n_326)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_209),
.Y(n_247)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_247),
.Y(n_332)
);

INVx3_ASAP7_75t_L g248 ( 
.A(n_157),
.Y(n_248)
);

AND2x2_ASAP7_75t_L g249 ( 
.A(n_152),
.B(n_123),
.Y(n_249)
);

CKINVDCx14_ASAP7_75t_R g289 ( 
.A(n_249),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_176),
.B(n_31),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_SL g317 ( 
.A(n_250),
.B(n_259),
.Y(n_317)
);

OAI22xp33_ASAP7_75t_SL g251 ( 
.A1(n_139),
.A2(n_117),
.B1(n_115),
.B2(n_111),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_180),
.Y(n_252)
);

BUFx3_ASAP7_75t_L g253 ( 
.A(n_154),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_253),
.B(n_254),
.Y(n_327)
);

INVx6_ASAP7_75t_L g254 ( 
.A(n_148),
.Y(n_254)
);

BUFx6f_ASAP7_75t_L g255 ( 
.A(n_161),
.Y(n_255)
);

AOI22xp33_ASAP7_75t_SL g284 ( 
.A1(n_255),
.A2(n_258),
.B1(n_269),
.B2(n_272),
.Y(n_284)
);

INVx2_ASAP7_75t_SL g256 ( 
.A(n_138),
.Y(n_256)
);

CKINVDCx16_ASAP7_75t_R g290 ( 
.A(n_256),
.Y(n_290)
);

HB1xp67_ASAP7_75t_L g257 ( 
.A(n_190),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_257),
.Y(n_304)
);

AOI22xp33_ASAP7_75t_SL g258 ( 
.A1(n_145),
.A2(n_108),
.B1(n_107),
.B2(n_49),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_137),
.B(n_20),
.Y(n_259)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_128),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_260),
.B(n_261),
.Y(n_336)
);

CKINVDCx16_ASAP7_75t_R g261 ( 
.A(n_143),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_178),
.B(n_44),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_130),
.B(n_44),
.Y(n_263)
);

NAND3xp33_ASAP7_75t_L g329 ( 
.A(n_263),
.B(n_266),
.C(n_275),
.Y(n_329)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_146),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_264),
.B(n_267),
.Y(n_337)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_166),
.A2(n_49),
.B1(n_1),
.B2(n_2),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_143),
.B(n_7),
.Y(n_266)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_169),
.Y(n_267)
);

INVx2_ASAP7_75t_SL g268 ( 
.A(n_171),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_268),
.Y(n_305)
);

AOI22xp33_ASAP7_75t_SL g269 ( 
.A1(n_145),
.A2(n_7),
.B1(n_16),
.B2(n_15),
.Y(n_269)
);

INVx3_ASAP7_75t_L g270 ( 
.A(n_205),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_270),
.Y(n_316)
);

INVx3_ASAP7_75t_L g271 ( 
.A(n_205),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_271),
.Y(n_322)
);

BUFx6f_ASAP7_75t_L g272 ( 
.A(n_161),
.Y(n_272)
);

OAI22xp33_ASAP7_75t_SL g273 ( 
.A1(n_189),
.A2(n_6),
.B1(n_16),
.B2(n_14),
.Y(n_273)
);

OA22x2_ASAP7_75t_L g338 ( 
.A1(n_273),
.A2(n_174),
.B1(n_11),
.B2(n_13),
.Y(n_338)
);

AOI22xp33_ASAP7_75t_SL g274 ( 
.A1(n_204),
.A2(n_6),
.B1(n_14),
.B2(n_13),
.Y(n_274)
);

OAI21xp33_ASAP7_75t_SL g275 ( 
.A1(n_195),
.A2(n_5),
.B(n_14),
.Y(n_275)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_162),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_276),
.Y(n_323)
);

INVx3_ASAP7_75t_L g277 ( 
.A(n_205),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_277),
.Y(n_325)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_126),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_278),
.B(n_279),
.Y(n_288)
);

BUFx2_ASAP7_75t_L g279 ( 
.A(n_167),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_177),
.B(n_5),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_SL g339 ( 
.A(n_280),
.B(n_17),
.Y(n_339)
);

BUFx2_ASAP7_75t_L g282 ( 
.A(n_167),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_282),
.B(n_135),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_SL g286 ( 
.A(n_229),
.B(n_192),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g371 ( 
.A(n_286),
.B(n_307),
.C(n_224),
.Y(n_371)
);

AOI22xp33_ASAP7_75t_L g287 ( 
.A1(n_223),
.A2(n_162),
.B1(n_133),
.B2(n_208),
.Y(n_287)
);

OAI21xp33_ASAP7_75t_SL g368 ( 
.A1(n_287),
.A2(n_294),
.B(n_328),
.Y(n_368)
);

AOI21xp33_ASAP7_75t_L g293 ( 
.A1(n_219),
.A2(n_172),
.B(n_135),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_293),
.B(n_238),
.Y(n_341)
);

AOI22xp33_ASAP7_75t_L g294 ( 
.A1(n_265),
.A2(n_133),
.B1(n_168),
.B2(n_208),
.Y(n_294)
);

A2O1A1Ixp33_ASAP7_75t_SL g367 ( 
.A1(n_295),
.A2(n_333),
.B(n_284),
.C(n_292),
.Y(n_367)
);

INVx1_ASAP7_75t_SL g361 ( 
.A(n_298),
.Y(n_361)
);

AOI21xp33_ASAP7_75t_SL g299 ( 
.A1(n_238),
.A2(n_141),
.B(n_151),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g363 ( 
.A(n_299),
.B(n_300),
.Y(n_363)
);

A2O1A1Ixp33_ASAP7_75t_L g306 ( 
.A1(n_222),
.A2(n_188),
.B(n_165),
.C(n_183),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_306),
.B(n_310),
.Y(n_350)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_281),
.B(n_196),
.C(n_126),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_218),
.B(n_168),
.Y(n_310)
);

NOR2x1_ASAP7_75t_L g313 ( 
.A(n_217),
.B(n_196),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_SL g378 ( 
.A(n_313),
.B(n_339),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_218),
.B(n_206),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_324),
.B(n_331),
.Y(n_356)
);

AOI22xp33_ASAP7_75t_L g328 ( 
.A1(n_244),
.A2(n_206),
.B1(n_182),
.B2(n_170),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_L g331 ( 
.A1(n_244),
.A2(n_182),
.B1(n_170),
.B2(n_163),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_L g358 ( 
.A1(n_331),
.A2(n_333),
.B1(n_249),
.B2(n_256),
.Y(n_358)
);

OAI22xp5_ASAP7_75t_L g333 ( 
.A1(n_220),
.A2(n_163),
.B1(n_174),
.B2(n_2),
.Y(n_333)
);

AND2x2_ASAP7_75t_L g366 ( 
.A(n_338),
.B(n_300),
.Y(n_366)
);

INVx3_ASAP7_75t_L g340 ( 
.A(n_291),
.Y(n_340)
);

INVx2_ASAP7_75t_L g393 ( 
.A(n_340),
.Y(n_393)
);

NAND3xp33_ASAP7_75t_L g402 ( 
.A(n_341),
.B(n_352),
.C(n_353),
.Y(n_402)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_288),
.Y(n_342)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_342),
.Y(n_391)
);

AOI21xp5_ASAP7_75t_L g343 ( 
.A1(n_295),
.A2(n_220),
.B(n_232),
.Y(n_343)
);

OAI21xp5_ASAP7_75t_SL g388 ( 
.A1(n_343),
.A2(n_367),
.B(n_372),
.Y(n_388)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_288),
.Y(n_344)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_344),
.Y(n_395)
);

CKINVDCx14_ASAP7_75t_R g345 ( 
.A(n_335),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_L g387 ( 
.A(n_345),
.B(n_349),
.Y(n_387)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_314),
.Y(n_346)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_346),
.Y(n_396)
);

MAJx2_ASAP7_75t_L g347 ( 
.A(n_286),
.B(n_213),
.C(n_281),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g400 ( 
.A(n_347),
.B(n_373),
.C(n_363),
.Y(n_400)
);

OR2x2_ASAP7_75t_L g348 ( 
.A(n_310),
.B(n_213),
.Y(n_348)
);

OAI21xp5_ASAP7_75t_L g389 ( 
.A1(n_348),
.A2(n_305),
.B(n_338),
.Y(n_389)
);

CKINVDCx20_ASAP7_75t_R g349 ( 
.A(n_303),
.Y(n_349)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_314),
.Y(n_351)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_351),
.Y(n_397)
);

INVxp67_ASAP7_75t_L g352 ( 
.A(n_336),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_297),
.B(n_238),
.Y(n_353)
);

OAI22xp5_ASAP7_75t_SL g354 ( 
.A1(n_292),
.A2(n_258),
.B1(n_269),
.B2(n_274),
.Y(n_354)
);

AOI22xp5_ASAP7_75t_L g408 ( 
.A1(n_354),
.A2(n_377),
.B1(n_379),
.B2(n_290),
.Y(n_408)
);

INVx2_ASAP7_75t_L g355 ( 
.A(n_283),
.Y(n_355)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_355),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_356),
.B(n_357),
.Y(n_392)
);

CKINVDCx20_ASAP7_75t_R g357 ( 
.A(n_337),
.Y(n_357)
);

OAI22xp5_ASAP7_75t_L g394 ( 
.A1(n_358),
.A2(n_364),
.B1(n_290),
.B2(n_302),
.Y(n_394)
);

INVx2_ASAP7_75t_SL g359 ( 
.A(n_291),
.Y(n_359)
);

AND2x2_ASAP7_75t_L g390 ( 
.A(n_359),
.B(n_363),
.Y(n_390)
);

INVxp67_ASAP7_75t_L g360 ( 
.A(n_335),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_360),
.B(n_362),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_L g362 ( 
.A(n_297),
.B(n_264),
.Y(n_362)
);

AOI22xp5_ASAP7_75t_L g364 ( 
.A1(n_324),
.A2(n_278),
.B1(n_228),
.B2(n_268),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g365 ( 
.A(n_313),
.B(n_236),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_365),
.B(n_370),
.Y(n_407)
);

AOI22xp5_ASAP7_75t_SL g384 ( 
.A1(n_366),
.A2(n_381),
.B1(n_383),
.B2(n_289),
.Y(n_384)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_314),
.Y(n_369)
);

INVx2_ASAP7_75t_SL g401 ( 
.A(n_369),
.Y(n_401)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_283),
.Y(n_370)
);

XNOR2xp5_ASAP7_75t_L g418 ( 
.A(n_371),
.B(n_309),
.Y(n_418)
);

AOI22xp5_ASAP7_75t_SL g372 ( 
.A1(n_300),
.A2(n_248),
.B1(n_215),
.B2(n_253),
.Y(n_372)
);

XOR2xp5_ASAP7_75t_L g373 ( 
.A(n_319),
.B(n_247),
.Y(n_373)
);

INVxp67_ASAP7_75t_L g374 ( 
.A(n_335),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_374),
.B(n_375),
.Y(n_411)
);

NOR2xp33_ASAP7_75t_L g375 ( 
.A(n_313),
.B(n_282),
.Y(n_375)
);

INVxp67_ASAP7_75t_L g376 ( 
.A(n_308),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_376),
.B(n_380),
.Y(n_412)
);

OAI22xp5_ASAP7_75t_L g377 ( 
.A1(n_317),
.A2(n_230),
.B1(n_254),
.B2(n_211),
.Y(n_377)
);

OAI22xp5_ASAP7_75t_SL g379 ( 
.A1(n_317),
.A2(n_233),
.B1(n_231),
.B2(n_255),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_339),
.B(n_242),
.Y(n_380)
);

OAI22xp33_ASAP7_75t_SL g381 ( 
.A1(n_306),
.A2(n_329),
.B1(n_285),
.B2(n_307),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_SL g382 ( 
.A(n_304),
.B(n_279),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_382),
.B(n_332),
.Y(n_420)
);

AOI22xp33_ASAP7_75t_SL g383 ( 
.A1(n_283),
.A2(n_277),
.B1(n_271),
.B2(n_270),
.Y(n_383)
);

OAI21xp5_ASAP7_75t_SL g426 ( 
.A1(n_384),
.A2(n_385),
.B(n_386),
.Y(n_426)
);

AOI22x1_ASAP7_75t_SL g385 ( 
.A1(n_354),
.A2(n_367),
.B1(n_343),
.B2(n_341),
.Y(n_385)
);

AOI32xp33_ASAP7_75t_L g386 ( 
.A1(n_350),
.A2(n_298),
.A3(n_299),
.B1(n_304),
.B2(n_305),
.Y(n_386)
);

INVxp67_ASAP7_75t_L g431 ( 
.A(n_389),
.Y(n_431)
);

AOI22xp5_ASAP7_75t_L g427 ( 
.A1(n_394),
.A2(n_398),
.B1(n_404),
.B2(n_413),
.Y(n_427)
);

OAI22xp5_ASAP7_75t_SL g398 ( 
.A1(n_356),
.A2(n_348),
.B1(n_350),
.B2(n_358),
.Y(n_398)
);

XOR2xp5_ASAP7_75t_L g437 ( 
.A(n_400),
.B(n_378),
.Y(n_437)
);

OAI22xp5_ASAP7_75t_SL g404 ( 
.A1(n_348),
.A2(n_338),
.B1(n_315),
.B2(n_326),
.Y(n_404)
);

AOI22xp5_ASAP7_75t_SL g405 ( 
.A1(n_366),
.A2(n_338),
.B1(n_325),
.B2(n_322),
.Y(n_405)
);

OAI21xp5_ASAP7_75t_SL g448 ( 
.A1(n_405),
.A2(n_406),
.B(n_409),
.Y(n_448)
);

AOI22xp5_ASAP7_75t_SL g406 ( 
.A1(n_366),
.A2(n_322),
.B1(n_316),
.B2(n_325),
.Y(n_406)
);

BUFx3_ASAP7_75t_L g429 ( 
.A(n_408),
.Y(n_429)
);

OA21x2_ASAP7_75t_L g409 ( 
.A1(n_365),
.A2(n_327),
.B(n_318),
.Y(n_409)
);

CKINVDCx20_ASAP7_75t_R g410 ( 
.A(n_382),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_L g433 ( 
.A(n_410),
.B(n_415),
.Y(n_433)
);

OAI22xp5_ASAP7_75t_L g413 ( 
.A1(n_342),
.A2(n_344),
.B1(n_367),
.B2(n_361),
.Y(n_413)
);

AND2x2_ASAP7_75t_L g414 ( 
.A(n_375),
.B(n_318),
.Y(n_414)
);

INVxp67_ASAP7_75t_L g434 ( 
.A(n_414),
.Y(n_434)
);

CKINVDCx20_ASAP7_75t_R g415 ( 
.A(n_353),
.Y(n_415)
);

OAI22xp5_ASAP7_75t_SL g416 ( 
.A1(n_367),
.A2(n_315),
.B1(n_326),
.B2(n_320),
.Y(n_416)
);

AOI22xp5_ASAP7_75t_L g428 ( 
.A1(n_416),
.A2(n_417),
.B1(n_377),
.B2(n_351),
.Y(n_428)
);

OAI22xp5_ASAP7_75t_SL g417 ( 
.A1(n_367),
.A2(n_320),
.B1(n_272),
.B2(n_221),
.Y(n_417)
);

MAJIxp5_ASAP7_75t_L g421 ( 
.A(n_418),
.B(n_371),
.C(n_373),
.Y(n_421)
);

AOI22xp5_ASAP7_75t_L g419 ( 
.A1(n_368),
.A2(n_321),
.B1(n_316),
.B2(n_332),
.Y(n_419)
);

OAI22xp5_ASAP7_75t_SL g440 ( 
.A1(n_419),
.A2(n_369),
.B1(n_346),
.B2(n_359),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_420),
.B(n_379),
.Y(n_423)
);

MAJIxp5_ASAP7_75t_L g469 ( 
.A(n_421),
.B(n_424),
.C(n_425),
.Y(n_469)
);

INVx8_ASAP7_75t_L g422 ( 
.A(n_393),
.Y(n_422)
);

INVx2_ASAP7_75t_L g467 ( 
.A(n_422),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_423),
.B(n_435),
.Y(n_456)
);

MAJIxp5_ASAP7_75t_L g424 ( 
.A(n_418),
.B(n_347),
.C(n_361),
.Y(n_424)
);

MAJIxp5_ASAP7_75t_L g425 ( 
.A(n_400),
.B(n_347),
.C(n_349),
.Y(n_425)
);

OAI22xp5_ASAP7_75t_L g468 ( 
.A1(n_428),
.A2(n_450),
.B1(n_453),
.B2(n_454),
.Y(n_468)
);

MAJIxp5_ASAP7_75t_L g430 ( 
.A(n_390),
.B(n_357),
.C(n_362),
.Y(n_430)
);

MAJIxp5_ASAP7_75t_L g476 ( 
.A(n_430),
.B(n_437),
.C(n_449),
.Y(n_476)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_396),
.Y(n_432)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_432),
.Y(n_479)
);

CKINVDCx20_ASAP7_75t_R g435 ( 
.A(n_420),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_SL g436 ( 
.A(n_415),
.B(n_378),
.Y(n_436)
);

CKINVDCx14_ASAP7_75t_R g473 ( 
.A(n_436),
.Y(n_473)
);

CKINVDCx20_ASAP7_75t_R g438 ( 
.A(n_392),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_438),
.B(n_452),
.Y(n_460)
);

OAI22xp5_ASAP7_75t_L g439 ( 
.A1(n_392),
.A2(n_364),
.B1(n_372),
.B2(n_380),
.Y(n_439)
);

AOI22xp5_ASAP7_75t_L g458 ( 
.A1(n_439),
.A2(n_440),
.B1(n_441),
.B2(n_446),
.Y(n_458)
);

OAI22xp5_ASAP7_75t_SL g441 ( 
.A1(n_405),
.A2(n_359),
.B1(n_340),
.B2(n_321),
.Y(n_441)
);

INVxp67_ASAP7_75t_SL g442 ( 
.A(n_387),
.Y(n_442)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_442),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_410),
.B(n_370),
.Y(n_443)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_443),
.Y(n_457)
);

AOI21xp5_ASAP7_75t_L g444 ( 
.A1(n_388),
.A2(n_318),
.B(n_355),
.Y(n_444)
);

HB1xp67_ASAP7_75t_L g474 ( 
.A(n_444),
.Y(n_474)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_396),
.Y(n_445)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_445),
.Y(n_461)
);

OAI22xp5_ASAP7_75t_L g446 ( 
.A1(n_385),
.A2(n_323),
.B1(n_302),
.B2(n_309),
.Y(n_446)
);

CKINVDCx16_ASAP7_75t_R g447 ( 
.A(n_414),
.Y(n_447)
);

NOR2xp33_ASAP7_75t_L g471 ( 
.A(n_447),
.B(n_414),
.Y(n_471)
);

XNOR2xp5_ASAP7_75t_L g449 ( 
.A(n_412),
.B(n_334),
.Y(n_449)
);

AOI22xp5_ASAP7_75t_L g450 ( 
.A1(n_413),
.A2(n_323),
.B1(n_312),
.B2(n_330),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_397),
.Y(n_451)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_451),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_391),
.B(n_296),
.Y(n_452)
);

AOI22xp5_ASAP7_75t_L g453 ( 
.A1(n_398),
.A2(n_312),
.B1(n_330),
.B2(n_296),
.Y(n_453)
);

AOI22xp5_ASAP7_75t_SL g454 ( 
.A1(n_416),
.A2(n_311),
.B1(n_301),
.B2(n_13),
.Y(n_454)
);

CKINVDCx16_ASAP7_75t_R g459 ( 
.A(n_443),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_SL g514 ( 
.A(n_459),
.B(n_401),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_438),
.B(n_395),
.Y(n_462)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_462),
.Y(n_487)
);

AOI22xp5_ASAP7_75t_L g463 ( 
.A1(n_429),
.A2(n_446),
.B1(n_441),
.B2(n_439),
.Y(n_463)
);

OAI22xp5_ASAP7_75t_SL g503 ( 
.A1(n_463),
.A2(n_480),
.B1(n_428),
.B2(n_450),
.Y(n_503)
);

NAND3xp33_ASAP7_75t_L g464 ( 
.A(n_436),
.B(n_433),
.C(n_412),
.Y(n_464)
);

NOR2xp33_ASAP7_75t_L g489 ( 
.A(n_464),
.B(n_478),
.Y(n_489)
);

OAI22xp5_ASAP7_75t_SL g465 ( 
.A1(n_427),
.A2(n_408),
.B1(n_384),
.B2(n_395),
.Y(n_465)
);

AOI22xp5_ASAP7_75t_L g490 ( 
.A1(n_465),
.A2(n_472),
.B1(n_429),
.B2(n_409),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_435),
.B(n_391),
.Y(n_466)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_466),
.Y(n_488)
);

AND2x2_ASAP7_75t_SL g470 ( 
.A(n_448),
.B(n_388),
.Y(n_470)
);

INVxp67_ASAP7_75t_L g501 ( 
.A(n_470),
.Y(n_501)
);

AND2x2_ASAP7_75t_L g512 ( 
.A(n_471),
.B(n_485),
.Y(n_512)
);

OAI22xp5_ASAP7_75t_SL g472 ( 
.A1(n_427),
.A2(n_389),
.B1(n_406),
.B2(n_419),
.Y(n_472)
);

XOR2xp5_ASAP7_75t_L g475 ( 
.A(n_437),
.B(n_390),
.Y(n_475)
);

XOR2xp5_ASAP7_75t_L g510 ( 
.A(n_475),
.B(n_482),
.Y(n_510)
);

INVx1_ASAP7_75t_SL g477 ( 
.A(n_432),
.Y(n_477)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_477),
.Y(n_504)
);

FAx1_ASAP7_75t_SL g478 ( 
.A(n_425),
.B(n_424),
.CI(n_430),
.CON(n_478),
.SN(n_478)
);

AOI22xp5_ASAP7_75t_L g480 ( 
.A1(n_429),
.A2(n_417),
.B1(n_394),
.B2(n_404),
.Y(n_480)
);

XOR2xp5_ASAP7_75t_L g482 ( 
.A(n_421),
.B(n_390),
.Y(n_482)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_422),
.Y(n_483)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_483),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_433),
.B(n_397),
.Y(n_484)
);

CKINVDCx20_ASAP7_75t_R g496 ( 
.A(n_484),
.Y(n_496)
);

INVx2_ASAP7_75t_SL g485 ( 
.A(n_445),
.Y(n_485)
);

OAI21xp33_ASAP7_75t_L g486 ( 
.A1(n_426),
.A2(n_411),
.B(n_403),
.Y(n_486)
);

CKINVDCx20_ASAP7_75t_R g498 ( 
.A(n_486),
.Y(n_498)
);

OAI22xp5_ASAP7_75t_SL g532 ( 
.A1(n_490),
.A2(n_485),
.B1(n_481),
.B2(n_461),
.Y(n_532)
);

MAJIxp5_ASAP7_75t_L g491 ( 
.A(n_482),
.B(n_469),
.C(n_475),
.Y(n_491)
);

MAJIxp5_ASAP7_75t_L g517 ( 
.A(n_491),
.B(n_492),
.C(n_493),
.Y(n_517)
);

MAJIxp5_ASAP7_75t_L g492 ( 
.A(n_469),
.B(n_447),
.C(n_449),
.Y(n_492)
);

MAJIxp5_ASAP7_75t_L g493 ( 
.A(n_476),
.B(n_434),
.C(n_431),
.Y(n_493)
);

NOR2xp33_ASAP7_75t_L g494 ( 
.A(n_455),
.B(n_403),
.Y(n_494)
);

NOR2xp33_ASAP7_75t_SL g538 ( 
.A(n_494),
.B(n_495),
.Y(n_538)
);

NOR2xp33_ASAP7_75t_L g495 ( 
.A(n_455),
.B(n_453),
.Y(n_495)
);

XNOR2xp5_ASAP7_75t_SL g497 ( 
.A(n_476),
.B(n_478),
.Y(n_497)
);

XOR2xp5_ASAP7_75t_L g524 ( 
.A(n_497),
.B(n_470),
.Y(n_524)
);

CKINVDCx20_ASAP7_75t_R g499 ( 
.A(n_460),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_499),
.B(n_500),
.Y(n_518)
);

CKINVDCx20_ASAP7_75t_R g500 ( 
.A(n_460),
.Y(n_500)
);

AOI21xp5_ASAP7_75t_L g502 ( 
.A1(n_474),
.A2(n_448),
.B(n_426),
.Y(n_502)
);

OAI21xp5_ASAP7_75t_L g519 ( 
.A1(n_502),
.A2(n_507),
.B(n_470),
.Y(n_519)
);

AOI22xp5_ASAP7_75t_L g525 ( 
.A1(n_503),
.A2(n_509),
.B1(n_468),
.B2(n_457),
.Y(n_525)
);

OAI22xp5_ASAP7_75t_L g505 ( 
.A1(n_473),
.A2(n_386),
.B1(n_454),
.B2(n_423),
.Y(n_505)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_505),
.Y(n_520)
);

A2O1A1Ixp33_ASAP7_75t_L g506 ( 
.A1(n_456),
.A2(n_411),
.B(n_407),
.C(n_402),
.Y(n_506)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_506),
.Y(n_522)
);

AOI21xp5_ASAP7_75t_SL g507 ( 
.A1(n_456),
.A2(n_444),
.B(n_407),
.Y(n_507)
);

MAJIxp5_ASAP7_75t_L g508 ( 
.A(n_478),
.B(n_451),
.C(n_409),
.Y(n_508)
);

MAJIxp5_ASAP7_75t_L g531 ( 
.A(n_508),
.B(n_480),
.C(n_477),
.Y(n_531)
);

OAI22xp5_ASAP7_75t_L g509 ( 
.A1(n_458),
.A2(n_452),
.B1(n_440),
.B2(n_409),
.Y(n_509)
);

CKINVDCx20_ASAP7_75t_R g513 ( 
.A(n_462),
.Y(n_513)
);

AOI22xp33_ASAP7_75t_L g523 ( 
.A1(n_513),
.A2(n_515),
.B1(n_457),
.B2(n_472),
.Y(n_523)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_514),
.Y(n_521)
);

CKINVDCx20_ASAP7_75t_R g515 ( 
.A(n_484),
.Y(n_515)
);

XNOR2xp5_ASAP7_75t_L g516 ( 
.A(n_493),
.B(n_465),
.Y(n_516)
);

XNOR2xp5_ASAP7_75t_L g546 ( 
.A(n_516),
.B(n_519),
.Y(n_546)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_523),
.Y(n_545)
);

XOR2xp5_ASAP7_75t_L g540 ( 
.A(n_524),
.B(n_510),
.Y(n_540)
);

OAI22xp5_ASAP7_75t_SL g556 ( 
.A1(n_525),
.A2(n_507),
.B1(n_488),
.B2(n_487),
.Y(n_556)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_504),
.Y(n_526)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_526),
.Y(n_554)
);

CKINVDCx14_ASAP7_75t_R g527 ( 
.A(n_512),
.Y(n_527)
);

OAI22xp5_ASAP7_75t_L g552 ( 
.A1(n_527),
.A2(n_528),
.B1(n_534),
.B2(n_513),
.Y(n_552)
);

AOI22xp5_ASAP7_75t_L g528 ( 
.A1(n_503),
.A2(n_466),
.B1(n_458),
.B2(n_463),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_504),
.Y(n_529)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_529),
.Y(n_555)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_512),
.Y(n_530)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_530),
.Y(n_547)
);

XNOR2xp5_ASAP7_75t_L g551 ( 
.A(n_531),
.B(n_535),
.Y(n_551)
);

AOI22xp5_ASAP7_75t_L g549 ( 
.A1(n_532),
.A2(n_536),
.B1(n_488),
.B2(n_487),
.Y(n_549)
);

OAI22xp5_ASAP7_75t_L g533 ( 
.A1(n_489),
.A2(n_485),
.B1(n_481),
.B2(n_461),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_SL g544 ( 
.A(n_533),
.B(n_515),
.Y(n_544)
);

AOI22xp5_ASAP7_75t_L g534 ( 
.A1(n_509),
.A2(n_479),
.B1(n_483),
.B2(n_467),
.Y(n_534)
);

XNOR2xp5_ASAP7_75t_L g535 ( 
.A(n_492),
.B(n_401),
.Y(n_535)
);

OAI22xp5_ASAP7_75t_SL g536 ( 
.A1(n_490),
.A2(n_467),
.B1(n_401),
.B2(n_422),
.Y(n_536)
);

HB1xp67_ASAP7_75t_L g537 ( 
.A(n_506),
.Y(n_537)
);

INVxp33_ASAP7_75t_L g557 ( 
.A(n_537),
.Y(n_557)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_512),
.Y(n_539)
);

NOR2xp33_ASAP7_75t_L g548 ( 
.A(n_539),
.B(n_531),
.Y(n_548)
);

XOR2xp5_ASAP7_75t_L g566 ( 
.A(n_540),
.B(n_502),
.Y(n_566)
);

CKINVDCx16_ASAP7_75t_R g541 ( 
.A(n_518),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_L g576 ( 
.A(n_541),
.B(n_543),
.Y(n_576)
);

FAx1_ASAP7_75t_SL g542 ( 
.A(n_518),
.B(n_508),
.CI(n_501),
.CON(n_542),
.SN(n_542)
);

NOR2xp33_ASAP7_75t_L g563 ( 
.A(n_542),
.B(n_553),
.Y(n_563)
);

CKINVDCx16_ASAP7_75t_R g543 ( 
.A(n_538),
.Y(n_543)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_544),
.Y(n_560)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_548),
.Y(n_562)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_549),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_SL g550 ( 
.A(n_517),
.B(n_491),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_SL g570 ( 
.A(n_550),
.B(n_559),
.Y(n_570)
);

AOI22xp5_ASAP7_75t_L g565 ( 
.A1(n_552),
.A2(n_556),
.B1(n_532),
.B2(n_500),
.Y(n_565)
);

BUFx4f_ASAP7_75t_SL g553 ( 
.A(n_536),
.Y(n_553)
);

XNOR2xp5_ASAP7_75t_L g558 ( 
.A(n_535),
.B(n_497),
.Y(n_558)
);

NOR2xp67_ASAP7_75t_SL g568 ( 
.A(n_558),
.B(n_524),
.Y(n_568)
);

MAJIxp5_ASAP7_75t_L g559 ( 
.A(n_517),
.B(n_510),
.C(n_501),
.Y(n_559)
);

XNOR2xp5_ASAP7_75t_L g561 ( 
.A(n_551),
.B(n_516),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_L g587 ( 
.A(n_561),
.B(n_565),
.Y(n_587)
);

AOI21xp5_ASAP7_75t_L g564 ( 
.A1(n_559),
.A2(n_519),
.B(n_522),
.Y(n_564)
);

AOI21xp5_ASAP7_75t_L g581 ( 
.A1(n_564),
.A2(n_575),
.B(n_547),
.Y(n_581)
);

XOR2xp5_ASAP7_75t_L g583 ( 
.A(n_566),
.B(n_568),
.Y(n_583)
);

XNOR2xp5_ASAP7_75t_L g567 ( 
.A(n_551),
.B(n_520),
.Y(n_567)
);

NOR2xp33_ASAP7_75t_L g579 ( 
.A(n_567),
.B(n_572),
.Y(n_579)
);

MAJIxp5_ASAP7_75t_L g569 ( 
.A(n_546),
.B(n_530),
.C(n_525),
.Y(n_569)
);

MAJIxp5_ASAP7_75t_L g577 ( 
.A(n_569),
.B(n_571),
.C(n_545),
.Y(n_577)
);

MAJIxp5_ASAP7_75t_L g571 ( 
.A(n_546),
.B(n_528),
.C(n_534),
.Y(n_571)
);

NOR2xp33_ASAP7_75t_L g572 ( 
.A(n_557),
.B(n_522),
.Y(n_572)
);

AOI22xp5_ASAP7_75t_L g573 ( 
.A1(n_557),
.A2(n_521),
.B1(n_499),
.B2(n_498),
.Y(n_573)
);

OAI22xp5_ASAP7_75t_L g582 ( 
.A1(n_573),
.A2(n_549),
.B1(n_547),
.B2(n_496),
.Y(n_582)
);

OAI21xp5_ASAP7_75t_L g575 ( 
.A1(n_556),
.A2(n_498),
.B(n_496),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_SL g590 ( 
.A(n_577),
.B(n_578),
.Y(n_590)
);

INVx11_ASAP7_75t_L g578 ( 
.A(n_576),
.Y(n_578)
);

NOR2xp33_ASAP7_75t_L g580 ( 
.A(n_570),
.B(n_542),
.Y(n_580)
);

NOR2xp33_ASAP7_75t_L g598 ( 
.A(n_580),
.B(n_585),
.Y(n_598)
);

OAI21xp5_ASAP7_75t_L g597 ( 
.A1(n_581),
.A2(n_566),
.B(n_399),
.Y(n_597)
);

AO21x1_ASAP7_75t_L g593 ( 
.A1(n_582),
.A2(n_586),
.B(n_563),
.Y(n_593)
);

AOI22xp33_ASAP7_75t_SL g584 ( 
.A1(n_560),
.A2(n_554),
.B1(n_555),
.B2(n_529),
.Y(n_584)
);

INVxp67_ASAP7_75t_L g591 ( 
.A(n_584),
.Y(n_591)
);

MAJIxp5_ASAP7_75t_L g585 ( 
.A(n_561),
.B(n_558),
.C(n_540),
.Y(n_585)
);

OAI21xp5_ASAP7_75t_L g586 ( 
.A1(n_575),
.A2(n_542),
.B(n_553),
.Y(n_586)
);

MAJIxp5_ASAP7_75t_L g588 ( 
.A(n_571),
.B(n_553),
.C(n_511),
.Y(n_588)
);

XNOR2xp5_ASAP7_75t_L g595 ( 
.A(n_588),
.B(n_589),
.Y(n_595)
);

MAJIxp5_ASAP7_75t_L g589 ( 
.A(n_569),
.B(n_511),
.C(n_393),
.Y(n_589)
);

XNOR2x2_ASAP7_75t_L g592 ( 
.A(n_585),
.B(n_567),
.Y(n_592)
);

AOI21xp33_ASAP7_75t_L g600 ( 
.A1(n_592),
.A2(n_597),
.B(n_578),
.Y(n_600)
);

AOI21xp5_ASAP7_75t_L g601 ( 
.A1(n_593),
.A2(n_594),
.B(n_596),
.Y(n_601)
);

MAJIxp5_ASAP7_75t_L g594 ( 
.A(n_577),
.B(n_562),
.C(n_574),
.Y(n_594)
);

AO21x1_ASAP7_75t_L g596 ( 
.A1(n_586),
.A2(n_573),
.B(n_565),
.Y(n_596)
);

XNOR2xp5_ASAP7_75t_L g599 ( 
.A(n_587),
.B(n_583),
.Y(n_599)
);

NOR2xp33_ASAP7_75t_SL g605 ( 
.A(n_599),
.B(n_311),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_SL g608 ( 
.A(n_600),
.B(n_604),
.Y(n_608)
);

AOI22xp5_ASAP7_75t_L g602 ( 
.A1(n_591),
.A2(n_588),
.B1(n_589),
.B2(n_583),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_L g607 ( 
.A(n_602),
.B(n_603),
.Y(n_607)
);

AOI22xp5_ASAP7_75t_SL g603 ( 
.A1(n_593),
.A2(n_581),
.B1(n_579),
.B2(n_399),
.Y(n_603)
);

NOR2xp33_ASAP7_75t_L g604 ( 
.A(n_595),
.B(n_598),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_SL g611 ( 
.A(n_605),
.B(n_606),
.Y(n_611)
);

NOR2xp33_ASAP7_75t_L g606 ( 
.A(n_598),
.B(n_301),
.Y(n_606)
);

OAI21xp5_ASAP7_75t_SL g609 ( 
.A1(n_601),
.A2(n_590),
.B(n_596),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_L g613 ( 
.A(n_609),
.B(n_0),
.Y(n_613)
);

NOR2xp33_ASAP7_75t_L g610 ( 
.A(n_603),
.B(n_13),
.Y(n_610)
);

NOR2xp33_ASAP7_75t_SL g612 ( 
.A(n_610),
.B(n_17),
.Y(n_612)
);

MAJIxp5_ASAP7_75t_L g614 ( 
.A(n_612),
.B(n_613),
.C(n_611),
.Y(n_614)
);

OAI22xp5_ASAP7_75t_L g615 ( 
.A1(n_614),
.A2(n_608),
.B1(n_607),
.B2(n_2),
.Y(n_615)
);

AOI21xp5_ASAP7_75t_L g616 ( 
.A1(n_615),
.A2(n_0),
.B(n_1),
.Y(n_616)
);

MAJx2_ASAP7_75t_L g617 ( 
.A(n_616),
.B(n_0),
.C(n_2),
.Y(n_617)
);

OAI21xp5_ASAP7_75t_L g618 ( 
.A1(n_617),
.A2(n_3),
.B(n_464),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_L g619 ( 
.A(n_618),
.B(n_3),
.Y(n_619)
);


endmodule