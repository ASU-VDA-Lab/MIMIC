module fake_aes_2826_n_41 (n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_41);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_41;
wire n_20;
wire n_38;
wire n_36;
wire n_37;
wire n_34;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_30;
wire n_13;
wire n_33;
wire n_26;
wire n_18;
wire n_32;
wire n_35;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_27;
wire n_21;
wire n_40;
wire n_29;
wire n_39;
INVx2_ASAP7_75t_L g11 ( .A(n_5), .Y(n_11) );
INVx1_ASAP7_75t_L g12 ( .A(n_1), .Y(n_12) );
NOR2xp67_ASAP7_75t_L g13 ( .A(n_9), .B(n_5), .Y(n_13) );
CKINVDCx5p33_ASAP7_75t_R g14 ( .A(n_1), .Y(n_14) );
INVx1_ASAP7_75t_L g15 ( .A(n_8), .Y(n_15) );
INVx1_ASAP7_75t_L g16 ( .A(n_9), .Y(n_16) );
AOI22xp5_ASAP7_75t_L g17 ( .A1(n_6), .A2(n_8), .B1(n_0), .B2(n_2), .Y(n_17) );
INVxp67_ASAP7_75t_SL g18 ( .A(n_12), .Y(n_18) );
HB1xp67_ASAP7_75t_L g19 ( .A(n_14), .Y(n_19) );
NAND2xp5_ASAP7_75t_L g20 ( .A(n_12), .B(n_0), .Y(n_20) );
NAND2xp33_ASAP7_75t_SL g21 ( .A(n_14), .B(n_2), .Y(n_21) );
CKINVDCx5p33_ASAP7_75t_R g22 ( .A(n_17), .Y(n_22) );
AOI22xp33_ASAP7_75t_L g23 ( .A1(n_18), .A2(n_16), .B1(n_15), .B2(n_11), .Y(n_23) );
AOI22xp33_ASAP7_75t_L g24 ( .A1(n_18), .A2(n_16), .B1(n_11), .B2(n_13), .Y(n_24) );
INVx3_ASAP7_75t_L g25 ( .A(n_20), .Y(n_25) );
BUFx2_ASAP7_75t_R g26 ( .A(n_22), .Y(n_26) );
OAI211xp5_ASAP7_75t_L g27 ( .A1(n_23), .A2(n_19), .B(n_20), .C(n_21), .Y(n_27) );
AOI211xp5_ASAP7_75t_L g28 ( .A1(n_25), .A2(n_19), .B(n_4), .C(n_6), .Y(n_28) );
AO21x2_ASAP7_75t_L g29 ( .A1(n_25), .A2(n_3), .B(n_4), .Y(n_29) );
INVx1_ASAP7_75t_L g30 ( .A(n_29), .Y(n_30) );
HB1xp67_ASAP7_75t_L g31 ( .A(n_29), .Y(n_31) );
OR2x2_ASAP7_75t_L g32 ( .A(n_30), .B(n_25), .Y(n_32) );
AND2x2_ASAP7_75t_L g33 ( .A(n_31), .B(n_24), .Y(n_33) );
NOR2x1_ASAP7_75t_L g34 ( .A(n_32), .B(n_29), .Y(n_34) );
AOI21xp33_ASAP7_75t_SL g35 ( .A1(n_33), .A2(n_26), .B(n_27), .Y(n_35) );
INVx1_ASAP7_75t_SL g36 ( .A(n_32), .Y(n_36) );
CKINVDCx5p33_ASAP7_75t_R g37 ( .A(n_36), .Y(n_37) );
OAI22x1_ASAP7_75t_L g38 ( .A1(n_34), .A2(n_30), .B1(n_28), .B2(n_7), .Y(n_38) );
INVx1_ASAP7_75t_L g39 ( .A(n_38), .Y(n_39) );
AOI31xp33_ASAP7_75t_L g40 ( .A1(n_37), .A2(n_35), .A3(n_7), .B(n_3), .Y(n_40) );
AOI22xp5_ASAP7_75t_L g41 ( .A1(n_39), .A2(n_10), .B1(n_38), .B2(n_40), .Y(n_41) );
endmodule