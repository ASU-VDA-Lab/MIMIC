module fake_netlist_1_8418_n_38 (n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_38);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_38;
wire n_20;
wire n_36;
wire n_37;
wire n_34;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_30;
wire n_33;
wire n_18;
wire n_32;
wire n_35;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_27;
NOR2xp33_ASAP7_75t_R g11 ( .A(n_0), .B(n_9), .Y(n_11) );
NAND2xp5_ASAP7_75t_L g12 ( .A(n_9), .B(n_4), .Y(n_12) );
INVx2_ASAP7_75t_L g13 ( .A(n_1), .Y(n_13) );
NOR2xp67_ASAP7_75t_L g14 ( .A(n_3), .B(n_10), .Y(n_14) );
CKINVDCx20_ASAP7_75t_R g15 ( .A(n_10), .Y(n_15) );
INVx1_ASAP7_75t_L g16 ( .A(n_2), .Y(n_16) );
BUFx6f_ASAP7_75t_L g17 ( .A(n_7), .Y(n_17) );
INVx6_ASAP7_75t_L g18 ( .A(n_17), .Y(n_18) );
OAI21x1_ASAP7_75t_L g19 ( .A1(n_13), .A2(n_0), .B(n_1), .Y(n_19) );
INVxp67_ASAP7_75t_L g20 ( .A(n_16), .Y(n_20) );
INVx2_ASAP7_75t_L g21 ( .A(n_13), .Y(n_21) );
NAND2xp5_ASAP7_75t_L g22 ( .A(n_16), .B(n_0), .Y(n_22) );
OAI22xp5_ASAP7_75t_L g23 ( .A1(n_20), .A2(n_13), .B1(n_12), .B2(n_15), .Y(n_23) );
AND2x2_ASAP7_75t_L g24 ( .A(n_22), .B(n_17), .Y(n_24) );
NOR2x1_ASAP7_75t_L g25 ( .A(n_22), .B(n_12), .Y(n_25) );
OR2x2_ASAP7_75t_L g26 ( .A(n_23), .B(n_1), .Y(n_26) );
OR2x2_ASAP7_75t_L g27 ( .A(n_24), .B(n_2), .Y(n_27) );
OR2x2_ASAP7_75t_L g28 ( .A(n_25), .B(n_2), .Y(n_28) );
NOR3xp33_ASAP7_75t_L g29 ( .A(n_26), .B(n_14), .C(n_19), .Y(n_29) );
OAI21xp5_ASAP7_75t_L g30 ( .A1(n_28), .A2(n_19), .B(n_21), .Y(n_30) );
OAI321xp33_ASAP7_75t_L g31 ( .A1(n_30), .A2(n_27), .A3(n_17), .B1(n_21), .B2(n_11), .C(n_29), .Y(n_31) );
AOI211xp5_ASAP7_75t_L g32 ( .A1(n_29), .A2(n_14), .B(n_17), .C(n_5), .Y(n_32) );
BUFx6f_ASAP7_75t_L g33 ( .A(n_31), .Y(n_33) );
NAND5xp2_ASAP7_75t_L g34 ( .A(n_32), .B(n_3), .C(n_4), .D(n_5), .E(n_6), .Y(n_34) );
HB1xp67_ASAP7_75t_L g35 ( .A(n_32), .Y(n_35) );
OAI22xp5_ASAP7_75t_L g36 ( .A1(n_35), .A2(n_17), .B1(n_18), .B2(n_8), .Y(n_36) );
OAI31xp33_ASAP7_75t_SL g37 ( .A1(n_34), .A2(n_6), .A3(n_7), .B(n_8), .Y(n_37) );
AOI222xp33_ASAP7_75t_L g38 ( .A1(n_36), .A2(n_17), .B1(n_18), .B2(n_33), .C1(n_37), .C2(n_35), .Y(n_38) );
endmodule