module fake_jpeg_26120_n_326 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_326);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_326;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_4),
.B(n_5),
.Y(n_16)
);

BUFx12_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

BUFx8_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_6),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_3),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_10),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_15),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_32),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_34),
.B(n_35),
.Y(n_47)
);

CKINVDCx16_ASAP7_75t_R g35 ( 
.A(n_27),
.Y(n_35)
);

AND2x2_ASAP7_75t_L g36 ( 
.A(n_18),
.B(n_0),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_SL g54 ( 
.A(n_36),
.B(n_38),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_18),
.Y(n_37)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

OR2x2_ASAP7_75t_L g38 ( 
.A(n_32),
.B(n_0),
.Y(n_38)
);

INVx11_ASAP7_75t_L g39 ( 
.A(n_27),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

INVx2_ASAP7_75t_SL g40 ( 
.A(n_28),
.Y(n_40)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_40),
.Y(n_50)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_18),
.Y(n_41)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_41),
.Y(n_48)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_18),
.Y(n_42)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_42),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_25),
.B(n_0),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_43),
.Y(n_44)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_39),
.Y(n_45)
);

INVx1_ASAP7_75t_SL g79 ( 
.A(n_45),
.Y(n_79)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_52),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_37),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_53),
.B(n_56),
.Y(n_70)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_55),
.Y(n_71)
);

INVx1_ASAP7_75t_SL g56 ( 
.A(n_38),
.Y(n_56)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_57),
.Y(n_69)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_43),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_58),
.B(n_38),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_43),
.A2(n_25),
.B1(n_33),
.B2(n_16),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_59),
.A2(n_60),
.B1(n_31),
.B2(n_29),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_L g60 ( 
.A1(n_43),
.A2(n_25),
.B1(n_33),
.B2(n_16),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_61),
.B(n_80),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_53),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_62),
.B(n_74),
.Y(n_91)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_48),
.Y(n_63)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_63),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_44),
.B(n_38),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_64),
.B(n_66),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_45),
.A2(n_29),
.B1(n_30),
.B2(n_31),
.Y(n_65)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_65),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g66 ( 
.A(n_44),
.B(n_36),
.C(n_41),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_58),
.A2(n_40),
.B1(n_36),
.B2(n_42),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_67),
.A2(n_77),
.B1(n_85),
.B2(n_86),
.Y(n_104)
);

AO22x1_ASAP7_75t_L g72 ( 
.A1(n_56),
.A2(n_36),
.B1(n_38),
.B2(n_40),
.Y(n_72)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_72),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_54),
.B(n_38),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_73),
.B(n_35),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_59),
.B(n_30),
.Y(n_74)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_51),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_75),
.B(n_82),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_57),
.Y(n_76)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_76),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_54),
.A2(n_40),
.B1(n_36),
.B2(n_42),
.Y(n_77)
);

BUFx2_ASAP7_75t_L g78 ( 
.A(n_51),
.Y(n_78)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_78),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_47),
.B(n_20),
.Y(n_80)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_48),
.Y(n_81)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_81),
.Y(n_111)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_51),
.Y(n_82)
);

BUFx2_ASAP7_75t_L g83 ( 
.A(n_46),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_83),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_47),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_84),
.B(n_87),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_46),
.A2(n_40),
.B1(n_36),
.B2(n_42),
.Y(n_85)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_49),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_46),
.A2(n_20),
.B1(n_40),
.B2(n_21),
.Y(n_88)
);

OAI21xp33_ASAP7_75t_SL g102 ( 
.A1(n_88),
.A2(n_35),
.B(n_50),
.Y(n_102)
);

BUFx3_ASAP7_75t_L g89 ( 
.A(n_49),
.Y(n_89)
);

BUFx2_ASAP7_75t_L g99 ( 
.A(n_89),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_61),
.A2(n_40),
.B1(n_52),
.B2(n_55),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_92),
.A2(n_102),
.B1(n_105),
.B2(n_83),
.Y(n_141)
);

CKINVDCx16_ASAP7_75t_R g93 ( 
.A(n_70),
.Y(n_93)
);

CKINVDCx16_ASAP7_75t_R g142 ( 
.A(n_93),
.Y(n_142)
);

OAI22x1_ASAP7_75t_SL g94 ( 
.A1(n_72),
.A2(n_36),
.B1(n_34),
.B2(n_39),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_94),
.A2(n_118),
.B1(n_79),
.B2(n_34),
.Y(n_129)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_69),
.Y(n_95)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_95),
.Y(n_132)
);

OR2x2_ASAP7_75t_L g98 ( 
.A(n_70),
.B(n_34),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_SL g133 ( 
.A1(n_98),
.A2(n_112),
.B(n_79),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_103),
.B(n_108),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_64),
.A2(n_50),
.B1(n_39),
.B2(n_26),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_66),
.B(n_37),
.Y(n_108)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_69),
.Y(n_109)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_109),
.Y(n_136)
);

AND2x2_ASAP7_75t_SL g112 ( 
.A(n_77),
.B(n_37),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_73),
.B(n_37),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_113),
.B(n_89),
.Y(n_124)
);

CKINVDCx16_ASAP7_75t_R g115 ( 
.A(n_80),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_115),
.B(n_22),
.Y(n_131)
);

INVx2_ASAP7_75t_SL g117 ( 
.A(n_69),
.Y(n_117)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_117),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_67),
.A2(n_50),
.B1(n_20),
.B2(n_21),
.Y(n_118)
);

AOI22x1_ASAP7_75t_SL g119 ( 
.A1(n_94),
.A2(n_84),
.B1(n_72),
.B2(n_85),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_SL g161 ( 
.A1(n_119),
.A2(n_121),
.B(n_128),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_95),
.A2(n_62),
.B1(n_75),
.B2(n_82),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_120),
.A2(n_127),
.B1(n_140),
.B2(n_117),
.Y(n_150)
);

AND2x2_ASAP7_75t_L g121 ( 
.A(n_105),
.B(n_81),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_99),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_123),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_124),
.B(n_126),
.Y(n_167)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_97),
.Y(n_125)
);

BUFx24_ASAP7_75t_L g153 ( 
.A(n_125),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_90),
.B(n_87),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_109),
.A2(n_68),
.B1(n_71),
.B2(n_21),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_110),
.A2(n_68),
.B1(n_71),
.B2(n_22),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_129),
.A2(n_134),
.B1(n_112),
.B2(n_116),
.Y(n_155)
);

AND2x2_ASAP7_75t_SL g130 ( 
.A(n_107),
.B(n_92),
.Y(n_130)
);

AOI21xp5_ASAP7_75t_L g148 ( 
.A1(n_130),
.A2(n_133),
.B(n_135),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_131),
.B(n_143),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_104),
.A2(n_63),
.B1(n_83),
.B2(n_34),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_L g135 ( 
.A1(n_107),
.A2(n_22),
.B(n_26),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_SL g137 ( 
.A1(n_98),
.A2(n_26),
.B(n_27),
.Y(n_137)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_137),
.B(n_114),
.Y(n_168)
);

MAJx2_ASAP7_75t_L g139 ( 
.A(n_96),
.B(n_27),
.C(n_32),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_139),
.B(n_103),
.Y(n_156)
);

INVx4_ASAP7_75t_L g140 ( 
.A(n_99),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_141),
.A2(n_112),
.B1(n_104),
.B2(n_118),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_90),
.B(n_37),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_99),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_144),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_96),
.B(n_76),
.C(n_18),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_145),
.B(n_18),
.C(n_32),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_112),
.A2(n_24),
.B1(n_28),
.B2(n_76),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_146),
.A2(n_100),
.B1(n_111),
.B2(n_78),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_108),
.B(n_113),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_SL g159 ( 
.A(n_147),
.B(n_98),
.Y(n_159)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_124),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_149),
.B(n_158),
.Y(n_185)
);

INVxp67_ASAP7_75t_L g203 ( 
.A(n_150),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_152),
.A2(n_174),
.B1(n_123),
.B2(n_136),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_141),
.A2(n_93),
.B1(n_116),
.B2(n_115),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_154),
.A2(n_155),
.B1(n_165),
.B2(n_179),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_SL g181 ( 
.A(n_156),
.B(n_157),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g157 ( 
.A(n_139),
.B(n_147),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_146),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_SL g209 ( 
.A(n_159),
.B(n_168),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_130),
.A2(n_129),
.B1(n_134),
.B2(n_119),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_160),
.A2(n_163),
.B1(n_171),
.B2(n_177),
.Y(n_189)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_143),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_162),
.B(n_170),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_130),
.A2(n_91),
.B1(n_101),
.B2(n_106),
.Y(n_163)
);

NOR2x1_ASAP7_75t_L g164 ( 
.A(n_142),
.B(n_91),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_164),
.B(n_172),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_130),
.A2(n_117),
.B1(n_101),
.B2(n_100),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_SL g169 ( 
.A(n_122),
.B(n_15),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g202 ( 
.A(n_169),
.B(n_175),
.Y(n_202)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_133),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_119),
.A2(n_114),
.B1(n_97),
.B2(n_111),
.Y(n_171)
);

INVx3_ASAP7_75t_L g172 ( 
.A(n_140),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_122),
.B(n_32),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_176),
.B(n_139),
.C(n_145),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_121),
.A2(n_78),
.B1(n_24),
.B2(n_28),
.Y(n_177)
);

CKINVDCx16_ASAP7_75t_R g178 ( 
.A(n_128),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_178),
.B(n_131),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_142),
.A2(n_24),
.B1(n_28),
.B2(n_32),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_126),
.A2(n_24),
.B1(n_23),
.B2(n_19),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_180),
.A2(n_17),
.B1(n_23),
.B2(n_19),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_182),
.B(n_192),
.C(n_194),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_SL g183 ( 
.A1(n_148),
.A2(n_121),
.B(n_137),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_SL g231 ( 
.A1(n_183),
.A2(n_184),
.B(n_199),
.Y(n_231)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_167),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_187),
.B(n_188),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_163),
.B(n_144),
.Y(n_188)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_190),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_157),
.B(n_159),
.C(n_156),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_L g193 ( 
.A1(n_148),
.A2(n_135),
.B(n_125),
.Y(n_193)
);

AOI21xp5_ASAP7_75t_L g237 ( 
.A1(n_193),
.A2(n_212),
.B(n_1),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_175),
.B(n_136),
.C(n_132),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_167),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_195),
.B(n_201),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_170),
.B(n_132),
.C(n_138),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_197),
.B(n_210),
.C(n_17),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_173),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_198),
.Y(n_216)
);

AOI22xp33_ASAP7_75t_SL g199 ( 
.A1(n_172),
.A2(n_138),
.B1(n_27),
.B2(n_2),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_200),
.A2(n_205),
.B1(n_164),
.B2(n_166),
.Y(n_227)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_174),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_173),
.Y(n_204)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_204),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_158),
.A2(n_23),
.B1(n_19),
.B2(n_17),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_171),
.Y(n_206)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_206),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_149),
.B(n_0),
.Y(n_207)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_207),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_168),
.B(n_17),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_208),
.B(n_176),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_160),
.B(n_17),
.C(n_14),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_151),
.Y(n_211)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_211),
.Y(n_223)
);

AOI21xp5_ASAP7_75t_L g212 ( 
.A1(n_161),
.A2(n_1),
.B(n_2),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_181),
.B(n_161),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_215),
.B(n_219),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_SL g238 ( 
.A(n_218),
.B(n_228),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_181),
.B(n_169),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_192),
.B(n_155),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_221),
.B(n_226),
.Y(n_256)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_185),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_224),
.B(n_229),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_209),
.B(n_162),
.Y(n_226)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_227),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_209),
.B(n_177),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_185),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_202),
.B(n_153),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_SL g247 ( 
.A(n_232),
.B(n_234),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_L g258 ( 
.A1(n_233),
.A2(n_237),
.B(n_2),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_202),
.B(n_153),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_182),
.B(n_153),
.C(n_14),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_235),
.B(n_208),
.C(n_212),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_194),
.B(n_13),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_SL g249 ( 
.A(n_236),
.B(n_207),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_213),
.A2(n_196),
.B1(n_203),
.B2(n_189),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_240),
.B(n_241),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_230),
.B(n_197),
.C(n_193),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_242),
.B(n_243),
.C(n_245),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_230),
.B(n_221),
.C(n_234),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_225),
.Y(n_244)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_244),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_232),
.B(n_191),
.C(n_183),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_217),
.A2(n_203),
.B1(n_189),
.B2(n_206),
.Y(n_248)
);

INVxp67_ASAP7_75t_L g263 ( 
.A(n_248),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_249),
.B(n_238),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_216),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_SL g268 ( 
.A(n_250),
.B(n_252),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_220),
.A2(n_201),
.B1(n_186),
.B2(n_195),
.Y(n_251)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_251),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_SL g252 ( 
.A(n_214),
.B(n_236),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_222),
.Y(n_253)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_253),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_218),
.B(n_191),
.C(n_187),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_255),
.B(n_233),
.C(n_228),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_223),
.A2(n_190),
.B1(n_211),
.B2(n_210),
.Y(n_257)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_257),
.Y(n_271)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_258),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_SL g282 ( 
.A(n_261),
.B(n_267),
.Y(n_282)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_246),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_262),
.B(n_264),
.Y(n_279)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_248),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_SL g267 ( 
.A(n_245),
.B(n_215),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_269),
.B(n_274),
.C(n_254),
.Y(n_283)
);

OAI22x1_ASAP7_75t_L g272 ( 
.A1(n_239),
.A2(n_237),
.B1(n_231),
.B2(n_227),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_272),
.A2(n_263),
.B1(n_264),
.B2(n_271),
.Y(n_276)
);

AOI21xp33_ASAP7_75t_L g274 ( 
.A1(n_255),
.A2(n_235),
.B(n_226),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_242),
.B(n_219),
.C(n_205),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_275),
.B(n_238),
.C(n_243),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_276),
.B(n_277),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_260),
.A2(n_241),
.B1(n_249),
.B2(n_247),
.Y(n_278)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_278),
.Y(n_299)
);

AND2x2_ASAP7_75t_L g280 ( 
.A(n_272),
.B(n_256),
.Y(n_280)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_280),
.Y(n_301)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_267),
.B(n_247),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_281),
.B(n_283),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_266),
.B(n_261),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g302 ( 
.A(n_284),
.B(n_285),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_268),
.B(n_254),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_262),
.B(n_259),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_286),
.B(n_287),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_270),
.B(n_13),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_273),
.B(n_12),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_288),
.B(n_289),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_265),
.B(n_12),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_266),
.B(n_12),
.C(n_4),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_290),
.B(n_277),
.C(n_282),
.Y(n_297)
);

OAI321xp33_ASAP7_75t_L g293 ( 
.A1(n_279),
.A2(n_263),
.A3(n_275),
.B1(n_269),
.B2(n_6),
.C(n_7),
.Y(n_293)
);

XOR2xp5_ASAP7_75t_L g306 ( 
.A(n_293),
.B(n_6),
.Y(n_306)
);

HB1xp67_ASAP7_75t_L g294 ( 
.A(n_290),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_294),
.B(n_281),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_280),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_SL g304 ( 
.A(n_295),
.B(n_297),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_284),
.B(n_4),
.C(n_5),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_300),
.B(n_282),
.C(n_8),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_303),
.B(n_305),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_298),
.B(n_5),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_306),
.B(n_307),
.C(n_308),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_291),
.B(n_292),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_297),
.B(n_7),
.C(n_8),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_309),
.B(n_310),
.C(n_311),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_292),
.B(n_7),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_SL g311 ( 
.A(n_302),
.B(n_7),
.Y(n_311)
);

NOR2xp67_ASAP7_75t_L g312 ( 
.A(n_306),
.B(n_296),
.Y(n_312)
);

INVxp67_ASAP7_75t_L g319 ( 
.A(n_312),
.Y(n_319)
);

OAI21xp5_ASAP7_75t_L g316 ( 
.A1(n_304),
.A2(n_301),
.B(n_299),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_316),
.B(n_9),
.C(n_10),
.Y(n_318)
);

A2O1A1O1Ixp25_ASAP7_75t_SL g317 ( 
.A1(n_307),
.A2(n_300),
.B(n_10),
.C(n_11),
.D(n_9),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_317),
.B(n_9),
.Y(n_320)
);

OAI21xp5_ASAP7_75t_SL g321 ( 
.A1(n_318),
.A2(n_320),
.B(n_317),
.Y(n_321)
);

OAI21xp5_ASAP7_75t_SL g322 ( 
.A1(n_321),
.A2(n_319),
.B(n_315),
.Y(n_322)
);

XNOR2xp5_ASAP7_75t_L g323 ( 
.A(n_322),
.B(n_313),
.Y(n_323)
);

AOI21xp5_ASAP7_75t_L g324 ( 
.A1(n_323),
.A2(n_314),
.B(n_11),
.Y(n_324)
);

AND2x2_ASAP7_75t_L g325 ( 
.A(n_324),
.B(n_11),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_325),
.B(n_11),
.Y(n_326)
);


endmodule