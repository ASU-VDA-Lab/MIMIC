module fake_aes_9598_n_36 (n_1, n_2, n_6, n_4, n_3, n_5, n_7, n_8, n_0, n_36);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_5;
input n_7;
input n_8;
input n_0;
output n_36;
wire n_20;
wire n_34;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_30;
wire n_33;
wire n_18;
wire n_32;
wire n_35;
wire n_12;
wire n_9;
wire n_17;
wire n_14;
wire n_10;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_27;
INVx1_ASAP7_75t_L g9 ( .A(n_6), .Y(n_9) );
CKINVDCx5p33_ASAP7_75t_R g10 ( .A(n_8), .Y(n_10) );
INVx1_ASAP7_75t_L g11 ( .A(n_6), .Y(n_11) );
INVx1_ASAP7_75t_L g12 ( .A(n_0), .Y(n_12) );
BUFx2_ASAP7_75t_L g13 ( .A(n_0), .Y(n_13) );
HB1xp67_ASAP7_75t_L g14 ( .A(n_0), .Y(n_14) );
CKINVDCx20_ASAP7_75t_R g15 ( .A(n_7), .Y(n_15) );
CKINVDCx5p33_ASAP7_75t_R g16 ( .A(n_3), .Y(n_16) );
AOI21xp5_ASAP7_75t_L g17 ( .A1(n_13), .A2(n_1), .B(n_2), .Y(n_17) );
INVx1_ASAP7_75t_L g18 ( .A(n_12), .Y(n_18) );
NAND2xp5_ASAP7_75t_SL g19 ( .A(n_13), .B(n_1), .Y(n_19) );
AOI21xp5_ASAP7_75t_L g20 ( .A1(n_13), .A2(n_1), .B(n_2), .Y(n_20) );
NAND2xp5_ASAP7_75t_L g21 ( .A(n_14), .B(n_2), .Y(n_21) );
BUFx4f_ASAP7_75t_SL g22 ( .A(n_15), .Y(n_22) );
OAI22xp5_ASAP7_75t_L g23 ( .A1(n_21), .A2(n_16), .B1(n_14), .B2(n_12), .Y(n_23) );
INVxp67_ASAP7_75t_L g24 ( .A(n_21), .Y(n_24) );
NAND2xp5_ASAP7_75t_L g25 ( .A(n_18), .B(n_16), .Y(n_25) );
OR2x2_ASAP7_75t_L g26 ( .A(n_24), .B(n_19), .Y(n_26) );
NAND2xp5_ASAP7_75t_L g27 ( .A(n_25), .B(n_18), .Y(n_27) );
NAND2xp5_ASAP7_75t_L g28 ( .A(n_26), .B(n_23), .Y(n_28) );
AOI22x1_ASAP7_75t_L g29 ( .A1(n_27), .A2(n_20), .B1(n_17), .B2(n_11), .Y(n_29) );
OAI22xp5_ASAP7_75t_L g30 ( .A1(n_28), .A2(n_15), .B1(n_22), .B2(n_10), .Y(n_30) );
AOI221xp5_ASAP7_75t_L g31 ( .A1(n_29), .A2(n_11), .B1(n_9), .B2(n_4), .C(n_3), .Y(n_31) );
AOI21xp5_ASAP7_75t_L g32 ( .A1(n_31), .A2(n_29), .B(n_9), .Y(n_32) );
XOR2xp5_ASAP7_75t_L g33 ( .A(n_30), .B(n_3), .Y(n_33) );
AOI21xp5_ASAP7_75t_L g34 ( .A1(n_32), .A2(n_4), .B(n_5), .Y(n_34) );
OAI21xp5_ASAP7_75t_SL g35 ( .A1(n_33), .A2(n_4), .B(n_5), .Y(n_35) );
AOI22xp33_ASAP7_75t_SL g36 ( .A1(n_34), .A2(n_7), .B1(n_8), .B2(n_35), .Y(n_36) );
endmodule