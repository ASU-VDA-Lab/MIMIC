module fake_ibex_531_n_883 (n_151, n_147, n_85, n_167, n_128, n_84, n_64, n_3, n_73, n_152, n_171, n_145, n_65, n_103, n_95, n_139, n_55, n_130, n_63, n_98, n_129, n_161, n_29, n_143, n_106, n_148, n_2, n_76, n_8, n_118, n_67, n_9, n_164, n_38, n_124, n_37, n_110, n_47, n_169, n_108, n_10, n_82, n_21, n_27, n_165, n_16, n_78, n_60, n_86, n_70, n_7, n_20, n_87, n_69, n_75, n_109, n_121, n_127, n_175, n_137, n_48, n_57, n_59, n_28, n_125, n_39, n_5, n_62, n_71, n_153, n_173, n_120, n_93, n_168, n_155, n_162, n_13, n_122, n_116, n_61, n_14, n_0, n_94, n_134, n_12, n_42, n_77, n_112, n_150, n_88, n_133, n_44, n_142, n_51, n_46, n_80, n_172, n_49, n_40, n_66, n_17, n_74, n_90, n_176, n_58, n_43, n_140, n_22, n_136, n_4, n_119, n_33, n_30, n_6, n_100, n_72, n_166, n_163, n_26, n_114, n_34, n_97, n_102, n_15, n_131, n_123, n_24, n_52, n_99, n_135, n_105, n_156, n_126, n_1, n_154, n_111, n_25, n_36, n_104, n_41, n_45, n_141, n_18, n_89, n_83, n_32, n_53, n_107, n_115, n_149, n_50, n_11, n_92, n_144, n_170, n_101, n_113, n_138, n_96, n_68, n_117, n_79, n_81, n_35, n_159, n_158, n_132, n_174, n_157, n_160, n_31, n_56, n_23, n_146, n_91, n_54, n_19, n_883);

input n_151;
input n_147;
input n_85;
input n_167;
input n_128;
input n_84;
input n_64;
input n_3;
input n_73;
input n_152;
input n_171;
input n_145;
input n_65;
input n_103;
input n_95;
input n_139;
input n_55;
input n_130;
input n_63;
input n_98;
input n_129;
input n_161;
input n_29;
input n_143;
input n_106;
input n_148;
input n_2;
input n_76;
input n_8;
input n_118;
input n_67;
input n_9;
input n_164;
input n_38;
input n_124;
input n_37;
input n_110;
input n_47;
input n_169;
input n_108;
input n_10;
input n_82;
input n_21;
input n_27;
input n_165;
input n_16;
input n_78;
input n_60;
input n_86;
input n_70;
input n_7;
input n_20;
input n_87;
input n_69;
input n_75;
input n_109;
input n_121;
input n_127;
input n_175;
input n_137;
input n_48;
input n_57;
input n_59;
input n_28;
input n_125;
input n_39;
input n_5;
input n_62;
input n_71;
input n_153;
input n_173;
input n_120;
input n_93;
input n_168;
input n_155;
input n_162;
input n_13;
input n_122;
input n_116;
input n_61;
input n_14;
input n_0;
input n_94;
input n_134;
input n_12;
input n_42;
input n_77;
input n_112;
input n_150;
input n_88;
input n_133;
input n_44;
input n_142;
input n_51;
input n_46;
input n_80;
input n_172;
input n_49;
input n_40;
input n_66;
input n_17;
input n_74;
input n_90;
input n_176;
input n_58;
input n_43;
input n_140;
input n_22;
input n_136;
input n_4;
input n_119;
input n_33;
input n_30;
input n_6;
input n_100;
input n_72;
input n_166;
input n_163;
input n_26;
input n_114;
input n_34;
input n_97;
input n_102;
input n_15;
input n_131;
input n_123;
input n_24;
input n_52;
input n_99;
input n_135;
input n_105;
input n_156;
input n_126;
input n_1;
input n_154;
input n_111;
input n_25;
input n_36;
input n_104;
input n_41;
input n_45;
input n_141;
input n_18;
input n_89;
input n_83;
input n_32;
input n_53;
input n_107;
input n_115;
input n_149;
input n_50;
input n_11;
input n_92;
input n_144;
input n_170;
input n_101;
input n_113;
input n_138;
input n_96;
input n_68;
input n_117;
input n_79;
input n_81;
input n_35;
input n_159;
input n_158;
input n_132;
input n_174;
input n_157;
input n_160;
input n_31;
input n_56;
input n_23;
input n_146;
input n_91;
input n_54;
input n_19;

output n_883;

wire n_599;
wire n_778;
wire n_822;
wire n_507;
wire n_743;
wire n_540;
wire n_754;
wire n_395;
wire n_756;
wire n_529;
wire n_389;
wire n_204;
wire n_626;
wire n_274;
wire n_387;
wire n_766;
wire n_688;
wire n_177;
wire n_707;
wire n_273;
wire n_330;
wire n_309;
wire n_328;
wire n_293;
wire n_341;
wire n_372;
wire n_418;
wire n_256;
wire n_510;
wire n_193;
wire n_845;
wire n_446;
wire n_350;
wire n_601;
wire n_621;
wire n_610;
wire n_790;
wire n_452;
wire n_664;
wire n_255;
wire n_586;
wire n_773;
wire n_638;
wire n_398;
wire n_304;
wire n_821;
wire n_191;
wire n_873;
wire n_593;
wire n_862;
wire n_545;
wire n_583;
wire n_678;
wire n_663;
wire n_194;
wire n_249;
wire n_334;
wire n_634;
wire n_733;
wire n_312;
wire n_622;
wire n_578;
wire n_478;
wire n_239;
wire n_432;
wire n_371;
wire n_403;
wire n_872;
wire n_423;
wire n_608;
wire n_864;
wire n_357;
wire n_412;
wire n_457;
wire n_494;
wire n_226;
wire n_336;
wire n_258;
wire n_861;
wire n_449;
wire n_547;
wire n_727;
wire n_216;
wire n_652;
wire n_781;
wire n_421;
wire n_828;
wire n_738;
wire n_475;
wire n_802;
wire n_753;
wire n_645;
wire n_500;
wire n_747;
wire n_542;
wire n_236;
wire n_376;
wire n_377;
wire n_584;
wire n_531;
wire n_647;
wire n_761;
wire n_556;
wire n_748;
wire n_189;
wire n_498;
wire n_708;
wire n_280;
wire n_375;
wire n_340;
wire n_317;
wire n_698;
wire n_187;
wire n_667;
wire n_682;
wire n_850;
wire n_182;
wire n_196;
wire n_327;
wire n_326;
wire n_879;
wire n_723;
wire n_270;
wire n_346;
wire n_383;
wire n_840;
wire n_561;
wire n_417;
wire n_471;
wire n_846;
wire n_739;
wire n_755;
wire n_265;
wire n_853;
wire n_504;
wire n_859;
wire n_259;
wire n_339;
wire n_276;
wire n_470;
wire n_770;
wire n_210;
wire n_348;
wire n_220;
wire n_875;
wire n_674;
wire n_481;
wire n_287;
wire n_243;
wire n_497;
wire n_671;
wire n_228;
wire n_711;
wire n_876;
wire n_552;
wire n_251;
wire n_384;
wire n_632;
wire n_373;
wire n_854;
wire n_458;
wire n_244;
wire n_343;
wire n_310;
wire n_714;
wire n_703;
wire n_426;
wire n_323;
wire n_469;
wire n_829;
wire n_598;
wire n_825;
wire n_740;
wire n_386;
wire n_549;
wire n_224;
wire n_183;
wire n_533;
wire n_508;
wire n_453;
wire n_591;
wire n_655;
wire n_333;
wire n_306;
wire n_400;
wire n_550;
wire n_736;
wire n_673;
wire n_798;
wire n_832;
wire n_732;
wire n_242;
wire n_278;
wire n_316;
wire n_404;
wire n_557;
wire n_641;
wire n_527;
wire n_590;
wire n_465;
wire n_325;
wire n_301;
wire n_496;
wire n_617;
wire n_434;
wire n_296;
wire n_690;
wire n_835;
wire n_526;
wire n_785;
wire n_824;
wire n_315;
wire n_441;
wire n_604;
wire n_637;
wire n_523;
wire n_694;
wire n_787;
wire n_614;
wire n_370;
wire n_431;
wire n_719;
wire n_574;
wire n_289;
wire n_716;
wire n_865;
wire n_515;
wire n_642;
wire n_286;
wire n_321;
wire n_569;
wire n_600;
wire n_215;
wire n_279;
wire n_374;
wire n_235;
wire n_464;
wire n_538;
wire n_669;
wire n_838;
wire n_750;
wire n_746;
wire n_261;
wire n_742;
wire n_521;
wire n_665;
wire n_459;
wire n_518;
wire n_367;
wire n_221;
wire n_852;
wire n_789;
wire n_880;
wire n_654;
wire n_656;
wire n_724;
wire n_437;
wire n_731;
wire n_602;
wire n_842;
wire n_355;
wire n_767;
wire n_474;
wire n_878;
wire n_758;
wire n_636;
wire n_594;
wire n_710;
wire n_720;
wire n_407;
wire n_490;
wire n_568;
wire n_813;
wire n_448;
wire n_646;
wire n_595;
wire n_466;
wire n_269;
wire n_570;
wire n_623;
wire n_585;
wire n_715;
wire n_791;
wire n_530;
wire n_356;
wire n_420;
wire n_483;
wire n_543;
wire n_580;
wire n_487;
wire n_769;
wire n_222;
wire n_660;
wire n_186;
wire n_524;
wire n_349;
wire n_765;
wire n_849;
wire n_857;
wire n_454;
wire n_777;
wire n_295;
wire n_730;
wire n_331;
wire n_576;
wire n_230;
wire n_759;
wire n_185;
wire n_388;
wire n_625;
wire n_619;
wire n_536;
wire n_611;
wire n_352;
wire n_290;
wire n_558;
wire n_666;
wire n_467;
wire n_427;
wire n_607;
wire n_827;
wire n_219;
wire n_246;
wire n_442;
wire n_207;
wire n_438;
wire n_851;
wire n_689;
wire n_793;
wire n_676;
wire n_253;
wire n_208;
wire n_234;
wire n_300;
wire n_358;
wire n_771;
wire n_205;
wire n_618;
wire n_488;
wire n_514;
wire n_705;
wire n_429;
wire n_560;
wire n_275;
wire n_541;
wire n_613;
wire n_659;
wire n_267;
wire n_662;
wire n_635;
wire n_844;
wire n_245;
wire n_648;
wire n_571;
wire n_229;
wire n_209;
wire n_472;
wire n_589;
wire n_783;
wire n_347;
wire n_847;
wire n_830;
wire n_473;
wire n_445;
wire n_629;
wire n_335;
wire n_413;
wire n_263;
wire n_573;
wire n_353;
wire n_359;
wire n_826;
wire n_299;
wire n_262;
wire n_433;
wire n_439;
wire n_704;
wire n_643;
wire n_679;
wire n_841;
wire n_772;
wire n_810;
wire n_839;
wire n_768;
wire n_338;
wire n_696;
wire n_837;
wire n_797;
wire n_796;
wire n_477;
wire n_640;
wire n_363;
wire n_402;
wire n_725;
wire n_180;
wire n_369;
wire n_596;
wire n_201;
wire n_699;
wire n_351;
wire n_368;
wire n_456;
wire n_834;
wire n_257;
wire n_869;
wire n_718;
wire n_801;
wire n_672;
wire n_722;
wire n_401;
wire n_553;
wire n_554;
wire n_735;
wire n_305;
wire n_882;
wire n_713;
wire n_307;
wire n_192;
wire n_804;
wire n_484;
wire n_566;
wire n_480;
wire n_416;
wire n_581;
wire n_651;
wire n_365;
wire n_721;
wire n_814;
wire n_605;
wire n_539;
wire n_179;
wire n_354;
wire n_392;
wire n_206;
wire n_630;
wire n_567;
wire n_548;
wire n_516;
wire n_763;
wire n_745;
wire n_329;
wire n_447;
wire n_188;
wire n_200;
wire n_444;
wire n_506;
wire n_562;
wire n_564;
wire n_868;
wire n_546;
wire n_199;
wire n_788;
wire n_795;
wire n_592;
wire n_495;
wire n_762;
wire n_410;
wire n_308;
wire n_675;
wire n_800;
wire n_463;
wire n_624;
wire n_706;
wire n_411;
wire n_520;
wire n_784;
wire n_684;
wire n_775;
wire n_658;
wire n_512;
wire n_615;
wire n_685;
wire n_283;
wire n_366;
wire n_397;
wire n_803;
wire n_692;
wire n_627;
wire n_709;
wire n_322;
wire n_227;
wire n_499;
wire n_757;
wire n_248;
wire n_702;
wire n_451;
wire n_712;
wire n_190;
wire n_650;
wire n_776;
wire n_409;
wire n_582;
wire n_818;
wire n_653;
wire n_238;
wire n_214;
wire n_579;
wire n_843;
wire n_332;
wire n_799;
wire n_517;
wire n_211;
wire n_744;
wire n_817;
wire n_218;
wire n_314;
wire n_691;
wire n_563;
wire n_277;
wire n_555;
wire n_337;
wire n_522;
wire n_700;
wire n_479;
wire n_534;
wire n_225;
wire n_360;
wire n_881;
wire n_272;
wire n_511;
wire n_734;
wire n_468;
wire n_223;
wire n_381;
wire n_525;
wire n_815;
wire n_780;
wire n_535;
wire n_382;
wire n_502;
wire n_681;
wire n_633;
wire n_532;
wire n_726;
wire n_405;
wire n_863;
wire n_415;
wire n_597;
wire n_288;
wire n_320;
wire n_247;
wire n_285;
wire n_379;
wire n_551;
wire n_612;
wire n_318;
wire n_291;
wire n_819;
wire n_237;
wire n_203;
wire n_268;
wire n_440;
wire n_858;
wire n_342;
wire n_233;
wire n_414;
wire n_385;
wire n_430;
wire n_729;
wire n_741;
wire n_603;
wire n_378;
wire n_486;
wire n_422;
wire n_264;
wire n_198;
wire n_616;
wire n_782;
wire n_833;
wire n_217;
wire n_324;
wire n_391;
wire n_831;
wire n_537;
wire n_728;
wire n_805;
wire n_670;
wire n_820;
wire n_390;
wire n_544;
wire n_178;
wire n_509;
wire n_695;
wire n_786;
wire n_639;
wire n_303;
wire n_362;
wire n_717;
wire n_505;
wire n_482;
wire n_240;
wire n_282;
wire n_680;
wire n_501;
wire n_809;
wire n_752;
wire n_856;
wire n_668;
wire n_779;
wire n_871;
wire n_266;
wire n_294;
wire n_485;
wire n_870;
wire n_284;
wire n_811;
wire n_808;
wire n_250;
wire n_493;
wire n_460;
wire n_609;
wire n_476;
wire n_792;
wire n_461;
wire n_575;
wire n_313;
wire n_519;
wire n_345;
wire n_408;
wire n_361;
wire n_455;
wire n_419;
wire n_774;
wire n_319;
wire n_195;
wire n_513;
wire n_212;
wire n_588;
wire n_877;
wire n_693;
wire n_311;
wire n_860;
wire n_661;
wire n_848;
wire n_406;
wire n_606;
wire n_737;
wire n_197;
wire n_528;
wire n_181;
wire n_631;
wire n_683;
wire n_260;
wire n_620;
wire n_794;
wire n_836;
wire n_462;
wire n_302;
wire n_450;
wire n_443;
wire n_686;
wire n_572;
wire n_867;
wire n_644;
wire n_577;
wire n_344;
wire n_393;
wire n_436;
wire n_428;
wire n_491;
wire n_297;
wire n_435;
wire n_628;
wire n_252;
wire n_396;
wire n_697;
wire n_816;
wire n_874;
wire n_489;
wire n_677;
wire n_399;
wire n_254;
wire n_213;
wire n_424;
wire n_565;
wire n_823;
wire n_701;
wire n_271;
wire n_241;
wire n_503;
wire n_292;
wire n_807;
wire n_394;
wire n_364;
wire n_687;
wire n_231;
wire n_202;
wire n_298;
wire n_587;
wire n_760;
wire n_751;
wire n_806;
wire n_657;
wire n_764;
wire n_184;
wire n_492;
wire n_649;
wire n_812;
wire n_855;
wire n_232;
wire n_380;
wire n_749;
wire n_281;
wire n_866;
wire n_559;
wire n_425;

INVx1_ASAP7_75t_SL g177 ( 
.A(n_155),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_0),
.Y(n_178)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_5),
.Y(n_179)
);

INVxp67_ASAP7_75t_SL g180 ( 
.A(n_114),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g181 ( 
.A(n_48),
.Y(n_181)
);

BUFx3_ASAP7_75t_L g182 ( 
.A(n_80),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_78),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_150),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_176),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_60),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_130),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_159),
.Y(n_188)
);

BUFx6f_ASAP7_75t_L g189 ( 
.A(n_112),
.Y(n_189)
);

INVxp67_ASAP7_75t_SL g190 ( 
.A(n_39),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_131),
.Y(n_191)
);

OR2x2_ASAP7_75t_L g192 ( 
.A(n_77),
.B(n_41),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_26),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_123),
.B(n_113),
.Y(n_194)
);

BUFx2_ASAP7_75t_L g195 ( 
.A(n_13),
.Y(n_195)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_55),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_29),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_14),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_103),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_71),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_53),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_156),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_29),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_162),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_146),
.B(n_49),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_70),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_81),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_128),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_20),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_62),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_139),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_153),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_167),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_65),
.Y(n_214)
);

CKINVDCx14_ASAP7_75t_R g215 ( 
.A(n_69),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_38),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_17),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_14),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_120),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_91),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_88),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_86),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_141),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_1),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_42),
.B(n_32),
.Y(n_225)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_54),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_72),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_106),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_33),
.Y(n_229)
);

INVx1_ASAP7_75t_SL g230 ( 
.A(n_26),
.Y(n_230)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_107),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_169),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_63),
.Y(n_233)
);

INVxp67_ASAP7_75t_L g234 ( 
.A(n_74),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_94),
.Y(n_235)
);

BUFx10_ASAP7_75t_L g236 ( 
.A(n_96),
.Y(n_236)
);

BUFx2_ASAP7_75t_L g237 ( 
.A(n_24),
.Y(n_237)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_35),
.Y(n_238)
);

BUFx2_ASAP7_75t_L g239 ( 
.A(n_68),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_61),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_15),
.Y(n_241)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_23),
.Y(n_242)
);

BUFx3_ASAP7_75t_L g243 ( 
.A(n_67),
.Y(n_243)
);

BUFx3_ASAP7_75t_L g244 ( 
.A(n_87),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_143),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_163),
.Y(n_246)
);

INVxp67_ASAP7_75t_L g247 ( 
.A(n_95),
.Y(n_247)
);

CKINVDCx14_ASAP7_75t_R g248 ( 
.A(n_101),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_73),
.Y(n_249)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_79),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_51),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_37),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_82),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_36),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_158),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_66),
.Y(n_256)
);

BUFx6f_ASAP7_75t_L g257 ( 
.A(n_110),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_52),
.Y(n_258)
);

CKINVDCx16_ASAP7_75t_R g259 ( 
.A(n_46),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_116),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_157),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_102),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_122),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_142),
.Y(n_264)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_36),
.Y(n_265)
);

BUFx6f_ASAP7_75t_L g266 ( 
.A(n_127),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_40),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_7),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_168),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_64),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_30),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_85),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_140),
.Y(n_273)
);

INVx1_ASAP7_75t_SL g274 ( 
.A(n_93),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_121),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_149),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_1),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_105),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_108),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_31),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_160),
.Y(n_281)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_98),
.Y(n_282)
);

BUFx10_ASAP7_75t_L g283 ( 
.A(n_148),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_59),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_144),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_18),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_6),
.Y(n_287)
);

BUFx5_ASAP7_75t_L g288 ( 
.A(n_58),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_50),
.Y(n_289)
);

BUFx5_ASAP7_75t_L g290 ( 
.A(n_90),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_75),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_76),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_195),
.B(n_0),
.Y(n_293)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_288),
.Y(n_294)
);

BUFx6f_ASAP7_75t_L g295 ( 
.A(n_181),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_239),
.Y(n_296)
);

AND2x4_ASAP7_75t_L g297 ( 
.A(n_179),
.B(n_2),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_225),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_179),
.Y(n_299)
);

INVx6_ASAP7_75t_L g300 ( 
.A(n_236),
.Y(n_300)
);

NOR2x1_ASAP7_75t_L g301 ( 
.A(n_265),
.B(n_43),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_237),
.B(n_3),
.Y(n_302)
);

OAI21x1_ASAP7_75t_L g303 ( 
.A1(n_196),
.A2(n_84),
.B(n_174),
.Y(n_303)
);

OA21x2_ASAP7_75t_L g304 ( 
.A1(n_196),
.A2(n_83),
.B(n_173),
.Y(n_304)
);

BUFx6f_ASAP7_75t_L g305 ( 
.A(n_181),
.Y(n_305)
);

AND2x2_ASAP7_75t_L g306 ( 
.A(n_259),
.B(n_4),
.Y(n_306)
);

INVx6_ASAP7_75t_L g307 ( 
.A(n_236),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_238),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_234),
.B(n_5),
.Y(n_309)
);

AND2x4_ASAP7_75t_L g310 ( 
.A(n_242),
.B(n_6),
.Y(n_310)
);

BUFx6f_ASAP7_75t_L g311 ( 
.A(n_181),
.Y(n_311)
);

HB1xp67_ASAP7_75t_L g312 ( 
.A(n_178),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_247),
.B(n_7),
.Y(n_313)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_288),
.Y(n_314)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_288),
.Y(n_315)
);

INVx3_ASAP7_75t_L g316 ( 
.A(n_283),
.Y(n_316)
);

BUFx6f_ASAP7_75t_L g317 ( 
.A(n_181),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_193),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_318)
);

AND2x2_ASAP7_75t_L g319 ( 
.A(n_215),
.B(n_8),
.Y(n_319)
);

BUFx2_ASAP7_75t_L g320 ( 
.A(n_197),
.Y(n_320)
);

AND2x2_ASAP7_75t_L g321 ( 
.A(n_215),
.B(n_10),
.Y(n_321)
);

INVx2_ASAP7_75t_SL g322 ( 
.A(n_283),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_217),
.Y(n_323)
);

BUFx12f_ASAP7_75t_L g324 ( 
.A(n_186),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_SL g325 ( 
.A1(n_198),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_325)
);

BUFx6f_ASAP7_75t_L g326 ( 
.A(n_189),
.Y(n_326)
);

BUFx6f_ASAP7_75t_L g327 ( 
.A(n_189),
.Y(n_327)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_288),
.Y(n_328)
);

INVx3_ASAP7_75t_L g329 ( 
.A(n_218),
.Y(n_329)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_288),
.Y(n_330)
);

BUFx8_ASAP7_75t_L g331 ( 
.A(n_290),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_282),
.B(n_11),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_224),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_268),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_277),
.B(n_12),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_226),
.B(n_15),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_280),
.Y(n_337)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_290),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_286),
.Y(n_339)
);

AOI22x1_ASAP7_75t_SL g340 ( 
.A1(n_203),
.A2(n_16),
.B1(n_17),
.B2(n_19),
.Y(n_340)
);

INVx3_ASAP7_75t_L g341 ( 
.A(n_226),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_SL g342 ( 
.A(n_290),
.B(n_16),
.Y(n_342)
);

AND2x2_ASAP7_75t_L g343 ( 
.A(n_248),
.B(n_19),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_183),
.Y(n_344)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_290),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_184),
.Y(n_346)
);

BUFx6f_ASAP7_75t_L g347 ( 
.A(n_189),
.Y(n_347)
);

INVx2_ASAP7_75t_L g348 ( 
.A(n_290),
.Y(n_348)
);

AOI22xp5_ASAP7_75t_L g349 ( 
.A1(n_248),
.A2(n_20),
.B1(n_21),
.B2(n_22),
.Y(n_349)
);

INVx2_ASAP7_75t_L g350 ( 
.A(n_231),
.Y(n_350)
);

INVx2_ASAP7_75t_SL g351 ( 
.A(n_182),
.Y(n_351)
);

BUFx12f_ASAP7_75t_L g352 ( 
.A(n_187),
.Y(n_352)
);

INVx3_ASAP7_75t_L g353 ( 
.A(n_231),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_199),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g355 ( 
.A(n_240),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_250),
.B(n_21),
.Y(n_356)
);

NOR2x1_ASAP7_75t_L g357 ( 
.A(n_185),
.B(n_188),
.Y(n_357)
);

AOI22xp5_ASAP7_75t_L g358 ( 
.A1(n_209),
.A2(n_22),
.B1(n_24),
.B2(n_25),
.Y(n_358)
);

INVx2_ASAP7_75t_L g359 ( 
.A(n_250),
.Y(n_359)
);

AND2x4_ASAP7_75t_L g360 ( 
.A(n_243),
.B(n_25),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_191),
.B(n_27),
.Y(n_361)
);

NAND2xp33_ASAP7_75t_R g362 ( 
.A(n_306),
.B(n_216),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_297),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_L g364 ( 
.A(n_316),
.B(n_201),
.Y(n_364)
);

INVx2_ASAP7_75t_L g365 ( 
.A(n_294),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_L g366 ( 
.A(n_316),
.B(n_202),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_297),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_297),
.Y(n_368)
);

HB1xp67_ASAP7_75t_L g369 ( 
.A(n_321),
.Y(n_369)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_294),
.Y(n_370)
);

AND2x6_ASAP7_75t_L g371 ( 
.A(n_360),
.B(n_244),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_310),
.Y(n_372)
);

BUFx3_ASAP7_75t_L g373 ( 
.A(n_331),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_SL g374 ( 
.A(n_331),
.B(n_204),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_310),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_316),
.B(n_229),
.Y(n_376)
);

NAND2xp33_ASAP7_75t_L g377 ( 
.A(n_319),
.B(n_292),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_296),
.B(n_241),
.Y(n_378)
);

INVx2_ASAP7_75t_L g379 ( 
.A(n_314),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_310),
.Y(n_380)
);

INVx4_ASAP7_75t_L g381 ( 
.A(n_360),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_329),
.Y(n_382)
);

INVx2_ASAP7_75t_L g383 ( 
.A(n_314),
.Y(n_383)
);

AND2x2_ASAP7_75t_L g384 ( 
.A(n_320),
.B(n_252),
.Y(n_384)
);

INVx2_ASAP7_75t_L g385 ( 
.A(n_315),
.Y(n_385)
);

AND3x2_ASAP7_75t_L g386 ( 
.A(n_343),
.B(n_190),
.C(n_180),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_344),
.B(n_346),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_354),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_341),
.Y(n_389)
);

AND3x2_ASAP7_75t_L g390 ( 
.A(n_312),
.B(n_190),
.C(n_180),
.Y(n_390)
);

OAI22xp33_ASAP7_75t_L g391 ( 
.A1(n_349),
.A2(n_230),
.B1(n_254),
.B2(n_287),
.Y(n_391)
);

NOR2xp33_ASAP7_75t_L g392 ( 
.A(n_300),
.B(n_207),
.Y(n_392)
);

CKINVDCx14_ASAP7_75t_R g393 ( 
.A(n_300),
.Y(n_393)
);

AND2x6_ASAP7_75t_L g394 ( 
.A(n_301),
.B(n_244),
.Y(n_394)
);

AND2x2_ASAP7_75t_L g395 ( 
.A(n_300),
.B(n_271),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_353),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_SL g397 ( 
.A(n_315),
.B(n_208),
.Y(n_397)
);

INVx2_ASAP7_75t_L g398 ( 
.A(n_328),
.Y(n_398)
);

AOI22xp33_ASAP7_75t_L g399 ( 
.A1(n_350),
.A2(n_245),
.B1(n_246),
.B2(n_235),
.Y(n_399)
);

AND3x2_ASAP7_75t_L g400 ( 
.A(n_340),
.B(n_205),
.C(n_210),
.Y(n_400)
);

AOI22xp33_ASAP7_75t_L g401 ( 
.A1(n_350),
.A2(n_359),
.B1(n_323),
.B2(n_333),
.Y(n_401)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_328),
.Y(n_402)
);

BUFx2_ASAP7_75t_L g403 ( 
.A(n_324),
.Y(n_403)
);

AOI21x1_ASAP7_75t_L g404 ( 
.A1(n_303),
.A2(n_213),
.B(n_212),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_359),
.Y(n_405)
);

AND2x2_ASAP7_75t_L g406 ( 
.A(n_307),
.B(n_200),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_351),
.Y(n_407)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_330),
.Y(n_408)
);

INVx3_ASAP7_75t_L g409 ( 
.A(n_330),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_SL g410 ( 
.A(n_338),
.B(n_219),
.Y(n_410)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_338),
.Y(n_411)
);

BUFx6f_ASAP7_75t_SL g412 ( 
.A(n_322),
.Y(n_412)
);

BUFx10_ASAP7_75t_L g413 ( 
.A(n_322),
.Y(n_413)
);

NAND3xp33_ASAP7_75t_L g414 ( 
.A(n_293),
.B(n_302),
.C(n_357),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_334),
.Y(n_415)
);

BUFx2_ASAP7_75t_L g416 ( 
.A(n_324),
.Y(n_416)
);

OR2x6_ASAP7_75t_L g417 ( 
.A(n_298),
.B(n_194),
.Y(n_417)
);

AND2x4_ASAP7_75t_L g418 ( 
.A(n_337),
.B(n_220),
.Y(n_418)
);

INVx2_ASAP7_75t_SL g419 ( 
.A(n_352),
.Y(n_419)
);

HB1xp67_ASAP7_75t_L g420 ( 
.A(n_356),
.Y(n_420)
);

NAND3xp33_ASAP7_75t_L g421 ( 
.A(n_309),
.B(n_232),
.C(n_227),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_339),
.B(n_206),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_299),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_308),
.Y(n_424)
);

INVx2_ASAP7_75t_L g425 ( 
.A(n_345),
.Y(n_425)
);

INVx2_ASAP7_75t_L g426 ( 
.A(n_345),
.Y(n_426)
);

AOI22xp33_ASAP7_75t_L g427 ( 
.A1(n_342),
.A2(n_272),
.B1(n_262),
.B2(n_263),
.Y(n_427)
);

INVx2_ASAP7_75t_L g428 ( 
.A(n_348),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_354),
.Y(n_429)
);

INVx2_ASAP7_75t_L g430 ( 
.A(n_348),
.Y(n_430)
);

NAND2xp33_ASAP7_75t_SL g431 ( 
.A(n_361),
.B(n_267),
.Y(n_431)
);

OR2x6_ASAP7_75t_L g432 ( 
.A(n_325),
.B(n_194),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_335),
.Y(n_433)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_295),
.Y(n_434)
);

AOI22xp5_ASAP7_75t_L g435 ( 
.A1(n_309),
.A2(n_261),
.B1(n_255),
.B2(n_256),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_SL g436 ( 
.A(n_332),
.B(n_258),
.Y(n_436)
);

NAND2xp33_ASAP7_75t_R g437 ( 
.A(n_304),
.B(n_211),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_336),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_SL g439 ( 
.A(n_313),
.B(n_264),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_313),
.B(n_214),
.Y(n_440)
);

INVx2_ASAP7_75t_L g441 ( 
.A(n_295),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_304),
.Y(n_442)
);

NAND2xp33_ASAP7_75t_SL g443 ( 
.A(n_355),
.B(n_192),
.Y(n_443)
);

HB1xp67_ASAP7_75t_L g444 ( 
.A(n_352),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_382),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_433),
.B(n_418),
.Y(n_446)
);

NOR2xp67_ASAP7_75t_SL g447 ( 
.A(n_373),
.B(n_221),
.Y(n_447)
);

NOR2x1p5_ASAP7_75t_L g448 ( 
.A(n_388),
.B(n_355),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_SL g449 ( 
.A(n_373),
.B(n_222),
.Y(n_449)
);

INVx2_ASAP7_75t_L g450 ( 
.A(n_409),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_418),
.B(n_223),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_369),
.B(n_228),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_369),
.B(n_233),
.Y(n_453)
);

INVxp67_ASAP7_75t_SL g454 ( 
.A(n_363),
.Y(n_454)
);

NAND2x1_ASAP7_75t_L g455 ( 
.A(n_381),
.B(n_304),
.Y(n_455)
);

AND2x2_ASAP7_75t_L g456 ( 
.A(n_393),
.B(n_318),
.Y(n_456)
);

NOR2xp33_ASAP7_75t_L g457 ( 
.A(n_376),
.B(n_269),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_415),
.B(n_249),
.Y(n_458)
);

BUFx4f_ASAP7_75t_L g459 ( 
.A(n_419),
.Y(n_459)
);

OAI22xp33_ASAP7_75t_L g460 ( 
.A1(n_417),
.A2(n_358),
.B1(n_276),
.B2(n_275),
.Y(n_460)
);

NOR2xp33_ASAP7_75t_R g461 ( 
.A(n_393),
.B(n_251),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_422),
.B(n_253),
.Y(n_462)
);

NOR2xp33_ASAP7_75t_L g463 ( 
.A(n_414),
.B(n_270),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_387),
.B(n_260),
.Y(n_464)
);

NOR2xp33_ASAP7_75t_L g465 ( 
.A(n_440),
.B(n_273),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_407),
.Y(n_466)
);

NOR2xp67_ASAP7_75t_L g467 ( 
.A(n_444),
.B(n_421),
.Y(n_467)
);

CKINVDCx11_ASAP7_75t_R g468 ( 
.A(n_403),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_438),
.B(n_278),
.Y(n_469)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_423),
.Y(n_470)
);

INVx2_ASAP7_75t_L g471 ( 
.A(n_424),
.Y(n_471)
);

AND2x2_ASAP7_75t_L g472 ( 
.A(n_384),
.B(n_395),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_364),
.B(n_285),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_SL g474 ( 
.A(n_374),
.B(n_289),
.Y(n_474)
);

NOR2xp33_ASAP7_75t_L g475 ( 
.A(n_439),
.B(n_279),
.Y(n_475)
);

INVx2_ASAP7_75t_SL g476 ( 
.A(n_413),
.Y(n_476)
);

NOR2xp33_ASAP7_75t_L g477 ( 
.A(n_439),
.B(n_281),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_364),
.B(n_291),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_366),
.B(n_177),
.Y(n_479)
);

AOI22xp33_ASAP7_75t_L g480 ( 
.A1(n_367),
.A2(n_284),
.B1(n_189),
.B2(n_257),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_366),
.B(n_274),
.Y(n_481)
);

AOI22xp5_ASAP7_75t_L g482 ( 
.A1(n_431),
.A2(n_205),
.B1(n_257),
.B2(n_266),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_405),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_389),
.Y(n_484)
);

OR2x6_ASAP7_75t_L g485 ( 
.A(n_416),
.B(n_266),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_SL g486 ( 
.A(n_365),
.B(n_266),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_436),
.B(n_392),
.Y(n_487)
);

HB1xp67_ASAP7_75t_L g488 ( 
.A(n_362),
.Y(n_488)
);

AOI22xp33_ASAP7_75t_L g489 ( 
.A1(n_368),
.A2(n_347),
.B1(n_327),
.B2(n_326),
.Y(n_489)
);

AND2x2_ASAP7_75t_L g490 ( 
.A(n_406),
.B(n_28),
.Y(n_490)
);

INVxp67_ASAP7_75t_L g491 ( 
.A(n_362),
.Y(n_491)
);

OR2x6_ASAP7_75t_L g492 ( 
.A(n_417),
.B(n_305),
.Y(n_492)
);

INVx3_ASAP7_75t_L g493 ( 
.A(n_396),
.Y(n_493)
);

NOR2xp33_ASAP7_75t_SL g494 ( 
.A(n_429),
.B(n_347),
.Y(n_494)
);

AOI22xp33_ASAP7_75t_L g495 ( 
.A1(n_372),
.A2(n_380),
.B1(n_375),
.B2(n_371),
.Y(n_495)
);

O2A1O1Ixp33_ASAP7_75t_L g496 ( 
.A1(n_391),
.A2(n_28),
.B(n_30),
.C(n_31),
.Y(n_496)
);

INVxp67_ASAP7_75t_SL g497 ( 
.A(n_401),
.Y(n_497)
);

AND2x4_ASAP7_75t_L g498 ( 
.A(n_386),
.B(n_32),
.Y(n_498)
);

AOI22xp33_ASAP7_75t_L g499 ( 
.A1(n_371),
.A2(n_347),
.B1(n_327),
.B2(n_326),
.Y(n_499)
);

OAI22xp5_ASAP7_75t_L g500 ( 
.A1(n_378),
.A2(n_347),
.B1(n_327),
.B2(n_326),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_397),
.Y(n_501)
);

NOR2xp33_ASAP7_75t_SL g502 ( 
.A(n_412),
.B(n_327),
.Y(n_502)
);

NOR2xp33_ASAP7_75t_L g503 ( 
.A(n_435),
.B(n_311),
.Y(n_503)
);

BUFx6f_ASAP7_75t_L g504 ( 
.A(n_404),
.Y(n_504)
);

INVx2_ASAP7_75t_SL g505 ( 
.A(n_390),
.Y(n_505)
);

AND2x2_ASAP7_75t_L g506 ( 
.A(n_401),
.B(n_33),
.Y(n_506)
);

OAI22xp33_ASAP7_75t_L g507 ( 
.A1(n_417),
.A2(n_326),
.B1(n_317),
.B2(n_37),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_397),
.Y(n_508)
);

OR2x6_ASAP7_75t_L g509 ( 
.A(n_432),
.B(n_317),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_399),
.B(n_34),
.Y(n_510)
);

AND3x1_ASAP7_75t_L g511 ( 
.A(n_400),
.B(n_34),
.C(n_35),
.Y(n_511)
);

NAND3xp33_ASAP7_75t_L g512 ( 
.A(n_427),
.B(n_44),
.C(n_45),
.Y(n_512)
);

A2O1A1Ixp33_ASAP7_75t_L g513 ( 
.A1(n_442),
.A2(n_365),
.B(n_370),
.C(n_379),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_454),
.B(n_390),
.Y(n_514)
);

AOI221xp5_ASAP7_75t_L g515 ( 
.A1(n_460),
.A2(n_391),
.B1(n_443),
.B2(n_412),
.C(n_377),
.Y(n_515)
);

O2A1O1Ixp33_ASAP7_75t_L g516 ( 
.A1(n_497),
.A2(n_432),
.B(n_410),
.C(n_383),
.Y(n_516)
);

INVx3_ASAP7_75t_L g517 ( 
.A(n_493),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_446),
.Y(n_518)
);

HB1xp67_ASAP7_75t_L g519 ( 
.A(n_485),
.Y(n_519)
);

AOI21xp5_ASAP7_75t_L g520 ( 
.A1(n_455),
.A2(n_411),
.B(n_379),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_SL g521 ( 
.A(n_476),
.B(n_495),
.Y(n_521)
);

OAI22xp5_ASAP7_75t_L g522 ( 
.A1(n_497),
.A2(n_425),
.B1(n_385),
.B2(n_402),
.Y(n_522)
);

AOI21xp5_ASAP7_75t_L g523 ( 
.A1(n_513),
.A2(n_426),
.B(n_385),
.Y(n_523)
);

AND2x2_ASAP7_75t_L g524 ( 
.A(n_472),
.B(n_383),
.Y(n_524)
);

O2A1O1Ixp33_ASAP7_75t_L g525 ( 
.A1(n_460),
.A2(n_428),
.B(n_411),
.C(n_430),
.Y(n_525)
);

HB1xp67_ASAP7_75t_L g526 ( 
.A(n_485),
.Y(n_526)
);

XOR2xp5_ASAP7_75t_L g527 ( 
.A(n_488),
.B(n_47),
.Y(n_527)
);

OAI21xp5_ASAP7_75t_L g528 ( 
.A1(n_487),
.A2(n_428),
.B(n_402),
.Y(n_528)
);

AND2x2_ASAP7_75t_L g529 ( 
.A(n_456),
.B(n_426),
.Y(n_529)
);

NOR2xp33_ASAP7_75t_R g530 ( 
.A(n_468),
.B(n_437),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_466),
.Y(n_531)
);

AO32x2_ASAP7_75t_L g532 ( 
.A1(n_500),
.A2(n_437),
.A3(n_394),
.B1(n_398),
.B2(n_408),
.Y(n_532)
);

CKINVDCx5p33_ASAP7_75t_R g533 ( 
.A(n_461),
.Y(n_533)
);

AOI21xp5_ASAP7_75t_L g534 ( 
.A1(n_469),
.A2(n_441),
.B(n_434),
.Y(n_534)
);

INVx4_ASAP7_75t_L g535 ( 
.A(n_459),
.Y(n_535)
);

AO21x1_ASAP7_75t_L g536 ( 
.A1(n_507),
.A2(n_56),
.B(n_57),
.Y(n_536)
);

NOR2xp33_ASAP7_75t_L g537 ( 
.A(n_505),
.B(n_491),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_470),
.Y(n_538)
);

O2A1O1Ixp33_ASAP7_75t_L g539 ( 
.A1(n_510),
.A2(n_175),
.B(n_92),
.C(n_97),
.Y(n_539)
);

O2A1O1Ixp33_ASAP7_75t_L g540 ( 
.A1(n_507),
.A2(n_89),
.B(n_99),
.C(n_100),
.Y(n_540)
);

OAI22xp5_ASAP7_75t_L g541 ( 
.A1(n_492),
.A2(n_104),
.B1(n_109),
.B2(n_111),
.Y(n_541)
);

AND2x2_ASAP7_75t_L g542 ( 
.A(n_459),
.B(n_115),
.Y(n_542)
);

OR2x6_ASAP7_75t_L g543 ( 
.A(n_492),
.B(n_117),
.Y(n_543)
);

INVx4_ASAP7_75t_L g544 ( 
.A(n_492),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_471),
.Y(n_545)
);

AOI21xp5_ASAP7_75t_L g546 ( 
.A1(n_501),
.A2(n_118),
.B(n_119),
.Y(n_546)
);

NOR2xp33_ASAP7_75t_L g547 ( 
.A(n_491),
.B(n_124),
.Y(n_547)
);

NOR2xp33_ASAP7_75t_L g548 ( 
.A(n_452),
.B(n_125),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_SL g549 ( 
.A(n_502),
.B(n_126),
.Y(n_549)
);

NOR2xp33_ASAP7_75t_L g550 ( 
.A(n_453),
.B(n_451),
.Y(n_550)
);

AOI21xp5_ASAP7_75t_L g551 ( 
.A1(n_508),
.A2(n_129),
.B(n_132),
.Y(n_551)
);

AOI21xp5_ASAP7_75t_L g552 ( 
.A1(n_445),
.A2(n_133),
.B(n_134),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_L g553 ( 
.A(n_475),
.B(n_172),
.Y(n_553)
);

NOR2xp33_ASAP7_75t_SL g554 ( 
.A(n_447),
.B(n_135),
.Y(n_554)
);

NOR3xp33_ASAP7_75t_L g555 ( 
.A(n_496),
.B(n_136),
.C(n_137),
.Y(n_555)
);

CKINVDCx6p67_ASAP7_75t_R g556 ( 
.A(n_509),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_SL g557 ( 
.A(n_461),
.B(n_138),
.Y(n_557)
);

AND2x4_ASAP7_75t_L g558 ( 
.A(n_509),
.B(n_467),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_SL g559 ( 
.A(n_464),
.B(n_145),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_L g560 ( 
.A(n_477),
.B(n_147),
.Y(n_560)
);

INVx6_ASAP7_75t_L g561 ( 
.A(n_498),
.Y(n_561)
);

BUFx12f_ASAP7_75t_L g562 ( 
.A(n_498),
.Y(n_562)
);

AOI22xp5_ASAP7_75t_L g563 ( 
.A1(n_509),
.A2(n_151),
.B1(n_152),
.B2(n_154),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_L g564 ( 
.A(n_477),
.B(n_161),
.Y(n_564)
);

HB1xp67_ASAP7_75t_L g565 ( 
.A(n_506),
.Y(n_565)
);

O2A1O1Ixp33_ASAP7_75t_L g566 ( 
.A1(n_479),
.A2(n_171),
.B(n_165),
.C(n_166),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_L g567 ( 
.A(n_465),
.B(n_164),
.Y(n_567)
);

OAI21xp33_ASAP7_75t_L g568 ( 
.A1(n_465),
.A2(n_457),
.B(n_481),
.Y(n_568)
);

OR2x2_ASAP7_75t_L g569 ( 
.A(n_463),
.B(n_170),
.Y(n_569)
);

O2A1O1Ixp5_ASAP7_75t_L g570 ( 
.A1(n_503),
.A2(n_474),
.B(n_457),
.C(n_463),
.Y(n_570)
);

AOI21xp5_ASAP7_75t_L g571 ( 
.A1(n_458),
.A2(n_473),
.B(n_478),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_L g572 ( 
.A(n_483),
.B(n_490),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_SL g573 ( 
.A(n_494),
.B(n_462),
.Y(n_573)
);

INVx3_ASAP7_75t_SL g574 ( 
.A(n_449),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_503),
.B(n_484),
.Y(n_575)
);

AO21x1_ASAP7_75t_L g576 ( 
.A1(n_486),
.A2(n_482),
.B(n_450),
.Y(n_576)
);

AOI21xp5_ASAP7_75t_L g577 ( 
.A1(n_504),
.A2(n_480),
.B(n_499),
.Y(n_577)
);

AO22x1_ASAP7_75t_L g578 ( 
.A1(n_511),
.A2(n_512),
.B1(n_499),
.B2(n_480),
.Y(n_578)
);

OAI21xp33_ASAP7_75t_L g579 ( 
.A1(n_489),
.A2(n_446),
.B(n_433),
.Y(n_579)
);

AOI21xp5_ASAP7_75t_L g580 ( 
.A1(n_489),
.A2(n_455),
.B(n_442),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_L g581 ( 
.A(n_446),
.B(n_433),
.Y(n_581)
);

AND2x2_ASAP7_75t_L g582 ( 
.A(n_446),
.B(n_420),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_581),
.Y(n_583)
);

BUFx3_ASAP7_75t_L g584 ( 
.A(n_562),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_518),
.Y(n_585)
);

A2O1A1Ixp33_ASAP7_75t_L g586 ( 
.A1(n_568),
.A2(n_570),
.B(n_550),
.C(n_571),
.Y(n_586)
);

INVx1_ASAP7_75t_SL g587 ( 
.A(n_561),
.Y(n_587)
);

OAI21xp5_ASAP7_75t_L g588 ( 
.A1(n_528),
.A2(n_577),
.B(n_525),
.Y(n_588)
);

O2A1O1Ixp5_ASAP7_75t_L g589 ( 
.A1(n_573),
.A2(n_559),
.B(n_576),
.C(n_548),
.Y(n_589)
);

AO31x2_ASAP7_75t_L g590 ( 
.A1(n_522),
.A2(n_536),
.A3(n_541),
.B(n_567),
.Y(n_590)
);

A2O1A1Ixp33_ASAP7_75t_L g591 ( 
.A1(n_516),
.A2(n_575),
.B(n_579),
.C(n_567),
.Y(n_591)
);

AOI21x1_ASAP7_75t_L g592 ( 
.A1(n_522),
.A2(n_560),
.B(n_564),
.Y(n_592)
);

AOI21x1_ASAP7_75t_L g593 ( 
.A1(n_560),
.A2(n_564),
.B(n_553),
.Y(n_593)
);

BUFx6f_ASAP7_75t_L g594 ( 
.A(n_543),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_L g595 ( 
.A(n_524),
.B(n_529),
.Y(n_595)
);

INVx5_ASAP7_75t_L g596 ( 
.A(n_543),
.Y(n_596)
);

BUFx6f_ASAP7_75t_L g597 ( 
.A(n_517),
.Y(n_597)
);

O2A1O1Ixp33_ASAP7_75t_SL g598 ( 
.A1(n_557),
.A2(n_569),
.B(n_541),
.C(n_549),
.Y(n_598)
);

AND2x2_ASAP7_75t_SL g599 ( 
.A(n_544),
.B(n_515),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_531),
.Y(n_600)
);

AND2x2_ASAP7_75t_L g601 ( 
.A(n_565),
.B(n_561),
.Y(n_601)
);

AOI21xp5_ASAP7_75t_L g602 ( 
.A1(n_534),
.A2(n_572),
.B(n_521),
.Y(n_602)
);

INVx5_ASAP7_75t_L g603 ( 
.A(n_535),
.Y(n_603)
);

HB1xp67_ASAP7_75t_L g604 ( 
.A(n_519),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_545),
.Y(n_605)
);

INVx1_ASAP7_75t_SL g606 ( 
.A(n_556),
.Y(n_606)
);

AO31x2_ASAP7_75t_L g607 ( 
.A1(n_546),
.A2(n_551),
.A3(n_547),
.B(n_552),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_514),
.B(n_537),
.Y(n_608)
);

OAI21x1_ASAP7_75t_SL g609 ( 
.A1(n_544),
.A2(n_540),
.B(n_563),
.Y(n_609)
);

NOR2xp33_ASAP7_75t_L g610 ( 
.A(n_514),
.B(n_535),
.Y(n_610)
);

BUFx4f_ASAP7_75t_SL g611 ( 
.A(n_574),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_SL g612 ( 
.A(n_530),
.B(n_526),
.Y(n_612)
);

NAND2xp33_ASAP7_75t_L g613 ( 
.A(n_533),
.B(n_542),
.Y(n_613)
);

INVx8_ASAP7_75t_L g614 ( 
.A(n_558),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_527),
.Y(n_615)
);

BUFx4_ASAP7_75t_SL g616 ( 
.A(n_554),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_L g617 ( 
.A(n_578),
.B(n_554),
.Y(n_617)
);

BUFx6f_ASAP7_75t_L g618 ( 
.A(n_532),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_L g619 ( 
.A(n_532),
.B(n_582),
.Y(n_619)
);

AND2x4_ASAP7_75t_L g620 ( 
.A(n_532),
.B(n_518),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_L g621 ( 
.A(n_582),
.B(n_581),
.Y(n_621)
);

INVxp67_ASAP7_75t_SL g622 ( 
.A(n_581),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_582),
.B(n_581),
.Y(n_623)
);

NOR2xp33_ASAP7_75t_L g624 ( 
.A(n_561),
.B(n_456),
.Y(n_624)
);

INVx1_ASAP7_75t_SL g625 ( 
.A(n_561),
.Y(n_625)
);

AOI21xp5_ASAP7_75t_L g626 ( 
.A1(n_580),
.A2(n_455),
.B(n_571),
.Y(n_626)
);

AOI21xp5_ASAP7_75t_L g627 ( 
.A1(n_580),
.A2(n_455),
.B(n_571),
.Y(n_627)
);

OAI22xp5_ASAP7_75t_L g628 ( 
.A1(n_565),
.A2(n_543),
.B1(n_572),
.B2(n_581),
.Y(n_628)
);

OAI22xp5_ASAP7_75t_L g629 ( 
.A1(n_565),
.A2(n_543),
.B1(n_572),
.B2(n_581),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_581),
.Y(n_630)
);

AOI21xp5_ASAP7_75t_L g631 ( 
.A1(n_580),
.A2(n_455),
.B(n_571),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_581),
.Y(n_632)
);

BUFx2_ASAP7_75t_L g633 ( 
.A(n_562),
.Y(n_633)
);

BUFx6f_ASAP7_75t_L g634 ( 
.A(n_543),
.Y(n_634)
);

O2A1O1Ixp5_ASAP7_75t_SL g635 ( 
.A1(n_541),
.A2(n_353),
.B(n_341),
.C(n_342),
.Y(n_635)
);

OAI21xp5_ASAP7_75t_L g636 ( 
.A1(n_570),
.A2(n_571),
.B(n_580),
.Y(n_636)
);

OR2x2_ASAP7_75t_L g637 ( 
.A(n_582),
.B(n_354),
.Y(n_637)
);

OR2x6_ASAP7_75t_L g638 ( 
.A(n_562),
.B(n_543),
.Y(n_638)
);

INVx4_ASAP7_75t_L g639 ( 
.A(n_543),
.Y(n_639)
);

NAND3x1_ASAP7_75t_L g640 ( 
.A(n_515),
.B(n_349),
.C(n_358),
.Y(n_640)
);

OAI21xp5_ASAP7_75t_L g641 ( 
.A1(n_570),
.A2(n_571),
.B(n_580),
.Y(n_641)
);

OAI22xp5_ASAP7_75t_L g642 ( 
.A1(n_565),
.A2(n_543),
.B1(n_572),
.B2(n_581),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_L g643 ( 
.A(n_582),
.B(n_581),
.Y(n_643)
);

O2A1O1Ixp33_ASAP7_75t_SL g644 ( 
.A1(n_567),
.A2(n_559),
.B(n_564),
.C(n_560),
.Y(n_644)
);

A2O1A1Ixp33_ASAP7_75t_L g645 ( 
.A1(n_568),
.A2(n_570),
.B(n_550),
.C(n_571),
.Y(n_645)
);

INVxp67_ASAP7_75t_SL g646 ( 
.A(n_581),
.Y(n_646)
);

AOI21xp5_ASAP7_75t_L g647 ( 
.A1(n_580),
.A2(n_455),
.B(n_571),
.Y(n_647)
);

AOI21xp5_ASAP7_75t_L g648 ( 
.A1(n_580),
.A2(n_455),
.B(n_571),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_581),
.Y(n_649)
);

NAND2x1_ASAP7_75t_L g650 ( 
.A(n_517),
.B(n_543),
.Y(n_650)
);

AO31x2_ASAP7_75t_L g651 ( 
.A1(n_522),
.A2(n_576),
.A3(n_536),
.B(n_523),
.Y(n_651)
);

OAI21x1_ASAP7_75t_SL g652 ( 
.A1(n_536),
.A2(n_544),
.B(n_541),
.Y(n_652)
);

A2O1A1Ixp33_ASAP7_75t_L g653 ( 
.A1(n_568),
.A2(n_570),
.B(n_550),
.C(n_571),
.Y(n_653)
);

OAI22xp5_ASAP7_75t_L g654 ( 
.A1(n_565),
.A2(n_543),
.B1(n_572),
.B2(n_581),
.Y(n_654)
);

AOI221x1_ASAP7_75t_L g655 ( 
.A1(n_555),
.A2(n_541),
.B1(n_522),
.B2(n_568),
.C(n_520),
.Y(n_655)
);

CKINVDCx5p33_ASAP7_75t_R g656 ( 
.A(n_562),
.Y(n_656)
);

OAI21xp5_ASAP7_75t_L g657 ( 
.A1(n_570),
.A2(n_571),
.B(n_580),
.Y(n_657)
);

AO31x2_ASAP7_75t_L g658 ( 
.A1(n_522),
.A2(n_576),
.A3(n_536),
.B(n_523),
.Y(n_658)
);

BUFx5_ASAP7_75t_L g659 ( 
.A(n_538),
.Y(n_659)
);

AOI221x1_ASAP7_75t_L g660 ( 
.A1(n_555),
.A2(n_541),
.B1(n_522),
.B2(n_568),
.C(n_520),
.Y(n_660)
);

OAI22x1_ASAP7_75t_L g661 ( 
.A1(n_527),
.A2(n_448),
.B1(n_354),
.B2(n_429),
.Y(n_661)
);

BUFx6f_ASAP7_75t_L g662 ( 
.A(n_543),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_581),
.Y(n_663)
);

AO21x1_ASAP7_75t_L g664 ( 
.A1(n_541),
.A2(n_566),
.B(n_539),
.Y(n_664)
);

AOI221xp5_ASAP7_75t_L g665 ( 
.A1(n_581),
.A2(n_460),
.B1(n_391),
.B2(n_443),
.C(n_518),
.Y(n_665)
);

INVx2_ASAP7_75t_L g666 ( 
.A(n_605),
.Y(n_666)
);

INVx3_ASAP7_75t_L g667 ( 
.A(n_650),
.Y(n_667)
);

AOI21xp5_ASAP7_75t_L g668 ( 
.A1(n_644),
.A2(n_627),
.B(n_626),
.Y(n_668)
);

AND2x2_ASAP7_75t_L g669 ( 
.A(n_583),
.B(n_630),
.Y(n_669)
);

OA21x2_ASAP7_75t_L g670 ( 
.A1(n_588),
.A2(n_641),
.B(n_636),
.Y(n_670)
);

HB1xp67_ASAP7_75t_L g671 ( 
.A(n_622),
.Y(n_671)
);

AO21x2_ASAP7_75t_L g672 ( 
.A1(n_652),
.A2(n_617),
.B(n_657),
.Y(n_672)
);

OAI21x1_ASAP7_75t_SL g673 ( 
.A1(n_639),
.A2(n_629),
.B(n_654),
.Y(n_673)
);

AOI21xp5_ASAP7_75t_L g674 ( 
.A1(n_631),
.A2(n_648),
.B(n_647),
.Y(n_674)
);

AO31x2_ASAP7_75t_L g675 ( 
.A1(n_591),
.A2(n_645),
.A3(n_586),
.B(n_653),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_632),
.B(n_649),
.Y(n_676)
);

BUFx3_ASAP7_75t_L g677 ( 
.A(n_603),
.Y(n_677)
);

INVx1_ASAP7_75t_SL g678 ( 
.A(n_621),
.Y(n_678)
);

AO21x1_ASAP7_75t_L g679 ( 
.A1(n_628),
.A2(n_642),
.B(n_639),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_585),
.Y(n_680)
);

BUFx12f_ASAP7_75t_L g681 ( 
.A(n_656),
.Y(n_681)
);

OA21x2_ASAP7_75t_L g682 ( 
.A1(n_655),
.A2(n_660),
.B(n_589),
.Y(n_682)
);

AOI21xp33_ASAP7_75t_SL g683 ( 
.A1(n_638),
.A2(n_661),
.B(n_599),
.Y(n_683)
);

OAI21xp5_ASAP7_75t_L g684 ( 
.A1(n_635),
.A2(n_619),
.B(n_602),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_600),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_663),
.Y(n_686)
);

AND2x2_ASAP7_75t_L g687 ( 
.A(n_623),
.B(n_643),
.Y(n_687)
);

OAI21x1_ASAP7_75t_SL g688 ( 
.A1(n_609),
.A2(n_616),
.B(n_664),
.Y(n_688)
);

INVx2_ASAP7_75t_SL g689 ( 
.A(n_603),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_595),
.Y(n_690)
);

CKINVDCx5p33_ASAP7_75t_R g691 ( 
.A(n_611),
.Y(n_691)
);

NOR2xp67_ASAP7_75t_L g692 ( 
.A(n_596),
.B(n_603),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_L g693 ( 
.A(n_665),
.B(n_608),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_601),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_604),
.Y(n_695)
);

OAI21xp5_ASAP7_75t_L g696 ( 
.A1(n_620),
.A2(n_640),
.B(n_598),
.Y(n_696)
);

OA21x2_ASAP7_75t_L g697 ( 
.A1(n_651),
.A2(n_658),
.B(n_618),
.Y(n_697)
);

NAND3xp33_ASAP7_75t_L g698 ( 
.A(n_610),
.B(n_662),
.C(n_634),
.Y(n_698)
);

INVx3_ASAP7_75t_L g699 ( 
.A(n_594),
.Y(n_699)
);

OA21x2_ASAP7_75t_L g700 ( 
.A1(n_651),
.A2(n_658),
.B(n_618),
.Y(n_700)
);

OAI21xp5_ASAP7_75t_L g701 ( 
.A1(n_624),
.A2(n_613),
.B(n_612),
.Y(n_701)
);

AO21x2_ASAP7_75t_L g702 ( 
.A1(n_590),
.A2(n_607),
.B(n_659),
.Y(n_702)
);

OR2x6_ASAP7_75t_L g703 ( 
.A(n_614),
.B(n_584),
.Y(n_703)
);

CKINVDCx6p67_ASAP7_75t_R g704 ( 
.A(n_633),
.Y(n_704)
);

AOI31xp33_ASAP7_75t_L g705 ( 
.A1(n_606),
.A2(n_615),
.A3(n_637),
.B(n_587),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_625),
.Y(n_706)
);

AOI21xp5_ASAP7_75t_L g707 ( 
.A1(n_597),
.A2(n_607),
.B(n_614),
.Y(n_707)
);

AND2x4_ASAP7_75t_L g708 ( 
.A(n_583),
.B(n_630),
.Y(n_708)
);

INVx2_ASAP7_75t_SL g709 ( 
.A(n_603),
.Y(n_709)
);

AOI21x1_ASAP7_75t_L g710 ( 
.A1(n_593),
.A2(n_617),
.B(n_592),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_622),
.Y(n_711)
);

BUFx2_ASAP7_75t_R g712 ( 
.A(n_656),
.Y(n_712)
);

NOR2xp33_ASAP7_75t_L g713 ( 
.A(n_621),
.B(n_623),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_622),
.Y(n_714)
);

INVxp67_ASAP7_75t_L g715 ( 
.A(n_622),
.Y(n_715)
);

OAI21xp5_ASAP7_75t_L g716 ( 
.A1(n_586),
.A2(n_653),
.B(n_645),
.Y(n_716)
);

OA21x2_ASAP7_75t_L g717 ( 
.A1(n_588),
.A2(n_641),
.B(n_636),
.Y(n_717)
);

NOR2xp67_ASAP7_75t_L g718 ( 
.A(n_596),
.B(n_562),
.Y(n_718)
);

CKINVDCx6p67_ASAP7_75t_R g719 ( 
.A(n_584),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_622),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_622),
.B(n_646),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_622),
.Y(n_722)
);

BUFx4_ASAP7_75t_SL g723 ( 
.A(n_638),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_622),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_622),
.Y(n_725)
);

HB1xp67_ASAP7_75t_L g726 ( 
.A(n_622),
.Y(n_726)
);

OA21x2_ASAP7_75t_L g727 ( 
.A1(n_588),
.A2(n_641),
.B(n_636),
.Y(n_727)
);

AND2x2_ASAP7_75t_L g728 ( 
.A(n_583),
.B(n_582),
.Y(n_728)
);

BUFx2_ASAP7_75t_L g729 ( 
.A(n_638),
.Y(n_729)
);

NOR2xp33_ASAP7_75t_L g730 ( 
.A(n_621),
.B(n_623),
.Y(n_730)
);

CKINVDCx11_ASAP7_75t_R g731 ( 
.A(n_638),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_669),
.Y(n_732)
);

INVx4_ASAP7_75t_L g733 ( 
.A(n_677),
.Y(n_733)
);

AND2x2_ASAP7_75t_L g734 ( 
.A(n_687),
.B(n_678),
.Y(n_734)
);

OAI21xp5_ASAP7_75t_L g735 ( 
.A1(n_721),
.A2(n_693),
.B(n_715),
.Y(n_735)
);

HB1xp67_ASAP7_75t_L g736 ( 
.A(n_671),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_686),
.Y(n_737)
);

OR2x2_ASAP7_75t_L g738 ( 
.A(n_678),
.B(n_721),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_713),
.B(n_730),
.Y(n_739)
);

AND2x2_ASAP7_75t_L g740 ( 
.A(n_713),
.B(n_730),
.Y(n_740)
);

AND2x2_ASAP7_75t_L g741 ( 
.A(n_726),
.B(n_715),
.Y(n_741)
);

AND2x2_ASAP7_75t_L g742 ( 
.A(n_726),
.B(n_666),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_676),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_666),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_685),
.Y(n_745)
);

INVxp67_ASAP7_75t_L g746 ( 
.A(n_728),
.Y(n_746)
);

INVx2_ASAP7_75t_SL g747 ( 
.A(n_677),
.Y(n_747)
);

AND2x2_ASAP7_75t_L g748 ( 
.A(n_708),
.B(n_711),
.Y(n_748)
);

INVx1_ASAP7_75t_SL g749 ( 
.A(n_704),
.Y(n_749)
);

HB1xp67_ASAP7_75t_L g750 ( 
.A(n_690),
.Y(n_750)
);

BUFx12f_ASAP7_75t_L g751 ( 
.A(n_731),
.Y(n_751)
);

CKINVDCx5p33_ASAP7_75t_R g752 ( 
.A(n_723),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_680),
.Y(n_753)
);

AOI21x1_ASAP7_75t_L g754 ( 
.A1(n_710),
.A2(n_668),
.B(n_674),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_714),
.Y(n_755)
);

HB1xp67_ASAP7_75t_L g756 ( 
.A(n_720),
.Y(n_756)
);

HB1xp67_ASAP7_75t_L g757 ( 
.A(n_722),
.Y(n_757)
);

BUFx2_ASAP7_75t_SL g758 ( 
.A(n_692),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_693),
.B(n_694),
.Y(n_759)
);

OR2x6_ASAP7_75t_L g760 ( 
.A(n_673),
.B(n_688),
.Y(n_760)
);

INVx2_ASAP7_75t_L g761 ( 
.A(n_670),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_724),
.Y(n_762)
);

NOR2xp33_ASAP7_75t_L g763 ( 
.A(n_705),
.B(n_683),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_725),
.Y(n_764)
);

AO21x2_ASAP7_75t_L g765 ( 
.A1(n_716),
.A2(n_684),
.B(n_696),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_717),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_727),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_695),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_706),
.Y(n_769)
);

AND2x2_ASAP7_75t_L g770 ( 
.A(n_702),
.B(n_700),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_707),
.Y(n_771)
);

OAI21xp5_ASAP7_75t_L g772 ( 
.A1(n_707),
.A2(n_705),
.B(n_698),
.Y(n_772)
);

HB1xp67_ASAP7_75t_L g773 ( 
.A(n_723),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_689),
.Y(n_774)
);

AND2x2_ASAP7_75t_L g775 ( 
.A(n_697),
.B(n_700),
.Y(n_775)
);

HB1xp67_ASAP7_75t_L g776 ( 
.A(n_709),
.Y(n_776)
);

INVx2_ASAP7_75t_L g777 ( 
.A(n_675),
.Y(n_777)
);

AND2x2_ASAP7_75t_L g778 ( 
.A(n_672),
.B(n_699),
.Y(n_778)
);

INVx2_ASAP7_75t_L g779 ( 
.A(n_761),
.Y(n_779)
);

AND2x2_ASAP7_75t_L g780 ( 
.A(n_770),
.B(n_682),
.Y(n_780)
);

AND2x2_ASAP7_75t_L g781 ( 
.A(n_770),
.B(n_682),
.Y(n_781)
);

AND2x4_ASAP7_75t_L g782 ( 
.A(n_771),
.B(n_775),
.Y(n_782)
);

OR2x2_ASAP7_75t_L g783 ( 
.A(n_738),
.B(n_736),
.Y(n_783)
);

AOI22xp33_ASAP7_75t_L g784 ( 
.A1(n_740),
.A2(n_731),
.B1(n_679),
.B2(n_729),
.Y(n_784)
);

HB1xp67_ASAP7_75t_L g785 ( 
.A(n_742),
.Y(n_785)
);

HB1xp67_ASAP7_75t_L g786 ( 
.A(n_742),
.Y(n_786)
);

NOR2x1_ASAP7_75t_L g787 ( 
.A(n_733),
.B(n_667),
.Y(n_787)
);

HB1xp67_ASAP7_75t_L g788 ( 
.A(n_741),
.Y(n_788)
);

BUFx3_ASAP7_75t_L g789 ( 
.A(n_733),
.Y(n_789)
);

AO21x2_ASAP7_75t_L g790 ( 
.A1(n_754),
.A2(n_701),
.B(n_718),
.Y(n_790)
);

INVxp67_ASAP7_75t_L g791 ( 
.A(n_735),
.Y(n_791)
);

AOI22xp33_ASAP7_75t_L g792 ( 
.A1(n_740),
.A2(n_763),
.B1(n_739),
.B2(n_734),
.Y(n_792)
);

CKINVDCx5p33_ASAP7_75t_R g793 ( 
.A(n_751),
.Y(n_793)
);

NAND4xp25_ASAP7_75t_L g794 ( 
.A(n_759),
.B(n_712),
.C(n_719),
.D(n_703),
.Y(n_794)
);

AND2x2_ASAP7_75t_L g795 ( 
.A(n_777),
.B(n_712),
.Y(n_795)
);

OR2x2_ASAP7_75t_L g796 ( 
.A(n_744),
.B(n_691),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_743),
.B(n_691),
.Y(n_797)
);

OR2x2_ASAP7_75t_L g798 ( 
.A(n_785),
.B(n_734),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_783),
.Y(n_799)
);

INVx2_ASAP7_75t_L g800 ( 
.A(n_779),
.Y(n_800)
);

AND2x2_ASAP7_75t_L g801 ( 
.A(n_780),
.B(n_778),
.Y(n_801)
);

AND2x2_ASAP7_75t_L g802 ( 
.A(n_780),
.B(n_765),
.Y(n_802)
);

AND2x2_ASAP7_75t_L g803 ( 
.A(n_780),
.B(n_765),
.Y(n_803)
);

INVx3_ASAP7_75t_L g804 ( 
.A(n_789),
.Y(n_804)
);

AND2x2_ASAP7_75t_L g805 ( 
.A(n_781),
.B(n_766),
.Y(n_805)
);

OR2x2_ASAP7_75t_L g806 ( 
.A(n_786),
.B(n_766),
.Y(n_806)
);

INVxp67_ASAP7_75t_L g807 ( 
.A(n_789),
.Y(n_807)
);

AND2x2_ASAP7_75t_L g808 ( 
.A(n_781),
.B(n_767),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_L g809 ( 
.A(n_788),
.B(n_750),
.Y(n_809)
);

NAND2x1p5_ASAP7_75t_L g810 ( 
.A(n_789),
.B(n_733),
.Y(n_810)
);

NOR2x1p5_ASAP7_75t_L g811 ( 
.A(n_804),
.B(n_794),
.Y(n_811)
);

AND2x2_ASAP7_75t_L g812 ( 
.A(n_801),
.B(n_782),
.Y(n_812)
);

NOR2x1p5_ASAP7_75t_L g813 ( 
.A(n_804),
.B(n_794),
.Y(n_813)
);

INVx2_ASAP7_75t_L g814 ( 
.A(n_800),
.Y(n_814)
);

AND2x4_ASAP7_75t_L g815 ( 
.A(n_804),
.B(n_782),
.Y(n_815)
);

AND2x2_ASAP7_75t_L g816 ( 
.A(n_801),
.B(n_782),
.Y(n_816)
);

NAND2x1p5_ASAP7_75t_L g817 ( 
.A(n_810),
.B(n_787),
.Y(n_817)
);

AND2x2_ASAP7_75t_L g818 ( 
.A(n_802),
.B(n_803),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_L g819 ( 
.A(n_799),
.B(n_791),
.Y(n_819)
);

NOR2x1_ASAP7_75t_L g820 ( 
.A(n_809),
.B(n_758),
.Y(n_820)
);

INVx2_ASAP7_75t_SL g821 ( 
.A(n_810),
.Y(n_821)
);

INVx3_ASAP7_75t_L g822 ( 
.A(n_810),
.Y(n_822)
);

INVx3_ASAP7_75t_SL g823 ( 
.A(n_806),
.Y(n_823)
);

INVx1_ASAP7_75t_SL g824 ( 
.A(n_798),
.Y(n_824)
);

OR2x2_ASAP7_75t_L g825 ( 
.A(n_824),
.B(n_805),
.Y(n_825)
);

AND2x2_ASAP7_75t_L g826 ( 
.A(n_818),
.B(n_805),
.Y(n_826)
);

INVx2_ASAP7_75t_L g827 ( 
.A(n_814),
.Y(n_827)
);

AND2x4_ASAP7_75t_L g828 ( 
.A(n_815),
.B(n_808),
.Y(n_828)
);

AND2x2_ASAP7_75t_L g829 ( 
.A(n_818),
.B(n_808),
.Y(n_829)
);

NAND2x1p5_ASAP7_75t_L g830 ( 
.A(n_822),
.B(n_821),
.Y(n_830)
);

BUFx3_ASAP7_75t_L g831 ( 
.A(n_817),
.Y(n_831)
);

INVx1_ASAP7_75t_SL g832 ( 
.A(n_823),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_819),
.B(n_791),
.Y(n_833)
);

INVxp67_ASAP7_75t_L g834 ( 
.A(n_820),
.Y(n_834)
);

OR2x6_ASAP7_75t_L g835 ( 
.A(n_831),
.B(n_811),
.Y(n_835)
);

AOI32xp33_ASAP7_75t_L g836 ( 
.A1(n_832),
.A2(n_822),
.A3(n_816),
.B1(n_812),
.B2(n_821),
.Y(n_836)
);

O2A1O1Ixp33_ASAP7_75t_SL g837 ( 
.A1(n_834),
.A2(n_773),
.B(n_749),
.C(n_822),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_826),
.B(n_823),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_825),
.Y(n_839)
);

INVxp67_ASAP7_75t_L g840 ( 
.A(n_833),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_825),
.Y(n_841)
);

INVx2_ASAP7_75t_L g842 ( 
.A(n_827),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_826),
.B(n_823),
.Y(n_843)
);

OAI22xp5_ASAP7_75t_L g844 ( 
.A1(n_831),
.A2(n_811),
.B1(n_813),
.B2(n_817),
.Y(n_844)
);

NOR2xp33_ASAP7_75t_L g845 ( 
.A(n_828),
.B(n_751),
.Y(n_845)
);

OAI21xp5_ASAP7_75t_L g846 ( 
.A1(n_830),
.A2(n_817),
.B(n_784),
.Y(n_846)
);

INVx3_ASAP7_75t_L g847 ( 
.A(n_831),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_L g848 ( 
.A(n_840),
.B(n_839),
.Y(n_848)
);

O2A1O1Ixp33_ASAP7_75t_L g849 ( 
.A1(n_837),
.A2(n_797),
.B(n_784),
.C(n_813),
.Y(n_849)
);

AOI22xp5_ASAP7_75t_SL g850 ( 
.A1(n_845),
.A2(n_752),
.B1(n_793),
.B2(n_830),
.Y(n_850)
);

AOI22xp5_ASAP7_75t_L g851 ( 
.A1(n_835),
.A2(n_828),
.B1(n_815),
.B2(n_816),
.Y(n_851)
);

AOI21xp5_ASAP7_75t_SL g852 ( 
.A1(n_844),
.A2(n_752),
.B(n_830),
.Y(n_852)
);

O2A1O1Ixp33_ASAP7_75t_L g853 ( 
.A1(n_835),
.A2(n_797),
.B(n_772),
.C(n_776),
.Y(n_853)
);

AOI21xp5_ASAP7_75t_L g854 ( 
.A1(n_852),
.A2(n_846),
.B(n_836),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_L g855 ( 
.A(n_848),
.B(n_841),
.Y(n_855)
);

OAI21xp33_ASAP7_75t_L g856 ( 
.A1(n_851),
.A2(n_843),
.B(n_838),
.Y(n_856)
);

OAI221xp5_ASAP7_75t_L g857 ( 
.A1(n_854),
.A2(n_849),
.B1(n_856),
.B2(n_850),
.C(n_853),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_L g858 ( 
.A(n_855),
.B(n_829),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_858),
.Y(n_859)
);

NOR2xp67_ASAP7_75t_L g860 ( 
.A(n_857),
.B(n_847),
.Y(n_860)
);

NAND2x1p5_ASAP7_75t_L g861 ( 
.A(n_860),
.B(n_847),
.Y(n_861)
);

AND2x2_ASAP7_75t_SL g862 ( 
.A(n_859),
.B(n_758),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_861),
.Y(n_863)
);

AOI22xp5_ASAP7_75t_L g864 ( 
.A1(n_862),
.A2(n_681),
.B1(n_795),
.B2(n_828),
.Y(n_864)
);

NOR2xp33_ASAP7_75t_R g865 ( 
.A(n_863),
.B(n_774),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_L g866 ( 
.A(n_864),
.B(n_842),
.Y(n_866)
);

AO22x2_ASAP7_75t_L g867 ( 
.A1(n_863),
.A2(n_768),
.B1(n_769),
.B2(n_746),
.Y(n_867)
);

AOI21xp5_ASAP7_75t_L g868 ( 
.A1(n_866),
.A2(n_867),
.B(n_865),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_867),
.Y(n_869)
);

AO221x2_ASAP7_75t_L g870 ( 
.A1(n_866),
.A2(n_732),
.B1(n_737),
.B2(n_745),
.C(n_753),
.Y(n_870)
);

OAI22xp5_ASAP7_75t_SL g871 ( 
.A1(n_866),
.A2(n_792),
.B1(n_747),
.B2(n_760),
.Y(n_871)
);

AOI21xp33_ASAP7_75t_SL g872 ( 
.A1(n_869),
.A2(n_747),
.B(n_796),
.Y(n_872)
);

O2A1O1Ixp33_ASAP7_75t_L g873 ( 
.A1(n_868),
.A2(n_753),
.B(n_745),
.C(n_757),
.Y(n_873)
);

OAI22x1_ASAP7_75t_SL g874 ( 
.A1(n_870),
.A2(n_755),
.B1(n_764),
.B2(n_762),
.Y(n_874)
);

OA21x2_ASAP7_75t_L g875 ( 
.A1(n_871),
.A2(n_792),
.B(n_807),
.Y(n_875)
);

XNOR2xp5_ASAP7_75t_L g876 ( 
.A(n_868),
.B(n_748),
.Y(n_876)
);

OAI21x1_ASAP7_75t_L g877 ( 
.A1(n_869),
.A2(n_787),
.B(n_796),
.Y(n_877)
);

HB1xp67_ASAP7_75t_L g878 ( 
.A(n_877),
.Y(n_878)
);

AOI21xp5_ASAP7_75t_L g879 ( 
.A1(n_873),
.A2(n_756),
.B(n_795),
.Y(n_879)
);

OAI22xp33_ASAP7_75t_L g880 ( 
.A1(n_878),
.A2(n_875),
.B1(n_872),
.B2(n_879),
.Y(n_880)
);

AOI31xp33_ASAP7_75t_L g881 ( 
.A1(n_878),
.A2(n_876),
.A3(n_874),
.B(n_796),
.Y(n_881)
);

OR2x6_ASAP7_75t_L g882 ( 
.A(n_881),
.B(n_880),
.Y(n_882)
);

AOI22xp33_ASAP7_75t_L g883 ( 
.A1(n_882),
.A2(n_828),
.B1(n_795),
.B2(n_790),
.Y(n_883)
);


endmodule