module fake_netlist_1_838_n_695 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_695);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_695;
wire n_117;
wire n_663;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_85;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_624;
wire n_255;
wire n_426;
wire n_108;
wire n_91;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_90;
wire n_357;
wire n_653;
wire n_260;
wire n_539;
wire n_201;
wire n_197;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_684;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_487;
wire n_451;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_84;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g79 ( .A(n_36), .Y(n_79) );
CKINVDCx14_ASAP7_75t_R g80 ( .A(n_27), .Y(n_80) );
INVx1_ASAP7_75t_L g81 ( .A(n_57), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_38), .Y(n_82) );
CKINVDCx20_ASAP7_75t_R g83 ( .A(n_53), .Y(n_83) );
INVx1_ASAP7_75t_L g84 ( .A(n_12), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_64), .Y(n_85) );
CKINVDCx5p33_ASAP7_75t_R g86 ( .A(n_73), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_13), .Y(n_87) );
CKINVDCx20_ASAP7_75t_R g88 ( .A(n_47), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_77), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_6), .Y(n_90) );
INVxp67_ASAP7_75t_SL g91 ( .A(n_6), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_9), .Y(n_92) );
CKINVDCx5p33_ASAP7_75t_R g93 ( .A(n_52), .Y(n_93) );
INVxp67_ASAP7_75t_SL g94 ( .A(n_15), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_19), .Y(n_95) );
INVx2_ASAP7_75t_L g96 ( .A(n_30), .Y(n_96) );
CKINVDCx5p33_ASAP7_75t_R g97 ( .A(n_20), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_37), .Y(n_98) );
INVxp33_ASAP7_75t_L g99 ( .A(n_24), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_59), .Y(n_100) );
CKINVDCx16_ASAP7_75t_R g101 ( .A(n_67), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_9), .Y(n_102) );
INVx2_ASAP7_75t_L g103 ( .A(n_70), .Y(n_103) );
INVxp67_ASAP7_75t_SL g104 ( .A(n_31), .Y(n_104) );
INVxp67_ASAP7_75t_SL g105 ( .A(n_13), .Y(n_105) );
BUFx6f_ASAP7_75t_L g106 ( .A(n_43), .Y(n_106) );
INVx2_ASAP7_75t_L g107 ( .A(n_55), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_33), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_58), .Y(n_109) );
BUFx3_ASAP7_75t_L g110 ( .A(n_46), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_34), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_42), .Y(n_112) );
INVxp67_ASAP7_75t_SL g113 ( .A(n_35), .Y(n_113) );
CKINVDCx5p33_ASAP7_75t_R g114 ( .A(n_26), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_8), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_56), .Y(n_116) );
INVxp67_ASAP7_75t_L g117 ( .A(n_8), .Y(n_117) );
CKINVDCx5p33_ASAP7_75t_R g118 ( .A(n_72), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_50), .Y(n_119) );
INVxp67_ASAP7_75t_SL g120 ( .A(n_65), .Y(n_120) );
INVxp67_ASAP7_75t_L g121 ( .A(n_48), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_0), .Y(n_122) );
INVxp33_ASAP7_75t_SL g123 ( .A(n_4), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_11), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_54), .Y(n_125) );
CKINVDCx20_ASAP7_75t_R g126 ( .A(n_4), .Y(n_126) );
BUFx6f_ASAP7_75t_L g127 ( .A(n_106), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_79), .Y(n_128) );
INVx1_ASAP7_75t_L g129 ( .A(n_79), .Y(n_129) );
NAND2xp5_ASAP7_75t_L g130 ( .A(n_117), .B(n_0), .Y(n_130) );
INVx1_ASAP7_75t_L g131 ( .A(n_81), .Y(n_131) );
AND2x4_ASAP7_75t_L g132 ( .A(n_84), .B(n_1), .Y(n_132) );
XOR2xp5_ASAP7_75t_L g133 ( .A(n_126), .B(n_1), .Y(n_133) );
INVx2_ASAP7_75t_L g134 ( .A(n_106), .Y(n_134) );
INVx1_ASAP7_75t_L g135 ( .A(n_81), .Y(n_135) );
HB1xp67_ASAP7_75t_L g136 ( .A(n_84), .Y(n_136) );
NAND2xp5_ASAP7_75t_L g137 ( .A(n_102), .B(n_2), .Y(n_137) );
INVx1_ASAP7_75t_L g138 ( .A(n_82), .Y(n_138) );
INVx1_ASAP7_75t_L g139 ( .A(n_82), .Y(n_139) );
BUFx6f_ASAP7_75t_L g140 ( .A(n_106), .Y(n_140) );
OAI21x1_ASAP7_75t_L g141 ( .A1(n_96), .A2(n_32), .B(n_76), .Y(n_141) );
INVx1_ASAP7_75t_L g142 ( .A(n_85), .Y(n_142) );
NAND2xp33_ASAP7_75t_SL g143 ( .A(n_99), .B(n_2), .Y(n_143) );
INVx2_ASAP7_75t_L g144 ( .A(n_106), .Y(n_144) );
INVx1_ASAP7_75t_L g145 ( .A(n_85), .Y(n_145) );
CKINVDCx8_ASAP7_75t_R g146 ( .A(n_101), .Y(n_146) );
INVx3_ASAP7_75t_L g147 ( .A(n_89), .Y(n_147) );
INVx2_ASAP7_75t_L g148 ( .A(n_106), .Y(n_148) );
INVx1_ASAP7_75t_SL g149 ( .A(n_83), .Y(n_149) );
INVx2_ASAP7_75t_L g150 ( .A(n_96), .Y(n_150) );
INVx1_ASAP7_75t_L g151 ( .A(n_89), .Y(n_151) );
NAND2xp5_ASAP7_75t_L g152 ( .A(n_103), .B(n_3), .Y(n_152) );
INVx1_ASAP7_75t_SL g153 ( .A(n_88), .Y(n_153) );
OA21x2_ASAP7_75t_L g154 ( .A1(n_98), .A2(n_39), .B(n_75), .Y(n_154) );
NAND2xp5_ASAP7_75t_L g155 ( .A(n_103), .B(n_3), .Y(n_155) );
AND2x4_ASAP7_75t_SL g156 ( .A(n_87), .B(n_29), .Y(n_156) );
INVxp67_ASAP7_75t_L g157 ( .A(n_87), .Y(n_157) );
INVx2_ASAP7_75t_L g158 ( .A(n_107), .Y(n_158) );
INVx1_ASAP7_75t_L g159 ( .A(n_98), .Y(n_159) );
INVx1_ASAP7_75t_L g160 ( .A(n_108), .Y(n_160) );
INVx1_ASAP7_75t_L g161 ( .A(n_108), .Y(n_161) );
INVx2_ASAP7_75t_L g162 ( .A(n_107), .Y(n_162) );
INVx2_ASAP7_75t_L g163 ( .A(n_109), .Y(n_163) );
OAI22xp5_ASAP7_75t_SL g164 ( .A1(n_123), .A2(n_5), .B1(n_7), .B2(n_10), .Y(n_164) );
INVx3_ASAP7_75t_L g165 ( .A(n_125), .Y(n_165) );
INVx2_ASAP7_75t_L g166 ( .A(n_109), .Y(n_166) );
INVx1_ASAP7_75t_L g167 ( .A(n_111), .Y(n_167) );
NOR2xp33_ASAP7_75t_L g168 ( .A(n_100), .B(n_125), .Y(n_168) );
BUFx2_ASAP7_75t_L g169 ( .A(n_80), .Y(n_169) );
AND2x2_ASAP7_75t_L g170 ( .A(n_169), .B(n_124), .Y(n_170) );
NAND2xp5_ASAP7_75t_L g171 ( .A(n_169), .B(n_86), .Y(n_171) );
NOR2xp33_ASAP7_75t_L g172 ( .A(n_157), .B(n_121), .Y(n_172) );
NAND2xp5_ASAP7_75t_SL g173 ( .A(n_128), .B(n_97), .Y(n_173) );
NAND2xp5_ASAP7_75t_L g174 ( .A(n_128), .B(n_118), .Y(n_174) );
NAND2xp5_ASAP7_75t_SL g175 ( .A(n_129), .B(n_93), .Y(n_175) );
INVx2_ASAP7_75t_SL g176 ( .A(n_136), .Y(n_176) );
BUFx6f_ASAP7_75t_SL g177 ( .A(n_132), .Y(n_177) );
NAND2xp5_ASAP7_75t_SL g178 ( .A(n_129), .B(n_114), .Y(n_178) );
INVx1_ASAP7_75t_L g179 ( .A(n_163), .Y(n_179) );
INVx1_ASAP7_75t_L g180 ( .A(n_163), .Y(n_180) );
NOR2xp33_ASAP7_75t_L g181 ( .A(n_168), .B(n_110), .Y(n_181) );
INVx1_ASAP7_75t_L g182 ( .A(n_163), .Y(n_182) );
OAI22xp5_ASAP7_75t_L g183 ( .A1(n_146), .A2(n_124), .B1(n_122), .B2(n_92), .Y(n_183) );
INVx1_ASAP7_75t_L g184 ( .A(n_166), .Y(n_184) );
NAND2xp5_ASAP7_75t_L g185 ( .A(n_131), .B(n_111), .Y(n_185) );
NAND2xp5_ASAP7_75t_SL g186 ( .A(n_131), .B(n_119), .Y(n_186) );
INVx2_ASAP7_75t_SL g187 ( .A(n_147), .Y(n_187) );
NAND3xp33_ASAP7_75t_L g188 ( .A(n_135), .B(n_112), .C(n_116), .Y(n_188) );
NAND2xp5_ASAP7_75t_SL g189 ( .A(n_135), .B(n_119), .Y(n_189) );
NAND2xp5_ASAP7_75t_L g190 ( .A(n_138), .B(n_112), .Y(n_190) );
NAND2xp5_ASAP7_75t_L g191 ( .A(n_138), .B(n_116), .Y(n_191) );
NAND2xp5_ASAP7_75t_L g192 ( .A(n_139), .B(n_110), .Y(n_192) );
INVx1_ASAP7_75t_L g193 ( .A(n_166), .Y(n_193) );
BUFx3_ASAP7_75t_L g194 ( .A(n_141), .Y(n_194) );
NAND2xp5_ASAP7_75t_SL g195 ( .A(n_139), .B(n_104), .Y(n_195) );
INVx1_ASAP7_75t_L g196 ( .A(n_166), .Y(n_196) );
NAND2xp5_ASAP7_75t_L g197 ( .A(n_142), .B(n_122), .Y(n_197) );
INVx3_ASAP7_75t_L g198 ( .A(n_132), .Y(n_198) );
INVx2_ASAP7_75t_L g199 ( .A(n_134), .Y(n_199) );
INVx1_ASAP7_75t_L g200 ( .A(n_147), .Y(n_200) );
NAND2x1p5_ASAP7_75t_L g201 ( .A(n_132), .B(n_95), .Y(n_201) );
NOR2xp33_ASAP7_75t_L g202 ( .A(n_146), .B(n_113), .Y(n_202) );
NAND2xp5_ASAP7_75t_L g203 ( .A(n_142), .B(n_90), .Y(n_203) );
AND2x4_ASAP7_75t_L g204 ( .A(n_132), .B(n_90), .Y(n_204) );
NOR2xp67_ASAP7_75t_L g205 ( .A(n_147), .B(n_165), .Y(n_205) );
AOI22xp33_ASAP7_75t_L g206 ( .A1(n_145), .A2(n_115), .B1(n_95), .B2(n_92), .Y(n_206) );
INVx2_ASAP7_75t_L g207 ( .A(n_134), .Y(n_207) );
NAND2xp5_ASAP7_75t_SL g208 ( .A(n_145), .B(n_120), .Y(n_208) );
AND2x2_ASAP7_75t_L g209 ( .A(n_151), .B(n_115), .Y(n_209) );
INVx4_ASAP7_75t_L g210 ( .A(n_156), .Y(n_210) );
BUFx3_ASAP7_75t_L g211 ( .A(n_141), .Y(n_211) );
NOR2xp33_ASAP7_75t_L g212 ( .A(n_151), .B(n_105), .Y(n_212) );
INVx2_ASAP7_75t_L g213 ( .A(n_134), .Y(n_213) );
AND2x4_ASAP7_75t_SL g214 ( .A(n_147), .B(n_94), .Y(n_214) );
NAND2xp5_ASAP7_75t_L g215 ( .A(n_159), .B(n_91), .Y(n_215) );
NOR2xp33_ASAP7_75t_L g216 ( .A(n_159), .B(n_40), .Y(n_216) );
INVx8_ASAP7_75t_L g217 ( .A(n_165), .Y(n_217) );
BUFx3_ASAP7_75t_L g218 ( .A(n_156), .Y(n_218) );
INVx1_ASAP7_75t_L g219 ( .A(n_165), .Y(n_219) );
NAND2xp5_ASAP7_75t_L g220 ( .A(n_160), .B(n_5), .Y(n_220) );
BUFx6f_ASAP7_75t_L g221 ( .A(n_127), .Y(n_221) );
BUFx3_ASAP7_75t_L g222 ( .A(n_156), .Y(n_222) );
NAND2xp5_ASAP7_75t_SL g223 ( .A(n_160), .B(n_41), .Y(n_223) );
AOI22xp33_ASAP7_75t_L g224 ( .A1(n_161), .A2(n_7), .B1(n_10), .B2(n_11), .Y(n_224) );
HB1xp67_ASAP7_75t_L g225 ( .A(n_149), .Y(n_225) );
INVx1_ASAP7_75t_L g226 ( .A(n_165), .Y(n_226) );
NAND2xp5_ASAP7_75t_L g227 ( .A(n_161), .B(n_12), .Y(n_227) );
NOR2x1p5_ASAP7_75t_L g228 ( .A(n_130), .B(n_14), .Y(n_228) );
INVx3_ASAP7_75t_L g229 ( .A(n_150), .Y(n_229) );
AOI22xp5_ASAP7_75t_L g230 ( .A1(n_176), .A2(n_143), .B1(n_164), .B2(n_167), .Y(n_230) );
NAND2xp5_ASAP7_75t_L g231 ( .A(n_176), .B(n_167), .Y(n_231) );
NOR2xp67_ASAP7_75t_L g232 ( .A(n_225), .B(n_162), .Y(n_232) );
INVx1_ASAP7_75t_L g233 ( .A(n_205), .Y(n_233) );
INVx1_ASAP7_75t_L g234 ( .A(n_205), .Y(n_234) );
INVx1_ASAP7_75t_L g235 ( .A(n_201), .Y(n_235) );
INVx2_ASAP7_75t_L g236 ( .A(n_179), .Y(n_236) );
NAND2xp5_ASAP7_75t_L g237 ( .A(n_172), .B(n_152), .Y(n_237) );
INVx2_ASAP7_75t_L g238 ( .A(n_179), .Y(n_238) );
BUFx2_ASAP7_75t_L g239 ( .A(n_218), .Y(n_239) );
NAND2xp5_ASAP7_75t_L g240 ( .A(n_174), .B(n_155), .Y(n_240) );
OR2x2_ASAP7_75t_L g241 ( .A(n_215), .B(n_153), .Y(n_241) );
BUFx6f_ASAP7_75t_L g242 ( .A(n_217), .Y(n_242) );
INVx1_ASAP7_75t_L g243 ( .A(n_201), .Y(n_243) );
NAND2xp5_ASAP7_75t_L g244 ( .A(n_217), .B(n_137), .Y(n_244) );
NAND2xp5_ASAP7_75t_L g245 ( .A(n_217), .B(n_162), .Y(n_245) );
INVx1_ASAP7_75t_L g246 ( .A(n_201), .Y(n_246) );
INVx2_ASAP7_75t_L g247 ( .A(n_180), .Y(n_247) );
NAND2xp5_ASAP7_75t_L g248 ( .A(n_217), .B(n_162), .Y(n_248) );
BUFx3_ASAP7_75t_L g249 ( .A(n_217), .Y(n_249) );
INVxp67_ASAP7_75t_L g250 ( .A(n_171), .Y(n_250) );
INVx5_ASAP7_75t_L g251 ( .A(n_198), .Y(n_251) );
INVx1_ASAP7_75t_L g252 ( .A(n_180), .Y(n_252) );
CKINVDCx14_ASAP7_75t_R g253 ( .A(n_210), .Y(n_253) );
NAND2xp5_ASAP7_75t_SL g254 ( .A(n_198), .B(n_158), .Y(n_254) );
AOI22xp5_ASAP7_75t_L g255 ( .A1(n_183), .A2(n_150), .B1(n_158), .B2(n_154), .Y(n_255) );
INVx2_ASAP7_75t_L g256 ( .A(n_182), .Y(n_256) );
CKINVDCx5p33_ASAP7_75t_R g257 ( .A(n_218), .Y(n_257) );
NOR2xp33_ASAP7_75t_L g258 ( .A(n_173), .B(n_158), .Y(n_258) );
NAND2xp5_ASAP7_75t_L g259 ( .A(n_170), .B(n_150), .Y(n_259) );
AOI21xp5_ASAP7_75t_L g260 ( .A1(n_198), .A2(n_154), .B(n_148), .Y(n_260) );
INVx1_ASAP7_75t_L g261 ( .A(n_182), .Y(n_261) );
INVx1_ASAP7_75t_L g262 ( .A(n_184), .Y(n_262) );
AND3x1_ASAP7_75t_SL g263 ( .A(n_228), .B(n_133), .C(n_15), .Y(n_263) );
INVx2_ASAP7_75t_L g264 ( .A(n_184), .Y(n_264) );
INVx1_ASAP7_75t_L g265 ( .A(n_193), .Y(n_265) );
NAND2xp5_ASAP7_75t_L g266 ( .A(n_170), .B(n_154), .Y(n_266) );
NAND2xp5_ASAP7_75t_L g267 ( .A(n_204), .B(n_154), .Y(n_267) );
INVx2_ASAP7_75t_L g268 ( .A(n_193), .Y(n_268) );
INVx2_ASAP7_75t_L g269 ( .A(n_196), .Y(n_269) );
AOI21xp5_ASAP7_75t_L g270 ( .A1(n_194), .A2(n_148), .B(n_144), .Y(n_270) );
BUFx2_ASAP7_75t_L g271 ( .A(n_222), .Y(n_271) );
INVx1_ASAP7_75t_L g272 ( .A(n_196), .Y(n_272) );
INVx1_ASAP7_75t_L g273 ( .A(n_209), .Y(n_273) );
INVx1_ASAP7_75t_L g274 ( .A(n_209), .Y(n_274) );
INVx1_ASAP7_75t_L g275 ( .A(n_200), .Y(n_275) );
CKINVDCx5p33_ASAP7_75t_R g276 ( .A(n_222), .Y(n_276) );
INVx1_ASAP7_75t_L g277 ( .A(n_200), .Y(n_277) );
BUFx12f_ASAP7_75t_L g278 ( .A(n_228), .Y(n_278) );
BUFx2_ASAP7_75t_L g279 ( .A(n_210), .Y(n_279) );
CKINVDCx20_ASAP7_75t_R g280 ( .A(n_214), .Y(n_280) );
NAND2xp5_ASAP7_75t_L g281 ( .A(n_204), .B(n_148), .Y(n_281) );
BUFx4f_ASAP7_75t_L g282 ( .A(n_204), .Y(n_282) );
HB1xp67_ASAP7_75t_L g283 ( .A(n_214), .Y(n_283) );
BUFx6f_ASAP7_75t_L g284 ( .A(n_194), .Y(n_284) );
INVx1_ASAP7_75t_L g285 ( .A(n_219), .Y(n_285) );
NAND2xp5_ASAP7_75t_L g286 ( .A(n_204), .B(n_144), .Y(n_286) );
HB1xp67_ASAP7_75t_L g287 ( .A(n_210), .Y(n_287) );
NOR2xp33_ASAP7_75t_L g288 ( .A(n_175), .B(n_144), .Y(n_288) );
INVx5_ASAP7_75t_L g289 ( .A(n_229), .Y(n_289) );
AND2x2_ASAP7_75t_L g290 ( .A(n_212), .B(n_133), .Y(n_290) );
INVx1_ASAP7_75t_L g291 ( .A(n_219), .Y(n_291) );
OR2x2_ASAP7_75t_L g292 ( .A(n_197), .B(n_14), .Y(n_292) );
NOR2xp67_ASAP7_75t_L g293 ( .A(n_188), .B(n_16), .Y(n_293) );
OAI21x1_ASAP7_75t_L g294 ( .A1(n_226), .A2(n_140), .B(n_127), .Y(n_294) );
INVx1_ASAP7_75t_L g295 ( .A(n_273), .Y(n_295) );
INVx1_ASAP7_75t_L g296 ( .A(n_274), .Y(n_296) );
BUFx2_ASAP7_75t_L g297 ( .A(n_249), .Y(n_297) );
BUFx3_ASAP7_75t_L g298 ( .A(n_242), .Y(n_298) );
INVx1_ASAP7_75t_L g299 ( .A(n_231), .Y(n_299) );
INVx1_ASAP7_75t_L g300 ( .A(n_236), .Y(n_300) );
AOI22xp5_ASAP7_75t_L g301 ( .A1(n_235), .A2(n_177), .B1(n_202), .B2(n_195), .Y(n_301) );
NAND2xp5_ASAP7_75t_L g302 ( .A(n_250), .B(n_208), .Y(n_302) );
AOI21xp5_ASAP7_75t_L g303 ( .A1(n_267), .A2(n_211), .B(n_187), .Y(n_303) );
NAND2xp5_ASAP7_75t_L g304 ( .A(n_232), .B(n_187), .Y(n_304) );
INVx2_ASAP7_75t_L g305 ( .A(n_236), .Y(n_305) );
INVx2_ASAP7_75t_SL g306 ( .A(n_249), .Y(n_306) );
INVx1_ASAP7_75t_L g307 ( .A(n_238), .Y(n_307) );
AOI21xp5_ASAP7_75t_L g308 ( .A1(n_266), .A2(n_211), .B(n_226), .Y(n_308) );
O2A1O1Ixp33_ASAP7_75t_L g309 ( .A1(n_259), .A2(n_220), .B(n_227), .C(n_189), .Y(n_309) );
OAI22xp5_ASAP7_75t_L g310 ( .A1(n_282), .A2(n_177), .B1(n_224), .B2(n_206), .Y(n_310) );
AOI21xp5_ASAP7_75t_L g311 ( .A1(n_270), .A2(n_178), .B(n_186), .Y(n_311) );
BUFx3_ASAP7_75t_L g312 ( .A(n_242), .Y(n_312) );
BUFx2_ASAP7_75t_L g313 ( .A(n_282), .Y(n_313) );
CKINVDCx5p33_ASAP7_75t_R g314 ( .A(n_253), .Y(n_314) );
AOI21x1_ASAP7_75t_L g315 ( .A1(n_260), .A2(n_185), .B(n_190), .Y(n_315) );
OR2x6_ASAP7_75t_SL g316 ( .A(n_257), .B(n_177), .Y(n_316) );
INVx2_ASAP7_75t_L g317 ( .A(n_238), .Y(n_317) );
AOI21xp5_ASAP7_75t_L g318 ( .A1(n_240), .A2(n_192), .B(n_191), .Y(n_318) );
INVx1_ASAP7_75t_L g319 ( .A(n_247), .Y(n_319) );
INVx3_ASAP7_75t_SL g320 ( .A(n_280), .Y(n_320) );
OA21x2_ASAP7_75t_L g321 ( .A1(n_294), .A2(n_188), .B(n_216), .Y(n_321) );
AND2x4_ASAP7_75t_L g322 ( .A(n_243), .B(n_203), .Y(n_322) );
AOI21xp5_ASAP7_75t_L g323 ( .A1(n_254), .A2(n_181), .B(n_223), .Y(n_323) );
INVx3_ASAP7_75t_L g324 ( .A(n_242), .Y(n_324) );
AOI21xp5_ASAP7_75t_L g325 ( .A1(n_254), .A2(n_244), .B(n_282), .Y(n_325) );
AOI21xp5_ASAP7_75t_L g326 ( .A1(n_275), .A2(n_229), .B(n_213), .Y(n_326) );
AND2x2_ASAP7_75t_L g327 ( .A(n_246), .B(n_229), .Y(n_327) );
AOI21xp5_ASAP7_75t_L g328 ( .A1(n_277), .A2(n_213), .B(n_207), .Y(n_328) );
AOI21xp5_ASAP7_75t_L g329 ( .A1(n_285), .A2(n_207), .B(n_199), .Y(n_329) );
AOI21xp5_ASAP7_75t_L g330 ( .A1(n_291), .A2(n_199), .B(n_221), .Y(n_330) );
AOI21xp5_ASAP7_75t_L g331 ( .A1(n_245), .A2(n_221), .B(n_140), .Y(n_331) );
AND2x2_ASAP7_75t_L g332 ( .A(n_241), .B(n_16), .Y(n_332) );
OAI22xp33_ASAP7_75t_L g333 ( .A1(n_280), .A2(n_241), .B1(n_230), .B2(n_292), .Y(n_333) );
NAND2xp5_ASAP7_75t_L g334 ( .A(n_237), .B(n_17), .Y(n_334) );
BUFx2_ASAP7_75t_L g335 ( .A(n_242), .Y(n_335) );
CKINVDCx5p33_ASAP7_75t_R g336 ( .A(n_253), .Y(n_336) );
O2A1O1Ixp33_ASAP7_75t_L g337 ( .A1(n_292), .A2(n_17), .B(n_18), .C(n_19), .Y(n_337) );
AND2x2_ASAP7_75t_L g338 ( .A(n_247), .B(n_18), .Y(n_338) );
NOR2xp67_ASAP7_75t_L g339 ( .A(n_278), .B(n_21), .Y(n_339) );
BUFx2_ASAP7_75t_L g340 ( .A(n_257), .Y(n_340) );
AND2x2_ASAP7_75t_L g341 ( .A(n_256), .B(n_140), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g342 ( .A(n_256), .B(n_140), .Y(n_342) );
CKINVDCx6p67_ASAP7_75t_R g343 ( .A(n_283), .Y(n_343) );
BUFx6f_ASAP7_75t_L g344 ( .A(n_284), .Y(n_344) );
AOI21xp5_ASAP7_75t_L g345 ( .A1(n_248), .A2(n_221), .B(n_140), .Y(n_345) );
INVx2_ASAP7_75t_L g346 ( .A(n_305), .Y(n_346) );
CKINVDCx5p33_ASAP7_75t_R g347 ( .A(n_320), .Y(n_347) );
INVx1_ASAP7_75t_L g348 ( .A(n_305), .Y(n_348) );
INVx1_ASAP7_75t_L g349 ( .A(n_317), .Y(n_349) );
INVx2_ASAP7_75t_L g350 ( .A(n_317), .Y(n_350) );
INVx2_ASAP7_75t_L g351 ( .A(n_315), .Y(n_351) );
INVx2_ASAP7_75t_L g352 ( .A(n_344), .Y(n_352) );
BUFx3_ASAP7_75t_L g353 ( .A(n_298), .Y(n_353) );
INVx1_ASAP7_75t_L g354 ( .A(n_300), .Y(n_354) );
AOI21xp5_ASAP7_75t_L g355 ( .A1(n_308), .A2(n_284), .B(n_286), .Y(n_355) );
INVx1_ASAP7_75t_L g356 ( .A(n_307), .Y(n_356) );
AOI221xp5_ASAP7_75t_L g357 ( .A1(n_333), .A2(n_290), .B1(n_258), .B2(n_233), .C(n_234), .Y(n_357) );
INVx2_ASAP7_75t_L g358 ( .A(n_344), .Y(n_358) );
OAI21x1_ASAP7_75t_L g359 ( .A1(n_303), .A2(n_294), .B(n_255), .Y(n_359) );
INVx2_ASAP7_75t_L g360 ( .A(n_344), .Y(n_360) );
AND2x2_ASAP7_75t_L g361 ( .A(n_299), .B(n_264), .Y(n_361) );
AND2x2_ASAP7_75t_L g362 ( .A(n_322), .B(n_264), .Y(n_362) );
AO21x1_ASAP7_75t_SL g363 ( .A1(n_319), .A2(n_265), .B(n_252), .Y(n_363) );
INVx1_ASAP7_75t_L g364 ( .A(n_338), .Y(n_364) );
INVx2_ASAP7_75t_L g365 ( .A(n_344), .Y(n_365) );
BUFx6f_ASAP7_75t_L g366 ( .A(n_298), .Y(n_366) );
BUFx2_ASAP7_75t_L g367 ( .A(n_297), .Y(n_367) );
HB1xp67_ASAP7_75t_L g368 ( .A(n_297), .Y(n_368) );
INVx1_ASAP7_75t_L g369 ( .A(n_338), .Y(n_369) );
INVx1_ASAP7_75t_L g370 ( .A(n_295), .Y(n_370) );
AND2x2_ASAP7_75t_SL g371 ( .A(n_332), .B(n_284), .Y(n_371) );
INVx2_ASAP7_75t_L g372 ( .A(n_341), .Y(n_372) );
INVx2_ASAP7_75t_L g373 ( .A(n_341), .Y(n_373) );
OR2x2_ASAP7_75t_L g374 ( .A(n_320), .B(n_290), .Y(n_374) );
INVx1_ASAP7_75t_L g375 ( .A(n_296), .Y(n_375) );
CKINVDCx5p33_ASAP7_75t_R g376 ( .A(n_314), .Y(n_376) );
AO21x2_ASAP7_75t_L g377 ( .A1(n_323), .A2(n_293), .B(n_261), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_348), .Y(n_378) );
INVx1_ASAP7_75t_L g379 ( .A(n_348), .Y(n_379) );
INVx1_ASAP7_75t_L g380 ( .A(n_349), .Y(n_380) );
BUFx2_ASAP7_75t_L g381 ( .A(n_367), .Y(n_381) );
BUFx2_ASAP7_75t_L g382 ( .A(n_367), .Y(n_382) );
AND2x4_ASAP7_75t_L g383 ( .A(n_362), .B(n_327), .Y(n_383) );
NOR2x1_ASAP7_75t_SL g384 ( .A(n_363), .B(n_284), .Y(n_384) );
AND2x2_ASAP7_75t_L g385 ( .A(n_361), .B(n_322), .Y(n_385) );
INVxp67_ASAP7_75t_SL g386 ( .A(n_351), .Y(n_386) );
INVx1_ASAP7_75t_L g387 ( .A(n_349), .Y(n_387) );
INVx2_ASAP7_75t_L g388 ( .A(n_351), .Y(n_388) );
INVx1_ASAP7_75t_L g389 ( .A(n_361), .Y(n_389) );
INVx1_ASAP7_75t_L g390 ( .A(n_346), .Y(n_390) );
AND2x2_ASAP7_75t_L g391 ( .A(n_362), .B(n_322), .Y(n_391) );
INVx2_ASAP7_75t_SL g392 ( .A(n_366), .Y(n_392) );
INVx1_ASAP7_75t_L g393 ( .A(n_346), .Y(n_393) );
NAND2xp5_ASAP7_75t_L g394 ( .A(n_364), .B(n_332), .Y(n_394) );
INVx2_ASAP7_75t_L g395 ( .A(n_351), .Y(n_395) );
AND2x2_ASAP7_75t_L g396 ( .A(n_354), .B(n_327), .Y(n_396) );
INVx1_ASAP7_75t_L g397 ( .A(n_346), .Y(n_397) );
AND2x4_ASAP7_75t_L g398 ( .A(n_354), .B(n_312), .Y(n_398) );
INVx1_ASAP7_75t_L g399 ( .A(n_350), .Y(n_399) );
HB1xp67_ASAP7_75t_L g400 ( .A(n_368), .Y(n_400) );
INVx1_ASAP7_75t_L g401 ( .A(n_350), .Y(n_401) );
NAND2xp5_ASAP7_75t_L g402 ( .A(n_364), .B(n_318), .Y(n_402) );
INVxp67_ASAP7_75t_SL g403 ( .A(n_350), .Y(n_403) );
BUFx2_ASAP7_75t_L g404 ( .A(n_368), .Y(n_404) );
OR2x2_ASAP7_75t_L g405 ( .A(n_356), .B(n_370), .Y(n_405) );
BUFx3_ASAP7_75t_L g406 ( .A(n_381), .Y(n_406) );
NOR3xp33_ASAP7_75t_L g407 ( .A(n_400), .B(n_357), .C(n_337), .Y(n_407) );
INVx2_ASAP7_75t_L g408 ( .A(n_390), .Y(n_408) );
BUFx2_ASAP7_75t_SL g409 ( .A(n_403), .Y(n_409) );
INVx3_ASAP7_75t_L g410 ( .A(n_398), .Y(n_410) );
BUFx2_ASAP7_75t_L g411 ( .A(n_403), .Y(n_411) );
OR2x2_ASAP7_75t_L g412 ( .A(n_381), .B(n_356), .Y(n_412) );
NAND2xp5_ASAP7_75t_L g413 ( .A(n_385), .B(n_357), .Y(n_413) );
INVx1_ASAP7_75t_SL g414 ( .A(n_382), .Y(n_414) );
OAI322xp33_ASAP7_75t_L g415 ( .A1(n_405), .A2(n_374), .A3(n_334), .B1(n_370), .B2(n_375), .C1(n_258), .C2(n_369), .Y(n_415) );
INVx1_ASAP7_75t_L g416 ( .A(n_378), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_378), .Y(n_417) );
NAND2xp5_ASAP7_75t_L g418 ( .A(n_385), .B(n_375), .Y(n_418) );
AOI221xp5_ASAP7_75t_L g419 ( .A1(n_394), .A2(n_302), .B1(n_374), .B2(n_340), .C(n_369), .Y(n_419) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_396), .B(n_340), .Y(n_420) );
INVx1_ASAP7_75t_L g421 ( .A(n_379), .Y(n_421) );
NAND2xp5_ASAP7_75t_L g422 ( .A(n_396), .B(n_343), .Y(n_422) );
OAI222xp33_ASAP7_75t_L g423 ( .A1(n_382), .A2(n_347), .B1(n_314), .B2(n_336), .C1(n_276), .C2(n_310), .Y(n_423) );
AOI221xp5_ASAP7_75t_SL g424 ( .A1(n_404), .A2(n_304), .B1(n_309), .B2(n_311), .C(n_288), .Y(n_424) );
INVx1_ASAP7_75t_L g425 ( .A(n_379), .Y(n_425) );
HB1xp67_ASAP7_75t_L g426 ( .A(n_404), .Y(n_426) );
AOI22xp33_ASAP7_75t_SL g427 ( .A1(n_384), .A2(n_371), .B1(n_336), .B2(n_276), .Y(n_427) );
NOR2x1_ASAP7_75t_L g428 ( .A(n_405), .B(n_339), .Y(n_428) );
INVx1_ASAP7_75t_L g429 ( .A(n_380), .Y(n_429) );
AO21x2_ASAP7_75t_L g430 ( .A1(n_386), .A2(n_359), .B(n_377), .Y(n_430) );
AO21x2_ASAP7_75t_L g431 ( .A1(n_386), .A2(n_359), .B(n_377), .Y(n_431) );
AOI22xp33_ASAP7_75t_L g432 ( .A1(n_383), .A2(n_371), .B1(n_363), .B2(n_278), .Y(n_432) );
INVx1_ASAP7_75t_L g433 ( .A(n_380), .Y(n_433) );
OAI33xp33_ASAP7_75t_L g434 ( .A1(n_402), .A2(n_263), .A3(n_376), .B1(n_281), .B2(n_272), .B3(n_262), .Y(n_434) );
INVx1_ASAP7_75t_SL g435 ( .A(n_391), .Y(n_435) );
INVx3_ASAP7_75t_L g436 ( .A(n_398), .Y(n_436) );
OAI22xp5_ASAP7_75t_L g437 ( .A1(n_394), .A2(n_371), .B1(n_316), .B2(n_372), .Y(n_437) );
NOR2xp33_ASAP7_75t_L g438 ( .A(n_391), .B(n_343), .Y(n_438) );
NAND4xp25_ASAP7_75t_L g439 ( .A(n_402), .B(n_288), .C(n_301), .D(n_271), .Y(n_439) );
OAI33xp33_ASAP7_75t_L g440 ( .A1(n_387), .A2(n_342), .A3(n_373), .B1(n_372), .B2(n_268), .B3(n_269), .Y(n_440) );
INVx1_ASAP7_75t_L g441 ( .A(n_416), .Y(n_441) );
INVx1_ASAP7_75t_L g442 ( .A(n_416), .Y(n_442) );
NOR3xp33_ASAP7_75t_L g443 ( .A(n_434), .B(n_389), .C(n_387), .Y(n_443) );
NAND2xp5_ASAP7_75t_L g444 ( .A(n_413), .B(n_389), .Y(n_444) );
AND2x2_ASAP7_75t_L g445 ( .A(n_408), .B(n_390), .Y(n_445) );
NAND2xp5_ASAP7_75t_L g446 ( .A(n_418), .B(n_401), .Y(n_446) );
INVx1_ASAP7_75t_L g447 ( .A(n_417), .Y(n_447) );
INVx2_ASAP7_75t_L g448 ( .A(n_408), .Y(n_448) );
NAND2xp5_ASAP7_75t_L g449 ( .A(n_435), .B(n_401), .Y(n_449) );
INVx1_ASAP7_75t_L g450 ( .A(n_417), .Y(n_450) );
INVx2_ASAP7_75t_L g451 ( .A(n_411), .Y(n_451) );
OR2x2_ASAP7_75t_L g452 ( .A(n_411), .B(n_395), .Y(n_452) );
INVx1_ASAP7_75t_L g453 ( .A(n_421), .Y(n_453) );
INVx2_ASAP7_75t_L g454 ( .A(n_421), .Y(n_454) );
INVxp67_ASAP7_75t_L g455 ( .A(n_409), .Y(n_455) );
AND2x4_ASAP7_75t_L g456 ( .A(n_410), .B(n_384), .Y(n_456) );
INVx1_ASAP7_75t_L g457 ( .A(n_425), .Y(n_457) );
OAI21xp5_ASAP7_75t_L g458 ( .A1(n_407), .A2(n_399), .B(n_393), .Y(n_458) );
INVx2_ASAP7_75t_L g459 ( .A(n_425), .Y(n_459) );
INVx1_ASAP7_75t_L g460 ( .A(n_429), .Y(n_460) );
OAI21xp33_ASAP7_75t_SL g461 ( .A1(n_432), .A2(n_399), .B(n_397), .Y(n_461) );
INVx3_ASAP7_75t_L g462 ( .A(n_410), .Y(n_462) );
INVx1_ASAP7_75t_L g463 ( .A(n_429), .Y(n_463) );
OR2x2_ASAP7_75t_L g464 ( .A(n_409), .B(n_395), .Y(n_464) );
AND2x2_ASAP7_75t_L g465 ( .A(n_433), .B(n_397), .Y(n_465) );
INVx1_ASAP7_75t_L g466 ( .A(n_433), .Y(n_466) );
BUFx3_ASAP7_75t_L g467 ( .A(n_406), .Y(n_467) );
NAND4xp25_ASAP7_75t_L g468 ( .A(n_419), .B(n_383), .C(n_398), .D(n_325), .Y(n_468) );
OAI21xp33_ASAP7_75t_SL g469 ( .A1(n_428), .A2(n_393), .B(n_392), .Y(n_469) );
AND2x4_ASAP7_75t_L g470 ( .A(n_410), .B(n_395), .Y(n_470) );
NAND2xp5_ASAP7_75t_R g471 ( .A(n_438), .B(n_392), .Y(n_471) );
OR2x2_ASAP7_75t_L g472 ( .A(n_414), .B(n_388), .Y(n_472) );
INVx1_ASAP7_75t_L g473 ( .A(n_412), .Y(n_473) );
AND2x4_ASAP7_75t_L g474 ( .A(n_436), .B(n_388), .Y(n_474) );
AND2x2_ASAP7_75t_L g475 ( .A(n_436), .B(n_388), .Y(n_475) );
AND2x2_ASAP7_75t_L g476 ( .A(n_436), .B(n_383), .Y(n_476) );
AND2x2_ASAP7_75t_L g477 ( .A(n_406), .B(n_383), .Y(n_477) );
OR2x2_ASAP7_75t_L g478 ( .A(n_412), .B(n_398), .Y(n_478) );
INVx1_ASAP7_75t_L g479 ( .A(n_426), .Y(n_479) );
INVx2_ASAP7_75t_L g480 ( .A(n_430), .Y(n_480) );
NAND2xp5_ASAP7_75t_L g481 ( .A(n_420), .B(n_373), .Y(n_481) );
INVx1_ASAP7_75t_L g482 ( .A(n_422), .Y(n_482) );
NAND2xp5_ASAP7_75t_L g483 ( .A(n_437), .B(n_373), .Y(n_483) );
NAND2xp5_ASAP7_75t_L g484 ( .A(n_439), .B(n_372), .Y(n_484) );
AOI21xp5_ASAP7_75t_L g485 ( .A1(n_440), .A2(n_392), .B(n_377), .Y(n_485) );
INVx1_ASAP7_75t_L g486 ( .A(n_415), .Y(n_486) );
NAND2xp5_ASAP7_75t_L g487 ( .A(n_427), .B(n_316), .Y(n_487) );
INVx1_ASAP7_75t_L g488 ( .A(n_430), .Y(n_488) );
INVx1_ASAP7_75t_L g489 ( .A(n_430), .Y(n_489) );
INVx1_ASAP7_75t_SL g490 ( .A(n_467), .Y(n_490) );
INVx1_ASAP7_75t_L g491 ( .A(n_441), .Y(n_491) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_473), .B(n_431), .Y(n_492) );
AND4x1_ASAP7_75t_L g493 ( .A(n_487), .B(n_423), .C(n_331), .D(n_345), .Y(n_493) );
NOR2x1_ASAP7_75t_SL g494 ( .A(n_464), .B(n_431), .Y(n_494) );
INVxp67_ASAP7_75t_L g495 ( .A(n_467), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_482), .B(n_431), .Y(n_496) );
INVx1_ASAP7_75t_L g497 ( .A(n_441), .Y(n_497) );
INVx1_ASAP7_75t_L g498 ( .A(n_454), .Y(n_498) );
INVx1_ASAP7_75t_L g499 ( .A(n_454), .Y(n_499) );
NOR2xp33_ASAP7_75t_L g500 ( .A(n_479), .B(n_239), .Y(n_500) );
BUFx2_ASAP7_75t_L g501 ( .A(n_455), .Y(n_501) );
INVx1_ASAP7_75t_L g502 ( .A(n_459), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_486), .B(n_424), .Y(n_503) );
NAND2xp5_ASAP7_75t_L g504 ( .A(n_444), .B(n_377), .Y(n_504) );
AND2x2_ASAP7_75t_L g505 ( .A(n_459), .B(n_127), .Y(n_505) );
CKINVDCx16_ASAP7_75t_R g506 ( .A(n_477), .Y(n_506) );
INVx1_ASAP7_75t_L g507 ( .A(n_442), .Y(n_507) );
INVx1_ASAP7_75t_L g508 ( .A(n_447), .Y(n_508) );
AND2x2_ASAP7_75t_L g509 ( .A(n_475), .B(n_127), .Y(n_509) );
AND2x2_ASAP7_75t_L g510 ( .A(n_475), .B(n_127), .Y(n_510) );
INVx1_ASAP7_75t_L g511 ( .A(n_450), .Y(n_511) );
AND2x2_ASAP7_75t_L g512 ( .A(n_448), .B(n_127), .Y(n_512) );
INVx1_ASAP7_75t_L g513 ( .A(n_453), .Y(n_513) );
NOR2xp33_ASAP7_75t_L g514 ( .A(n_481), .B(n_313), .Y(n_514) );
INVx1_ASAP7_75t_L g515 ( .A(n_457), .Y(n_515) );
INVxp67_ASAP7_75t_SL g516 ( .A(n_464), .Y(n_516) );
AND2x2_ASAP7_75t_L g517 ( .A(n_448), .B(n_140), .Y(n_517) );
CKINVDCx16_ASAP7_75t_R g518 ( .A(n_477), .Y(n_518) );
INVx2_ASAP7_75t_L g519 ( .A(n_452), .Y(n_519) );
NOR3xp33_ASAP7_75t_L g520 ( .A(n_484), .B(n_324), .C(n_313), .Y(n_520) );
INVx2_ASAP7_75t_L g521 ( .A(n_452), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_465), .B(n_353), .Y(n_522) );
NOR2xp33_ASAP7_75t_L g523 ( .A(n_478), .B(n_353), .Y(n_523) );
INVx1_ASAP7_75t_L g524 ( .A(n_460), .Y(n_524) );
OR2x2_ASAP7_75t_L g525 ( .A(n_451), .B(n_359), .Y(n_525) );
AND2x2_ASAP7_75t_L g526 ( .A(n_463), .B(n_365), .Y(n_526) );
INVx1_ASAP7_75t_L g527 ( .A(n_466), .Y(n_527) );
INVx1_ASAP7_75t_SL g528 ( .A(n_472), .Y(n_528) );
AND2x2_ASAP7_75t_L g529 ( .A(n_451), .B(n_365), .Y(n_529) );
INVx1_ASAP7_75t_L g530 ( .A(n_465), .Y(n_530) );
AND2x2_ASAP7_75t_L g531 ( .A(n_488), .B(n_365), .Y(n_531) );
INVx2_ASAP7_75t_L g532 ( .A(n_445), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_445), .B(n_353), .Y(n_533) );
NOR2xp33_ASAP7_75t_L g534 ( .A(n_478), .B(n_289), .Y(n_534) );
AOI22xp33_ASAP7_75t_L g535 ( .A1(n_468), .A2(n_366), .B1(n_335), .B2(n_358), .Y(n_535) );
HB1xp67_ASAP7_75t_L g536 ( .A(n_472), .Y(n_536) );
AND2x2_ASAP7_75t_L g537 ( .A(n_489), .B(n_360), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_446), .B(n_449), .Y(n_538) );
INVx1_ASAP7_75t_L g539 ( .A(n_480), .Y(n_539) );
AND2x2_ASAP7_75t_L g540 ( .A(n_470), .B(n_360), .Y(n_540) );
NOR2xp33_ASAP7_75t_L g541 ( .A(n_476), .B(n_289), .Y(n_541) );
INVx1_ASAP7_75t_L g542 ( .A(n_480), .Y(n_542) );
AND2x2_ASAP7_75t_L g543 ( .A(n_470), .B(n_360), .Y(n_543) );
INVx1_ASAP7_75t_L g544 ( .A(n_470), .Y(n_544) );
INVx2_ASAP7_75t_SL g545 ( .A(n_456), .Y(n_545) );
INVx1_ASAP7_75t_L g546 ( .A(n_458), .Y(n_546) );
AND2x2_ASAP7_75t_L g547 ( .A(n_474), .B(n_476), .Y(n_547) );
INVx1_ASAP7_75t_L g548 ( .A(n_497), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g549 ( .A(n_530), .B(n_483), .Y(n_549) );
OAI21xp5_ASAP7_75t_SL g550 ( .A1(n_535), .A2(n_456), .B(n_471), .Y(n_550) );
INVx1_ASAP7_75t_L g551 ( .A(n_497), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g552 ( .A(n_506), .B(n_443), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_518), .B(n_462), .Y(n_553) );
OAI211xp5_ASAP7_75t_L g554 ( .A1(n_503), .A2(n_469), .B(n_461), .C(n_462), .Y(n_554) );
INVx1_ASAP7_75t_L g555 ( .A(n_507), .Y(n_555) );
INVx1_ASAP7_75t_L g556 ( .A(n_507), .Y(n_556) );
INVx1_ASAP7_75t_SL g557 ( .A(n_490), .Y(n_557) );
INVx1_ASAP7_75t_L g558 ( .A(n_508), .Y(n_558) );
INVx1_ASAP7_75t_L g559 ( .A(n_508), .Y(n_559) );
OAI21xp33_ASAP7_75t_L g560 ( .A1(n_496), .A2(n_471), .B(n_485), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_536), .B(n_462), .Y(n_561) );
NAND2x1p5_ASAP7_75t_L g562 ( .A(n_501), .B(n_456), .Y(n_562) );
NAND2xp5_ASAP7_75t_SL g563 ( .A(n_495), .B(n_474), .Y(n_563) );
INVx2_ASAP7_75t_L g564 ( .A(n_498), .Y(n_564) );
INVx2_ASAP7_75t_L g565 ( .A(n_498), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g566 ( .A(n_538), .B(n_474), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_528), .B(n_366), .Y(n_567) );
INVx1_ASAP7_75t_L g568 ( .A(n_511), .Y(n_568) );
INVx1_ASAP7_75t_L g569 ( .A(n_511), .Y(n_569) );
NOR2xp33_ASAP7_75t_L g570 ( .A(n_501), .B(n_366), .Y(n_570) );
NAND2xp5_ASAP7_75t_L g571 ( .A(n_532), .B(n_366), .Y(n_571) );
INVxp67_ASAP7_75t_SL g572 ( .A(n_494), .Y(n_572) );
AND2x2_ASAP7_75t_L g573 ( .A(n_547), .B(n_532), .Y(n_573) );
OR2x2_ASAP7_75t_L g574 ( .A(n_516), .B(n_366), .Y(n_574) );
NOR2xp33_ASAP7_75t_L g575 ( .A(n_546), .B(n_22), .Y(n_575) );
AND2x2_ASAP7_75t_L g576 ( .A(n_547), .B(n_358), .Y(n_576) );
INVx1_ASAP7_75t_L g577 ( .A(n_513), .Y(n_577) );
XNOR2xp5_ASAP7_75t_L g578 ( .A(n_493), .B(n_287), .Y(n_578) );
INVx1_ASAP7_75t_L g579 ( .A(n_513), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g580 ( .A(n_527), .B(n_355), .Y(n_580) );
NAND2xp5_ASAP7_75t_L g581 ( .A(n_515), .B(n_355), .Y(n_581) );
INVx1_ASAP7_75t_L g582 ( .A(n_515), .Y(n_582) );
INVx1_ASAP7_75t_L g583 ( .A(n_524), .Y(n_583) );
INVx1_ASAP7_75t_L g584 ( .A(n_524), .Y(n_584) );
INVx1_ASAP7_75t_L g585 ( .A(n_491), .Y(n_585) );
NAND2x1p5_ASAP7_75t_L g586 ( .A(n_509), .B(n_312), .Y(n_586) );
BUFx2_ASAP7_75t_L g587 ( .A(n_545), .Y(n_587) );
INVx1_ASAP7_75t_L g588 ( .A(n_499), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g589 ( .A(n_519), .B(n_358), .Y(n_589) );
INVxp67_ASAP7_75t_L g590 ( .A(n_494), .Y(n_590) );
INVx1_ASAP7_75t_L g591 ( .A(n_499), .Y(n_591) );
INVx1_ASAP7_75t_L g592 ( .A(n_502), .Y(n_592) );
INVx1_ASAP7_75t_L g593 ( .A(n_502), .Y(n_593) );
NOR2xp33_ASAP7_75t_SL g594 ( .A(n_545), .B(n_352), .Y(n_594) );
INVx2_ASAP7_75t_L g595 ( .A(n_539), .Y(n_595) );
INVx1_ASAP7_75t_L g596 ( .A(n_519), .Y(n_596) );
NOR2xp33_ASAP7_75t_L g597 ( .A(n_500), .B(n_23), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g598 ( .A(n_521), .B(n_352), .Y(n_598) );
OAI21xp5_ASAP7_75t_L g599 ( .A1(n_520), .A2(n_335), .B(n_269), .Y(n_599) );
INVx1_ASAP7_75t_L g600 ( .A(n_521), .Y(n_600) );
NOR3xp33_ASAP7_75t_L g601 ( .A(n_597), .B(n_541), .C(n_534), .Y(n_601) );
NOR2xp67_ASAP7_75t_L g602 ( .A(n_590), .B(n_492), .Y(n_602) );
INVx1_ASAP7_75t_L g603 ( .A(n_555), .Y(n_603) );
NOR2xp33_ASAP7_75t_L g604 ( .A(n_557), .B(n_504), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g605 ( .A(n_549), .B(n_510), .Y(n_605) );
NOR3xp33_ASAP7_75t_L g606 ( .A(n_597), .B(n_509), .C(n_510), .Y(n_606) );
AOI221x1_ASAP7_75t_L g607 ( .A1(n_560), .A2(n_539), .B1(n_542), .B2(n_505), .C(n_544), .Y(n_607) );
AND2x2_ASAP7_75t_L g608 ( .A(n_573), .B(n_544), .Y(n_608) );
NAND4xp25_ASAP7_75t_SL g609 ( .A(n_554), .B(n_522), .C(n_533), .D(n_540), .Y(n_609) );
NOR2x1_ASAP7_75t_L g610 ( .A(n_550), .B(n_542), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g611 ( .A(n_566), .B(n_526), .Y(n_611) );
O2A1O1Ixp5_ASAP7_75t_L g612 ( .A1(n_572), .A2(n_523), .B(n_514), .C(n_526), .Y(n_612) );
OAI21xp33_ASAP7_75t_SL g613 ( .A1(n_572), .A2(n_543), .B(n_540), .Y(n_613) );
AND2x2_ASAP7_75t_L g614 ( .A(n_587), .B(n_543), .Y(n_614) );
NAND3xp33_ASAP7_75t_SL g615 ( .A(n_562), .B(n_505), .C(n_517), .Y(n_615) );
NOR3xp33_ASAP7_75t_L g616 ( .A(n_575), .B(n_517), .C(n_512), .Y(n_616) );
NOR3x1_ASAP7_75t_L g617 ( .A(n_552), .B(n_525), .C(n_306), .Y(n_617) );
OR2x2_ASAP7_75t_L g618 ( .A(n_596), .B(n_525), .Y(n_618) );
AND2x2_ASAP7_75t_L g619 ( .A(n_576), .B(n_537), .Y(n_619) );
AOI22xp5_ASAP7_75t_L g620 ( .A1(n_578), .A2(n_531), .B1(n_537), .B2(n_529), .Y(n_620) );
AND2x4_ASAP7_75t_L g621 ( .A(n_590), .B(n_531), .Y(n_621) );
AOI221x1_ASAP7_75t_L g622 ( .A1(n_575), .A2(n_512), .B1(n_529), .B2(n_352), .C(n_330), .Y(n_622) );
NAND2xp5_ASAP7_75t_SL g623 ( .A(n_562), .B(n_594), .Y(n_623) );
HB1xp67_ASAP7_75t_L g624 ( .A(n_595), .Y(n_624) );
AOI21xp33_ASAP7_75t_SL g625 ( .A1(n_563), .A2(n_553), .B(n_586), .Y(n_625) );
INVx1_ASAP7_75t_L g626 ( .A(n_556), .Y(n_626) );
NAND2xp5_ASAP7_75t_L g627 ( .A(n_600), .B(n_268), .Y(n_627) );
CKINVDCx20_ASAP7_75t_R g628 ( .A(n_561), .Y(n_628) );
OAI21xp5_ASAP7_75t_SL g629 ( .A1(n_563), .A2(n_599), .B(n_586), .Y(n_629) );
NOR2xp33_ASAP7_75t_L g630 ( .A(n_585), .B(n_25), .Y(n_630) );
HB1xp67_ASAP7_75t_L g631 ( .A(n_595), .Y(n_631) );
AND2x2_ASAP7_75t_L g632 ( .A(n_558), .B(n_28), .Y(n_632) );
NOR2x1_ASAP7_75t_L g633 ( .A(n_570), .B(n_324), .Y(n_633) );
XNOR2xp5_ASAP7_75t_L g634 ( .A(n_559), .B(n_324), .Y(n_634) );
NAND2xp5_ASAP7_75t_L g635 ( .A(n_568), .B(n_44), .Y(n_635) );
INVx1_ASAP7_75t_L g636 ( .A(n_569), .Y(n_636) );
NAND4xp25_ASAP7_75t_L g637 ( .A(n_570), .B(n_279), .C(n_326), .D(n_328), .Y(n_637) );
NAND2xp5_ASAP7_75t_SL g638 ( .A(n_564), .B(n_306), .Y(n_638) );
AO22x2_ASAP7_75t_L g639 ( .A1(n_607), .A2(n_577), .B1(n_579), .B2(n_582), .Y(n_639) );
AOI322xp5_ASAP7_75t_L g640 ( .A1(n_613), .A2(n_610), .A3(n_606), .B1(n_615), .B2(n_601), .C1(n_616), .C2(n_623), .Y(n_640) );
OAI221xp5_ASAP7_75t_SL g641 ( .A1(n_629), .A2(n_583), .B1(n_584), .B2(n_574), .C(n_548), .Y(n_641) );
INVxp67_ASAP7_75t_L g642 ( .A(n_604), .Y(n_642) );
NAND2xp5_ASAP7_75t_L g643 ( .A(n_605), .B(n_551), .Y(n_643) );
OAI21xp5_ASAP7_75t_L g644 ( .A1(n_612), .A2(n_580), .B(n_581), .Y(n_644) );
INVx1_ASAP7_75t_SL g645 ( .A(n_628), .Y(n_645) );
AOI221xp5_ASAP7_75t_L g646 ( .A1(n_609), .A2(n_593), .B1(n_592), .B2(n_591), .C(n_588), .Y(n_646) );
NAND3xp33_ASAP7_75t_L g647 ( .A(n_612), .B(n_564), .C(n_565), .Y(n_647) );
INVx1_ASAP7_75t_L g648 ( .A(n_603), .Y(n_648) );
AND2x2_ASAP7_75t_L g649 ( .A(n_614), .B(n_565), .Y(n_649) );
AOI21xp5_ASAP7_75t_L g650 ( .A1(n_625), .A2(n_567), .B(n_571), .Y(n_650) );
AOI221xp5_ASAP7_75t_L g651 ( .A1(n_626), .A2(n_598), .B1(n_589), .B2(n_221), .C(n_329), .Y(n_651) );
NAND3xp33_ASAP7_75t_L g652 ( .A(n_622), .B(n_221), .C(n_321), .Y(n_652) );
NAND2xp5_ASAP7_75t_L g653 ( .A(n_620), .B(n_45), .Y(n_653) );
CKINVDCx6p67_ASAP7_75t_R g654 ( .A(n_638), .Y(n_654) );
INVx1_ASAP7_75t_L g655 ( .A(n_636), .Y(n_655) );
OAI211xp5_ASAP7_75t_L g656 ( .A1(n_606), .A2(n_289), .B(n_321), .C(n_251), .Y(n_656) );
INVx1_ASAP7_75t_L g657 ( .A(n_624), .Y(n_657) );
NOR2xp33_ASAP7_75t_L g658 ( .A(n_608), .B(n_49), .Y(n_658) );
NOR2x1_ASAP7_75t_L g659 ( .A(n_637), .B(n_321), .Y(n_659) );
AO21x1_ASAP7_75t_L g660 ( .A1(n_616), .A2(n_51), .B(n_60), .Y(n_660) );
NOR3xp33_ASAP7_75t_L g661 ( .A(n_630), .B(n_61), .C(n_62), .Y(n_661) );
AND2x4_ASAP7_75t_L g662 ( .A(n_647), .B(n_602), .Y(n_662) );
NAND4xp25_ASAP7_75t_L g663 ( .A(n_640), .B(n_617), .C(n_601), .D(n_633), .Y(n_663) );
NOR3xp33_ASAP7_75t_L g664 ( .A(n_641), .B(n_635), .C(n_627), .Y(n_664) );
AND2x2_ASAP7_75t_L g665 ( .A(n_649), .B(n_621), .Y(n_665) );
NOR3x1_ASAP7_75t_L g666 ( .A(n_640), .B(n_611), .C(n_618), .Y(n_666) );
INVx3_ASAP7_75t_SL g667 ( .A(n_645), .Y(n_667) );
NOR2x1_ASAP7_75t_L g668 ( .A(n_656), .B(n_632), .Y(n_668) );
INVx4_ASAP7_75t_L g669 ( .A(n_654), .Y(n_669) );
INVx1_ASAP7_75t_L g670 ( .A(n_648), .Y(n_670) );
AND2x4_ASAP7_75t_L g671 ( .A(n_644), .B(n_621), .Y(n_671) );
NAND4xp75_ASAP7_75t_L g672 ( .A(n_660), .B(n_619), .C(n_634), .D(n_624), .Y(n_672) );
NAND2xp5_ASAP7_75t_L g673 ( .A(n_646), .B(n_631), .Y(n_673) );
INVxp33_ASAP7_75t_L g674 ( .A(n_658), .Y(n_674) );
INVx1_ASAP7_75t_L g675 ( .A(n_655), .Y(n_675) );
INVx2_ASAP7_75t_L g676 ( .A(n_670), .Y(n_676) );
OAI22xp5_ASAP7_75t_L g677 ( .A1(n_669), .A2(n_642), .B1(n_639), .B2(n_643), .Y(n_677) );
AOI221xp5_ASAP7_75t_L g678 ( .A1(n_663), .A2(n_669), .B1(n_673), .B2(n_662), .C(n_671), .Y(n_678) );
INVx1_ASAP7_75t_L g679 ( .A(n_675), .Y(n_679) );
INVx2_ASAP7_75t_L g680 ( .A(n_665), .Y(n_680) );
INVx2_ASAP7_75t_L g681 ( .A(n_671), .Y(n_681) );
OAI21xp33_ASAP7_75t_SL g682 ( .A1(n_672), .A2(n_657), .B(n_659), .Y(n_682) );
OAI21x1_ASAP7_75t_SL g683 ( .A1(n_668), .A2(n_650), .B(n_639), .Y(n_683) );
AOI211xp5_ASAP7_75t_L g684 ( .A1(n_678), .A2(n_667), .B(n_674), .C(n_666), .Y(n_684) );
AOI211xp5_ASAP7_75t_L g685 ( .A1(n_682), .A2(n_664), .B(n_662), .C(n_653), .Y(n_685) );
AND3x1_ASAP7_75t_L g686 ( .A(n_681), .B(n_668), .C(n_661), .Y(n_686) );
OR2x2_ASAP7_75t_L g687 ( .A(n_676), .B(n_679), .Y(n_687) );
AOI211xp5_ASAP7_75t_L g688 ( .A1(n_677), .A2(n_652), .B(n_651), .C(n_631), .Y(n_688) );
NAND4xp25_ASAP7_75t_SL g689 ( .A(n_684), .B(n_683), .C(n_680), .D(n_679), .Y(n_689) );
NOR3xp33_ASAP7_75t_L g690 ( .A(n_685), .B(n_63), .C(n_66), .Y(n_690) );
OAI221xp5_ASAP7_75t_L g691 ( .A1(n_686), .A2(n_251), .B1(n_289), .B2(n_71), .C(n_74), .Y(n_691) );
AOI221x1_ASAP7_75t_L g692 ( .A1(n_690), .A2(n_688), .B1(n_687), .B2(n_78), .C(n_69), .Y(n_692) );
AOI22xp5_ASAP7_75t_L g693 ( .A1(n_689), .A2(n_289), .B1(n_251), .B2(n_68), .Y(n_693) );
HB1xp67_ASAP7_75t_L g694 ( .A(n_693), .Y(n_694) );
AOI221xp5_ASAP7_75t_L g695 ( .A1(n_694), .A2(n_251), .B1(n_691), .B2(n_692), .C(n_689), .Y(n_695) );
endmodule