module fake_jpeg_11587_n_483 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_483);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_483;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx10_ASAP7_75t_L g17 ( 
.A(n_15),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_8),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_11),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_3),
.Y(n_23)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

CKINVDCx16_ASAP7_75t_R g25 ( 
.A(n_12),
.Y(n_25)
);

INVx6_ASAP7_75t_SL g26 ( 
.A(n_2),
.Y(n_26)
);

INVx11_ASAP7_75t_SL g27 ( 
.A(n_13),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_3),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_11),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_1),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_12),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_12),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_8),
.Y(n_39)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_5),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_7),
.Y(n_41)
);

CKINVDCx14_ASAP7_75t_R g42 ( 
.A(n_12),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_16),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_4),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_13),
.Y(n_45)
);

BUFx24_ASAP7_75t_L g46 ( 
.A(n_14),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_11),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_15),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_14),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_9),
.Y(n_50)
);

INVx13_ASAP7_75t_L g51 ( 
.A(n_7),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_16),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_8),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_11),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_7),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_0),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_3),
.Y(n_57)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_22),
.Y(n_58)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_58),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_48),
.B(n_16),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_59),
.B(n_76),
.Y(n_120)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_43),
.Y(n_60)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_60),
.Y(n_119)
);

INVx6_ASAP7_75t_SL g61 ( 
.A(n_26),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_61),
.B(n_64),
.Y(n_128)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_45),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g152 ( 
.A(n_62),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_39),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_63),
.Y(n_121)
);

CKINVDCx14_ASAP7_75t_R g64 ( 
.A(n_26),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_17),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_65),
.B(n_71),
.Y(n_131)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_21),
.Y(n_66)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_66),
.Y(n_140)
);

BUFx12f_ASAP7_75t_L g67 ( 
.A(n_26),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g166 ( 
.A(n_67),
.Y(n_166)
);

BUFx12f_ASAP7_75t_L g68 ( 
.A(n_21),
.Y(n_68)
);

INVx1_ASAP7_75t_SL g178 ( 
.A(n_68),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_39),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_69),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_39),
.Y(n_70)
);

INVx6_ASAP7_75t_L g132 ( 
.A(n_70),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_48),
.B(n_15),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_52),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_72),
.A2(n_42),
.B1(n_25),
.B2(n_57),
.Y(n_135)
);

INVx5_ASAP7_75t_L g73 ( 
.A(n_22),
.Y(n_73)
);

INVx2_ASAP7_75t_SL g156 ( 
.A(n_73),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_39),
.Y(n_74)
);

INVx6_ASAP7_75t_L g133 ( 
.A(n_74),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_43),
.B(n_0),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_75),
.B(n_77),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_18),
.B(n_57),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_17),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_53),
.Y(n_78)
);

INVx6_ASAP7_75t_L g137 ( 
.A(n_78),
.Y(n_137)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_22),
.Y(n_79)
);

INVx3_ASAP7_75t_L g144 ( 
.A(n_79),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_18),
.B(n_1),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_80),
.B(n_84),
.Y(n_155)
);

INVx5_ASAP7_75t_L g81 ( 
.A(n_24),
.Y(n_81)
);

INVx5_ASAP7_75t_L g118 ( 
.A(n_81),
.Y(n_118)
);

BUFx3_ASAP7_75t_L g82 ( 
.A(n_45),
.Y(n_82)
);

INVx5_ASAP7_75t_L g134 ( 
.A(n_82),
.Y(n_134)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_21),
.Y(n_83)
);

INVx3_ASAP7_75t_L g161 ( 
.A(n_83),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_19),
.B(n_1),
.Y(n_84)
);

INVx8_ASAP7_75t_L g85 ( 
.A(n_46),
.Y(n_85)
);

INVx5_ASAP7_75t_L g141 ( 
.A(n_85),
.Y(n_141)
);

INVx5_ASAP7_75t_L g86 ( 
.A(n_24),
.Y(n_86)
);

INVx5_ASAP7_75t_L g160 ( 
.A(n_86),
.Y(n_160)
);

AND2x2_ASAP7_75t_SL g87 ( 
.A(n_17),
.B(n_2),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_87),
.B(n_98),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_19),
.B(n_2),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_88),
.B(n_104),
.Y(n_147)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_20),
.Y(n_89)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_89),
.Y(n_126)
);

INVx5_ASAP7_75t_L g90 ( 
.A(n_24),
.Y(n_90)
);

INVx5_ASAP7_75t_L g177 ( 
.A(n_90),
.Y(n_177)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_45),
.Y(n_91)
);

INVx3_ASAP7_75t_L g162 ( 
.A(n_91),
.Y(n_162)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_32),
.Y(n_92)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_92),
.Y(n_146)
);

BUFx4f_ASAP7_75t_L g93 ( 
.A(n_46),
.Y(n_93)
);

INVx3_ASAP7_75t_L g169 ( 
.A(n_93),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_53),
.Y(n_94)
);

INVx6_ASAP7_75t_L g170 ( 
.A(n_94),
.Y(n_170)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_20),
.Y(n_95)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_95),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_53),
.Y(n_96)
);

INVx6_ASAP7_75t_L g172 ( 
.A(n_96),
.Y(n_172)
);

INVx4_ASAP7_75t_SL g97 ( 
.A(n_46),
.Y(n_97)
);

INVx4_ASAP7_75t_L g122 ( 
.A(n_97),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_23),
.B(n_3),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_53),
.Y(n_99)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_99),
.Y(n_127)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_32),
.Y(n_100)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_100),
.Y(n_159)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_28),
.Y(n_101)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_101),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_33),
.Y(n_102)
);

INVx4_ASAP7_75t_L g139 ( 
.A(n_102),
.Y(n_139)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_45),
.Y(n_103)
);

INVx4_ASAP7_75t_L g143 ( 
.A(n_103),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_23),
.B(n_4),
.Y(n_104)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_45),
.Y(n_105)
);

INVx4_ASAP7_75t_L g173 ( 
.A(n_105),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_17),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_106),
.B(n_107),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_17),
.Y(n_107)
);

BUFx3_ASAP7_75t_L g108 ( 
.A(n_49),
.Y(n_108)
);

INVx4_ASAP7_75t_L g175 ( 
.A(n_108),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_29),
.B(n_4),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_109),
.B(n_6),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_33),
.Y(n_110)
);

INVx4_ASAP7_75t_L g180 ( 
.A(n_110),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_29),
.B(n_6),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_111),
.B(n_115),
.Y(n_183)
);

INVx8_ASAP7_75t_L g112 ( 
.A(n_46),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_112),
.Y(n_151)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_28),
.Y(n_113)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_113),
.Y(n_154)
);

INVx5_ASAP7_75t_L g114 ( 
.A(n_49),
.Y(n_114)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_114),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_37),
.B(n_6),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_33),
.Y(n_116)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_116),
.Y(n_176)
);

CKINVDCx16_ASAP7_75t_R g117 ( 
.A(n_17),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_117),
.B(n_68),
.Y(n_186)
);

INVx11_ASAP7_75t_L g123 ( 
.A(n_97),
.Y(n_123)
);

INVx11_ASAP7_75t_L g198 ( 
.A(n_123),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_102),
.A2(n_116),
.B1(n_110),
.B2(n_52),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_124),
.A2(n_27),
.B1(n_78),
.B2(n_42),
.Y(n_210)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_85),
.A2(n_46),
.B1(n_49),
.B2(n_40),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_129),
.A2(n_135),
.B1(n_136),
.B2(n_142),
.Y(n_211)
);

AOI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_112),
.A2(n_40),
.B1(n_56),
.B2(n_52),
.Y(n_136)
);

NAND2xp33_ASAP7_75t_SL g138 ( 
.A(n_87),
.B(n_25),
.Y(n_138)
);

NAND2x1_ASAP7_75t_SL g213 ( 
.A(n_138),
.B(n_51),
.Y(n_213)
);

AOI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_67),
.A2(n_40),
.B1(n_56),
.B2(n_52),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_L g149 ( 
.A1(n_63),
.A2(n_35),
.B1(n_54),
.B2(n_47),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_149),
.A2(n_150),
.B1(n_167),
.B2(n_171),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_69),
.A2(n_55),
.B1(n_50),
.B2(n_44),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_158),
.B(n_164),
.Y(n_192)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_79),
.Y(n_163)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_163),
.Y(n_196)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_91),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_103),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_165),
.B(n_174),
.Y(n_203)
);

AOI22xp33_ASAP7_75t_L g167 ( 
.A1(n_70),
.A2(n_36),
.B1(n_54),
.B2(n_47),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_SL g171 ( 
.A1(n_67),
.A2(n_35),
.B1(n_41),
.B2(n_38),
.Y(n_171)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_105),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_L g179 ( 
.A1(n_74),
.A2(n_34),
.B1(n_41),
.B2(n_38),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g249 ( 
.A1(n_179),
.A2(n_184),
.B1(n_178),
.B2(n_151),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_73),
.B(n_50),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_SL g199 ( 
.A(n_182),
.B(n_187),
.Y(n_199)
);

AOI22xp33_ASAP7_75t_SL g184 ( 
.A1(n_66),
.A2(n_83),
.B1(n_81),
.B2(n_86),
.Y(n_184)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_90),
.Y(n_185)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_185),
.Y(n_190)
);

INVxp67_ASAP7_75t_L g245 ( 
.A(n_186),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_68),
.B(n_55),
.Y(n_187)
);

AOI22xp33_ASAP7_75t_SL g188 ( 
.A1(n_122),
.A2(n_30),
.B1(n_36),
.B2(n_34),
.Y(n_188)
);

INVxp67_ASAP7_75t_L g268 ( 
.A(n_188),
.Y(n_268)
);

INVx3_ASAP7_75t_L g189 ( 
.A(n_122),
.Y(n_189)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_189),
.Y(n_277)
);

CKINVDCx14_ASAP7_75t_R g191 ( 
.A(n_123),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_191),
.B(n_229),
.Y(n_253)
);

INVx5_ASAP7_75t_L g193 ( 
.A(n_175),
.Y(n_193)
);

HB1xp67_ASAP7_75t_L g262 ( 
.A(n_193),
.Y(n_262)
);

INVx2_ASAP7_75t_SL g194 ( 
.A(n_169),
.Y(n_194)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_194),
.Y(n_300)
);

AND2x2_ASAP7_75t_L g195 ( 
.A(n_157),
.B(n_62),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_195),
.B(n_172),
.C(n_245),
.Y(n_282)
);

BUFx6f_ASAP7_75t_L g197 ( 
.A(n_121),
.Y(n_197)
);

BUFx6f_ASAP7_75t_L g287 ( 
.A(n_197),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_147),
.B(n_31),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_200),
.B(n_216),
.Y(n_266)
);

INVx5_ASAP7_75t_L g201 ( 
.A(n_175),
.Y(n_201)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_201),
.Y(n_290)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_176),
.Y(n_202)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_202),
.Y(n_257)
);

BUFx6f_ASAP7_75t_L g204 ( 
.A(n_121),
.Y(n_204)
);

BUFx6f_ASAP7_75t_L g288 ( 
.A(n_204),
.Y(n_288)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_140),
.Y(n_205)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_205),
.Y(n_279)
);

AOI22xp33_ASAP7_75t_SL g206 ( 
.A1(n_126),
.A2(n_31),
.B1(n_30),
.B2(n_114),
.Y(n_206)
);

INVxp67_ASAP7_75t_L g269 ( 
.A(n_206),
.Y(n_269)
);

INVx4_ASAP7_75t_L g207 ( 
.A(n_134),
.Y(n_207)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_207),
.Y(n_280)
);

INVx3_ASAP7_75t_L g208 ( 
.A(n_118),
.Y(n_208)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_208),
.Y(n_291)
);

OAI22xp33_ASAP7_75t_SL g209 ( 
.A1(n_142),
.A2(n_99),
.B1(n_96),
.B2(n_94),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_209),
.A2(n_224),
.B1(n_248),
.B2(n_249),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_L g265 ( 
.A1(n_210),
.A2(n_231),
.B1(n_132),
.B2(n_170),
.Y(n_265)
);

INVx3_ASAP7_75t_L g212 ( 
.A(n_160),
.Y(n_212)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_212),
.Y(n_295)
);

AND2x2_ASAP7_75t_L g256 ( 
.A(n_213),
.B(n_221),
.Y(n_256)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_161),
.Y(n_214)
);

BUFx6f_ASAP7_75t_L g297 ( 
.A(n_214),
.Y(n_297)
);

INVx4_ASAP7_75t_L g215 ( 
.A(n_177),
.Y(n_215)
);

CKINVDCx16_ASAP7_75t_R g267 ( 
.A(n_215),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_120),
.B(n_44),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_130),
.B(n_37),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_217),
.B(n_225),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_153),
.B(n_131),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_218),
.B(n_220),
.Y(n_261)
);

AOI22xp33_ASAP7_75t_SL g219 ( 
.A1(n_145),
.A2(n_108),
.B1(n_82),
.B2(n_27),
.Y(n_219)
);

INVxp67_ASAP7_75t_L g272 ( 
.A(n_219),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_155),
.B(n_7),
.Y(n_220)
);

INVx4_ASAP7_75t_L g221 ( 
.A(n_143),
.Y(n_221)
);

INVx4_ASAP7_75t_L g222 ( 
.A(n_143),
.Y(n_222)
);

AND2x2_ASAP7_75t_L g264 ( 
.A(n_222),
.B(n_227),
.Y(n_264)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_154),
.Y(n_223)
);

INVxp67_ASAP7_75t_L g286 ( 
.A(n_223),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_136),
.A2(n_51),
.B1(n_93),
.B2(n_10),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_119),
.B(n_8),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_183),
.B(n_9),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_226),
.B(n_233),
.Y(n_274)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_146),
.Y(n_227)
);

BUFx3_ASAP7_75t_L g228 ( 
.A(n_166),
.Y(n_228)
);

INVxp67_ASAP7_75t_L g298 ( 
.A(n_228),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_181),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_162),
.Y(n_230)
);

AND2x2_ASAP7_75t_L g285 ( 
.A(n_230),
.B(n_232),
.Y(n_285)
);

AOI22xp33_ASAP7_75t_L g231 ( 
.A1(n_149),
.A2(n_51),
.B1(n_10),
.B2(n_13),
.Y(n_231)
);

BUFx3_ASAP7_75t_L g232 ( 
.A(n_166),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_128),
.Y(n_233)
);

INVx5_ASAP7_75t_L g234 ( 
.A(n_141),
.Y(n_234)
);

AOI22xp33_ASAP7_75t_SL g260 ( 
.A1(n_234),
.A2(n_241),
.B1(n_242),
.B2(n_243),
.Y(n_260)
);

BUFx2_ASAP7_75t_L g235 ( 
.A(n_168),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_235),
.Y(n_251)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_127),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_236),
.B(n_237),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_159),
.B(n_9),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_173),
.B(n_14),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_238),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_167),
.B(n_14),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_239),
.B(n_247),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_SL g241 ( 
.A(n_171),
.B(n_173),
.Y(n_241)
);

BUFx6f_ASAP7_75t_L g242 ( 
.A(n_148),
.Y(n_242)
);

AOI22xp33_ASAP7_75t_SL g243 ( 
.A1(n_178),
.A2(n_125),
.B1(n_129),
.B2(n_144),
.Y(n_243)
);

CKINVDCx16_ASAP7_75t_R g244 ( 
.A(n_184),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_244),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_179),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_246),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_127),
.B(n_180),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_139),
.A2(n_180),
.B1(n_133),
.B2(n_137),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_156),
.Y(n_250)
);

CKINVDCx12_ASAP7_75t_R g254 ( 
.A(n_250),
.Y(n_254)
);

FAx1_ASAP7_75t_L g252 ( 
.A(n_213),
.B(n_151),
.CI(n_156),
.CON(n_252),
.SN(n_252)
);

OR2x2_ASAP7_75t_L g305 ( 
.A(n_252),
.B(n_193),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_239),
.A2(n_139),
.B1(n_133),
.B2(n_137),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_258),
.A2(n_265),
.B1(n_293),
.B2(n_299),
.Y(n_301)
);

CKINVDCx12_ASAP7_75t_R g259 ( 
.A(n_198),
.Y(n_259)
);

CKINVDCx14_ASAP7_75t_R g329 ( 
.A(n_259),
.Y(n_329)
);

OAI21xp5_ASAP7_75t_L g263 ( 
.A1(n_217),
.A2(n_152),
.B(n_148),
.Y(n_263)
);

OAI21xp5_ASAP7_75t_L g322 ( 
.A1(n_263),
.A2(n_194),
.B(n_208),
.Y(n_322)
);

OAI21xp5_ASAP7_75t_SL g276 ( 
.A1(n_195),
.A2(n_152),
.B(n_132),
.Y(n_276)
);

AOI21xp5_ASAP7_75t_L g308 ( 
.A1(n_276),
.A2(n_278),
.B(n_296),
.Y(n_308)
);

OAI21xp5_ASAP7_75t_SL g278 ( 
.A1(n_195),
.A2(n_170),
.B(n_172),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g334 ( 
.A(n_282),
.B(n_278),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_225),
.B(n_200),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_284),
.B(n_289),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_216),
.B(n_192),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_245),
.B(n_223),
.C(n_203),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_292),
.B(n_282),
.C(n_256),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_L g293 ( 
.A1(n_210),
.A2(n_199),
.B1(n_211),
.B2(n_240),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_247),
.B(n_227),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_294),
.B(n_202),
.Y(n_309)
);

AOI21xp5_ASAP7_75t_L g296 ( 
.A1(n_198),
.A2(n_189),
.B(n_234),
.Y(n_296)
);

OAI22xp33_ASAP7_75t_SL g299 ( 
.A1(n_205),
.A2(n_214),
.B1(n_224),
.B2(n_236),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_SL g302 ( 
.A(n_289),
.B(n_196),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_SL g368 ( 
.A(n_302),
.B(n_304),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_SL g304 ( 
.A(n_266),
.B(n_230),
.Y(n_304)
);

OAI21xp5_ASAP7_75t_L g342 ( 
.A1(n_305),
.A2(n_313),
.B(n_330),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_255),
.B(n_235),
.Y(n_306)
);

INVxp67_ASAP7_75t_L g348 ( 
.A(n_306),
.Y(n_348)
);

OAI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_281),
.A2(n_283),
.B1(n_271),
.B2(n_273),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_L g339 ( 
.A1(n_307),
.A2(n_324),
.B1(n_338),
.B2(n_264),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_309),
.B(n_315),
.Y(n_341)
);

INVx2_ASAP7_75t_L g310 ( 
.A(n_300),
.Y(n_310)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_310),
.Y(n_343)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_283),
.A2(n_248),
.B1(n_242),
.B2(n_197),
.Y(n_311)
);

AND2x2_ASAP7_75t_L g349 ( 
.A(n_311),
.B(n_322),
.Y(n_349)
);

AOI22xp33_ASAP7_75t_SL g312 ( 
.A1(n_272),
.A2(n_207),
.B1(n_228),
.B2(n_232),
.Y(n_312)
);

INVxp67_ASAP7_75t_L g367 ( 
.A(n_312),
.Y(n_367)
);

AOI21xp5_ASAP7_75t_L g313 ( 
.A1(n_269),
.A2(n_270),
.B(n_268),
.Y(n_313)
);

XOR2xp5_ASAP7_75t_L g314 ( 
.A(n_284),
.B(n_190),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g363 ( 
.A(n_314),
.B(n_331),
.C(n_277),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_SL g315 ( 
.A(n_273),
.B(n_190),
.Y(n_315)
);

HB1xp67_ASAP7_75t_L g316 ( 
.A(n_291),
.Y(n_316)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_316),
.Y(n_344)
);

INVxp67_ASAP7_75t_L g317 ( 
.A(n_285),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_317),
.B(n_320),
.Y(n_346)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_300),
.Y(n_318)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_318),
.Y(n_345)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_294),
.Y(n_319)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_319),
.Y(n_347)
);

INVxp67_ASAP7_75t_L g320 ( 
.A(n_285),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_255),
.B(n_222),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_321),
.B(n_323),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_292),
.B(n_221),
.Y(n_323)
);

OAI22xp5_ASAP7_75t_SL g324 ( 
.A1(n_281),
.A2(n_204),
.B1(n_194),
.B2(n_212),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_L g325 ( 
.A1(n_258),
.A2(n_201),
.B1(n_215),
.B2(n_271),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_325),
.B(n_332),
.Y(n_355)
);

AND2x2_ASAP7_75t_L g326 ( 
.A(n_256),
.B(n_276),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_L g340 ( 
.A(n_326),
.B(n_327),
.Y(n_340)
);

BUFx6f_ASAP7_75t_L g328 ( 
.A(n_287),
.Y(n_328)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_328),
.Y(n_351)
);

O2A1O1Ixp33_ASAP7_75t_L g330 ( 
.A1(n_269),
.A2(n_268),
.B(n_252),
.C(n_256),
.Y(n_330)
);

XOR2xp5_ASAP7_75t_L g331 ( 
.A(n_266),
.B(n_275),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_L g332 ( 
.A1(n_270),
.A2(n_263),
.B1(n_272),
.B2(n_252),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_257),
.Y(n_333)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_333),
.Y(n_359)
);

XOR2xp5_ASAP7_75t_L g350 ( 
.A(n_334),
.B(n_327),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_SL g335 ( 
.A(n_253),
.B(n_274),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_335),
.B(n_337),
.Y(n_357)
);

BUFx24_ASAP7_75t_L g336 ( 
.A(n_254),
.Y(n_336)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_336),
.Y(n_365)
);

AOI22xp5_ASAP7_75t_L g337 ( 
.A1(n_260),
.A2(n_286),
.B1(n_295),
.B2(n_291),
.Y(n_337)
);

OAI22xp5_ASAP7_75t_L g338 ( 
.A1(n_286),
.A2(n_296),
.B1(n_261),
.B2(n_251),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_339),
.B(n_360),
.Y(n_374)
);

MAJIxp5_ASAP7_75t_L g391 ( 
.A(n_350),
.B(n_363),
.C(n_290),
.Y(n_391)
);

OAI21xp5_ASAP7_75t_L g352 ( 
.A1(n_305),
.A2(n_285),
.B(n_298),
.Y(n_352)
);

OAI21xp5_ASAP7_75t_L g381 ( 
.A1(n_352),
.A2(n_362),
.B(n_366),
.Y(n_381)
);

AOI22xp5_ASAP7_75t_SL g354 ( 
.A1(n_326),
.A2(n_298),
.B1(n_295),
.B2(n_280),
.Y(n_354)
);

INVxp67_ASAP7_75t_L g378 ( 
.A(n_354),
.Y(n_378)
);

AOI22xp5_ASAP7_75t_L g356 ( 
.A1(n_307),
.A2(n_280),
.B1(n_267),
.B2(n_264),
.Y(n_356)
);

OAI22xp5_ASAP7_75t_SL g373 ( 
.A1(n_356),
.A2(n_358),
.B1(n_361),
.B2(n_325),
.Y(n_373)
);

AOI22xp5_ASAP7_75t_L g358 ( 
.A1(n_324),
.A2(n_264),
.B1(n_279),
.B2(n_251),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_303),
.B(n_257),
.Y(n_360)
);

AOI22xp5_ASAP7_75t_L g361 ( 
.A1(n_319),
.A2(n_279),
.B1(n_287),
.B2(n_288),
.Y(n_361)
);

OAI21xp5_ASAP7_75t_L g362 ( 
.A1(n_305),
.A2(n_277),
.B(n_262),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_303),
.B(n_297),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_364),
.B(n_310),
.Y(n_383)
);

OAI21xp5_ASAP7_75t_L g366 ( 
.A1(n_330),
.A2(n_313),
.B(n_322),
.Y(n_366)
);

AND2x2_ASAP7_75t_L g369 ( 
.A(n_362),
.B(n_308),
.Y(n_369)
);

OAI21xp5_ASAP7_75t_SL g394 ( 
.A1(n_369),
.A2(n_384),
.B(n_386),
.Y(n_394)
);

AOI322xp5_ASAP7_75t_L g370 ( 
.A1(n_357),
.A2(n_338),
.A3(n_315),
.B1(n_304),
.B2(n_301),
.C1(n_332),
.C2(n_331),
.Y(n_370)
);

NOR4xp25_ASAP7_75t_L g397 ( 
.A(n_370),
.B(n_380),
.C(n_383),
.D(n_385),
.Y(n_397)
);

AOI22xp5_ASAP7_75t_L g371 ( 
.A1(n_349),
.A2(n_355),
.B1(n_357),
.B2(n_347),
.Y(n_371)
);

OAI22xp5_ASAP7_75t_SL g393 ( 
.A1(n_371),
.A2(n_372),
.B1(n_389),
.B2(n_339),
.Y(n_393)
);

AOI22xp5_ASAP7_75t_L g372 ( 
.A1(n_349),
.A2(n_301),
.B1(n_314),
.B2(n_309),
.Y(n_372)
);

AOI22xp5_ASAP7_75t_L g399 ( 
.A1(n_373),
.A2(n_349),
.B1(n_353),
.B2(n_348),
.Y(n_399)
);

INVx2_ASAP7_75t_SL g375 ( 
.A(n_359),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_375),
.B(n_379),
.Y(n_395)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_345),
.Y(n_376)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_376),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_L g377 ( 
.A(n_368),
.B(n_329),
.Y(n_377)
);

CKINVDCx14_ASAP7_75t_R g402 ( 
.A(n_377),
.Y(n_402)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_345),
.Y(n_379)
);

FAx1_ASAP7_75t_SL g380 ( 
.A(n_342),
.B(n_334),
.CI(n_326),
.CON(n_380),
.SN(n_380)
);

NOR2xp33_ASAP7_75t_L g382 ( 
.A(n_368),
.B(n_318),
.Y(n_382)
);

INVxp67_ASAP7_75t_L g405 ( 
.A(n_382),
.Y(n_405)
);

CKINVDCx20_ASAP7_75t_R g384 ( 
.A(n_364),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_360),
.B(n_333),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_359),
.Y(n_386)
);

OAI22x1_ASAP7_75t_L g387 ( 
.A1(n_342),
.A2(n_337),
.B1(n_311),
.B2(n_308),
.Y(n_387)
);

OAI21xp5_ASAP7_75t_SL g400 ( 
.A1(n_387),
.A2(n_367),
.B(n_354),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_341),
.B(n_317),
.Y(n_388)
);

XNOR2xp5_ASAP7_75t_L g406 ( 
.A(n_388),
.B(n_346),
.Y(n_406)
);

AOI22xp5_ASAP7_75t_L g389 ( 
.A1(n_349),
.A2(n_320),
.B1(n_328),
.B2(n_288),
.Y(n_389)
);

OAI21xp5_ASAP7_75t_L g390 ( 
.A1(n_366),
.A2(n_352),
.B(n_355),
.Y(n_390)
);

OAI21xp5_ASAP7_75t_L g411 ( 
.A1(n_390),
.A2(n_365),
.B(n_336),
.Y(n_411)
);

MAJIxp5_ASAP7_75t_L g403 ( 
.A(n_391),
.B(n_350),
.C(n_340),
.Y(n_403)
);

INVx2_ASAP7_75t_SL g392 ( 
.A(n_351),
.Y(n_392)
);

OAI21xp5_ASAP7_75t_SL g413 ( 
.A1(n_392),
.A2(n_290),
.B(n_336),
.Y(n_413)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_393),
.Y(n_424)
);

OAI22xp5_ASAP7_75t_SL g396 ( 
.A1(n_372),
.A2(n_347),
.B1(n_341),
.B2(n_356),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_396),
.B(n_398),
.Y(n_416)
);

OAI22xp5_ASAP7_75t_SL g398 ( 
.A1(n_374),
.A2(n_371),
.B1(n_384),
.B2(n_378),
.Y(n_398)
);

OAI22xp5_ASAP7_75t_L g425 ( 
.A1(n_399),
.A2(n_404),
.B1(n_409),
.B2(n_410),
.Y(n_425)
);

OAI31xp33_ASAP7_75t_L g430 ( 
.A1(n_400),
.A2(n_380),
.A3(n_370),
.B(n_389),
.Y(n_430)
);

OAI22xp5_ASAP7_75t_SL g401 ( 
.A1(n_374),
.A2(n_363),
.B1(n_358),
.B2(n_354),
.Y(n_401)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_401),
.Y(n_428)
);

MAJIxp5_ASAP7_75t_L g418 ( 
.A(n_403),
.B(n_407),
.C(n_412),
.Y(n_418)
);

AOI22xp5_ASAP7_75t_L g404 ( 
.A1(n_373),
.A2(n_353),
.B1(n_350),
.B2(n_363),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_SL g414 ( 
.A(n_406),
.B(n_413),
.Y(n_414)
);

MAJIxp5_ASAP7_75t_L g407 ( 
.A(n_391),
.B(n_340),
.C(n_346),
.Y(n_407)
);

AOI22xp5_ASAP7_75t_L g409 ( 
.A1(n_390),
.A2(n_344),
.B1(n_343),
.B2(n_351),
.Y(n_409)
);

AOI22xp5_ASAP7_75t_L g410 ( 
.A1(n_369),
.A2(n_344),
.B1(n_343),
.B2(n_361),
.Y(n_410)
);

AOI21xp33_ASAP7_75t_L g427 ( 
.A1(n_411),
.A2(n_388),
.B(n_385),
.Y(n_427)
);

XNOR2xp5_ASAP7_75t_L g412 ( 
.A(n_391),
.B(n_365),
.Y(n_412)
);

CKINVDCx20_ASAP7_75t_R g415 ( 
.A(n_395),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_415),
.B(n_417),
.Y(n_443)
);

CKINVDCx20_ASAP7_75t_R g417 ( 
.A(n_395),
.Y(n_417)
);

CKINVDCx14_ASAP7_75t_R g419 ( 
.A(n_402),
.Y(n_419)
);

OAI22xp5_ASAP7_75t_L g441 ( 
.A1(n_419),
.A2(n_410),
.B1(n_408),
.B2(n_376),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_SL g420 ( 
.A(n_405),
.B(n_377),
.Y(n_420)
);

CKINVDCx20_ASAP7_75t_R g431 ( 
.A(n_420),
.Y(n_431)
);

XNOR2xp5_ASAP7_75t_L g421 ( 
.A(n_403),
.B(n_381),
.Y(n_421)
);

MAJIxp5_ASAP7_75t_L g440 ( 
.A(n_421),
.B(n_422),
.C(n_423),
.Y(n_440)
);

XNOR2xp5_ASAP7_75t_L g422 ( 
.A(n_403),
.B(n_381),
.Y(n_422)
);

MAJIxp5_ASAP7_75t_L g423 ( 
.A(n_407),
.B(n_369),
.C(n_387),
.Y(n_423)
);

MAJIxp5_ASAP7_75t_L g426 ( 
.A(n_412),
.B(n_369),
.C(n_387),
.Y(n_426)
);

OR2x2_ASAP7_75t_L g444 ( 
.A(n_426),
.B(n_429),
.Y(n_444)
);

AOI21xp5_ASAP7_75t_L g442 ( 
.A1(n_427),
.A2(n_430),
.B(n_400),
.Y(n_442)
);

CKINVDCx20_ASAP7_75t_R g429 ( 
.A(n_402),
.Y(n_429)
);

OAI21xp33_ASAP7_75t_L g432 ( 
.A1(n_430),
.A2(n_397),
.B(n_380),
.Y(n_432)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_432),
.Y(n_452)
);

AOI22xp5_ASAP7_75t_L g433 ( 
.A1(n_424),
.A2(n_393),
.B1(n_398),
.B2(n_401),
.Y(n_433)
);

OAI22xp5_ASAP7_75t_L g451 ( 
.A1(n_433),
.A2(n_436),
.B1(n_442),
.B2(n_414),
.Y(n_451)
);

OAI322xp33_ASAP7_75t_L g434 ( 
.A1(n_421),
.A2(n_382),
.A3(n_397),
.B1(n_380),
.B2(n_406),
.C1(n_411),
.C2(n_383),
.Y(n_434)
);

NOR2xp33_ASAP7_75t_L g449 ( 
.A(n_434),
.B(n_438),
.Y(n_449)
);

OAI22xp5_ASAP7_75t_SL g435 ( 
.A1(n_424),
.A2(n_399),
.B1(n_404),
.B2(n_409),
.Y(n_435)
);

AOI22xp5_ASAP7_75t_L g448 ( 
.A1(n_435),
.A2(n_441),
.B1(n_396),
.B2(n_425),
.Y(n_448)
);

NOR3xp33_ASAP7_75t_SL g436 ( 
.A(n_428),
.B(n_408),
.C(n_379),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_416),
.Y(n_437)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_437),
.Y(n_445)
);

BUFx24_ASAP7_75t_SL g438 ( 
.A(n_429),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_416),
.Y(n_439)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_439),
.Y(n_447)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_437),
.Y(n_446)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_446),
.Y(n_461)
);

OAI22xp5_ASAP7_75t_SL g463 ( 
.A1(n_448),
.A2(n_450),
.B1(n_439),
.B2(n_443),
.Y(n_463)
);

OAI22xp33_ASAP7_75t_L g450 ( 
.A1(n_443),
.A2(n_417),
.B1(n_415),
.B2(n_428),
.Y(n_450)
);

XNOR2xp5_ASAP7_75t_L g459 ( 
.A(n_451),
.B(n_425),
.Y(n_459)
);

MAJIxp5_ASAP7_75t_L g453 ( 
.A(n_440),
.B(n_418),
.C(n_422),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_SL g460 ( 
.A(n_453),
.B(n_454),
.Y(n_460)
);

MAJIxp5_ASAP7_75t_L g454 ( 
.A(n_440),
.B(n_418),
.C(n_444),
.Y(n_454)
);

XOR2xp5_ASAP7_75t_L g455 ( 
.A(n_448),
.B(n_426),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_455),
.B(n_457),
.Y(n_465)
);

NOR2xp33_ASAP7_75t_L g456 ( 
.A(n_454),
.B(n_431),
.Y(n_456)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_456),
.Y(n_464)
);

MAJIxp5_ASAP7_75t_L g457 ( 
.A(n_453),
.B(n_444),
.C(n_433),
.Y(n_457)
);

MAJIxp5_ASAP7_75t_L g458 ( 
.A(n_450),
.B(n_423),
.C(n_435),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_458),
.B(n_459),
.Y(n_466)
);

NOR2xp33_ASAP7_75t_SL g462 ( 
.A(n_449),
.B(n_442),
.Y(n_462)
);

CKINVDCx16_ASAP7_75t_R g467 ( 
.A(n_462),
.Y(n_467)
);

OAI22xp5_ASAP7_75t_L g468 ( 
.A1(n_463),
.A2(n_447),
.B1(n_445),
.B2(n_446),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_468),
.B(n_469),
.Y(n_471)
);

OAI22xp5_ASAP7_75t_L g469 ( 
.A1(n_457),
.A2(n_447),
.B1(n_445),
.B2(n_452),
.Y(n_469)
);

OAI21xp5_ASAP7_75t_SL g470 ( 
.A1(n_460),
.A2(n_458),
.B(n_461),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_470),
.B(n_459),
.Y(n_474)
);

AOI31xp33_ASAP7_75t_L g472 ( 
.A1(n_464),
.A2(n_414),
.A3(n_436),
.B(n_463),
.Y(n_472)
);

MAJIxp5_ASAP7_75t_L g475 ( 
.A(n_472),
.B(n_470),
.C(n_467),
.Y(n_475)
);

INVxp67_ASAP7_75t_L g473 ( 
.A(n_466),
.Y(n_473)
);

OAI21xp5_ASAP7_75t_L g476 ( 
.A1(n_473),
.A2(n_465),
.B(n_466),
.Y(n_476)
);

O2A1O1Ixp33_ASAP7_75t_SL g477 ( 
.A1(n_474),
.A2(n_465),
.B(n_455),
.C(n_394),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_475),
.B(n_476),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_SL g478 ( 
.A(n_477),
.B(n_471),
.Y(n_478)
);

AOI321xp33_ASAP7_75t_L g480 ( 
.A1(n_478),
.A2(n_386),
.A3(n_394),
.B1(n_413),
.B2(n_375),
.C(n_336),
.Y(n_480)
);

AOI22xp33_ASAP7_75t_L g481 ( 
.A1(n_480),
.A2(n_375),
.B1(n_392),
.B2(n_479),
.Y(n_481)
);

AOI221xp5_ASAP7_75t_L g482 ( 
.A1(n_481),
.A2(n_375),
.B1(n_392),
.B2(n_328),
.C(n_297),
.Y(n_482)
);

XOR2xp5_ASAP7_75t_L g483 ( 
.A(n_482),
.B(n_392),
.Y(n_483)
);


endmodule