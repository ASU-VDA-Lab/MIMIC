module fake_jpeg_27094_n_69 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_69);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_69;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_23;
wire n_10;
wire n_27;
wire n_55;
wire n_64;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_59;
wire n_35;
wire n_48;
wire n_68;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_65;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_44;
wire n_26;
wire n_38;
wire n_9;
wire n_36;
wire n_11;
wire n_62;
wire n_17;
wire n_25;
wire n_31;
wire n_56;
wire n_67;
wire n_29;
wire n_37;
wire n_50;
wire n_43;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_66;

CKINVDCx20_ASAP7_75t_R g8 ( 
.A(n_6),
.Y(n_8)
);

INVx1_ASAP7_75t_L g9 ( 
.A(n_2),
.Y(n_9)
);

BUFx12_ASAP7_75t_L g10 ( 
.A(n_4),
.Y(n_10)
);

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_2),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_7),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_7),
.Y(n_13)
);

INVx2_ASAP7_75t_L g14 ( 
.A(n_6),
.Y(n_14)
);

BUFx12f_ASAP7_75t_L g15 ( 
.A(n_4),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_14),
.B(n_0),
.Y(n_18)
);

AND2x2_ASAP7_75t_L g26 ( 
.A(n_18),
.B(n_17),
.Y(n_26)
);

AOI22xp33_ASAP7_75t_L g19 ( 
.A1(n_14),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_19),
.B(n_21),
.Y(n_25)
);

INVx11_ASAP7_75t_L g20 ( 
.A(n_15),
.Y(n_20)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_20),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_22),
.B(n_23),
.Y(n_29)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_17),
.Y(n_23)
);

AOI21xp5_ASAP7_75t_L g24 ( 
.A1(n_18),
.A2(n_19),
.B(n_21),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g37 ( 
.A(n_24),
.B(n_25),
.C(n_26),
.Y(n_37)
);

OR2x2_ASAP7_75t_L g42 ( 
.A(n_26),
.B(n_30),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_18),
.B(n_12),
.Y(n_27)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_27),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_SL g30 ( 
.A(n_22),
.B(n_11),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_29),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_31),
.B(n_33),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_29),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_32),
.B(n_36),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_30),
.B(n_12),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_L g34 ( 
.A1(n_26),
.A2(n_23),
.B1(n_22),
.B2(n_20),
.Y(n_34)
);

AOI22xp5_ASAP7_75t_L g47 ( 
.A1(n_34),
.A2(n_40),
.B1(n_21),
.B2(n_10),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g35 ( 
.A1(n_24),
.A2(n_23),
.B1(n_11),
.B2(n_16),
.Y(n_35)
);

AOI22xp5_ASAP7_75t_L g46 ( 
.A1(n_35),
.A2(n_9),
.B1(n_13),
.B2(n_20),
.Y(n_46)
);

INVxp67_ASAP7_75t_L g36 ( 
.A(n_28),
.Y(n_36)
);

AND2x2_ASAP7_75t_L g50 ( 
.A(n_37),
.B(n_1),
.Y(n_50)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_28),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_39),
.B(n_1),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g40 ( 
.A1(n_25),
.A2(n_20),
.B1(n_16),
.B2(n_9),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_30),
.B(n_8),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_41),
.B(n_3),
.Y(n_49)
);

INVxp67_ASAP7_75t_L g45 ( 
.A(n_40),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_45),
.B(n_48),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_46),
.B(n_47),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_49),
.B(n_50),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_43),
.Y(n_54)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_54),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_45),
.A2(n_37),
.B1(n_34),
.B2(n_42),
.Y(n_55)
);

AOI21xp5_ASAP7_75t_L g57 ( 
.A1(n_55),
.A2(n_50),
.B(n_42),
.Y(n_57)
);

HB1xp67_ASAP7_75t_L g56 ( 
.A(n_54),
.Y(n_56)
);

INVxp67_ASAP7_75t_L g61 ( 
.A(n_56),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_57),
.A2(n_52),
.B1(n_51),
.B2(n_44),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_55),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_59),
.B(n_51),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_60),
.B(n_62),
.Y(n_64)
);

OAI21xp5_ASAP7_75t_L g63 ( 
.A1(n_61),
.A2(n_58),
.B(n_53),
.Y(n_63)
);

O2A1O1Ixp33_ASAP7_75t_SL g65 ( 
.A1(n_63),
.A2(n_61),
.B(n_31),
.C(n_38),
.Y(n_65)
);

OAI21xp5_ASAP7_75t_L g67 ( 
.A1(n_65),
.A2(n_66),
.B(n_5),
.Y(n_67)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_64),
.B(n_3),
.Y(n_66)
);

OAI21xp5_ASAP7_75t_SL g68 ( 
.A1(n_67),
.A2(n_36),
.B(n_47),
.Y(n_68)
);

XNOR2xp5_ASAP7_75t_L g69 ( 
.A(n_68),
.B(n_10),
.Y(n_69)
);


endmodule