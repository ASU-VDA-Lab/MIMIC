module fake_jpeg_15816_n_188 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_188);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_188;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

INVx11_ASAP7_75t_SL g17 ( 
.A(n_0),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_13),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_7),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_10),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

INVxp67_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

CKINVDCx16_ASAP7_75t_R g25 ( 
.A(n_0),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_5),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_2),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

OR2x4_ASAP7_75t_L g32 ( 
.A(n_17),
.B(n_1),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_SL g49 ( 
.A(n_32),
.B(n_25),
.Y(n_49)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_23),
.Y(n_33)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_33),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_34),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_22),
.B(n_3),
.Y(n_35)
);

AND2x2_ASAP7_75t_L g48 ( 
.A(n_35),
.B(n_19),
.Y(n_48)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_15),
.Y(n_36)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_36),
.Y(n_44)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_23),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

BUFx12_ASAP7_75t_L g38 ( 
.A(n_23),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_15),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_39),
.B(n_42),
.Y(n_52)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_16),
.Y(n_40)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_16),
.Y(n_41)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_41),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_16),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_35),
.B(n_31),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_43),
.B(n_45),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_32),
.B(n_31),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_40),
.A2(n_25),
.B1(n_29),
.B2(n_22),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_46),
.A2(n_54),
.B1(n_58),
.B2(n_30),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_48),
.B(n_28),
.Y(n_67)
);

CKINVDCx14_ASAP7_75t_R g64 ( 
.A(n_49),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_39),
.A2(n_24),
.B1(n_19),
.B2(n_27),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_50),
.A2(n_60),
.B1(n_37),
.B2(n_20),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_36),
.A2(n_29),
.B1(n_26),
.B2(n_21),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_38),
.B(n_21),
.Y(n_55)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_55),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_L g58 ( 
.A1(n_33),
.A2(n_27),
.B1(n_26),
.B2(n_18),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g60 ( 
.A(n_34),
.B(n_3),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_38),
.B(n_18),
.Y(n_61)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_61),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_62),
.B(n_67),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g63 ( 
.A(n_50),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_63),
.B(n_73),
.Y(n_84)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_44),
.Y(n_68)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_68),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_57),
.A2(n_20),
.B1(n_28),
.B2(n_30),
.Y(n_69)
);

OAI22x1_ASAP7_75t_L g82 ( 
.A1(n_69),
.A2(n_71),
.B1(n_80),
.B2(n_20),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_43),
.B(n_42),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_70),
.B(n_52),
.Y(n_91)
);

OAI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_47),
.A2(n_42),
.B1(n_41),
.B2(n_34),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_72),
.A2(n_47),
.B1(n_52),
.B2(n_44),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_61),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_59),
.Y(n_74)
);

INVx1_ASAP7_75t_SL g89 ( 
.A(n_74),
.Y(n_89)
);

A2O1A1Ixp33_ASAP7_75t_L g75 ( 
.A1(n_45),
.A2(n_4),
.B(n_5),
.C(n_6),
.Y(n_75)
);

CKINVDCx14_ASAP7_75t_R g97 ( 
.A(n_75),
.Y(n_97)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_57),
.Y(n_77)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_77),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g78 ( 
.A(n_55),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_78),
.B(n_53),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_60),
.A2(n_48),
.B1(n_49),
.B2(n_51),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_79),
.A2(n_51),
.B1(n_47),
.B2(n_28),
.Y(n_93)
);

AOI21xp5_ASAP7_75t_L g80 ( 
.A1(n_60),
.A2(n_4),
.B(n_6),
.Y(n_80)
);

BUFx2_ASAP7_75t_SL g81 ( 
.A(n_77),
.Y(n_81)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_81),
.Y(n_101)
);

OA22x2_ASAP7_75t_L g105 ( 
.A1(n_82),
.A2(n_87),
.B1(n_59),
.B2(n_30),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_85),
.B(n_88),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_73),
.B(n_53),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_91),
.B(n_92),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_70),
.B(n_48),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_93),
.B(n_98),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_63),
.A2(n_41),
.B1(n_59),
.B2(n_53),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_94),
.A2(n_96),
.B1(n_80),
.B2(n_65),
.Y(n_104)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_68),
.Y(n_95)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_95),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_67),
.A2(n_78),
.B1(n_62),
.B2(n_64),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_74),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_76),
.B(n_56),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_99),
.B(n_100),
.Y(n_103)
);

OR2x2_ASAP7_75t_L g100 ( 
.A(n_79),
.B(n_65),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_104),
.A2(n_105),
.B1(n_114),
.B2(n_115),
.Y(n_133)
);

A2O1A1O1Ixp25_ASAP7_75t_L g106 ( 
.A1(n_100),
.A2(n_76),
.B(n_75),
.C(n_66),
.D(n_38),
.Y(n_106)
);

XOR2xp5_ASAP7_75t_SL g127 ( 
.A(n_106),
.B(n_4),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_83),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_108),
.B(n_95),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_91),
.B(n_66),
.C(n_56),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_SL g128 ( 
.A(n_109),
.B(n_9),
.Y(n_128)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_90),
.Y(n_110)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_110),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_82),
.A2(n_97),
.B1(n_98),
.B2(n_89),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_111),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_92),
.B(n_74),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_113),
.B(n_116),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_84),
.A2(n_100),
.B1(n_86),
.B2(n_93),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_84),
.A2(n_56),
.B1(n_6),
.B2(n_7),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_99),
.B(n_96),
.Y(n_116)
);

AOI21xp5_ASAP7_75t_L g118 ( 
.A1(n_86),
.A2(n_56),
.B(n_8),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_SL g122 ( 
.A1(n_118),
.A2(n_83),
.B(n_87),
.Y(n_122)
);

AOI21xp5_ASAP7_75t_L g120 ( 
.A1(n_103),
.A2(n_86),
.B(n_90),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_SL g147 ( 
.A1(n_120),
.A2(n_122),
.B(n_124),
.Y(n_147)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_121),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_107),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_123),
.B(n_134),
.Y(n_142)
);

OAI32xp33_ASAP7_75t_L g124 ( 
.A1(n_116),
.A2(n_94),
.A3(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_101),
.B(n_89),
.Y(n_126)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_126),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_L g135 ( 
.A(n_127),
.B(n_128),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_102),
.B(n_9),
.Y(n_130)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_130),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_102),
.B(n_10),
.Y(n_131)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_131),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_103),
.B(n_11),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_132),
.B(n_115),
.Y(n_136)
);

CKINVDCx16_ASAP7_75t_R g134 ( 
.A(n_107),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_136),
.B(n_141),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_129),
.B(n_113),
.Y(n_137)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_137),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_L g138 ( 
.A(n_120),
.B(n_109),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_138),
.B(n_128),
.C(n_114),
.Y(n_149)
);

CKINVDCx16_ASAP7_75t_R g139 ( 
.A(n_125),
.Y(n_139)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_139),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_129),
.B(n_101),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_130),
.B(n_108),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_SL g152 ( 
.A(n_143),
.B(n_132),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_123),
.B(n_110),
.Y(n_148)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_148),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_149),
.B(n_159),
.C(n_147),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_137),
.A2(n_119),
.B1(n_133),
.B2(n_117),
.Y(n_150)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_150),
.Y(n_160)
);

XOR2xp5_ASAP7_75t_L g151 ( 
.A(n_138),
.B(n_133),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_151),
.B(n_152),
.Y(n_167)
);

OA21x2_ASAP7_75t_SL g153 ( 
.A1(n_135),
.A2(n_127),
.B(n_106),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_L g165 ( 
.A1(n_153),
.A2(n_131),
.B(n_142),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_147),
.A2(n_119),
.B1(n_105),
.B2(n_124),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_157),
.A2(n_146),
.B1(n_140),
.B2(n_143),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_SL g159 ( 
.A(n_135),
.B(n_118),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_161),
.B(n_162),
.C(n_104),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_151),
.B(n_146),
.C(n_140),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_163),
.A2(n_164),
.B1(n_160),
.B2(n_166),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_156),
.A2(n_136),
.B1(n_145),
.B2(n_144),
.Y(n_164)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_165),
.Y(n_173)
);

INVxp67_ASAP7_75t_L g166 ( 
.A(n_155),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_166),
.A2(n_156),
.B1(n_154),
.B2(n_158),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_168),
.A2(n_170),
.B1(n_171),
.B2(n_173),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_169),
.B(n_11),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_162),
.A2(n_150),
.B1(n_149),
.B2(n_157),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_161),
.A2(n_105),
.B1(n_112),
.B2(n_152),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_167),
.A2(n_159),
.B1(n_105),
.B2(n_122),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_172),
.B(n_12),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_174),
.B(n_167),
.C(n_125),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_175),
.B(n_177),
.Y(n_180)
);

INVxp67_ASAP7_75t_L g181 ( 
.A(n_176),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_SL g182 ( 
.A(n_178),
.B(n_179),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_174),
.B(n_13),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g183 ( 
.A(n_180),
.B(n_170),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_L g185 ( 
.A1(n_183),
.A2(n_184),
.B(n_181),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_SL g184 ( 
.A1(n_182),
.A2(n_177),
.B(n_169),
.Y(n_184)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_185),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_L g187 ( 
.A1(n_186),
.A2(n_172),
.B(n_14),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_187),
.B(n_14),
.Y(n_188)
);


endmodule