module fake_jpeg_11879_n_641 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_641);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_641;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_19;
wire n_182;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_620;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_638;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_637;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_639;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_92;
wire n_332;
wire n_640;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_615;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_384;
wire n_296;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_599;
wire n_239;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_587;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx12_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

BUFx8_ASAP7_75t_L g20 ( 
.A(n_16),
.Y(n_20)
);

INVx4_ASAP7_75t_L g21 ( 
.A(n_16),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_10),
.B(n_5),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_16),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_6),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_3),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_4),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_11),
.Y(n_36)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_13),
.Y(n_37)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_15),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_14),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_3),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_4),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_3),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_0),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_17),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_12),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_10),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_17),
.Y(n_47)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_6),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_4),
.B(n_3),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_11),
.Y(n_50)
);

INVx11_ASAP7_75t_L g51 ( 
.A(n_18),
.Y(n_51)
);

BUFx24_ASAP7_75t_L g52 ( 
.A(n_11),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_17),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_13),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_7),
.Y(n_55)
);

CKINVDCx16_ASAP7_75t_R g56 ( 
.A(n_9),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_14),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_11),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_18),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_33),
.Y(n_60)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_60),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_26),
.B(n_9),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_61),
.B(n_113),
.Y(n_149)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_21),
.Y(n_62)
);

INVx3_ASAP7_75t_L g162 ( 
.A(n_62),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_22),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_63),
.Y(n_135)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_33),
.Y(n_64)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_64),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_22),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_65),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_22),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_66),
.Y(n_157)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_25),
.Y(n_67)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_67),
.Y(n_130)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_21),
.Y(n_68)
);

INVx3_ASAP7_75t_L g170 ( 
.A(n_68),
.Y(n_170)
);

BUFx8_ASAP7_75t_L g69 ( 
.A(n_52),
.Y(n_69)
);

BUFx12f_ASAP7_75t_L g184 ( 
.A(n_69),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_19),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_70),
.B(n_72),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_26),
.B(n_9),
.C(n_17),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_71),
.B(n_104),
.C(n_43),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_19),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_22),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_73),
.Y(n_166)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_21),
.Y(n_74)
);

INVx3_ASAP7_75t_L g192 ( 
.A(n_74),
.Y(n_192)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_28),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g177 ( 
.A(n_75),
.Y(n_177)
);

BUFx12f_ASAP7_75t_L g76 ( 
.A(n_20),
.Y(n_76)
);

BUFx3_ASAP7_75t_L g174 ( 
.A(n_76),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_28),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g181 ( 
.A(n_77),
.Y(n_181)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_28),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g182 ( 
.A(n_78),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_19),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_79),
.B(n_92),
.Y(n_138)
);

BUFx12f_ASAP7_75t_L g80 ( 
.A(n_20),
.Y(n_80)
);

BUFx3_ASAP7_75t_L g206 ( 
.A(n_80),
.Y(n_206)
);

BUFx2_ASAP7_75t_L g81 ( 
.A(n_27),
.Y(n_81)
);

INVx1_ASAP7_75t_SL g165 ( 
.A(n_81),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_28),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g186 ( 
.A(n_82),
.Y(n_186)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_20),
.Y(n_83)
);

INVx3_ASAP7_75t_L g198 ( 
.A(n_83),
.Y(n_198)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_34),
.Y(n_84)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_84),
.Y(n_158)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_34),
.Y(n_85)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_85),
.Y(n_188)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_25),
.Y(n_86)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_86),
.Y(n_132)
);

BUFx5_ASAP7_75t_L g87 ( 
.A(n_27),
.Y(n_87)
);

BUFx5_ASAP7_75t_L g168 ( 
.A(n_87),
.Y(n_168)
);

BUFx3_ASAP7_75t_L g88 ( 
.A(n_27),
.Y(n_88)
);

BUFx12f_ASAP7_75t_L g190 ( 
.A(n_88),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_49),
.B(n_9),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_89),
.B(n_109),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_53),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g195 ( 
.A(n_90),
.Y(n_195)
);

BUFx5_ASAP7_75t_L g91 ( 
.A(n_37),
.Y(n_91)
);

BUFx12f_ASAP7_75t_L g196 ( 
.A(n_91),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_19),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_49),
.B(n_8),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_93),
.B(n_94),
.Y(n_146)
);

BUFx12f_ASAP7_75t_SL g94 ( 
.A(n_52),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_53),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g210 ( 
.A(n_95),
.Y(n_210)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_53),
.Y(n_96)
);

INVx6_ASAP7_75t_L g140 ( 
.A(n_96),
.Y(n_140)
);

BUFx2_ASAP7_75t_L g97 ( 
.A(n_37),
.Y(n_97)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_97),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_53),
.Y(n_98)
);

INVx6_ASAP7_75t_L g180 ( 
.A(n_98),
.Y(n_180)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_29),
.Y(n_99)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_99),
.Y(n_155)
);

BUFx12f_ASAP7_75t_L g100 ( 
.A(n_20),
.Y(n_100)
);

INVx5_ASAP7_75t_L g167 ( 
.A(n_100),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_30),
.Y(n_101)
);

INVx8_ASAP7_75t_L g176 ( 
.A(n_101),
.Y(n_176)
);

INVx11_ASAP7_75t_L g102 ( 
.A(n_52),
.Y(n_102)
);

CKINVDCx14_ASAP7_75t_R g160 ( 
.A(n_102),
.Y(n_160)
);

BUFx3_ASAP7_75t_L g103 ( 
.A(n_37),
.Y(n_103)
);

INVx5_ASAP7_75t_L g200 ( 
.A(n_103),
.Y(n_200)
);

AOI21xp5_ASAP7_75t_L g104 ( 
.A1(n_52),
.A2(n_18),
.B(n_8),
.Y(n_104)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_29),
.Y(n_105)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_105),
.Y(n_163)
);

INVx5_ASAP7_75t_L g106 ( 
.A(n_48),
.Y(n_106)
);

INVx2_ASAP7_75t_SL g152 ( 
.A(n_106),
.Y(n_152)
);

INVx11_ASAP7_75t_L g107 ( 
.A(n_52),
.Y(n_107)
);

INVx4_ASAP7_75t_L g143 ( 
.A(n_107),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_30),
.Y(n_108)
);

INVx5_ASAP7_75t_L g217 ( 
.A(n_108),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_32),
.B(n_8),
.Y(n_109)
);

BUFx3_ASAP7_75t_L g110 ( 
.A(n_42),
.Y(n_110)
);

INVx4_ASAP7_75t_L g134 ( 
.A(n_110),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_30),
.Y(n_111)
);

INVx4_ASAP7_75t_L g204 ( 
.A(n_111),
.Y(n_204)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_57),
.Y(n_112)
);

INVx4_ASAP7_75t_L g205 ( 
.A(n_112),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_32),
.B(n_10),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_35),
.B(n_7),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_114),
.B(n_41),
.Y(n_179)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_20),
.Y(n_115)
);

INVx3_ASAP7_75t_L g202 ( 
.A(n_115),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_35),
.B(n_18),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_116),
.B(n_56),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_57),
.Y(n_117)
);

INVx4_ASAP7_75t_L g209 ( 
.A(n_117),
.Y(n_209)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_57),
.Y(n_118)
);

INVx3_ASAP7_75t_L g213 ( 
.A(n_118),
.Y(n_213)
);

BUFx12f_ASAP7_75t_L g119 ( 
.A(n_51),
.Y(n_119)
);

INVx4_ASAP7_75t_L g211 ( 
.A(n_119),
.Y(n_211)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_23),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_120),
.B(n_123),
.Y(n_153)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_42),
.Y(n_121)
);

INVx3_ASAP7_75t_L g214 ( 
.A(n_121),
.Y(n_214)
);

BUFx16f_ASAP7_75t_L g122 ( 
.A(n_42),
.Y(n_122)
);

INVx13_ASAP7_75t_L g187 ( 
.A(n_122),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_19),
.Y(n_123)
);

INVx5_ASAP7_75t_L g124 ( 
.A(n_48),
.Y(n_124)
);

INVx2_ASAP7_75t_SL g189 ( 
.A(n_124),
.Y(n_189)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_36),
.Y(n_125)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_125),
.Y(n_197)
);

BUFx5_ASAP7_75t_L g126 ( 
.A(n_51),
.Y(n_126)
);

AND2x2_ASAP7_75t_L g151 ( 
.A(n_126),
.B(n_46),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_38),
.Y(n_127)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_127),
.Y(n_175)
);

INVx11_ASAP7_75t_L g128 ( 
.A(n_51),
.Y(n_128)
);

HB1xp67_ASAP7_75t_L g137 ( 
.A(n_128),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_38),
.Y(n_129)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_129),
.Y(n_191)
);

OAI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_101),
.A2(n_48),
.B1(n_29),
.B2(n_23),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_133),
.A2(n_178),
.B1(n_151),
.B2(n_160),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_142),
.B(n_156),
.Y(n_234)
);

HB1xp67_ASAP7_75t_L g144 ( 
.A(n_62),
.Y(n_144)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_144),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_SL g145 ( 
.A(n_94),
.B(n_40),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_SL g223 ( 
.A(n_145),
.B(n_154),
.Y(n_223)
);

AOI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_76),
.A2(n_100),
.B1(n_80),
.B2(n_83),
.Y(n_148)
);

AOI21xp5_ASAP7_75t_L g256 ( 
.A1(n_148),
.A2(n_24),
.B(n_119),
.Y(n_256)
);

CKINVDCx16_ASAP7_75t_R g270 ( 
.A(n_151),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_122),
.B(n_40),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_120),
.B(n_45),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_76),
.B(n_45),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_159),
.B(n_161),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_80),
.B(n_58),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_100),
.B(n_58),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_164),
.B(n_172),
.Y(n_248)
);

HB1xp67_ASAP7_75t_L g169 ( 
.A(n_68),
.Y(n_169)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_169),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_108),
.A2(n_38),
.B1(n_54),
.B2(n_50),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g252 ( 
.A1(n_171),
.A2(n_194),
.B1(n_43),
.B2(n_31),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_74),
.B(n_39),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_110),
.B(n_39),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_173),
.B(n_179),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_88),
.A2(n_56),
.B1(n_42),
.B2(n_46),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_128),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_183),
.B(n_201),
.Y(n_220)
);

AND2x2_ASAP7_75t_L g241 ( 
.A(n_185),
.B(n_69),
.Y(n_241)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_121),
.Y(n_193)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_193),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_111),
.A2(n_47),
.B1(n_41),
.B2(n_54),
.Y(n_194)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_127),
.Y(n_199)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_199),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_102),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_115),
.B(n_47),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g277 ( 
.A(n_203),
.B(n_46),
.Y(n_277)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_129),
.Y(n_207)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_207),
.Y(n_258)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_106),
.Y(n_208)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_208),
.Y(n_260)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_124),
.Y(n_212)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_212),
.Y(n_265)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_69),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_215),
.B(n_184),
.Y(n_227)
);

BUFx12_ASAP7_75t_L g216 ( 
.A(n_107),
.Y(n_216)
);

INVx13_ASAP7_75t_L g226 ( 
.A(n_216),
.Y(n_226)
);

INVx3_ASAP7_75t_L g218 ( 
.A(n_184),
.Y(n_218)
);

BUFx2_ASAP7_75t_L g314 ( 
.A(n_218),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_144),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_219),
.B(n_225),
.Y(n_299)
);

BUFx6f_ASAP7_75t_L g221 ( 
.A(n_135),
.Y(n_221)
);

INVx5_ASAP7_75t_L g320 ( 
.A(n_221),
.Y(n_320)
);

INVx6_ASAP7_75t_L g222 ( 
.A(n_176),
.Y(n_222)
);

INVx4_ASAP7_75t_L g302 ( 
.A(n_222),
.Y(n_302)
);

AND2x4_ASAP7_75t_L g224 ( 
.A(n_130),
.B(n_132),
.Y(n_224)
);

AND2x2_ASAP7_75t_L g327 ( 
.A(n_224),
.B(n_264),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_169),
.Y(n_225)
);

CKINVDCx14_ASAP7_75t_R g330 ( 
.A(n_227),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_136),
.A2(n_112),
.B1(n_118),
.B2(n_117),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_229),
.A2(n_252),
.B1(n_140),
.B2(n_180),
.Y(n_295)
);

AOI22xp33_ASAP7_75t_SL g230 ( 
.A1(n_165),
.A2(n_81),
.B1(n_97),
.B2(n_36),
.Y(n_230)
);

AOI22xp33_ASAP7_75t_SL g350 ( 
.A1(n_230),
.A2(n_232),
.B1(n_239),
.B2(n_249),
.Y(n_350)
);

AOI22xp33_ASAP7_75t_SL g232 ( 
.A1(n_198),
.A2(n_44),
.B1(n_59),
.B2(n_55),
.Y(n_232)
);

INVx2_ASAP7_75t_SL g235 ( 
.A(n_184),
.Y(n_235)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_235),
.Y(n_298)
);

INVx13_ASAP7_75t_L g236 ( 
.A(n_187),
.Y(n_236)
);

BUFx3_ASAP7_75t_L g297 ( 
.A(n_236),
.Y(n_297)
);

INVx5_ASAP7_75t_L g237 ( 
.A(n_190),
.Y(n_237)
);

INVx3_ASAP7_75t_L g322 ( 
.A(n_237),
.Y(n_322)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_139),
.Y(n_238)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_238),
.Y(n_352)
);

AOI22xp33_ASAP7_75t_SL g239 ( 
.A1(n_202),
.A2(n_44),
.B1(n_59),
.B2(n_55),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_149),
.B(n_50),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_SL g301 ( 
.A(n_240),
.B(n_254),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_241),
.B(n_210),
.C(n_157),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_131),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_242),
.B(n_247),
.Y(n_300)
);

INVx2_ASAP7_75t_SL g243 ( 
.A(n_167),
.Y(n_243)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_243),
.Y(n_318)
);

OAI22xp33_ASAP7_75t_SL g244 ( 
.A1(n_133),
.A2(n_77),
.B1(n_65),
.B2(n_98),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_244),
.A2(n_256),
.B1(n_196),
.B2(n_189),
.Y(n_294)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_141),
.Y(n_246)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_246),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_138),
.Y(n_247)
);

AOI22xp33_ASAP7_75t_SL g249 ( 
.A1(n_147),
.A2(n_103),
.B1(n_31),
.B2(n_24),
.Y(n_249)
);

NOR2x1_ASAP7_75t_L g250 ( 
.A(n_146),
.B(n_87),
.Y(n_250)
);

NOR2x1_ASAP7_75t_L g338 ( 
.A(n_250),
.B(n_177),
.Y(n_338)
);

AOI22xp33_ASAP7_75t_L g251 ( 
.A1(n_213),
.A2(n_82),
.B1(n_96),
.B2(n_95),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_L g307 ( 
.A1(n_251),
.A2(n_261),
.B1(n_279),
.B2(n_280),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_153),
.B(n_46),
.Y(n_254)
);

INVx2_ASAP7_75t_SL g255 ( 
.A(n_217),
.Y(n_255)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_255),
.Y(n_321)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_158),
.Y(n_257)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_257),
.Y(n_313)
);

INVx3_ASAP7_75t_L g259 ( 
.A(n_174),
.Y(n_259)
);

INVx4_ASAP7_75t_L g348 ( 
.A(n_259),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_188),
.B(n_0),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_262),
.B(n_276),
.Y(n_304)
);

INVx4_ASAP7_75t_SL g264 ( 
.A(n_187),
.Y(n_264)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_197),
.Y(n_266)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_266),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_155),
.B(n_163),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_267),
.B(n_273),
.Y(n_312)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_214),
.Y(n_268)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_268),
.Y(n_324)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_175),
.Y(n_269)
);

INVx2_ASAP7_75t_L g333 ( 
.A(n_269),
.Y(n_333)
);

INVx4_ASAP7_75t_L g271 ( 
.A(n_190),
.Y(n_271)
);

INVx3_ASAP7_75t_L g325 ( 
.A(n_271),
.Y(n_325)
);

BUFx2_ASAP7_75t_L g272 ( 
.A(n_200),
.Y(n_272)
);

INVx2_ASAP7_75t_L g341 ( 
.A(n_272),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_134),
.B(n_46),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_204),
.Y(n_274)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_274),
.Y(n_347)
);

CKINVDCx12_ASAP7_75t_R g275 ( 
.A(n_174),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_275),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_191),
.B(n_0),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_277),
.B(n_278),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_152),
.B(n_42),
.Y(n_278)
);

AOI22xp33_ASAP7_75t_SL g279 ( 
.A1(n_162),
.A2(n_119),
.B1(n_90),
.B2(n_78),
.Y(n_279)
);

AOI22xp33_ASAP7_75t_L g280 ( 
.A1(n_204),
.A2(n_75),
.B1(n_73),
.B2(n_66),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_SL g281 ( 
.A(n_170),
.B(n_63),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_281),
.B(n_289),
.Y(n_335)
);

CKINVDCx9p33_ASAP7_75t_R g282 ( 
.A(n_206),
.Y(n_282)
);

OR2x2_ASAP7_75t_L g296 ( 
.A(n_282),
.B(n_290),
.Y(n_296)
);

INVx6_ASAP7_75t_L g283 ( 
.A(n_176),
.Y(n_283)
);

INVx3_ASAP7_75t_L g326 ( 
.A(n_283),
.Y(n_326)
);

INVx8_ASAP7_75t_L g284 ( 
.A(n_135),
.Y(n_284)
);

INVx3_ASAP7_75t_L g339 ( 
.A(n_284),
.Y(n_339)
);

INVx4_ASAP7_75t_SL g285 ( 
.A(n_206),
.Y(n_285)
);

AND2x2_ASAP7_75t_L g329 ( 
.A(n_285),
.B(n_291),
.Y(n_329)
);

AOI22xp33_ASAP7_75t_L g286 ( 
.A1(n_205),
.A2(n_7),
.B1(n_15),
.B2(n_14),
.Y(n_286)
);

OAI22xp33_ASAP7_75t_L g309 ( 
.A1(n_286),
.A2(n_157),
.B1(n_210),
.B2(n_195),
.Y(n_309)
);

BUFx2_ASAP7_75t_L g287 ( 
.A(n_205),
.Y(n_287)
);

INVx2_ASAP7_75t_L g346 ( 
.A(n_287),
.Y(n_346)
);

INVx6_ASAP7_75t_L g288 ( 
.A(n_150),
.Y(n_288)
);

INVx3_ASAP7_75t_L g351 ( 
.A(n_288),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_152),
.B(n_6),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_160),
.Y(n_290)
);

INVx3_ASAP7_75t_L g291 ( 
.A(n_211),
.Y(n_291)
);

INVx4_ASAP7_75t_L g292 ( 
.A(n_190),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_292),
.B(n_235),
.Y(n_343)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_209),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_293),
.B(n_189),
.Y(n_319)
);

OAI22xp33_ASAP7_75t_SL g353 ( 
.A1(n_294),
.A2(n_282),
.B1(n_272),
.B2(n_218),
.Y(n_353)
);

OAI22xp5_ASAP7_75t_L g354 ( 
.A1(n_295),
.A2(n_332),
.B1(n_342),
.B2(n_284),
.Y(n_354)
);

FAx1_ASAP7_75t_SL g303 ( 
.A(n_262),
.B(n_137),
.CI(n_148),
.CON(n_303),
.SN(n_303)
);

NOR2xp33_ASAP7_75t_SL g362 ( 
.A(n_303),
.B(n_306),
.Y(n_362)
);

AOI32xp33_ASAP7_75t_L g306 ( 
.A1(n_248),
.A2(n_245),
.A3(n_290),
.B1(n_263),
.B2(n_250),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_261),
.A2(n_209),
.B1(n_180),
.B2(n_140),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g371 ( 
.A1(n_308),
.A2(n_309),
.B1(n_315),
.B2(n_337),
.Y(n_371)
);

OR2x2_ASAP7_75t_L g310 ( 
.A(n_223),
.B(n_192),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_SL g357 ( 
.A(n_310),
.B(n_338),
.Y(n_357)
);

AOI21xp5_ASAP7_75t_SL g311 ( 
.A1(n_241),
.A2(n_137),
.B(n_216),
.Y(n_311)
);

OAI21xp5_ASAP7_75t_L g360 ( 
.A1(n_311),
.A2(n_323),
.B(n_331),
.Y(n_360)
);

OAI22xp33_ASAP7_75t_L g315 ( 
.A1(n_256),
.A2(n_150),
.B1(n_195),
.B2(n_186),
.Y(n_315)
);

CKINVDCx16_ASAP7_75t_R g386 ( 
.A(n_319),
.Y(n_386)
);

OAI21xp5_ASAP7_75t_L g323 ( 
.A1(n_241),
.A2(n_143),
.B(n_196),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_L g359 ( 
.A(n_328),
.B(n_255),
.Y(n_359)
);

AOI22xp5_ASAP7_75t_SL g331 ( 
.A1(n_270),
.A2(n_196),
.B1(n_143),
.B2(n_182),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_L g332 ( 
.A1(n_229),
.A2(n_186),
.B1(n_182),
.B2(n_181),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_276),
.B(n_181),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_336),
.B(n_344),
.Y(n_385)
);

OAI22xp5_ASAP7_75t_SL g337 ( 
.A1(n_234),
.A2(n_166),
.B1(n_177),
.B2(n_168),
.Y(n_337)
);

OAI22xp5_ASAP7_75t_SL g340 ( 
.A1(n_220),
.A2(n_166),
.B1(n_1),
.B2(n_2),
.Y(n_340)
);

AOI22xp5_ASAP7_75t_L g389 ( 
.A1(n_340),
.A2(n_345),
.B1(n_243),
.B2(n_293),
.Y(n_389)
);

AOI22xp5_ASAP7_75t_L g342 ( 
.A1(n_224),
.A2(n_12),
.B1(n_15),
.B2(n_14),
.Y(n_342)
);

CKINVDCx16_ASAP7_75t_R g398 ( 
.A(n_343),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_224),
.B(n_0),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_SL g345 ( 
.A1(n_238),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_345)
);

OAI22xp33_ASAP7_75t_SL g349 ( 
.A1(n_246),
.A2(n_5),
.B1(n_12),
.B2(n_13),
.Y(n_349)
);

AOI22xp5_ASAP7_75t_SL g380 ( 
.A1(n_349),
.A2(n_235),
.B1(n_255),
.B2(n_243),
.Y(n_380)
);

AOI22xp5_ASAP7_75t_L g422 ( 
.A1(n_353),
.A2(n_354),
.B1(n_377),
.B2(n_309),
.Y(n_422)
);

AND2x6_ASAP7_75t_L g355 ( 
.A(n_338),
.B(n_242),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_L g404 ( 
.A(n_355),
.B(n_366),
.Y(n_404)
);

INVx1_ASAP7_75t_SL g356 ( 
.A(n_327),
.Y(n_356)
);

INVx1_ASAP7_75t_SL g401 ( 
.A(n_356),
.Y(n_401)
);

AND2x2_ASAP7_75t_L g358 ( 
.A(n_327),
.B(n_224),
.Y(n_358)
);

INVxp67_ASAP7_75t_L g426 ( 
.A(n_358),
.Y(n_426)
);

XOR2xp5_ASAP7_75t_L g411 ( 
.A(n_359),
.B(n_312),
.Y(n_411)
);

CKINVDCx12_ASAP7_75t_R g361 ( 
.A(n_329),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_361),
.Y(n_432)
);

INVx2_ASAP7_75t_L g363 ( 
.A(n_321),
.Y(n_363)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_363),
.Y(n_409)
);

AOI22xp33_ASAP7_75t_SL g364 ( 
.A1(n_308),
.A2(n_287),
.B1(n_259),
.B2(n_292),
.Y(n_364)
);

BUFx3_ASAP7_75t_L g408 ( 
.A(n_364),
.Y(n_408)
);

INVx2_ASAP7_75t_L g365 ( 
.A(n_321),
.Y(n_365)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_365),
.Y(n_410)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_299),
.Y(n_366)
);

INVx13_ASAP7_75t_L g367 ( 
.A(n_297),
.Y(n_367)
);

BUFx2_ASAP7_75t_SL g406 ( 
.A(n_367),
.Y(n_406)
);

INVx5_ASAP7_75t_L g368 ( 
.A(n_302),
.Y(n_368)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_368),
.Y(n_414)
);

NOR2xp33_ASAP7_75t_L g369 ( 
.A(n_330),
.B(n_247),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_SL g434 ( 
.A(n_369),
.B(n_375),
.Y(n_434)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_305),
.Y(n_370)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_370),
.Y(n_420)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_313),
.Y(n_372)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_372),
.Y(n_424)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_328),
.B(n_311),
.C(n_323),
.Y(n_373)
);

MAJIxp5_ASAP7_75t_L g400 ( 
.A(n_373),
.B(n_397),
.C(n_344),
.Y(n_400)
);

INVx2_ASAP7_75t_L g374 ( 
.A(n_318),
.Y(n_374)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_374),
.Y(n_436)
);

NOR2xp33_ASAP7_75t_L g375 ( 
.A(n_301),
.B(n_266),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_L g376 ( 
.A(n_300),
.B(n_257),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_SL g437 ( 
.A(n_376),
.B(n_382),
.Y(n_437)
);

OAI22xp5_ASAP7_75t_SL g377 ( 
.A1(n_295),
.A2(n_253),
.B1(n_258),
.B2(n_269),
.Y(n_377)
);

AND2x2_ASAP7_75t_L g378 ( 
.A(n_327),
.B(n_225),
.Y(n_378)
);

XNOR2xp5_ASAP7_75t_L g412 ( 
.A(n_378),
.B(n_342),
.Y(n_412)
);

BUFx12f_ASAP7_75t_L g379 ( 
.A(n_297),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_L g407 ( 
.A(n_379),
.B(n_390),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_380),
.B(n_389),
.Y(n_405)
);

INVx13_ASAP7_75t_L g381 ( 
.A(n_334),
.Y(n_381)
);

CKINVDCx20_ASAP7_75t_R g417 ( 
.A(n_381),
.Y(n_417)
);

NOR2xp33_ASAP7_75t_L g382 ( 
.A(n_310),
.B(n_219),
.Y(n_382)
);

CKINVDCx12_ASAP7_75t_R g383 ( 
.A(n_329),
.Y(n_383)
);

CKINVDCx20_ASAP7_75t_R g429 ( 
.A(n_383),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_SL g384 ( 
.A(n_335),
.B(n_231),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_SL g416 ( 
.A(n_384),
.B(n_387),
.Y(n_416)
);

AO22x1_ASAP7_75t_L g387 ( 
.A1(n_315),
.A2(n_231),
.B1(n_228),
.B2(n_268),
.Y(n_387)
);

BUFx8_ASAP7_75t_L g388 ( 
.A(n_296),
.Y(n_388)
);

CKINVDCx20_ASAP7_75t_R g431 ( 
.A(n_388),
.Y(n_431)
);

AND2x6_ASAP7_75t_L g390 ( 
.A(n_316),
.B(n_226),
.Y(n_390)
);

CKINVDCx20_ASAP7_75t_R g391 ( 
.A(n_319),
.Y(n_391)
);

NOR2xp33_ASAP7_75t_L g428 ( 
.A(n_391),
.B(n_333),
.Y(n_428)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_317),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_392),
.B(n_394),
.Y(n_413)
);

INVx13_ASAP7_75t_L g393 ( 
.A(n_298),
.Y(n_393)
);

CKINVDCx20_ASAP7_75t_R g433 ( 
.A(n_393),
.Y(n_433)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_352),
.Y(n_394)
);

OAI21xp5_ASAP7_75t_L g395 ( 
.A1(n_296),
.A2(n_228),
.B(n_233),
.Y(n_395)
);

AOI21xp5_ASAP7_75t_SL g419 ( 
.A1(n_395),
.A2(n_329),
.B(n_324),
.Y(n_419)
);

AOI22xp5_ASAP7_75t_L g396 ( 
.A1(n_307),
.A2(n_253),
.B1(n_258),
.B2(n_274),
.Y(n_396)
);

OAI22xp5_ASAP7_75t_L g421 ( 
.A1(n_396),
.A2(n_347),
.B1(n_333),
.B2(n_318),
.Y(n_421)
);

MAJIxp5_ASAP7_75t_L g397 ( 
.A(n_304),
.B(n_233),
.C(n_265),
.Y(n_397)
);

OAI22xp5_ASAP7_75t_SL g399 ( 
.A1(n_371),
.A2(n_294),
.B1(n_332),
.B2(n_350),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_399),
.B(n_402),
.Y(n_448)
);

MAJIxp5_ASAP7_75t_L g452 ( 
.A(n_400),
.B(n_425),
.C(n_435),
.Y(n_452)
);

OAI22xp5_ASAP7_75t_SL g402 ( 
.A1(n_371),
.A2(n_304),
.B1(n_336),
.B2(n_303),
.Y(n_402)
);

AOI21xp5_ASAP7_75t_L g403 ( 
.A1(n_360),
.A2(n_303),
.B(n_331),
.Y(n_403)
);

AOI21xp5_ASAP7_75t_L g442 ( 
.A1(n_403),
.A2(n_360),
.B(n_395),
.Y(n_442)
);

XNOR2xp5_ASAP7_75t_SL g445 ( 
.A(n_411),
.B(n_415),
.Y(n_445)
);

AND2x2_ASAP7_75t_L g446 ( 
.A(n_412),
.B(n_421),
.Y(n_446)
);

XNOR2xp5_ASAP7_75t_L g415 ( 
.A(n_359),
.B(n_337),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_391),
.B(n_340),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_418),
.B(n_427),
.Y(n_453)
);

OAI21xp5_ASAP7_75t_L g438 ( 
.A1(n_419),
.A2(n_358),
.B(n_356),
.Y(n_438)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_422),
.Y(n_449)
);

AOI22xp33_ASAP7_75t_L g423 ( 
.A1(n_366),
.A2(n_326),
.B1(n_302),
.B2(n_339),
.Y(n_423)
);

AOI22xp33_ASAP7_75t_SL g467 ( 
.A1(n_423),
.A2(n_298),
.B1(n_379),
.B2(n_377),
.Y(n_467)
);

MAJIxp5_ASAP7_75t_L g425 ( 
.A(n_373),
.B(n_260),
.C(n_265),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_386),
.B(n_385),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_428),
.B(n_430),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_386),
.B(n_345),
.Y(n_430)
);

XNOR2xp5_ASAP7_75t_L g435 ( 
.A(n_385),
.B(n_325),
.Y(n_435)
);

AO22x1_ASAP7_75t_L g484 ( 
.A1(n_438),
.A2(n_426),
.B1(n_419),
.B2(n_401),
.Y(n_484)
);

XOR2xp5_ASAP7_75t_L g439 ( 
.A(n_411),
.B(n_397),
.Y(n_439)
);

MAJIxp5_ASAP7_75t_L g500 ( 
.A(n_439),
.B(n_440),
.C(n_447),
.Y(n_500)
);

XNOR2xp5_ASAP7_75t_L g440 ( 
.A(n_400),
.B(n_427),
.Y(n_440)
);

NOR2x1_ASAP7_75t_L g441 ( 
.A(n_432),
.B(n_362),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_SL g478 ( 
.A(n_441),
.B(n_412),
.Y(n_478)
);

AOI21xp5_ASAP7_75t_L g505 ( 
.A1(n_442),
.A2(n_461),
.B(n_383),
.Y(n_505)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_409),
.Y(n_443)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_443),
.Y(n_483)
);

OAI22xp5_ASAP7_75t_L g444 ( 
.A1(n_418),
.A2(n_396),
.B1(n_389),
.B2(n_362),
.Y(n_444)
);

AOI22xp5_ASAP7_75t_L g486 ( 
.A1(n_444),
.A2(n_463),
.B1(n_464),
.B2(n_471),
.Y(n_486)
);

XNOR2xp5_ASAP7_75t_L g447 ( 
.A(n_425),
.B(n_378),
.Y(n_447)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_413),
.Y(n_450)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_450),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_SL g451 ( 
.A(n_434),
.B(n_398),
.Y(n_451)
);

NAND3xp33_ASAP7_75t_L g481 ( 
.A(n_451),
.B(n_460),
.C(n_470),
.Y(n_481)
);

HB1xp67_ASAP7_75t_L g454 ( 
.A(n_406),
.Y(n_454)
);

CKINVDCx20_ASAP7_75t_R g479 ( 
.A(n_454),
.Y(n_479)
);

INVx13_ASAP7_75t_L g455 ( 
.A(n_432),
.Y(n_455)
);

CKINVDCx16_ASAP7_75t_R g499 ( 
.A(n_455),
.Y(n_499)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_413),
.Y(n_456)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_456),
.Y(n_492)
);

CKINVDCx20_ASAP7_75t_R g457 ( 
.A(n_416),
.Y(n_457)
);

NOR2xp33_ASAP7_75t_L g473 ( 
.A(n_457),
.B(n_458),
.Y(n_473)
);

CKINVDCx16_ASAP7_75t_R g458 ( 
.A(n_437),
.Y(n_458)
);

AND2x6_ASAP7_75t_L g459 ( 
.A(n_404),
.B(n_355),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_459),
.B(n_465),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_SL g460 ( 
.A(n_437),
.B(n_398),
.Y(n_460)
);

AOI21xp5_ASAP7_75t_L g461 ( 
.A1(n_403),
.A2(n_357),
.B(n_388),
.Y(n_461)
);

OAI22xp5_ASAP7_75t_L g463 ( 
.A1(n_422),
.A2(n_354),
.B1(n_387),
.B2(n_380),
.Y(n_463)
);

OAI22xp5_ASAP7_75t_SL g464 ( 
.A1(n_405),
.A2(n_387),
.B1(n_390),
.B2(n_392),
.Y(n_464)
);

AND2x6_ASAP7_75t_L g465 ( 
.A(n_407),
.B(n_388),
.Y(n_465)
);

CKINVDCx20_ASAP7_75t_R g466 ( 
.A(n_416),
.Y(n_466)
);

NOR2xp33_ASAP7_75t_L g485 ( 
.A(n_466),
.B(n_469),
.Y(n_485)
);

INVxp67_ASAP7_75t_L g482 ( 
.A(n_467),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_431),
.B(n_388),
.Y(n_468)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_468),
.Y(n_503)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_420),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_SL g470 ( 
.A(n_417),
.B(n_394),
.Y(n_470)
);

OAI22xp5_ASAP7_75t_L g471 ( 
.A1(n_405),
.A2(n_372),
.B1(n_370),
.B2(n_358),
.Y(n_471)
);

NOR2xp33_ASAP7_75t_L g472 ( 
.A(n_417),
.B(n_314),
.Y(n_472)
);

NOR2xp33_ASAP7_75t_SL g488 ( 
.A(n_472),
.B(n_379),
.Y(n_488)
);

NOR2xp33_ASAP7_75t_L g474 ( 
.A(n_458),
.B(n_440),
.Y(n_474)
);

NOR2xp33_ASAP7_75t_SL g520 ( 
.A(n_474),
.B(n_493),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_457),
.B(n_431),
.Y(n_476)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_476),
.Y(n_509)
);

XOR2xp5_ASAP7_75t_L g477 ( 
.A(n_439),
.B(n_445),
.Y(n_477)
);

XOR2xp5_ASAP7_75t_L g532 ( 
.A(n_477),
.B(n_490),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_L g511 ( 
.A(n_478),
.B(n_489),
.Y(n_511)
);

OR2x2_ASAP7_75t_L g480 ( 
.A(n_468),
.B(n_402),
.Y(n_480)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_480),
.Y(n_517)
);

XNOR2x1_ASAP7_75t_L g512 ( 
.A(n_484),
.B(n_471),
.Y(n_512)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_488),
.Y(n_535)
);

INVxp67_ASAP7_75t_L g489 ( 
.A(n_441),
.Y(n_489)
);

XNOR2xp5_ASAP7_75t_L g490 ( 
.A(n_452),
.B(n_435),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_SL g491 ( 
.A(n_466),
.B(n_430),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_491),
.B(n_502),
.Y(n_530)
);

NOR2xp33_ASAP7_75t_SL g493 ( 
.A(n_450),
.B(n_429),
.Y(n_493)
);

AOI22xp33_ASAP7_75t_SL g494 ( 
.A1(n_449),
.A2(n_408),
.B1(n_399),
.B2(n_429),
.Y(n_494)
);

OAI22xp5_ASAP7_75t_SL g514 ( 
.A1(n_494),
.A2(n_461),
.B1(n_448),
.B2(n_455),
.Y(n_514)
);

OAI22xp5_ASAP7_75t_L g495 ( 
.A1(n_449),
.A2(n_408),
.B1(n_426),
.B2(n_401),
.Y(n_495)
);

OAI22xp5_ASAP7_75t_L g510 ( 
.A1(n_495),
.A2(n_501),
.B1(n_469),
.B2(n_443),
.Y(n_510)
);

NOR2xp33_ASAP7_75t_SL g496 ( 
.A(n_456),
.B(n_420),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_SL g518 ( 
.A(n_496),
.B(n_504),
.Y(n_518)
);

OAI21xp5_ASAP7_75t_L g497 ( 
.A1(n_442),
.A2(n_378),
.B(n_424),
.Y(n_497)
);

INVxp67_ASAP7_75t_L g521 ( 
.A(n_497),
.Y(n_521)
);

AOI22xp5_ASAP7_75t_L g498 ( 
.A1(n_463),
.A2(n_421),
.B1(n_415),
.B2(n_424),
.Y(n_498)
);

OAI22xp5_ASAP7_75t_SL g516 ( 
.A1(n_498),
.A2(n_462),
.B1(n_453),
.B2(n_446),
.Y(n_516)
);

OAI22xp5_ASAP7_75t_L g501 ( 
.A1(n_448),
.A2(n_433),
.B1(n_414),
.B2(n_436),
.Y(n_501)
);

INVxp67_ASAP7_75t_L g502 ( 
.A(n_444),
.Y(n_502)
);

NOR2xp33_ASAP7_75t_L g504 ( 
.A(n_453),
.B(n_433),
.Y(n_504)
);

INVxp67_ASAP7_75t_L g525 ( 
.A(n_505),
.Y(n_525)
);

FAx1_ASAP7_75t_L g506 ( 
.A(n_438),
.B(n_361),
.CI(n_381),
.CON(n_506),
.SN(n_506)
);

NOR2xp33_ASAP7_75t_L g522 ( 
.A(n_506),
.B(n_464),
.Y(n_522)
);

MAJIxp5_ASAP7_75t_L g507 ( 
.A(n_500),
.B(n_452),
.C(n_447),
.Y(n_507)
);

MAJIxp5_ASAP7_75t_L g538 ( 
.A(n_507),
.B(n_508),
.C(n_523),
.Y(n_538)
);

MAJIxp5_ASAP7_75t_L g508 ( 
.A(n_500),
.B(n_490),
.C(n_477),
.Y(n_508)
);

AOI22xp5_ASAP7_75t_L g540 ( 
.A1(n_510),
.A2(n_514),
.B1(n_516),
.B2(n_519),
.Y(n_540)
);

XNOR2x1_ASAP7_75t_SL g556 ( 
.A(n_512),
.B(n_506),
.Y(n_556)
);

XNOR2xp5_ASAP7_75t_L g513 ( 
.A(n_484),
.B(n_445),
.Y(n_513)
);

XNOR2xp5_ASAP7_75t_L g539 ( 
.A(n_513),
.B(n_533),
.Y(n_539)
);

XNOR2xp5_ASAP7_75t_SL g515 ( 
.A(n_478),
.B(n_473),
.Y(n_515)
);

XOR2xp5_ASAP7_75t_L g552 ( 
.A(n_515),
.B(n_485),
.Y(n_552)
);

OAI22xp5_ASAP7_75t_SL g519 ( 
.A1(n_486),
.A2(n_462),
.B1(n_446),
.B2(n_465),
.Y(n_519)
);

AOI21x1_ASAP7_75t_L g561 ( 
.A1(n_522),
.A2(n_488),
.B(n_479),
.Y(n_561)
);

MAJIxp5_ASAP7_75t_L g523 ( 
.A(n_497),
.B(n_446),
.C(n_414),
.Y(n_523)
);

MAJIxp5_ASAP7_75t_L g524 ( 
.A(n_505),
.B(n_436),
.C(n_410),
.Y(n_524)
);

MAJIxp5_ASAP7_75t_L g542 ( 
.A(n_524),
.B(n_527),
.C(n_529),
.Y(n_542)
);

OAI22xp5_ASAP7_75t_SL g526 ( 
.A1(n_486),
.A2(n_459),
.B1(n_410),
.B2(n_409),
.Y(n_526)
);

AOI22xp5_ASAP7_75t_L g543 ( 
.A1(n_526),
.A2(n_528),
.B1(n_495),
.B2(n_509),
.Y(n_543)
);

MAJIxp5_ASAP7_75t_L g527 ( 
.A(n_498),
.B(n_325),
.C(n_322),
.Y(n_527)
);

OAI22xp5_ASAP7_75t_SL g528 ( 
.A1(n_480),
.A2(n_368),
.B1(n_326),
.B2(n_374),
.Y(n_528)
);

MAJIxp5_ASAP7_75t_L g529 ( 
.A(n_487),
.B(n_322),
.C(n_365),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_SL g531 ( 
.A(n_475),
.B(n_363),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_531),
.B(n_473),
.Y(n_537)
);

XNOR2xp5_ASAP7_75t_L g533 ( 
.A(n_484),
.B(n_339),
.Y(n_533)
);

XNOR2xp5_ASAP7_75t_L g534 ( 
.A(n_476),
.B(n_291),
.Y(n_534)
);

XNOR2xp5_ASAP7_75t_L g551 ( 
.A(n_534),
.B(n_483),
.Y(n_551)
);

MAJIxp5_ASAP7_75t_L g536 ( 
.A(n_487),
.B(n_314),
.C(n_341),
.Y(n_536)
);

MAJIxp5_ASAP7_75t_L g544 ( 
.A(n_536),
.B(n_499),
.C(n_483),
.Y(n_544)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_537),
.Y(n_573)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_518),
.Y(n_541)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_541),
.Y(n_576)
);

INVxp67_ASAP7_75t_L g566 ( 
.A(n_543),
.Y(n_566)
);

XNOR2xp5_ASAP7_75t_L g578 ( 
.A(n_544),
.B(n_529),
.Y(n_578)
);

MAJIxp5_ASAP7_75t_L g545 ( 
.A(n_507),
.B(n_503),
.C(n_475),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_L g562 ( 
.A(n_545),
.B(n_547),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_L g546 ( 
.A(n_535),
.B(n_481),
.Y(n_546)
);

CKINVDCx14_ASAP7_75t_R g568 ( 
.A(n_546),
.Y(n_568)
);

MAJIxp5_ASAP7_75t_L g547 ( 
.A(n_532),
.B(n_503),
.C(n_501),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_534),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_L g570 ( 
.A(n_548),
.B(n_550),
.Y(n_570)
);

NOR2xp33_ASAP7_75t_SL g549 ( 
.A(n_511),
.B(n_493),
.Y(n_549)
);

NOR2xp33_ASAP7_75t_L g575 ( 
.A(n_549),
.B(n_555),
.Y(n_575)
);

HB1xp67_ASAP7_75t_L g550 ( 
.A(n_536),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g571 ( 
.A(n_551),
.B(n_553),
.Y(n_571)
);

XNOR2xp5_ASAP7_75t_SL g574 ( 
.A(n_552),
.B(n_556),
.Y(n_574)
);

CKINVDCx20_ASAP7_75t_R g553 ( 
.A(n_530),
.Y(n_553)
);

AOI22xp5_ASAP7_75t_L g554 ( 
.A1(n_526),
.A2(n_492),
.B1(n_482),
.B2(n_496),
.Y(n_554)
);

HB1xp67_ASAP7_75t_L g577 ( 
.A(n_554),
.Y(n_577)
);

OAI211xp5_ASAP7_75t_L g555 ( 
.A1(n_521),
.A2(n_485),
.B(n_504),
.C(n_492),
.Y(n_555)
);

NOR2xp33_ASAP7_75t_L g557 ( 
.A(n_520),
.B(n_479),
.Y(n_557)
);

CKINVDCx20_ASAP7_75t_R g565 ( 
.A(n_557),
.Y(n_565)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_517),
.Y(n_558)
);

NOR2xp33_ASAP7_75t_L g579 ( 
.A(n_558),
.B(n_533),
.Y(n_579)
);

OAI22xp5_ASAP7_75t_SL g559 ( 
.A1(n_521),
.A2(n_480),
.B1(n_491),
.B2(n_506),
.Y(n_559)
);

AOI22xp5_ASAP7_75t_SL g572 ( 
.A1(n_559),
.A2(n_525),
.B1(n_528),
.B2(n_516),
.Y(n_572)
);

MAJIxp5_ASAP7_75t_L g560 ( 
.A(n_532),
.B(n_499),
.C(n_506),
.Y(n_560)
);

MAJIxp5_ASAP7_75t_L g564 ( 
.A(n_560),
.B(n_524),
.C(n_523),
.Y(n_564)
);

OAI21xp5_ASAP7_75t_L g581 ( 
.A1(n_561),
.A2(n_525),
.B(n_512),
.Y(n_581)
);

XOR2xp5_ASAP7_75t_L g563 ( 
.A(n_547),
.B(n_508),
.Y(n_563)
);

XNOR2xp5_ASAP7_75t_L g585 ( 
.A(n_563),
.B(n_564),
.Y(n_585)
);

MAJIxp5_ASAP7_75t_L g567 ( 
.A(n_538),
.B(n_527),
.C(n_519),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_L g586 ( 
.A(n_567),
.B(n_578),
.Y(n_586)
);

XOR2xp5_ASAP7_75t_L g569 ( 
.A(n_539),
.B(n_513),
.Y(n_569)
);

XOR2xp5_ASAP7_75t_L g594 ( 
.A(n_569),
.B(n_572),
.Y(n_594)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_579),
.Y(n_583)
);

XNOR2xp5_ASAP7_75t_L g580 ( 
.A(n_538),
.B(n_515),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_L g595 ( 
.A(n_580),
.B(n_581),
.Y(n_595)
);

MAJIxp5_ASAP7_75t_L g582 ( 
.A(n_567),
.B(n_545),
.C(n_542),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_L g601 ( 
.A(n_582),
.B(n_589),
.Y(n_601)
);

OAI21x1_ASAP7_75t_SL g584 ( 
.A1(n_575),
.A2(n_554),
.B(n_540),
.Y(n_584)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_584),
.Y(n_604)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_576),
.Y(n_587)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_587),
.Y(n_607)
);

NOR2xp33_ASAP7_75t_SL g588 ( 
.A(n_565),
.B(n_552),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_SL g603 ( 
.A(n_588),
.B(n_590),
.Y(n_603)
);

FAx1_ASAP7_75t_SL g589 ( 
.A(n_581),
.B(n_560),
.CI(n_559),
.CON(n_589),
.SN(n_589)
);

MAJIxp5_ASAP7_75t_L g590 ( 
.A(n_578),
.B(n_542),
.C(n_540),
.Y(n_590)
);

BUFx2_ASAP7_75t_L g591 ( 
.A(n_573),
.Y(n_591)
);

NOR2xp33_ASAP7_75t_L g606 ( 
.A(n_591),
.B(n_593),
.Y(n_606)
);

NOR2xp33_ASAP7_75t_L g592 ( 
.A(n_568),
.B(n_543),
.Y(n_592)
);

XNOR2xp5_ASAP7_75t_L g609 ( 
.A(n_592),
.B(n_596),
.Y(n_609)
);

BUFx24_ASAP7_75t_SL g593 ( 
.A(n_580),
.Y(n_593)
);

MAJIxp5_ASAP7_75t_L g596 ( 
.A(n_563),
.B(n_544),
.C(n_551),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_571),
.Y(n_597)
);

AOI22xp5_ASAP7_75t_L g600 ( 
.A1(n_597),
.A2(n_577),
.B1(n_570),
.B2(n_566),
.Y(n_600)
);

OA22x2_ASAP7_75t_L g598 ( 
.A1(n_572),
.A2(n_556),
.B1(n_539),
.B2(n_351),
.Y(n_598)
);

INVxp67_ASAP7_75t_L g605 ( 
.A(n_598),
.Y(n_605)
);

MAJIxp5_ASAP7_75t_L g599 ( 
.A(n_586),
.B(n_590),
.C(n_582),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_L g613 ( 
.A(n_599),
.B(n_600),
.Y(n_613)
);

OAI21xp5_ASAP7_75t_L g602 ( 
.A1(n_595),
.A2(n_562),
.B(n_564),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_L g614 ( 
.A(n_602),
.B(n_608),
.Y(n_614)
);

MAJIxp5_ASAP7_75t_L g608 ( 
.A(n_585),
.B(n_566),
.C(n_569),
.Y(n_608)
);

MAJIxp5_ASAP7_75t_L g610 ( 
.A(n_585),
.B(n_574),
.C(n_351),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_SL g615 ( 
.A(n_610),
.B(n_611),
.Y(n_615)
);

MAJIxp5_ASAP7_75t_L g611 ( 
.A(n_596),
.B(n_574),
.C(n_341),
.Y(n_611)
);

XNOR2xp5_ASAP7_75t_L g612 ( 
.A(n_594),
.B(n_346),
.Y(n_612)
);

NOR2xp33_ASAP7_75t_L g622 ( 
.A(n_612),
.B(n_379),
.Y(n_622)
);

NOR2xp33_ASAP7_75t_L g616 ( 
.A(n_599),
.B(n_591),
.Y(n_616)
);

AOI21xp5_ASAP7_75t_L g627 ( 
.A1(n_616),
.A2(n_617),
.B(n_618),
.Y(n_627)
);

OAI21xp5_ASAP7_75t_SL g617 ( 
.A1(n_601),
.A2(n_583),
.B(n_589),
.Y(n_617)
);

OAI21x1_ASAP7_75t_L g618 ( 
.A1(n_606),
.A2(n_598),
.B(n_594),
.Y(n_618)
);

NOR2xp33_ASAP7_75t_L g619 ( 
.A(n_609),
.B(n_598),
.Y(n_619)
);

XNOR2xp5_ASAP7_75t_L g625 ( 
.A(n_619),
.B(n_620),
.Y(n_625)
);

OAI21x1_ASAP7_75t_L g620 ( 
.A1(n_603),
.A2(n_393),
.B(n_367),
.Y(n_620)
);

XNOR2xp5_ASAP7_75t_L g621 ( 
.A(n_611),
.B(n_608),
.Y(n_621)
);

MAJIxp5_ASAP7_75t_L g626 ( 
.A(n_621),
.B(n_605),
.C(n_607),
.Y(n_626)
);

MAJIxp5_ASAP7_75t_L g623 ( 
.A(n_622),
.B(n_610),
.C(n_612),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_L g631 ( 
.A(n_623),
.B(n_626),
.Y(n_631)
);

OAI21xp5_ASAP7_75t_L g624 ( 
.A1(n_614),
.A2(n_613),
.B(n_604),
.Y(n_624)
);

AOI21xp5_ASAP7_75t_L g630 ( 
.A1(n_624),
.A2(n_628),
.B(n_629),
.Y(n_630)
);

OAI21xp5_ASAP7_75t_SL g628 ( 
.A1(n_615),
.A2(n_605),
.B(n_622),
.Y(n_628)
);

MAJIxp5_ASAP7_75t_L g629 ( 
.A(n_614),
.B(n_221),
.C(n_346),
.Y(n_629)
);

AOI21x1_ASAP7_75t_L g632 ( 
.A1(n_627),
.A2(n_236),
.B(n_260),
.Y(n_632)
);

AOI21xp5_ASAP7_75t_L g635 ( 
.A1(n_632),
.A2(n_633),
.B(n_271),
.Y(n_635)
);

OAI21xp5_ASAP7_75t_SL g633 ( 
.A1(n_623),
.A2(n_226),
.B(n_348),
.Y(n_633)
);

AOI322xp5_ASAP7_75t_L g634 ( 
.A1(n_630),
.A2(n_625),
.A3(n_320),
.B1(n_237),
.B2(n_348),
.C1(n_283),
.C2(n_222),
.Y(n_634)
);

O2A1O1Ixp33_ASAP7_75t_SL g637 ( 
.A1(n_634),
.A2(n_264),
.B(n_285),
.C(n_320),
.Y(n_637)
);

NOR2xp33_ASAP7_75t_L g636 ( 
.A(n_635),
.B(n_631),
.Y(n_636)
);

AOI22xp33_ASAP7_75t_SL g638 ( 
.A1(n_636),
.A2(n_637),
.B1(n_288),
.B2(n_5),
.Y(n_638)
);

AOI21xp5_ASAP7_75t_SL g639 ( 
.A1(n_638),
.A2(n_16),
.B(n_5),
.Y(n_639)
);

XNOR2xp5_ASAP7_75t_L g640 ( 
.A(n_639),
.B(n_12),
.Y(n_640)
);

AOI21xp5_ASAP7_75t_L g641 ( 
.A1(n_640),
.A2(n_1),
.B(n_2),
.Y(n_641)
);


endmodule