module fake_jpeg_14884_n_91 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_91);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_91;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_44;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_36;
wire n_62;
wire n_43;
wire n_82;

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_5),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_32),
.Y(n_35)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_15),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_2),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_11),
.Y(n_38)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_5),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_10),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_2),
.Y(n_41)
);

INVx1_ASAP7_75t_SL g42 ( 
.A(n_4),
.Y(n_42)
);

BUFx24_ASAP7_75t_L g43 ( 
.A(n_1),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_20),
.Y(n_44)
);

BUFx24_ASAP7_75t_L g45 ( 
.A(n_43),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_45),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_41),
.B(n_0),
.Y(n_46)
);

OR2x2_ASAP7_75t_L g58 ( 
.A(n_46),
.B(n_33),
.Y(n_58)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_43),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_47),
.B(n_48),
.Y(n_53)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_34),
.Y(n_49)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_49),
.Y(n_57)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_39),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_50),
.B(n_51),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_35),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_52),
.B(n_0),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_49),
.A2(n_42),
.B1(n_44),
.B2(n_35),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_54),
.A2(n_55),
.B1(n_63),
.B2(n_7),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_L g55 ( 
.A1(n_52),
.A2(n_44),
.B1(n_34),
.B2(n_37),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_58),
.B(n_6),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_45),
.B(n_38),
.Y(n_59)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_59),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_60),
.B(n_62),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_46),
.B(n_3),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_50),
.A2(n_40),
.B1(n_4),
.B2(n_3),
.Y(n_63)
);

OR2x2_ASAP7_75t_L g74 ( 
.A(n_64),
.B(n_71),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_65),
.A2(n_61),
.B1(n_22),
.B2(n_23),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_58),
.B(n_8),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_67),
.B(n_70),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_L g68 ( 
.A1(n_57),
.A2(n_9),
.B1(n_12),
.B2(n_13),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_68),
.A2(n_17),
.B1(n_18),
.B2(n_19),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_56),
.B(n_14),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_53),
.B(n_16),
.Y(n_71)
);

NAND3xp33_ASAP7_75t_L g72 ( 
.A(n_69),
.B(n_55),
.C(n_54),
.Y(n_72)
);

XNOR2x2_ASAP7_75t_SL g78 ( 
.A(n_72),
.B(n_68),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_73),
.B(n_75),
.Y(n_77)
);

XOR2xp5_ASAP7_75t_L g81 ( 
.A(n_78),
.B(n_69),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_74),
.B(n_66),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_79),
.Y(n_80)
);

OAI21xp5_ASAP7_75t_L g82 ( 
.A1(n_81),
.A2(n_77),
.B(n_76),
.Y(n_82)
);

AOI21xp5_ASAP7_75t_SL g84 ( 
.A1(n_82),
.A2(n_83),
.B(n_76),
.Y(n_84)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_80),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_84),
.B(n_21),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_85),
.B(n_24),
.Y(n_86)
);

AOI21xp33_ASAP7_75t_L g87 ( 
.A1(n_86),
.A2(n_25),
.B(n_26),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_87),
.B(n_27),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_SL g89 ( 
.A1(n_88),
.A2(n_28),
.B(n_29),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_89),
.B(n_30),
.Y(n_90)
);

XOR2xp5_ASAP7_75t_L g91 ( 
.A(n_90),
.B(n_31),
.Y(n_91)
);


endmodule