module fake_jpeg_19731_n_170 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_170);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_170;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_93;
wire n_54;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_38),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_44),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_2),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_15),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_8),
.Y(n_55)
);

BUFx2_ASAP7_75t_L g56 ( 
.A(n_17),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_37),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_6),
.Y(n_58)
);

BUFx5_ASAP7_75t_L g59 ( 
.A(n_21),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_35),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_2),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_16),
.Y(n_62)
);

BUFx12_ASAP7_75t_L g63 ( 
.A(n_24),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_47),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_8),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_19),
.Y(n_66)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_1),
.Y(n_67)
);

BUFx5_ASAP7_75t_L g68 ( 
.A(n_18),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_46),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_12),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_32),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_41),
.Y(n_72)
);

INVx13_ASAP7_75t_L g73 ( 
.A(n_40),
.Y(n_73)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_50),
.Y(n_74)
);

BUFx24_ASAP7_75t_L g75 ( 
.A(n_22),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_13),
.Y(n_76)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_45),
.Y(n_77)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_43),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_42),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_0),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_53),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_81),
.B(n_82),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_55),
.Y(n_82)
);

INVx2_ASAP7_75t_R g83 ( 
.A(n_75),
.Y(n_83)
);

AOI21xp33_ASAP7_75t_L g98 ( 
.A1(n_83),
.A2(n_63),
.B(n_65),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_61),
.B(n_0),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_84),
.B(n_86),
.Y(n_91)
);

BUFx2_ASAP7_75t_L g85 ( 
.A(n_75),
.Y(n_85)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_85),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_58),
.Y(n_86)
);

INVx6_ASAP7_75t_L g87 ( 
.A(n_75),
.Y(n_87)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_87),
.Y(n_88)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_87),
.Y(n_89)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_89),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_83),
.A2(n_67),
.B1(n_77),
.B2(n_74),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_92),
.A2(n_63),
.B1(n_78),
.B2(n_64),
.Y(n_111)
);

BUFx3_ASAP7_75t_L g93 ( 
.A(n_83),
.Y(n_93)
);

CKINVDCx16_ASAP7_75t_R g103 ( 
.A(n_93),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_81),
.B(n_56),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_94),
.B(n_95),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_86),
.B(n_56),
.Y(n_95)
);

INVx5_ASAP7_75t_L g97 ( 
.A(n_85),
.Y(n_97)
);

HB1xp67_ASAP7_75t_L g110 ( 
.A(n_97),
.Y(n_110)
);

OR2x2_ASAP7_75t_L g100 ( 
.A(n_98),
.B(n_67),
.Y(n_100)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_93),
.Y(n_99)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_99),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_100),
.A2(n_73),
.B1(n_78),
.B2(n_68),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_94),
.A2(n_77),
.B1(n_74),
.B2(n_82),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_101),
.A2(n_105),
.B1(n_109),
.B2(n_111),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_95),
.B(n_80),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_104),
.B(n_1),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_90),
.A2(n_66),
.B1(n_52),
.B2(n_76),
.Y(n_105)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_96),
.Y(n_106)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_106),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_96),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_107),
.B(n_97),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_L g109 ( 
.A1(n_88),
.A2(n_54),
.B1(n_70),
.B2(n_63),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_100),
.A2(n_91),
.B1(n_71),
.B2(n_89),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_113),
.A2(n_119),
.B1(n_122),
.B2(n_10),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_114),
.B(n_115),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_102),
.B(n_51),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_116),
.B(n_123),
.Y(n_137)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_110),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_117),
.B(n_120),
.Y(n_139)
);

AOI21xp5_ASAP7_75t_L g118 ( 
.A1(n_101),
.A2(n_57),
.B(n_79),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_SL g131 ( 
.A1(n_118),
.A2(n_59),
.B(n_26),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_103),
.B(n_54),
.C(n_70),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_119),
.B(n_121),
.C(n_122),
.Y(n_130)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_108),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_105),
.B(n_60),
.Y(n_123)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_108),
.Y(n_124)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_124),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_109),
.B(n_62),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_125),
.B(n_127),
.Y(n_138)
);

OAI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_101),
.A2(n_88),
.B1(n_72),
.B2(n_69),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_126),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_140)
);

BUFx3_ASAP7_75t_L g128 ( 
.A(n_108),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_105),
.B(n_73),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_129),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_130),
.B(n_141),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_131),
.B(n_28),
.Y(n_144)
);

AND2x2_ASAP7_75t_L g133 ( 
.A(n_121),
.B(n_3),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_SL g146 ( 
.A1(n_133),
.A2(n_9),
.B(n_10),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_L g135 ( 
.A1(n_112),
.A2(n_3),
.B(n_4),
.Y(n_135)
);

AOI21xp5_ASAP7_75t_L g145 ( 
.A1(n_135),
.A2(n_136),
.B(n_7),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_L g136 ( 
.A1(n_126),
.A2(n_4),
.B(n_5),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_140),
.A2(n_9),
.B1(n_11),
.B2(n_20),
.Y(n_148)
);

FAx1_ASAP7_75t_SL g143 ( 
.A(n_130),
.B(n_29),
.CI(n_49),
.CON(n_143),
.SN(n_143)
);

HAxp5_ASAP7_75t_SL g155 ( 
.A(n_143),
.B(n_146),
.CON(n_155),
.SN(n_155)
);

CKINVDCx14_ASAP7_75t_R g156 ( 
.A(n_144),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_145),
.A2(n_147),
.B1(n_148),
.B2(n_151),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_138),
.A2(n_128),
.B1(n_30),
.B2(n_14),
.Y(n_147)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_139),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_150),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_134),
.B(n_33),
.Y(n_151)
);

AO21x2_ASAP7_75t_L g154 ( 
.A1(n_145),
.A2(n_136),
.B(n_133),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_154),
.A2(n_140),
.B1(n_147),
.B2(n_149),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_L g159 ( 
.A1(n_157),
.A2(n_158),
.B(n_142),
.Y(n_159)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_153),
.Y(n_158)
);

NOR3xp33_ASAP7_75t_L g160 ( 
.A(n_159),
.B(n_135),
.C(n_154),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g161 ( 
.A(n_160),
.B(n_154),
.Y(n_161)
);

HB1xp67_ASAP7_75t_L g162 ( 
.A(n_161),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_SL g163 ( 
.A(n_162),
.B(n_137),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_163),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_164),
.B(n_156),
.Y(n_165)
);

AOI321xp33_ASAP7_75t_L g166 ( 
.A1(n_165),
.A2(n_132),
.A3(n_155),
.B1(n_152),
.B2(n_143),
.C(n_148),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_166),
.B(n_34),
.C(n_23),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_167),
.B(n_36),
.C(n_25),
.Y(n_168)
);

MAJx2_ASAP7_75t_L g169 ( 
.A(n_168),
.B(n_27),
.C(n_31),
.Y(n_169)
);

AOI21xp5_ASAP7_75t_L g170 ( 
.A1(n_169),
.A2(n_39),
.B(n_48),
.Y(n_170)
);


endmodule