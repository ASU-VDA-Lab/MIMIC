module real_aes_4526_n_8 (n_4, n_0, n_3, n_5, n_2, n_7, n_6, n_1, n_8);
input n_4;
input n_0;
input n_3;
input n_5;
input n_2;
input n_7;
input n_6;
input n_1;
output n_8;
wire n_17;
wire n_22;
wire n_24;
wire n_13;
wire n_12;
wire n_19;
wire n_14;
wire n_11;
wire n_16;
wire n_15;
wire n_23;
wire n_9;
wire n_20;
wire n_18;
wire n_21;
wire n_10;
AOI21xp5_ASAP7_75t_L g8 ( .A1(n_0), .A2(n_9), .B(n_23), .Y(n_8) );
HB1xp67_ASAP7_75t_L g22 ( .A(n_1), .Y(n_22) );
OAI321xp33_ASAP7_75t_L g9 ( .A1(n_2), .A2(n_10), .A3(n_11), .B1(n_12), .B2(n_14), .C(n_21), .Y(n_9) );
HB1xp67_ASAP7_75t_L g10 ( .A(n_3), .Y(n_10) );
BUFx6f_ASAP7_75t_L g18 ( .A(n_4), .Y(n_18) );
CKINVDCx5p33_ASAP7_75t_R g20 ( .A(n_5), .Y(n_20) );
CKINVDCx5p33_ASAP7_75t_R g19 ( .A(n_6), .Y(n_19) );
INVx1_ASAP7_75t_L g13 ( .A(n_7), .Y(n_13) );
NOR2xp33_ASAP7_75t_L g23 ( .A(n_9), .B(n_24), .Y(n_23) );
NOR2xp33_ASAP7_75t_L g24 ( .A(n_11), .B(n_22), .Y(n_24) );
CKINVDCx5p33_ASAP7_75t_R g11 ( .A(n_12), .Y(n_11) );
HB1xp67_ASAP7_75t_L g12 ( .A(n_13), .Y(n_12) );
AOI22xp5_ASAP7_75t_L g14 ( .A1(n_15), .A2(n_16), .B1(n_19), .B2(n_20), .Y(n_14) );
INVx2_ASAP7_75t_SL g15 ( .A(n_16), .Y(n_15) );
BUFx2_ASAP7_75t_L g16 ( .A(n_17), .Y(n_16) );
HB1xp67_ASAP7_75t_L g17 ( .A(n_18), .Y(n_17) );
CKINVDCx20_ASAP7_75t_R g21 ( .A(n_22), .Y(n_21) );
endmodule