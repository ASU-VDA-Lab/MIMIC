module fake_ariane_340_n_199 (n_8, n_24, n_7, n_22, n_1, n_6, n_13, n_20, n_27, n_29, n_17, n_4, n_2, n_18, n_28, n_9, n_11, n_26, n_3, n_14, n_0, n_19, n_30, n_31, n_16, n_5, n_12, n_15, n_21, n_23, n_10, n_25, n_199);

input n_8;
input n_24;
input n_7;
input n_22;
input n_1;
input n_6;
input n_13;
input n_20;
input n_27;
input n_29;
input n_17;
input n_4;
input n_2;
input n_18;
input n_28;
input n_9;
input n_11;
input n_26;
input n_3;
input n_14;
input n_0;
input n_19;
input n_30;
input n_31;
input n_16;
input n_5;
input n_12;
input n_15;
input n_21;
input n_23;
input n_10;
input n_25;

output n_199;

wire n_83;
wire n_56;
wire n_60;
wire n_170;
wire n_190;
wire n_160;
wire n_64;
wire n_179;
wire n_180;
wire n_119;
wire n_124;
wire n_167;
wire n_90;
wire n_195;
wire n_38;
wire n_47;
wire n_110;
wire n_153;
wire n_197;
wire n_86;
wire n_75;
wire n_89;
wire n_67;
wire n_176;
wire n_149;
wire n_34;
wire n_158;
wire n_172;
wire n_69;
wire n_95;
wire n_175;
wire n_92;
wire n_143;
wire n_183;
wire n_150;
wire n_98;
wire n_74;
wire n_113;
wire n_114;
wire n_33;
wire n_40;
wire n_181;
wire n_152;
wire n_120;
wire n_169;
wire n_106;
wire n_53;
wire n_173;
wire n_111;
wire n_115;
wire n_133;
wire n_66;
wire n_71;
wire n_109;
wire n_96;
wire n_156;
wire n_49;
wire n_174;
wire n_100;
wire n_50;
wire n_187;
wire n_132;
wire n_62;
wire n_147;
wire n_51;
wire n_166;
wire n_76;
wire n_103;
wire n_79;
wire n_46;
wire n_84;
wire n_36;
wire n_91;
wire n_159;
wire n_107;
wire n_189;
wire n_72;
wire n_105;
wire n_128;
wire n_44;
wire n_82;
wire n_178;
wire n_42;
wire n_57;
wire n_131;
wire n_70;
wire n_117;
wire n_139;
wire n_165;
wire n_85;
wire n_144;
wire n_130;
wire n_48;
wire n_101;
wire n_94;
wire n_134;
wire n_188;
wire n_185;
wire n_32;
wire n_37;
wire n_58;
wire n_65;
wire n_123;
wire n_138;
wire n_112;
wire n_45;
wire n_162;
wire n_129;
wire n_126;
wire n_137;
wire n_122;
wire n_198;
wire n_148;
wire n_164;
wire n_52;
wire n_157;
wire n_184;
wire n_177;
wire n_135;
wire n_73;
wire n_77;
wire n_171;
wire n_121;
wire n_93;
wire n_118;
wire n_61;
wire n_108;
wire n_102;
wire n_182;
wire n_196;
wire n_125;
wire n_168;
wire n_43;
wire n_81;
wire n_87;
wire n_41;
wire n_140;
wire n_55;
wire n_191;
wire n_151;
wire n_136;
wire n_192;
wire n_80;
wire n_146;
wire n_194;
wire n_97;
wire n_154;
wire n_142;
wire n_161;
wire n_163;
wire n_88;
wire n_186;
wire n_141;
wire n_68;
wire n_116;
wire n_104;
wire n_145;
wire n_78;
wire n_193;
wire n_39;
wire n_63;
wire n_59;
wire n_99;
wire n_155;
wire n_127;
wire n_35;
wire n_54;

CKINVDCx5p33_ASAP7_75t_R g32 ( 
.A(n_9),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_17),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_20),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_25),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_23),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_13),
.Y(n_39)
);

INVxp67_ASAP7_75t_SL g40 ( 
.A(n_19),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_7),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_27),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_29),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_30),
.Y(n_44)
);

CKINVDCx5p33_ASAP7_75t_R g45 ( 
.A(n_2),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_10),
.Y(n_46)
);

CKINVDCx5p33_ASAP7_75t_R g47 ( 
.A(n_11),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_15),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_0),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_13),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_7),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_22),
.Y(n_52)
);

INVxp67_ASAP7_75t_SL g53 ( 
.A(n_14),
.Y(n_53)
);

INVxp33_ASAP7_75t_SL g54 ( 
.A(n_11),
.Y(n_54)
);

CKINVDCx5p33_ASAP7_75t_R g55 ( 
.A(n_37),
.Y(n_55)
);

CKINVDCx5p33_ASAP7_75t_R g56 ( 
.A(n_38),
.Y(n_56)
);

BUFx2_ASAP7_75t_L g57 ( 
.A(n_33),
.Y(n_57)
);

CKINVDCx5p33_ASAP7_75t_R g58 ( 
.A(n_32),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_41),
.Y(n_59)
);

CKINVDCx5p33_ASAP7_75t_R g60 ( 
.A(n_54),
.Y(n_60)
);

CKINVDCx5p33_ASAP7_75t_R g61 ( 
.A(n_45),
.Y(n_61)
);

CKINVDCx5p33_ASAP7_75t_R g62 ( 
.A(n_47),
.Y(n_62)
);

CKINVDCx5p33_ASAP7_75t_R g63 ( 
.A(n_34),
.Y(n_63)
);

CKINVDCx5p33_ASAP7_75t_R g64 ( 
.A(n_34),
.Y(n_64)
);

CKINVDCx5p33_ASAP7_75t_R g65 ( 
.A(n_35),
.Y(n_65)
);

CKINVDCx5p33_ASAP7_75t_R g66 ( 
.A(n_35),
.Y(n_66)
);

CKINVDCx5p33_ASAP7_75t_R g67 ( 
.A(n_44),
.Y(n_67)
);

CKINVDCx5p33_ASAP7_75t_R g68 ( 
.A(n_42),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_33),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_36),
.Y(n_70)
);

CKINVDCx5p33_ASAP7_75t_R g71 ( 
.A(n_42),
.Y(n_71)
);

CKINVDCx5p33_ASAP7_75t_R g72 ( 
.A(n_43),
.Y(n_72)
);

CKINVDCx5p33_ASAP7_75t_R g73 ( 
.A(n_43),
.Y(n_73)
);

CKINVDCx5p33_ASAP7_75t_R g74 ( 
.A(n_52),
.Y(n_74)
);

CKINVDCx5p33_ASAP7_75t_R g75 ( 
.A(n_53),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_57),
.Y(n_76)
);

HB1xp67_ASAP7_75t_L g77 ( 
.A(n_61),
.Y(n_77)
);

AO22x2_ASAP7_75t_L g78 ( 
.A1(n_69),
.A2(n_51),
.B1(n_50),
.B2(n_49),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_57),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_69),
.A2(n_51),
.B1(n_50),
.B2(n_49),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_63),
.B(n_40),
.Y(n_81)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_64),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_65),
.B(n_68),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_74),
.B(n_46),
.Y(n_84)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_67),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_66),
.Y(n_86)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_67),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_71),
.B(n_48),
.Y(n_88)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_72),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_73),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_62),
.B(n_48),
.Y(n_91)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_75),
.Y(n_92)
);

A2O1A1Ixp33_ASAP7_75t_L g93 ( 
.A1(n_85),
.A2(n_39),
.B(n_36),
.C(n_58),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_92),
.B(n_58),
.Y(n_94)
);

NOR3xp33_ASAP7_75t_SL g95 ( 
.A(n_80),
.B(n_60),
.C(n_39),
.Y(n_95)
);

A2O1A1Ixp33_ASAP7_75t_L g96 ( 
.A1(n_85),
.A2(n_70),
.B(n_56),
.C(n_55),
.Y(n_96)
);

OR2x6_ASAP7_75t_L g97 ( 
.A(n_78),
.B(n_80),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_84),
.Y(n_98)
);

INVx3_ASAP7_75t_SL g99 ( 
.A(n_92),
.Y(n_99)
);

AOI21xp5_ASAP7_75t_L g100 ( 
.A1(n_81),
.A2(n_31),
.B(n_28),
.Y(n_100)
);

INVx1_ASAP7_75t_SL g101 ( 
.A(n_83),
.Y(n_101)
);

NOR2x1_ASAP7_75t_L g102 ( 
.A(n_92),
.B(n_70),
.Y(n_102)
);

AOI21xp5_ASAP7_75t_L g103 ( 
.A1(n_81),
.A2(n_26),
.B(n_24),
.Y(n_103)
);

BUFx4f_ASAP7_75t_L g104 ( 
.A(n_82),
.Y(n_104)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_98),
.Y(n_105)
);

OAI21x1_ASAP7_75t_L g106 ( 
.A1(n_100),
.A2(n_85),
.B(n_87),
.Y(n_106)
);

BUFx8_ASAP7_75t_L g107 ( 
.A(n_101),
.Y(n_107)
);

OAI21x1_ASAP7_75t_L g108 ( 
.A1(n_103),
.A2(n_87),
.B(n_88),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_93),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_104),
.A2(n_87),
.B1(n_89),
.B2(n_90),
.Y(n_110)
);

AOI21xp5_ASAP7_75t_L g111 ( 
.A1(n_104),
.A2(n_89),
.B(n_90),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_101),
.Y(n_112)
);

AO31x2_ASAP7_75t_L g113 ( 
.A1(n_109),
.A2(n_96),
.A3(n_89),
.B(n_82),
.Y(n_113)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_105),
.Y(n_114)
);

OR2x2_ASAP7_75t_L g115 ( 
.A(n_112),
.B(n_97),
.Y(n_115)
);

AND2x4_ASAP7_75t_L g116 ( 
.A(n_105),
.B(n_111),
.Y(n_116)
);

NAND2xp33_ASAP7_75t_R g117 ( 
.A(n_107),
.B(n_83),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_R g118 ( 
.A(n_107),
.B(n_59),
.Y(n_118)
);

AND2x2_ASAP7_75t_L g119 ( 
.A(n_110),
.B(n_97),
.Y(n_119)
);

INVx2_ASAP7_75t_SL g120 ( 
.A(n_116),
.Y(n_120)
);

HB1xp67_ASAP7_75t_L g121 ( 
.A(n_116),
.Y(n_121)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_114),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g123 ( 
.A(n_119),
.B(n_97),
.Y(n_123)
);

OA21x2_ASAP7_75t_L g124 ( 
.A1(n_116),
.A2(n_106),
.B(n_108),
.Y(n_124)
);

INVxp67_ASAP7_75t_SL g125 ( 
.A(n_121),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_122),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_122),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_121),
.B(n_114),
.Y(n_128)
);

OR2x2_ASAP7_75t_L g129 ( 
.A(n_121),
.B(n_115),
.Y(n_129)
);

AND2x2_ASAP7_75t_L g130 ( 
.A(n_123),
.B(n_119),
.Y(n_130)
);

OR2x2_ASAP7_75t_L g131 ( 
.A(n_120),
.B(n_115),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_123),
.B(n_59),
.Y(n_132)
);

AND2x4_ASAP7_75t_L g133 ( 
.A(n_120),
.B(n_116),
.Y(n_133)
);

HB1xp67_ASAP7_75t_L g134 ( 
.A(n_120),
.Y(n_134)
);

AND2x2_ASAP7_75t_L g135 ( 
.A(n_123),
.B(n_113),
.Y(n_135)
);

OR2x2_ASAP7_75t_L g136 ( 
.A(n_129),
.B(n_123),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g137 ( 
.A(n_132),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_126),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_133),
.A2(n_117),
.B1(n_107),
.B2(n_102),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_133),
.B(n_120),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_126),
.Y(n_141)
);

BUFx2_ASAP7_75t_L g142 ( 
.A(n_125),
.Y(n_142)
);

AOI33xp33_ASAP7_75t_L g143 ( 
.A1(n_127),
.A2(n_91),
.A3(n_86),
.B1(n_79),
.B2(n_76),
.B3(n_95),
.Y(n_143)
);

NAND2x1_ASAP7_75t_L g144 ( 
.A(n_142),
.B(n_127),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_136),
.B(n_128),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_138),
.B(n_128),
.Y(n_146)
);

INVx1_ASAP7_75t_SL g147 ( 
.A(n_139),
.Y(n_147)
);

AOI21xp33_ASAP7_75t_SL g148 ( 
.A1(n_137),
.A2(n_77),
.B(n_86),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_141),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_140),
.B(n_125),
.Y(n_150)
);

NAND2x1_ASAP7_75t_L g151 ( 
.A(n_140),
.B(n_133),
.Y(n_151)
);

OAI32xp33_ASAP7_75t_L g152 ( 
.A1(n_143),
.A2(n_92),
.A3(n_94),
.B1(n_91),
.B2(n_134),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_149),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_146),
.Y(n_154)
);

INVx3_ASAP7_75t_L g155 ( 
.A(n_144),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_145),
.B(n_134),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_150),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_148),
.A2(n_78),
.B1(n_129),
.B2(n_120),
.Y(n_158)
);

OAI221xp5_ASAP7_75t_L g159 ( 
.A1(n_147),
.A2(n_76),
.B1(n_79),
.B2(n_131),
.C(n_78),
.Y(n_159)
);

HB1xp67_ASAP7_75t_L g160 ( 
.A(n_150),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_152),
.B(n_151),
.Y(n_161)
);

INVx6_ASAP7_75t_L g162 ( 
.A(n_144),
.Y(n_162)
);

O2A1O1Ixp33_ASAP7_75t_L g163 ( 
.A1(n_158),
.A2(n_99),
.B(n_78),
.C(n_143),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_161),
.A2(n_78),
.B1(n_135),
.B2(n_130),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_157),
.B(n_135),
.Y(n_165)
);

NOR5xp2_ASAP7_75t_L g166 ( 
.A(n_160),
.B(n_122),
.C(n_113),
.D(n_118),
.E(n_3),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_L g167 ( 
.A1(n_159),
.A2(n_123),
.B1(n_130),
.B2(n_131),
.Y(n_167)
);

AOI21xp5_ASAP7_75t_L g168 ( 
.A1(n_161),
.A2(n_160),
.B(n_133),
.Y(n_168)
);

NOR4xp25_ASAP7_75t_L g169 ( 
.A(n_154),
.B(n_122),
.C(n_113),
.D(n_2),
.Y(n_169)
);

A2O1A1Ixp33_ASAP7_75t_L g170 ( 
.A1(n_153),
.A2(n_108),
.B(n_113),
.C(n_106),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_156),
.Y(n_171)
);

AND2x2_ASAP7_75t_L g172 ( 
.A(n_171),
.B(n_155),
.Y(n_172)
);

INVx2_ASAP7_75t_SL g173 ( 
.A(n_165),
.Y(n_173)
);

NAND3xp33_ASAP7_75t_SL g174 ( 
.A(n_168),
.B(n_162),
.C(n_155),
.Y(n_174)
);

NOR4xp75_ASAP7_75t_L g175 ( 
.A(n_169),
.B(n_162),
.C(n_1),
.D(n_3),
.Y(n_175)
);

NOR2x1_ASAP7_75t_L g176 ( 
.A(n_170),
.B(n_162),
.Y(n_176)
);

AND2x2_ASAP7_75t_L g177 ( 
.A(n_164),
.B(n_124),
.Y(n_177)
);

OAI211xp5_ASAP7_75t_L g178 ( 
.A1(n_163),
.A2(n_0),
.B(n_1),
.C(n_4),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_167),
.A2(n_113),
.B1(n_124),
.B2(n_6),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_L g180 ( 
.A1(n_176),
.A2(n_167),
.B(n_166),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_172),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_178),
.A2(n_177),
.B1(n_179),
.B2(n_174),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_173),
.Y(n_183)
);

AOI22xp33_ASAP7_75t_L g184 ( 
.A1(n_179),
.A2(n_175),
.B1(n_124),
.B2(n_6),
.Y(n_184)
);

INVx1_ASAP7_75t_SL g185 ( 
.A(n_172),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_183),
.Y(n_186)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_185),
.Y(n_187)
);

NOR2x1p5_ASAP7_75t_L g188 ( 
.A(n_181),
.B(n_4),
.Y(n_188)
);

NAND4xp25_ASAP7_75t_L g189 ( 
.A(n_184),
.B(n_5),
.C(n_8),
.D(n_9),
.Y(n_189)
);

INVx1_ASAP7_75t_SL g190 ( 
.A(n_181),
.Y(n_190)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_190),
.Y(n_191)
);

OAI22x1_ASAP7_75t_L g192 ( 
.A1(n_188),
.A2(n_182),
.B1(n_187),
.B2(n_186),
.Y(n_192)
);

OAI22x1_ASAP7_75t_L g193 ( 
.A1(n_187),
.A2(n_180),
.B1(n_124),
.B2(n_10),
.Y(n_193)
);

AOI221xp5_ASAP7_75t_L g194 ( 
.A1(n_189),
.A2(n_5),
.B1(n_8),
.B2(n_12),
.C(n_14),
.Y(n_194)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_191),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_192),
.B(n_12),
.Y(n_196)
);

OAI211xp5_ASAP7_75t_L g197 ( 
.A1(n_194),
.A2(n_16),
.B(n_124),
.C(n_21),
.Y(n_197)
);

AOI22xp33_ASAP7_75t_SL g198 ( 
.A1(n_197),
.A2(n_193),
.B1(n_124),
.B2(n_18),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_198),
.A2(n_196),
.B1(n_195),
.B2(n_124),
.Y(n_199)
);


endmodule