module fake_netlist_1_6388_n_939 (n_107, n_103, n_52, n_50, n_7, n_3, n_34, n_25, n_9, n_96, n_72, n_77, n_90, n_99, n_43, n_73, n_62, n_97, n_33, n_4, n_59, n_76, n_6, n_74, n_8, n_61, n_44, n_66, n_88, n_46, n_108, n_37, n_18, n_65, n_87, n_5, n_81, n_85, n_102, n_47, n_1, n_16, n_78, n_95, n_40, n_68, n_105, n_36, n_11, n_15, n_71, n_70, n_94, n_2, n_17, n_58, n_20, n_84, n_12, n_56, n_80, n_67, n_22, n_19, n_26, n_39, n_101, n_98, n_38, n_104, n_100, n_24, n_35, n_91, n_32, n_93, n_48, n_63, n_54, n_41, n_55, n_29, n_60, n_10, n_30, n_13, n_92, n_75, n_82, n_53, n_64, n_69, n_83, n_23, n_0, n_57, n_51, n_106, n_45, n_42, n_21, n_86, n_27, n_89, n_28, n_79, n_49, n_14, n_31, n_939, n_940);
input n_107;
input n_103;
input n_52;
input n_50;
input n_7;
input n_3;
input n_34;
input n_25;
input n_9;
input n_96;
input n_72;
input n_77;
input n_90;
input n_99;
input n_43;
input n_73;
input n_62;
input n_97;
input n_33;
input n_4;
input n_59;
input n_76;
input n_6;
input n_74;
input n_8;
input n_61;
input n_44;
input n_66;
input n_88;
input n_46;
input n_108;
input n_37;
input n_18;
input n_65;
input n_87;
input n_5;
input n_81;
input n_85;
input n_102;
input n_47;
input n_1;
input n_16;
input n_78;
input n_95;
input n_40;
input n_68;
input n_105;
input n_36;
input n_11;
input n_15;
input n_71;
input n_70;
input n_94;
input n_2;
input n_17;
input n_58;
input n_20;
input n_84;
input n_12;
input n_56;
input n_80;
input n_67;
input n_22;
input n_19;
input n_26;
input n_39;
input n_101;
input n_98;
input n_38;
input n_104;
input n_100;
input n_24;
input n_35;
input n_91;
input n_32;
input n_93;
input n_48;
input n_63;
input n_54;
input n_41;
input n_55;
input n_29;
input n_60;
input n_10;
input n_30;
input n_13;
input n_92;
input n_75;
input n_82;
input n_53;
input n_64;
input n_69;
input n_83;
input n_23;
input n_0;
input n_57;
input n_51;
input n_106;
input n_45;
input n_42;
input n_21;
input n_86;
input n_27;
input n_89;
input n_28;
input n_79;
input n_49;
input n_14;
input n_31;
output n_939;
output n_940;
wire n_890;
wire n_107;
wire n_646;
wire n_759;
wire n_658;
wire n_673;
wire n_156;
wire n_154;
wire n_239;
wire n_7;
wire n_309;
wire n_356;
wire n_895;
wire n_327;
wire n_25;
wire n_204;
wire n_592;
wire n_769;
wire n_929;
wire n_169;
wire n_370;
wire n_384;
wire n_439;
wire n_545;
wire n_180;
wire n_604;
wire n_99;
wire n_43;
wire n_73;
wire n_440;
wire n_199;
wire n_279;
wire n_786;
wire n_831;
wire n_357;
wire n_74;
wire n_729;
wire n_308;
wire n_518;
wire n_394;
wire n_44;
wire n_189;
wire n_681;
wire n_226;
wire n_352;
wire n_447;
wire n_66;
wire n_379;
wire n_903;
wire n_535;
wire n_689;
wire n_886;
wire n_595;
wire n_875;
wire n_626;
wire n_316;
wire n_285;
wire n_564;
wire n_586;
wire n_471;
wire n_47;
wire n_766;
wire n_475;
wire n_744;
wire n_850;
wire n_281;
wire n_645;
wire n_497;
wire n_399;
wire n_11;
wire n_295;
wire n_371;
wire n_579;
wire n_516;
wire n_608;
wire n_368;
wire n_805;
wire n_373;
wire n_139;
wire n_342;
wire n_151;
wire n_71;
wire n_288;
wire n_557;
wire n_176;
wire n_753;
wire n_859;
wire n_436;
wire n_438;
wire n_900;
wire n_869;
wire n_931;
wire n_935;
wire n_359;
wire n_195;
wire n_300;
wire n_487;
wire n_461;
wire n_723;
wire n_223;
wire n_833;
wire n_405;
wire n_830;
wire n_562;
wire n_19;
wire n_409;
wire n_482;
wire n_838;
wire n_569;
wire n_534;
wire n_707;
wire n_526;
wire n_261;
wire n_423;
wire n_483;
wire n_220;
wire n_353;
wire n_410;
wire n_104;
wire n_709;
wire n_303;
wire n_502;
wire n_821;
wire n_468;
wire n_159;
wire n_566;
wire n_91;
wire n_301;
wire n_340;
wire n_148;
wire n_149;
wire n_567;
wire n_378;
wire n_752;
wire n_246;
wire n_676;
wire n_823;
wire n_191;
wire n_143;
wire n_780;
wire n_864;
wire n_629;
wire n_446;
wire n_63;
wire n_402;
wire n_54;
wire n_876;
wire n_387;
wire n_125;
wire n_145;
wire n_166;
wire n_558;
wire n_596;
wire n_492;
wire n_181;
wire n_123;
wire n_219;
wire n_343;
wire n_494;
wire n_553;
wire n_555;
wire n_135;
wire n_481;
wire n_621;
wire n_817;
wire n_776;
wire n_315;
wire n_397;
wire n_53;
wire n_880;
wire n_213;
wire n_196;
wire n_293;
wire n_797;
wire n_836;
wire n_127;
wire n_312;
wire n_742;
wire n_424;
wire n_23;
wire n_110;
wire n_182;
wire n_269;
wire n_663;
wire n_529;
wire n_656;
wire n_751;
wire n_887;
wire n_186;
wire n_137;
wire n_507;
wire n_334;
wire n_164;
wire n_433;
wire n_660;
wire n_120;
wire n_392;
wire n_650;
wire n_806;
wire n_155;
wire n_162;
wire n_114;
wire n_772;
wire n_50;
wire n_816;
wire n_789;
wire n_3;
wire n_331;
wire n_651;
wire n_574;
wire n_882;
wire n_636;
wire n_330;
wire n_614;
wire n_231;
wire n_884;
wire n_9;
wire n_737;
wire n_428;
wire n_178;
wire n_478;
wire n_814;
wire n_652;
wire n_678;
wire n_708;
wire n_229;
wire n_97;
wire n_133;
wire n_324;
wire n_442;
wire n_422;
wire n_192;
wire n_699;
wire n_857;
wire n_329;
wire n_6;
wire n_8;
wire n_578;
wire n_928;
wire n_883;
wire n_187;
wire n_548;
wire n_188;
wire n_443;
wire n_304;
wire n_18;
wire n_682;
wire n_801;
wire n_441;
wire n_868;
wire n_628;
wire n_425;
wire n_920;
wire n_912;
wire n_314;
wire n_824;
wire n_601;
wire n_307;
wire n_517;
wire n_215;
wire n_736;
wire n_172;
wire n_905;
wire n_109;
wire n_332;
wire n_198;
wire n_386;
wire n_934;
wire n_653;
wire n_351;
wire n_1;
wire n_16;
wire n_670;
wire n_95;
wire n_40;
wire n_210;
wire n_426;
wire n_755;
wire n_716;
wire n_228;
wire n_863;
wire n_671;
wire n_892;
wire n_278;
wire n_115;
wire n_270;
wire n_476;
wire n_765;
wire n_829;
wire n_599;
wire n_715;
wire n_849;
wire n_179;
wire n_289;
wire n_404;
wire n_366;
wire n_721;
wire n_362;
wire n_617;
wire n_688;
wire n_837;
wire n_485;
wire n_396;
wire n_549;
wire n_354;
wire n_720;
wire n_152;
wire n_851;
wire n_70;
wire n_588;
wire n_458;
wire n_375;
wire n_855;
wire n_17;
wire n_322;
wire n_911;
wire n_317;
wire n_221;
wire n_328;
wire n_506;
wire n_711;
wire n_491;
wire n_800;
wire n_388;
wire n_773;
wire n_266;
wire n_763;
wire n_80;
wire n_632;
wire n_793;
wire n_906;
wire n_679;
wire n_522;
wire n_546;
wire n_615;
wire n_684;
wire n_701;
wire n_326;
wire n_532;
wire n_756;
wire n_635;
wire n_544;
wire n_879;
wire n_888;
wire n_576;
wire n_275;
wire n_691;
wire n_622;
wire n_661;
wire n_909;
wire n_493;
wire n_274;
wire n_910;
wire n_150;
wire n_235;
wire n_690;
wire n_38;
wire n_533;
wire n_272;
wire n_686;
wire n_299;
wire n_100;
wire n_561;
wire n_581;
wire n_280;
wire n_141;
wire n_509;
wire n_160;
wire n_499;
wire n_377;
wire n_263;
wire n_757;
wire n_844;
wire n_695;
wire n_193;
wire n_232;
wire n_344;
wire n_878;
wire n_783;
wire n_812;
wire n_147;
wire n_185;
wire n_367;
wire n_795;
wire n_267;
wire n_687;
wire n_171;
wire n_638;
wire n_873;
wire n_899;
wire n_450;
wire n_585;
wire n_140;
wire n_644;
wire n_111;
wire n_746;
wire n_212;
wire n_779;
wire n_30;
wire n_634;
wire n_13;
wire n_254;
wire n_559;
wire n_704;
wire n_435;
wire n_728;
wire n_583;
wire n_841;
wire n_64;
wire n_69;
wire n_248;
wire n_866;
wire n_407;
wire n_527;
wire n_83;
wire n_200;
wire n_603;
wire n_262;
wire n_921;
wire n_119;
wire n_667;
wire n_503;
wire n_856;
wire n_927;
wire n_339;
wire n_347;
wire n_124;
wire n_696;
wire n_748;
wire n_79;
wire n_129;
wire n_904;
wire n_611;
wire n_521;
wire n_157;
wire n_774;
wire n_103;
wire n_808;
wire n_421;
wire n_52;
wire n_253;
wire n_434;
wire n_677;
wire n_624;
wire n_273;
wire n_325;
wire n_571;
wire n_524;
wire n_692;
wire n_530;
wire n_743;
wire n_163;
wire n_348;
wire n_96;
wire n_685;
wire n_762;
wire n_77;
wire n_72;
wire n_90;
wire n_594;
wire n_669;
wire n_214;
wire n_787;
wire n_770;
wire n_167;
wire n_861;
wire n_809;
wire n_364;
wire n_33;
wire n_908;
wire n_464;
wire n_76;
wire n_470;
wire n_590;
wire n_61;
wire n_463;
wire n_216;
wire n_153;
wire n_355;
wire n_609;
wire n_121;
wire n_286;
wire n_408;
wire n_247;
wire n_431;
wire n_224;
wire n_161;
wire n_484;
wire n_165;
wire n_860;
wire n_413;
wire n_65;
wire n_537;
wire n_710;
wire n_525;
wire n_560;
wire n_5;
wire n_496;
wire n_393;
wire n_843;
wire n_211;
wire n_85;
wire n_320;
wire n_264;
wire n_102;
wire n_283;
wire n_733;
wire n_846;
wire n_290;
wire n_217;
wire n_201;
wire n_791;
wire n_792;
wire n_277;
wire n_932;
wire n_259;
wire n_885;
wire n_612;
wire n_244;
wire n_666;
wire n_771;
wire n_827;
wire n_276;
wire n_297;
wire n_225;
wire n_631;
wire n_350;
wire n_747;
wire n_208;
wire n_616;
wire n_854;
wire n_523;
wire n_815;
wire n_901;
wire n_528;
wire n_419;
wire n_252;
wire n_922;
wire n_519;
wire n_168;
wire n_839;
wire n_271;
wire n_693;
wire n_785;
wire n_896;
wire n_739;
wire n_94;
wire n_194;
wire n_858;
wire n_758;
wire n_825;
wire n_282;
wire n_58;
wire n_775;
wire n_113;
wire n_242;
wire n_498;
wire n_501;
wire n_284;
wire n_321;
wire n_302;
wire n_538;
wire n_703;
wire n_811;
wire n_116;
wire n_734;
wire n_292;
wire n_547;
wire n_593;
wire n_118;
wire n_587;
wire n_233;
wire n_554;
wire n_597;
wire n_698;
wire n_741;
wire n_257;
wire n_705;
wire n_828;
wire n_722;
wire n_203;
wire n_26;
wire n_477;
wire n_460;
wire n_243;
wire n_318;
wire n_346;
wire n_98;
wire n_345;
wire n_230;
wire n_452;
wire n_714;
wire n_146;
wire n_337;
wire n_32;
wire n_637;
wire n_641;
wire n_726;
wire n_531;
wire n_872;
wire n_93;
wire n_539;
wire n_847;
wire n_406;
wire n_372;
wire n_842;
wire n_820;
wire n_713;
wire n_467;
wire n_923;
wire n_702;
wire n_41;
wire n_760;
wire n_826;
wire n_918;
wire n_623;
wire n_417;
wire n_451;
wire n_665;
wire n_898;
wire n_647;
wire n_445;
wire n_500;
wire n_732;
wire n_926;
wire n_845;
wire n_575;
wire n_10;
wire n_390;
wire n_600;
wire n_818;
wire n_75;
wire n_82;
wire n_183;
wire n_731;
wire n_550;
wire n_132;
wire n_643;
wire n_761;
wire n_778;
wire n_582;
wire n_784;
wire n_170;
wire n_925;
wire n_205;
wire n_158;
wire n_915;
wire n_126;
wire n_473;
wire n_249;
wire n_389;
wire n_834;
wire n_510;
wire n_360;
wire n_363;
wire n_749;
wire n_427;
wire n_724;
wire n_106;
wire n_296;
wire n_605;
wire n_42;
wire n_21;
wire n_835;
wire n_437;
wire n_871;
wire n_620;
wire n_89;
wire n_480;
wire n_939;
wire n_130;
wire n_310;
wire n_341;
wire n_700;
wire n_640;
wire n_14;
wire n_236;
wire n_639;
wire n_727;
wire n_136;
wire n_260;
wire n_891;
wire n_580;
wire n_610;
wire n_222;
wire n_657;
wire n_822;
wire n_381;
wire n_142;
wire n_34;
wire n_853;
wire n_754;
wire n_385;
wire n_798;
wire n_227;
wire n_395;
wire n_454;
wire n_453;
wire n_250;
wire n_551;
wire n_268;
wire n_190;
wire n_606;
wire n_62;
wire n_712;
wire n_777;
wire n_4;
wire n_59;
wire n_323;
wire n_565;
wire n_781;
wire n_914;
wire n_852;
wire n_376;
wire n_902;
wire n_694;
wire n_240;
wire n_459;
wire n_768;
wire n_88;
wire n_568;
wire n_46;
wire n_174;
wire n_717;
wire n_807;
wire n_108;
wire n_335;
wire n_37;
wire n_122;
wire n_374;
wire n_613;
wire n_380;
wire n_515;
wire n_802;
wire n_865;
wire n_672;
wire n_867;
wire n_466;
wire n_87;
wire n_207;
wire n_197;
wire n_81;
wire n_572;
wire n_541;
wire n_298;
wire n_112;
wire n_630;
wire n_735;
wire n_649;
wire n_602;
wire n_78;
wire n_552;
wire n_68;
wire n_919;
wire n_444;
wire n_105;
wire n_251;
wire n_598;
wire n_810;
wire n_36;
wire n_416;
wire n_916;
wire n_870;
wire n_889;
wire n_432;
wire n_913;
wire n_917;
wire n_465;
wire n_414;
wire n_680;
wire n_730;
wire n_369;
wire n_469;
wire n_361;
wire n_767;
wire n_237;
wire n_881;
wire n_654;
wire n_15;
wire n_520;
wire n_633;
wire n_429;
wire n_803;
wire n_256;
wire n_398;
wire n_668;
wire n_117;
wire n_238;
wire n_365;
wire n_577;
wire n_796;
wire n_804;
wire n_294;
wire n_2;
wire n_338;
wire n_662;
wire n_907;
wire n_591;
wire n_391;
wire n_209;
wire n_241;
wire n_874;
wire n_84;
wire n_20;
wire n_782;
wire n_449;
wire n_832;
wire n_12;
wire n_56;
wire n_412;
wire n_455;
wire n_67;
wire n_504;
wire n_618;
wire n_790;
wire n_456;
wire n_22;
wire n_683;
wire n_479;
wire n_584;
wire n_311;
wire n_401;
wire n_877;
wire n_383;
wire n_813;
wire n_202;
wire n_319;
wire n_542;
wire n_725;
wire n_819;
wire n_862;
wire n_930;
wire n_39;
wire n_101;
wire n_291;
wire n_489;
wire n_245;
wire n_664;
wire n_933;
wire n_508;
wire n_764;
wire n_719;
wire n_486;
wire n_788;
wire n_24;
wire n_35;
wire n_655;
wire n_472;
wire n_490;
wire n_540;
wire n_840;
wire n_400;
wire n_794;
wire n_457;
wire n_659;
wire n_134;
wire n_48;
wire n_255;
wire n_563;
wire n_513;
wire n_55;
wire n_718;
wire n_543;
wire n_336;
wire n_29;
wire n_218;
wire n_893;
wire n_173;
wire n_488;
wire n_556;
wire n_648;
wire n_382;
wire n_799;
wire n_894;
wire n_138;
wire n_60;
wire n_936;
wire n_937;
wire n_462;
wire n_573;
wire n_536;
wire n_474;
wire n_924;
wire n_745;
wire n_305;
wire n_495;
wire n_505;
wire n_430;
wire n_418;
wire n_92;
wire n_313;
wire n_358;
wire n_333;
wire n_627;
wire n_740;
wire n_706;
wire n_589;
wire n_750;
wire n_175;
wire n_897;
wire n_128;
wire n_306;
wire n_31;
wire n_415;
wire n_697;
wire n_0;
wire n_512;
wire n_258;
wire n_619;
wire n_642;
wire n_675;
wire n_234;
wire n_607;
wire n_848;
wire n_184;
wire n_265;
wire n_57;
wire n_674;
wire n_51;
wire n_570;
wire n_411;
wire n_514;
wire n_287;
wire n_144;
wire n_403;
wire n_625;
wire n_45;
wire n_131;
wire n_420;
wire n_86;
wire n_27;
wire n_738;
wire n_177;
wire n_28;
wire n_511;
wire n_448;
wire n_49;
wire n_206;
wire n_349;
INVx2_ASAP7_75t_L g109 ( .A(n_23), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_46), .Y(n_110) );
CKINVDCx5p33_ASAP7_75t_R g111 ( .A(n_62), .Y(n_111) );
CKINVDCx5p33_ASAP7_75t_R g112 ( .A(n_92), .Y(n_112) );
NOR2xp67_ASAP7_75t_L g113 ( .A(n_22), .B(n_29), .Y(n_113) );
CKINVDCx20_ASAP7_75t_R g114 ( .A(n_49), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_18), .Y(n_115) );
CKINVDCx5p33_ASAP7_75t_R g116 ( .A(n_36), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_93), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_81), .Y(n_118) );
CKINVDCx5p33_ASAP7_75t_R g119 ( .A(n_94), .Y(n_119) );
INVx2_ASAP7_75t_L g120 ( .A(n_77), .Y(n_120) );
CKINVDCx5p33_ASAP7_75t_R g121 ( .A(n_7), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_84), .Y(n_122) );
CKINVDCx20_ASAP7_75t_R g123 ( .A(n_98), .Y(n_123) );
INVx1_ASAP7_75t_SL g124 ( .A(n_0), .Y(n_124) );
CKINVDCx5p33_ASAP7_75t_R g125 ( .A(n_48), .Y(n_125) );
HB1xp67_ASAP7_75t_L g126 ( .A(n_24), .Y(n_126) );
INVx1_ASAP7_75t_L g127 ( .A(n_76), .Y(n_127) );
CKINVDCx5p33_ASAP7_75t_R g128 ( .A(n_68), .Y(n_128) );
INVx1_ASAP7_75t_L g129 ( .A(n_55), .Y(n_129) );
INVx1_ASAP7_75t_L g130 ( .A(n_97), .Y(n_130) );
INVx1_ASAP7_75t_L g131 ( .A(n_2), .Y(n_131) );
CKINVDCx5p33_ASAP7_75t_R g132 ( .A(n_12), .Y(n_132) );
INVx3_ASAP7_75t_L g133 ( .A(n_101), .Y(n_133) );
CKINVDCx5p33_ASAP7_75t_R g134 ( .A(n_71), .Y(n_134) );
INVx1_ASAP7_75t_L g135 ( .A(n_83), .Y(n_135) );
INVx1_ASAP7_75t_L g136 ( .A(n_64), .Y(n_136) );
CKINVDCx20_ASAP7_75t_R g137 ( .A(n_91), .Y(n_137) );
CKINVDCx5p33_ASAP7_75t_R g138 ( .A(n_58), .Y(n_138) );
INVx1_ASAP7_75t_L g139 ( .A(n_65), .Y(n_139) );
INVx1_ASAP7_75t_L g140 ( .A(n_57), .Y(n_140) );
CKINVDCx5p33_ASAP7_75t_R g141 ( .A(n_88), .Y(n_141) );
CKINVDCx5p33_ASAP7_75t_R g142 ( .A(n_8), .Y(n_142) );
CKINVDCx5p33_ASAP7_75t_R g143 ( .A(n_69), .Y(n_143) );
CKINVDCx11_ASAP7_75t_R g144 ( .A(n_61), .Y(n_144) );
INVx1_ASAP7_75t_L g145 ( .A(n_21), .Y(n_145) );
INVx1_ASAP7_75t_L g146 ( .A(n_25), .Y(n_146) );
BUFx10_ASAP7_75t_L g147 ( .A(n_19), .Y(n_147) );
CKINVDCx20_ASAP7_75t_R g148 ( .A(n_11), .Y(n_148) );
INVx2_ASAP7_75t_L g149 ( .A(n_20), .Y(n_149) );
AND2x2_ASAP7_75t_L g150 ( .A(n_126), .B(n_0), .Y(n_150) );
INVx2_ASAP7_75t_L g151 ( .A(n_133), .Y(n_151) );
INVx5_ASAP7_75t_L g152 ( .A(n_133), .Y(n_152) );
AND2x4_ASAP7_75t_L g153 ( .A(n_133), .B(n_1), .Y(n_153) );
OAI22x1_ASAP7_75t_R g154 ( .A1(n_148), .A2(n_1), .B1(n_2), .B2(n_3), .Y(n_154) );
CKINVDCx6p67_ASAP7_75t_R g155 ( .A(n_147), .Y(n_155) );
OA21x2_ASAP7_75t_L g156 ( .A1(n_109), .A2(n_51), .B(n_107), .Y(n_156) );
INVx3_ASAP7_75t_L g157 ( .A(n_147), .Y(n_157) );
BUFx6f_ASAP7_75t_L g158 ( .A(n_109), .Y(n_158) );
INVx2_ASAP7_75t_L g159 ( .A(n_120), .Y(n_159) );
INVx1_ASAP7_75t_L g160 ( .A(n_110), .Y(n_160) );
OA21x2_ASAP7_75t_L g161 ( .A1(n_120), .A2(n_50), .B(n_106), .Y(n_161) );
INVx1_ASAP7_75t_L g162 ( .A(n_115), .Y(n_162) );
AOI22xp5_ASAP7_75t_L g163 ( .A1(n_148), .A2(n_3), .B1(n_4), .B2(n_5), .Y(n_163) );
INVx1_ASAP7_75t_L g164 ( .A(n_117), .Y(n_164) );
NAND2xp5_ASAP7_75t_SL g165 ( .A(n_147), .B(n_4), .Y(n_165) );
INVx5_ASAP7_75t_L g166 ( .A(n_149), .Y(n_166) );
AND2x2_ASAP7_75t_L g167 ( .A(n_131), .B(n_5), .Y(n_167) );
BUFx8_ASAP7_75t_L g168 ( .A(n_149), .Y(n_168) );
HB1xp67_ASAP7_75t_L g169 ( .A(n_121), .Y(n_169) );
CKINVDCx5p33_ASAP7_75t_R g170 ( .A(n_144), .Y(n_170) );
BUFx6f_ASAP7_75t_L g171 ( .A(n_118), .Y(n_171) );
INVx4_ASAP7_75t_L g172 ( .A(n_112), .Y(n_172) );
NOR2xp33_ASAP7_75t_L g173 ( .A(n_122), .B(n_6), .Y(n_173) );
AND2x4_ASAP7_75t_L g174 ( .A(n_127), .B(n_6), .Y(n_174) );
BUFx10_ASAP7_75t_L g175 ( .A(n_153), .Y(n_175) );
NAND2xp5_ASAP7_75t_SL g176 ( .A(n_172), .B(n_112), .Y(n_176) );
INVx2_ASAP7_75t_L g177 ( .A(n_158), .Y(n_177) );
INVx2_ASAP7_75t_L g178 ( .A(n_158), .Y(n_178) );
INVx3_ASAP7_75t_L g179 ( .A(n_153), .Y(n_179) );
NOR2xp33_ASAP7_75t_L g180 ( .A(n_157), .B(n_129), .Y(n_180) );
INVx2_ASAP7_75t_SL g181 ( .A(n_168), .Y(n_181) );
INVx2_ASAP7_75t_L g182 ( .A(n_158), .Y(n_182) );
INVx2_ASAP7_75t_L g183 ( .A(n_158), .Y(n_183) );
INVx2_ASAP7_75t_SL g184 ( .A(n_168), .Y(n_184) );
AND2x2_ASAP7_75t_L g185 ( .A(n_155), .B(n_116), .Y(n_185) );
INVx1_ASAP7_75t_L g186 ( .A(n_151), .Y(n_186) );
INVx1_ASAP7_75t_L g187 ( .A(n_151), .Y(n_187) );
INVxp33_ASAP7_75t_SL g188 ( .A(n_170), .Y(n_188) );
NOR2xp33_ASAP7_75t_L g189 ( .A(n_157), .B(n_130), .Y(n_189) );
INVx2_ASAP7_75t_L g190 ( .A(n_158), .Y(n_190) );
INVx2_ASAP7_75t_L g191 ( .A(n_158), .Y(n_191) );
INVx2_ASAP7_75t_SL g192 ( .A(n_168), .Y(n_192) );
INVx2_ASAP7_75t_L g193 ( .A(n_152), .Y(n_193) );
INVx2_ASAP7_75t_L g194 ( .A(n_152), .Y(n_194) );
INVx2_ASAP7_75t_L g195 ( .A(n_152), .Y(n_195) );
INVx4_ASAP7_75t_L g196 ( .A(n_152), .Y(n_196) );
NAND2xp5_ASAP7_75t_L g197 ( .A(n_172), .B(n_116), .Y(n_197) );
INVx2_ASAP7_75t_L g198 ( .A(n_152), .Y(n_198) );
NAND2xp5_ASAP7_75t_L g199 ( .A(n_172), .B(n_138), .Y(n_199) );
INVx2_ASAP7_75t_L g200 ( .A(n_152), .Y(n_200) );
NOR2x1p5_ASAP7_75t_L g201 ( .A(n_155), .B(n_138), .Y(n_201) );
INVx2_ASAP7_75t_L g202 ( .A(n_152), .Y(n_202) );
INVx1_ASAP7_75t_SL g203 ( .A(n_169), .Y(n_203) );
AND2x2_ASAP7_75t_L g204 ( .A(n_155), .B(n_141), .Y(n_204) );
INVx2_ASAP7_75t_L g205 ( .A(n_171), .Y(n_205) );
INVx2_ASAP7_75t_L g206 ( .A(n_171), .Y(n_206) );
NOR2xp33_ASAP7_75t_L g207 ( .A(n_157), .B(n_135), .Y(n_207) );
NOR2x1p5_ASAP7_75t_L g208 ( .A(n_157), .B(n_141), .Y(n_208) );
BUFx6f_ASAP7_75t_L g209 ( .A(n_156), .Y(n_209) );
INVx1_ASAP7_75t_L g210 ( .A(n_151), .Y(n_210) );
INVx2_ASAP7_75t_L g211 ( .A(n_171), .Y(n_211) );
AND2x4_ASAP7_75t_L g212 ( .A(n_153), .B(n_136), .Y(n_212) );
INVx1_ASAP7_75t_L g213 ( .A(n_153), .Y(n_213) );
INVx1_ASAP7_75t_L g214 ( .A(n_171), .Y(n_214) );
NAND2xp5_ASAP7_75t_L g215 ( .A(n_172), .B(n_132), .Y(n_215) );
INVx3_ASAP7_75t_L g216 ( .A(n_171), .Y(n_216) );
NAND2xp5_ASAP7_75t_L g217 ( .A(n_160), .B(n_142), .Y(n_217) );
NAND2xp33_ASAP7_75t_SL g218 ( .A(n_150), .B(n_114), .Y(n_218) );
INVx2_ASAP7_75t_L g219 ( .A(n_171), .Y(n_219) );
INVx2_ASAP7_75t_L g220 ( .A(n_159), .Y(n_220) );
INVx2_ASAP7_75t_L g221 ( .A(n_159), .Y(n_221) );
INVx2_ASAP7_75t_SL g222 ( .A(n_168), .Y(n_222) );
BUFx10_ASAP7_75t_L g223 ( .A(n_169), .Y(n_223) );
INVx1_ASAP7_75t_L g224 ( .A(n_159), .Y(n_224) );
INVx2_ASAP7_75t_L g225 ( .A(n_156), .Y(n_225) );
INVx2_ASAP7_75t_L g226 ( .A(n_166), .Y(n_226) );
INVx2_ASAP7_75t_L g227 ( .A(n_186), .Y(n_227) );
NAND2xp5_ASAP7_75t_L g228 ( .A(n_215), .B(n_150), .Y(n_228) );
BUFx6f_ASAP7_75t_L g229 ( .A(n_181), .Y(n_229) );
NOR3xp33_ASAP7_75t_L g230 ( .A(n_218), .B(n_165), .C(n_163), .Y(n_230) );
INVx1_ASAP7_75t_L g231 ( .A(n_186), .Y(n_231) );
NAND2xp5_ASAP7_75t_L g232 ( .A(n_197), .B(n_160), .Y(n_232) );
NAND2xp5_ASAP7_75t_L g233 ( .A(n_199), .B(n_162), .Y(n_233) );
NAND2xp5_ASAP7_75t_L g234 ( .A(n_217), .B(n_162), .Y(n_234) );
AND2x2_ASAP7_75t_L g235 ( .A(n_203), .B(n_167), .Y(n_235) );
INVx2_ASAP7_75t_L g236 ( .A(n_187), .Y(n_236) );
INVx2_ASAP7_75t_L g237 ( .A(n_187), .Y(n_237) );
NAND2xp5_ASAP7_75t_L g238 ( .A(n_212), .B(n_164), .Y(n_238) );
NAND2xp5_ASAP7_75t_L g239 ( .A(n_212), .B(n_164), .Y(n_239) );
INVx2_ASAP7_75t_L g240 ( .A(n_210), .Y(n_240) );
NAND2xp5_ASAP7_75t_L g241 ( .A(n_212), .B(n_174), .Y(n_241) );
AND2x2_ASAP7_75t_L g242 ( .A(n_203), .B(n_223), .Y(n_242) );
INVxp67_ASAP7_75t_L g243 ( .A(n_185), .Y(n_243) );
NAND2xp5_ASAP7_75t_L g244 ( .A(n_212), .B(n_174), .Y(n_244) );
NAND2xp5_ASAP7_75t_SL g245 ( .A(n_181), .B(n_174), .Y(n_245) );
INVx1_ASAP7_75t_L g246 ( .A(n_210), .Y(n_246) );
NAND2xp5_ASAP7_75t_L g247 ( .A(n_185), .B(n_174), .Y(n_247) );
AND2x2_ASAP7_75t_L g248 ( .A(n_223), .B(n_204), .Y(n_248) );
NAND2xp5_ASAP7_75t_SL g249 ( .A(n_184), .B(n_166), .Y(n_249) );
NOR2xp67_ASAP7_75t_L g250 ( .A(n_224), .B(n_163), .Y(n_250) );
INVx2_ASAP7_75t_L g251 ( .A(n_179), .Y(n_251) );
INVx2_ASAP7_75t_L g252 ( .A(n_179), .Y(n_252) );
HB1xp67_ASAP7_75t_L g253 ( .A(n_204), .Y(n_253) );
INVxp67_ASAP7_75t_L g254 ( .A(n_223), .Y(n_254) );
NAND2xp5_ASAP7_75t_L g255 ( .A(n_184), .B(n_167), .Y(n_255) );
NAND2xp5_ASAP7_75t_L g256 ( .A(n_192), .B(n_173), .Y(n_256) );
BUFx6f_ASAP7_75t_SL g257 ( .A(n_223), .Y(n_257) );
NAND2xp5_ASAP7_75t_L g258 ( .A(n_192), .B(n_166), .Y(n_258) );
INVx1_ASAP7_75t_L g259 ( .A(n_224), .Y(n_259) );
NOR2xp33_ASAP7_75t_SL g260 ( .A(n_222), .B(n_114), .Y(n_260) );
NAND2xp5_ASAP7_75t_L g261 ( .A(n_222), .B(n_166), .Y(n_261) );
NAND2xp5_ASAP7_75t_L g262 ( .A(n_180), .B(n_166), .Y(n_262) );
NAND2xp5_ASAP7_75t_SL g263 ( .A(n_175), .B(n_166), .Y(n_263) );
NAND2xp5_ASAP7_75t_L g264 ( .A(n_189), .B(n_166), .Y(n_264) );
NAND2xp5_ASAP7_75t_L g265 ( .A(n_207), .B(n_208), .Y(n_265) );
NAND2xp5_ASAP7_75t_L g266 ( .A(n_208), .B(n_111), .Y(n_266) );
NAND2xp5_ASAP7_75t_L g267 ( .A(n_176), .B(n_119), .Y(n_267) );
NAND3xp33_ASAP7_75t_L g268 ( .A(n_213), .B(n_156), .C(n_161), .Y(n_268) );
NAND2xp33_ASAP7_75t_L g269 ( .A(n_209), .B(n_125), .Y(n_269) );
AOI22xp5_ASAP7_75t_L g270 ( .A1(n_201), .A2(n_137), .B1(n_123), .B2(n_124), .Y(n_270) );
INVxp67_ASAP7_75t_L g271 ( .A(n_201), .Y(n_271) );
OR2x2_ASAP7_75t_L g272 ( .A(n_220), .B(n_7), .Y(n_272) );
INVx1_ASAP7_75t_L g273 ( .A(n_179), .Y(n_273) );
INVx1_ASAP7_75t_L g274 ( .A(n_213), .Y(n_274) );
INVx2_ASAP7_75t_L g275 ( .A(n_179), .Y(n_275) );
INVx1_ASAP7_75t_L g276 ( .A(n_220), .Y(n_276) );
NAND2xp5_ASAP7_75t_SL g277 ( .A(n_175), .B(n_139), .Y(n_277) );
NOR2xp33_ASAP7_75t_L g278 ( .A(n_175), .B(n_128), .Y(n_278) );
INVx2_ASAP7_75t_L g279 ( .A(n_205), .Y(n_279) );
NAND2xp33_ASAP7_75t_L g280 ( .A(n_209), .B(n_134), .Y(n_280) );
NAND2xp5_ASAP7_75t_L g281 ( .A(n_175), .B(n_143), .Y(n_281) );
NAND2xp5_ASAP7_75t_L g282 ( .A(n_221), .B(n_140), .Y(n_282) );
NOR3xp33_ASAP7_75t_L g283 ( .A(n_221), .B(n_145), .C(n_146), .Y(n_283) );
INVx1_ASAP7_75t_SL g284 ( .A(n_188), .Y(n_284) );
AOI22xp33_ASAP7_75t_L g285 ( .A1(n_225), .A2(n_137), .B1(n_123), .B2(n_156), .Y(n_285) );
NAND2xp5_ASAP7_75t_L g286 ( .A(n_193), .B(n_156), .Y(n_286) );
INVx3_ASAP7_75t_L g287 ( .A(n_196), .Y(n_287) );
INVx1_ASAP7_75t_L g288 ( .A(n_226), .Y(n_288) );
INVx1_ASAP7_75t_L g289 ( .A(n_193), .Y(n_289) );
NAND2xp5_ASAP7_75t_L g290 ( .A(n_235), .B(n_225), .Y(n_290) );
INVx1_ASAP7_75t_L g291 ( .A(n_273), .Y(n_291) );
OAI21x1_ASAP7_75t_L g292 ( .A1(n_286), .A2(n_225), .B(n_268), .Y(n_292) );
O2A1O1Ixp33_ASAP7_75t_L g293 ( .A1(n_230), .A2(n_226), .B(n_195), .C(n_198), .Y(n_293) );
INVx3_ASAP7_75t_L g294 ( .A(n_227), .Y(n_294) );
O2A1O1Ixp33_ASAP7_75t_SL g295 ( .A1(n_245), .A2(n_249), .B(n_265), .C(n_258), .Y(n_295) );
INVx3_ASAP7_75t_L g296 ( .A(n_227), .Y(n_296) );
NAND2xp5_ASAP7_75t_SL g297 ( .A(n_242), .B(n_196), .Y(n_297) );
NAND2x1p5_ASAP7_75t_L g298 ( .A(n_242), .B(n_248), .Y(n_298) );
NAND2xp5_ASAP7_75t_L g299 ( .A(n_235), .B(n_209), .Y(n_299) );
O2A1O1Ixp33_ASAP7_75t_L g300 ( .A1(n_247), .A2(n_195), .B(n_202), .C(n_198), .Y(n_300) );
O2A1O1Ixp33_ASAP7_75t_L g301 ( .A1(n_243), .A2(n_200), .B(n_202), .C(n_194), .Y(n_301) );
BUFx4f_ASAP7_75t_L g302 ( .A(n_248), .Y(n_302) );
A2O1A1Ixp33_ASAP7_75t_L g303 ( .A1(n_274), .A2(n_209), .B(n_200), .C(n_194), .Y(n_303) );
AO21x1_ASAP7_75t_L g304 ( .A1(n_262), .A2(n_214), .B(n_191), .Y(n_304) );
NAND2xp5_ASAP7_75t_SL g305 ( .A(n_254), .B(n_196), .Y(n_305) );
AO21x1_ASAP7_75t_L g306 ( .A1(n_264), .A2(n_214), .B(n_191), .Y(n_306) );
NAND2xp5_ASAP7_75t_SL g307 ( .A(n_229), .B(n_196), .Y(n_307) );
INVx2_ASAP7_75t_L g308 ( .A(n_251), .Y(n_308) );
OAI21xp5_ASAP7_75t_L g309 ( .A1(n_273), .A2(n_193), .B(n_194), .Y(n_309) );
BUFx6f_ASAP7_75t_L g310 ( .A(n_229), .Y(n_310) );
BUFx12f_ASAP7_75t_L g311 ( .A(n_272), .Y(n_311) );
AOI21xp5_ASAP7_75t_L g312 ( .A1(n_245), .A2(n_209), .B(n_161), .Y(n_312) );
NAND2xp5_ASAP7_75t_L g313 ( .A(n_228), .B(n_161), .Y(n_313) );
INVx1_ASAP7_75t_L g314 ( .A(n_236), .Y(n_314) );
INVxp67_ASAP7_75t_L g315 ( .A(n_260), .Y(n_315) );
OAI21xp5_ASAP7_75t_L g316 ( .A1(n_241), .A2(n_161), .B(n_219), .Y(n_316) );
NAND2xp5_ASAP7_75t_L g317 ( .A(n_234), .B(n_216), .Y(n_317) );
AND2x4_ASAP7_75t_SL g318 ( .A(n_253), .B(n_154), .Y(n_318) );
NAND2xp5_ASAP7_75t_SL g319 ( .A(n_229), .B(n_113), .Y(n_319) );
CKINVDCx10_ASAP7_75t_R g320 ( .A(n_257), .Y(n_320) );
INVx1_ASAP7_75t_L g321 ( .A(n_236), .Y(n_321) );
INVx1_ASAP7_75t_L g322 ( .A(n_237), .Y(n_322) );
NAND2xp5_ASAP7_75t_L g323 ( .A(n_255), .B(n_216), .Y(n_323) );
AOI21xp5_ASAP7_75t_L g324 ( .A1(n_277), .A2(n_219), .B(n_211), .Y(n_324) );
AO21x1_ASAP7_75t_L g325 ( .A1(n_269), .A2(n_190), .B(n_191), .Y(n_325) );
NAND2xp5_ASAP7_75t_L g326 ( .A(n_238), .B(n_216), .Y(n_326) );
INVxp67_ASAP7_75t_L g327 ( .A(n_284), .Y(n_327) );
NOR2xp33_ASAP7_75t_SL g328 ( .A(n_257), .B(n_154), .Y(n_328) );
INVxp67_ASAP7_75t_L g329 ( .A(n_257), .Y(n_329) );
INVx2_ASAP7_75t_L g330 ( .A(n_251), .Y(n_330) );
INVx2_ASAP7_75t_SL g331 ( .A(n_272), .Y(n_331) );
O2A1O1Ixp33_ASAP7_75t_L g332 ( .A1(n_239), .A2(n_216), .B(n_211), .C(n_206), .Y(n_332) );
AOI21xp5_ASAP7_75t_L g333 ( .A1(n_277), .A2(n_206), .B(n_205), .Y(n_333) );
OAI21xp5_ASAP7_75t_L g334 ( .A1(n_244), .A2(n_190), .B(n_183), .Y(n_334) );
HB1xp67_ASAP7_75t_L g335 ( .A(n_237), .Y(n_335) );
AOI21xp5_ASAP7_75t_L g336 ( .A1(n_232), .A2(n_183), .B(n_182), .Y(n_336) );
AOI21xp5_ASAP7_75t_L g337 ( .A1(n_233), .A2(n_182), .B(n_178), .Y(n_337) );
INVxp67_ASAP7_75t_L g338 ( .A(n_270), .Y(n_338) );
AOI22xp5_ASAP7_75t_L g339 ( .A1(n_250), .A2(n_178), .B1(n_177), .B2(n_190), .Y(n_339) );
NAND2xp5_ASAP7_75t_L g340 ( .A(n_298), .B(n_285), .Y(n_340) );
OAI22xp5_ASAP7_75t_L g341 ( .A1(n_331), .A2(n_335), .B1(n_290), .B2(n_302), .Y(n_341) );
OAI21xp5_ASAP7_75t_L g342 ( .A1(n_312), .A2(n_275), .B(n_252), .Y(n_342) );
NAND2xp5_ASAP7_75t_L g343 ( .A(n_298), .B(n_240), .Y(n_343) );
AND2x4_ASAP7_75t_L g344 ( .A(n_329), .B(n_271), .Y(n_344) );
NAND2xp5_ASAP7_75t_L g345 ( .A(n_302), .B(n_240), .Y(n_345) );
O2A1O1Ixp5_ASAP7_75t_L g346 ( .A1(n_325), .A2(n_249), .B(n_256), .C(n_261), .Y(n_346) );
INVx1_ASAP7_75t_L g347 ( .A(n_290), .Y(n_347) );
AOI21xp5_ASAP7_75t_L g348 ( .A1(n_313), .A2(n_263), .B(n_269), .Y(n_348) );
NOR2xp33_ASAP7_75t_SL g349 ( .A(n_328), .B(n_278), .Y(n_349) );
OAI21xp5_ASAP7_75t_L g350 ( .A1(n_303), .A2(n_275), .B(n_252), .Y(n_350) );
BUFx2_ASAP7_75t_R g351 ( .A(n_320), .Y(n_351) );
NOR2xp67_ASAP7_75t_L g352 ( .A(n_327), .B(n_266), .Y(n_352) );
AOI21xp5_ASAP7_75t_L g353 ( .A1(n_295), .A2(n_263), .B(n_280), .Y(n_353) );
OAI22xp33_ASAP7_75t_L g354 ( .A1(n_328), .A2(n_259), .B1(n_231), .B2(n_246), .Y(n_354) );
AND2x4_ASAP7_75t_L g355 ( .A(n_318), .B(n_283), .Y(n_355) );
INVx3_ASAP7_75t_SL g356 ( .A(n_319), .Y(n_356) );
AO31x2_ASAP7_75t_L g357 ( .A1(n_304), .A2(n_177), .A3(n_282), .B(n_276), .Y(n_357) );
CKINVDCx5p33_ASAP7_75t_R g358 ( .A(n_311), .Y(n_358) );
OR2x6_ASAP7_75t_L g359 ( .A(n_315), .B(n_289), .Y(n_359) );
OR2x6_ASAP7_75t_L g360 ( .A(n_338), .B(n_289), .Y(n_360) );
AOI21xp5_ASAP7_75t_L g361 ( .A1(n_316), .A2(n_280), .B(n_281), .Y(n_361) );
AOI21xp5_ASAP7_75t_L g362 ( .A1(n_316), .A2(n_229), .B(n_267), .Y(n_362) );
AOI21xp5_ASAP7_75t_L g363 ( .A1(n_334), .A2(n_229), .B(n_287), .Y(n_363) );
O2A1O1Ixp5_ASAP7_75t_L g364 ( .A1(n_306), .A2(n_307), .B(n_334), .C(n_299), .Y(n_364) );
AOI21xp33_ASAP7_75t_L g365 ( .A1(n_299), .A2(n_288), .B(n_287), .Y(n_365) );
AOI21xp5_ASAP7_75t_L g366 ( .A1(n_336), .A2(n_287), .B(n_279), .Y(n_366) );
AOI21x1_ASAP7_75t_SL g367 ( .A1(n_323), .A2(n_54), .B(n_108), .Y(n_367) );
NAND2xp5_ASAP7_75t_L g368 ( .A(n_314), .B(n_8), .Y(n_368) );
AOI21xp33_ASAP7_75t_L g369 ( .A1(n_301), .A2(n_279), .B(n_10), .Y(n_369) );
AO31x2_ASAP7_75t_L g370 ( .A1(n_321), .A2(n_9), .A3(n_10), .B(n_11), .Y(n_370) );
OAI21x1_ASAP7_75t_L g371 ( .A1(n_367), .A2(n_292), .B(n_332), .Y(n_371) );
BUFx2_ASAP7_75t_R g372 ( .A(n_358), .Y(n_372) );
HB1xp67_ASAP7_75t_L g373 ( .A(n_360), .Y(n_373) );
OAI21x1_ASAP7_75t_L g374 ( .A1(n_362), .A2(n_300), .B(n_293), .Y(n_374) );
NAND2xp5_ASAP7_75t_L g375 ( .A(n_347), .B(n_291), .Y(n_375) );
AO21x2_ASAP7_75t_L g376 ( .A1(n_361), .A2(n_309), .B(n_337), .Y(n_376) );
OA21x2_ASAP7_75t_L g377 ( .A1(n_342), .A2(n_309), .B(n_322), .Y(n_377) );
OAI21xp5_ASAP7_75t_L g378 ( .A1(n_364), .A2(n_339), .B(n_317), .Y(n_378) );
NAND2x1p5_ASAP7_75t_L g379 ( .A(n_343), .B(n_294), .Y(n_379) );
INVx2_ASAP7_75t_L g380 ( .A(n_357), .Y(n_380) );
NAND2xp5_ASAP7_75t_L g381 ( .A(n_340), .B(n_294), .Y(n_381) );
OAI21x1_ASAP7_75t_L g382 ( .A1(n_348), .A2(n_333), .B(n_324), .Y(n_382) );
OAI21x1_ASAP7_75t_L g383 ( .A1(n_353), .A2(n_296), .B(n_308), .Y(n_383) );
BUFx4f_ASAP7_75t_L g384 ( .A(n_360), .Y(n_384) );
OAI21x1_ASAP7_75t_L g385 ( .A1(n_363), .A2(n_296), .B(n_330), .Y(n_385) );
AO21x2_ASAP7_75t_L g386 ( .A1(n_369), .A2(n_297), .B(n_326), .Y(n_386) );
BUFx6f_ASAP7_75t_L g387 ( .A(n_359), .Y(n_387) );
NAND2x1p5_ASAP7_75t_L g388 ( .A(n_345), .B(n_310), .Y(n_388) );
NOR2xp33_ASAP7_75t_L g389 ( .A(n_355), .B(n_305), .Y(n_389) );
AND2x4_ASAP7_75t_L g390 ( .A(n_359), .B(n_310), .Y(n_390) );
INVx1_ASAP7_75t_L g391 ( .A(n_368), .Y(n_391) );
INVx2_ASAP7_75t_L g392 ( .A(n_357), .Y(n_392) );
NOR2x1_ASAP7_75t_R g393 ( .A(n_351), .B(n_344), .Y(n_393) );
OR2x2_ASAP7_75t_L g394 ( .A(n_341), .B(n_310), .Y(n_394) );
AO21x2_ASAP7_75t_L g395 ( .A1(n_350), .A2(n_9), .B(n_12), .Y(n_395) );
OAI21x1_ASAP7_75t_L g396 ( .A1(n_346), .A2(n_59), .B(n_104), .Y(n_396) );
INVx1_ASAP7_75t_L g397 ( .A(n_370), .Y(n_397) );
OAI21x1_ASAP7_75t_L g398 ( .A1(n_366), .A2(n_56), .B(n_103), .Y(n_398) );
OAI21x1_ASAP7_75t_L g399 ( .A1(n_357), .A2(n_53), .B(n_102), .Y(n_399) );
NOR2xp33_ASAP7_75t_L g400 ( .A(n_354), .B(n_13), .Y(n_400) );
AND2x2_ASAP7_75t_L g401 ( .A(n_375), .B(n_370), .Y(n_401) );
OAI21x1_ASAP7_75t_L g402 ( .A1(n_371), .A2(n_365), .B(n_352), .Y(n_402) );
AND2x4_ASAP7_75t_L g403 ( .A(n_390), .B(n_370), .Y(n_403) );
INVx2_ASAP7_75t_L g404 ( .A(n_380), .Y(n_404) );
BUFx2_ASAP7_75t_L g405 ( .A(n_394), .Y(n_405) );
HB1xp67_ASAP7_75t_L g406 ( .A(n_384), .Y(n_406) );
OAI21x1_ASAP7_75t_L g407 ( .A1(n_371), .A2(n_349), .B(n_356), .Y(n_407) );
AOI21xp5_ASAP7_75t_L g408 ( .A1(n_380), .A2(n_344), .B(n_52), .Y(n_408) );
INVx2_ASAP7_75t_L g409 ( .A(n_380), .Y(n_409) );
INVx1_ASAP7_75t_L g410 ( .A(n_397), .Y(n_410) );
INVx2_ASAP7_75t_L g411 ( .A(n_392), .Y(n_411) );
BUFx10_ASAP7_75t_L g412 ( .A(n_390), .Y(n_412) );
BUFx12f_ASAP7_75t_L g413 ( .A(n_393), .Y(n_413) );
INVx3_ASAP7_75t_L g414 ( .A(n_390), .Y(n_414) );
AO21x2_ASAP7_75t_L g415 ( .A1(n_397), .A2(n_13), .B(n_14), .Y(n_415) );
INVx2_ASAP7_75t_L g416 ( .A(n_392), .Y(n_416) );
INVx4_ASAP7_75t_L g417 ( .A(n_384), .Y(n_417) );
BUFx6f_ASAP7_75t_L g418 ( .A(n_385), .Y(n_418) );
HB1xp67_ASAP7_75t_L g419 ( .A(n_384), .Y(n_419) );
INVx1_ASAP7_75t_L g420 ( .A(n_392), .Y(n_420) );
INVx2_ASAP7_75t_L g421 ( .A(n_385), .Y(n_421) );
OAI22xp5_ASAP7_75t_L g422 ( .A1(n_384), .A2(n_14), .B1(n_15), .B2(n_16), .Y(n_422) );
AOI22xp33_ASAP7_75t_L g423 ( .A1(n_391), .A2(n_15), .B1(n_16), .B2(n_17), .Y(n_423) );
INVx1_ASAP7_75t_L g424 ( .A(n_381), .Y(n_424) );
INVx2_ASAP7_75t_L g425 ( .A(n_383), .Y(n_425) );
OR2x6_ASAP7_75t_L g426 ( .A(n_387), .B(n_17), .Y(n_426) );
BUFx2_ASAP7_75t_L g427 ( .A(n_394), .Y(n_427) );
OA21x2_ASAP7_75t_L g428 ( .A1(n_399), .A2(n_26), .B(n_27), .Y(n_428) );
AND2x2_ASAP7_75t_L g429 ( .A(n_375), .B(n_391), .Y(n_429) );
INVx2_ASAP7_75t_L g430 ( .A(n_383), .Y(n_430) );
INVx1_ASAP7_75t_L g431 ( .A(n_381), .Y(n_431) );
OR2x2_ASAP7_75t_L g432 ( .A(n_373), .B(n_28), .Y(n_432) );
INVx1_ASAP7_75t_L g433 ( .A(n_395), .Y(n_433) );
INVx3_ASAP7_75t_L g434 ( .A(n_390), .Y(n_434) );
INVx2_ASAP7_75t_SL g435 ( .A(n_387), .Y(n_435) );
AND2x4_ASAP7_75t_L g436 ( .A(n_387), .B(n_376), .Y(n_436) );
INVx1_ASAP7_75t_L g437 ( .A(n_395), .Y(n_437) );
INVx1_ASAP7_75t_L g438 ( .A(n_395), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_377), .Y(n_439) );
HB1xp67_ASAP7_75t_L g440 ( .A(n_387), .Y(n_440) );
HB1xp67_ASAP7_75t_L g441 ( .A(n_387), .Y(n_441) );
INVx2_ASAP7_75t_L g442 ( .A(n_377), .Y(n_442) );
AND2x4_ASAP7_75t_L g443 ( .A(n_387), .B(n_30), .Y(n_443) );
CKINVDCx20_ASAP7_75t_R g444 ( .A(n_372), .Y(n_444) );
INVx1_ASAP7_75t_L g445 ( .A(n_377), .Y(n_445) );
INVx2_ASAP7_75t_SL g446 ( .A(n_379), .Y(n_446) );
INVx1_ASAP7_75t_L g447 ( .A(n_377), .Y(n_447) );
INVx1_ASAP7_75t_L g448 ( .A(n_399), .Y(n_448) );
INVx1_ASAP7_75t_L g449 ( .A(n_376), .Y(n_449) );
INVx1_ASAP7_75t_L g450 ( .A(n_410), .Y(n_450) );
INVx1_ASAP7_75t_L g451 ( .A(n_410), .Y(n_451) );
AND2x2_ASAP7_75t_L g452 ( .A(n_401), .B(n_376), .Y(n_452) );
INVx2_ASAP7_75t_L g453 ( .A(n_404), .Y(n_453) );
AND2x2_ASAP7_75t_L g454 ( .A(n_401), .B(n_379), .Y(n_454) );
INVx2_ASAP7_75t_L g455 ( .A(n_404), .Y(n_455) );
AND2x2_ASAP7_75t_L g456 ( .A(n_403), .B(n_379), .Y(n_456) );
NOR2x1_ASAP7_75t_L g457 ( .A(n_417), .B(n_400), .Y(n_457) );
INVx2_ASAP7_75t_L g458 ( .A(n_404), .Y(n_458) );
NAND2xp5_ASAP7_75t_L g459 ( .A(n_429), .B(n_389), .Y(n_459) );
INVx2_ASAP7_75t_L g460 ( .A(n_409), .Y(n_460) );
INVx1_ASAP7_75t_L g461 ( .A(n_420), .Y(n_461) );
INVx1_ASAP7_75t_L g462 ( .A(n_420), .Y(n_462) );
INVx1_ASAP7_75t_L g463 ( .A(n_409), .Y(n_463) );
OR2x2_ASAP7_75t_L g464 ( .A(n_405), .B(n_388), .Y(n_464) );
AND2x2_ASAP7_75t_L g465 ( .A(n_403), .B(n_378), .Y(n_465) );
HB1xp67_ASAP7_75t_L g466 ( .A(n_429), .Y(n_466) );
INVx2_ASAP7_75t_SL g467 ( .A(n_412), .Y(n_467) );
NAND2xp5_ASAP7_75t_L g468 ( .A(n_424), .B(n_393), .Y(n_468) );
INVx1_ASAP7_75t_L g469 ( .A(n_409), .Y(n_469) );
AND2x2_ASAP7_75t_L g470 ( .A(n_403), .B(n_378), .Y(n_470) );
AND2x4_ASAP7_75t_L g471 ( .A(n_436), .B(n_398), .Y(n_471) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_424), .B(n_386), .Y(n_472) );
AND2x2_ASAP7_75t_L g473 ( .A(n_403), .B(n_388), .Y(n_473) );
INVx1_ASAP7_75t_L g474 ( .A(n_411), .Y(n_474) );
NAND2xp5_ASAP7_75t_L g475 ( .A(n_431), .B(n_386), .Y(n_475) );
AND2x2_ASAP7_75t_L g476 ( .A(n_431), .B(n_388), .Y(n_476) );
AND2x2_ASAP7_75t_L g477 ( .A(n_405), .B(n_386), .Y(n_477) );
AND2x2_ASAP7_75t_L g478 ( .A(n_427), .B(n_374), .Y(n_478) );
INVx2_ASAP7_75t_L g479 ( .A(n_411), .Y(n_479) );
INVx1_ASAP7_75t_L g480 ( .A(n_411), .Y(n_480) );
NOR2xp33_ASAP7_75t_L g481 ( .A(n_413), .B(n_372), .Y(n_481) );
INVx1_ASAP7_75t_L g482 ( .A(n_416), .Y(n_482) );
NAND2xp5_ASAP7_75t_L g483 ( .A(n_406), .B(n_374), .Y(n_483) );
OAI22xp5_ASAP7_75t_L g484 ( .A1(n_426), .A2(n_398), .B1(n_396), .B2(n_382), .Y(n_484) );
INVx2_ASAP7_75t_L g485 ( .A(n_416), .Y(n_485) );
INVx2_ASAP7_75t_L g486 ( .A(n_416), .Y(n_486) );
INVx3_ASAP7_75t_L g487 ( .A(n_417), .Y(n_487) );
AND2x2_ASAP7_75t_L g488 ( .A(n_427), .B(n_396), .Y(n_488) );
INVx1_ASAP7_75t_L g489 ( .A(n_449), .Y(n_489) );
OR2x2_ASAP7_75t_L g490 ( .A(n_449), .B(n_382), .Y(n_490) );
AND2x2_ASAP7_75t_L g491 ( .A(n_436), .B(n_31), .Y(n_491) );
INVx1_ASAP7_75t_L g492 ( .A(n_439), .Y(n_492) );
OR2x2_ASAP7_75t_L g493 ( .A(n_414), .B(n_32), .Y(n_493) );
NOR2xp33_ASAP7_75t_L g494 ( .A(n_413), .B(n_33), .Y(n_494) );
INVx1_ASAP7_75t_L g495 ( .A(n_415), .Y(n_495) );
INVx1_ASAP7_75t_L g496 ( .A(n_415), .Y(n_496) );
INVx2_ASAP7_75t_L g497 ( .A(n_442), .Y(n_497) );
INVx1_ASAP7_75t_L g498 ( .A(n_439), .Y(n_498) );
AOI22xp33_ASAP7_75t_L g499 ( .A1(n_417), .A2(n_34), .B1(n_35), .B2(n_37), .Y(n_499) );
AND2x2_ASAP7_75t_L g500 ( .A(n_436), .B(n_38), .Y(n_500) );
INVx1_ASAP7_75t_L g501 ( .A(n_445), .Y(n_501) );
INVx1_ASAP7_75t_L g502 ( .A(n_445), .Y(n_502) );
INVx2_ASAP7_75t_L g503 ( .A(n_442), .Y(n_503) );
INVx1_ASAP7_75t_L g504 ( .A(n_447), .Y(n_504) );
INVx2_ASAP7_75t_L g505 ( .A(n_442), .Y(n_505) );
INVx2_ASAP7_75t_L g506 ( .A(n_447), .Y(n_506) );
INVx1_ASAP7_75t_L g507 ( .A(n_436), .Y(n_507) );
AND2x2_ASAP7_75t_L g508 ( .A(n_414), .B(n_39), .Y(n_508) );
INVx1_ASAP7_75t_L g509 ( .A(n_433), .Y(n_509) );
BUFx3_ASAP7_75t_L g510 ( .A(n_412), .Y(n_510) );
AND2x2_ASAP7_75t_L g511 ( .A(n_414), .B(n_40), .Y(n_511) );
INVx1_ASAP7_75t_L g512 ( .A(n_433), .Y(n_512) );
AOI22xp33_ASAP7_75t_L g513 ( .A1(n_417), .A2(n_41), .B1(n_42), .B2(n_43), .Y(n_513) );
AND2x2_ASAP7_75t_L g514 ( .A(n_414), .B(n_44), .Y(n_514) );
INVxp67_ASAP7_75t_SL g515 ( .A(n_440), .Y(n_515) );
INVx4_ASAP7_75t_L g516 ( .A(n_426), .Y(n_516) );
INVx2_ASAP7_75t_L g517 ( .A(n_421), .Y(n_517) );
INVx1_ASAP7_75t_L g518 ( .A(n_437), .Y(n_518) );
INVx2_ASAP7_75t_L g519 ( .A(n_421), .Y(n_519) );
AND2x2_ASAP7_75t_L g520 ( .A(n_434), .B(n_45), .Y(n_520) );
INVx1_ASAP7_75t_L g521 ( .A(n_437), .Y(n_521) );
INVx1_ASAP7_75t_L g522 ( .A(n_438), .Y(n_522) );
INVx1_ASAP7_75t_L g523 ( .A(n_438), .Y(n_523) );
AND2x4_ASAP7_75t_L g524 ( .A(n_434), .B(n_47), .Y(n_524) );
OR2x2_ASAP7_75t_L g525 ( .A(n_434), .B(n_60), .Y(n_525) );
AND2x2_ASAP7_75t_L g526 ( .A(n_434), .B(n_63), .Y(n_526) );
INVx2_ASAP7_75t_L g527 ( .A(n_421), .Y(n_527) );
INVx1_ASAP7_75t_L g528 ( .A(n_415), .Y(n_528) );
NOR2xp33_ASAP7_75t_L g529 ( .A(n_419), .B(n_105), .Y(n_529) );
AND2x2_ASAP7_75t_L g530 ( .A(n_441), .B(n_66), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_466), .B(n_435), .Y(n_531) );
INVx1_ASAP7_75t_L g532 ( .A(n_450), .Y(n_532) );
OR2x2_ASAP7_75t_L g533 ( .A(n_459), .B(n_435), .Y(n_533) );
OAI221xp5_ASAP7_75t_SL g534 ( .A1(n_468), .A2(n_426), .B1(n_432), .B2(n_423), .C(n_408), .Y(n_534) );
AOI22xp33_ASAP7_75t_L g535 ( .A1(n_516), .A2(n_422), .B1(n_426), .B2(n_444), .Y(n_535) );
OR2x2_ASAP7_75t_L g536 ( .A(n_454), .B(n_446), .Y(n_536) );
OR2x2_ASAP7_75t_L g537 ( .A(n_454), .B(n_446), .Y(n_537) );
AND2x2_ASAP7_75t_L g538 ( .A(n_476), .B(n_412), .Y(n_538) );
NAND3xp33_ASAP7_75t_L g539 ( .A(n_495), .B(n_426), .C(n_432), .Y(n_539) );
AND2x2_ASAP7_75t_L g540 ( .A(n_476), .B(n_412), .Y(n_540) );
NOR2x1_ASAP7_75t_SL g541 ( .A(n_510), .B(n_443), .Y(n_541) );
INVx4_ASAP7_75t_L g542 ( .A(n_516), .Y(n_542) );
NOR2xp33_ASAP7_75t_L g543 ( .A(n_457), .B(n_443), .Y(n_543) );
HB1xp67_ASAP7_75t_L g544 ( .A(n_463), .Y(n_544) );
AND2x4_ASAP7_75t_L g545 ( .A(n_507), .B(n_407), .Y(n_545) );
INVx2_ASAP7_75t_L g546 ( .A(n_497), .Y(n_546) );
NAND2xp5_ASAP7_75t_SL g547 ( .A(n_516), .B(n_443), .Y(n_547) );
INVx2_ASAP7_75t_L g548 ( .A(n_497), .Y(n_548) );
INVxp67_ASAP7_75t_SL g549 ( .A(n_453), .Y(n_549) );
INVx1_ASAP7_75t_L g550 ( .A(n_450), .Y(n_550) );
AND2x2_ASAP7_75t_L g551 ( .A(n_452), .B(n_443), .Y(n_551) );
INVx1_ASAP7_75t_L g552 ( .A(n_451), .Y(n_552) );
AND2x2_ASAP7_75t_L g553 ( .A(n_452), .B(n_402), .Y(n_553) );
BUFx2_ASAP7_75t_L g554 ( .A(n_510), .Y(n_554) );
INVx3_ASAP7_75t_L g555 ( .A(n_487), .Y(n_555) );
BUFx3_ASAP7_75t_L g556 ( .A(n_467), .Y(n_556) );
AND2x2_ASAP7_75t_L g557 ( .A(n_465), .B(n_402), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g558 ( .A(n_451), .B(n_448), .Y(n_558) );
INVx5_ASAP7_75t_L g559 ( .A(n_487), .Y(n_559) );
AOI22xp33_ASAP7_75t_L g560 ( .A1(n_481), .A2(n_448), .B1(n_428), .B2(n_425), .Y(n_560) );
INVx2_ASAP7_75t_L g561 ( .A(n_503), .Y(n_561) );
AND2x2_ASAP7_75t_L g562 ( .A(n_465), .B(n_407), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g563 ( .A(n_461), .B(n_425), .Y(n_563) );
BUFx2_ASAP7_75t_L g564 ( .A(n_467), .Y(n_564) );
INVx1_ASAP7_75t_L g565 ( .A(n_461), .Y(n_565) );
INVx2_ASAP7_75t_L g566 ( .A(n_503), .Y(n_566) );
OR2x2_ASAP7_75t_L g567 ( .A(n_464), .B(n_425), .Y(n_567) );
AND2x2_ASAP7_75t_L g568 ( .A(n_470), .B(n_428), .Y(n_568) );
INVx2_ASAP7_75t_L g569 ( .A(n_505), .Y(n_569) );
BUFx2_ASAP7_75t_L g570 ( .A(n_515), .Y(n_570) );
INVx2_ASAP7_75t_L g571 ( .A(n_505), .Y(n_571) );
BUFx2_ASAP7_75t_L g572 ( .A(n_487), .Y(n_572) );
INVx1_ASAP7_75t_L g573 ( .A(n_462), .Y(n_573) );
OR2x2_ASAP7_75t_L g574 ( .A(n_464), .B(n_430), .Y(n_574) );
INVx1_ASAP7_75t_L g575 ( .A(n_462), .Y(n_575) );
INVx1_ASAP7_75t_L g576 ( .A(n_492), .Y(n_576) );
INVx1_ASAP7_75t_L g577 ( .A(n_492), .Y(n_577) );
AND2x2_ASAP7_75t_L g578 ( .A(n_470), .B(n_428), .Y(n_578) );
AND2x2_ASAP7_75t_L g579 ( .A(n_456), .B(n_428), .Y(n_579) );
INVx1_ASAP7_75t_L g580 ( .A(n_498), .Y(n_580) );
OAI22xp5_ASAP7_75t_L g581 ( .A1(n_493), .A2(n_418), .B1(n_430), .B2(n_72), .Y(n_581) );
AND2x2_ASAP7_75t_L g582 ( .A(n_456), .B(n_418), .Y(n_582) );
INVx2_ASAP7_75t_L g583 ( .A(n_506), .Y(n_583) );
INVx1_ASAP7_75t_L g584 ( .A(n_498), .Y(n_584) );
INVx1_ASAP7_75t_L g585 ( .A(n_501), .Y(n_585) );
BUFx2_ASAP7_75t_L g586 ( .A(n_491), .Y(n_586) );
INVx2_ASAP7_75t_L g587 ( .A(n_506), .Y(n_587) );
AND2x2_ASAP7_75t_L g588 ( .A(n_473), .B(n_418), .Y(n_588) );
AND2x2_ASAP7_75t_L g589 ( .A(n_473), .B(n_418), .Y(n_589) );
AOI22xp33_ASAP7_75t_L g590 ( .A1(n_494), .A2(n_418), .B1(n_70), .B2(n_73), .Y(n_590) );
INVx2_ASAP7_75t_L g591 ( .A(n_453), .Y(n_591) );
INVx3_ASAP7_75t_L g592 ( .A(n_463), .Y(n_592) );
INVx2_ASAP7_75t_L g593 ( .A(n_455), .Y(n_593) );
INVx1_ASAP7_75t_L g594 ( .A(n_501), .Y(n_594) );
AND2x4_ASAP7_75t_SL g595 ( .A(n_524), .B(n_418), .Y(n_595) );
INVx1_ASAP7_75t_L g596 ( .A(n_502), .Y(n_596) );
OR2x2_ASAP7_75t_L g597 ( .A(n_469), .B(n_67), .Y(n_597) );
INVxp67_ASAP7_75t_SL g598 ( .A(n_455), .Y(n_598) );
BUFx2_ASAP7_75t_L g599 ( .A(n_491), .Y(n_599) );
AND2x2_ASAP7_75t_L g600 ( .A(n_500), .B(n_74), .Y(n_600) );
OAI22xp5_ASAP7_75t_L g601 ( .A1(n_493), .A2(n_75), .B1(n_78), .B2(n_79), .Y(n_601) );
INVxp67_ASAP7_75t_L g602 ( .A(n_528), .Y(n_602) );
AND2x2_ASAP7_75t_L g603 ( .A(n_500), .B(n_80), .Y(n_603) );
INVx1_ASAP7_75t_L g604 ( .A(n_502), .Y(n_604) );
INVx1_ASAP7_75t_SL g605 ( .A(n_530), .Y(n_605) );
INVx1_ASAP7_75t_L g606 ( .A(n_504), .Y(n_606) );
INVx2_ASAP7_75t_L g607 ( .A(n_458), .Y(n_607) );
AND2x4_ASAP7_75t_L g608 ( .A(n_507), .B(n_82), .Y(n_608) );
INVx1_ASAP7_75t_L g609 ( .A(n_504), .Y(n_609) );
INVx1_ASAP7_75t_L g610 ( .A(n_489), .Y(n_610) );
INVx2_ASAP7_75t_L g611 ( .A(n_458), .Y(n_611) );
BUFx3_ASAP7_75t_L g612 ( .A(n_469), .Y(n_612) );
NAND2xp5_ASAP7_75t_SL g613 ( .A(n_524), .B(n_471), .Y(n_613) );
INVx1_ASAP7_75t_L g614 ( .A(n_489), .Y(n_614) );
OR2x2_ASAP7_75t_L g615 ( .A(n_474), .B(n_85), .Y(n_615) );
INVx2_ASAP7_75t_L g616 ( .A(n_460), .Y(n_616) );
INVx1_ASAP7_75t_L g617 ( .A(n_509), .Y(n_617) );
INVx1_ASAP7_75t_L g618 ( .A(n_509), .Y(n_618) );
INVx1_ASAP7_75t_SL g619 ( .A(n_530), .Y(n_619) );
AND2x4_ASAP7_75t_L g620 ( .A(n_512), .B(n_86), .Y(n_620) );
OR2x2_ASAP7_75t_L g621 ( .A(n_474), .B(n_87), .Y(n_621) );
AND2x4_ASAP7_75t_L g622 ( .A(n_512), .B(n_89), .Y(n_622) );
NAND2xp5_ASAP7_75t_L g623 ( .A(n_477), .B(n_90), .Y(n_623) );
HB1xp67_ASAP7_75t_L g624 ( .A(n_480), .Y(n_624) );
AND2x2_ASAP7_75t_L g625 ( .A(n_478), .B(n_95), .Y(n_625) );
INVx1_ASAP7_75t_L g626 ( .A(n_518), .Y(n_626) );
AOI22xp33_ASAP7_75t_SL g627 ( .A1(n_508), .A2(n_96), .B1(n_99), .B2(n_100), .Y(n_627) );
AND2x2_ASAP7_75t_L g628 ( .A(n_478), .B(n_477), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g629 ( .A(n_480), .B(n_482), .Y(n_629) );
NOR2x1_ASAP7_75t_L g630 ( .A(n_525), .B(n_524), .Y(n_630) );
NAND2xp5_ASAP7_75t_SL g631 ( .A(n_471), .B(n_525), .Y(n_631) );
INVxp67_ASAP7_75t_L g632 ( .A(n_528), .Y(n_632) );
OAI22xp5_ASAP7_75t_L g633 ( .A1(n_529), .A2(n_499), .B1(n_513), .B2(n_520), .Y(n_633) );
INVx3_ASAP7_75t_L g634 ( .A(n_482), .Y(n_634) );
AND2x2_ASAP7_75t_L g635 ( .A(n_508), .B(n_520), .Y(n_635) );
AND2x2_ASAP7_75t_L g636 ( .A(n_511), .B(n_514), .Y(n_636) );
AND2x2_ASAP7_75t_L g637 ( .A(n_511), .B(n_514), .Y(n_637) );
OR2x2_ASAP7_75t_L g638 ( .A(n_570), .B(n_628), .Y(n_638) );
INVx1_ASAP7_75t_L g639 ( .A(n_532), .Y(n_639) );
AND2x2_ASAP7_75t_L g640 ( .A(n_586), .B(n_518), .Y(n_640) );
INVx2_ASAP7_75t_L g641 ( .A(n_583), .Y(n_641) );
INVx1_ASAP7_75t_L g642 ( .A(n_550), .Y(n_642) );
NOR2xp33_ASAP7_75t_L g643 ( .A(n_533), .B(n_521), .Y(n_643) );
INVx2_ASAP7_75t_L g644 ( .A(n_583), .Y(n_644) );
AND2x2_ASAP7_75t_L g645 ( .A(n_599), .B(n_521), .Y(n_645) );
AND2x2_ASAP7_75t_L g646 ( .A(n_553), .B(n_523), .Y(n_646) );
INVxp67_ASAP7_75t_L g647 ( .A(n_554), .Y(n_647) );
AND2x2_ASAP7_75t_L g648 ( .A(n_562), .B(n_523), .Y(n_648) );
AND2x2_ASAP7_75t_L g649 ( .A(n_557), .B(n_522), .Y(n_649) );
AND2x2_ASAP7_75t_L g650 ( .A(n_551), .B(n_522), .Y(n_650) );
NAND2xp5_ASAP7_75t_L g651 ( .A(n_552), .B(n_472), .Y(n_651) );
NAND2xp5_ASAP7_75t_L g652 ( .A(n_565), .B(n_475), .Y(n_652) );
AND2x4_ASAP7_75t_L g653 ( .A(n_542), .B(n_471), .Y(n_653) );
AND2x2_ASAP7_75t_L g654 ( .A(n_588), .B(n_488), .Y(n_654) );
AND2x2_ASAP7_75t_L g655 ( .A(n_589), .B(n_488), .Y(n_655) );
INVx2_ASAP7_75t_L g656 ( .A(n_587), .Y(n_656) );
NAND2xp5_ASAP7_75t_L g657 ( .A(n_573), .B(n_496), .Y(n_657) );
INVx2_ASAP7_75t_L g658 ( .A(n_587), .Y(n_658) );
HB1xp67_ASAP7_75t_L g659 ( .A(n_544), .Y(n_659) );
NAND2xp5_ASAP7_75t_L g660 ( .A(n_575), .B(n_576), .Y(n_660) );
INVx1_ASAP7_75t_L g661 ( .A(n_577), .Y(n_661) );
AND2x2_ASAP7_75t_L g662 ( .A(n_582), .B(n_490), .Y(n_662) );
NAND2xp5_ASAP7_75t_L g663 ( .A(n_580), .B(n_490), .Y(n_663) );
NAND2xp5_ASAP7_75t_L g664 ( .A(n_584), .B(n_460), .Y(n_664) );
AND2x2_ASAP7_75t_L g665 ( .A(n_605), .B(n_479), .Y(n_665) );
INVx2_ASAP7_75t_L g666 ( .A(n_546), .Y(n_666) );
BUFx3_ASAP7_75t_L g667 ( .A(n_556), .Y(n_667) );
INVx1_ASAP7_75t_L g668 ( .A(n_585), .Y(n_668) );
NAND2xp5_ASAP7_75t_L g669 ( .A(n_594), .B(n_479), .Y(n_669) );
OR2x2_ASAP7_75t_L g670 ( .A(n_536), .B(n_486), .Y(n_670) );
AND2x2_ASAP7_75t_L g671 ( .A(n_568), .B(n_486), .Y(n_671) );
INVx2_ASAP7_75t_SL g672 ( .A(n_559), .Y(n_672) );
NAND2xp5_ASAP7_75t_L g673 ( .A(n_596), .B(n_485), .Y(n_673) );
AND2x2_ASAP7_75t_L g674 ( .A(n_578), .B(n_485), .Y(n_674) );
INVx2_ASAP7_75t_L g675 ( .A(n_546), .Y(n_675) );
AND2x2_ASAP7_75t_L g676 ( .A(n_579), .B(n_483), .Y(n_676) );
INVxp67_ASAP7_75t_SL g677 ( .A(n_612), .Y(n_677) );
INVx2_ASAP7_75t_L g678 ( .A(n_548), .Y(n_678) );
INVx1_ASAP7_75t_L g679 ( .A(n_604), .Y(n_679) );
AND2x4_ASAP7_75t_SL g680 ( .A(n_542), .B(n_526), .Y(n_680) );
HB1xp67_ASAP7_75t_L g681 ( .A(n_544), .Y(n_681) );
OR2x2_ASAP7_75t_L g682 ( .A(n_537), .B(n_517), .Y(n_682) );
INVx2_ASAP7_75t_L g683 ( .A(n_548), .Y(n_683) );
AND2x4_ASAP7_75t_SL g684 ( .A(n_542), .B(n_526), .Y(n_684) );
AND2x2_ASAP7_75t_L g685 ( .A(n_619), .B(n_517), .Y(n_685) );
NOR2xp33_ASAP7_75t_SL g686 ( .A(n_556), .B(n_527), .Y(n_686) );
INVx1_ASAP7_75t_L g687 ( .A(n_606), .Y(n_687) );
BUFx2_ASAP7_75t_L g688 ( .A(n_564), .Y(n_688) );
AND2x2_ASAP7_75t_L g689 ( .A(n_635), .B(n_519), .Y(n_689) );
INVx2_ASAP7_75t_L g690 ( .A(n_561), .Y(n_690) );
OR2x2_ASAP7_75t_L g691 ( .A(n_612), .B(n_527), .Y(n_691) );
NAND2xp5_ASAP7_75t_L g692 ( .A(n_609), .B(n_519), .Y(n_692) );
AND2x4_ASAP7_75t_L g693 ( .A(n_613), .B(n_484), .Y(n_693) );
NOR2xp33_ASAP7_75t_SL g694 ( .A(n_559), .B(n_630), .Y(n_694) );
AND2x2_ASAP7_75t_L g695 ( .A(n_636), .B(n_637), .Y(n_695) );
INVx2_ASAP7_75t_L g696 ( .A(n_561), .Y(n_696) );
INVx1_ASAP7_75t_L g697 ( .A(n_610), .Y(n_697) );
NAND2xp5_ASAP7_75t_L g698 ( .A(n_614), .B(n_626), .Y(n_698) );
INVx1_ASAP7_75t_L g699 ( .A(n_617), .Y(n_699) );
INVx1_ASAP7_75t_L g700 ( .A(n_618), .Y(n_700) );
NAND2xp5_ASAP7_75t_L g701 ( .A(n_624), .B(n_531), .Y(n_701) );
INVx1_ASAP7_75t_L g702 ( .A(n_624), .Y(n_702) );
INVx1_ASAP7_75t_L g703 ( .A(n_592), .Y(n_703) );
INVx2_ASAP7_75t_SL g704 ( .A(n_559), .Y(n_704) );
NAND2xp5_ASAP7_75t_L g705 ( .A(n_592), .B(n_634), .Y(n_705) );
INVx1_ASAP7_75t_L g706 ( .A(n_634), .Y(n_706) );
AND2x2_ASAP7_75t_L g707 ( .A(n_538), .B(n_540), .Y(n_707) );
OR2x2_ASAP7_75t_L g708 ( .A(n_629), .B(n_549), .Y(n_708) );
AND2x2_ASAP7_75t_L g709 ( .A(n_549), .B(n_598), .Y(n_709) );
INVx2_ASAP7_75t_L g710 ( .A(n_566), .Y(n_710) );
INVx1_ASAP7_75t_L g711 ( .A(n_558), .Y(n_711) );
AND2x2_ASAP7_75t_L g712 ( .A(n_598), .B(n_566), .Y(n_712) );
NAND2xp5_ASAP7_75t_L g713 ( .A(n_572), .B(n_571), .Y(n_713) );
AND2x2_ASAP7_75t_L g714 ( .A(n_569), .B(n_571), .Y(n_714) );
AND2x2_ASAP7_75t_L g715 ( .A(n_569), .B(n_607), .Y(n_715) );
INVx1_ASAP7_75t_L g716 ( .A(n_563), .Y(n_716) );
NAND2xp5_ASAP7_75t_L g717 ( .A(n_602), .B(n_632), .Y(n_717) );
INVx2_ASAP7_75t_L g718 ( .A(n_591), .Y(n_718) );
NAND2xp5_ASAP7_75t_L g719 ( .A(n_602), .B(n_632), .Y(n_719) );
INVx1_ASAP7_75t_L g720 ( .A(n_620), .Y(n_720) );
AND2x2_ASAP7_75t_L g721 ( .A(n_591), .B(n_607), .Y(n_721) );
HB1xp67_ASAP7_75t_L g722 ( .A(n_593), .Y(n_722) );
AND2x2_ASAP7_75t_L g723 ( .A(n_593), .B(n_616), .Y(n_723) );
INVx2_ASAP7_75t_L g724 ( .A(n_611), .Y(n_724) );
AND2x2_ASAP7_75t_L g725 ( .A(n_611), .B(n_616), .Y(n_725) );
INVx1_ASAP7_75t_L g726 ( .A(n_620), .Y(n_726) );
BUFx2_ASAP7_75t_L g727 ( .A(n_559), .Y(n_727) );
INVx1_ASAP7_75t_L g728 ( .A(n_620), .Y(n_728) );
AND2x2_ASAP7_75t_L g729 ( .A(n_613), .B(n_545), .Y(n_729) );
INVx2_ASAP7_75t_L g730 ( .A(n_567), .Y(n_730) );
INVx1_ASAP7_75t_L g731 ( .A(n_622), .Y(n_731) );
INVx2_ASAP7_75t_SL g732 ( .A(n_555), .Y(n_732) );
INVx1_ASAP7_75t_L g733 ( .A(n_622), .Y(n_733) );
AND2x2_ASAP7_75t_L g734 ( .A(n_545), .B(n_574), .Y(n_734) );
INVx4_ASAP7_75t_L g735 ( .A(n_555), .Y(n_735) );
INVx1_ASAP7_75t_L g736 ( .A(n_622), .Y(n_736) );
INVx1_ASAP7_75t_L g737 ( .A(n_555), .Y(n_737) );
INVx1_ASAP7_75t_L g738 ( .A(n_608), .Y(n_738) );
INVx1_ASAP7_75t_SL g739 ( .A(n_600), .Y(n_739) );
OR2x2_ASAP7_75t_L g740 ( .A(n_631), .B(n_539), .Y(n_740) );
AND2x2_ASAP7_75t_L g741 ( .A(n_625), .B(n_543), .Y(n_741) );
AND2x2_ASAP7_75t_L g742 ( .A(n_545), .B(n_631), .Y(n_742) );
NAND2xp5_ASAP7_75t_L g743 ( .A(n_543), .B(n_535), .Y(n_743) );
NAND2xp5_ASAP7_75t_L g744 ( .A(n_535), .B(n_623), .Y(n_744) );
AND2x2_ASAP7_75t_L g745 ( .A(n_695), .B(n_595), .Y(n_745) );
AND2x4_ASAP7_75t_L g746 ( .A(n_735), .B(n_541), .Y(n_746) );
INVx1_ASAP7_75t_L g747 ( .A(n_701), .Y(n_747) );
NAND2xp5_ASAP7_75t_L g748 ( .A(n_716), .B(n_560), .Y(n_748) );
INVx1_ASAP7_75t_L g749 ( .A(n_639), .Y(n_749) );
INVx2_ASAP7_75t_L g750 ( .A(n_709), .Y(n_750) );
INVx2_ASAP7_75t_L g751 ( .A(n_709), .Y(n_751) );
INVx2_ASAP7_75t_L g752 ( .A(n_712), .Y(n_752) );
INVx3_ASAP7_75t_L g753 ( .A(n_735), .Y(n_753) );
INVx2_ASAP7_75t_L g754 ( .A(n_712), .Y(n_754) );
NAND2xp5_ASAP7_75t_L g755 ( .A(n_711), .B(n_560), .Y(n_755) );
AND2x4_ASAP7_75t_L g756 ( .A(n_735), .B(n_595), .Y(n_756) );
OR2x2_ASAP7_75t_L g757 ( .A(n_638), .B(n_547), .Y(n_757) );
INVx1_ASAP7_75t_L g758 ( .A(n_642), .Y(n_758) );
OR2x2_ASAP7_75t_L g759 ( .A(n_708), .B(n_547), .Y(n_759) );
NAND2xp5_ASAP7_75t_L g760 ( .A(n_646), .B(n_649), .Y(n_760) );
INVx1_ASAP7_75t_L g761 ( .A(n_661), .Y(n_761) );
AOI31xp33_ASAP7_75t_L g762 ( .A1(n_672), .A2(n_627), .A3(n_633), .B(n_590), .Y(n_762) );
INVx1_ASAP7_75t_L g763 ( .A(n_668), .Y(n_763) );
INVx2_ASAP7_75t_L g764 ( .A(n_691), .Y(n_764) );
NAND2xp5_ASAP7_75t_L g765 ( .A(n_646), .B(n_608), .Y(n_765) );
INVx1_ASAP7_75t_L g766 ( .A(n_679), .Y(n_766) );
NOR2xp33_ASAP7_75t_L g767 ( .A(n_743), .B(n_534), .Y(n_767) );
INVx1_ASAP7_75t_L g768 ( .A(n_687), .Y(n_768) );
AND2x2_ASAP7_75t_L g769 ( .A(n_734), .B(n_608), .Y(n_769) );
NAND2x1p5_ASAP7_75t_L g770 ( .A(n_667), .B(n_603), .Y(n_770) );
INVx2_ASAP7_75t_L g771 ( .A(n_722), .Y(n_771) );
AND2x2_ASAP7_75t_L g772 ( .A(n_734), .B(n_597), .Y(n_772) );
AND2x2_ASAP7_75t_L g773 ( .A(n_662), .B(n_615), .Y(n_773) );
AND2x4_ASAP7_75t_L g774 ( .A(n_729), .B(n_621), .Y(n_774) );
AOI21xp33_ASAP7_75t_SL g775 ( .A1(n_647), .A2(n_534), .B(n_627), .Y(n_775) );
AND2x2_ASAP7_75t_SL g776 ( .A(n_680), .B(n_590), .Y(n_776) );
NOR2x1_ASAP7_75t_L g777 ( .A(n_727), .B(n_601), .Y(n_777) );
INVx1_ASAP7_75t_L g778 ( .A(n_697), .Y(n_778) );
AND2x2_ASAP7_75t_L g779 ( .A(n_662), .B(n_581), .Y(n_779) );
BUFx2_ASAP7_75t_L g780 ( .A(n_667), .Y(n_780) );
OR2x2_ASAP7_75t_L g781 ( .A(n_649), .B(n_730), .Y(n_781) );
INVx1_ASAP7_75t_L g782 ( .A(n_699), .Y(n_782) );
NAND2xp5_ASAP7_75t_L g783 ( .A(n_702), .B(n_648), .Y(n_783) );
HB1xp67_ASAP7_75t_L g784 ( .A(n_659), .Y(n_784) );
INVx1_ASAP7_75t_L g785 ( .A(n_700), .Y(n_785) );
HB1xp67_ASAP7_75t_L g786 ( .A(n_659), .Y(n_786) );
INVx1_ASAP7_75t_L g787 ( .A(n_660), .Y(n_787) );
OR2x2_ASAP7_75t_L g788 ( .A(n_730), .B(n_648), .Y(n_788) );
INVx1_ASAP7_75t_L g789 ( .A(n_698), .Y(n_789) );
AND2x2_ASAP7_75t_L g790 ( .A(n_688), .B(n_654), .Y(n_790) );
OR2x2_ASAP7_75t_L g791 ( .A(n_670), .B(n_676), .Y(n_791) );
NAND5xp2_ASAP7_75t_L g792 ( .A(n_694), .B(n_744), .C(n_686), .D(n_731), .E(n_736), .Y(n_792) );
INVx1_ASAP7_75t_L g793 ( .A(n_681), .Y(n_793) );
OR2x2_ASAP7_75t_L g794 ( .A(n_676), .B(n_682), .Y(n_794) );
OAI22xp5_ASAP7_75t_L g795 ( .A1(n_680), .A2(n_684), .B1(n_739), .B2(n_677), .Y(n_795) );
INVx1_ASAP7_75t_L g796 ( .A(n_681), .Y(n_796) );
INVx1_ASAP7_75t_L g797 ( .A(n_717), .Y(n_797) );
NAND3xp33_ASAP7_75t_L g798 ( .A(n_740), .B(n_719), .C(n_706), .Y(n_798) );
INVx1_ASAP7_75t_L g799 ( .A(n_643), .Y(n_799) );
AND2x2_ASAP7_75t_L g800 ( .A(n_654), .B(n_655), .Y(n_800) );
INVx1_ASAP7_75t_L g801 ( .A(n_643), .Y(n_801) );
NAND5xp2_ASAP7_75t_SL g802 ( .A(n_729), .B(n_742), .C(n_741), .D(n_640), .E(n_645), .Y(n_802) );
AND2x2_ASAP7_75t_L g803 ( .A(n_655), .B(n_689), .Y(n_803) );
AND2x2_ASAP7_75t_L g804 ( .A(n_650), .B(n_707), .Y(n_804) );
INVx4_ASAP7_75t_L g805 ( .A(n_684), .Y(n_805) );
BUFx2_ASAP7_75t_L g806 ( .A(n_672), .Y(n_806) );
INVx1_ASAP7_75t_L g807 ( .A(n_663), .Y(n_807) );
HB1xp67_ASAP7_75t_L g808 ( .A(n_722), .Y(n_808) );
INVx2_ASAP7_75t_L g809 ( .A(n_641), .Y(n_809) );
NAND2xp5_ASAP7_75t_L g810 ( .A(n_651), .B(n_652), .Y(n_810) );
AND2x2_ASAP7_75t_L g811 ( .A(n_650), .B(n_742), .Y(n_811) );
OR2x2_ASAP7_75t_L g812 ( .A(n_671), .B(n_674), .Y(n_812) );
AND2x2_ASAP7_75t_L g813 ( .A(n_665), .B(n_671), .Y(n_813) );
INVx1_ASAP7_75t_L g814 ( .A(n_657), .Y(n_814) );
INVx2_ASAP7_75t_L g815 ( .A(n_641), .Y(n_815) );
NAND2xp5_ASAP7_75t_L g816 ( .A(n_714), .B(n_715), .Y(n_816) );
OAI22xp5_ASAP7_75t_L g817 ( .A1(n_693), .A2(n_704), .B1(n_738), .B2(n_728), .Y(n_817) );
INVx1_ASAP7_75t_L g818 ( .A(n_664), .Y(n_818) );
AND2x4_ASAP7_75t_L g819 ( .A(n_653), .B(n_693), .Y(n_819) );
INVx2_ASAP7_75t_L g820 ( .A(n_644), .Y(n_820) );
INVx2_ASAP7_75t_L g821 ( .A(n_644), .Y(n_821) );
OR2x2_ASAP7_75t_L g822 ( .A(n_674), .B(n_713), .Y(n_822) );
AND2x2_ASAP7_75t_L g823 ( .A(n_685), .B(n_693), .Y(n_823) );
NAND2xp5_ASAP7_75t_L g824 ( .A(n_714), .B(n_721), .Y(n_824) );
INVxp67_ASAP7_75t_L g825 ( .A(n_737), .Y(n_825) );
INVx1_ASAP7_75t_L g826 ( .A(n_783), .Y(n_826) );
A2O1A1O1Ixp25_ASAP7_75t_L g827 ( .A1(n_762), .A2(n_733), .B(n_726), .C(n_720), .D(n_703), .Y(n_827) );
OR2x2_ASAP7_75t_L g828 ( .A(n_812), .B(n_723), .Y(n_828) );
NAND2xp5_ASAP7_75t_L g829 ( .A(n_814), .B(n_723), .Y(n_829) );
INVxp67_ASAP7_75t_L g830 ( .A(n_780), .Y(n_830) );
NAND4xp25_ASAP7_75t_L g831 ( .A(n_767), .B(n_705), .C(n_653), .D(n_673), .Y(n_831) );
INVx1_ASAP7_75t_L g832 ( .A(n_783), .Y(n_832) );
INVx1_ASAP7_75t_L g833 ( .A(n_791), .Y(n_833) );
INVx1_ASAP7_75t_L g834 ( .A(n_794), .Y(n_834) );
AOI22xp5_ASAP7_75t_L g835 ( .A1(n_767), .A2(n_653), .B1(n_732), .B2(n_704), .Y(n_835) );
AOI32xp33_ASAP7_75t_L g836 ( .A1(n_777), .A2(n_732), .A3(n_725), .B1(n_721), .B2(n_715), .Y(n_836) );
NAND2xp5_ASAP7_75t_L g837 ( .A(n_755), .B(n_725), .Y(n_837) );
INVx1_ASAP7_75t_L g838 ( .A(n_749), .Y(n_838) );
INVx1_ASAP7_75t_L g839 ( .A(n_758), .Y(n_839) );
INVx1_ASAP7_75t_L g840 ( .A(n_761), .Y(n_840) );
NAND3xp33_ASAP7_75t_L g841 ( .A(n_798), .B(n_692), .C(n_669), .Y(n_841) );
OAI33xp33_ASAP7_75t_L g842 ( .A1(n_817), .A2(n_656), .A3(n_658), .B1(n_666), .B2(n_675), .B3(n_678), .Y(n_842) );
INVx1_ASAP7_75t_L g843 ( .A(n_763), .Y(n_843) );
AND2x2_ASAP7_75t_L g844 ( .A(n_823), .B(n_656), .Y(n_844) );
INVx1_ASAP7_75t_L g845 ( .A(n_766), .Y(n_845) );
AND2x2_ASAP7_75t_L g846 ( .A(n_790), .B(n_658), .Y(n_846) );
AND2x2_ASAP7_75t_L g847 ( .A(n_811), .B(n_666), .Y(n_847) );
AOI21xp33_ASAP7_75t_L g848 ( .A1(n_762), .A2(n_675), .B(n_678), .Y(n_848) );
INVx1_ASAP7_75t_L g849 ( .A(n_768), .Y(n_849) );
AOI211xp5_ASAP7_75t_L g850 ( .A1(n_795), .A2(n_683), .B(n_690), .C(n_696), .Y(n_850) );
INVx1_ASAP7_75t_L g851 ( .A(n_778), .Y(n_851) );
INVx1_ASAP7_75t_L g852 ( .A(n_782), .Y(n_852) );
AND2x2_ASAP7_75t_L g853 ( .A(n_819), .B(n_683), .Y(n_853) );
AOI321xp33_ASAP7_75t_L g854 ( .A1(n_775), .A2(n_690), .A3(n_696), .B1(n_710), .B2(n_718), .C(n_724), .Y(n_854) );
INVx2_ASAP7_75t_L g855 ( .A(n_808), .Y(n_855) );
INVx2_ASAP7_75t_L g856 ( .A(n_808), .Y(n_856) );
AND2x2_ASAP7_75t_L g857 ( .A(n_819), .B(n_710), .Y(n_857) );
INVx1_ASAP7_75t_L g858 ( .A(n_785), .Y(n_858) );
INVx1_ASAP7_75t_L g859 ( .A(n_818), .Y(n_859) );
INVx1_ASAP7_75t_L g860 ( .A(n_760), .Y(n_860) );
NOR4xp25_ASAP7_75t_L g861 ( .A(n_798), .B(n_718), .C(n_724), .D(n_797), .Y(n_861) );
INVx1_ASAP7_75t_L g862 ( .A(n_760), .Y(n_862) );
INVx2_ASAP7_75t_SL g863 ( .A(n_805), .Y(n_863) );
INVx1_ASAP7_75t_L g864 ( .A(n_793), .Y(n_864) );
AOI211x1_ASAP7_75t_SL g865 ( .A1(n_817), .A2(n_795), .B(n_755), .C(n_748), .Y(n_865) );
NAND2xp5_ASAP7_75t_L g866 ( .A(n_748), .B(n_796), .Y(n_866) );
INVx1_ASAP7_75t_L g867 ( .A(n_816), .Y(n_867) );
INVx1_ASAP7_75t_L g868 ( .A(n_816), .Y(n_868) );
AND2x2_ASAP7_75t_L g869 ( .A(n_800), .B(n_813), .Y(n_869) );
NAND2xp5_ASAP7_75t_L g870 ( .A(n_807), .B(n_789), .Y(n_870) );
NOR2xp67_ASAP7_75t_L g871 ( .A(n_805), .B(n_792), .Y(n_871) );
OAI22xp33_ASAP7_75t_L g872 ( .A1(n_770), .A2(n_753), .B1(n_802), .B2(n_806), .Y(n_872) );
INVx1_ASAP7_75t_L g873 ( .A(n_824), .Y(n_873) );
OAI211xp5_ASAP7_75t_SL g874 ( .A1(n_865), .A2(n_747), .B(n_801), .C(n_799), .Y(n_874) );
AOI221xp5_ASAP7_75t_L g875 ( .A1(n_848), .A2(n_787), .B1(n_810), .B2(n_825), .C(n_784), .Y(n_875) );
OAI31xp33_ASAP7_75t_L g876 ( .A1(n_848), .A2(n_792), .A3(n_770), .B(n_746), .Y(n_876) );
INVx1_ASAP7_75t_L g877 ( .A(n_829), .Y(n_877) );
OR2x2_ASAP7_75t_L g878 ( .A(n_837), .B(n_824), .Y(n_878) );
AND2x2_ASAP7_75t_L g879 ( .A(n_863), .B(n_803), .Y(n_879) );
INVx1_ASAP7_75t_L g880 ( .A(n_829), .Y(n_880) );
INVx1_ASAP7_75t_L g881 ( .A(n_870), .Y(n_881) );
INVx1_ASAP7_75t_SL g882 ( .A(n_870), .Y(n_882) );
OAI322xp33_ASAP7_75t_L g883 ( .A1(n_872), .A2(n_810), .A3(n_757), .B1(n_759), .B2(n_750), .C1(n_751), .C2(n_825), .Y(n_883) );
NOR3xp33_ASAP7_75t_L g884 ( .A(n_831), .B(n_784), .C(n_786), .Y(n_884) );
OAI31xp33_ASAP7_75t_L g885 ( .A1(n_831), .A2(n_746), .A3(n_753), .B(n_786), .Y(n_885) );
NAND2xp5_ASAP7_75t_L g886 ( .A(n_866), .B(n_804), .Y(n_886) );
INVx1_ASAP7_75t_L g887 ( .A(n_867), .Y(n_887) );
OAI221xp5_ASAP7_75t_L g888 ( .A1(n_836), .A2(n_765), .B1(n_764), .B2(n_754), .C(n_752), .Y(n_888) );
NAND2xp5_ASAP7_75t_L g889 ( .A(n_866), .B(n_773), .Y(n_889) );
INVx1_ASAP7_75t_L g890 ( .A(n_868), .Y(n_890) );
AOI21xp33_ASAP7_75t_L g891 ( .A1(n_830), .A2(n_776), .B(n_779), .Y(n_891) );
OAI21xp33_ASAP7_75t_SL g892 ( .A1(n_871), .A2(n_745), .B(n_765), .Y(n_892) );
OR2x2_ASAP7_75t_L g893 ( .A(n_837), .B(n_788), .Y(n_893) );
INVx1_ASAP7_75t_L g894 ( .A(n_873), .Y(n_894) );
AOI21xp33_ASAP7_75t_L g895 ( .A1(n_859), .A2(n_771), .B(n_774), .Y(n_895) );
AOI22xp33_ASAP7_75t_L g896 ( .A1(n_860), .A2(n_862), .B1(n_832), .B2(n_826), .Y(n_896) );
INVx1_ASAP7_75t_L g897 ( .A(n_864), .Y(n_897) );
OAI21xp5_ASAP7_75t_L g898 ( .A1(n_827), .A2(n_781), .B(n_756), .Y(n_898) );
INVxp67_ASAP7_75t_L g899 ( .A(n_841), .Y(n_899) );
INVx2_ASAP7_75t_L g900 ( .A(n_879), .Y(n_900) );
OAI221xp5_ASAP7_75t_SL g901 ( .A1(n_885), .A2(n_835), .B1(n_854), .B2(n_850), .C(n_861), .Y(n_901) );
OAI32xp33_ASAP7_75t_L g902 ( .A1(n_892), .A2(n_834), .A3(n_833), .B1(n_828), .B2(n_855), .Y(n_902) );
NAND2xp5_ASAP7_75t_SL g903 ( .A(n_876), .B(n_861), .Y(n_903) );
NAND3xp33_ASAP7_75t_L g904 ( .A(n_899), .B(n_856), .C(n_839), .Y(n_904) );
AOI221x1_ASAP7_75t_L g905 ( .A1(n_874), .A2(n_843), .B1(n_858), .B2(n_838), .C(n_840), .Y(n_905) );
AOI211xp5_ASAP7_75t_L g906 ( .A1(n_883), .A2(n_842), .B(n_756), .C(n_845), .Y(n_906) );
OAI221xp5_ASAP7_75t_L g907 ( .A1(n_898), .A2(n_852), .B1(n_851), .B2(n_849), .C(n_857), .Y(n_907) );
OAI211xp5_ASAP7_75t_L g908 ( .A1(n_899), .A2(n_853), .B(n_769), .C(n_869), .Y(n_908) );
NOR2xp33_ASAP7_75t_L g909 ( .A(n_874), .B(n_822), .Y(n_909) );
OAI21xp33_ASAP7_75t_SL g910 ( .A1(n_875), .A2(n_846), .B(n_844), .Y(n_910) );
NAND2xp5_ASAP7_75t_L g911 ( .A(n_881), .B(n_847), .Y(n_911) );
OAI222xp33_ASAP7_75t_L g912 ( .A1(n_888), .A2(n_774), .B1(n_772), .B2(n_809), .C1(n_815), .C2(n_820), .Y(n_912) );
OR2x2_ASAP7_75t_L g913 ( .A(n_878), .B(n_821), .Y(n_913) );
NOR3xp33_ASAP7_75t_L g914 ( .A(n_903), .B(n_891), .C(n_884), .Y(n_914) );
INVx2_ASAP7_75t_L g915 ( .A(n_913), .Y(n_915) );
INVx1_ASAP7_75t_L g916 ( .A(n_911), .Y(n_916) );
NOR3xp33_ASAP7_75t_L g917 ( .A(n_907), .B(n_884), .C(n_882), .Y(n_917) );
INVx1_ASAP7_75t_L g918 ( .A(n_911), .Y(n_918) );
NOR2xp33_ASAP7_75t_L g919 ( .A(n_909), .B(n_877), .Y(n_919) );
NAND3xp33_ASAP7_75t_SL g920 ( .A(n_906), .B(n_896), .C(n_880), .Y(n_920) );
NAND2xp5_ASAP7_75t_L g921 ( .A(n_914), .B(n_905), .Y(n_921) );
INVx1_ASAP7_75t_L g922 ( .A(n_916), .Y(n_922) );
AOI211x1_ASAP7_75t_L g923 ( .A1(n_920), .A2(n_902), .B(n_912), .C(n_908), .Y(n_923) );
NOR2x1_ASAP7_75t_L g924 ( .A(n_918), .B(n_904), .Y(n_924) );
HB1xp67_ASAP7_75t_L g925 ( .A(n_922), .Y(n_925) );
INVx1_ASAP7_75t_L g926 ( .A(n_924), .Y(n_926) );
NAND4xp75_ASAP7_75t_L g927 ( .A(n_923), .B(n_910), .C(n_919), .D(n_915), .Y(n_927) );
INVx2_ASAP7_75t_L g928 ( .A(n_926), .Y(n_928) );
NAND4xp75_ASAP7_75t_L g929 ( .A(n_927), .B(n_921), .C(n_917), .D(n_900), .Y(n_929) );
INVx1_ASAP7_75t_L g930 ( .A(n_928), .Y(n_930) );
OR2x2_ASAP7_75t_L g931 ( .A(n_929), .B(n_925), .Y(n_931) );
CKINVDCx20_ASAP7_75t_R g932 ( .A(n_931), .Y(n_932) );
INVx1_ASAP7_75t_L g933 ( .A(n_930), .Y(n_933) );
INVx1_ASAP7_75t_L g934 ( .A(n_933), .Y(n_934) );
OAI22xp33_ASAP7_75t_SL g935 ( .A1(n_934), .A2(n_932), .B1(n_901), .B2(n_894), .Y(n_935) );
OAI22xp5_ASAP7_75t_L g936 ( .A1(n_935), .A2(n_886), .B1(n_887), .B2(n_890), .Y(n_936) );
NAND2xp5_ASAP7_75t_L g937 ( .A(n_936), .B(n_897), .Y(n_937) );
OR2x6_ASAP7_75t_L g938 ( .A(n_937), .B(n_893), .Y(n_938) );
UNKNOWN g939 ( );
AOI21xp5_ASAP7_75t_L g940 ( .A1(n_939), .A2(n_889), .B(n_895), .Y(n_940) );
endmodule