module fake_jpeg_1930_n_94 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_94);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_94;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

INVx1_ASAP7_75t_L g11 ( 
.A(n_4),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_5),
.Y(n_12)
);

INVx1_ASAP7_75t_SL g13 ( 
.A(n_7),
.Y(n_13)
);

HB1xp67_ASAP7_75t_L g14 ( 
.A(n_10),
.Y(n_14)
);

BUFx12f_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g16 ( 
.A(n_9),
.B(n_10),
.Y(n_16)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_8),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_4),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_4),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_16),
.B(n_0),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_SL g41 ( 
.A(n_23),
.B(n_33),
.Y(n_41)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_24),
.Y(n_45)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_17),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_25),
.Y(n_37)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_17),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_26),
.Y(n_43)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_27),
.Y(n_34)
);

INVx5_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_28),
.B(n_29),
.Y(n_40)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_18),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_30),
.B(n_31),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_18),
.Y(n_31)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_22),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_32),
.B(n_21),
.Y(n_44)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

AOI22xp33_ASAP7_75t_SL g35 ( 
.A1(n_33),
.A2(n_13),
.B1(n_22),
.B2(n_12),
.Y(n_35)
);

INVxp67_ASAP7_75t_L g59 ( 
.A(n_35),
.Y(n_59)
);

MAJIxp5_ASAP7_75t_L g36 ( 
.A(n_30),
.B(n_16),
.C(n_14),
.Y(n_36)
);

MAJIxp5_ASAP7_75t_L g49 ( 
.A(n_36),
.B(n_38),
.C(n_21),
.Y(n_49)
);

MAJIxp5_ASAP7_75t_L g38 ( 
.A(n_24),
.B(n_13),
.C(n_12),
.Y(n_38)
);

NOR2x1_ASAP7_75t_L g39 ( 
.A(n_32),
.B(n_11),
.Y(n_39)
);

OR2x2_ASAP7_75t_L g52 ( 
.A(n_39),
.B(n_44),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_31),
.B(n_19),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_46),
.B(n_47),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_28),
.B(n_19),
.Y(n_47)
);

MAJIxp5_ASAP7_75t_L g69 ( 
.A(n_49),
.B(n_55),
.C(n_34),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_41),
.B(n_20),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_50),
.B(n_57),
.Y(n_63)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_51),
.Y(n_61)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_53),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_41),
.A2(n_29),
.B1(n_20),
.B2(n_2),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_54),
.A2(n_37),
.B1(n_43),
.B2(n_45),
.Y(n_64)
);

OR2x2_ASAP7_75t_SL g55 ( 
.A(n_36),
.B(n_0),
.Y(n_55)
);

OAI21xp5_ASAP7_75t_L g56 ( 
.A1(n_39),
.A2(n_1),
.B(n_2),
.Y(n_56)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_56),
.B(n_60),
.C(n_45),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_38),
.B(n_6),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_42),
.B(n_7),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_58),
.B(n_8),
.Y(n_62)
);

OR2x4_ASAP7_75t_L g60 ( 
.A(n_40),
.B(n_1),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_62),
.B(n_67),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_64),
.A2(n_59),
.B1(n_53),
.B2(n_51),
.Y(n_75)
);

NOR3xp33_ASAP7_75t_L g70 ( 
.A(n_65),
.B(n_69),
.C(n_60),
.Y(n_70)
);

MAJIxp5_ASAP7_75t_L g66 ( 
.A(n_49),
.B(n_43),
.C(n_34),
.Y(n_66)
);

XOR2xp5_ASAP7_75t_L g74 ( 
.A(n_66),
.B(n_59),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_48),
.B(n_43),
.Y(n_67)
);

XOR2xp5_ASAP7_75t_L g80 ( 
.A(n_70),
.B(n_73),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_63),
.B(n_52),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_72),
.B(n_74),
.Y(n_79)
);

XNOR2xp5_ASAP7_75t_SL g73 ( 
.A(n_66),
.B(n_55),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_75),
.A2(n_68),
.B1(n_54),
.B2(n_56),
.Y(n_78)
);

HB1xp67_ASAP7_75t_L g76 ( 
.A(n_61),
.Y(n_76)
);

CKINVDCx16_ASAP7_75t_R g77 ( 
.A(n_76),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_78),
.A2(n_82),
.B1(n_3),
.B2(n_5),
.Y(n_85)
);

INVx13_ASAP7_75t_L g81 ( 
.A(n_74),
.Y(n_81)
);

HB1xp67_ASAP7_75t_L g83 ( 
.A(n_81),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_73),
.A2(n_65),
.B1(n_52),
.B2(n_5),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_80),
.B(n_71),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_84),
.B(n_85),
.Y(n_88)
);

NAND3xp33_ASAP7_75t_L g86 ( 
.A(n_82),
.B(n_9),
.C(n_3),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_L g87 ( 
.A1(n_86),
.A2(n_79),
.B(n_78),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_SL g90 ( 
.A1(n_87),
.A2(n_81),
.B(n_77),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_83),
.B(n_80),
.C(n_79),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_L g91 ( 
.A1(n_89),
.A2(n_77),
.B(n_81),
.Y(n_91)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_90),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_92),
.B(n_91),
.C(n_88),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_93),
.B(n_3),
.Y(n_94)
);


endmodule