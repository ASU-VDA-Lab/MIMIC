module real_jpeg_24581_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_249;
wire n_215;
wire n_166;
wire n_176;
wire n_221;
wire n_288;
wire n_286;
wire n_292;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_280;
wire n_64;
wire n_177;
wire n_291;
wire n_236;
wire n_47;
wire n_131;
wire n_271;
wire n_281;
wire n_276;
wire n_163;
wire n_22;
wire n_287;
wire n_237;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_299;
wire n_173;
wire n_243;
wire n_115;
wire n_255;
wire n_98;
wire n_27;
wire n_56;
wire n_293;
wire n_48;
wire n_164;
wire n_184;
wire n_200;
wire n_275;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_13;
wire n_113;
wire n_155;
wire n_120;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_267;
wire n_208;
wire n_62;
wire n_239;
wire n_290;
wire n_162;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_172;
wire n_211;
wire n_285;
wire n_45;
wire n_160;
wire n_112;
wire n_42;
wire n_268;
wire n_145;
wire n_18;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_294;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_298;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_296;
wire n_134;
wire n_270;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_203;
wire n_192;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_110;
wire n_61;
wire n_195;
wire n_205;
wire n_258;
wire n_289;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_150;
wire n_74;
wire n_32;
wire n_20;
wire n_228;
wire n_80;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_225;
wire n_103;
wire n_259;
wire n_232;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_284;
wire n_226;
wire n_277;
wire n_185;
wire n_240;
wire n_125;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_297;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_169;
wire n_88;
wire n_59;
wire n_279;
wire n_128;
wire n_167;
wire n_213;
wire n_179;
wire n_295;
wire n_202;
wire n_133;
wire n_216;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_210;
wire n_206;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_283;
wire n_181;
wire n_101;
wire n_274;
wire n_256;
wire n_182;
wire n_253;
wire n_96;
wire n_269;
wire n_273;
wire n_89;
wire n_16;

INVx3_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_1),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_2),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_L g33 ( 
.A1(n_3),
.A2(n_19),
.B1(n_22),
.B2(n_34),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_3),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_L g51 ( 
.A1(n_3),
.A2(n_26),
.B1(n_27),
.B2(n_34),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_3),
.A2(n_34),
.B1(n_60),
.B2(n_63),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_3),
.A2(n_34),
.B1(n_44),
.B2(n_46),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g38 ( 
.A1(n_4),
.A2(n_26),
.B1(n_27),
.B2(n_39),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_4),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_4),
.A2(n_39),
.B1(n_56),
.B2(n_57),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_4),
.A2(n_39),
.B1(n_44),
.B2(n_46),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_4),
.A2(n_19),
.B1(n_22),
.B2(n_39),
.Y(n_101)
);

O2A1O1Ixp33_ASAP7_75t_L g184 ( 
.A1(n_4),
.A2(n_62),
.B(n_185),
.C(n_186),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_4),
.B(n_65),
.Y(n_200)
);

O2A1O1Ixp33_ASAP7_75t_L g210 ( 
.A1(n_4),
.A2(n_22),
.B(n_25),
.C(n_211),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_4),
.B(n_43),
.C(n_44),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_4),
.B(n_23),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_4),
.B(n_145),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g255 ( 
.A(n_4),
.B(n_41),
.Y(n_255)
);

BUFx10_ASAP7_75t_L g62 ( 
.A(n_5),
.Y(n_62)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

INVx13_ASAP7_75t_L g57 ( 
.A(n_7),
.Y(n_57)
);

OAI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_8),
.A2(n_57),
.B1(n_60),
.B2(n_129),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_8),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_8),
.A2(n_19),
.B1(n_22),
.B2(n_129),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_8),
.A2(n_26),
.B1(n_27),
.B2(n_129),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_8),
.A2(n_44),
.B1(n_46),
.B2(n_129),
.Y(n_240)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_SL g18 ( 
.A1(n_10),
.A2(n_19),
.B1(n_21),
.B2(n_22),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_10),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_10),
.A2(n_21),
.B1(n_26),
.B2(n_27),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_10),
.A2(n_21),
.B1(n_64),
.B2(n_104),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_10),
.A2(n_21),
.B1(n_44),
.B2(n_46),
.Y(n_141)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_11),
.Y(n_81)
);

INVx6_ASAP7_75t_L g82 ( 
.A(n_11),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_11),
.B(n_119),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_11),
.B(n_240),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_110),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_SL g13 ( 
.A(n_14),
.B(n_109),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_93),
.Y(n_14)
);

OR2x2_ASAP7_75t_L g109 ( 
.A(n_15),
.B(n_93),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_15),
.B(n_298),
.Y(n_297)
);

OR2x2_ASAP7_75t_L g299 ( 
.A(n_15),
.B(n_298),
.Y(n_299)
);

FAx1_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_52),
.CI(n_78),
.CON(n_15),
.SN(n_15)
);

OAI21xp5_ASAP7_75t_SL g157 ( 
.A1(n_16),
.A2(n_17),
.B(n_35),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_35),
.Y(n_16)
);

AOI21xp5_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_23),
.B(n_30),
.Y(n_17)
);

AOI21xp5_ASAP7_75t_L g70 ( 
.A1(n_18),
.A2(n_71),
.B(n_72),
.Y(n_70)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_19),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_L g32 ( 
.A1(n_19),
.A2(n_22),
.B1(n_25),
.B2(n_29),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_19),
.A2(n_22),
.B1(n_61),
.B2(n_62),
.Y(n_65)
);

INVx8_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

OAI21xp33_ASAP7_75t_L g185 ( 
.A1(n_22),
.A2(n_39),
.B(n_61),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_23),
.B(n_172),
.Y(n_171)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_24),
.B(n_32),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_SL g72 ( 
.A(n_24),
.B(n_33),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_24),
.B(n_100),
.Y(n_99)
);

AOI21xp5_ASAP7_75t_L g148 ( 
.A1(n_24),
.A2(n_31),
.B(n_100),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_26),
.B1(n_27),
.B2(n_29),
.Y(n_24)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_25),
.Y(n_29)
);

AOI22xp33_ASAP7_75t_L g50 ( 
.A1(n_26),
.A2(n_27),
.B1(n_42),
.B2(n_43),
.Y(n_50)
);

OAI21xp33_ASAP7_75t_L g211 ( 
.A1(n_26),
.A2(n_29),
.B(n_39),
.Y(n_211)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_27),
.B(n_228),
.Y(n_227)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_30),
.B(n_99),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g169 ( 
.A(n_30),
.B(n_170),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_SL g30 ( 
.A(n_31),
.B(n_33),
.Y(n_30)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_31),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g178 ( 
.A(n_31),
.B(n_179),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_36),
.B(n_47),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_36),
.B(n_213),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_SL g36 ( 
.A(n_37),
.B(n_40),
.Y(n_36)
);

AOI21xp5_ASAP7_75t_SL g74 ( 
.A1(n_37),
.A2(n_40),
.B(n_75),
.Y(n_74)
);

CKINVDCx16_ASAP7_75t_R g37 ( 
.A(n_38),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_38),
.B(n_49),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_L g122 ( 
.A1(n_40),
.A2(n_48),
.B(n_86),
.Y(n_122)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_41),
.B(n_50),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_41),
.B(n_51),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_41),
.B(n_215),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g41 ( 
.A1(n_42),
.A2(n_43),
.B1(n_44),
.B2(n_46),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx6_ASAP7_75t_SL g46 ( 
.A(n_44),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_44),
.B(n_81),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_44),
.B(n_251),
.Y(n_250)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVxp33_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_48),
.B(n_225),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_49),
.B(n_51),
.Y(n_48)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_49),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_49),
.B(n_215),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_L g52 ( 
.A1(n_53),
.A2(n_68),
.B1(n_76),
.B2(n_77),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_53),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_53),
.A2(n_76),
.B1(n_95),
.B2(n_107),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_53),
.B(n_70),
.C(n_73),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_54),
.B(n_66),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_54),
.B(n_150),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_55),
.B(n_58),
.Y(n_54)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_55),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_55),
.B(n_65),
.Y(n_126)
);

INVx11_ASAP7_75t_L g104 ( 
.A(n_56),
.Y(n_104)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx11_ASAP7_75t_L g60 ( 
.A(n_57),
.Y(n_60)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_57),
.Y(n_64)
);

INVx6_ASAP7_75t_L g187 ( 
.A(n_57),
.Y(n_187)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_58),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_58),
.B(n_67),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_58),
.B(n_128),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_59),
.B(n_65),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_L g59 ( 
.A1(n_60),
.A2(n_61),
.B1(n_62),
.B2(n_63),
.Y(n_59)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_65),
.B(n_67),
.Y(n_66)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_65),
.Y(n_91)
);

AOI21xp5_ASAP7_75t_L g102 ( 
.A1(n_65),
.A2(n_103),
.B(n_105),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_65),
.B(n_128),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_66),
.B(n_127),
.Y(n_180)
);

CKINVDCx16_ASAP7_75t_R g77 ( 
.A(n_68),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_69),
.A2(n_70),
.B1(n_73),
.B2(n_74),
.Y(n_68)
);

CKINVDCx16_ASAP7_75t_R g69 ( 
.A(n_70),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_71),
.B(n_101),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_72),
.B(n_132),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_72),
.B(n_178),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_73),
.A2(n_74),
.B1(n_97),
.B2(n_98),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_73),
.B(n_167),
.C(n_169),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_73),
.A2(n_74),
.B1(n_169),
.B2(n_196),
.Y(n_195)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

OAI21xp5_ASAP7_75t_SL g85 ( 
.A1(n_75),
.A2(n_86),
.B(n_87),
.Y(n_85)
);

AOI21xp33_ASAP7_75t_L g78 ( 
.A1(n_79),
.A2(n_84),
.B(n_88),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_79),
.B(n_85),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_79),
.A2(n_85),
.B1(n_135),
.B2(n_136),
.Y(n_134)
);

CKINVDCx16_ASAP7_75t_R g136 ( 
.A(n_79),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_79),
.A2(n_88),
.B1(n_89),
.B2(n_136),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_79),
.B(n_210),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_L g266 ( 
.A1(n_79),
.A2(n_136),
.B1(n_210),
.B2(n_267),
.Y(n_266)
);

AOI21xp5_ASAP7_75t_L g79 ( 
.A1(n_80),
.A2(n_82),
.B(n_83),
.Y(n_79)
);

OR2x2_ASAP7_75t_L g120 ( 
.A(n_80),
.B(n_121),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_SL g140 ( 
.A1(n_80),
.A2(n_141),
.B(n_142),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g202 ( 
.A(n_80),
.B(n_83),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_SL g238 ( 
.A(n_80),
.B(n_239),
.Y(n_238)
);

BUFx2_ASAP7_75t_L g189 ( 
.A(n_81),
.Y(n_189)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_82),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_83),
.Y(n_119)
);

XOR2xp5_ASAP7_75t_L g154 ( 
.A(n_84),
.B(n_155),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_85),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_87),
.B(n_147),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_87),
.B(n_214),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_89),
.Y(n_88)
);

AOI21xp5_ASAP7_75t_SL g89 ( 
.A1(n_90),
.A2(n_91),
.B(n_92),
.Y(n_89)
);

XNOR2xp5_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_108),
.Y(n_93)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_95),
.Y(n_107)
);

XNOR2xp5_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_102),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_98),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g177 ( 
.A(n_99),
.B(n_178),
.Y(n_177)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

CKINVDCx14_ASAP7_75t_R g105 ( 
.A(n_106),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_106),
.B(n_150),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_SL g110 ( 
.A1(n_111),
.A2(n_296),
.B(n_299),
.Y(n_110)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_L g112 ( 
.A1(n_113),
.A2(n_159),
.B(n_295),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_151),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g295 ( 
.A(n_114),
.B(n_151),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_134),
.C(n_137),
.Y(n_114)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_115),
.B(n_134),
.Y(n_293)
);

XOR2xp5_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_123),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_116),
.B(n_124),
.C(n_131),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_122),
.Y(n_116)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_117),
.B(n_122),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_118),
.B(n_120),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_118),
.B(n_237),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_L g188 ( 
.A1(n_120),
.A2(n_141),
.B(n_189),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_120),
.B(n_245),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_121),
.B(n_144),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_124),
.A2(n_125),
.B1(n_130),
.B2(n_131),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_125),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_127),
.Y(n_125)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

CKINVDCx14_ASAP7_75t_R g132 ( 
.A(n_133),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_133),
.B(n_171),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g292 ( 
.A(n_137),
.B(n_293),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_148),
.C(n_149),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_138),
.A2(n_139),
.B1(n_282),
.B2(n_283),
.Y(n_281)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_146),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_140),
.B(n_146),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_143),
.B(n_202),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_143),
.B(n_238),
.Y(n_256)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_147),
.B(n_225),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_148),
.A2(n_149),
.B1(n_284),
.B2(n_285),
.Y(n_283)
);

CKINVDCx14_ASAP7_75t_R g284 ( 
.A(n_148),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_149),
.Y(n_285)
);

XOR2xp5_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_158),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_153),
.A2(n_154),
.B1(n_156),
.B2(n_157),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_153),
.B(n_157),
.C(n_158),
.Y(n_298)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_157),
.Y(n_156)
);

AOI21xp5_ASAP7_75t_L g159 ( 
.A1(n_160),
.A2(n_290),
.B(n_294),
.Y(n_159)
);

A2O1A1Ixp33_ASAP7_75t_SL g160 ( 
.A1(n_161),
.A2(n_203),
.B(n_276),
.C(n_289),
.Y(n_160)
);

OR2x2_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_191),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_162),
.B(n_191),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_163),
.A2(n_164),
.B1(n_175),
.B2(n_190),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_165),
.A2(n_166),
.B1(n_173),
.B2(n_174),
.Y(n_164)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_165),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_165),
.B(n_174),
.C(n_190),
.Y(n_277)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_166),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_167),
.A2(n_168),
.B1(n_194),
.B2(n_195),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_168),
.Y(n_167)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_169),
.Y(n_196)
);

CKINVDCx16_ASAP7_75t_R g170 ( 
.A(n_171),
.Y(n_170)
);

INVxp67_ASAP7_75t_SL g179 ( 
.A(n_172),
.Y(n_179)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_175),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_183),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_177),
.A2(n_180),
.B1(n_181),
.B2(n_182),
.Y(n_176)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_177),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_177),
.B(n_182),
.C(n_183),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_180),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_188),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_184),
.B(n_188),
.Y(n_197)
);

INVx8_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_197),
.C(n_198),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_192),
.A2(n_193),
.B1(n_217),
.B2(n_218),
.Y(n_216)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_197),
.B(n_198),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_200),
.C(n_201),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_199),
.B(n_208),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_200),
.B(n_201),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_202),
.B(n_253),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_204),
.B(n_275),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_L g204 ( 
.A1(n_205),
.A2(n_219),
.B(n_274),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_216),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_206),
.B(n_216),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_209),
.C(n_212),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_207),
.B(n_272),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_209),
.B(n_212),
.Y(n_272)
);

CKINVDCx16_ASAP7_75t_R g267 ( 
.A(n_210),
.Y(n_267)
);

INVxp33_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

AOI21xp5_ASAP7_75t_L g219 ( 
.A1(n_220),
.A2(n_269),
.B(n_273),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_SL g220 ( 
.A1(n_221),
.A2(n_260),
.B(n_268),
.Y(n_220)
);

AOI21xp5_ASAP7_75t_L g221 ( 
.A1(n_222),
.A2(n_242),
.B(n_259),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_229),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_SL g259 ( 
.A(n_223),
.B(n_229),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_224),
.B(n_226),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_224),
.A2(n_226),
.B1(n_227),
.B2(n_247),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_224),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_227),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_230),
.A2(n_231),
.B1(n_236),
.B2(n_241),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_232),
.A2(n_233),
.B1(n_234),
.B2(n_235),
.Y(n_231)
);

CKINVDCx14_ASAP7_75t_R g234 ( 
.A(n_232),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_232),
.B(n_235),
.C(n_241),
.Y(n_261)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_233),
.Y(n_235)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_236),
.Y(n_241)
);

INVxp67_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

CKINVDCx16_ASAP7_75t_R g239 ( 
.A(n_240),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_SL g242 ( 
.A1(n_243),
.A2(n_248),
.B(n_258),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_246),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_244),
.B(n_246),
.Y(n_258)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_245),
.Y(n_253)
);

AOI21xp5_ASAP7_75t_L g248 ( 
.A1(n_249),
.A2(n_254),
.B(n_257),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_252),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_256),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_SL g257 ( 
.A(n_255),
.B(n_256),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_262),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_SL g268 ( 
.A(n_261),
.B(n_262),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_263),
.B(n_266),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_264),
.B(n_265),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_264),
.B(n_265),
.C(n_266),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_270),
.B(n_271),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_SL g273 ( 
.A(n_270),
.B(n_271),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_278),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g289 ( 
.A(n_277),
.B(n_278),
.Y(n_289)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_279),
.B(n_288),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_280),
.A2(n_281),
.B1(n_286),
.B2(n_287),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_280),
.B(n_287),
.C(n_288),
.Y(n_291)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

CKINVDCx16_ASAP7_75t_R g286 ( 
.A(n_287),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_291),
.B(n_292),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_SL g294 ( 
.A(n_291),
.B(n_292),
.Y(n_294)
);

INVxp67_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);


endmodule