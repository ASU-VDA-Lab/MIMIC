module fake_jpeg_15950_n_275 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_275);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_275;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_228;
wire n_178;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_223;
wire n_187;
wire n_21;
wire n_57;
wire n_175;
wire n_234;
wire n_272;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_139;
wire n_45;
wire n_61;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_140;
wire n_82;
wire n_128;
wire n_100;
wire n_258;
wire n_96;

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_13),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

INVx5_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

INVx1_ASAP7_75t_SL g22 ( 
.A(n_6),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

INVx8_ASAP7_75t_SL g24 ( 
.A(n_7),
.Y(n_24)
);

INVx11_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_14),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

BUFx16f_ASAP7_75t_L g34 ( 
.A(n_26),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_26),
.Y(n_35)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_35),
.Y(n_53)
);

INVx13_ASAP7_75t_L g36 ( 
.A(n_24),
.Y(n_36)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_36),
.Y(n_43)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g38 ( 
.A1(n_21),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_38),
.A2(n_22),
.B1(n_25),
.B2(n_21),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_22),
.B(n_8),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_39),
.B(n_20),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_17),
.Y(n_40)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_26),
.Y(n_41)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g42 ( 
.A(n_39),
.B(n_31),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_42),
.B(n_51),
.Y(n_71)
);

AND2x2_ASAP7_75t_SL g44 ( 
.A(n_34),
.B(n_26),
.Y(n_44)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_44),
.B(n_46),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_39),
.B(n_31),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_L g47 ( 
.A1(n_36),
.A2(n_30),
.B1(n_21),
.B2(n_22),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_47),
.A2(n_41),
.B1(n_34),
.B2(n_17),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_48),
.A2(n_30),
.B1(n_36),
.B2(n_38),
.Y(n_73)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_34),
.Y(n_49)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_49),
.Y(n_61)
);

AOI21xp33_ASAP7_75t_SL g50 ( 
.A1(n_34),
.A2(n_24),
.B(n_32),
.Y(n_50)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_50),
.B(n_54),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_40),
.Y(n_51)
);

MAJIxp5_ASAP7_75t_L g54 ( 
.A(n_35),
.B(n_32),
.C(n_18),
.Y(n_54)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_55),
.Y(n_83)
);

OAI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_36),
.A2(n_25),
.B1(n_19),
.B2(n_29),
.Y(n_56)
);

OAI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_56),
.A2(n_17),
.B1(n_33),
.B2(n_27),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g57 ( 
.A(n_34),
.B(n_0),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_57),
.B(n_60),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_58),
.Y(n_62)
);

INVx11_ASAP7_75t_L g115 ( 
.A(n_62),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_42),
.B(n_60),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_63),
.B(n_74),
.Y(n_96)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_58),
.Y(n_64)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_64),
.Y(n_97)
);

BUFx24_ASAP7_75t_L g65 ( 
.A(n_43),
.Y(n_65)
);

INVx13_ASAP7_75t_L g93 ( 
.A(n_65),
.Y(n_93)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_53),
.Y(n_68)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_68),
.Y(n_105)
);

OR2x2_ASAP7_75t_L g69 ( 
.A(n_46),
.B(n_36),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_69),
.B(n_70),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_57),
.B(n_37),
.Y(n_70)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_53),
.Y(n_72)
);

INVxp67_ASAP7_75t_SL g100 ( 
.A(n_72),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_73),
.A2(n_40),
.B1(n_23),
.B2(n_27),
.Y(n_102)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_59),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_59),
.B(n_29),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_75),
.B(n_77),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_L g76 ( 
.A1(n_48),
.A2(n_25),
.B1(n_41),
.B2(n_19),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_76),
.A2(n_85),
.B1(n_55),
.B2(n_52),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_43),
.B(n_20),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_44),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_78),
.B(n_82),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_50),
.A2(n_38),
.B1(n_41),
.B2(n_37),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_79),
.A2(n_81),
.B1(n_86),
.B2(n_55),
.Y(n_94)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_57),
.Y(n_80)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_80),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_43),
.A2(n_41),
.B1(n_37),
.B2(n_34),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_57),
.B(n_32),
.Y(n_82)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_52),
.Y(n_84)
);

INVx13_ASAP7_75t_L g104 ( 
.A(n_84),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_52),
.A2(n_17),
.B1(n_33),
.B2(n_23),
.Y(n_86)
);

OAI21xp33_ASAP7_75t_SL g112 ( 
.A1(n_87),
.A2(n_18),
.B(n_32),
.Y(n_112)
);

BUFx12f_ASAP7_75t_L g89 ( 
.A(n_45),
.Y(n_89)
);

INVx6_ASAP7_75t_SL g90 ( 
.A(n_89),
.Y(n_90)
);

OA22x2_ASAP7_75t_L g91 ( 
.A1(n_78),
.A2(n_51),
.B1(n_44),
.B2(n_40),
.Y(n_91)
);

AO22x1_ASAP7_75t_L g135 ( 
.A1(n_91),
.A2(n_84),
.B1(n_62),
.B2(n_64),
.Y(n_135)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_94),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_SL g98 ( 
.A1(n_88),
.A2(n_44),
.B(n_54),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_98),
.B(n_99),
.C(n_109),
.Y(n_142)
);

AND2x2_ASAP7_75t_SL g99 ( 
.A(n_70),
.B(n_45),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_101),
.A2(n_102),
.B1(n_106),
.B2(n_112),
.Y(n_118)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_82),
.B(n_0),
.Y(n_103)
);

XNOR2x1_ASAP7_75t_L g127 ( 
.A(n_103),
.B(n_69),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_73),
.A2(n_23),
.B1(n_27),
.B2(n_33),
.Y(n_106)
);

AOI21xp5_ASAP7_75t_L g107 ( 
.A1(n_88),
.A2(n_32),
.B(n_1),
.Y(n_107)
);

CKINVDCx16_ASAP7_75t_R g122 ( 
.A(n_107),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_67),
.B(n_49),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_108),
.B(n_111),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_80),
.B(n_35),
.C(n_45),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_67),
.B(n_49),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_67),
.B(n_35),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_113),
.B(n_69),
.Y(n_124)
);

OAI211xp5_ASAP7_75t_L g116 ( 
.A1(n_66),
.A2(n_35),
.B(n_18),
.C(n_28),
.Y(n_116)
);

A2O1A1O1Ixp25_ASAP7_75t_L g133 ( 
.A1(n_116),
.A2(n_85),
.B(n_28),
.C(n_62),
.D(n_65),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_97),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_119),
.B(n_125),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_L g120 ( 
.A(n_98),
.B(n_66),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_120),
.B(n_121),
.C(n_140),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g121 ( 
.A(n_113),
.B(n_88),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_110),
.B(n_72),
.Y(n_123)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_123),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_SL g145 ( 
.A1(n_124),
.A2(n_126),
.B(n_107),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_97),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_96),
.Y(n_126)
);

OAI21xp33_ASAP7_75t_SL g149 ( 
.A1(n_127),
.A2(n_133),
.B(n_116),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_92),
.B(n_71),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_128),
.B(n_138),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_110),
.B(n_74),
.Y(n_129)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_129),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_96),
.B(n_114),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g166 ( 
.A(n_130),
.B(n_144),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_90),
.B(n_68),
.Y(n_131)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_131),
.Y(n_164)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_105),
.Y(n_134)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_134),
.Y(n_157)
);

OA21x2_ASAP7_75t_L g153 ( 
.A1(n_135),
.A2(n_112),
.B(n_91),
.Y(n_153)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_105),
.Y(n_136)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_136),
.Y(n_171)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_91),
.Y(n_137)
);

CKINVDCx16_ASAP7_75t_R g172 ( 
.A(n_137),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_92),
.B(n_65),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_91),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_139),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_SL g140 ( 
.A(n_108),
.B(n_11),
.Y(n_140)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_104),
.Y(n_141)
);

INVx3_ASAP7_75t_L g156 ( 
.A(n_141),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_111),
.B(n_61),
.C(n_65),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_143),
.B(n_99),
.C(n_95),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_103),
.B(n_61),
.Y(n_144)
);

CKINVDCx14_ASAP7_75t_R g177 ( 
.A(n_145),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_141),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g197 ( 
.A(n_148),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_149),
.A2(n_150),
.B1(n_132),
.B2(n_133),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_118),
.A2(n_101),
.B1(n_114),
.B2(n_106),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_137),
.A2(n_95),
.B1(n_91),
.B2(n_109),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_151),
.A2(n_168),
.B1(n_117),
.B2(n_138),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_152),
.B(n_154),
.C(n_160),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_L g181 ( 
.A1(n_153),
.A2(n_163),
.B(n_132),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_142),
.B(n_99),
.C(n_102),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_142),
.B(n_99),
.C(n_103),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_128),
.B(n_103),
.Y(n_161)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_161),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_121),
.B(n_89),
.C(n_83),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_162),
.B(n_165),
.C(n_169),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_L g163 ( 
.A1(n_139),
.A2(n_100),
.B(n_28),
.Y(n_163)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_120),
.B(n_100),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_118),
.A2(n_115),
.B1(n_104),
.B2(n_93),
.Y(n_168)
);

MAJx2_ASAP7_75t_L g169 ( 
.A(n_127),
.B(n_90),
.C(n_104),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_117),
.B(n_93),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_170),
.B(n_173),
.Y(n_178)
);

NOR3xp33_ASAP7_75t_L g173 ( 
.A(n_126),
.B(n_11),
.C(n_15),
.Y(n_173)
);

CKINVDCx16_ASAP7_75t_R g174 ( 
.A(n_155),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_174),
.B(n_188),
.Y(n_201)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_157),
.Y(n_176)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_176),
.Y(n_198)
);

CKINVDCx14_ASAP7_75t_R g209 ( 
.A(n_179),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_156),
.B(n_135),
.Y(n_180)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_180),
.Y(n_207)
);

XOR2x1_ASAP7_75t_L g205 ( 
.A(n_181),
.B(n_195),
.Y(n_205)
);

A2O1A1Ixp33_ASAP7_75t_L g182 ( 
.A1(n_145),
.A2(n_122),
.B(n_124),
.C(n_135),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_182),
.B(n_151),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_156),
.B(n_143),
.Y(n_183)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_183),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_184),
.B(n_193),
.Y(n_213)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_157),
.Y(n_185)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_185),
.Y(n_206)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_171),
.Y(n_186)
);

CKINVDCx16_ASAP7_75t_R g199 ( 
.A(n_186),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_SL g187 ( 
.A(n_166),
.B(n_140),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_SL g215 ( 
.A(n_187),
.B(n_196),
.Y(n_215)
);

INVxp67_ASAP7_75t_L g188 ( 
.A(n_168),
.Y(n_188)
);

INVx13_ASAP7_75t_L g189 ( 
.A(n_148),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_189),
.B(n_194),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_172),
.A2(n_167),
.B1(n_154),
.B2(n_159),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_190),
.A2(n_152),
.B1(n_160),
.B2(n_159),
.Y(n_208)
);

AOI21xp5_ASAP7_75t_L g193 ( 
.A1(n_163),
.A2(n_89),
.B(n_136),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_158),
.Y(n_194)
);

AND2x4_ASAP7_75t_L g195 ( 
.A(n_169),
.B(n_134),
.Y(n_195)
);

BUFx2_ASAP7_75t_L g196 ( 
.A(n_164),
.Y(n_196)
);

BUFx24_ASAP7_75t_SL g200 ( 
.A(n_194),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_200),
.B(n_187),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g202 ( 
.A(n_192),
.B(n_165),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_202),
.B(n_204),
.C(n_191),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_192),
.B(n_147),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g223 ( 
.A1(n_208),
.A2(n_214),
.B1(n_216),
.B2(n_195),
.Y(n_223)
);

NOR2xp67_ASAP7_75t_SL g210 ( 
.A(n_195),
.B(n_162),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_SL g230 ( 
.A1(n_210),
.A2(n_185),
.B(n_186),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_SL g221 ( 
.A(n_212),
.B(n_179),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_188),
.A2(n_153),
.B1(n_146),
.B2(n_161),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_177),
.A2(n_153),
.B1(n_170),
.B2(n_147),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_176),
.B(n_115),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_217),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_217),
.Y(n_219)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_219),
.Y(n_239)
);

HB1xp67_ASAP7_75t_L g220 ( 
.A(n_199),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_220),
.B(n_224),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_SL g237 ( 
.A(n_221),
.B(n_230),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_216),
.B(n_191),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_222),
.B(n_223),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_205),
.A2(n_195),
.B1(n_181),
.B2(n_184),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_225),
.A2(n_213),
.B1(n_207),
.B2(n_206),
.Y(n_233)
);

AOI21xp5_ASAP7_75t_L g226 ( 
.A1(n_205),
.A2(n_182),
.B(n_193),
.Y(n_226)
);

AOI22xp33_ASAP7_75t_SL g242 ( 
.A1(n_226),
.A2(n_197),
.B1(n_89),
.B2(n_93),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_SL g235 ( 
.A(n_227),
.B(n_228),
.Y(n_235)
);

AOI322xp5_ASAP7_75t_L g228 ( 
.A1(n_215),
.A2(n_209),
.A3(n_212),
.B1(n_201),
.B2(n_211),
.C1(n_178),
.C2(n_175),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_202),
.B(n_190),
.C(n_175),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_229),
.B(n_231),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_208),
.B(n_213),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_L g232 ( 
.A1(n_214),
.A2(n_196),
.B1(n_115),
.B2(n_197),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_232),
.A2(n_206),
.B1(n_198),
.B2(n_203),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_233),
.B(n_10),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_L g246 ( 
.A1(n_234),
.A2(n_236),
.B1(n_242),
.B2(n_243),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_218),
.A2(n_196),
.B1(n_189),
.B2(n_204),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_231),
.B(n_197),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_240),
.B(n_229),
.C(n_230),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_221),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_245),
.B(n_248),
.C(n_238),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_239),
.B(n_226),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g255 ( 
.A(n_247),
.B(n_250),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_241),
.B(n_224),
.C(n_222),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_SL g249 ( 
.A1(n_242),
.A2(n_225),
.B(n_10),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_249),
.B(n_251),
.Y(n_261)
);

OAI21xp5_ASAP7_75t_SL g251 ( 
.A1(n_235),
.A2(n_9),
.B(n_16),
.Y(n_251)
);

NOR2xp67_ASAP7_75t_L g252 ( 
.A(n_237),
.B(n_11),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_SL g257 ( 
.A(n_252),
.B(n_253),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_237),
.A2(n_240),
.B1(n_244),
.B2(n_238),
.Y(n_253)
);

NOR2x1_ASAP7_75t_SL g254 ( 
.A(n_244),
.B(n_6),
.Y(n_254)
);

AO21x1_ASAP7_75t_L g256 ( 
.A1(n_254),
.A2(n_12),
.B(n_16),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_256),
.B(n_258),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_253),
.B(n_83),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_SL g264 ( 
.A(n_259),
.B(n_260),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_248),
.B(n_5),
.Y(n_260)
);

OAI21xp5_ASAP7_75t_SL g263 ( 
.A1(n_257),
.A2(n_245),
.B(n_246),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_263),
.B(n_265),
.Y(n_270)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_255),
.Y(n_265)
);

AOI221xp5_ASAP7_75t_L g266 ( 
.A1(n_261),
.A2(n_5),
.B1(n_15),
.B2(n_3),
.C(n_4),
.Y(n_266)
);

AOI322xp5_ASAP7_75t_L g268 ( 
.A1(n_266),
.A2(n_256),
.A3(n_12),
.B1(n_3),
.B2(n_4),
.C1(n_5),
.C2(n_16),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_262),
.B(n_264),
.Y(n_267)
);

OAI21xp5_ASAP7_75t_L g271 ( 
.A1(n_267),
.A2(n_268),
.B(n_269),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g269 ( 
.A(n_262),
.B(n_258),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_L g272 ( 
.A1(n_270),
.A2(n_3),
.B(n_13),
.Y(n_272)
);

OAI21xp5_ASAP7_75t_L g273 ( 
.A1(n_272),
.A2(n_1),
.B(n_2),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_273),
.B(n_271),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_274),
.B(n_13),
.Y(n_275)
);


endmodule