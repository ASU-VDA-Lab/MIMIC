module fake_jpeg_17011_n_62 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_62);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_62;

wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_23;
wire n_27;
wire n_55;
wire n_22;
wire n_51;
wire n_47;
wire n_40;
wire n_19;
wire n_20;
wire n_18;
wire n_59;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_31;
wire n_25;
wire n_56;
wire n_37;
wire n_29;
wire n_50;
wire n_43;
wire n_32;

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_1),
.B(n_0),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_0),
.B(n_3),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_16),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_15),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_13),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_12),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_14),
.Y(n_29)
);

BUFx8_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_17),
.B(n_7),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

INVx5_ASAP7_75t_L g34 ( 
.A(n_32),
.Y(n_34)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_34),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g35 ( 
.A(n_27),
.B(n_8),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_35),
.B(n_36),
.Y(n_47)
);

INVx13_ASAP7_75t_L g36 ( 
.A(n_30),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_32),
.Y(n_37)
);

CKINVDCx6p67_ASAP7_75t_R g50 ( 
.A(n_37),
.Y(n_50)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_30),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_38),
.A2(n_39),
.B1(n_40),
.B2(n_41),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g39 ( 
.A1(n_21),
.A2(n_24),
.B1(n_22),
.B2(n_23),
.Y(n_39)
);

NAND3xp33_ASAP7_75t_L g40 ( 
.A(n_19),
.B(n_20),
.C(n_31),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_18),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_25),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_29),
.B(n_26),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_28),
.B(n_19),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_19),
.B(n_26),
.Y(n_46)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_50),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_51),
.B(n_52),
.Y(n_53)
);

INVxp67_ASAP7_75t_L g52 ( 
.A(n_50),
.Y(n_52)
);

MAJIxp5_ASAP7_75t_SL g54 ( 
.A(n_52),
.B(n_47),
.C(n_45),
.Y(n_54)
);

AOI21xp5_ASAP7_75t_L g55 ( 
.A1(n_54),
.A2(n_46),
.B(n_49),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_55),
.Y(n_56)
);

AOI21xp33_ASAP7_75t_L g57 ( 
.A1(n_56),
.A2(n_53),
.B(n_48),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_57),
.B(n_58),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_56),
.Y(n_58)
);

AO21x1_ASAP7_75t_L g60 ( 
.A1(n_59),
.A2(n_44),
.B(n_42),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_60),
.Y(n_61)
);

XNOR2xp5_ASAP7_75t_L g62 ( 
.A(n_61),
.B(n_43),
.Y(n_62)
);


endmodule