module fake_jpeg_21132_n_284 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_284);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_284;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_265;
wire n_272;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_273;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

INVx8_ASAP7_75t_L g19 ( 
.A(n_17),
.Y(n_19)
);

INVx11_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

BUFx10_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_14),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_16),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_5),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_16),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_2),
.B(n_12),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

BUFx12_ASAP7_75t_L g35 ( 
.A(n_5),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_11),
.Y(n_36)
);

BUFx4f_ASAP7_75t_SL g37 ( 
.A(n_12),
.Y(n_37)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_8),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_15),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_1),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_6),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_2),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_13),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_32),
.B(n_18),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_44),
.B(n_45),
.Y(n_68)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_27),
.Y(n_45)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_27),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_46),
.B(n_53),
.Y(n_82)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_27),
.Y(n_47)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_47),
.Y(n_73)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_29),
.Y(n_48)
);

INVx6_ASAP7_75t_L g90 ( 
.A(n_48),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_29),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_49),
.Y(n_81)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_29),
.Y(n_50)
);

NAND2xp33_ASAP7_75t_SL g93 ( 
.A(n_50),
.B(n_65),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_31),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_51),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_31),
.Y(n_52)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_52),
.Y(n_78)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_34),
.Y(n_53)
);

INVx4_ASAP7_75t_SL g54 ( 
.A(n_31),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_54),
.B(n_56),
.Y(n_91)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_34),
.Y(n_55)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_55),
.Y(n_80)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_33),
.Y(n_56)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_33),
.Y(n_57)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_57),
.Y(n_88)
);

NOR2xp67_ASAP7_75t_R g58 ( 
.A(n_35),
.B(n_0),
.Y(n_58)
);

HAxp5_ASAP7_75t_SL g83 ( 
.A(n_58),
.B(n_35),
.CON(n_83),
.SN(n_83)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_33),
.Y(n_59)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_59),
.Y(n_70)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_34),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_60),
.B(n_63),
.Y(n_79)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_39),
.Y(n_61)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_61),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_62),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_32),
.B(n_18),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_39),
.Y(n_64)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_64),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_26),
.Y(n_65)
);

INVx2_ASAP7_75t_SL g66 ( 
.A(n_35),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_66),
.B(n_67),
.Y(n_84)
);

INVx4_ASAP7_75t_SL g67 ( 
.A(n_35),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_57),
.A2(n_28),
.B1(n_26),
.B2(n_19),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_69),
.A2(n_92),
.B1(n_47),
.B2(n_22),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_56),
.A2(n_28),
.B1(n_19),
.B2(n_20),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_71),
.A2(n_72),
.B1(n_37),
.B2(n_61),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_48),
.A2(n_19),
.B1(n_38),
.B2(n_20),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_66),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_75),
.B(n_85),
.Y(n_101)
);

BUFx8_ASAP7_75t_L g77 ( 
.A(n_67),
.Y(n_77)
);

INVx1_ASAP7_75t_SL g110 ( 
.A(n_77),
.Y(n_110)
);

OR2x2_ASAP7_75t_SL g129 ( 
.A(n_83),
.B(n_37),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_53),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_65),
.B(n_21),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_89),
.B(n_52),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_50),
.A2(n_20),
.B1(n_38),
.B2(n_25),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_94),
.B(n_118),
.Y(n_136)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_81),
.Y(n_95)
);

INVx4_ASAP7_75t_L g139 ( 
.A(n_95),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_68),
.B(n_24),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_96),
.B(n_97),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_68),
.B(n_24),
.Y(n_97)
);

BUFx3_ASAP7_75t_L g98 ( 
.A(n_73),
.Y(n_98)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_98),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_79),
.B(n_23),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_99),
.B(n_100),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_84),
.B(n_23),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_75),
.B(n_30),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_102),
.B(n_104),
.Y(n_155)
);

BUFx4f_ASAP7_75t_L g103 ( 
.A(n_81),
.Y(n_103)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_103),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_82),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_90),
.A2(n_38),
.B1(n_54),
.B2(n_55),
.Y(n_105)
);

INVxp67_ASAP7_75t_L g153 ( 
.A(n_105),
.Y(n_153)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_70),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_106),
.Y(n_131)
);

OR2x2_ASAP7_75t_L g107 ( 
.A(n_82),
.B(n_25),
.Y(n_107)
);

OR2x2_ASAP7_75t_L g132 ( 
.A(n_107),
.B(n_116),
.Y(n_132)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_81),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_108),
.B(n_109),
.Y(n_143)
);

CKINVDCx16_ASAP7_75t_R g109 ( 
.A(n_91),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_91),
.Y(n_111)
);

INVx5_ASAP7_75t_L g140 ( 
.A(n_111),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_85),
.B(n_30),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_112),
.B(n_114),
.Y(n_152)
);

AND2x2_ASAP7_75t_L g154 ( 
.A(n_113),
.B(n_117),
.Y(n_154)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_87),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_90),
.A2(n_40),
.B1(n_36),
.B2(n_43),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_115),
.A2(n_121),
.B1(n_86),
.B2(n_78),
.Y(n_142)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_87),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_70),
.Y(n_117)
);

INVx4_ASAP7_75t_L g118 ( 
.A(n_73),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_77),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_119),
.B(n_120),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_76),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_89),
.A2(n_59),
.B1(n_51),
.B2(n_49),
.Y(n_121)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_87),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_122),
.B(n_124),
.Y(n_149)
);

NAND2xp33_ASAP7_75t_SL g123 ( 
.A(n_93),
.B(n_64),
.Y(n_123)
);

AOI32xp33_ASAP7_75t_L g137 ( 
.A1(n_123),
.A2(n_88),
.A3(n_86),
.B1(n_76),
.B2(n_74),
.Y(n_137)
);

OR2x2_ASAP7_75t_L g124 ( 
.A(n_80),
.B(n_35),
.Y(n_124)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_77),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_125),
.B(n_126),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_80),
.B(n_37),
.Y(n_126)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_77),
.Y(n_127)
);

A2O1A1Ixp33_ASAP7_75t_L g135 ( 
.A1(n_127),
.A2(n_129),
.B(n_78),
.C(n_37),
.Y(n_135)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_90),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_128),
.A2(n_130),
.B1(n_74),
.B2(n_41),
.Y(n_144)
);

AO22x1_ASAP7_75t_SL g134 ( 
.A1(n_123),
.A2(n_93),
.B1(n_88),
.B2(n_69),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_134),
.B(n_121),
.Y(n_162)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_135),
.B(n_111),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_137),
.B(n_129),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_142),
.A2(n_144),
.B1(n_147),
.B2(n_148),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_94),
.A2(n_92),
.B1(n_62),
.B2(n_43),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_104),
.A2(n_41),
.B1(n_40),
.B2(n_36),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_113),
.A2(n_42),
.B1(n_22),
.B2(n_21),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_151),
.A2(n_120),
.B1(n_108),
.B2(n_114),
.Y(n_168)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_139),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g175 ( 
.A(n_156),
.Y(n_175)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_146),
.Y(n_157)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_157),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_155),
.B(n_101),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_158),
.B(n_159),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_136),
.B(n_101),
.C(n_124),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_160),
.B(n_132),
.C(n_149),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_141),
.B(n_102),
.Y(n_161)
);

CKINVDCx16_ASAP7_75t_R g185 ( 
.A(n_161),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_162),
.B(n_165),
.Y(n_176)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_139),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_163),
.B(n_171),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_152),
.B(n_107),
.Y(n_166)
);

INVxp67_ASAP7_75t_L g184 ( 
.A(n_166),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_140),
.Y(n_167)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_167),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_168),
.B(n_169),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_136),
.A2(n_106),
.B1(n_117),
.B2(n_128),
.Y(n_169)
);

INVx3_ASAP7_75t_L g170 ( 
.A(n_138),
.Y(n_170)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_170),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_SL g171 ( 
.A(n_155),
.B(n_42),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_140),
.B(n_125),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_172),
.B(n_173),
.Y(n_182)
);

BUFx12_ASAP7_75t_L g173 ( 
.A(n_138),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_146),
.Y(n_174)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_174),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_180),
.B(n_164),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_162),
.A2(n_153),
.B1(n_154),
.B2(n_134),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_181),
.A2(n_144),
.B1(n_147),
.B2(n_151),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_167),
.B(n_143),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_187),
.B(n_193),
.Y(n_197)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_169),
.Y(n_190)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_190),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_157),
.B(n_154),
.Y(n_191)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_191),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_174),
.B(n_149),
.C(n_150),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_192),
.B(n_132),
.C(n_148),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_160),
.B(n_154),
.Y(n_193)
);

AND2x6_ASAP7_75t_L g194 ( 
.A(n_165),
.B(n_137),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_194),
.B(n_164),
.Y(n_200)
);

HB1xp67_ASAP7_75t_L g195 ( 
.A(n_192),
.Y(n_195)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_195),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_SL g196 ( 
.A1(n_194),
.A2(n_176),
.B(n_153),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_SL g213 ( 
.A1(n_196),
.A2(n_200),
.B(n_210),
.Y(n_213)
);

NOR3xp33_ASAP7_75t_L g198 ( 
.A(n_184),
.B(n_171),
.C(n_131),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_198),
.B(n_205),
.Y(n_218)
);

CKINVDCx16_ASAP7_75t_R g199 ( 
.A(n_177),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_199),
.B(n_207),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_202),
.B(n_209),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_190),
.A2(n_134),
.B1(n_142),
.B2(n_168),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_204),
.A2(n_206),
.B1(n_131),
.B2(n_179),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_188),
.A2(n_176),
.B1(n_189),
.B2(n_178),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_182),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_185),
.B(n_173),
.Y(n_208)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_208),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g209 ( 
.A(n_193),
.B(n_150),
.Y(n_209)
);

AOI21xp5_ASAP7_75t_L g210 ( 
.A1(n_181),
.A2(n_191),
.B(n_189),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_211),
.B(n_180),
.C(n_186),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_214),
.B(n_216),
.C(n_220),
.Y(n_237)
);

AND2x2_ASAP7_75t_L g215 ( 
.A(n_197),
.B(n_132),
.Y(n_215)
);

AOI21xp5_ASAP7_75t_L g231 ( 
.A1(n_215),
.A2(n_199),
.B(n_203),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_202),
.B(n_178),
.C(n_188),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_196),
.B(n_184),
.C(n_133),
.Y(n_220)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_221),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_209),
.B(n_170),
.C(n_173),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_222),
.B(n_175),
.C(n_118),
.Y(n_238)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_201),
.Y(n_223)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_223),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_SL g224 ( 
.A(n_211),
.B(n_135),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_224),
.B(n_210),
.Y(n_230)
);

HB1xp67_ASAP7_75t_L g227 ( 
.A(n_225),
.Y(n_227)
);

INVx1_ASAP7_75t_SL g241 ( 
.A(n_227),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_219),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_228),
.B(n_239),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_218),
.A2(n_204),
.B1(n_206),
.B2(n_207),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_L g246 ( 
.A1(n_229),
.A2(n_163),
.B1(n_156),
.B2(n_145),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_230),
.B(n_233),
.Y(n_245)
);

AOI21xp5_ASAP7_75t_SL g250 ( 
.A1(n_231),
.A2(n_175),
.B(n_98),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_212),
.B(n_205),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_212),
.B(n_203),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_234),
.B(n_235),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_SL g235 ( 
.A(n_214),
.B(n_201),
.Y(n_235)
);

OAI21xp5_ASAP7_75t_L g236 ( 
.A1(n_213),
.A2(n_179),
.B(n_173),
.Y(n_236)
);

AOI21xp5_ASAP7_75t_L g249 ( 
.A1(n_236),
.A2(n_119),
.B(n_127),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_238),
.B(n_234),
.C(n_237),
.Y(n_251)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_215),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_L g240 ( 
.A1(n_238),
.A2(n_217),
.B(n_216),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_240),
.B(n_246),
.C(n_248),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_226),
.A2(n_224),
.B1(n_183),
.B2(n_222),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_243),
.B(n_251),
.C(n_21),
.Y(n_260)
);

AOI21x1_ASAP7_75t_SL g244 ( 
.A1(n_232),
.A2(n_145),
.B(n_183),
.Y(n_244)
);

HB1xp67_ASAP7_75t_L g254 ( 
.A(n_244),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_L g248 ( 
.A1(n_237),
.A2(n_230),
.B1(n_233),
.B2(n_235),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_SL g253 ( 
.A1(n_249),
.A2(n_250),
.B(n_110),
.Y(n_253)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_253),
.Y(n_262)
);

MAJx2_ASAP7_75t_L g255 ( 
.A(n_251),
.B(n_17),
.C(n_15),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_255),
.B(n_260),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_247),
.B(n_175),
.C(n_103),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_256),
.B(n_257),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_247),
.B(n_245),
.C(n_242),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_245),
.B(n_103),
.C(n_21),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_258),
.B(n_259),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_244),
.B(n_21),
.C(n_14),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_252),
.B(n_241),
.Y(n_261)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_261),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_254),
.B(n_241),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_266),
.B(n_267),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_254),
.A2(n_250),
.B1(n_122),
.B2(n_116),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_264),
.B(n_95),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_268),
.B(n_273),
.Y(n_277)
);

CKINVDCx16_ASAP7_75t_R g269 ( 
.A(n_261),
.Y(n_269)
);

AOI21xp33_ASAP7_75t_L g274 ( 
.A1(n_269),
.A2(n_270),
.B(n_263),
.Y(n_274)
);

AOI322xp5_ASAP7_75t_L g270 ( 
.A1(n_262),
.A2(n_0),
.A3(n_1),
.B1(n_3),
.B2(n_4),
.C1(n_5),
.C2(n_6),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_265),
.B(n_0),
.Y(n_273)
);

OR2x2_ASAP7_75t_L g279 ( 
.A(n_274),
.B(n_268),
.Y(n_279)
);

AOI21xp5_ASAP7_75t_L g275 ( 
.A1(n_271),
.A2(n_1),
.B(n_7),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_275),
.B(n_276),
.C(n_273),
.Y(n_278)
);

OAI21xp5_ASAP7_75t_L g276 ( 
.A1(n_272),
.A2(n_7),
.B(n_8),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_SL g281 ( 
.A(n_278),
.B(n_279),
.Y(n_281)
);

AOI321xp33_ASAP7_75t_L g280 ( 
.A1(n_279),
.A2(n_277),
.A3(n_9),
.B1(n_10),
.B2(n_11),
.C(n_13),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_280),
.A2(n_110),
.B1(n_9),
.B2(n_10),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_SL g283 ( 
.A(n_282),
.B(n_281),
.Y(n_283)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_283),
.B(n_7),
.Y(n_284)
);


endmodule