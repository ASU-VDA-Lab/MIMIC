module real_jpeg_10607_n_11 (n_5, n_4, n_8, n_0, n_250, n_1, n_2, n_6, n_7, n_3, n_10, n_9, n_11);

input n_5;
input n_4;
input n_8;
input n_0;
input n_250;
input n_1;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_11;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_201;
wire n_114;
wire n_68;
wire n_247;
wire n_146;
wire n_78;
wire n_83;
wire n_215;
wire n_166;
wire n_221;
wire n_176;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_173;
wire n_105;
wire n_243;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_200;
wire n_48;
wire n_164;
wire n_184;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_13;
wire n_120;
wire n_155;
wire n_113;
wire n_199;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_188;
wire n_139;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_208;
wire n_62;
wire n_239;
wire n_162;
wire n_245;
wire n_121;
wire n_234;
wire n_106;
wire n_172;
wire n_211;
wire n_160;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_222;
wire n_148;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_195;
wire n_110;
wire n_205;
wire n_117;
wire n_193;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_228;
wire n_150;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_225;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_240;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_191;
wire n_52;
wire n_58;
wire n_63;
wire n_12;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_244;
wire n_167;
wire n_179;
wire n_202;
wire n_213;
wire n_133;
wire n_216;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_210;
wire n_127;
wire n_206;
wire n_224;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;
wire n_16;

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_0),
.A2(n_1),
.B1(n_22),
.B2(n_23),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_0),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_L g41 ( 
.A1(n_0),
.A2(n_10),
.B1(n_16),
.B2(n_22),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_L g47 ( 
.A1(n_0),
.A2(n_8),
.B1(n_22),
.B2(n_25),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_0),
.A2(n_38),
.B1(n_94),
.B2(n_95),
.Y(n_93)
);

A2O1A1Ixp33_ASAP7_75t_L g19 ( 
.A1(n_1),
.A2(n_17),
.B(n_20),
.C(n_21),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_1),
.B(n_17),
.Y(n_20)
);

INVx2_ASAP7_75t_SL g23 ( 
.A(n_1),
.Y(n_23)
);

INVx2_ASAP7_75t_SL g85 ( 
.A(n_2),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_2),
.B(n_193),
.Y(n_192)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_3),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g49 ( 
.A1(n_4),
.A2(n_50),
.B1(n_51),
.B2(n_52),
.Y(n_49)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_4),
.Y(n_52)
);

AOI21xp33_ASAP7_75t_L g118 ( 
.A1(n_4),
.A2(n_9),
.B(n_51),
.Y(n_118)
);

O2A1O1Ixp33_ASAP7_75t_L g42 ( 
.A1(n_5),
.A2(n_22),
.B(n_43),
.C(n_44),
.Y(n_42)
);

NAND2xp33_ASAP7_75t_SL g43 ( 
.A(n_5),
.B(n_22),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g44 ( 
.A1(n_5),
.A2(n_6),
.B1(n_45),
.B2(n_46),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_5),
.Y(n_45)
);

OAI32xp33_ASAP7_75t_L g139 ( 
.A1(n_5),
.A2(n_6),
.A3(n_22),
.B1(n_140),
.B2(n_141),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_6),
.Y(n_46)
);

A2O1A1Ixp33_ASAP7_75t_L g53 ( 
.A1(n_6),
.A2(n_49),
.B(n_52),
.C(n_54),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g54 ( 
.A(n_6),
.B(n_52),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_6),
.A2(n_8),
.B1(n_25),
.B2(n_46),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_6),
.A2(n_9),
.B1(n_39),
.B2(n_46),
.Y(n_72)
);

A2O1A1Ixp33_ASAP7_75t_L g117 ( 
.A1(n_6),
.A2(n_39),
.B(n_52),
.C(n_118),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g195 ( 
.A1(n_6),
.A2(n_10),
.B1(n_16),
.B2(n_46),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g15 ( 
.A1(n_7),
.A2(n_10),
.B1(n_16),
.B2(n_17),
.Y(n_15)
);

INVx2_ASAP7_75t_SL g17 ( 
.A(n_7),
.Y(n_17)
);

OAI22xp5_ASAP7_75t_L g24 ( 
.A1(n_7),
.A2(n_8),
.B1(n_17),
.B2(n_25),
.Y(n_24)
);

HAxp5_ASAP7_75t_SL g38 ( 
.A(n_7),
.B(n_39),
.CON(n_38),
.SN(n_38)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_8),
.Y(n_25)
);

AOI22xp33_ASAP7_75t_L g173 ( 
.A1(n_8),
.A2(n_25),
.B1(n_50),
.B2(n_51),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_9),
.Y(n_39)
);

AOI21xp5_ASAP7_75t_L g77 ( 
.A1(n_9),
.A2(n_22),
.B(n_78),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_9),
.B(n_22),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_9),
.A2(n_39),
.B1(n_50),
.B2(n_51),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_9),
.B(n_26),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_9),
.B(n_44),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_10),
.Y(n_16)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_10),
.A2(n_16),
.B1(n_50),
.B2(n_51),
.Y(n_87)
);

XOR2xp5_ASAP7_75t_L g11 ( 
.A(n_12),
.B(n_32),
.Y(n_11)
);

NAND2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_30),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_27),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_14),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_14),
.B(n_34),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_14),
.B(n_34),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g14 ( 
.A1(n_15),
.A2(n_18),
.B1(n_24),
.B2(n_26),
.Y(n_14)
);

AOI22xp5_ASAP7_75t_L g56 ( 
.A1(n_15),
.A2(n_18),
.B1(n_26),
.B2(n_38),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_19),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_SL g29 ( 
.A(n_19),
.B(n_21),
.Y(n_29)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_20),
.Y(n_95)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_21),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_22),
.B(n_23),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_24),
.B(n_29),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_28),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_28),
.B(n_31),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_SL g37 ( 
.A(n_29),
.B(n_38),
.Y(n_37)
);

OAI21xp5_ASAP7_75t_L g32 ( 
.A1(n_33),
.A2(n_61),
.B(n_248),
.Y(n_32)
);

MAJIxp5_ASAP7_75t_L g34 ( 
.A(n_35),
.B(n_56),
.C(n_57),
.Y(n_34)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_35),
.A2(n_36),
.B1(n_244),
.B2(n_246),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_36),
.Y(n_35)
);

MAJIxp5_ASAP7_75t_L g36 ( 
.A(n_37),
.B(n_40),
.C(n_48),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_37),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_37),
.B(n_75),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_37),
.A2(n_73),
.B1(n_75),
.B2(n_76),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_37),
.A2(n_73),
.B1(n_101),
.B2(n_102),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_37),
.B(n_75),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_37),
.A2(n_73),
.B1(n_190),
.B2(n_191),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_37),
.A2(n_73),
.B1(n_218),
.B2(n_219),
.Y(n_217)
);

AOI21xp5_ASAP7_75t_L g225 ( 
.A1(n_37),
.A2(n_191),
.B(n_207),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_37),
.A2(n_73),
.B1(n_228),
.B2(n_232),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_37),
.A2(n_73),
.B1(n_229),
.B2(n_230),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_39),
.B(n_49),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_39),
.B(n_85),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_40),
.A2(n_48),
.B1(n_220),
.B2(n_231),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_40),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g40 ( 
.A1(n_41),
.A2(n_42),
.B1(n_44),
.B2(n_47),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_41),
.A2(n_42),
.B1(n_44),
.B2(n_223),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_42),
.B(n_44),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_45),
.B(n_46),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_47),
.B(n_59),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_48),
.A2(n_220),
.B1(n_221),
.B2(n_222),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_48),
.Y(n_220)
);

AOI21xp5_ASAP7_75t_SL g48 ( 
.A1(n_49),
.A2(n_53),
.B(n_55),
.Y(n_48)
);

AOI21xp5_ASAP7_75t_SL g71 ( 
.A1(n_49),
.A2(n_53),
.B(n_72),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_49),
.A2(n_53),
.B1(n_72),
.B2(n_195),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_49),
.A2(n_53),
.B1(n_55),
.B2(n_195),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_SL g129 ( 
.A(n_50),
.B(n_130),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_51),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_51),
.B(n_85),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_56),
.A2(n_57),
.B1(n_58),
.B2(n_245),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_56),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_58),
.Y(n_57)
);

INVxp67_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_60),
.B(n_77),
.Y(n_76)
);

AOI21xp5_ASAP7_75t_L g61 ( 
.A1(n_62),
.A2(n_241),
.B(n_247),
.Y(n_61)
);

OAI321xp33_ASAP7_75t_L g62 ( 
.A1(n_63),
.A2(n_215),
.A3(n_234),
.B1(n_239),
.B2(n_240),
.C(n_250),
.Y(n_62)
);

AOI21xp5_ASAP7_75t_L g63 ( 
.A1(n_64),
.A2(n_201),
.B(n_214),
.Y(n_63)
);

OAI21xp5_ASAP7_75t_SL g64 ( 
.A1(n_65),
.A2(n_182),
.B(n_200),
.Y(n_64)
);

O2A1O1Ixp33_ASAP7_75t_SL g65 ( 
.A1(n_66),
.A2(n_110),
.B(n_166),
.C(n_181),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_67),
.B(n_98),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_67),
.B(n_98),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g67 ( 
.A(n_68),
.B(n_89),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_69),
.A2(n_70),
.B1(n_81),
.B2(n_82),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_69),
.B(n_82),
.C(n_89),
.Y(n_167)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

AOI211xp5_ASAP7_75t_SL g70 ( 
.A1(n_71),
.A2(n_73),
.B(n_74),
.C(n_80),
.Y(n_70)
);

CKINVDCx16_ASAP7_75t_R g79 ( 
.A(n_71),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_71),
.A2(n_79),
.B1(n_83),
.B2(n_88),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_71),
.A2(n_75),
.B1(n_76),
.B2(n_79),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_71),
.A2(n_79),
.B1(n_121),
.B2(n_122),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_71),
.A2(n_79),
.B1(n_117),
.B2(n_133),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_71),
.B(n_96),
.C(n_121),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_71),
.A2(n_79),
.B1(n_155),
.B2(n_156),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_71),
.B(n_149),
.C(n_155),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_71),
.A2(n_79),
.B1(n_171),
.B2(n_172),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_71),
.B(n_83),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_71),
.B(n_172),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_73),
.B(n_220),
.C(n_222),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_73),
.B(n_232),
.C(n_233),
.Y(n_242)
);

INVxp67_ASAP7_75t_L g147 ( 
.A(n_74),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_75),
.B(n_79),
.Y(n_74)
);

A2O1A1Ixp33_ASAP7_75t_L g146 ( 
.A1(n_75),
.A2(n_79),
.B(n_143),
.C(n_147),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_75),
.A2(n_76),
.B1(n_151),
.B2(n_152),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_76),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_76),
.B(n_96),
.C(n_108),
.Y(n_107)
);

AOI21xp5_ASAP7_75t_L g209 ( 
.A1(n_76),
.A2(n_210),
.B(n_211),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_76),
.B(n_210),
.Y(n_211)
);

INVxp67_ASAP7_75t_L g223 ( 
.A(n_77),
.Y(n_223)
);

CKINVDCx16_ASAP7_75t_R g140 ( 
.A(n_78),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_79),
.B(n_117),
.Y(n_116)
);

AOI21xp5_ASAP7_75t_L g179 ( 
.A1(n_80),
.A2(n_97),
.B(n_180),
.Y(n_179)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_80),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_82),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_83),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_84),
.A2(n_85),
.B1(n_86),
.B2(n_87),
.Y(n_83)
);

AOI21xp5_ASAP7_75t_SL g96 ( 
.A1(n_84),
.A2(n_85),
.B(n_86),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_84),
.A2(n_85),
.B1(n_87),
.B2(n_173),
.Y(n_172)
);

INVxp33_ASAP7_75t_L g193 ( 
.A(n_84),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_90),
.A2(n_91),
.B1(n_92),
.B2(n_97),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_90),
.A2(n_91),
.B1(n_175),
.B2(n_176),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_90),
.A2(n_91),
.B1(n_187),
.B2(n_188),
.Y(n_186)
);

CKINVDCx14_ASAP7_75t_R g90 ( 
.A(n_91),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_92),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_96),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_93),
.A2(n_96),
.B1(n_105),
.B2(n_106),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_93),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_96),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_96),
.A2(n_105),
.B1(n_120),
.B2(n_123),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_96),
.B(n_127),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_96),
.B(n_129),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_96),
.A2(n_105),
.B1(n_139),
.B2(n_142),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_96),
.A2(n_105),
.B1(n_108),
.B2(n_109),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_96),
.B(n_139),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_103),
.C(n_107),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_99),
.A2(n_100),
.B1(n_161),
.B2(n_163),
.Y(n_160)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_101),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_101),
.A2(n_102),
.B1(n_138),
.B2(n_143),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_103),
.A2(n_104),
.B1(n_107),
.B2(n_162),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_104),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_105),
.B(n_132),
.Y(n_131)
);

CKINVDCx14_ASAP7_75t_R g162 ( 
.A(n_107),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_109),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_111),
.B(n_165),
.Y(n_110)
);

AOI21xp5_ASAP7_75t_L g111 ( 
.A1(n_112),
.A2(n_158),
.B(n_164),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_SL g112 ( 
.A1(n_113),
.A2(n_145),
.B(n_157),
.Y(n_112)
);

AOI21xp5_ASAP7_75t_L g113 ( 
.A1(n_114),
.A2(n_135),
.B(n_144),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_SL g114 ( 
.A1(n_115),
.A2(n_124),
.B(n_134),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_119),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_116),
.B(n_119),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_117),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_120),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_122),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_131),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_128),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_137),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_136),
.B(n_137),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_138),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_139),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_148),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_146),
.B(n_148),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_149),
.A2(n_150),
.B1(n_153),
.B2(n_154),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_152),
.Y(n_151)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_156),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_160),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_SL g164 ( 
.A(n_159),
.B(n_160),
.Y(n_164)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_161),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_168),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_SL g181 ( 
.A(n_167),
.B(n_168),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_179),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_170),
.A2(n_174),
.B1(n_177),
.B2(n_178),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_170),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_170),
.B(n_178),
.C(n_179),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_172),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_SL g191 ( 
.A(n_173),
.B(n_192),
.Y(n_191)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_174),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_175),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_SL g197 ( 
.A1(n_175),
.A2(n_198),
.B(n_199),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_180),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_184),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_183),
.B(n_184),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_197),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_189),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_186),
.B(n_189),
.C(n_197),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_187),
.Y(n_188)
);

OAI21xp33_ASAP7_75t_SL g212 ( 
.A1(n_187),
.A2(n_198),
.B(n_199),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_190),
.A2(n_191),
.B1(n_194),
.B2(n_196),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_191),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_191),
.B(n_194),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_194),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_203),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_SL g214 ( 
.A(n_202),
.B(n_203),
.Y(n_214)
);

AOI22xp33_ASAP7_75t_SL g203 ( 
.A1(n_204),
.A2(n_205),
.B1(n_212),
.B2(n_213),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_205),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_209),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_206),
.B(n_209),
.C(n_213),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_208),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_211),
.B(n_217),
.C(n_224),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_211),
.B(n_217),
.Y(n_237)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_212),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_226),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_216),
.B(n_226),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_219),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_222),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_224),
.A2(n_225),
.B1(n_237),
.B2(n_238),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_225),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_233),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_228),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_230),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_235),
.B(n_236),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_235),
.B(n_236),
.Y(n_239)
);

CKINVDCx16_ASAP7_75t_R g238 ( 
.A(n_237),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_242),
.B(n_243),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_242),
.B(n_243),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_244),
.Y(n_246)
);


endmodule