module fake_netlist_5_1741_n_1273 (n_137, n_91, n_82, n_122, n_142, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_60, n_155, n_152, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_125, n_35, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_157, n_29, n_79, n_131, n_151, n_47, n_25, n_53, n_160, n_8, n_158, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_159, n_95, n_119, n_59, n_26, n_133, n_55, n_99, n_2, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_27, n_64, n_77, n_102, n_106, n_161, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_134, n_32, n_41, n_104, n_103, n_56, n_51, n_63, n_97, n_141, n_11, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_1273);

input n_137;
input n_91;
input n_82;
input n_122;
input n_142;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_60;
input n_155;
input n_152;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_125;
input n_35;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_157;
input n_29;
input n_79;
input n_131;
input n_151;
input n_47;
input n_25;
input n_53;
input n_160;
input n_8;
input n_158;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_159;
input n_95;
input n_119;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_27;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_134;
input n_32;
input n_41;
input n_104;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_11;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_1273;

wire n_924;
wire n_1263;
wire n_977;
wire n_611;
wire n_1126;
wire n_1166;
wire n_469;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1150;
wire n_226;
wire n_667;
wire n_790;
wire n_1055;
wire n_880;
wire n_544;
wire n_1007;
wire n_552;
wire n_1198;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1021;
wire n_551;
wire n_688;
wire n_800;
wire n_671;
wire n_819;
wire n_1022;
wire n_915;
wire n_864;
wire n_173;
wire n_859;
wire n_951;
wire n_1264;
wire n_447;
wire n_247;
wire n_292;
wire n_625;
wire n_854;
wire n_674;
wire n_417;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_606;
wire n_275;
wire n_877;
wire n_755;
wire n_1118;
wire n_947;
wire n_373;
wire n_307;
wire n_530;
wire n_1107;
wire n_556;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_929;
wire n_1124;
wire n_902;
wire n_191;
wire n_1104;
wire n_659;
wire n_1257;
wire n_171;
wire n_1182;
wire n_579;
wire n_1261;
wire n_938;
wire n_1098;
wire n_320;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_406;
wire n_519;
wire n_1016;
wire n_1243;
wire n_546;
wire n_281;
wire n_240;
wire n_291;
wire n_231;
wire n_257;
wire n_731;
wire n_371;
wire n_709;
wire n_317;
wire n_1236;
wire n_569;
wire n_227;
wire n_920;
wire n_335;
wire n_370;
wire n_976;
wire n_343;
wire n_308;
wire n_297;
wire n_1078;
wire n_775;
wire n_219;
wire n_600;
wire n_223;
wire n_264;
wire n_955;
wire n_163;
wire n_339;
wire n_1146;
wire n_882;
wire n_183;
wire n_243;
wire n_1036;
wire n_1097;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_215;
wire n_350;
wire n_196;
wire n_798;
wire n_646;
wire n_436;
wire n_1216;
wire n_290;
wire n_580;
wire n_1040;
wire n_578;
wire n_926;
wire n_344;
wire n_1218;
wire n_422;
wire n_475;
wire n_777;
wire n_1070;
wire n_1030;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_496;
wire n_958;
wire n_1034;
wire n_670;
wire n_521;
wire n_663;
wire n_845;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_680;
wire n_395;
wire n_164;
wire n_553;
wire n_901;
wire n_813;
wire n_214;
wire n_675;
wire n_888;
wire n_1167;
wire n_637;
wire n_184;
wire n_446;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_468;
wire n_213;
wire n_342;
wire n_464;
wire n_363;
wire n_197;
wire n_1069;
wire n_1075;
wire n_460;
wire n_889;
wire n_973;
wire n_477;
wire n_571;
wire n_461;
wire n_1211;
wire n_1197;
wire n_907;
wire n_190;
wire n_989;
wire n_1039;
wire n_228;
wire n_283;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1002;
wire n_310;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1248;
wire n_230;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_440;
wire n_793;
wire n_478;
wire n_476;
wire n_534;
wire n_884;
wire n_345;
wire n_944;
wire n_182;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_832;
wire n_857;
wire n_207;
wire n_561;
wire n_1027;
wire n_971;
wire n_1156;
wire n_326;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_596;
wire n_558;
wire n_702;
wire n_822;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1199;
wire n_352;
wire n_1038;
wire n_520;
wire n_409;
wire n_887;
wire n_300;
wire n_809;
wire n_870;
wire n_931;
wire n_599;
wire n_434;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_965;
wire n_935;
wire n_1175;
wire n_817;
wire n_360;
wire n_759;
wire n_806;
wire n_324;
wire n_187;
wire n_1189;
wire n_1259;
wire n_706;
wire n_746;
wire n_747;
wire n_784;
wire n_1244;
wire n_431;
wire n_1194;
wire n_615;
wire n_851;
wire n_843;
wire n_523;
wire n_913;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_776;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_649;
wire n_547;
wire n_1191;
wire n_284;
wire n_1128;
wire n_744;
wire n_590;
wire n_629;
wire n_254;
wire n_1233;
wire n_526;
wire n_372;
wire n_293;
wire n_677;
wire n_244;
wire n_1121;
wire n_368;
wire n_314;
wire n_433;
wire n_604;
wire n_949;
wire n_1008;
wire n_946;
wire n_1001;
wire n_498;
wire n_689;
wire n_738;
wire n_640;
wire n_624;
wire n_252;
wire n_295;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1195;
wire n_610;
wire n_936;
wire n_568;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_259;
wire n_448;
wire n_758;
wire n_999;
wire n_1158;
wire n_563;
wire n_1145;
wire n_878;
wire n_524;
wire n_204;
wire n_394;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1068;
wire n_331;
wire n_906;
wire n_1163;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_658;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_592;
wire n_1169;
wire n_1017;
wire n_978;
wire n_1054;
wire n_1269;
wire n_1095;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_484;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1009;
wire n_1148;
wire n_750;
wire n_742;
wire n_995;
wire n_454;
wire n_374;
wire n_185;
wire n_396;
wire n_1073;
wire n_255;
wire n_662;
wire n_459;
wire n_218;
wire n_962;
wire n_1215;
wire n_1171;
wire n_723;
wire n_1065;
wire n_473;
wire n_1043;
wire n_355;
wire n_486;
wire n_614;
wire n_337;
wire n_1177;
wire n_168;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_208;
wire n_743;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_1240;
wire n_829;
wire n_361;
wire n_1237;
wire n_700;
wire n_573;
wire n_1132;
wire n_388;
wire n_1127;
wire n_761;
wire n_1006;
wire n_329;
wire n_274;
wire n_1270;
wire n_582;
wire n_309;
wire n_512;
wire n_322;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_224;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_239;
wire n_630;
wire n_504;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_987;
wire n_261;
wire n_174;
wire n_767;
wire n_993;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_729;
wire n_1131;
wire n_1084;
wire n_970;
wire n_911;
wire n_513;
wire n_1094;
wire n_560;
wire n_340;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_495;
wire n_602;
wire n_574;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_490;
wire n_996;
wire n_921;
wire n_233;
wire n_572;
wire n_366;
wire n_815;
wire n_327;
wire n_1037;
wire n_1080;
wire n_426;
wire n_1082;
wire n_589;
wire n_716;
wire n_562;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_531;
wire n_890;
wire n_764;
wire n_1056;
wire n_162;
wire n_960;
wire n_222;
wire n_1123;
wire n_1047;
wire n_634;
wire n_199;
wire n_1252;
wire n_348;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_256;
wire n_950;
wire n_380;
wire n_419;
wire n_444;
wire n_1060;
wire n_1141;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_912;
wire n_315;
wire n_968;
wire n_451;
wire n_619;
wire n_408;
wire n_376;
wire n_967;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_483;
wire n_683;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_983;
wire n_280;
wire n_873;
wire n_378;
wire n_1112;
wire n_762;
wire n_690;
wire n_583;
wire n_302;
wire n_1203;
wire n_821;
wire n_321;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_212;
wire n_385;
wire n_507;
wire n_330;
wire n_1228;
wire n_972;
wire n_692;
wire n_820;
wire n_1200;
wire n_1185;
wire n_991;
wire n_828;
wire n_779;
wire n_576;
wire n_1143;
wire n_804;
wire n_537;
wire n_945;
wire n_492;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_286;
wire n_883;
wire n_470;
wire n_325;
wire n_449;
wire n_1214;
wire n_900;
wire n_856;
wire n_918;
wire n_942;
wire n_189;
wire n_1147;
wire n_1077;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_195;
wire n_356;
wire n_894;
wire n_831;
wire n_964;
wire n_1096;
wire n_234;
wire n_833;
wire n_225;
wire n_988;
wire n_814;
wire n_192;
wire n_1201;
wire n_1114;
wire n_655;
wire n_669;
wire n_472;
wire n_1176;
wire n_387;
wire n_1149;
wire n_398;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_211;
wire n_1219;
wire n_1204;
wire n_178;
wire n_1035;
wire n_287;
wire n_555;
wire n_783;
wire n_1188;
wire n_661;
wire n_849;
wire n_336;
wire n_584;
wire n_681;
wire n_430;
wire n_510;
wire n_216;
wire n_311;
wire n_830;
wire n_801;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_445;
wire n_749;
wire n_1134;
wire n_717;
wire n_165;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1019;
wire n_1105;
wire n_249;
wire n_304;
wire n_577;
wire n_338;
wire n_693;
wire n_836;
wire n_990;
wire n_975;
wire n_1256;
wire n_567;
wire n_778;
wire n_1122;
wire n_306;
wire n_458;
wire n_770;
wire n_1102;
wire n_711;
wire n_1187;
wire n_1164;
wire n_489;
wire n_1174;
wire n_617;
wire n_876;
wire n_1190;
wire n_601;
wire n_917;
wire n_966;
wire n_253;
wire n_1116;
wire n_1212;
wire n_172;
wire n_206;
wire n_217;
wire n_726;
wire n_982;
wire n_818;
wire n_861;
wire n_1183;
wire n_899;
wire n_1253;
wire n_210;
wire n_774;
wire n_1059;
wire n_176;
wire n_1133;
wire n_557;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_1168;
wire n_707;
wire n_937;
wire n_393;
wire n_487;
wire n_665;
wire n_177;
wire n_421;
wire n_910;
wire n_768;
wire n_205;
wire n_1136;
wire n_754;
wire n_179;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_735;
wire n_232;
wire n_1109;
wire n_895;
wire n_202;
wire n_427;
wire n_791;
wire n_732;
wire n_193;
wire n_808;
wire n_797;
wire n_1025;
wire n_500;
wire n_1067;
wire n_435;
wire n_766;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_594;
wire n_200;
wire n_1155;
wire n_1184;
wire n_1011;
wire n_985;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_626;
wire n_1144;
wire n_1137;
wire n_1170;
wire n_305;
wire n_676;
wire n_294;
wire n_318;
wire n_653;
wire n_642;
wire n_194;
wire n_855;
wire n_1178;
wire n_850;
wire n_684;
wire n_268;
wire n_664;
wire n_503;
wire n_235;
wire n_605;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_780;
wire n_998;
wire n_467;
wire n_1227;
wire n_840;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_672;
wire n_581;
wire n_382;
wire n_554;
wire n_898;
wire n_1013;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_198;
wire n_714;
wire n_909;
wire n_997;
wire n_932;
wire n_612;
wire n_788;
wire n_1268;
wire n_559;
wire n_825;
wire n_508;
wire n_506;
wire n_737;
wire n_986;
wire n_509;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_209;
wire n_733;
wire n_941;
wire n_981;
wire n_867;
wire n_186;
wire n_587;
wire n_792;
wire n_756;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_518;
wire n_505;
wire n_282;
wire n_752;
wire n_905;
wire n_1108;
wire n_782;
wire n_1100;
wire n_862;
wire n_760;
wire n_381;
wire n_220;
wire n_390;
wire n_481;
wire n_769;
wire n_1046;
wire n_271;
wire n_934;
wire n_826;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_167;
wire n_379;
wire n_428;
wire n_570;
wire n_853;
wire n_377;
wire n_751;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_704;
wire n_787;
wire n_961;
wire n_771;
wire n_276;
wire n_1225;
wire n_169;
wire n_522;
wire n_1262;
wire n_400;
wire n_930;
wire n_181;
wire n_221;
wire n_622;
wire n_1087;
wire n_386;
wire n_994;
wire n_848;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1247;
wire n_922;
wire n_816;
wire n_591;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_432;
wire n_839;
wire n_1210;
wire n_328;
wire n_1250;
wire n_369;
wire n_871;
wire n_598;
wire n_685;
wire n_608;
wire n_928;
wire n_772;
wire n_499;
wire n_517;
wire n_402;
wire n_413;
wire n_1086;
wire n_796;
wire n_236;
wire n_1012;
wire n_903;
wire n_740;
wire n_203;
wire n_384;
wire n_277;
wire n_1061;
wire n_333;
wire n_462;
wire n_1193;
wire n_1255;
wire n_258;
wire n_1113;
wire n_1226;
wire n_722;
wire n_188;
wire n_844;
wire n_201;
wire n_471;
wire n_852;
wire n_1028;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_632;
wire n_699;
wire n_979;
wire n_1245;
wire n_846;
wire n_465;
wire n_362;
wire n_170;
wire n_273;
wire n_585;
wire n_270;
wire n_616;
wire n_745;
wire n_1103;
wire n_648;
wire n_312;
wire n_1076;
wire n_1091;
wire n_494;
wire n_641;
wire n_730;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_180;
wire n_656;
wire n_1220;
wire n_229;
wire n_437;
wire n_453;
wire n_403;
wire n_1130;
wire n_720;
wire n_863;
wire n_805;
wire n_712;
wire n_246;
wire n_1042;
wire n_269;
wire n_285;
wire n_412;
wire n_657;
wire n_644;
wire n_1160;
wire n_491;
wire n_1258;
wire n_1074;
wire n_251;
wire n_566;
wire n_565;
wire n_597;
wire n_1181;
wire n_1196;
wire n_651;
wire n_334;
wire n_811;
wire n_807;
wire n_835;
wire n_175;
wire n_666;
wire n_262;
wire n_1254;
wire n_1026;
wire n_1234;
wire n_319;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_1004;
wire n_1186;
wire n_242;
wire n_1032;
wire n_1018;
wire n_438;
wire n_713;
wire n_904;
wire n_166;
wire n_1180;
wire n_1271;
wire n_533;
wire n_1251;
wire n_278;

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_51),
.Y(n_162)
);

HB1xp67_ASAP7_75t_L g163 ( 
.A(n_38),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_37),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_137),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_133),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_152),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_37),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_93),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_28),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_138),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_135),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_39),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_56),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_156),
.Y(n_175)
);

BUFx8_ASAP7_75t_SL g176 ( 
.A(n_46),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g177 ( 
.A(n_52),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_115),
.Y(n_178)
);

BUFx10_ASAP7_75t_L g179 ( 
.A(n_35),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_39),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_94),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_126),
.Y(n_182)
);

INVx1_ASAP7_75t_SL g183 ( 
.A(n_124),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_30),
.Y(n_184)
);

BUFx8_ASAP7_75t_SL g185 ( 
.A(n_19),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_100),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_40),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_18),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_143),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_62),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_90),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_24),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_159),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_58),
.Y(n_194)
);

INVx1_ASAP7_75t_SL g195 ( 
.A(n_136),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_123),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_0),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_117),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_134),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_95),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_147),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_63),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_131),
.Y(n_203)
);

INVx1_ASAP7_75t_SL g204 ( 
.A(n_127),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_142),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_57),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_76),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_0),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_157),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_149),
.Y(n_210)
);

BUFx6f_ASAP7_75t_L g211 ( 
.A(n_81),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_53),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_60),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_107),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_132),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_114),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_153),
.Y(n_217)
);

BUFx10_ASAP7_75t_L g218 ( 
.A(n_67),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_108),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_3),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_50),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_116),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_84),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_160),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_2),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_121),
.Y(n_226)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_106),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_68),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_45),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_8),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_7),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_15),
.Y(n_232)
);

INVxp67_ASAP7_75t_L g233 ( 
.A(n_144),
.Y(n_233)
);

CKINVDCx16_ASAP7_75t_R g234 ( 
.A(n_129),
.Y(n_234)
);

BUFx3_ASAP7_75t_L g235 ( 
.A(n_111),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_140),
.Y(n_236)
);

INVx2_ASAP7_75t_SL g237 ( 
.A(n_18),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_158),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_150),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_92),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_89),
.Y(n_241)
);

BUFx3_ASAP7_75t_L g242 ( 
.A(n_145),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_9),
.Y(n_243)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_120),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_110),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_148),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_139),
.Y(n_247)
);

INVx1_ASAP7_75t_SL g248 ( 
.A(n_22),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_19),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_4),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_25),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_82),
.Y(n_252)
);

BUFx5_ASAP7_75t_L g253 ( 
.A(n_128),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_12),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_118),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_48),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_49),
.Y(n_257)
);

INVx1_ASAP7_75t_SL g258 ( 
.A(n_32),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_154),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_112),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_14),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_146),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_130),
.Y(n_263)
);

BUFx3_ASAP7_75t_L g264 ( 
.A(n_99),
.Y(n_264)
);

BUFx10_ASAP7_75t_L g265 ( 
.A(n_11),
.Y(n_265)
);

INVx1_ASAP7_75t_SL g266 ( 
.A(n_122),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_24),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_59),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_155),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_141),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_25),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_2),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_70),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_73),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_113),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_125),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_119),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_151),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_75),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_54),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_35),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_4),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_173),
.Y(n_283)
);

INVxp67_ASAP7_75t_L g284 ( 
.A(n_163),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_184),
.Y(n_285)
);

NOR2xp67_ASAP7_75t_L g286 ( 
.A(n_237),
.B(n_1),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_229),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_176),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_243),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_249),
.Y(n_290)
);

INVx1_ASAP7_75t_SL g291 ( 
.A(n_185),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_187),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_225),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_254),
.Y(n_294)
);

NOR2xp67_ASAP7_75t_L g295 ( 
.A(n_237),
.B(n_1),
.Y(n_295)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_253),
.Y(n_296)
);

INVxp67_ASAP7_75t_SL g297 ( 
.A(n_235),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_180),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_235),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_242),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_188),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_192),
.Y(n_302)
);

BUFx6f_ASAP7_75t_SL g303 ( 
.A(n_218),
.Y(n_303)
);

INVxp67_ASAP7_75t_L g304 ( 
.A(n_179),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_242),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_264),
.Y(n_306)
);

INVxp33_ASAP7_75t_SL g307 ( 
.A(n_164),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_164),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_181),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_168),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_264),
.Y(n_311)
);

INVx3_ASAP7_75t_L g312 ( 
.A(n_227),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_168),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_182),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_186),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_177),
.B(n_3),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_165),
.Y(n_317)
);

INVxp67_ASAP7_75t_SL g318 ( 
.A(n_233),
.Y(n_318)
);

BUFx3_ASAP7_75t_L g319 ( 
.A(n_218),
.Y(n_319)
);

INVx1_ASAP7_75t_SL g320 ( 
.A(n_179),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_197),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_167),
.Y(n_322)
);

INVxp67_ASAP7_75t_L g323 ( 
.A(n_179),
.Y(n_323)
);

INVxp67_ASAP7_75t_L g324 ( 
.A(n_265),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_172),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_178),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_208),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_189),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_190),
.Y(n_329)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_253),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_191),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_196),
.Y(n_332)
);

INVxp67_ASAP7_75t_L g333 ( 
.A(n_265),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_202),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_193),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_194),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_170),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_227),
.B(n_5),
.Y(n_338)
);

HB1xp67_ASAP7_75t_L g339 ( 
.A(n_170),
.Y(n_339)
);

INVx2_ASAP7_75t_L g340 ( 
.A(n_253),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_205),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_212),
.Y(n_342)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_253),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_244),
.B(n_253),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g345 ( 
.A(n_281),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_213),
.Y(n_346)
);

CKINVDCx16_ASAP7_75t_R g347 ( 
.A(n_234),
.Y(n_347)
);

BUFx2_ASAP7_75t_L g348 ( 
.A(n_281),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_221),
.Y(n_349)
);

INVxp67_ASAP7_75t_SL g350 ( 
.A(n_223),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_198),
.Y(n_351)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_282),
.Y(n_352)
);

CKINVDCx20_ASAP7_75t_R g353 ( 
.A(n_282),
.Y(n_353)
);

OR2x2_ASAP7_75t_L g354 ( 
.A(n_248),
.B(n_5),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_245),
.Y(n_355)
);

INVxp33_ASAP7_75t_SL g356 ( 
.A(n_220),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_230),
.Y(n_357)
);

INVxp67_ASAP7_75t_L g358 ( 
.A(n_265),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_231),
.Y(n_359)
);

BUFx6f_ASAP7_75t_L g360 ( 
.A(n_211),
.Y(n_360)
);

BUFx2_ASAP7_75t_L g361 ( 
.A(n_232),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_199),
.Y(n_362)
);

CKINVDCx20_ASAP7_75t_R g363 ( 
.A(n_250),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_247),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_200),
.Y(n_365)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_251),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_259),
.Y(n_367)
);

INVx1_ASAP7_75t_SL g368 ( 
.A(n_258),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_263),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_269),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_201),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_203),
.Y(n_372)
);

INVxp67_ASAP7_75t_SL g373 ( 
.A(n_274),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_360),
.Y(n_374)
);

AND2x2_ASAP7_75t_L g375 ( 
.A(n_297),
.B(n_218),
.Y(n_375)
);

BUFx6f_ASAP7_75t_L g376 ( 
.A(n_360),
.Y(n_376)
);

INVx3_ASAP7_75t_L g377 ( 
.A(n_360),
.Y(n_377)
);

HB1xp67_ASAP7_75t_L g378 ( 
.A(n_368),
.Y(n_378)
);

AND2x2_ASAP7_75t_L g379 ( 
.A(n_299),
.B(n_183),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_360),
.Y(n_380)
);

INVx2_ASAP7_75t_L g381 ( 
.A(n_360),
.Y(n_381)
);

BUFx6f_ASAP7_75t_L g382 ( 
.A(n_296),
.Y(n_382)
);

INVx2_ASAP7_75t_L g383 ( 
.A(n_296),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_312),
.Y(n_384)
);

AND2x4_ASAP7_75t_L g385 ( 
.A(n_350),
.B(n_373),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_312),
.Y(n_386)
);

AND2x4_ASAP7_75t_L g387 ( 
.A(n_317),
.B(n_244),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_312),
.Y(n_388)
);

BUFx6f_ASAP7_75t_L g389 ( 
.A(n_330),
.Y(n_389)
);

INVx1_ASAP7_75t_SL g390 ( 
.A(n_320),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_283),
.Y(n_391)
);

NOR2xp33_ASAP7_75t_L g392 ( 
.A(n_356),
.B(n_195),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_285),
.Y(n_393)
);

INVx5_ASAP7_75t_L g394 ( 
.A(n_330),
.Y(n_394)
);

INVx3_ASAP7_75t_L g395 ( 
.A(n_340),
.Y(n_395)
);

AND2x2_ASAP7_75t_L g396 ( 
.A(n_300),
.B(n_204),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_322),
.B(n_162),
.Y(n_397)
);

INVx3_ASAP7_75t_L g398 ( 
.A(n_340),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_287),
.Y(n_399)
);

INVx3_ASAP7_75t_L g400 ( 
.A(n_343),
.Y(n_400)
);

INVx2_ASAP7_75t_L g401 ( 
.A(n_343),
.Y(n_401)
);

BUFx6f_ASAP7_75t_L g402 ( 
.A(n_344),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_325),
.B(n_326),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_289),
.Y(n_404)
);

BUFx6f_ASAP7_75t_L g405 ( 
.A(n_331),
.Y(n_405)
);

AND2x4_ASAP7_75t_L g406 ( 
.A(n_332),
.B(n_211),
.Y(n_406)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_334),
.Y(n_407)
);

BUFx6f_ASAP7_75t_L g408 ( 
.A(n_341),
.Y(n_408)
);

BUFx6f_ASAP7_75t_L g409 ( 
.A(n_342),
.Y(n_409)
);

INVx2_ASAP7_75t_SL g410 ( 
.A(n_319),
.Y(n_410)
);

BUFx6f_ASAP7_75t_L g411 ( 
.A(n_346),
.Y(n_411)
);

BUFx6f_ASAP7_75t_L g412 ( 
.A(n_349),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_290),
.Y(n_413)
);

BUFx6f_ASAP7_75t_L g414 ( 
.A(n_355),
.Y(n_414)
);

AND2x4_ASAP7_75t_L g415 ( 
.A(n_364),
.B(n_211),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_294),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_367),
.B(n_369),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_370),
.Y(n_418)
);

AND2x2_ASAP7_75t_L g419 ( 
.A(n_305),
.B(n_306),
.Y(n_419)
);

AND2x2_ASAP7_75t_L g420 ( 
.A(n_311),
.B(n_266),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_338),
.B(n_162),
.Y(n_421)
);

INVx2_ASAP7_75t_L g422 ( 
.A(n_316),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_286),
.Y(n_423)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_318),
.Y(n_424)
);

BUFx2_ASAP7_75t_L g425 ( 
.A(n_308),
.Y(n_425)
);

INVx2_ASAP7_75t_L g426 ( 
.A(n_319),
.Y(n_426)
);

BUFx3_ASAP7_75t_L g427 ( 
.A(n_309),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_295),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_354),
.Y(n_429)
);

BUFx2_ASAP7_75t_L g430 ( 
.A(n_308),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_314),
.B(n_315),
.Y(n_431)
);

INVx3_ASAP7_75t_L g432 ( 
.A(n_328),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_361),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_329),
.Y(n_434)
);

BUFx6f_ASAP7_75t_L g435 ( 
.A(n_335),
.Y(n_435)
);

BUFx6f_ASAP7_75t_L g436 ( 
.A(n_336),
.Y(n_436)
);

INVx2_ASAP7_75t_L g437 ( 
.A(n_351),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_362),
.B(n_365),
.Y(n_438)
);

BUFx6f_ASAP7_75t_L g439 ( 
.A(n_371),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_372),
.Y(n_440)
);

OAI22xp5_ASAP7_75t_SL g441 ( 
.A1(n_310),
.A2(n_261),
.B1(n_271),
.B2(n_267),
.Y(n_441)
);

BUFx6f_ASAP7_75t_L g442 ( 
.A(n_348),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_284),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_383),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_378),
.Y(n_445)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_383),
.Y(n_446)
);

AOI22xp33_ASAP7_75t_L g447 ( 
.A1(n_422),
.A2(n_402),
.B1(n_424),
.B2(n_385),
.Y(n_447)
);

INVx4_ASAP7_75t_L g448 ( 
.A(n_394),
.Y(n_448)
);

AND2x2_ASAP7_75t_L g449 ( 
.A(n_424),
.B(n_339),
.Y(n_449)
);

INVx2_ASAP7_75t_SL g450 ( 
.A(n_378),
.Y(n_450)
);

INVx1_ASAP7_75t_SL g451 ( 
.A(n_390),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_SL g452 ( 
.A(n_392),
.B(n_347),
.Y(n_452)
);

INVx3_ASAP7_75t_L g453 ( 
.A(n_382),
.Y(n_453)
);

NAND3xp33_ASAP7_75t_L g454 ( 
.A(n_422),
.B(n_211),
.C(n_210),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_402),
.B(n_298),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_383),
.Y(n_456)
);

AND2x4_ASAP7_75t_L g457 ( 
.A(n_419),
.B(n_211),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_401),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_401),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_402),
.B(n_385),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_402),
.B(n_298),
.Y(n_461)
);

AO21x2_ASAP7_75t_L g462 ( 
.A1(n_421),
.A2(n_323),
.B(n_304),
.Y(n_462)
);

AND2x2_ASAP7_75t_L g463 ( 
.A(n_424),
.B(n_301),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_401),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_402),
.B(n_385),
.Y(n_465)
);

NAND2xp33_ASAP7_75t_SL g466 ( 
.A(n_441),
.B(n_363),
.Y(n_466)
);

NOR2xp33_ASAP7_75t_L g467 ( 
.A(n_434),
.B(n_356),
.Y(n_467)
);

NOR2xp33_ASAP7_75t_L g468 ( 
.A(n_434),
.B(n_307),
.Y(n_468)
);

BUFx6f_ASAP7_75t_SL g469 ( 
.A(n_435),
.Y(n_469)
);

AO21x2_ASAP7_75t_L g470 ( 
.A1(n_421),
.A2(n_333),
.B(n_324),
.Y(n_470)
);

AND2x6_ASAP7_75t_L g471 ( 
.A(n_402),
.B(n_291),
.Y(n_471)
);

INVx2_ASAP7_75t_L g472 ( 
.A(n_395),
.Y(n_472)
);

AO21x2_ASAP7_75t_L g473 ( 
.A1(n_431),
.A2(n_358),
.B(n_253),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_385),
.B(n_301),
.Y(n_474)
);

BUFx10_ASAP7_75t_L g475 ( 
.A(n_435),
.Y(n_475)
);

BUFx3_ASAP7_75t_L g476 ( 
.A(n_419),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_422),
.B(n_302),
.Y(n_477)
);

INVx2_ASAP7_75t_L g478 ( 
.A(n_395),
.Y(n_478)
);

NOR3xp33_ASAP7_75t_L g479 ( 
.A(n_390),
.B(n_321),
.C(n_302),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_395),
.Y(n_480)
);

AOI22xp33_ASAP7_75t_L g481 ( 
.A1(n_429),
.A2(n_307),
.B1(n_303),
.B2(n_253),
.Y(n_481)
);

NOR2xp33_ASAP7_75t_L g482 ( 
.A(n_440),
.B(n_321),
.Y(n_482)
);

BUFx3_ASAP7_75t_L g483 ( 
.A(n_426),
.Y(n_483)
);

OR2x6_ASAP7_75t_L g484 ( 
.A(n_437),
.B(n_206),
.Y(n_484)
);

NOR2xp33_ASAP7_75t_L g485 ( 
.A(n_440),
.B(n_327),
.Y(n_485)
);

INVx2_ASAP7_75t_L g486 ( 
.A(n_395),
.Y(n_486)
);

NOR2xp33_ASAP7_75t_L g487 ( 
.A(n_437),
.B(n_327),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_398),
.Y(n_488)
);

INVx2_ASAP7_75t_L g489 ( 
.A(n_398),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_410),
.B(n_357),
.Y(n_490)
);

BUFx6f_ASAP7_75t_L g491 ( 
.A(n_376),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_410),
.B(n_357),
.Y(n_492)
);

AOI22xp5_ASAP7_75t_L g493 ( 
.A1(n_441),
.A2(n_214),
.B1(n_209),
.B2(n_345),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_398),
.Y(n_494)
);

INVx2_ASAP7_75t_L g495 ( 
.A(n_398),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_400),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_400),
.Y(n_497)
);

INVx2_ASAP7_75t_L g498 ( 
.A(n_400),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_400),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_407),
.Y(n_500)
);

INVx4_ASAP7_75t_L g501 ( 
.A(n_394),
.Y(n_501)
);

AND2x2_ASAP7_75t_L g502 ( 
.A(n_379),
.B(n_396),
.Y(n_502)
);

CKINVDCx5p33_ASAP7_75t_R g503 ( 
.A(n_427),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_407),
.Y(n_504)
);

XOR2x2_ASAP7_75t_L g505 ( 
.A(n_425),
.B(n_292),
.Y(n_505)
);

NAND3xp33_ASAP7_75t_L g506 ( 
.A(n_387),
.B(n_215),
.C(n_207),
.Y(n_506)
);

NOR2xp33_ASAP7_75t_L g507 ( 
.A(n_437),
.B(n_431),
.Y(n_507)
);

AND2x2_ASAP7_75t_L g508 ( 
.A(n_379),
.B(n_359),
.Y(n_508)
);

NOR2xp33_ASAP7_75t_SL g509 ( 
.A(n_427),
.B(n_288),
.Y(n_509)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_382),
.Y(n_510)
);

AOI22xp33_ASAP7_75t_L g511 ( 
.A1(n_429),
.A2(n_387),
.B1(n_420),
.B2(n_396),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_SL g512 ( 
.A(n_442),
.B(n_359),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_SL g513 ( 
.A(n_442),
.B(n_363),
.Y(n_513)
);

AOI22xp33_ASAP7_75t_L g514 ( 
.A1(n_387),
.A2(n_303),
.B1(n_253),
.B2(n_352),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_483),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_447),
.B(n_432),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_507),
.B(n_432),
.Y(n_517)
);

INVx2_ASAP7_75t_L g518 ( 
.A(n_446),
.Y(n_518)
);

NOR2xp33_ASAP7_75t_L g519 ( 
.A(n_451),
.B(n_438),
.Y(n_519)
);

NAND2x1_ASAP7_75t_L g520 ( 
.A(n_453),
.B(n_377),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_460),
.B(n_432),
.Y(n_521)
);

INVx2_ASAP7_75t_SL g522 ( 
.A(n_450),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_SL g523 ( 
.A(n_465),
.B(n_442),
.Y(n_523)
);

INVx2_ASAP7_75t_L g524 ( 
.A(n_446),
.Y(n_524)
);

OR2x2_ASAP7_75t_L g525 ( 
.A(n_450),
.B(n_433),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_483),
.Y(n_526)
);

BUFx3_ASAP7_75t_L g527 ( 
.A(n_476),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_483),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_SL g529 ( 
.A(n_502),
.B(n_442),
.Y(n_529)
);

HB1xp67_ASAP7_75t_L g530 ( 
.A(n_445),
.Y(n_530)
);

NOR2xp33_ASAP7_75t_L g531 ( 
.A(n_487),
.B(n_438),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_SL g532 ( 
.A(n_502),
.B(n_442),
.Y(n_532)
);

INVx2_ASAP7_75t_L g533 ( 
.A(n_446),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_476),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_476),
.Y(n_535)
);

INVx2_ASAP7_75t_SL g536 ( 
.A(n_449),
.Y(n_536)
);

AOI22xp33_ASAP7_75t_L g537 ( 
.A1(n_473),
.A2(n_442),
.B1(n_375),
.B2(n_439),
.Y(n_537)
);

HB1xp67_ASAP7_75t_L g538 ( 
.A(n_455),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_461),
.B(n_432),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_500),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_L g541 ( 
.A(n_463),
.B(n_436),
.Y(n_541)
);

OAI22xp5_ASAP7_75t_L g542 ( 
.A1(n_474),
.A2(n_439),
.B1(n_436),
.B2(n_435),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_463),
.B(n_436),
.Y(n_543)
);

NOR2xp33_ASAP7_75t_L g544 ( 
.A(n_477),
.B(n_436),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_L g545 ( 
.A(n_457),
.B(n_436),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_SL g546 ( 
.A(n_475),
.B(n_442),
.Y(n_546)
);

AND2x2_ASAP7_75t_L g547 ( 
.A(n_449),
.B(n_375),
.Y(n_547)
);

INVxp67_ASAP7_75t_L g548 ( 
.A(n_508),
.Y(n_548)
);

NOR2xp33_ASAP7_75t_L g549 ( 
.A(n_468),
.B(n_436),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_L g550 ( 
.A(n_457),
.B(n_436),
.Y(n_550)
);

OR2x2_ASAP7_75t_L g551 ( 
.A(n_508),
.B(n_433),
.Y(n_551)
);

INVxp67_ASAP7_75t_L g552 ( 
.A(n_467),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_L g553 ( 
.A(n_457),
.B(n_439),
.Y(n_553)
);

INVx3_ASAP7_75t_L g554 ( 
.A(n_510),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_500),
.Y(n_555)
);

INVx2_ASAP7_75t_SL g556 ( 
.A(n_457),
.Y(n_556)
);

INVxp67_ASAP7_75t_SL g557 ( 
.A(n_453),
.Y(n_557)
);

BUFx6f_ASAP7_75t_SL g558 ( 
.A(n_484),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_SL g559 ( 
.A(n_475),
.B(n_439),
.Y(n_559)
);

BUFx6f_ASAP7_75t_SL g560 ( 
.A(n_484),
.Y(n_560)
);

OAI21xp5_ASAP7_75t_L g561 ( 
.A1(n_454),
.A2(n_397),
.B(n_420),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_504),
.Y(n_562)
);

BUFx6f_ASAP7_75t_SL g563 ( 
.A(n_484),
.Y(n_563)
);

INVx3_ASAP7_75t_L g564 ( 
.A(n_510),
.Y(n_564)
);

NOR2xp67_ASAP7_75t_L g565 ( 
.A(n_454),
.B(n_410),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_L g566 ( 
.A(n_511),
.B(n_439),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_504),
.Y(n_567)
);

AND2x4_ASAP7_75t_L g568 ( 
.A(n_506),
.B(n_426),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_444),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_480),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_SL g571 ( 
.A(n_475),
.B(n_439),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_SL g572 ( 
.A(n_475),
.B(n_439),
.Y(n_572)
);

NOR2xp33_ASAP7_75t_L g573 ( 
.A(n_482),
.B(n_435),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_L g574 ( 
.A(n_462),
.B(n_435),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_480),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_488),
.Y(n_576)
);

NOR2xp67_ASAP7_75t_L g577 ( 
.A(n_506),
.B(n_503),
.Y(n_577)
);

BUFx6f_ASAP7_75t_L g578 ( 
.A(n_491),
.Y(n_578)
);

INVx2_ASAP7_75t_SL g579 ( 
.A(n_473),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_488),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_L g581 ( 
.A(n_462),
.B(n_435),
.Y(n_581)
);

NOR2xp33_ASAP7_75t_L g582 ( 
.A(n_485),
.B(n_366),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_444),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_SL g584 ( 
.A(n_514),
.B(n_427),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_SL g585 ( 
.A(n_481),
.B(n_426),
.Y(n_585)
);

INVx1_ASAP7_75t_SL g586 ( 
.A(n_505),
.Y(n_586)
);

NOR2xp33_ASAP7_75t_L g587 ( 
.A(n_490),
.B(n_366),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_L g588 ( 
.A(n_462),
.B(n_423),
.Y(n_588)
);

NAND3xp33_ASAP7_75t_L g589 ( 
.A(n_479),
.B(n_492),
.C(n_452),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_494),
.Y(n_590)
);

INVx3_ASAP7_75t_L g591 ( 
.A(n_491),
.Y(n_591)
);

NOR2xp33_ASAP7_75t_SL g592 ( 
.A(n_509),
.B(n_469),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_L g593 ( 
.A(n_470),
.B(n_423),
.Y(n_593)
);

INVx2_ASAP7_75t_SL g594 ( 
.A(n_473),
.Y(n_594)
);

NOR2xp33_ASAP7_75t_L g595 ( 
.A(n_470),
.B(n_512),
.Y(n_595)
);

NAND2xp33_ASAP7_75t_L g596 ( 
.A(n_471),
.B(n_382),
.Y(n_596)
);

HB1xp67_ASAP7_75t_L g597 ( 
.A(n_484),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_L g598 ( 
.A(n_470),
.B(n_428),
.Y(n_598)
);

AND2x2_ASAP7_75t_L g599 ( 
.A(n_484),
.B(n_428),
.Y(n_599)
);

AOI22xp33_ASAP7_75t_L g600 ( 
.A1(n_471),
.A2(n_415),
.B1(n_406),
.B2(n_387),
.Y(n_600)
);

AOI22xp33_ASAP7_75t_L g601 ( 
.A1(n_471),
.A2(n_456),
.B1(n_459),
.B2(n_458),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_494),
.Y(n_602)
);

NAND2xp33_ASAP7_75t_L g603 ( 
.A(n_471),
.B(n_382),
.Y(n_603)
);

INVx2_ASAP7_75t_L g604 ( 
.A(n_456),
.Y(n_604)
);

INVx2_ASAP7_75t_L g605 ( 
.A(n_458),
.Y(n_605)
);

AND2x2_ASAP7_75t_L g606 ( 
.A(n_513),
.B(n_443),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_496),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_453),
.B(n_405),
.Y(n_608)
);

AND2x2_ASAP7_75t_L g609 ( 
.A(n_496),
.B(n_443),
.Y(n_609)
);

NOR3xp33_ASAP7_75t_L g610 ( 
.A(n_466),
.B(n_430),
.C(n_425),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_499),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_499),
.Y(n_612)
);

O2A1O1Ixp33_ASAP7_75t_SL g613 ( 
.A1(n_516),
.A2(n_397),
.B(n_464),
.C(n_459),
.Y(n_613)
);

INVx2_ASAP7_75t_L g614 ( 
.A(n_567),
.Y(n_614)
);

INVx2_ASAP7_75t_L g615 ( 
.A(n_567),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_534),
.Y(n_616)
);

CKINVDCx5p33_ASAP7_75t_R g617 ( 
.A(n_519),
.Y(n_617)
);

AOI21xp5_ASAP7_75t_L g618 ( 
.A1(n_596),
.A2(n_491),
.B(n_453),
.Y(n_618)
);

AOI21xp5_ASAP7_75t_L g619 ( 
.A1(n_596),
.A2(n_491),
.B(n_448),
.Y(n_619)
);

OAI21xp5_ASAP7_75t_L g620 ( 
.A1(n_521),
.A2(n_471),
.B(n_464),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_L g621 ( 
.A(n_531),
.B(n_471),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_535),
.Y(n_622)
);

O2A1O1Ixp5_ASAP7_75t_L g623 ( 
.A1(n_585),
.A2(n_486),
.B(n_478),
.C(n_498),
.Y(n_623)
);

AOI21x1_ASAP7_75t_L g624 ( 
.A1(n_545),
.A2(n_486),
.B(n_478),
.Y(n_624)
);

NOR2xp33_ASAP7_75t_L g625 ( 
.A(n_552),
.B(n_493),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_L g626 ( 
.A(n_573),
.B(n_471),
.Y(n_626)
);

CKINVDCx8_ASAP7_75t_R g627 ( 
.A(n_582),
.Y(n_627)
);

AOI21xp5_ASAP7_75t_L g628 ( 
.A1(n_603),
.A2(n_491),
.B(n_448),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_517),
.B(n_472),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_L g630 ( 
.A(n_549),
.B(n_472),
.Y(n_630)
);

BUFx6f_ASAP7_75t_L g631 ( 
.A(n_578),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g632 ( 
.A(n_538),
.B(n_544),
.Y(n_632)
);

NOR2xp33_ASAP7_75t_L g633 ( 
.A(n_548),
.B(n_493),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_L g634 ( 
.A(n_541),
.B(n_472),
.Y(n_634)
);

AOI21xp5_ASAP7_75t_L g635 ( 
.A1(n_603),
.A2(n_501),
.B(n_448),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_SL g636 ( 
.A(n_543),
.B(n_489),
.Y(n_636)
);

O2A1O1Ixp33_ASAP7_75t_L g637 ( 
.A1(n_588),
.A2(n_418),
.B(n_417),
.C(n_403),
.Y(n_637)
);

AND2x2_ASAP7_75t_L g638 ( 
.A(n_547),
.B(n_430),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_L g639 ( 
.A(n_547),
.B(n_489),
.Y(n_639)
);

AOI21xp5_ASAP7_75t_L g640 ( 
.A1(n_550),
.A2(n_501),
.B(n_448),
.Y(n_640)
);

BUFx2_ASAP7_75t_L g641 ( 
.A(n_530),
.Y(n_641)
);

AOI21xp5_ASAP7_75t_L g642 ( 
.A1(n_553),
.A2(n_501),
.B(n_394),
.Y(n_642)
);

BUFx3_ASAP7_75t_L g643 ( 
.A(n_527),
.Y(n_643)
);

INVx2_ASAP7_75t_L g644 ( 
.A(n_569),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_L g645 ( 
.A(n_536),
.B(n_489),
.Y(n_645)
);

INVx2_ASAP7_75t_L g646 ( 
.A(n_569),
.Y(n_646)
);

O2A1O1Ixp33_ASAP7_75t_L g647 ( 
.A1(n_593),
.A2(n_418),
.B(n_403),
.C(n_417),
.Y(n_647)
);

AOI21xp5_ASAP7_75t_L g648 ( 
.A1(n_559),
.A2(n_501),
.B(n_394),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_570),
.Y(n_649)
);

AOI22xp33_ASAP7_75t_L g650 ( 
.A1(n_579),
.A2(n_469),
.B1(n_310),
.B2(n_313),
.Y(n_650)
);

AND2x2_ASAP7_75t_SL g651 ( 
.A(n_592),
.B(n_469),
.Y(n_651)
);

INVx1_ASAP7_75t_SL g652 ( 
.A(n_525),
.Y(n_652)
);

AOI21xp5_ASAP7_75t_L g653 ( 
.A1(n_559),
.A2(n_394),
.B(n_389),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_L g654 ( 
.A(n_536),
.B(n_495),
.Y(n_654)
);

OAI321xp33_ASAP7_75t_L g655 ( 
.A1(n_561),
.A2(n_393),
.A3(n_416),
.B1(n_404),
.B2(n_399),
.C(n_391),
.Y(n_655)
);

AOI21x1_ASAP7_75t_L g656 ( 
.A1(n_520),
.A2(n_497),
.B(n_495),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_L g657 ( 
.A(n_539),
.B(n_495),
.Y(n_657)
);

AOI21xp5_ASAP7_75t_L g658 ( 
.A1(n_571),
.A2(n_394),
.B(n_389),
.Y(n_658)
);

A2O1A1Ixp33_ASAP7_75t_L g659 ( 
.A1(n_595),
.A2(n_391),
.B(n_416),
.C(n_399),
.Y(n_659)
);

AND2x2_ASAP7_75t_L g660 ( 
.A(n_522),
.B(n_313),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_L g661 ( 
.A(n_598),
.B(n_497),
.Y(n_661)
);

BUFx4f_ASAP7_75t_L g662 ( 
.A(n_551),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_L g663 ( 
.A(n_529),
.B(n_497),
.Y(n_663)
);

AND2x2_ASAP7_75t_L g664 ( 
.A(n_522),
.B(n_337),
.Y(n_664)
);

AOI22xp5_ASAP7_75t_L g665 ( 
.A1(n_566),
.A2(n_353),
.B1(n_352),
.B2(n_345),
.Y(n_665)
);

AOI21xp5_ASAP7_75t_L g666 ( 
.A1(n_571),
.A2(n_394),
.B(n_389),
.Y(n_666)
);

INVx2_ASAP7_75t_L g667 ( 
.A(n_583),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_SL g668 ( 
.A(n_574),
.B(n_581),
.Y(n_668)
);

AOI21xp5_ASAP7_75t_L g669 ( 
.A1(n_572),
.A2(n_389),
.B(n_382),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_575),
.Y(n_670)
);

OAI21xp33_ASAP7_75t_L g671 ( 
.A1(n_525),
.A2(n_353),
.B(n_337),
.Y(n_671)
);

INVx2_ASAP7_75t_L g672 ( 
.A(n_583),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_529),
.B(n_498),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_SL g674 ( 
.A(n_537),
.B(n_498),
.Y(n_674)
);

AND2x2_ASAP7_75t_L g675 ( 
.A(n_606),
.B(n_505),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_532),
.B(n_405),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_576),
.Y(n_677)
);

AOI21xp5_ASAP7_75t_L g678 ( 
.A1(n_572),
.A2(n_389),
.B(n_382),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_L g679 ( 
.A(n_532),
.B(n_405),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_580),
.Y(n_680)
);

AOI21xp5_ASAP7_75t_L g681 ( 
.A1(n_601),
.A2(n_389),
.B(n_382),
.Y(n_681)
);

A2O1A1Ixp33_ASAP7_75t_L g682 ( 
.A1(n_587),
.A2(n_393),
.B(n_404),
.C(n_413),
.Y(n_682)
);

O2A1O1Ixp33_ASAP7_75t_L g683 ( 
.A1(n_584),
.A2(n_585),
.B(n_523),
.C(n_542),
.Y(n_683)
);

AOI21xp5_ASAP7_75t_L g684 ( 
.A1(n_523),
.A2(n_389),
.B(n_376),
.Y(n_684)
);

INVx3_ASAP7_75t_L g685 ( 
.A(n_527),
.Y(n_685)
);

AOI22xp5_ASAP7_75t_L g686 ( 
.A1(n_568),
.A2(n_405),
.B1(n_408),
.B2(n_409),
.Y(n_686)
);

NAND2xp33_ASAP7_75t_L g687 ( 
.A(n_556),
.B(n_216),
.Y(n_687)
);

INVx3_ASAP7_75t_L g688 ( 
.A(n_554),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_L g689 ( 
.A(n_609),
.B(n_405),
.Y(n_689)
);

AOI21xp5_ASAP7_75t_L g690 ( 
.A1(n_556),
.A2(n_376),
.B(n_377),
.Y(n_690)
);

CKINVDCx5p33_ASAP7_75t_R g691 ( 
.A(n_558),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_L g692 ( 
.A(n_609),
.B(n_405),
.Y(n_692)
);

OR2x2_ASAP7_75t_L g693 ( 
.A(n_551),
.B(n_413),
.Y(n_693)
);

OAI21xp5_ASAP7_75t_L g694 ( 
.A1(n_579),
.A2(n_380),
.B(n_374),
.Y(n_694)
);

AOI21xp5_ASAP7_75t_L g695 ( 
.A1(n_600),
.A2(n_376),
.B(n_377),
.Y(n_695)
);

BUFx6f_ASAP7_75t_L g696 ( 
.A(n_578),
.Y(n_696)
);

INVx3_ASAP7_75t_L g697 ( 
.A(n_554),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_L g698 ( 
.A(n_606),
.B(n_408),
.Y(n_698)
);

OAI21xp5_ASAP7_75t_L g699 ( 
.A1(n_594),
.A2(n_568),
.B(n_526),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_SL g700 ( 
.A(n_568),
.B(n_409),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_590),
.Y(n_701)
);

AOI21xp5_ASAP7_75t_L g702 ( 
.A1(n_557),
.A2(n_376),
.B(n_377),
.Y(n_702)
);

NAND2x1p5_ASAP7_75t_L g703 ( 
.A(n_546),
.B(n_384),
.Y(n_703)
);

OR2x2_ASAP7_75t_L g704 ( 
.A(n_586),
.B(n_292),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_L g705 ( 
.A(n_515),
.B(n_408),
.Y(n_705)
);

INVx4_ASAP7_75t_L g706 ( 
.A(n_578),
.Y(n_706)
);

OR2x2_ASAP7_75t_L g707 ( 
.A(n_589),
.B(n_293),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_SL g708 ( 
.A(n_594),
.B(n_409),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_602),
.Y(n_709)
);

NOR3xp33_ASAP7_75t_SL g710 ( 
.A(n_617),
.B(n_584),
.C(n_272),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_L g711 ( 
.A(n_632),
.B(n_577),
.Y(n_711)
);

A2O1A1Ixp33_ASAP7_75t_SL g712 ( 
.A1(n_621),
.A2(n_610),
.B(n_599),
.C(n_591),
.Y(n_712)
);

AND2x4_ASAP7_75t_L g713 ( 
.A(n_643),
.B(n_599),
.Y(n_713)
);

AOI22xp33_ASAP7_75t_L g714 ( 
.A1(n_625),
.A2(n_558),
.B1(n_560),
.B2(n_563),
.Y(n_714)
);

AND2x2_ASAP7_75t_L g715 ( 
.A(n_662),
.B(n_597),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_668),
.B(n_565),
.Y(n_716)
);

AOI221xp5_ASAP7_75t_L g717 ( 
.A1(n_625),
.A2(n_256),
.B1(n_558),
.B2(n_560),
.C(n_563),
.Y(n_717)
);

BUFx6f_ASAP7_75t_L g718 ( 
.A(n_631),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_SL g719 ( 
.A(n_662),
.B(n_546),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_SL g720 ( 
.A(n_651),
.B(n_578),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_614),
.Y(n_721)
);

AO32x1_ASAP7_75t_L g722 ( 
.A1(n_614),
.A2(n_540),
.A3(n_555),
.B1(n_562),
.B2(n_604),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_646),
.Y(n_723)
);

INVx2_ASAP7_75t_L g724 ( 
.A(n_646),
.Y(n_724)
);

INVx3_ASAP7_75t_L g725 ( 
.A(n_631),
.Y(n_725)
);

BUFx2_ASAP7_75t_L g726 ( 
.A(n_641),
.Y(n_726)
);

OAI22xp5_ASAP7_75t_L g727 ( 
.A1(n_651),
.A2(n_560),
.B1(n_563),
.B2(n_528),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_SL g728 ( 
.A(n_652),
.B(n_607),
.Y(n_728)
);

NOR2xp33_ASAP7_75t_L g729 ( 
.A(n_627),
.B(n_293),
.Y(n_729)
);

NAND3xp33_ASAP7_75t_SL g730 ( 
.A(n_665),
.B(n_169),
.C(n_166),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_SL g731 ( 
.A(n_650),
.B(n_611),
.Y(n_731)
);

OAI22xp5_ASAP7_75t_L g732 ( 
.A1(n_626),
.A2(n_699),
.B1(n_685),
.B2(n_668),
.Y(n_732)
);

A2O1A1Ixp33_ASAP7_75t_L g733 ( 
.A1(n_683),
.A2(n_612),
.B(n_604),
.C(n_605),
.Y(n_733)
);

NOR2xp33_ASAP7_75t_L g734 ( 
.A(n_671),
.B(n_303),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_615),
.Y(n_735)
);

AND2x2_ASAP7_75t_L g736 ( 
.A(n_638),
.B(n_407),
.Y(n_736)
);

HB1xp67_ASAP7_75t_L g737 ( 
.A(n_643),
.Y(n_737)
);

A2O1A1Ixp33_ASAP7_75t_L g738 ( 
.A1(n_633),
.A2(n_605),
.B(n_554),
.C(n_564),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_649),
.B(n_670),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_644),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_SL g741 ( 
.A(n_650),
.B(n_591),
.Y(n_741)
);

AO32x2_ASAP7_75t_L g742 ( 
.A1(n_706),
.A2(n_659),
.A3(n_655),
.B1(n_613),
.B2(n_682),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_SL g743 ( 
.A(n_660),
.B(n_591),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_SL g744 ( 
.A(n_664),
.B(n_564),
.Y(n_744)
);

O2A1O1Ixp33_ASAP7_75t_L g745 ( 
.A1(n_682),
.A2(n_608),
.B(n_533),
.C(n_524),
.Y(n_745)
);

A2O1A1Ixp33_ASAP7_75t_L g746 ( 
.A1(n_633),
.A2(n_564),
.B(n_533),
.C(n_524),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_SL g747 ( 
.A(n_685),
.B(n_518),
.Y(n_747)
);

INVx2_ASAP7_75t_L g748 ( 
.A(n_667),
.Y(n_748)
);

CKINVDCx8_ASAP7_75t_R g749 ( 
.A(n_691),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_672),
.Y(n_750)
);

AOI21xp5_ASAP7_75t_L g751 ( 
.A1(n_694),
.A2(n_630),
.B(n_661),
.Y(n_751)
);

CKINVDCx5p33_ASAP7_75t_R g752 ( 
.A(n_707),
.Y(n_752)
);

INVx3_ASAP7_75t_L g753 ( 
.A(n_631),
.Y(n_753)
);

HB1xp67_ASAP7_75t_L g754 ( 
.A(n_631),
.Y(n_754)
);

AND2x2_ASAP7_75t_L g755 ( 
.A(n_675),
.B(n_406),
.Y(n_755)
);

AOI21xp5_ASAP7_75t_L g756 ( 
.A1(n_634),
.A2(n_518),
.B(n_376),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_SL g757 ( 
.A(n_693),
.B(n_166),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_L g758 ( 
.A(n_677),
.B(n_406),
.Y(n_758)
);

HB1xp67_ASAP7_75t_L g759 ( 
.A(n_696),
.Y(n_759)
);

NOR3xp33_ASAP7_75t_SL g760 ( 
.A(n_659),
.B(n_171),
.C(n_169),
.Y(n_760)
);

OR2x6_ASAP7_75t_L g761 ( 
.A(n_704),
.B(n_406),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_680),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_701),
.B(n_415),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_L g764 ( 
.A(n_709),
.B(n_415),
.Y(n_764)
);

OAI22xp5_ASAP7_75t_L g765 ( 
.A1(n_698),
.A2(n_171),
.B1(n_174),
.B2(n_175),
.Y(n_765)
);

BUFx3_ASAP7_75t_L g766 ( 
.A(n_616),
.Y(n_766)
);

INVx2_ASAP7_75t_L g767 ( 
.A(n_688),
.Y(n_767)
);

BUFx6f_ASAP7_75t_L g768 ( 
.A(n_696),
.Y(n_768)
);

NOR2xp33_ASAP7_75t_L g769 ( 
.A(n_622),
.B(n_174),
.Y(n_769)
);

AOI22xp5_ASAP7_75t_L g770 ( 
.A1(n_687),
.A2(n_270),
.B1(n_217),
.B2(n_219),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_645),
.Y(n_771)
);

OAI22xp5_ASAP7_75t_L g772 ( 
.A1(n_689),
.A2(n_175),
.B1(n_277),
.B2(n_278),
.Y(n_772)
);

A2O1A1Ixp33_ASAP7_75t_L g773 ( 
.A1(n_637),
.A2(n_415),
.B(n_277),
.C(n_278),
.Y(n_773)
);

INVx2_ASAP7_75t_L g774 ( 
.A(n_688),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_SL g775 ( 
.A(n_647),
.B(n_279),
.Y(n_775)
);

AOI21xp5_ASAP7_75t_L g776 ( 
.A1(n_674),
.A2(n_376),
.B(n_374),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_L g777 ( 
.A(n_639),
.B(n_384),
.Y(n_777)
);

HB1xp67_ASAP7_75t_L g778 ( 
.A(n_696),
.Y(n_778)
);

NOR2xp33_ASAP7_75t_L g779 ( 
.A(n_654),
.B(n_279),
.Y(n_779)
);

AOI22xp5_ASAP7_75t_L g780 ( 
.A1(n_729),
.A2(n_752),
.B1(n_755),
.B2(n_730),
.Y(n_780)
);

BUFx8_ASAP7_75t_L g781 ( 
.A(n_726),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_L g782 ( 
.A(n_736),
.B(n_692),
.Y(n_782)
);

NAND3xp33_ASAP7_75t_SL g783 ( 
.A(n_717),
.B(n_280),
.C(n_224),
.Y(n_783)
);

CKINVDCx11_ASAP7_75t_R g784 ( 
.A(n_749),
.Y(n_784)
);

AOI21xp5_ASAP7_75t_L g785 ( 
.A1(n_751),
.A2(n_620),
.B(n_674),
.Y(n_785)
);

AOI21xp5_ASAP7_75t_L g786 ( 
.A1(n_732),
.A2(n_657),
.B(n_629),
.Y(n_786)
);

O2A1O1Ixp5_ASAP7_75t_L g787 ( 
.A1(n_775),
.A2(n_700),
.B(n_708),
.C(n_636),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_762),
.Y(n_788)
);

BUFx2_ASAP7_75t_L g789 ( 
.A(n_737),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_739),
.Y(n_790)
);

AOI21xp5_ASAP7_75t_L g791 ( 
.A1(n_716),
.A2(n_733),
.B(n_738),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_771),
.B(n_663),
.Y(n_792)
);

AO31x2_ASAP7_75t_L g793 ( 
.A1(n_773),
.A2(n_679),
.A3(n_676),
.B(n_618),
.Y(n_793)
);

OR2x2_ASAP7_75t_L g794 ( 
.A(n_729),
.B(n_700),
.Y(n_794)
);

OA21x2_ASAP7_75t_L g795 ( 
.A1(n_746),
.A2(n_623),
.B(n_624),
.Y(n_795)
);

INVx3_ASAP7_75t_SL g796 ( 
.A(n_713),
.Y(n_796)
);

OAI22xp33_ASAP7_75t_L g797 ( 
.A1(n_711),
.A2(n_766),
.B1(n_761),
.B2(n_757),
.Y(n_797)
);

AO22x1_ASAP7_75t_L g798 ( 
.A1(n_734),
.A2(n_280),
.B1(n_226),
.B2(n_228),
.Y(n_798)
);

INVx2_ASAP7_75t_L g799 ( 
.A(n_724),
.Y(n_799)
);

AOI21xp5_ASAP7_75t_L g800 ( 
.A1(n_719),
.A2(n_635),
.B(n_636),
.Y(n_800)
);

BUFx2_ASAP7_75t_L g801 ( 
.A(n_737),
.Y(n_801)
);

A2O1A1Ixp33_ASAP7_75t_L g802 ( 
.A1(n_710),
.A2(n_686),
.B(n_695),
.C(n_623),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_721),
.Y(n_803)
);

INVx2_ASAP7_75t_L g804 ( 
.A(n_723),
.Y(n_804)
);

INVx1_ASAP7_75t_SL g805 ( 
.A(n_715),
.Y(n_805)
);

CKINVDCx5p33_ASAP7_75t_R g806 ( 
.A(n_710),
.Y(n_806)
);

AOI221xp5_ASAP7_75t_SL g807 ( 
.A1(n_731),
.A2(n_708),
.B1(n_673),
.B2(n_681),
.C(n_705),
.Y(n_807)
);

AOI21xp5_ASAP7_75t_L g808 ( 
.A1(n_777),
.A2(n_613),
.B(n_619),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_735),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_740),
.Y(n_810)
);

NAND2xp33_ASAP7_75t_L g811 ( 
.A(n_718),
.B(n_696),
.Y(n_811)
);

AOI21xp5_ASAP7_75t_L g812 ( 
.A1(n_756),
.A2(n_628),
.B(n_706),
.Y(n_812)
);

BUFx2_ASAP7_75t_L g813 ( 
.A(n_713),
.Y(n_813)
);

INVx2_ASAP7_75t_SL g814 ( 
.A(n_728),
.Y(n_814)
);

INVx1_ASAP7_75t_SL g815 ( 
.A(n_754),
.Y(n_815)
);

AOI21xp5_ASAP7_75t_L g816 ( 
.A1(n_712),
.A2(n_640),
.B(n_669),
.Y(n_816)
);

BUFx10_ASAP7_75t_L g817 ( 
.A(n_769),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_750),
.Y(n_818)
);

AOI21xp5_ASAP7_75t_L g819 ( 
.A1(n_720),
.A2(n_678),
.B(n_684),
.Y(n_819)
);

OAI21x1_ASAP7_75t_L g820 ( 
.A1(n_776),
.A2(n_656),
.B(n_653),
.Y(n_820)
);

AOI21x1_ASAP7_75t_L g821 ( 
.A1(n_741),
.A2(n_666),
.B(n_658),
.Y(n_821)
);

INVx2_ASAP7_75t_L g822 ( 
.A(n_748),
.Y(n_822)
);

AOI21xp5_ASAP7_75t_L g823 ( 
.A1(n_745),
.A2(n_763),
.B(n_758),
.Y(n_823)
);

O2A1O1Ixp33_ASAP7_75t_L g824 ( 
.A1(n_743),
.A2(n_703),
.B(n_697),
.C(n_690),
.Y(n_824)
);

OAI21x1_ASAP7_75t_L g825 ( 
.A1(n_747),
.A2(n_702),
.B(n_642),
.Y(n_825)
);

OAI221xp5_ASAP7_75t_L g826 ( 
.A1(n_761),
.A2(n_703),
.B1(n_697),
.B2(n_273),
.C(n_268),
.Y(n_826)
);

OAI21x1_ASAP7_75t_L g827 ( 
.A1(n_727),
.A2(n_648),
.B(n_381),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_L g828 ( 
.A(n_779),
.B(n_386),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_L g829 ( 
.A(n_779),
.B(n_386),
.Y(n_829)
);

OAI22xp5_ASAP7_75t_L g830 ( 
.A1(n_714),
.A2(n_257),
.B1(n_236),
.B2(n_238),
.Y(n_830)
);

AO31x2_ASAP7_75t_L g831 ( 
.A1(n_722),
.A2(n_388),
.A3(n_381),
.B(n_380),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_L g832 ( 
.A(n_767),
.B(n_388),
.Y(n_832)
);

OAI21x1_ASAP7_75t_L g833 ( 
.A1(n_764),
.A2(n_381),
.B(n_97),
.Y(n_833)
);

NOR2xp33_ASAP7_75t_SL g834 ( 
.A(n_754),
.B(n_222),
.Y(n_834)
);

AO31x2_ASAP7_75t_L g835 ( 
.A1(n_722),
.A2(n_414),
.A3(n_412),
.B(n_411),
.Y(n_835)
);

INVxp67_ASAP7_75t_L g836 ( 
.A(n_761),
.Y(n_836)
);

INVx2_ASAP7_75t_SL g837 ( 
.A(n_759),
.Y(n_837)
);

AND2x4_ASAP7_75t_L g838 ( 
.A(n_744),
.B(n_55),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_774),
.Y(n_839)
);

AOI22xp5_ASAP7_75t_L g840 ( 
.A1(n_714),
.A2(n_262),
.B1(n_240),
.B2(n_241),
.Y(n_840)
);

NAND2x1p5_ASAP7_75t_L g841 ( 
.A(n_718),
.B(n_408),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_SL g842 ( 
.A(n_765),
.B(n_239),
.Y(n_842)
);

NOR2xp33_ASAP7_75t_L g843 ( 
.A(n_772),
.B(n_246),
.Y(n_843)
);

CKINVDCx5p33_ASAP7_75t_R g844 ( 
.A(n_784),
.Y(n_844)
);

INVx2_ASAP7_75t_L g845 ( 
.A(n_822),
.Y(n_845)
);

INVx2_ASAP7_75t_L g846 ( 
.A(n_804),
.Y(n_846)
);

AOI22xp33_ASAP7_75t_SL g847 ( 
.A1(n_806),
.A2(n_760),
.B1(n_742),
.B2(n_260),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_788),
.Y(n_848)
);

CKINVDCx5p33_ASAP7_75t_R g849 ( 
.A(n_781),
.Y(n_849)
);

CKINVDCx11_ASAP7_75t_R g850 ( 
.A(n_796),
.Y(n_850)
);

AOI22xp33_ASAP7_75t_L g851 ( 
.A1(n_783),
.A2(n_778),
.B1(n_759),
.B2(n_408),
.Y(n_851)
);

HB1xp67_ASAP7_75t_L g852 ( 
.A(n_815),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_809),
.Y(n_853)
);

AOI22xp5_ASAP7_75t_L g854 ( 
.A1(n_780),
.A2(n_770),
.B1(n_760),
.B2(n_255),
.Y(n_854)
);

AOI22xp33_ASAP7_75t_L g855 ( 
.A1(n_817),
.A2(n_778),
.B1(n_408),
.B2(n_412),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_810),
.Y(n_856)
);

AOI22xp33_ASAP7_75t_L g857 ( 
.A1(n_843),
.A2(n_753),
.B1(n_725),
.B2(n_275),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_818),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_803),
.Y(n_859)
);

INVx2_ASAP7_75t_L g860 ( 
.A(n_799),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_790),
.Y(n_861)
);

INVx1_ASAP7_75t_SL g862 ( 
.A(n_805),
.Y(n_862)
);

AOI22xp5_ASAP7_75t_L g863 ( 
.A1(n_797),
.A2(n_252),
.B1(n_276),
.B2(n_753),
.Y(n_863)
);

AOI22xp33_ASAP7_75t_L g864 ( 
.A1(n_794),
.A2(n_725),
.B1(n_718),
.B2(n_768),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_839),
.Y(n_865)
);

AOI22xp33_ASAP7_75t_L g866 ( 
.A1(n_838),
.A2(n_768),
.B1(n_718),
.B2(n_414),
.Y(n_866)
);

AOI22xp33_ASAP7_75t_SL g867 ( 
.A1(n_817),
.A2(n_742),
.B1(n_768),
.B2(n_8),
.Y(n_867)
);

BUFx3_ASAP7_75t_L g868 ( 
.A(n_781),
.Y(n_868)
);

INVxp67_ASAP7_75t_SL g869 ( 
.A(n_811),
.Y(n_869)
);

BUFx3_ASAP7_75t_L g870 ( 
.A(n_789),
.Y(n_870)
);

CKINVDCx11_ASAP7_75t_R g871 ( 
.A(n_805),
.Y(n_871)
);

BUFx10_ASAP7_75t_L g872 ( 
.A(n_814),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_832),
.Y(n_873)
);

BUFx10_ASAP7_75t_L g874 ( 
.A(n_838),
.Y(n_874)
);

INVx8_ASAP7_75t_L g875 ( 
.A(n_815),
.Y(n_875)
);

INVx3_ASAP7_75t_SL g876 ( 
.A(n_837),
.Y(n_876)
);

INVx6_ASAP7_75t_L g877 ( 
.A(n_801),
.Y(n_877)
);

INVx1_ASAP7_75t_SL g878 ( 
.A(n_813),
.Y(n_878)
);

BUFx6f_ASAP7_75t_L g879 ( 
.A(n_841),
.Y(n_879)
);

CKINVDCx20_ASAP7_75t_R g880 ( 
.A(n_836),
.Y(n_880)
);

INVx1_ASAP7_75t_SL g881 ( 
.A(n_834),
.Y(n_881)
);

CKINVDCx11_ASAP7_75t_R g882 ( 
.A(n_830),
.Y(n_882)
);

BUFx8_ASAP7_75t_L g883 ( 
.A(n_834),
.Y(n_883)
);

BUFx12f_ASAP7_75t_L g884 ( 
.A(n_841),
.Y(n_884)
);

BUFx2_ASAP7_75t_L g885 ( 
.A(n_832),
.Y(n_885)
);

INVx5_ASAP7_75t_L g886 ( 
.A(n_826),
.Y(n_886)
);

INVx6_ASAP7_75t_L g887 ( 
.A(n_798),
.Y(n_887)
);

INVx2_ASAP7_75t_L g888 ( 
.A(n_792),
.Y(n_888)
);

BUFx4_ASAP7_75t_R g889 ( 
.A(n_840),
.Y(n_889)
);

INVx2_ASAP7_75t_L g890 ( 
.A(n_821),
.Y(n_890)
);

AOI22xp5_ASAP7_75t_L g891 ( 
.A1(n_842),
.A2(n_768),
.B1(n_414),
.B2(n_412),
.Y(n_891)
);

OAI22xp5_ASAP7_75t_L g892 ( 
.A1(n_782),
.A2(n_742),
.B1(n_414),
.B2(n_412),
.Y(n_892)
);

CKINVDCx6p67_ASAP7_75t_R g893 ( 
.A(n_828),
.Y(n_893)
);

AOI22xp33_ASAP7_75t_L g894 ( 
.A1(n_828),
.A2(n_414),
.B1(n_412),
.B2(n_411),
.Y(n_894)
);

CKINVDCx6p67_ASAP7_75t_R g895 ( 
.A(n_829),
.Y(n_895)
);

CKINVDCx5p33_ASAP7_75t_R g896 ( 
.A(n_830),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_829),
.Y(n_897)
);

INVx6_ASAP7_75t_L g898 ( 
.A(n_824),
.Y(n_898)
);

OAI22xp33_ASAP7_75t_L g899 ( 
.A1(n_791),
.A2(n_742),
.B1(n_414),
.B2(n_412),
.Y(n_899)
);

OAI22xp5_ASAP7_75t_L g900 ( 
.A1(n_802),
.A2(n_414),
.B1(n_412),
.B2(n_411),
.Y(n_900)
);

BUFx4f_ASAP7_75t_SL g901 ( 
.A(n_787),
.Y(n_901)
);

CKINVDCx20_ASAP7_75t_R g902 ( 
.A(n_819),
.Y(n_902)
);

AOI22xp33_ASAP7_75t_SL g903 ( 
.A1(n_785),
.A2(n_6),
.B1(n_7),
.B2(n_9),
.Y(n_903)
);

INVx6_ASAP7_75t_L g904 ( 
.A(n_807),
.Y(n_904)
);

INVx2_ASAP7_75t_L g905 ( 
.A(n_795),
.Y(n_905)
);

CKINVDCx6p67_ASAP7_75t_R g906 ( 
.A(n_807),
.Y(n_906)
);

AOI22xp33_ASAP7_75t_L g907 ( 
.A1(n_823),
.A2(n_411),
.B1(n_409),
.B2(n_722),
.Y(n_907)
);

AOI22xp33_ASAP7_75t_L g908 ( 
.A1(n_786),
.A2(n_411),
.B1(n_409),
.B2(n_11),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_831),
.Y(n_909)
);

NAND2x1p5_ASAP7_75t_L g910 ( 
.A(n_827),
.B(n_409),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_909),
.Y(n_911)
);

AOI22xp5_ASAP7_75t_L g912 ( 
.A1(n_896),
.A2(n_882),
.B1(n_893),
.B2(n_895),
.Y(n_912)
);

INVx4_ASAP7_75t_L g913 ( 
.A(n_898),
.Y(n_913)
);

OA21x2_ASAP7_75t_L g914 ( 
.A1(n_905),
.A2(n_816),
.B(n_808),
.Y(n_914)
);

INVx2_ASAP7_75t_L g915 ( 
.A(n_890),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_L g916 ( 
.A(n_897),
.B(n_831),
.Y(n_916)
);

OR2x6_ASAP7_75t_L g917 ( 
.A(n_898),
.B(n_812),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_904),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_L g919 ( 
.A(n_888),
.B(n_831),
.Y(n_919)
);

BUFx3_ASAP7_75t_L g920 ( 
.A(n_902),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_L g921 ( 
.A(n_861),
.B(n_835),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_904),
.Y(n_922)
);

INVx2_ASAP7_75t_L g923 ( 
.A(n_904),
.Y(n_923)
);

INVx2_ASAP7_75t_L g924 ( 
.A(n_859),
.Y(n_924)
);

OA21x2_ASAP7_75t_L g925 ( 
.A1(n_907),
.A2(n_833),
.B(n_820),
.Y(n_925)
);

AOI22xp33_ASAP7_75t_SL g926 ( 
.A1(n_883),
.A2(n_800),
.B1(n_795),
.B2(n_825),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_906),
.Y(n_927)
);

AND2x2_ASAP7_75t_L g928 ( 
.A(n_867),
.B(n_835),
.Y(n_928)
);

HB1xp67_ASAP7_75t_L g929 ( 
.A(n_852),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_848),
.Y(n_930)
);

BUFx2_ASAP7_75t_L g931 ( 
.A(n_901),
.Y(n_931)
);

BUFx6f_ASAP7_75t_SL g932 ( 
.A(n_874),
.Y(n_932)
);

INVx1_ASAP7_75t_L g933 ( 
.A(n_853),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_856),
.Y(n_934)
);

INVx1_ASAP7_75t_L g935 ( 
.A(n_858),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_898),
.Y(n_936)
);

AND2x2_ASAP7_75t_L g937 ( 
.A(n_867),
.B(n_835),
.Y(n_937)
);

BUFx6f_ASAP7_75t_L g938 ( 
.A(n_910),
.Y(n_938)
);

INVx2_ASAP7_75t_L g939 ( 
.A(n_910),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_865),
.Y(n_940)
);

BUFx2_ASAP7_75t_L g941 ( 
.A(n_901),
.Y(n_941)
);

INVx1_ASAP7_75t_L g942 ( 
.A(n_846),
.Y(n_942)
);

INVx2_ASAP7_75t_L g943 ( 
.A(n_860),
.Y(n_943)
);

BUFx3_ASAP7_75t_L g944 ( 
.A(n_883),
.Y(n_944)
);

INVx1_ASAP7_75t_L g945 ( 
.A(n_873),
.Y(n_945)
);

AND2x2_ASAP7_75t_L g946 ( 
.A(n_847),
.B(n_793),
.Y(n_946)
);

OR2x2_ASAP7_75t_L g947 ( 
.A(n_852),
.B(n_793),
.Y(n_947)
);

BUFx3_ASAP7_75t_L g948 ( 
.A(n_875),
.Y(n_948)
);

INVx2_ASAP7_75t_L g949 ( 
.A(n_845),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_899),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_SL g951 ( 
.A(n_886),
.B(n_409),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_899),
.Y(n_952)
);

BUFx2_ASAP7_75t_L g953 ( 
.A(n_869),
.Y(n_953)
);

INVx5_ASAP7_75t_L g954 ( 
.A(n_886),
.Y(n_954)
);

INVx2_ASAP7_75t_L g955 ( 
.A(n_885),
.Y(n_955)
);

INVx2_ASAP7_75t_SL g956 ( 
.A(n_875),
.Y(n_956)
);

OAI21x1_ASAP7_75t_L g957 ( 
.A1(n_900),
.A2(n_793),
.B(n_411),
.Y(n_957)
);

OR2x2_ASAP7_75t_L g958 ( 
.A(n_955),
.B(n_862),
.Y(n_958)
);

A2O1A1Ixp33_ASAP7_75t_L g959 ( 
.A1(n_954),
.A2(n_886),
.B(n_908),
.C(n_903),
.Y(n_959)
);

HB1xp67_ASAP7_75t_L g960 ( 
.A(n_929),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_L g961 ( 
.A(n_955),
.B(n_870),
.Y(n_961)
);

AO21x2_ASAP7_75t_L g962 ( 
.A1(n_951),
.A2(n_892),
.B(n_863),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_L g963 ( 
.A(n_955),
.B(n_881),
.Y(n_963)
);

INVx4_ASAP7_75t_L g964 ( 
.A(n_913),
.Y(n_964)
);

OAI21x1_ASAP7_75t_L g965 ( 
.A1(n_957),
.A2(n_908),
.B(n_869),
.Y(n_965)
);

AND2x2_ASAP7_75t_L g966 ( 
.A(n_920),
.B(n_877),
.Y(n_966)
);

OAI21xp5_ASAP7_75t_L g967 ( 
.A1(n_951),
.A2(n_854),
.B(n_903),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_L g968 ( 
.A(n_929),
.B(n_877),
.Y(n_968)
);

A2O1A1Ixp33_ASAP7_75t_L g969 ( 
.A1(n_954),
.A2(n_886),
.B(n_847),
.C(n_866),
.Y(n_969)
);

AND2x2_ASAP7_75t_L g970 ( 
.A(n_946),
.B(n_877),
.Y(n_970)
);

AND2x4_ASAP7_75t_L g971 ( 
.A(n_924),
.B(n_879),
.Y(n_971)
);

OAI21xp5_ASAP7_75t_L g972 ( 
.A1(n_936),
.A2(n_857),
.B(n_851),
.Y(n_972)
);

AND2x2_ASAP7_75t_L g973 ( 
.A(n_946),
.B(n_924),
.Y(n_973)
);

AND2x4_ASAP7_75t_L g974 ( 
.A(n_924),
.B(n_879),
.Y(n_974)
);

AND2x4_ASAP7_75t_L g975 ( 
.A(n_930),
.B(n_879),
.Y(n_975)
);

AOI221xp5_ASAP7_75t_L g976 ( 
.A1(n_946),
.A2(n_878),
.B1(n_851),
.B2(n_875),
.C(n_880),
.Y(n_976)
);

AND2x2_ASAP7_75t_L g977 ( 
.A(n_947),
.B(n_871),
.Y(n_977)
);

AO32x2_ASAP7_75t_L g978 ( 
.A1(n_913),
.A2(n_889),
.A3(n_876),
.B1(n_887),
.B2(n_874),
.Y(n_978)
);

AND2x2_ASAP7_75t_L g979 ( 
.A(n_920),
.B(n_876),
.Y(n_979)
);

OR2x6_ASAP7_75t_L g980 ( 
.A(n_917),
.B(n_887),
.Y(n_980)
);

AND2x2_ASAP7_75t_L g981 ( 
.A(n_947),
.B(n_864),
.Y(n_981)
);

AND2x2_ASAP7_75t_L g982 ( 
.A(n_947),
.B(n_872),
.Y(n_982)
);

AND2x4_ASAP7_75t_L g983 ( 
.A(n_930),
.B(n_879),
.Y(n_983)
);

BUFx4f_ASAP7_75t_L g984 ( 
.A(n_927),
.Y(n_984)
);

HB1xp67_ASAP7_75t_L g985 ( 
.A(n_953),
.Y(n_985)
);

NOR2x1p5_ASAP7_75t_L g986 ( 
.A(n_944),
.B(n_868),
.Y(n_986)
);

AO32x2_ASAP7_75t_L g987 ( 
.A1(n_913),
.A2(n_887),
.A3(n_872),
.B1(n_855),
.B2(n_13),
.Y(n_987)
);

AO21x1_ASAP7_75t_L g988 ( 
.A1(n_936),
.A2(n_891),
.B(n_10),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_L g989 ( 
.A(n_945),
.B(n_844),
.Y(n_989)
);

AND2x2_ASAP7_75t_L g990 ( 
.A(n_928),
.B(n_855),
.Y(n_990)
);

O2A1O1Ixp33_ASAP7_75t_L g991 ( 
.A1(n_927),
.A2(n_894),
.B(n_10),
.C(n_12),
.Y(n_991)
);

A2O1A1Ixp33_ASAP7_75t_L g992 ( 
.A1(n_954),
.A2(n_920),
.B(n_953),
.C(n_922),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_L g993 ( 
.A(n_945),
.B(n_850),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_L g994 ( 
.A(n_920),
.B(n_849),
.Y(n_994)
);

AND2x2_ASAP7_75t_L g995 ( 
.A(n_928),
.B(n_894),
.Y(n_995)
);

OR2x6_ASAP7_75t_L g996 ( 
.A(n_917),
.B(n_884),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_L g997 ( 
.A(n_942),
.B(n_940),
.Y(n_997)
);

HB1xp67_ASAP7_75t_L g998 ( 
.A(n_953),
.Y(n_998)
);

OAI21xp5_ASAP7_75t_L g999 ( 
.A1(n_918),
.A2(n_86),
.B(n_161),
.Y(n_999)
);

AND2x2_ASAP7_75t_L g1000 ( 
.A(n_928),
.B(n_6),
.Y(n_1000)
);

OAI22xp5_ASAP7_75t_SL g1001 ( 
.A1(n_912),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_1001)
);

NOR2xp33_ASAP7_75t_L g1002 ( 
.A(n_918),
.B(n_16),
.Y(n_1002)
);

AND2x2_ASAP7_75t_L g1003 ( 
.A(n_931),
.B(n_16),
.Y(n_1003)
);

AND2x2_ASAP7_75t_L g1004 ( 
.A(n_973),
.B(n_914),
.Y(n_1004)
);

INVx2_ASAP7_75t_L g1005 ( 
.A(n_973),
.Y(n_1005)
);

INVx3_ASAP7_75t_L g1006 ( 
.A(n_971),
.Y(n_1006)
);

OR2x2_ASAP7_75t_L g1007 ( 
.A(n_960),
.B(n_911),
.Y(n_1007)
);

AND2x2_ASAP7_75t_L g1008 ( 
.A(n_970),
.B(n_911),
.Y(n_1008)
);

BUFx3_ASAP7_75t_L g1009 ( 
.A(n_984),
.Y(n_1009)
);

INVx2_ASAP7_75t_L g1010 ( 
.A(n_997),
.Y(n_1010)
);

AND2x4_ASAP7_75t_L g1011 ( 
.A(n_971),
.B(n_917),
.Y(n_1011)
);

AND2x2_ASAP7_75t_L g1012 ( 
.A(n_970),
.B(n_914),
.Y(n_1012)
);

NOR2x1p5_ASAP7_75t_L g1013 ( 
.A(n_964),
.B(n_944),
.Y(n_1013)
);

OR2x2_ASAP7_75t_L g1014 ( 
.A(n_985),
.B(n_914),
.Y(n_1014)
);

OR2x2_ASAP7_75t_L g1015 ( 
.A(n_998),
.B(n_914),
.Y(n_1015)
);

AND2x4_ASAP7_75t_L g1016 ( 
.A(n_971),
.B(n_917),
.Y(n_1016)
);

INVx1_ASAP7_75t_L g1017 ( 
.A(n_974),
.Y(n_1017)
);

INVx2_ASAP7_75t_L g1018 ( 
.A(n_974),
.Y(n_1018)
);

INVx1_ASAP7_75t_L g1019 ( 
.A(n_974),
.Y(n_1019)
);

AND2x2_ASAP7_75t_L g1020 ( 
.A(n_1000),
.B(n_937),
.Y(n_1020)
);

BUFx3_ASAP7_75t_L g1021 ( 
.A(n_984),
.Y(n_1021)
);

AOI22xp33_ASAP7_75t_L g1022 ( 
.A1(n_1001),
.A2(n_922),
.B1(n_931),
.B2(n_941),
.Y(n_1022)
);

INVx2_ASAP7_75t_L g1023 ( 
.A(n_975),
.Y(n_1023)
);

AND2x2_ASAP7_75t_L g1024 ( 
.A(n_1000),
.B(n_937),
.Y(n_1024)
);

AND2x2_ASAP7_75t_L g1025 ( 
.A(n_990),
.B(n_937),
.Y(n_1025)
);

HB1xp67_ASAP7_75t_L g1026 ( 
.A(n_982),
.Y(n_1026)
);

NAND2xp5_ASAP7_75t_L g1027 ( 
.A(n_982),
.B(n_933),
.Y(n_1027)
);

AND2x2_ASAP7_75t_L g1028 ( 
.A(n_990),
.B(n_914),
.Y(n_1028)
);

NOR2xp33_ASAP7_75t_L g1029 ( 
.A(n_963),
.B(n_913),
.Y(n_1029)
);

AND2x2_ASAP7_75t_L g1030 ( 
.A(n_995),
.B(n_926),
.Y(n_1030)
);

NOR2xp67_ASAP7_75t_L g1031 ( 
.A(n_964),
.B(n_954),
.Y(n_1031)
);

OAI33xp33_ASAP7_75t_L g1032 ( 
.A1(n_1007),
.A2(n_991),
.A3(n_958),
.B1(n_961),
.B2(n_968),
.B3(n_989),
.Y(n_1032)
);

OAI33xp33_ASAP7_75t_L g1033 ( 
.A1(n_1007),
.A2(n_935),
.A3(n_934),
.B1(n_933),
.B2(n_993),
.B3(n_940),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_L g1034 ( 
.A(n_1010),
.B(n_1025),
.Y(n_1034)
);

INVx1_ASAP7_75t_L g1035 ( 
.A(n_1005),
.Y(n_1035)
);

AOI22xp33_ASAP7_75t_L g1036 ( 
.A1(n_1022),
.A2(n_967),
.B1(n_980),
.B2(n_941),
.Y(n_1036)
);

BUFx2_ASAP7_75t_L g1037 ( 
.A(n_1006),
.Y(n_1037)
);

AND2x2_ASAP7_75t_L g1038 ( 
.A(n_1005),
.B(n_992),
.Y(n_1038)
);

HB1xp67_ASAP7_75t_L g1039 ( 
.A(n_1005),
.Y(n_1039)
);

INVx2_ASAP7_75t_L g1040 ( 
.A(n_1005),
.Y(n_1040)
);

INVx1_ASAP7_75t_L g1041 ( 
.A(n_1007),
.Y(n_1041)
);

AND2x2_ASAP7_75t_L g1042 ( 
.A(n_1004),
.B(n_992),
.Y(n_1042)
);

OAI21x1_ASAP7_75t_L g1043 ( 
.A1(n_1014),
.A2(n_965),
.B(n_957),
.Y(n_1043)
);

INVx1_ASAP7_75t_L g1044 ( 
.A(n_1010),
.Y(n_1044)
);

INVx1_ASAP7_75t_L g1045 ( 
.A(n_1010),
.Y(n_1045)
);

AOI22xp33_ASAP7_75t_L g1046 ( 
.A1(n_1022),
.A2(n_980),
.B1(n_931),
.B2(n_941),
.Y(n_1046)
);

AND2x2_ASAP7_75t_L g1047 ( 
.A(n_1004),
.B(n_981),
.Y(n_1047)
);

AND2x2_ASAP7_75t_L g1048 ( 
.A(n_1004),
.B(n_981),
.Y(n_1048)
);

AND2x2_ASAP7_75t_L g1049 ( 
.A(n_1004),
.B(n_995),
.Y(n_1049)
);

BUFx2_ASAP7_75t_L g1050 ( 
.A(n_1006),
.Y(n_1050)
);

AND2x2_ASAP7_75t_L g1051 ( 
.A(n_1012),
.B(n_980),
.Y(n_1051)
);

INVx2_ASAP7_75t_L g1052 ( 
.A(n_1014),
.Y(n_1052)
);

INVx2_ASAP7_75t_L g1053 ( 
.A(n_1014),
.Y(n_1053)
);

INVxp67_ASAP7_75t_L g1054 ( 
.A(n_1026),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_L g1055 ( 
.A(n_1047),
.B(n_1027),
.Y(n_1055)
);

AND2x2_ASAP7_75t_L g1056 ( 
.A(n_1047),
.B(n_1018),
.Y(n_1056)
);

INVx1_ASAP7_75t_L g1057 ( 
.A(n_1041),
.Y(n_1057)
);

INVx2_ASAP7_75t_SL g1058 ( 
.A(n_1037),
.Y(n_1058)
);

OR2x6_ASAP7_75t_L g1059 ( 
.A(n_1043),
.B(n_980),
.Y(n_1059)
);

NOR4xp25_ASAP7_75t_SL g1060 ( 
.A(n_1037),
.B(n_969),
.C(n_959),
.D(n_1019),
.Y(n_1060)
);

INVx2_ASAP7_75t_L g1061 ( 
.A(n_1040),
.Y(n_1061)
);

INVx2_ASAP7_75t_L g1062 ( 
.A(n_1040),
.Y(n_1062)
);

AOI22xp33_ASAP7_75t_SL g1063 ( 
.A1(n_1042),
.A2(n_1030),
.B1(n_984),
.B2(n_954),
.Y(n_1063)
);

INVx1_ASAP7_75t_L g1064 ( 
.A(n_1041),
.Y(n_1064)
);

HB1xp67_ASAP7_75t_L g1065 ( 
.A(n_1054),
.Y(n_1065)
);

AND2x2_ASAP7_75t_L g1066 ( 
.A(n_1047),
.B(n_1018),
.Y(n_1066)
);

AND2x4_ASAP7_75t_L g1067 ( 
.A(n_1051),
.B(n_1031),
.Y(n_1067)
);

OR2x2_ASAP7_75t_L g1068 ( 
.A(n_1034),
.B(n_1027),
.Y(n_1068)
);

NAND2x1_ASAP7_75t_L g1069 ( 
.A(n_1067),
.B(n_1050),
.Y(n_1069)
);

HB1xp67_ASAP7_75t_L g1070 ( 
.A(n_1065),
.Y(n_1070)
);

INVx1_ASAP7_75t_L g1071 ( 
.A(n_1057),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_L g1072 ( 
.A(n_1055),
.B(n_1048),
.Y(n_1072)
);

NAND2xp5_ASAP7_75t_L g1073 ( 
.A(n_1057),
.B(n_1048),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_L g1074 ( 
.A(n_1068),
.B(n_1048),
.Y(n_1074)
);

INVx1_ASAP7_75t_L g1075 ( 
.A(n_1064),
.Y(n_1075)
);

INVx4_ASAP7_75t_L g1076 ( 
.A(n_1067),
.Y(n_1076)
);

INVx1_ASAP7_75t_L g1077 ( 
.A(n_1064),
.Y(n_1077)
);

NOR3xp33_ASAP7_75t_L g1078 ( 
.A(n_1070),
.B(n_1032),
.C(n_994),
.Y(n_1078)
);

AND2x2_ASAP7_75t_L g1079 ( 
.A(n_1076),
.B(n_1067),
.Y(n_1079)
);

NAND2xp5_ASAP7_75t_L g1080 ( 
.A(n_1071),
.B(n_1068),
.Y(n_1080)
);

OR2x2_ASAP7_75t_L g1081 ( 
.A(n_1074),
.B(n_1034),
.Y(n_1081)
);

INVx1_ASAP7_75t_L g1082 ( 
.A(n_1075),
.Y(n_1082)
);

AND2x4_ASAP7_75t_L g1083 ( 
.A(n_1079),
.B(n_1076),
.Y(n_1083)
);

NOR2xp33_ASAP7_75t_L g1084 ( 
.A(n_1078),
.B(n_1072),
.Y(n_1084)
);

INVx2_ASAP7_75t_SL g1085 ( 
.A(n_1082),
.Y(n_1085)
);

INVxp67_ASAP7_75t_SL g1086 ( 
.A(n_1080),
.Y(n_1086)
);

AOI22xp5_ASAP7_75t_L g1087 ( 
.A1(n_1080),
.A2(n_1032),
.B1(n_1063),
.B2(n_1067),
.Y(n_1087)
);

INVxp67_ASAP7_75t_SL g1088 ( 
.A(n_1081),
.Y(n_1088)
);

OAI22xp5_ASAP7_75t_L g1089 ( 
.A1(n_1078),
.A2(n_1060),
.B1(n_1036),
.B2(n_1069),
.Y(n_1089)
);

AOI22xp5_ASAP7_75t_L g1090 ( 
.A1(n_1078),
.A2(n_1059),
.B1(n_1033),
.B2(n_1042),
.Y(n_1090)
);

AOI221xp5_ASAP7_75t_L g1091 ( 
.A1(n_1078),
.A2(n_1002),
.B1(n_1033),
.B2(n_1077),
.C(n_1073),
.Y(n_1091)
);

NOR2xp33_ASAP7_75t_SL g1092 ( 
.A(n_1079),
.B(n_944),
.Y(n_1092)
);

AND2x2_ASAP7_75t_L g1093 ( 
.A(n_1079),
.B(n_1056),
.Y(n_1093)
);

NAND2xp5_ASAP7_75t_L g1094 ( 
.A(n_1078),
.B(n_1073),
.Y(n_1094)
);

INVxp33_ASAP7_75t_L g1095 ( 
.A(n_1092),
.Y(n_1095)
);

NAND2xp5_ASAP7_75t_L g1096 ( 
.A(n_1086),
.B(n_1061),
.Y(n_1096)
);

INVxp67_ASAP7_75t_SL g1097 ( 
.A(n_1088),
.Y(n_1097)
);

OR2x2_ASAP7_75t_L g1098 ( 
.A(n_1094),
.B(n_1056),
.Y(n_1098)
);

NAND2xp5_ASAP7_75t_L g1099 ( 
.A(n_1085),
.B(n_1084),
.Y(n_1099)
);

NAND2xp5_ASAP7_75t_SL g1100 ( 
.A(n_1089),
.B(n_1058),
.Y(n_1100)
);

OAI222xp33_ASAP7_75t_L g1101 ( 
.A1(n_1090),
.A2(n_1059),
.B1(n_1046),
.B2(n_1058),
.C1(n_912),
.C2(n_1054),
.Y(n_1101)
);

AND2x4_ASAP7_75t_L g1102 ( 
.A(n_1083),
.B(n_986),
.Y(n_1102)
);

OAI22xp5_ASAP7_75t_L g1103 ( 
.A1(n_1087),
.A2(n_1002),
.B1(n_959),
.B2(n_944),
.Y(n_1103)
);

INVx2_ASAP7_75t_L g1104 ( 
.A(n_1083),
.Y(n_1104)
);

NOR4xp25_ASAP7_75t_SL g1105 ( 
.A(n_1091),
.B(n_1050),
.C(n_969),
.D(n_976),
.Y(n_1105)
);

INVx1_ASAP7_75t_L g1106 ( 
.A(n_1093),
.Y(n_1106)
);

NAND3xp33_ASAP7_75t_L g1107 ( 
.A(n_1091),
.B(n_1003),
.C(n_972),
.Y(n_1107)
);

INVx1_ASAP7_75t_L g1108 ( 
.A(n_1085),
.Y(n_1108)
);

OAI21xp5_ASAP7_75t_SL g1109 ( 
.A1(n_1089),
.A2(n_977),
.B(n_979),
.Y(n_1109)
);

AOI21xp5_ASAP7_75t_L g1110 ( 
.A1(n_1089),
.A2(n_1059),
.B(n_999),
.Y(n_1110)
);

AND2x2_ASAP7_75t_L g1111 ( 
.A(n_1083),
.B(n_1066),
.Y(n_1111)
);

INVx2_ASAP7_75t_L g1112 ( 
.A(n_1104),
.Y(n_1112)
);

NAND2xp5_ASAP7_75t_L g1113 ( 
.A(n_1097),
.B(n_1061),
.Y(n_1113)
);

XOR2x2_ASAP7_75t_L g1114 ( 
.A(n_1100),
.B(n_977),
.Y(n_1114)
);

AND2x2_ASAP7_75t_L g1115 ( 
.A(n_1102),
.B(n_1066),
.Y(n_1115)
);

INVx1_ASAP7_75t_L g1116 ( 
.A(n_1106),
.Y(n_1116)
);

OAI21xp5_ASAP7_75t_SL g1117 ( 
.A1(n_1109),
.A2(n_966),
.B(n_1042),
.Y(n_1117)
);

OAI211xp5_ASAP7_75t_SL g1118 ( 
.A1(n_1099),
.A2(n_926),
.B(n_20),
.C(n_21),
.Y(n_1118)
);

OAI22xp5_ASAP7_75t_L g1119 ( 
.A1(n_1107),
.A2(n_1059),
.B1(n_1038),
.B2(n_1013),
.Y(n_1119)
);

INVx2_ASAP7_75t_L g1120 ( 
.A(n_1111),
.Y(n_1120)
);

AOI22xp5_ASAP7_75t_L g1121 ( 
.A1(n_1103),
.A2(n_1059),
.B1(n_1013),
.B2(n_1009),
.Y(n_1121)
);

INVx1_ASAP7_75t_L g1122 ( 
.A(n_1108),
.Y(n_1122)
);

AND2x2_ASAP7_75t_L g1123 ( 
.A(n_1102),
.B(n_1049),
.Y(n_1123)
);

INVx1_ASAP7_75t_L g1124 ( 
.A(n_1096),
.Y(n_1124)
);

OAI21xp5_ASAP7_75t_L g1125 ( 
.A1(n_1103),
.A2(n_1038),
.B(n_1031),
.Y(n_1125)
);

XOR2x2_ASAP7_75t_L g1126 ( 
.A(n_1110),
.B(n_1098),
.Y(n_1126)
);

INVx2_ASAP7_75t_L g1127 ( 
.A(n_1096),
.Y(n_1127)
);

INVxp33_ASAP7_75t_L g1128 ( 
.A(n_1095),
.Y(n_1128)
);

INVx1_ASAP7_75t_L g1129 ( 
.A(n_1105),
.Y(n_1129)
);

NAND2xp5_ASAP7_75t_L g1130 ( 
.A(n_1101),
.B(n_1062),
.Y(n_1130)
);

INVx1_ASAP7_75t_L g1131 ( 
.A(n_1112),
.Y(n_1131)
);

OAI211xp5_ASAP7_75t_SL g1132 ( 
.A1(n_1129),
.A2(n_1062),
.B(n_1053),
.C(n_1052),
.Y(n_1132)
);

NOR4xp25_ASAP7_75t_L g1133 ( 
.A(n_1112),
.B(n_1038),
.C(n_1052),
.D(n_1053),
.Y(n_1133)
);

NOR2xp67_ASAP7_75t_L g1134 ( 
.A(n_1127),
.B(n_1122),
.Y(n_1134)
);

NOR2xp67_ASAP7_75t_L g1135 ( 
.A(n_1113),
.B(n_17),
.Y(n_1135)
);

NOR3xp33_ASAP7_75t_L g1136 ( 
.A(n_1116),
.B(n_913),
.C(n_956),
.Y(n_1136)
);

NOR3x1_ASAP7_75t_L g1137 ( 
.A(n_1124),
.B(n_956),
.C(n_1017),
.Y(n_1137)
);

INVx1_ASAP7_75t_L g1138 ( 
.A(n_1113),
.Y(n_1138)
);

NOR4xp25_ASAP7_75t_L g1139 ( 
.A(n_1120),
.B(n_1053),
.C(n_1052),
.D(n_1045),
.Y(n_1139)
);

O2A1O1Ixp33_ASAP7_75t_SL g1140 ( 
.A1(n_1118),
.A2(n_956),
.B(n_1039),
.C(n_1026),
.Y(n_1140)
);

NOR2x1_ASAP7_75t_L g1141 ( 
.A(n_1118),
.B(n_1013),
.Y(n_1141)
);

AOI21x1_ASAP7_75t_L g1142 ( 
.A1(n_1130),
.A2(n_1031),
.B(n_988),
.Y(n_1142)
);

NAND2xp33_ASAP7_75t_SL g1143 ( 
.A(n_1128),
.B(n_932),
.Y(n_1143)
);

NAND3xp33_ASAP7_75t_SL g1144 ( 
.A(n_1128),
.B(n_923),
.C(n_1030),
.Y(n_1144)
);

NOR2x1_ASAP7_75t_L g1145 ( 
.A(n_1130),
.B(n_1009),
.Y(n_1145)
);

AOI22xp33_ASAP7_75t_SL g1146 ( 
.A1(n_1119),
.A2(n_1009),
.B1(n_1021),
.B2(n_1030),
.Y(n_1146)
);

NAND2xp5_ASAP7_75t_L g1147 ( 
.A(n_1126),
.B(n_1049),
.Y(n_1147)
);

AOI221xp5_ASAP7_75t_SL g1148 ( 
.A1(n_1147),
.A2(n_1125),
.B1(n_1115),
.B2(n_1123),
.C(n_1114),
.Y(n_1148)
);

AOI221x1_ASAP7_75t_L g1149 ( 
.A1(n_1131),
.A2(n_1121),
.B1(n_1117),
.B2(n_1045),
.C(n_1044),
.Y(n_1149)
);

INVx1_ASAP7_75t_L g1150 ( 
.A(n_1135),
.Y(n_1150)
);

NOR2x1p5_ASAP7_75t_L g1151 ( 
.A(n_1138),
.B(n_1009),
.Y(n_1151)
);

INVxp67_ASAP7_75t_L g1152 ( 
.A(n_1145),
.Y(n_1152)
);

NOR2xp33_ASAP7_75t_SL g1153 ( 
.A(n_1134),
.B(n_1021),
.Y(n_1153)
);

NAND4xp25_ASAP7_75t_L g1154 ( 
.A(n_1146),
.B(n_1021),
.C(n_948),
.D(n_1029),
.Y(n_1154)
);

NAND2xp5_ASAP7_75t_SL g1155 ( 
.A(n_1141),
.B(n_1021),
.Y(n_1155)
);

NAND2xp5_ASAP7_75t_L g1156 ( 
.A(n_1137),
.B(n_1049),
.Y(n_1156)
);

OAI211xp5_ASAP7_75t_SL g1157 ( 
.A1(n_1140),
.A2(n_1136),
.B(n_1143),
.C(n_1132),
.Y(n_1157)
);

AOI222xp33_ASAP7_75t_L g1158 ( 
.A1(n_1144),
.A2(n_1030),
.B1(n_1024),
.B2(n_1020),
.C1(n_954),
.C2(n_1025),
.Y(n_1158)
);

OAI21xp5_ASAP7_75t_L g1159 ( 
.A1(n_1142),
.A2(n_1029),
.B(n_954),
.Y(n_1159)
);

NAND3xp33_ASAP7_75t_SL g1160 ( 
.A(n_1133),
.B(n_923),
.C(n_1051),
.Y(n_1160)
);

OR2x2_ASAP7_75t_L g1161 ( 
.A(n_1139),
.B(n_1039),
.Y(n_1161)
);

O2A1O1Ixp33_ASAP7_75t_L g1162 ( 
.A1(n_1140),
.A2(n_923),
.B(n_20),
.C(n_21),
.Y(n_1162)
);

NAND3xp33_ASAP7_75t_SL g1163 ( 
.A(n_1146),
.B(n_1051),
.C(n_978),
.Y(n_1163)
);

OAI211xp5_ASAP7_75t_SL g1164 ( 
.A1(n_1146),
.A2(n_17),
.B(n_22),
.C(n_23),
.Y(n_1164)
);

OAI21xp5_ASAP7_75t_L g1165 ( 
.A1(n_1135),
.A2(n_954),
.B(n_1043),
.Y(n_1165)
);

AOI221xp5_ASAP7_75t_L g1166 ( 
.A1(n_1140),
.A2(n_1044),
.B1(n_1025),
.B2(n_1019),
.C(n_1017),
.Y(n_1166)
);

AOI221xp5_ASAP7_75t_L g1167 ( 
.A1(n_1140),
.A2(n_1017),
.B1(n_1019),
.B2(n_1035),
.C(n_1020),
.Y(n_1167)
);

OAI221xp5_ASAP7_75t_L g1168 ( 
.A1(n_1146),
.A2(n_948),
.B1(n_996),
.B2(n_917),
.C(n_964),
.Y(n_1168)
);

OAI221xp5_ASAP7_75t_L g1169 ( 
.A1(n_1146),
.A2(n_948),
.B1(n_996),
.B2(n_917),
.C(n_1035),
.Y(n_1169)
);

INVx1_ASAP7_75t_L g1170 ( 
.A(n_1131),
.Y(n_1170)
);

AOI211xp5_ASAP7_75t_L g1171 ( 
.A1(n_1140),
.A2(n_23),
.B(n_26),
.C(n_27),
.Y(n_1171)
);

NAND3xp33_ASAP7_75t_L g1172 ( 
.A(n_1153),
.B(n_26),
.C(n_27),
.Y(n_1172)
);

OAI22x1_ASAP7_75t_L g1173 ( 
.A1(n_1150),
.A2(n_1152),
.B1(n_1151),
.B2(n_1170),
.Y(n_1173)
);

AOI221xp5_ASAP7_75t_L g1174 ( 
.A1(n_1162),
.A2(n_1020),
.B1(n_1024),
.B2(n_1040),
.C(n_932),
.Y(n_1174)
);

AND2x2_ASAP7_75t_L g1175 ( 
.A(n_1148),
.B(n_1155),
.Y(n_1175)
);

OAI22xp33_ASAP7_75t_SL g1176 ( 
.A1(n_1161),
.A2(n_996),
.B1(n_942),
.B2(n_935),
.Y(n_1176)
);

AOI222xp33_ASAP7_75t_L g1177 ( 
.A1(n_1163),
.A2(n_1024),
.B1(n_932),
.B2(n_1043),
.C1(n_31),
.C2(n_32),
.Y(n_1177)
);

NAND3xp33_ASAP7_75t_L g1178 ( 
.A(n_1171),
.B(n_28),
.C(n_29),
.Y(n_1178)
);

AOI21xp33_ASAP7_75t_L g1179 ( 
.A1(n_1157),
.A2(n_29),
.B(n_30),
.Y(n_1179)
);

INVx1_ASAP7_75t_L g1180 ( 
.A(n_1156),
.Y(n_1180)
);

INVx2_ASAP7_75t_SL g1181 ( 
.A(n_1149),
.Y(n_1181)
);

O2A1O1Ixp33_ASAP7_75t_L g1182 ( 
.A1(n_1164),
.A2(n_31),
.B(n_33),
.C(n_34),
.Y(n_1182)
);

AOI211xp5_ASAP7_75t_L g1183 ( 
.A1(n_1154),
.A2(n_1168),
.B(n_1169),
.C(n_1160),
.Y(n_1183)
);

OAI211xp5_ASAP7_75t_SL g1184 ( 
.A1(n_1158),
.A2(n_33),
.B(n_34),
.C(n_36),
.Y(n_1184)
);

OAI321xp33_ASAP7_75t_L g1185 ( 
.A1(n_1165),
.A2(n_996),
.A3(n_934),
.B1(n_1028),
.B2(n_1015),
.C(n_1012),
.Y(n_1185)
);

OAI211xp5_ASAP7_75t_SL g1186 ( 
.A1(n_1159),
.A2(n_36),
.B(n_38),
.C(n_40),
.Y(n_1186)
);

NOR3xp33_ASAP7_75t_L g1187 ( 
.A(n_1166),
.B(n_1167),
.C(n_42),
.Y(n_1187)
);

OAI221xp5_ASAP7_75t_L g1188 ( 
.A1(n_1148),
.A2(n_1023),
.B1(n_1006),
.B2(n_1010),
.C(n_1018),
.Y(n_1188)
);

OAI222xp33_ASAP7_75t_L g1189 ( 
.A1(n_1155),
.A2(n_1023),
.B1(n_1006),
.B2(n_1018),
.C1(n_978),
.C2(n_987),
.Y(n_1189)
);

OAI21xp33_ASAP7_75t_SL g1190 ( 
.A1(n_1155),
.A2(n_1023),
.B(n_1008),
.Y(n_1190)
);

INVx2_ASAP7_75t_SL g1191 ( 
.A(n_1151),
.Y(n_1191)
);

INVxp33_ASAP7_75t_SL g1192 ( 
.A(n_1150),
.Y(n_1192)
);

AOI22xp5_ASAP7_75t_L g1193 ( 
.A1(n_1148),
.A2(n_932),
.B1(n_1023),
.B2(n_1006),
.Y(n_1193)
);

OAI211xp5_ASAP7_75t_SL g1194 ( 
.A1(n_1150),
.A2(n_41),
.B(n_42),
.C(n_43),
.Y(n_1194)
);

A2O1A1Ixp33_ASAP7_75t_L g1195 ( 
.A1(n_1164),
.A2(n_965),
.B(n_1006),
.C(n_44),
.Y(n_1195)
);

OAI22xp5_ASAP7_75t_L g1196 ( 
.A1(n_1193),
.A2(n_932),
.B1(n_983),
.B2(n_975),
.Y(n_1196)
);

NOR2x1p5_ASAP7_75t_L g1197 ( 
.A(n_1178),
.B(n_41),
.Y(n_1197)
);

NAND4xp75_ASAP7_75t_L g1198 ( 
.A(n_1175),
.B(n_43),
.C(n_44),
.D(n_45),
.Y(n_1198)
);

XOR2xp5_ASAP7_75t_L g1199 ( 
.A(n_1192),
.B(n_46),
.Y(n_1199)
);

INVx1_ASAP7_75t_L g1200 ( 
.A(n_1173),
.Y(n_1200)
);

INVxp67_ASAP7_75t_L g1201 ( 
.A(n_1172),
.Y(n_1201)
);

NOR2x1_ASAP7_75t_L g1202 ( 
.A(n_1194),
.B(n_47),
.Y(n_1202)
);

NOR2x1p5_ASAP7_75t_L g1203 ( 
.A(n_1180),
.B(n_47),
.Y(n_1203)
);

NOR2x1_ASAP7_75t_L g1204 ( 
.A(n_1186),
.B(n_48),
.Y(n_1204)
);

OR2x2_ASAP7_75t_L g1205 ( 
.A(n_1181),
.B(n_1008),
.Y(n_1205)
);

AND2x2_ASAP7_75t_L g1206 ( 
.A(n_1191),
.B(n_978),
.Y(n_1206)
);

INVx2_ASAP7_75t_L g1207 ( 
.A(n_1188),
.Y(n_1207)
);

OAI22xp33_ASAP7_75t_L g1208 ( 
.A1(n_1179),
.A2(n_978),
.B1(n_1015),
.B2(n_987),
.Y(n_1208)
);

NAND4xp75_ASAP7_75t_L g1209 ( 
.A(n_1174),
.B(n_1008),
.C(n_1028),
.D(n_1012),
.Y(n_1209)
);

INVx2_ASAP7_75t_L g1210 ( 
.A(n_1190),
.Y(n_1210)
);

NOR2x1_ASAP7_75t_L g1211 ( 
.A(n_1184),
.B(n_411),
.Y(n_1211)
);

XOR2xp5_ASAP7_75t_L g1212 ( 
.A(n_1176),
.B(n_61),
.Y(n_1212)
);

INVx1_ASAP7_75t_L g1213 ( 
.A(n_1182),
.Y(n_1213)
);

NOR2x1_ASAP7_75t_L g1214 ( 
.A(n_1195),
.B(n_975),
.Y(n_1214)
);

NAND4xp75_ASAP7_75t_L g1215 ( 
.A(n_1177),
.B(n_1187),
.C(n_1183),
.D(n_1189),
.Y(n_1215)
);

AND2x4_ASAP7_75t_L g1216 ( 
.A(n_1185),
.B(n_1011),
.Y(n_1216)
);

AND2x4_ASAP7_75t_L g1217 ( 
.A(n_1191),
.B(n_983),
.Y(n_1217)
);

NOR2xp33_ASAP7_75t_L g1218 ( 
.A(n_1198),
.B(n_64),
.Y(n_1218)
);

NOR3xp33_ASAP7_75t_L g1219 ( 
.A(n_1200),
.B(n_949),
.C(n_943),
.Y(n_1219)
);

NAND2x1p5_ASAP7_75t_L g1220 ( 
.A(n_1203),
.B(n_983),
.Y(n_1220)
);

AND3x1_ASAP7_75t_L g1221 ( 
.A(n_1202),
.B(n_1028),
.C(n_1012),
.Y(n_1221)
);

NAND3xp33_ASAP7_75t_L g1222 ( 
.A(n_1213),
.B(n_1201),
.C(n_1211),
.Y(n_1222)
);

INVx1_ASAP7_75t_L g1223 ( 
.A(n_1199),
.Y(n_1223)
);

AND2x4_ASAP7_75t_L g1224 ( 
.A(n_1217),
.B(n_1011),
.Y(n_1224)
);

NOR3xp33_ASAP7_75t_L g1225 ( 
.A(n_1215),
.B(n_949),
.C(n_943),
.Y(n_1225)
);

NOR2xp33_ASAP7_75t_L g1226 ( 
.A(n_1210),
.B(n_65),
.Y(n_1226)
);

OR3x1_ASAP7_75t_L g1227 ( 
.A(n_1212),
.B(n_1197),
.C(n_1204),
.Y(n_1227)
);

AND2x4_ASAP7_75t_L g1228 ( 
.A(n_1217),
.B(n_1011),
.Y(n_1228)
);

NOR2x1p5_ASAP7_75t_L g1229 ( 
.A(n_1207),
.B(n_943),
.Y(n_1229)
);

AOI211xp5_ASAP7_75t_L g1230 ( 
.A1(n_1205),
.A2(n_1016),
.B(n_1011),
.C(n_1015),
.Y(n_1230)
);

NOR3xp33_ASAP7_75t_L g1231 ( 
.A(n_1196),
.B(n_949),
.C(n_919),
.Y(n_1231)
);

NAND4xp75_ASAP7_75t_L g1232 ( 
.A(n_1214),
.B(n_1206),
.C(n_1209),
.D(n_1208),
.Y(n_1232)
);

XNOR2xp5_ASAP7_75t_L g1233 ( 
.A(n_1227),
.B(n_1232),
.Y(n_1233)
);

XNOR2x1_ASAP7_75t_L g1234 ( 
.A(n_1223),
.B(n_1216),
.Y(n_1234)
);

INVx1_ASAP7_75t_L g1235 ( 
.A(n_1222),
.Y(n_1235)
);

INVx2_ASAP7_75t_L g1236 ( 
.A(n_1220),
.Y(n_1236)
);

XNOR2x1_ASAP7_75t_L g1237 ( 
.A(n_1229),
.B(n_66),
.Y(n_1237)
);

BUFx2_ASAP7_75t_L g1238 ( 
.A(n_1221),
.Y(n_1238)
);

NAND2xp5_ASAP7_75t_L g1239 ( 
.A(n_1218),
.B(n_962),
.Y(n_1239)
);

OAI21xp5_ASAP7_75t_L g1240 ( 
.A1(n_1226),
.A2(n_1016),
.B(n_1011),
.Y(n_1240)
);

NOR4xp25_ASAP7_75t_L g1241 ( 
.A(n_1219),
.B(n_69),
.C(n_71),
.D(n_72),
.Y(n_1241)
);

AND2x2_ASAP7_75t_L g1242 ( 
.A(n_1224),
.B(n_1016),
.Y(n_1242)
);

NAND2xp5_ASAP7_75t_L g1243 ( 
.A(n_1228),
.B(n_962),
.Y(n_1243)
);

INVx2_ASAP7_75t_L g1244 ( 
.A(n_1225),
.Y(n_1244)
);

NAND2xp5_ASAP7_75t_L g1245 ( 
.A(n_1231),
.B(n_1016),
.Y(n_1245)
);

AOI22xp5_ASAP7_75t_L g1246 ( 
.A1(n_1230),
.A2(n_1016),
.B1(n_1011),
.B2(n_938),
.Y(n_1246)
);

AOI221xp5_ASAP7_75t_L g1247 ( 
.A1(n_1226),
.A2(n_1016),
.B1(n_919),
.B2(n_938),
.C(n_916),
.Y(n_1247)
);

AOI22xp5_ASAP7_75t_L g1248 ( 
.A1(n_1233),
.A2(n_938),
.B1(n_939),
.B2(n_952),
.Y(n_1248)
);

AO22x2_ASAP7_75t_L g1249 ( 
.A1(n_1234),
.A2(n_987),
.B1(n_939),
.B2(n_950),
.Y(n_1249)
);

AOI22xp5_ASAP7_75t_L g1250 ( 
.A1(n_1238),
.A2(n_938),
.B1(n_939),
.B2(n_952),
.Y(n_1250)
);

INVx1_ASAP7_75t_L g1251 ( 
.A(n_1236),
.Y(n_1251)
);

AOI22xp5_ASAP7_75t_L g1252 ( 
.A1(n_1235),
.A2(n_938),
.B1(n_950),
.B2(n_921),
.Y(n_1252)
);

AOI22xp5_ASAP7_75t_L g1253 ( 
.A1(n_1235),
.A2(n_938),
.B1(n_921),
.B2(n_916),
.Y(n_1253)
);

AOI22xp33_ASAP7_75t_SL g1254 ( 
.A1(n_1244),
.A2(n_1239),
.B1(n_1237),
.B2(n_1242),
.Y(n_1254)
);

AOI22xp5_ASAP7_75t_L g1255 ( 
.A1(n_1243),
.A2(n_938),
.B1(n_915),
.B2(n_925),
.Y(n_1255)
);

AOI22xp5_ASAP7_75t_L g1256 ( 
.A1(n_1246),
.A2(n_915),
.B1(n_925),
.B2(n_987),
.Y(n_1256)
);

AOI22xp5_ASAP7_75t_L g1257 ( 
.A1(n_1245),
.A2(n_915),
.B1(n_925),
.B2(n_957),
.Y(n_1257)
);

INVx3_ASAP7_75t_L g1258 ( 
.A(n_1251),
.Y(n_1258)
);

INVx2_ASAP7_75t_L g1259 ( 
.A(n_1249),
.Y(n_1259)
);

AOI22xp5_ASAP7_75t_L g1260 ( 
.A1(n_1254),
.A2(n_1241),
.B1(n_1247),
.B2(n_1240),
.Y(n_1260)
);

OAI22xp5_ASAP7_75t_L g1261 ( 
.A1(n_1248),
.A2(n_925),
.B1(n_77),
.B2(n_78),
.Y(n_1261)
);

OR2x2_ASAP7_75t_L g1262 ( 
.A(n_1250),
.B(n_74),
.Y(n_1262)
);

OAI22xp33_ASAP7_75t_L g1263 ( 
.A1(n_1252),
.A2(n_925),
.B1(n_80),
.B2(n_83),
.Y(n_1263)
);

OAI22xp5_ASAP7_75t_SL g1264 ( 
.A1(n_1258),
.A2(n_1253),
.B1(n_1256),
.B2(n_1255),
.Y(n_1264)
);

BUFx2_ASAP7_75t_L g1265 ( 
.A(n_1259),
.Y(n_1265)
);

AOI31xp33_ASAP7_75t_L g1266 ( 
.A1(n_1260),
.A2(n_1257),
.A3(n_85),
.B(n_87),
.Y(n_1266)
);

OAI22x1_ASAP7_75t_L g1267 ( 
.A1(n_1262),
.A2(n_79),
.B1(n_88),
.B2(n_91),
.Y(n_1267)
);

NAND2xp5_ASAP7_75t_SL g1268 ( 
.A(n_1265),
.B(n_1263),
.Y(n_1268)
);

NAND2xp33_ASAP7_75t_SL g1269 ( 
.A(n_1268),
.B(n_1267),
.Y(n_1269)
);

NAND3xp33_ASAP7_75t_L g1270 ( 
.A(n_1269),
.B(n_1266),
.C(n_1261),
.Y(n_1270)
);

AO21x2_ASAP7_75t_L g1271 ( 
.A1(n_1270),
.A2(n_1264),
.B(n_98),
.Y(n_1271)
);

OAI221xp5_ASAP7_75t_R g1272 ( 
.A1(n_1271),
.A2(n_96),
.B1(n_101),
.B2(n_102),
.C(n_103),
.Y(n_1272)
);

AOI211xp5_ASAP7_75t_L g1273 ( 
.A1(n_1272),
.A2(n_104),
.B(n_105),
.C(n_109),
.Y(n_1273)
);


endmodule