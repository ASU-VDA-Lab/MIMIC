module fake_jpeg_12791_n_344 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_344);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_344;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx11_ASAP7_75t_SL g17 ( 
.A(n_4),
.Y(n_17)
);

INVx6_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_11),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_16),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

INVx5_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

BUFx16f_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_0),
.B(n_16),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_11),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_16),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_8),
.B(n_0),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_5),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_6),
.B(n_15),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_13),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_2),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_12),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_3),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_SL g40 ( 
.A(n_8),
.B(n_14),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_10),
.Y(n_41)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_2),
.Y(n_42)
);

INVx11_ASAP7_75t_L g43 ( 
.A(n_17),
.Y(n_43)
);

INVx11_ASAP7_75t_L g112 ( 
.A(n_43),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_28),
.B(n_1),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_44),
.B(n_1),
.Y(n_70)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_42),
.Y(n_45)
);

INVx5_ASAP7_75t_L g79 ( 
.A(n_45),
.Y(n_79)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_25),
.Y(n_46)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_46),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_32),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_47),
.Y(n_93)
);

INVx11_ASAP7_75t_L g48 ( 
.A(n_17),
.Y(n_48)
);

BUFx5_ASAP7_75t_L g104 ( 
.A(n_48),
.Y(n_104)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_42),
.Y(n_49)
);

INVx5_ASAP7_75t_L g83 ( 
.A(n_49),
.Y(n_83)
);

BUFx5_ASAP7_75t_L g50 ( 
.A(n_42),
.Y(n_50)
);

BUFx2_ASAP7_75t_L g96 ( 
.A(n_50),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_40),
.B(n_9),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_51),
.B(n_65),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_32),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_52),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_32),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_53),
.Y(n_113)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_27),
.Y(n_54)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_54),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_28),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_55),
.B(n_33),
.Y(n_69)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_19),
.Y(n_56)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_56),
.Y(n_84)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_25),
.Y(n_57)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_57),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_40),
.B(n_9),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_58),
.B(n_62),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_22),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_59),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_22),
.Y(n_60)
);

INVx6_ASAP7_75t_L g90 ( 
.A(n_60),
.Y(n_90)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_22),
.Y(n_61)
);

INVx5_ASAP7_75t_L g87 ( 
.A(n_61),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_35),
.B(n_7),
.Y(n_62)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_18),
.Y(n_63)
);

INVx5_ASAP7_75t_L g98 ( 
.A(n_63),
.Y(n_98)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_27),
.Y(n_64)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_64),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g65 ( 
.A(n_35),
.B(n_7),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_22),
.Y(n_66)
);

INVx5_ASAP7_75t_L g103 ( 
.A(n_66),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_18),
.Y(n_67)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_67),
.Y(n_109)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_37),
.Y(n_68)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_68),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_69),
.B(n_73),
.Y(n_136)
);

NAND3xp33_ASAP7_75t_L g139 ( 
.A(n_70),
.B(n_10),
.C(n_15),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_55),
.B(n_33),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_44),
.B(n_39),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_74),
.B(n_75),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_56),
.B(n_39),
.Y(n_75)
);

CKINVDCx12_ASAP7_75t_R g76 ( 
.A(n_43),
.Y(n_76)
);

CKINVDCx16_ASAP7_75t_R g140 ( 
.A(n_76),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_65),
.A2(n_21),
.B1(n_20),
.B2(n_36),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_77),
.A2(n_10),
.B1(n_14),
.B2(n_3),
.Y(n_150)
);

CKINVDCx9p33_ASAP7_75t_R g78 ( 
.A(n_48),
.Y(n_78)
);

OR2x2_ASAP7_75t_L g130 ( 
.A(n_78),
.B(n_26),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_47),
.A2(n_52),
.B1(n_53),
.B2(n_68),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_80),
.A2(n_66),
.B1(n_60),
.B2(n_67),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_46),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_81),
.B(n_86),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_54),
.B(n_37),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_85),
.B(n_70),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_51),
.B(n_20),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_L g88 ( 
.A1(n_47),
.A2(n_18),
.B1(n_36),
.B2(n_34),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_88),
.A2(n_91),
.B1(n_52),
.B2(n_53),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_45),
.A2(n_24),
.B1(n_38),
.B2(n_30),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_89),
.A2(n_26),
.B1(n_23),
.B2(n_19),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_64),
.A2(n_24),
.B1(n_38),
.B2(n_30),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_57),
.B(n_34),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_95),
.B(n_101),
.Y(n_138)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_63),
.Y(n_99)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_99),
.Y(n_117)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_49),
.Y(n_100)
);

INVx4_ASAP7_75t_L g141 ( 
.A(n_100),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_49),
.B(n_31),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_49),
.B(n_21),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_102),
.B(n_105),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_50),
.B(n_29),
.Y(n_105)
);

INVx4_ASAP7_75t_SL g106 ( 
.A(n_59),
.Y(n_106)
);

INVx4_ASAP7_75t_L g155 ( 
.A(n_106),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_45),
.B(n_29),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_107),
.B(n_115),
.Y(n_152)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_61),
.Y(n_111)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_111),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g115 ( 
.A(n_59),
.B(n_31),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_63),
.B(n_41),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_116),
.Y(n_127)
);

AND2x2_ASAP7_75t_SL g118 ( 
.A(n_75),
.B(n_85),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_118),
.B(n_82),
.C(n_112),
.Y(n_178)
);

AND2x4_ASAP7_75t_L g119 ( 
.A(n_72),
.B(n_24),
.Y(n_119)
);

INVx1_ASAP7_75t_SL g180 ( 
.A(n_119),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_121),
.A2(n_126),
.B1(n_129),
.B2(n_132),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_123),
.B(n_150),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_74),
.B(n_41),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_125),
.B(n_108),
.Y(n_164)
);

INVxp67_ASAP7_75t_L g160 ( 
.A(n_128),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_80),
.A2(n_67),
.B1(n_66),
.B2(n_60),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g176 ( 
.A(n_130),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_93),
.Y(n_131)
);

INVx3_ASAP7_75t_L g161 ( 
.A(n_131),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_91),
.A2(n_23),
.B1(n_25),
.B2(n_3),
.Y(n_132)
);

HB1xp67_ASAP7_75t_L g133 ( 
.A(n_84),
.Y(n_133)
);

HB1xp67_ASAP7_75t_L g185 ( 
.A(n_133),
.Y(n_185)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_87),
.Y(n_134)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_134),
.Y(n_192)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_93),
.Y(n_135)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_135),
.Y(n_165)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_84),
.Y(n_137)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_137),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_139),
.B(n_142),
.Y(n_163)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_96),
.Y(n_142)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_87),
.Y(n_143)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_143),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_78),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_144),
.B(n_145),
.Y(n_186)
);

NAND2xp33_ASAP7_75t_SL g145 ( 
.A(n_92),
.B(n_25),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_112),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_146),
.B(n_104),
.Y(n_189)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_97),
.Y(n_147)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_147),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_L g148 ( 
.A1(n_109),
.A2(n_113),
.B1(n_110),
.B2(n_99),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_148),
.A2(n_153),
.B1(n_113),
.B2(n_110),
.Y(n_162)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_109),
.Y(n_149)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_149),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_90),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_71),
.Y(n_154)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_154),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_SL g156 ( 
.A(n_136),
.B(n_94),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_SL g207 ( 
.A(n_156),
.B(n_140),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_162),
.A2(n_172),
.B1(n_177),
.B2(n_188),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_164),
.B(n_138),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_122),
.B(n_90),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_167),
.B(n_169),
.Y(n_204)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_117),
.Y(n_168)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_168),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_122),
.B(n_71),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_SL g170 ( 
.A1(n_132),
.A2(n_96),
.B1(n_100),
.B2(n_83),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_SL g205 ( 
.A1(n_170),
.A2(n_174),
.B1(n_175),
.B2(n_155),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_123),
.A2(n_114),
.B1(n_111),
.B2(n_98),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_SL g174 ( 
.A1(n_127),
.A2(n_83),
.B1(n_79),
.B2(n_82),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_SL g175 ( 
.A1(n_127),
.A2(n_144),
.B1(n_137),
.B2(n_129),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_125),
.A2(n_114),
.B1(n_98),
.B2(n_103),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_178),
.B(n_182),
.Y(n_202)
);

AOI21xp5_ASAP7_75t_L g179 ( 
.A1(n_130),
.A2(n_79),
.B(n_103),
.Y(n_179)
);

AOI21xp5_ASAP7_75t_L g223 ( 
.A1(n_179),
.A2(n_182),
.B(n_178),
.Y(n_223)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_117),
.Y(n_181)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_181),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_118),
.B(n_106),
.C(n_104),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_118),
.B(n_4),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_184),
.B(n_191),
.Y(n_208)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_147),
.Y(n_187)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_187),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_150),
.A2(n_6),
.B1(n_12),
.B2(n_13),
.Y(n_188)
);

CKINVDCx14_ASAP7_75t_R g215 ( 
.A(n_189),
.Y(n_215)
);

AO22x2_ASAP7_75t_SL g190 ( 
.A1(n_126),
.A2(n_15),
.B1(n_12),
.B2(n_13),
.Y(n_190)
);

OA22x2_ASAP7_75t_L g203 ( 
.A1(n_190),
.A2(n_153),
.B1(n_155),
.B2(n_131),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_152),
.B(n_6),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_191),
.B(n_120),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_193),
.B(n_194),
.Y(n_243)
);

INVx8_ASAP7_75t_L g195 ( 
.A(n_161),
.Y(n_195)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_195),
.Y(n_235)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_157),
.Y(n_196)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_196),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_164),
.B(n_151),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_198),
.B(n_207),
.Y(n_248)
);

OR2x6_ASAP7_75t_L g199 ( 
.A(n_180),
.B(n_119),
.Y(n_199)
);

BUFx24_ASAP7_75t_L g233 ( 
.A(n_199),
.Y(n_233)
);

OAI21xp33_ASAP7_75t_SL g200 ( 
.A1(n_176),
.A2(n_119),
.B(n_146),
.Y(n_200)
);

OAI21xp33_ASAP7_75t_L g241 ( 
.A1(n_200),
.A2(n_173),
.B(n_171),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_SL g201 ( 
.A1(n_180),
.A2(n_119),
.B(n_154),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_201),
.B(n_206),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_203),
.B(n_210),
.Y(n_234)
);

CKINVDCx16_ASAP7_75t_R g231 ( 
.A(n_205),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_SL g206 ( 
.A1(n_186),
.A2(n_176),
.B(n_160),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_183),
.A2(n_124),
.B1(n_149),
.B2(n_135),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_209),
.A2(n_214),
.B1(n_218),
.B2(n_162),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_167),
.B(n_124),
.Y(n_210)
);

CKINVDCx16_ASAP7_75t_R g211 ( 
.A(n_185),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_211),
.B(n_219),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_183),
.A2(n_134),
.B1(n_143),
.B2(n_142),
.Y(n_214)
);

INVx1_ASAP7_75t_SL g216 ( 
.A(n_166),
.Y(n_216)
);

INVx13_ASAP7_75t_L g242 ( 
.A(n_216),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_169),
.B(n_141),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_217),
.B(n_226),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_158),
.A2(n_14),
.B1(n_141),
.B2(n_160),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_159),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_166),
.Y(n_220)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_220),
.Y(n_229)
);

CKINVDCx16_ASAP7_75t_R g221 ( 
.A(n_179),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_221),
.B(n_222),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_SL g222 ( 
.A(n_163),
.B(n_184),
.Y(n_222)
);

CKINVDCx16_ASAP7_75t_R g238 ( 
.A(n_223),
.Y(n_238)
);

BUFx12f_ASAP7_75t_L g225 ( 
.A(n_192),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_225),
.B(n_171),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_173),
.B(n_172),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_217),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_236),
.B(n_247),
.Y(n_257)
);

BUFx2_ASAP7_75t_L g260 ( 
.A(n_239),
.Y(n_260)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_220),
.Y(n_240)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_240),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_241),
.B(n_201),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_213),
.A2(n_190),
.B1(n_177),
.B2(n_165),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_244),
.B(n_249),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_245),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_215),
.B(n_192),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_246),
.B(n_253),
.Y(n_273)
);

AND2x6_ASAP7_75t_L g247 ( 
.A(n_202),
.B(n_190),
.Y(n_247)
);

CKINVDCx14_ASAP7_75t_R g249 ( 
.A(n_199),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_197),
.Y(n_250)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_250),
.Y(n_268)
);

AND2x6_ASAP7_75t_L g251 ( 
.A(n_202),
.B(n_223),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_251),
.B(n_199),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_204),
.B(n_210),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_252),
.B(n_208),
.C(n_224),
.Y(n_265)
);

NOR2xp67_ASAP7_75t_L g253 ( 
.A(n_218),
.B(n_188),
.Y(n_253)
);

OAI21xp5_ASAP7_75t_SL g279 ( 
.A1(n_254),
.A2(n_259),
.B(n_263),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_234),
.A2(n_213),
.B1(n_204),
.B2(n_226),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_255),
.A2(n_261),
.B1(n_250),
.B2(n_203),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_227),
.B(n_206),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_258),
.B(n_262),
.C(n_265),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_234),
.A2(n_199),
.B1(n_203),
.B2(n_190),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_227),
.B(n_208),
.Y(n_262)
);

AOI21xp5_ASAP7_75t_L g263 ( 
.A1(n_233),
.A2(n_199),
.B(n_197),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_236),
.B(n_216),
.Y(n_264)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_264),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_237),
.B(n_212),
.Y(n_269)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_269),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_L g270 ( 
.A1(n_233),
.A2(n_209),
.B(n_212),
.Y(n_270)
);

OAI21xp5_ASAP7_75t_L g290 ( 
.A1(n_270),
.A2(n_228),
.B(n_242),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_237),
.B(n_196),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_271),
.B(n_272),
.Y(n_285)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_229),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_230),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_274),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_233),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_275),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_260),
.A2(n_239),
.B1(n_231),
.B2(n_247),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_277),
.A2(n_284),
.B1(n_286),
.B2(n_261),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_274),
.B(n_248),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_SL g293 ( 
.A(n_281),
.B(n_292),
.Y(n_293)
);

OAI21xp5_ASAP7_75t_SL g283 ( 
.A1(n_263),
.A2(n_233),
.B(n_231),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_SL g299 ( 
.A(n_283),
.B(n_289),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_L g284 ( 
.A1(n_260),
.A2(n_238),
.B1(n_252),
.B2(n_244),
.Y(n_284)
);

OAI22xp33_ASAP7_75t_SL g286 ( 
.A1(n_273),
.A2(n_203),
.B1(n_240),
.B2(n_229),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_258),
.B(n_251),
.C(n_232),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_287),
.B(n_276),
.C(n_259),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_288),
.A2(n_256),
.B1(n_264),
.B2(n_270),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_290),
.B(n_289),
.Y(n_298)
);

XOR2xp5_ASAP7_75t_L g291 ( 
.A(n_262),
.B(n_243),
.Y(n_291)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_291),
.B(n_254),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_267),
.B(n_225),
.Y(n_292)
);

XOR2xp5_ASAP7_75t_L g308 ( 
.A(n_294),
.B(n_295),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_276),
.B(n_265),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_285),
.Y(n_296)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_296),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_SL g315 ( 
.A(n_297),
.B(n_303),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_298),
.B(n_299),
.Y(n_311)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_285),
.Y(n_300)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_300),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_301),
.A2(n_278),
.B1(n_280),
.B2(n_277),
.Y(n_307)
);

HB1xp67_ASAP7_75t_L g314 ( 
.A(n_302),
.Y(n_314)
);

XOR2xp5_ASAP7_75t_L g303 ( 
.A(n_287),
.B(n_257),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_291),
.B(n_256),
.C(n_275),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_304),
.B(n_305),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_279),
.B(n_269),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g306 ( 
.A(n_284),
.B(n_255),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_306),
.B(n_288),
.Y(n_312)
);

INVxp67_ASAP7_75t_L g321 ( 
.A(n_307),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_SL g319 ( 
.A(n_312),
.B(n_282),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_293),
.B(n_282),
.Y(n_313)
);

NAND3xp33_ASAP7_75t_L g320 ( 
.A(n_313),
.B(n_280),
.C(n_278),
.Y(n_320)
);

BUFx6f_ASAP7_75t_L g317 ( 
.A(n_303),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_SL g325 ( 
.A(n_317),
.B(n_306),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_308),
.B(n_295),
.C(n_294),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_318),
.B(n_319),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_320),
.B(n_322),
.Y(n_331)
);

OAI21xp5_ASAP7_75t_SL g322 ( 
.A1(n_311),
.A2(n_304),
.B(n_267),
.Y(n_322)
);

CKINVDCx14_ASAP7_75t_R g323 ( 
.A(n_311),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_323),
.B(n_325),
.Y(n_329)
);

OAI21xp5_ASAP7_75t_L g324 ( 
.A1(n_310),
.A2(n_279),
.B(n_290),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_L g328 ( 
.A1(n_324),
.A2(n_309),
.B1(n_316),
.B2(n_297),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_308),
.B(n_315),
.C(n_317),
.Y(n_326)
);

OAI21xp5_ASAP7_75t_SL g332 ( 
.A1(n_326),
.A2(n_271),
.B(n_235),
.Y(n_332)
);

AOI21xp5_ASAP7_75t_L g327 ( 
.A1(n_321),
.A2(n_307),
.B(n_314),
.Y(n_327)
);

XNOR2xp5_ASAP7_75t_L g334 ( 
.A(n_327),
.B(n_272),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_SL g336 ( 
.A(n_328),
.B(n_332),
.Y(n_336)
);

XNOR2xp5_ASAP7_75t_L g333 ( 
.A(n_323),
.B(n_283),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_SL g337 ( 
.A(n_333),
.B(n_329),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_334),
.B(n_335),
.C(n_337),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_327),
.B(n_330),
.C(n_331),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_335),
.B(n_333),
.C(n_266),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_SL g340 ( 
.A(n_339),
.B(n_336),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_340),
.B(n_338),
.C(n_266),
.Y(n_341)
);

OAI331xp33_ASAP7_75t_L g342 ( 
.A1(n_341),
.A2(n_268),
.A3(n_228),
.B1(n_242),
.B2(n_235),
.B3(n_165),
.C1(n_195),
.Y(n_342)
);

OAI21xp5_ASAP7_75t_SL g343 ( 
.A1(n_342),
.A2(n_268),
.B(n_225),
.Y(n_343)
);

XOR2xp5_ASAP7_75t_L g344 ( 
.A(n_343),
.B(n_161),
.Y(n_344)
);


endmodule