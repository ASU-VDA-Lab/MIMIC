module fake_jpeg_17415_n_150 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_150);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_150;

wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g40 ( 
.A(n_27),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_11),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_38),
.Y(n_42)
);

BUFx12_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_10),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_2),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_39),
.Y(n_47)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_29),
.Y(n_48)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_13),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_18),
.Y(n_50)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_24),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_3),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_28),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_19),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_5),
.Y(n_55)
);

INVxp67_ASAP7_75t_L g56 ( 
.A(n_23),
.Y(n_56)
);

BUFx5_ASAP7_75t_L g57 ( 
.A(n_21),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_16),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_59),
.Y(n_72)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_50),
.Y(n_60)
);

INVx8_ASAP7_75t_L g73 ( 
.A(n_60),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_61),
.Y(n_70)
);

INVx3_ASAP7_75t_SL g62 ( 
.A(n_44),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_62),
.B(n_64),
.Y(n_67)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_50),
.Y(n_63)
);

INVx5_ASAP7_75t_L g68 ( 
.A(n_63),
.Y(n_68)
);

CKINVDCx16_ASAP7_75t_R g64 ( 
.A(n_40),
.Y(n_64)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_46),
.Y(n_65)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_65),
.Y(n_69)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_46),
.Y(n_66)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_66),
.Y(n_74)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_59),
.Y(n_71)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_71),
.Y(n_84)
);

INVx2_ASAP7_75t_SL g75 ( 
.A(n_62),
.Y(n_75)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_75),
.Y(n_87)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_61),
.Y(n_76)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_76),
.Y(n_86)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_60),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_77),
.B(n_78),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_59),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_62),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_79),
.B(n_81),
.Y(n_85)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_59),
.Y(n_80)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_80),
.Y(n_95)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_65),
.Y(n_81)
);

INVx6_ASAP7_75t_L g82 ( 
.A(n_59),
.Y(n_82)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_82),
.Y(n_99)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_65),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_83),
.B(n_52),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_72),
.Y(n_88)
);

INVx1_ASAP7_75t_SL g114 ( 
.A(n_88),
.Y(n_114)
);

BUFx2_ASAP7_75t_L g90 ( 
.A(n_68),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_90),
.B(n_100),
.Y(n_104)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_91),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_L g92 ( 
.A1(n_70),
.A2(n_69),
.B1(n_74),
.B2(n_51),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_L g106 ( 
.A1(n_92),
.A2(n_102),
.B1(n_54),
.B2(n_43),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_73),
.A2(n_55),
.B1(n_49),
.B2(n_56),
.Y(n_93)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_93),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_67),
.B(n_0),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_94),
.B(n_103),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_78),
.Y(n_96)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_96),
.Y(n_113)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_67),
.B(n_0),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_97),
.B(n_1),
.Y(n_111)
);

AND2x2_ASAP7_75t_SL g98 ( 
.A(n_75),
.B(n_42),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_98),
.B(n_45),
.C(n_57),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_72),
.Y(n_100)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_71),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_101),
.B(n_43),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_L g102 ( 
.A1(n_82),
.A2(n_48),
.B1(n_58),
.B2(n_54),
.Y(n_102)
);

OR2x2_ASAP7_75t_L g103 ( 
.A(n_67),
.B(n_53),
.Y(n_103)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_105),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_106),
.A2(n_110),
.B1(n_87),
.B2(n_85),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_107),
.B(n_111),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_99),
.A2(n_47),
.B1(n_56),
.B2(n_3),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_94),
.B(n_97),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_115),
.B(n_98),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_109),
.A2(n_89),
.B1(n_106),
.B2(n_84),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_118),
.A2(n_110),
.B1(n_89),
.B2(n_104),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_119),
.B(n_120),
.Y(n_126)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_113),
.Y(n_121)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_121),
.Y(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_117),
.Y(n_123)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_123),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_118),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_SL g130 ( 
.A1(n_124),
.A2(n_122),
.B(n_112),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_125),
.A2(n_114),
.B1(n_2),
.B2(n_4),
.Y(n_132)
);

AOI21xp5_ASAP7_75t_L g127 ( 
.A1(n_126),
.A2(n_119),
.B(n_116),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_127),
.A2(n_128),
.B1(n_130),
.B2(n_132),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_L g128 ( 
.A1(n_125),
.A2(n_114),
.B1(n_95),
.B2(n_86),
.Y(n_128)
);

XOR2xp5_ASAP7_75t_L g131 ( 
.A(n_126),
.B(n_108),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_131),
.B(n_1),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_129),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_SL g137 ( 
.A1(n_134),
.A2(n_136),
.B(n_4),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_135),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_128),
.A2(n_17),
.B1(n_37),
.B2(n_36),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_137),
.A2(n_133),
.B1(n_5),
.B2(n_6),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_139),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g141 ( 
.A(n_140),
.B(n_138),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_141),
.A2(n_20),
.B1(n_34),
.B2(n_32),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_142),
.B(n_14),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_143),
.B(n_15),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_144),
.B(n_12),
.C(n_31),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_145),
.B(n_9),
.Y(n_146)
);

CKINVDCx16_ASAP7_75t_R g147 ( 
.A(n_146),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_L g148 ( 
.A1(n_147),
.A2(n_22),
.B(n_30),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_L g149 ( 
.A1(n_148),
.A2(n_8),
.B(n_26),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_L g150 ( 
.A1(n_149),
.A2(n_7),
.B(n_25),
.Y(n_150)
);


endmodule