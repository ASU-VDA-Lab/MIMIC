module fake_jpeg_16889_n_293 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_293);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_293;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_223;
wire n_187;
wire n_57;
wire n_21;
wire n_175;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_125;
wire n_80;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_212;
wire n_131;
wire n_56;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_270;
wire n_260;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

BUFx12f_ASAP7_75t_L g14 ( 
.A(n_9),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_8),
.Y(n_15)
);

INVx4_ASAP7_75t_L g16 ( 
.A(n_12),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_6),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_5),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_8),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

INVx6_ASAP7_75t_SL g26 ( 
.A(n_1),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_4),
.Y(n_27)
);

INVx11_ASAP7_75t_SL g28 ( 
.A(n_0),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_18),
.Y(n_30)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_30),
.Y(n_42)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_18),
.Y(n_31)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_31),
.Y(n_52)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_32),
.Y(n_47)
);

CKINVDCx16_ASAP7_75t_R g33 ( 
.A(n_28),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_33),
.B(n_35),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_18),
.Y(n_34)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_34),
.Y(n_48)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_14),
.Y(n_36)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_36),
.Y(n_40)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_18),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_37),
.B(n_19),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_14),
.Y(n_38)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_38),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_30),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_43),
.B(n_44),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_30),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_SL g45 ( 
.A(n_33),
.B(n_15),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_45),
.B(n_53),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_30),
.B(n_14),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_46),
.B(n_49),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_34),
.B(n_14),
.Y(n_49)
);

MAJIxp5_ASAP7_75t_L g50 ( 
.A(n_36),
.B(n_29),
.C(n_25),
.Y(n_50)
);

OAI21xp5_ASAP7_75t_L g59 ( 
.A1(n_50),
.A2(n_51),
.B(n_54),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_31),
.A2(n_16),
.B1(n_26),
.B2(n_20),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_31),
.A2(n_16),
.B1(n_26),
.B2(n_20),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_55),
.Y(n_79)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_42),
.Y(n_56)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_56),
.Y(n_81)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_52),
.Y(n_57)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_57),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_46),
.B(n_35),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_60),
.B(n_61),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_46),
.B(n_38),
.Y(n_61)
);

OR2x2_ASAP7_75t_L g62 ( 
.A(n_51),
.B(n_22),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_62),
.B(n_75),
.Y(n_84)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

INVx5_ASAP7_75t_L g80 ( 
.A(n_63),
.Y(n_80)
);

INVxp67_ASAP7_75t_L g66 ( 
.A(n_39),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_66),
.B(n_71),
.Y(n_91)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_52),
.Y(n_67)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_67),
.Y(n_86)
);

INVx4_ASAP7_75t_SL g68 ( 
.A(n_52),
.Y(n_68)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_68),
.Y(n_90)
);

INVx2_ASAP7_75t_SL g69 ( 
.A(n_42),
.Y(n_69)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_69),
.Y(n_93)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_48),
.Y(n_70)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_70),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_45),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_51),
.A2(n_16),
.B1(n_26),
.B2(n_20),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_72),
.A2(n_54),
.B1(n_23),
.B2(n_37),
.Y(n_88)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_48),
.Y(n_73)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_73),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_39),
.Y(n_74)
);

OR2x2_ASAP7_75t_L g82 ( 
.A(n_74),
.B(n_54),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_49),
.B(n_24),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_49),
.B(n_35),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_76),
.B(n_38),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_41),
.A2(n_21),
.B1(n_24),
.B2(n_23),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_77),
.A2(n_78),
.B1(n_21),
.B2(n_22),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_41),
.A2(n_24),
.B1(n_21),
.B2(n_23),
.Y(n_78)
);

OAI21xp5_ASAP7_75t_L g114 ( 
.A1(n_82),
.A2(n_65),
.B(n_28),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_87),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_88),
.B(n_62),
.Y(n_111)
);

XNOR2xp5_ASAP7_75t_SL g89 ( 
.A(n_58),
.B(n_50),
.Y(n_89)
);

XNOR2xp5_ASAP7_75t_SL g128 ( 
.A(n_89),
.B(n_29),
.Y(n_128)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_56),
.Y(n_92)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_92),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_SL g94 ( 
.A1(n_60),
.A2(n_53),
.B(n_50),
.Y(n_94)
);

AOI21xp5_ASAP7_75t_L g116 ( 
.A1(n_94),
.A2(n_57),
.B(n_67),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_58),
.A2(n_37),
.B1(n_43),
.B2(n_44),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_96),
.A2(n_101),
.B1(n_63),
.B2(n_69),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_97),
.B(n_100),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_59),
.A2(n_48),
.B1(n_32),
.B2(n_47),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_98),
.A2(n_72),
.B1(n_74),
.B2(n_68),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_76),
.B(n_36),
.C(n_38),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_99),
.B(n_36),
.C(n_38),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_75),
.B(n_47),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_59),
.A2(n_32),
.B1(n_47),
.B2(n_34),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_61),
.B(n_40),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_102),
.B(n_62),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_64),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_104),
.B(n_105),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_64),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_107),
.A2(n_122),
.B1(n_124),
.B2(n_126),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_108),
.B(n_109),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_83),
.B(n_65),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_111),
.A2(n_84),
.B1(n_82),
.B2(n_88),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_112),
.B(n_128),
.C(n_99),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_SL g132 ( 
.A1(n_114),
.A2(n_116),
.B(n_117),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_83),
.B(n_71),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_115),
.B(n_119),
.Y(n_153)
);

A2O1A1O1Ixp25_ASAP7_75t_L g117 ( 
.A1(n_89),
.A2(n_68),
.B(n_36),
.C(n_41),
.D(n_40),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_93),
.Y(n_118)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_118),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_104),
.B(n_73),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_81),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_120),
.B(n_93),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_105),
.B(n_55),
.Y(n_121)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_121),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_96),
.A2(n_63),
.B1(n_69),
.B2(n_70),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_91),
.B(n_55),
.Y(n_125)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_125),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_97),
.A2(n_34),
.B1(n_15),
.B2(n_17),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_100),
.B(n_27),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_127),
.B(n_130),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_102),
.B(n_17),
.Y(n_129)
);

CKINVDCx14_ASAP7_75t_R g151 ( 
.A(n_129),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_90),
.B(n_27),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_90),
.B(n_22),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_131),
.B(n_103),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_135),
.B(n_144),
.C(n_112),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_118),
.A2(n_80),
.B1(n_79),
.B2(n_85),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_136),
.A2(n_146),
.B1(n_147),
.B2(n_120),
.Y(n_162)
);

AO21x2_ASAP7_75t_L g137 ( 
.A1(n_113),
.A2(n_101),
.B(n_98),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_137),
.A2(n_141),
.B1(n_147),
.B2(n_146),
.Y(n_167)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_139),
.Y(n_173)
);

INVx4_ASAP7_75t_L g140 ( 
.A(n_110),
.Y(n_140)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_140),
.Y(n_187)
);

OA22x2_ASAP7_75t_L g141 ( 
.A1(n_122),
.A2(n_82),
.B1(n_87),
.B2(n_80),
.Y(n_141)
);

INVx1_ASAP7_75t_SL g142 ( 
.A(n_117),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_142),
.B(n_145),
.Y(n_182)
);

OAI32xp33_ASAP7_75t_L g183 ( 
.A1(n_143),
.A2(n_153),
.A3(n_134),
.B1(n_141),
.B2(n_160),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_128),
.B(n_94),
.C(n_84),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_125),
.B(n_85),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g146 ( 
.A(n_121),
.Y(n_146)
);

INVxp67_ASAP7_75t_L g147 ( 
.A(n_124),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_SL g149 ( 
.A(n_113),
.B(n_86),
.Y(n_149)
);

CKINVDCx16_ASAP7_75t_R g164 ( 
.A(n_149),
.Y(n_164)
);

INVx13_ASAP7_75t_L g150 ( 
.A(n_110),
.Y(n_150)
);

INVxp67_ASAP7_75t_L g181 ( 
.A(n_150),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_123),
.A2(n_86),
.B1(n_79),
.B2(n_81),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_152),
.A2(n_107),
.B1(n_95),
.B2(n_103),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_130),
.B(n_92),
.Y(n_154)
);

CKINVDCx16_ASAP7_75t_R g190 ( 
.A(n_154),
.Y(n_190)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_156),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_119),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_157),
.Y(n_170)
);

AND2x6_ASAP7_75t_L g158 ( 
.A(n_116),
.B(n_10),
.Y(n_158)
);

A2O1A1O1Ixp25_ASAP7_75t_L g166 ( 
.A1(n_158),
.A2(n_114),
.B(n_137),
.C(n_151),
.D(n_155),
.Y(n_166)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_106),
.Y(n_159)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_159),
.Y(n_175)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_106),
.Y(n_160)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_160),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_162),
.A2(n_171),
.B1(n_177),
.B2(n_178),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_163),
.B(n_165),
.C(n_184),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_144),
.B(n_108),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_166),
.A2(n_167),
.B1(n_168),
.B2(n_174),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_161),
.A2(n_111),
.B1(n_129),
.B2(n_115),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_133),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_172),
.B(n_176),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_137),
.A2(n_127),
.B1(n_109),
.B2(n_126),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_133),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_161),
.A2(n_131),
.B1(n_95),
.B2(n_19),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_137),
.A2(n_142),
.B1(n_141),
.B2(n_159),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_137),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_179)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_179),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_141),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_180)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_180),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_183),
.B(n_158),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_135),
.B(n_29),
.C(n_25),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_138),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_SL g198 ( 
.A(n_186),
.B(n_189),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_148),
.A2(n_19),
.B1(n_25),
.B2(n_7),
.Y(n_188)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_188),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_153),
.Y(n_189)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_156),
.Y(n_191)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_191),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_165),
.B(n_132),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_192),
.B(n_199),
.C(n_213),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_170),
.B(n_152),
.Y(n_193)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_193),
.Y(n_215)
);

BUFx24_ASAP7_75t_SL g194 ( 
.A(n_164),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_194),
.B(n_201),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_169),
.B(n_134),
.Y(n_196)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_196),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_169),
.B(n_155),
.Y(n_197)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_197),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_163),
.B(n_132),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_173),
.B(n_140),
.Y(n_200)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_200),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_187),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_190),
.B(n_150),
.Y(n_203)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_203),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_205),
.B(n_168),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_174),
.B(n_19),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_209),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_191),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_212),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_178),
.B(n_6),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_SL g214 ( 
.A(n_182),
.B(n_7),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_214),
.B(n_11),
.Y(n_226)
);

XNOR2x1_ASAP7_75t_L g216 ( 
.A(n_199),
.B(n_183),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_216),
.A2(n_223),
.B1(n_211),
.B2(n_195),
.Y(n_237)
);

A2O1A1Ixp33_ASAP7_75t_L g217 ( 
.A1(n_196),
.A2(n_166),
.B(n_185),
.C(n_175),
.Y(n_217)
);

CKINVDCx16_ASAP7_75t_R g247 ( 
.A(n_217),
.Y(n_247)
);

HB1xp67_ASAP7_75t_L g219 ( 
.A(n_197),
.Y(n_219)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_219),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_208),
.B(n_184),
.C(n_185),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_220),
.B(n_192),
.C(n_213),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_204),
.A2(n_202),
.B1(n_211),
.B2(n_195),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_SL g238 ( 
.A(n_226),
.B(n_198),
.Y(n_238)
);

HB1xp67_ASAP7_75t_L g228 ( 
.A(n_206),
.Y(n_228)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_228),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_231),
.B(n_207),
.Y(n_242)
);

AOI21xp5_ASAP7_75t_L g232 ( 
.A1(n_205),
.A2(n_167),
.B(n_180),
.Y(n_232)
);

OAI21xp5_ASAP7_75t_L g236 ( 
.A1(n_232),
.A2(n_204),
.B(n_202),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_222),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_233),
.B(n_234),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_220),
.B(n_208),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_235),
.B(n_240),
.C(n_242),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_236),
.B(n_237),
.Y(n_248)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_238),
.Y(n_254)
);

HB1xp67_ASAP7_75t_L g239 ( 
.A(n_225),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_239),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_218),
.B(n_175),
.C(n_207),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_218),
.B(n_210),
.C(n_179),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_243),
.B(n_245),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_L g244 ( 
.A1(n_215),
.A2(n_181),
.B1(n_9),
.B2(n_10),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_244),
.A2(n_226),
.B1(n_224),
.B2(n_230),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_216),
.B(n_181),
.C(n_1),
.Y(n_245)
);

HB1xp67_ASAP7_75t_L g249 ( 
.A(n_246),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_249),
.B(n_13),
.Y(n_269)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_250),
.Y(n_260)
);

INVxp67_ASAP7_75t_L g252 ( 
.A(n_237),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_252),
.B(n_259),
.Y(n_263)
);

NAND2xp33_ASAP7_75t_SL g255 ( 
.A(n_247),
.B(n_217),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_255),
.A2(n_257),
.B1(n_232),
.B2(n_252),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_243),
.A2(n_227),
.B1(n_221),
.B2(n_223),
.Y(n_257)
);

INVxp67_ASAP7_75t_L g259 ( 
.A(n_245),
.Y(n_259)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_254),
.Y(n_261)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_261),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_259),
.B(n_229),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_262),
.B(n_264),
.Y(n_273)
);

AND2x2_ASAP7_75t_L g264 ( 
.A(n_248),
.B(n_242),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g276 ( 
.A(n_265),
.B(n_266),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_258),
.B(n_240),
.C(n_235),
.Y(n_266)
);

OAI21xp5_ASAP7_75t_L g267 ( 
.A1(n_248),
.A2(n_241),
.B(n_231),
.Y(n_267)
);

A2O1A1Ixp33_ASAP7_75t_SL g275 ( 
.A1(n_267),
.A2(n_0),
.B(n_2),
.C(n_3),
.Y(n_275)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_251),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_268),
.B(n_269),
.Y(n_277)
);

HB1xp67_ASAP7_75t_L g270 ( 
.A(n_263),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_270),
.B(n_274),
.Y(n_278)
);

OAI21xp5_ASAP7_75t_SL g271 ( 
.A1(n_260),
.A2(n_256),
.B(n_253),
.Y(n_271)
);

OAI21xp5_ASAP7_75t_SL g284 ( 
.A1(n_271),
.A2(n_11),
.B(n_12),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_SL g274 ( 
.A(n_266),
.B(n_258),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_275),
.B(n_2),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_276),
.B(n_267),
.C(n_264),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_279),
.B(n_11),
.C(n_12),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_277),
.B(n_10),
.Y(n_280)
);

AO21x1_ASAP7_75t_L g287 ( 
.A1(n_280),
.A2(n_284),
.B(n_13),
.Y(n_287)
);

INVxp67_ASAP7_75t_L g281 ( 
.A(n_273),
.Y(n_281)
);

OAI21xp5_ASAP7_75t_L g285 ( 
.A1(n_281),
.A2(n_283),
.B(n_272),
.Y(n_285)
);

AOI21x1_ASAP7_75t_SL g288 ( 
.A1(n_282),
.A2(n_5),
.B(n_3),
.Y(n_288)
);

INVxp67_ASAP7_75t_L g283 ( 
.A(n_275),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_285),
.B(n_286),
.Y(n_289)
);

INVxp67_ASAP7_75t_L g290 ( 
.A(n_287),
.Y(n_290)
);

AOI322xp5_ASAP7_75t_L g291 ( 
.A1(n_289),
.A2(n_278),
.A3(n_281),
.B1(n_288),
.B2(n_3),
.C1(n_4),
.C2(n_5),
.Y(n_291)
);

AO21x2_ASAP7_75t_L g292 ( 
.A1(n_291),
.A2(n_290),
.B(n_4),
.Y(n_292)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_292),
.B(n_5),
.Y(n_293)
);


endmodule