module fake_jpeg_6854_n_341 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_341);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_341;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g16 ( 
.A(n_13),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_5),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_1),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

INVx11_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_0),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_10),
.Y(n_26)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_6),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

INVx1_ASAP7_75t_SL g31 ( 
.A(n_0),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_10),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

INVx11_ASAP7_75t_L g34 ( 
.A(n_19),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_34),
.A2(n_36),
.B1(n_42),
.B2(n_27),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_22),
.Y(n_35)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_35),
.Y(n_63)
);

INVx11_ASAP7_75t_L g36 ( 
.A(n_19),
.Y(n_36)
);

CKINVDCx16_ASAP7_75t_R g37 ( 
.A(n_31),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_37),
.B(n_38),
.Y(n_46)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_24),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_33),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_39),
.B(n_43),
.Y(n_50)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_24),
.Y(n_40)
);

INVx5_ASAP7_75t_L g68 ( 
.A(n_40),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_19),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

INVx11_ASAP7_75t_L g42 ( 
.A(n_19),
.Y(n_42)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_24),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_44),
.B(n_45),
.Y(n_64)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_33),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g47 ( 
.A1(n_36),
.A2(n_25),
.B1(n_18),
.B2(n_17),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_L g86 ( 
.A1(n_47),
.A2(n_54),
.B1(n_72),
.B2(n_73),
.Y(n_86)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_40),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_48),
.B(n_51),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_37),
.A2(n_27),
.B1(n_26),
.B2(n_32),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_49),
.A2(n_58),
.B1(n_59),
.B2(n_62),
.Y(n_76)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_52),
.B(n_60),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_53),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_L g54 ( 
.A1(n_36),
.A2(n_27),
.B1(n_18),
.B2(n_29),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_37),
.B(n_21),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_56),
.B(n_57),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_35),
.B(n_21),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_36),
.A2(n_42),
.B1(n_43),
.B2(n_38),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_42),
.A2(n_25),
.B1(n_18),
.B2(n_17),
.Y(n_59)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_39),
.Y(n_60)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_38),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_61),
.B(n_69),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_42),
.A2(n_25),
.B1(n_29),
.B2(n_17),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_34),
.A2(n_26),
.B1(n_32),
.B2(n_29),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_65),
.A2(n_16),
.B1(n_32),
.B2(n_28),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_38),
.B(n_16),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_66),
.B(n_67),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_43),
.B(n_16),
.Y(n_67)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_43),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_39),
.Y(n_70)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_70),
.Y(n_83)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_39),
.Y(n_71)
);

INVx11_ASAP7_75t_L g96 ( 
.A(n_71),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_L g72 ( 
.A1(n_34),
.A2(n_45),
.B1(n_44),
.B2(n_28),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_34),
.A2(n_21),
.B1(n_28),
.B2(n_26),
.Y(n_73)
);

AO22x1_ASAP7_75t_SL g74 ( 
.A1(n_68),
.A2(n_41),
.B1(n_34),
.B2(n_45),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_74),
.A2(n_58),
.B1(n_72),
.B2(n_48),
.Y(n_106)
);

HB1xp67_ASAP7_75t_L g75 ( 
.A(n_68),
.Y(n_75)
);

CKINVDCx16_ASAP7_75t_R g108 ( 
.A(n_75),
.Y(n_108)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_68),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_77),
.B(n_81),
.Y(n_98)
);

BUFx4f_ASAP7_75t_SL g79 ( 
.A(n_63),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_79),
.Y(n_119)
);

AOI21xp5_ASAP7_75t_L g103 ( 
.A1(n_80),
.A2(n_59),
.B(n_62),
.Y(n_103)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_63),
.Y(n_81)
);

BUFx12f_ASAP7_75t_L g82 ( 
.A(n_63),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_82),
.Y(n_111)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_61),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_84),
.B(n_89),
.Y(n_102)
);

FAx1_ASAP7_75t_SL g85 ( 
.A(n_56),
.B(n_35),
.CI(n_45),
.CON(n_85),
.SN(n_85)
);

NOR2xp33_ASAP7_75t_SL g105 ( 
.A(n_85),
.B(n_49),
.Y(n_105)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_66),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_67),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_90),
.B(n_91),
.Y(n_121)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_69),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_55),
.Y(n_95)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_95),
.Y(n_120)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_71),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_97),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_92),
.B(n_57),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_99),
.B(n_93),
.Y(n_125)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_94),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_100),
.B(n_101),
.Y(n_130)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_78),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_SL g127 ( 
.A1(n_103),
.A2(n_104),
.B(n_114),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_92),
.B(n_64),
.C(n_70),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_105),
.B(n_112),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_106),
.A2(n_110),
.B1(n_31),
.B2(n_91),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_88),
.A2(n_49),
.B1(n_65),
.B2(n_48),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_107),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_L g109 ( 
.A1(n_85),
.A2(n_65),
.B(n_46),
.Y(n_109)
);

AOI21xp5_ASAP7_75t_L g141 ( 
.A1(n_109),
.A2(n_33),
.B(n_20),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_76),
.A2(n_88),
.B1(n_86),
.B2(n_85),
.Y(n_110)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_87),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_74),
.A2(n_51),
.B1(n_52),
.B2(n_47),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_113),
.A2(n_54),
.B1(n_97),
.B2(n_84),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_SL g114 ( 
.A1(n_89),
.A2(n_46),
.B(n_64),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_L g115 ( 
.A1(n_74),
.A2(n_52),
.B1(n_44),
.B2(n_60),
.Y(n_115)
);

OAI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_115),
.A2(n_96),
.B1(n_79),
.B2(n_55),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_83),
.B(n_50),
.C(n_35),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_SL g134 ( 
.A1(n_116),
.A2(n_117),
.B(n_77),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_83),
.B(n_50),
.C(n_35),
.Y(n_117)
);

AOI32xp33_ASAP7_75t_L g118 ( 
.A1(n_74),
.A2(n_44),
.A3(n_35),
.B1(n_53),
.B2(n_60),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_SL g137 ( 
.A(n_118),
.B(n_79),
.C(n_35),
.Y(n_137)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_93),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_122),
.B(n_31),
.Y(n_153)
);

BUFx24_ASAP7_75t_SL g124 ( 
.A(n_90),
.Y(n_124)
);

INVxp67_ASAP7_75t_L g139 ( 
.A(n_124),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_125),
.B(n_131),
.Y(n_173)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_102),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_126),
.B(n_128),
.Y(n_160)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_102),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_99),
.B(n_104),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_121),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_132),
.B(n_135),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_122),
.B(n_73),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_133),
.B(n_144),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_134),
.B(n_148),
.C(n_141),
.Y(n_181)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_121),
.Y(n_135)
);

INVx4_ASAP7_75t_L g136 ( 
.A(n_120),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_SL g174 ( 
.A1(n_136),
.A2(n_138),
.B1(n_120),
.B2(n_111),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_137),
.B(n_117),
.Y(n_165)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_123),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_140),
.A2(n_150),
.B1(n_113),
.B2(n_105),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_SL g159 ( 
.A1(n_141),
.A2(n_149),
.B(n_116),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_98),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_142),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_143),
.A2(n_123),
.B1(n_41),
.B2(n_23),
.Y(n_182)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_98),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_110),
.A2(n_96),
.B1(n_79),
.B2(n_41),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_145),
.A2(n_108),
.B1(n_119),
.B2(n_111),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g147 ( 
.A(n_115),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_147),
.B(n_152),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_104),
.B(n_35),
.Y(n_148)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_148),
.Y(n_154)
);

INVx2_ASAP7_75t_R g149 ( 
.A(n_114),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_109),
.B(n_22),
.Y(n_151)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_151),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_SL g152 ( 
.A(n_107),
.B(n_81),
.Y(n_152)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_153),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_L g155 ( 
.A1(n_149),
.A2(n_103),
.B1(n_118),
.B2(n_106),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g201 ( 
.A(n_155),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_157),
.A2(n_169),
.B1(n_177),
.B2(n_178),
.Y(n_188)
);

OA21x2_ASAP7_75t_L g158 ( 
.A1(n_149),
.A2(n_107),
.B(n_117),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_158),
.B(n_163),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_L g204 ( 
.A1(n_159),
.A2(n_176),
.B(n_181),
.Y(n_204)
);

BUFx12_ASAP7_75t_L g162 ( 
.A(n_138),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_162),
.Y(n_193)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_130),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_SL g197 ( 
.A(n_165),
.B(n_140),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g166 ( 
.A(n_131),
.B(n_116),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_166),
.B(n_180),
.C(n_181),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_129),
.A2(n_112),
.B1(n_101),
.B2(n_100),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_SL g170 ( 
.A(n_130),
.B(n_108),
.Y(n_170)
);

CKINVDCx14_ASAP7_75t_R g190 ( 
.A(n_170),
.Y(n_190)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_133),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_172),
.B(n_175),
.Y(n_187)
);

CKINVDCx16_ASAP7_75t_R g208 ( 
.A(n_174),
.Y(n_208)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_143),
.Y(n_175)
);

AOI21xp5_ASAP7_75t_SL g176 ( 
.A1(n_149),
.A2(n_151),
.B(n_127),
.Y(n_176)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_143),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_178),
.B(n_179),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_142),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g180 ( 
.A(n_127),
.B(n_22),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_182),
.A2(n_145),
.B1(n_140),
.B2(n_128),
.Y(n_198)
);

AOI22x1_ASAP7_75t_R g185 ( 
.A1(n_176),
.A2(n_137),
.B1(n_141),
.B2(n_152),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_SL g221 ( 
.A(n_185),
.B(n_154),
.Y(n_221)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_160),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_186),
.B(n_189),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_L g219 ( 
.A1(n_188),
.A2(n_156),
.B1(n_154),
.B2(n_158),
.Y(n_219)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_164),
.Y(n_189)
);

AOI21xp5_ASAP7_75t_SL g191 ( 
.A1(n_159),
.A2(n_134),
.B(n_125),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_191),
.B(n_196),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_173),
.B(n_146),
.Y(n_192)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_192),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_173),
.B(n_146),
.Y(n_194)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_194),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_172),
.B(n_132),
.Y(n_195)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_195),
.Y(n_218)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_182),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_197),
.B(n_207),
.C(n_163),
.Y(n_222)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_198),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_161),
.B(n_126),
.Y(n_200)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_200),
.Y(n_227)
);

INVxp33_ASAP7_75t_L g202 ( 
.A(n_177),
.Y(n_202)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_202),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_SL g203 ( 
.A(n_167),
.B(n_153),
.Y(n_203)
);

CKINVDCx16_ASAP7_75t_R g217 ( 
.A(n_203),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_204),
.B(n_180),
.Y(n_220)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_168),
.Y(n_205)
);

AOI22xp33_ASAP7_75t_SL g230 ( 
.A1(n_205),
.A2(n_209),
.B1(n_210),
.B2(n_136),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_161),
.B(n_135),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_206),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_SL g207 ( 
.A(n_166),
.B(n_145),
.Y(n_207)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_162),
.Y(n_209)
);

CKINVDCx14_ASAP7_75t_R g210 ( 
.A(n_162),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_207),
.B(n_165),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_212),
.B(n_221),
.Y(n_240)
);

OAI22x1_ASAP7_75t_L g214 ( 
.A1(n_185),
.A2(n_171),
.B1(n_158),
.B2(n_175),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_L g248 ( 
.A1(n_214),
.A2(n_191),
.B1(n_184),
.B2(n_187),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_208),
.A2(n_156),
.B1(n_179),
.B2(n_167),
.Y(n_216)
);

INVxp67_ASAP7_75t_L g258 ( 
.A(n_216),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_219),
.A2(n_224),
.B1(n_232),
.B2(n_235),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_220),
.B(n_222),
.C(n_226),
.Y(n_246)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_209),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_223),
.B(n_228),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_188),
.A2(n_150),
.B1(n_138),
.B2(n_139),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_199),
.B(n_82),
.Y(n_226)
);

BUFx6f_ASAP7_75t_L g228 ( 
.A(n_193),
.Y(n_228)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_230),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_183),
.A2(n_201),
.B1(n_184),
.B2(n_191),
.Y(n_232)
);

BUFx5_ASAP7_75t_L g233 ( 
.A(n_193),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_233),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_183),
.A2(n_136),
.B1(n_41),
.B2(n_95),
.Y(n_235)
);

AO22x2_ASAP7_75t_SL g236 ( 
.A1(n_187),
.A2(n_55),
.B1(n_22),
.B2(n_23),
.Y(n_236)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_236),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_217),
.B(n_194),
.Y(n_239)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_239),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_211),
.B(n_186),
.Y(n_244)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_244),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_225),
.A2(n_232),
.B1(n_229),
.B2(n_234),
.Y(n_245)
);

CKINVDCx14_ASAP7_75t_R g266 ( 
.A(n_245),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_229),
.A2(n_198),
.B1(n_204),
.B2(n_208),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_247),
.A2(n_250),
.B1(n_251),
.B2(n_255),
.Y(n_262)
);

FAx1_ASAP7_75t_SL g265 ( 
.A(n_248),
.B(n_221),
.CI(n_236),
.CON(n_265),
.SN(n_265)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_233),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_249),
.B(n_252),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_231),
.A2(n_196),
.B1(n_205),
.B2(n_190),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_214),
.A2(n_199),
.B1(n_192),
.B2(n_200),
.Y(n_251)
);

CKINVDCx16_ASAP7_75t_R g252 ( 
.A(n_235),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_228),
.B(n_189),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_253),
.Y(n_260)
);

XNOR2x1_ASAP7_75t_L g254 ( 
.A(n_220),
.B(n_197),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_254),
.B(n_256),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_L g255 ( 
.A1(n_218),
.A2(n_203),
.B1(n_195),
.B2(n_206),
.Y(n_255)
);

XNOR2x1_ASAP7_75t_L g256 ( 
.A(n_222),
.B(n_82),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_212),
.B(n_82),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_257),
.B(n_30),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_227),
.B(n_0),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_259),
.B(n_213),
.Y(n_263)
);

OAI21xp5_ASAP7_75t_L g261 ( 
.A1(n_258),
.A2(n_216),
.B(n_215),
.Y(n_261)
);

AOI21xp5_ASAP7_75t_L g291 ( 
.A1(n_261),
.A2(n_268),
.B(n_277),
.Y(n_291)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_263),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_265),
.B(n_275),
.Y(n_283)
);

OAI21xp5_ASAP7_75t_L g268 ( 
.A1(n_258),
.A2(n_236),
.B(n_226),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_237),
.A2(n_223),
.B1(n_95),
.B2(n_55),
.Y(n_270)
);

OAI21xp5_ASAP7_75t_L g296 ( 
.A1(n_270),
.A2(n_274),
.B(n_279),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_241),
.Y(n_272)
);

OAI21xp5_ASAP7_75t_SL g295 ( 
.A1(n_272),
.A2(n_278),
.B(n_2),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_246),
.B(n_22),
.C(n_23),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_273),
.B(n_247),
.C(n_238),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_242),
.A2(n_23),
.B1(n_22),
.B2(n_30),
.Y(n_274)
);

AOI322xp5_ASAP7_75t_L g275 ( 
.A1(n_256),
.A2(n_8),
.A3(n_15),
.B1(n_14),
.B2(n_13),
.C1(n_12),
.C2(n_11),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_276),
.B(n_246),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_239),
.B(n_0),
.Y(n_277)
);

INVxp67_ASAP7_75t_L g278 ( 
.A(n_245),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_238),
.A2(n_30),
.B1(n_20),
.B2(n_3),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_260),
.B(n_243),
.Y(n_280)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_280),
.Y(n_306)
);

AND2x2_ASAP7_75t_L g300 ( 
.A(n_281),
.B(n_276),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_282),
.B(n_284),
.C(n_289),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_273),
.B(n_251),
.C(n_254),
.Y(n_284)
);

INVx3_ASAP7_75t_L g285 ( 
.A(n_266),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_285),
.B(n_261),
.Y(n_301)
);

INVxp33_ASAP7_75t_L g287 ( 
.A(n_263),
.Y(n_287)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_287),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_267),
.B(n_259),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_SL g309 ( 
.A(n_288),
.B(n_290),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_262),
.B(n_257),
.C(n_240),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_270),
.B(n_262),
.Y(n_290)
);

XOR2xp5_ASAP7_75t_L g292 ( 
.A(n_269),
.B(n_240),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_292),
.B(n_269),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_264),
.B(n_20),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_293),
.B(n_294),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_277),
.B(n_1),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_295),
.B(n_274),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_298),
.B(n_300),
.C(n_292),
.Y(n_311)
);

INVx6_ASAP7_75t_L g299 ( 
.A(n_287),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_299),
.B(n_284),
.Y(n_318)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_301),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_302),
.B(n_307),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_L g303 ( 
.A1(n_291),
.A2(n_278),
.B1(n_285),
.B2(n_271),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g319 ( 
.A1(n_303),
.A2(n_308),
.B1(n_310),
.B2(n_9),
.Y(n_319)
);

NAND3xp33_ASAP7_75t_L g304 ( 
.A(n_291),
.B(n_268),
.C(n_265),
.Y(n_304)
);

AND2x2_ASAP7_75t_L g314 ( 
.A(n_304),
.B(n_289),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_282),
.A2(n_279),
.B1(n_265),
.B2(n_9),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_L g310 ( 
.A1(n_286),
.A2(n_8),
.B1(n_14),
.B2(n_12),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_311),
.B(n_297),
.C(n_15),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_SL g312 ( 
.A(n_309),
.B(n_283),
.Y(n_312)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_312),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_SL g313 ( 
.A(n_306),
.B(n_296),
.Y(n_313)
);

OAI21xp5_ASAP7_75t_SL g322 ( 
.A1(n_313),
.A2(n_318),
.B(n_321),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_314),
.B(n_317),
.Y(n_323)
);

OR2x2_ASAP7_75t_L g315 ( 
.A(n_304),
.B(n_296),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_315),
.B(n_319),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_SL g320 ( 
.A1(n_299),
.A2(n_281),
.B1(n_9),
.B2(n_11),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_320),
.B(n_14),
.Y(n_328)
);

OAI21xp5_ASAP7_75t_SL g321 ( 
.A1(n_305),
.A2(n_300),
.B(n_298),
.Y(n_321)
);

XOR2xp5_ASAP7_75t_L g326 ( 
.A(n_318),
.B(n_305),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_326),
.B(n_327),
.C(n_2),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_328),
.B(n_323),
.Y(n_335)
);

A2O1A1Ixp33_ASAP7_75t_L g329 ( 
.A1(n_315),
.A2(n_12),
.B(n_3),
.C(n_4),
.Y(n_329)
);

AOI21xp5_ASAP7_75t_L g332 ( 
.A1(n_329),
.A2(n_316),
.B(n_3),
.Y(n_332)
);

AND2x2_ASAP7_75t_L g330 ( 
.A(n_326),
.B(n_314),
.Y(n_330)
);

A2O1A1O1Ixp25_ASAP7_75t_L g336 ( 
.A1(n_330),
.A2(n_331),
.B(n_322),
.C(n_329),
.D(n_5),
.Y(n_336)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_324),
.Y(n_331)
);

A2O1A1Ixp33_ASAP7_75t_SL g337 ( 
.A1(n_332),
.A2(n_333),
.B(n_334),
.C(n_335),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_SL g334 ( 
.A(n_325),
.B(n_2),
.Y(n_334)
);

OAI31xp33_ASAP7_75t_SL g338 ( 
.A1(n_336),
.A2(n_3),
.A3(n_4),
.B(n_5),
.Y(n_338)
);

OAI321xp33_ASAP7_75t_L g339 ( 
.A1(n_338),
.A2(n_4),
.A3(n_6),
.B1(n_7),
.B2(n_337),
.C(n_332),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_339),
.B(n_4),
.C(n_6),
.Y(n_340)
);

NOR3xp33_ASAP7_75t_SL g341 ( 
.A(n_340),
.B(n_7),
.C(n_338),
.Y(n_341)
);


endmodule