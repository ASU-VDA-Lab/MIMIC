module real_jpeg_27688_n_11 (n_5, n_4, n_8, n_0, n_1, n_2, n_262, n_6, n_7, n_3, n_10, n_9, n_11);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_2;
input n_262;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_11;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_247;
wire n_146;
wire n_83;
wire n_78;
wire n_249;
wire n_215;
wire n_176;
wire n_221;
wire n_166;
wire n_194;
wire n_153;
wire n_104;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_237;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_243;
wire n_173;
wire n_255;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_13;
wire n_120;
wire n_155;
wire n_113;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_242;
wire n_141;
wire n_65;
wire n_33;
wire n_188;
wire n_139;
wire n_142;
wire n_175;
wire n_238;
wire n_76;
wire n_67;
wire n_178;
wire n_79;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_222;
wire n_148;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_258;
wire n_205;
wire n_195;
wire n_110;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_204;
wire n_158;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_241;
wire n_259;
wire n_103;
wire n_225;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_12;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_187;
wire n_97;
wire n_34;
wire n_230;
wire n_190;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_244;
wire n_167;
wire n_202;
wire n_179;
wire n_213;
wire n_133;
wire n_216;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_256;
wire n_101;
wire n_182;
wire n_253;
wire n_96;
wire n_89;
wire n_16;

OAI22xp5_ASAP7_75t_L g29 ( 
.A1(n_0),
.A2(n_17),
.B1(n_18),
.B2(n_30),
.Y(n_29)
);

CKINVDCx16_ASAP7_75t_R g30 ( 
.A(n_0),
.Y(n_30)
);

OAI22xp33_ASAP7_75t_SL g44 ( 
.A1(n_0),
.A2(n_25),
.B1(n_26),
.B2(n_30),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_0),
.A2(n_30),
.B1(n_59),
.B2(n_60),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g209 ( 
.A1(n_0),
.A2(n_30),
.B1(n_49),
.B2(n_50),
.Y(n_209)
);

INVx11_ASAP7_75t_L g95 ( 
.A(n_1),
.Y(n_95)
);

INVx5_ASAP7_75t_L g143 ( 
.A(n_1),
.Y(n_143)
);

BUFx12_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_3),
.Y(n_50)
);

BUFx2_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

OAI22xp5_ASAP7_75t_L g40 ( 
.A1(n_5),
.A2(n_17),
.B1(n_18),
.B2(n_41),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_5),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_5),
.A2(n_41),
.B1(n_49),
.B2(n_50),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_5),
.A2(n_25),
.B1(n_26),
.B2(n_41),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_5),
.A2(n_41),
.B1(n_59),
.B2(n_60),
.Y(n_97)
);

AOI21xp33_ASAP7_75t_SL g106 ( 
.A1(n_5),
.A2(n_22),
.B(n_26),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_5),
.B(n_32),
.Y(n_120)
);

AOI21xp33_ASAP7_75t_L g129 ( 
.A1(n_5),
.A2(n_6),
.B(n_60),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_5),
.B(n_134),
.Y(n_133)
);

O2A1O1Ixp33_ASAP7_75t_L g152 ( 
.A1(n_5),
.A2(n_8),
.B(n_25),
.C(n_153),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g58 ( 
.A1(n_6),
.A2(n_59),
.B1(n_60),
.B2(n_62),
.Y(n_58)
);

INVx11_ASAP7_75t_L g62 ( 
.A(n_6),
.Y(n_62)
);

BUFx24_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_8),
.Y(n_48)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_8),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g15 ( 
.A1(n_9),
.A2(n_16),
.B1(n_17),
.B2(n_18),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_9),
.Y(n_16)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_9),
.A2(n_16),
.B1(n_25),
.B2(n_26),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_9),
.A2(n_16),
.B1(n_49),
.B2(n_50),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g190 ( 
.A1(n_9),
.A2(n_16),
.B1(n_59),
.B2(n_60),
.Y(n_190)
);

INVx11_ASAP7_75t_SL g61 ( 
.A(n_10),
.Y(n_61)
);

XOR2xp5_ASAP7_75t_L g11 ( 
.A(n_12),
.B(n_35),
.Y(n_11)
);

NAND2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_33),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_27),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_14),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_19),
.Y(n_14)
);

AOI22xp5_ASAP7_75t_L g28 ( 
.A1(n_15),
.A2(n_29),
.B1(n_31),
.B2(n_32),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_17),
.Y(n_18)
);

OAI22xp5_ASAP7_75t_L g21 ( 
.A1(n_17),
.A2(n_18),
.B1(n_22),
.B2(n_23),
.Y(n_21)
);

A2O1A1Ixp33_ASAP7_75t_L g105 ( 
.A1(n_17),
.A2(n_23),
.B(n_41),
.C(n_106),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g39 ( 
.A(n_19),
.B(n_40),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_24),
.Y(n_19)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_20),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_24),
.Y(n_20)
);

CKINVDCx14_ASAP7_75t_R g23 ( 
.A(n_22),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_SL g24 ( 
.A1(n_22),
.A2(n_23),
.B1(n_25),
.B2(n_26),
.Y(n_24)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_24),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_25),
.A2(n_26),
.B1(n_47),
.B2(n_51),
.Y(n_52)
);

INVx8_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_28),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_28),
.B(n_34),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_28),
.B(n_37),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_28),
.B(n_37),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_29),
.A2(n_31),
.B1(n_32),
.B2(n_40),
.Y(n_67)
);

OAI21xp5_ASAP7_75t_L g35 ( 
.A1(n_36),
.A2(n_72),
.B(n_259),
.Y(n_35)
);

MAJIxp5_ASAP7_75t_L g37 ( 
.A(n_38),
.B(n_67),
.C(n_68),
.Y(n_37)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_38),
.B(n_256),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g38 ( 
.A(n_39),
.B(n_42),
.C(n_54),
.Y(n_38)
);

AOI211xp5_ASAP7_75t_L g81 ( 
.A1(n_39),
.A2(n_82),
.B(n_84),
.C(n_89),
.Y(n_81)
);

CKINVDCx16_ASAP7_75t_R g90 ( 
.A(n_39),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_39),
.A2(n_85),
.B1(n_86),
.B2(n_90),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_39),
.A2(n_90),
.B1(n_114),
.B2(n_115),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_39),
.A2(n_90),
.B1(n_204),
.B2(n_205),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_39),
.A2(n_90),
.B1(n_234),
.B2(n_235),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_L g239 ( 
.A1(n_39),
.A2(n_204),
.B(n_224),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_39),
.A2(n_90),
.B1(n_242),
.B2(n_246),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_39),
.A2(n_90),
.B1(n_243),
.B2(n_244),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_39),
.B(n_54),
.C(n_237),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_39),
.B(n_246),
.C(n_247),
.Y(n_254)
);

A2O1A1Ixp33_ASAP7_75t_L g128 ( 
.A1(n_41),
.A2(n_50),
.B(n_62),
.C(n_129),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g139 ( 
.A(n_41),
.B(n_58),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_41),
.B(n_143),
.Y(n_142)
);

OAI21xp33_ASAP7_75t_L g153 ( 
.A1(n_41),
.A2(n_49),
.B(n_51),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_42),
.A2(n_54),
.B1(n_55),
.B2(n_245),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_42),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_L g42 ( 
.A1(n_43),
.A2(n_45),
.B1(n_46),
.B2(n_53),
.Y(n_42)
);

CKINVDCx16_ASAP7_75t_R g43 ( 
.A(n_44),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_44),
.A2(n_87),
.B1(n_134),
.B2(n_238),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_45),
.B(n_46),
.Y(n_71)
);

INVxp67_ASAP7_75t_L g238 ( 
.A(n_45),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_46),
.B(n_52),
.Y(n_45)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_46),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g46 ( 
.A1(n_47),
.A2(n_49),
.B1(n_50),
.B2(n_51),
.Y(n_46)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_49),
.A2(n_50),
.B1(n_62),
.B2(n_65),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_50),
.Y(n_49)
);

CKINVDCx16_ASAP7_75t_R g70 ( 
.A(n_53),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_54),
.A2(n_55),
.B1(n_236),
.B2(n_237),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_55),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g55 ( 
.A(n_56),
.B(n_66),
.Y(n_55)
);

INVxp33_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

AND2x2_ASAP7_75t_SL g82 ( 
.A(n_57),
.B(n_83),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_58),
.B(n_63),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_58),
.B(n_64),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_58),
.A2(n_63),
.B1(n_208),
.B2(n_209),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_58),
.A2(n_63),
.B1(n_66),
.B2(n_209),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_SL g141 ( 
.A(n_59),
.B(n_142),
.Y(n_141)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_60),
.B(n_95),
.Y(n_94)
);

INVx5_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx11_ASAP7_75t_L g65 ( 
.A(n_62),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g256 ( 
.A1(n_67),
.A2(n_68),
.B1(n_69),
.B2(n_257),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_67),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_69),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_70),
.B(n_71),
.Y(n_69)
);

AND2x2_ASAP7_75t_SL g86 ( 
.A(n_71),
.B(n_87),
.Y(n_86)
);

AOI21xp5_ASAP7_75t_L g72 ( 
.A1(n_73),
.A2(n_253),
.B(n_258),
.Y(n_72)
);

OAI321xp33_ASAP7_75t_L g73 ( 
.A1(n_74),
.A2(n_231),
.A3(n_248),
.B1(n_251),
.B2(n_252),
.C(n_262),
.Y(n_73)
);

AOI21xp5_ASAP7_75t_L g74 ( 
.A1(n_75),
.A2(n_215),
.B(n_230),
.Y(n_74)
);

OAI21xp5_ASAP7_75t_SL g75 ( 
.A1(n_76),
.A2(n_196),
.B(n_214),
.Y(n_75)
);

O2A1O1Ixp33_ASAP7_75t_SL g76 ( 
.A1(n_77),
.A2(n_121),
.B(n_178),
.C(n_195),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_111),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_78),
.B(n_111),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_100),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_80),
.A2(n_81),
.B1(n_91),
.B2(n_92),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_80),
.B(n_92),
.C(n_100),
.Y(n_179)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_82),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_82),
.A2(n_88),
.B1(n_93),
.B2(n_99),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_82),
.A2(n_85),
.B1(n_86),
.B2(n_88),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_82),
.A2(n_88),
.B1(n_132),
.B2(n_133),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_82),
.A2(n_88),
.B1(n_128),
.B2(n_146),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_82),
.B(n_107),
.C(n_132),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_82),
.A2(n_88),
.B1(n_167),
.B2(n_168),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_82),
.B(n_161),
.C(n_167),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_82),
.B(n_93),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_82),
.A2(n_88),
.B1(n_186),
.B2(n_187),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_82),
.B(n_187),
.Y(n_201)
);

INVxp67_ASAP7_75t_L g208 ( 
.A(n_83),
.Y(n_208)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_84),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_88),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_85),
.B(n_90),
.Y(n_89)
);

A2O1A1Ixp33_ASAP7_75t_L g158 ( 
.A1(n_85),
.A2(n_88),
.B(n_155),
.C(n_159),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_85),
.A2(n_86),
.B1(n_163),
.B2(n_164),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_85),
.B(n_90),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_86),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_86),
.B(n_107),
.C(n_119),
.Y(n_118)
);

AOI21xp5_ASAP7_75t_L g220 ( 
.A1(n_86),
.A2(n_221),
.B(n_222),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_86),
.B(n_221),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_88),
.B(n_128),
.Y(n_127)
);

AOI21xp5_ASAP7_75t_L g193 ( 
.A1(n_89),
.A2(n_110),
.B(n_194),
.Y(n_193)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_89),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_92),
.Y(n_91)
);

CKINVDCx14_ASAP7_75t_R g99 ( 
.A(n_93),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_94),
.A2(n_95),
.B1(n_96),
.B2(n_98),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_94),
.B(n_95),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_94),
.A2(n_98),
.B1(n_188),
.B2(n_190),
.Y(n_187)
);

INVx11_ASAP7_75t_L g189 ( 
.A(n_95),
.Y(n_189)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_97),
.B(n_109),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_101),
.A2(n_102),
.B1(n_103),
.B2(n_110),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_101),
.A2(n_102),
.B1(n_183),
.B2(n_184),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_101),
.A2(n_102),
.B1(n_201),
.B2(n_202),
.Y(n_200)
);

CKINVDCx16_ASAP7_75t_R g101 ( 
.A(n_102),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_103),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_107),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_104),
.A2(n_105),
.B1(n_107),
.B2(n_108),
.Y(n_117)
);

CKINVDCx16_ASAP7_75t_R g104 ( 
.A(n_105),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_107),
.A2(n_108),
.B1(n_131),
.B2(n_135),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_107),
.B(n_139),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_107),
.B(n_141),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_107),
.A2(n_108),
.B1(n_152),
.B2(n_154),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_107),
.A2(n_108),
.B1(n_119),
.B2(n_120),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_107),
.B(n_152),
.Y(n_168)
);

INVx1_ASAP7_75t_SL g107 ( 
.A(n_108),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g144 ( 
.A(n_108),
.B(n_145),
.Y(n_144)
);

INVxp33_ASAP7_75t_L g206 ( 
.A(n_109),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_112),
.B(n_116),
.C(n_118),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_112),
.A2(n_113),
.B1(n_173),
.B2(n_175),
.Y(n_172)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

CKINVDCx16_ASAP7_75t_R g115 ( 
.A(n_114),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_114),
.A2(n_115),
.B1(n_151),
.B2(n_155),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_116),
.A2(n_117),
.B1(n_118),
.B2(n_174),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_117),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_118),
.Y(n_174)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g121 ( 
.A(n_122),
.B(n_177),
.Y(n_121)
);

AOI21xp5_ASAP7_75t_L g122 ( 
.A1(n_123),
.A2(n_170),
.B(n_176),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_SL g123 ( 
.A1(n_124),
.A2(n_157),
.B(n_169),
.Y(n_123)
);

AOI21xp5_ASAP7_75t_L g124 ( 
.A1(n_125),
.A2(n_148),
.B(n_156),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_SL g125 ( 
.A1(n_126),
.A2(n_136),
.B(n_147),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_130),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_127),
.B(n_130),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_128),
.Y(n_146)
);

CKINVDCx16_ASAP7_75t_R g135 ( 
.A(n_131),
.Y(n_135)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_144),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_140),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_150),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_149),
.B(n_150),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_151),
.Y(n_155)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_152),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_160),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_158),
.B(n_160),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_161),
.A2(n_162),
.B1(n_165),
.B2(n_166),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_164),
.Y(n_163)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_168),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_172),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_171),
.B(n_172),
.Y(n_176)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_173),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_180),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_SL g195 ( 
.A(n_179),
.B(n_180),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_193),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_182),
.A2(n_185),
.B1(n_191),
.B2(n_192),
.Y(n_181)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_182),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_183),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_L g211 ( 
.A1(n_183),
.A2(n_212),
.B(n_213),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_185),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_185),
.B(n_191),
.C(n_193),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_187),
.Y(n_186)
);

INVx11_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_190),
.B(n_206),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_194),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_198),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_197),
.B(n_198),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_211),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_203),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_200),
.B(n_203),
.C(n_211),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_201),
.Y(n_202)
);

OAI21xp33_ASAP7_75t_L g228 ( 
.A1(n_201),
.A2(n_212),
.B(n_213),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_204),
.A2(n_205),
.B1(n_207),
.B2(n_210),
.Y(n_203)
);

CKINVDCx16_ASAP7_75t_R g204 ( 
.A(n_205),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_205),
.B(n_207),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_207),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_217),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_SL g230 ( 
.A(n_216),
.B(n_217),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_218),
.A2(n_219),
.B1(n_228),
.B2(n_229),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_223),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_220),
.B(n_223),
.C(n_229),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_222),
.B(n_233),
.C(n_239),
.Y(n_232)
);

FAx1_ASAP7_75t_SL g250 ( 
.A(n_222),
.B(n_233),
.CI(n_239),
.CON(n_250),
.SN(n_250)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_224),
.A2(n_225),
.B1(n_226),
.B2(n_227),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_225),
.Y(n_224)
);

CKINVDCx16_ASAP7_75t_R g227 ( 
.A(n_226),
.Y(n_227)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_228),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_240),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_232),
.B(n_240),
.Y(n_252)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_237),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_247),
.Y(n_240)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_242),
.Y(n_246)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_250),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_249),
.B(n_250),
.Y(n_251)
);

BUFx24_ASAP7_75t_SL g260 ( 
.A(n_250),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_254),
.B(n_255),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_254),
.B(n_255),
.Y(n_258)
);


endmodule