module fake_jpeg_3019_n_29 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_29);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_29;

wire n_13;
wire n_21;
wire n_23;
wire n_10;
wire n_27;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_11;
wire n_17;
wire n_25;
wire n_12;
wire n_15;

NOR2xp33_ASAP7_75t_SL g10 ( 
.A(n_6),
.B(n_3),
.Y(n_10)
);

NOR2xp33_ASAP7_75t_SL g11 ( 
.A(n_5),
.B(n_3),
.Y(n_11)
);

INVx6_ASAP7_75t_SL g12 ( 
.A(n_4),
.Y(n_12)
);

INVx2_ASAP7_75t_L g13 ( 
.A(n_2),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_4),
.Y(n_14)
);

BUFx12f_ASAP7_75t_SL g15 ( 
.A(n_7),
.Y(n_15)
);

INVx8_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_0),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_13),
.B(n_0),
.Y(n_18)
);

AOI22xp33_ASAP7_75t_L g22 ( 
.A1(n_18),
.A2(n_20),
.B1(n_21),
.B2(n_12),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_SL g19 ( 
.A1(n_13),
.A2(n_1),
.B1(n_2),
.B2(n_8),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_SL g23 ( 
.A1(n_19),
.A2(n_17),
.B1(n_14),
.B2(n_16),
.Y(n_23)
);

INVx1_ASAP7_75t_SL g20 ( 
.A(n_12),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_22),
.Y(n_24)
);

AOI21xp5_ASAP7_75t_SL g25 ( 
.A1(n_24),
.A2(n_21),
.B(n_15),
.Y(n_25)
);

OAI21xp5_ASAP7_75t_L g26 ( 
.A1(n_25),
.A2(n_20),
.B(n_23),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_26),
.B(n_1),
.Y(n_28)
);

MAJIxp5_ASAP7_75t_L g27 ( 
.A(n_26),
.B(n_23),
.C(n_17),
.Y(n_27)
);

O2A1O1Ixp33_ASAP7_75t_SL g29 ( 
.A1(n_27),
.A2(n_28),
.B(n_10),
.C(n_11),
.Y(n_29)
);


endmodule