module fake_jpeg_11594_n_50 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_50);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_50;

wire n_13;
wire n_21;
wire n_33;
wire n_45;
wire n_23;
wire n_10;
wire n_27;
wire n_22;
wire n_47;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_12;
wire n_32;
wire n_8;
wire n_15;

BUFx6f_ASAP7_75t_L g8 ( 
.A(n_6),
.Y(n_8)
);

CKINVDCx20_ASAP7_75t_R g9 ( 
.A(n_5),
.Y(n_9)
);

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_0),
.Y(n_10)
);

NOR2xp33_ASAP7_75t_L g11 ( 
.A(n_3),
.B(n_4),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_6),
.Y(n_12)
);

INVx3_ASAP7_75t_L g13 ( 
.A(n_2),
.Y(n_13)
);

INVx6_ASAP7_75t_L g14 ( 
.A(n_3),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_2),
.Y(n_15)
);

BUFx3_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

INVx3_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_11),
.B(n_15),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_SL g36 ( 
.A(n_18),
.B(n_27),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_SL g19 ( 
.A1(n_17),
.A2(n_0),
.B1(n_1),
.B2(n_4),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_L g33 ( 
.A1(n_19),
.A2(n_25),
.B1(n_26),
.B2(n_29),
.Y(n_33)
);

AND2x2_ASAP7_75t_L g20 ( 
.A(n_17),
.B(n_0),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_20),
.B(n_23),
.Y(n_37)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_21),
.Y(n_32)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_22),
.Y(n_35)
);

INVxp67_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

INVx11_ASAP7_75t_L g24 ( 
.A(n_16),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_24),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_L g25 ( 
.A1(n_14),
.A2(n_1),
.B1(n_7),
.B2(n_8),
.Y(n_25)
);

OA22x2_ASAP7_75t_L g26 ( 
.A1(n_8),
.A2(n_7),
.B1(n_10),
.B2(n_9),
.Y(n_26)
);

INVxp67_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_16),
.Y(n_28)
);

OAI21xp5_ASAP7_75t_L g34 ( 
.A1(n_28),
.A2(n_30),
.B(n_24),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_SL g29 ( 
.A1(n_14),
.A2(n_8),
.B1(n_10),
.B2(n_12),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_12),
.B(n_9),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_34),
.B(n_20),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_38),
.B(n_40),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_L g39 ( 
.A1(n_33),
.A2(n_20),
.B1(n_26),
.B2(n_28),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g42 ( 
.A1(n_39),
.A2(n_34),
.B1(n_26),
.B2(n_37),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_SL g40 ( 
.A(n_36),
.B(n_27),
.Y(n_40)
);

MAJIxp5_ASAP7_75t_L g45 ( 
.A(n_42),
.B(n_26),
.C(n_32),
.Y(n_45)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_39),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g44 ( 
.A1(n_43),
.A2(n_32),
.B1(n_35),
.B2(n_23),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_44),
.B(n_31),
.Y(n_47)
);

MAJIxp5_ASAP7_75t_L g46 ( 
.A(n_45),
.B(n_42),
.C(n_43),
.Y(n_46)
);

OAI21xp5_ASAP7_75t_SL g48 ( 
.A1(n_46),
.A2(n_47),
.B(n_41),
.Y(n_48)
);

INVxp67_ASAP7_75t_L g49 ( 
.A(n_48),
.Y(n_49)
);

XNOR2xp5_ASAP7_75t_L g50 ( 
.A(n_49),
.B(n_31),
.Y(n_50)
);


endmodule