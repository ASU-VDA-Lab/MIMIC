module fake_jpeg_5663_n_328 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_328);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_328;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_13;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_145;
wire n_18;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_5),
.Y(n_13)
);

INVx6_ASAP7_75t_SL g14 ( 
.A(n_11),
.Y(n_14)
);

INVx2_ASAP7_75t_L g15 ( 
.A(n_10),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_4),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_7),
.Y(n_19)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_1),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

INVx11_ASAP7_75t_SL g26 ( 
.A(n_0),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_26),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_28),
.B(n_29),
.Y(n_43)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_26),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_30),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_13),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_SL g42 ( 
.A(n_31),
.B(n_32),
.Y(n_42)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_33),
.B(n_34),
.Y(n_48)
);

INVx13_ASAP7_75t_L g34 ( 
.A(n_22),
.Y(n_34)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_35),
.B(n_36),
.Y(n_53)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_13),
.Y(n_37)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_37),
.Y(n_41)
);

INVxp67_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_38),
.Y(n_44)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

INVx11_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_38),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_45),
.B(n_54),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_30),
.Y(n_46)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_46),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_47),
.Y(n_60)
);

BUFx2_ASAP7_75t_L g49 ( 
.A(n_30),
.Y(n_49)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_49),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_50),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_29),
.Y(n_51)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_51),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_35),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_52),
.Y(n_62)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_29),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_34),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_55),
.B(n_34),
.Y(n_76)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_36),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_56),
.B(n_36),
.Y(n_71)
);

A2O1A1Ixp33_ASAP7_75t_L g58 ( 
.A1(n_42),
.A2(n_37),
.B(n_31),
.C(n_23),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_58),
.B(n_59),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_42),
.Y(n_59)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_51),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_63),
.B(n_74),
.Y(n_91)
);

OR2x2_ASAP7_75t_SL g64 ( 
.A(n_41),
.B(n_37),
.Y(n_64)
);

OAI21xp33_ASAP7_75t_L g79 ( 
.A1(n_64),
.A2(n_72),
.B(n_32),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_43),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_66),
.Y(n_83)
);

AOI21xp33_ASAP7_75t_SL g70 ( 
.A1(n_44),
.A2(n_15),
.B(n_36),
.Y(n_70)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_70),
.B(n_53),
.C(n_32),
.Y(n_81)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_71),
.Y(n_87)
);

NOR2xp67_ASAP7_75t_L g72 ( 
.A(n_44),
.B(n_31),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_47),
.Y(n_73)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_73),
.Y(n_101)
);

CKINVDCx16_ASAP7_75t_R g74 ( 
.A(n_48),
.Y(n_74)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_49),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_75),
.B(n_52),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_76),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_41),
.B(n_15),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_77),
.B(n_78),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_43),
.B(n_15),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g103 ( 
.A(n_79),
.B(n_80),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_78),
.B(n_40),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_81),
.B(n_89),
.C(n_28),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_60),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_82),
.Y(n_104)
);

OAI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_72),
.A2(n_39),
.B1(n_36),
.B2(n_56),
.Y(n_84)
);

CKINVDCx16_ASAP7_75t_R g106 ( 
.A(n_84),
.Y(n_106)
);

INVx1_ASAP7_75t_SL g85 ( 
.A(n_70),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_85),
.B(n_90),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_74),
.A2(n_39),
.B1(n_45),
.B2(n_32),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_86),
.A2(n_61),
.B1(n_57),
.B2(n_75),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_64),
.B(n_55),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_88),
.B(n_69),
.Y(n_111)
);

AOI32xp33_ASAP7_75t_L g89 ( 
.A1(n_66),
.A2(n_39),
.A3(n_49),
.B1(n_46),
.B2(n_33),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_77),
.Y(n_90)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_92),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_59),
.A2(n_20),
.B1(n_23),
.B2(n_33),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_94),
.A2(n_96),
.B1(n_57),
.B2(n_20),
.Y(n_110)
);

INVx5_ASAP7_75t_L g95 ( 
.A(n_68),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_95),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_58),
.A2(n_71),
.B1(n_20),
.B2(n_23),
.Y(n_96)
);

HB1xp67_ASAP7_75t_L g97 ( 
.A(n_61),
.Y(n_97)
);

CKINVDCx16_ASAP7_75t_R g119 ( 
.A(n_97),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_76),
.B(n_34),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g105 ( 
.A(n_98),
.B(n_69),
.Y(n_105)
);

BUFx24_ASAP7_75t_SL g102 ( 
.A(n_83),
.Y(n_102)
);

CKINVDCx16_ASAP7_75t_R g147 ( 
.A(n_102),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_105),
.B(n_118),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_107),
.A2(n_124),
.B1(n_54),
.B2(n_101),
.Y(n_138)
);

BUFx3_ASAP7_75t_L g108 ( 
.A(n_95),
.Y(n_108)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_108),
.Y(n_131)
);

BUFx12f_ASAP7_75t_L g109 ( 
.A(n_97),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_109),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_110),
.A2(n_93),
.B1(n_91),
.B2(n_89),
.Y(n_135)
);

OAI21xp33_ASAP7_75t_L g144 ( 
.A1(n_111),
.A2(n_34),
.B(n_22),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_100),
.B(n_65),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_112),
.B(n_115),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_L g140 ( 
.A1(n_113),
.A2(n_94),
.B(n_98),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_100),
.B(n_65),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_90),
.B(n_63),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_116),
.B(n_87),
.Y(n_133)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_92),
.Y(n_118)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_80),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_120),
.B(n_123),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_93),
.B(n_68),
.Y(n_122)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_122),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_83),
.B(n_19),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_87),
.A2(n_20),
.B1(n_23),
.B2(n_22),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_120),
.B(n_81),
.C(n_85),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_125),
.B(n_140),
.C(n_28),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_106),
.A2(n_99),
.B1(n_96),
.B2(n_80),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_128),
.B(n_150),
.Y(n_159)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_112),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_129),
.B(n_130),
.Y(n_154)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_115),
.Y(n_130)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_133),
.Y(n_152)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_116),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_134),
.B(n_136),
.Y(n_160)
);

CKINVDCx14_ASAP7_75t_R g175 ( 
.A(n_135),
.Y(n_175)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_110),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_117),
.B(n_99),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_137),
.B(n_139),
.Y(n_156)
);

INVxp67_ASAP7_75t_L g167 ( 
.A(n_138),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_111),
.B(n_88),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_103),
.B(n_91),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_143),
.B(n_17),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_144),
.B(n_24),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_114),
.B(n_62),
.Y(n_145)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_145),
.Y(n_161)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_105),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_146),
.B(n_119),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_106),
.A2(n_28),
.B1(n_101),
.B2(n_13),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_148),
.A2(n_121),
.B1(n_60),
.B2(n_67),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_114),
.B(n_62),
.Y(n_149)
);

CKINVDCx16_ASAP7_75t_R g153 ( 
.A(n_149),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_113),
.A2(n_103),
.B1(n_118),
.B2(n_123),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_142),
.B(n_24),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_151),
.B(n_164),
.Y(n_188)
);

AND2x2_ASAP7_75t_L g155 ( 
.A(n_143),
.B(n_19),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_SL g189 ( 
.A1(n_155),
.A2(n_157),
.B(n_158),
.Y(n_189)
);

NAND2xp33_ASAP7_75t_SL g157 ( 
.A(n_135),
.B(n_140),
.Y(n_157)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_162),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_133),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_163),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_SL g164 ( 
.A(n_142),
.B(n_24),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_L g165 ( 
.A1(n_136),
.A2(n_119),
.B1(n_19),
.B2(n_17),
.Y(n_165)
);

OAI22xp33_ASAP7_75t_SL g190 ( 
.A1(n_165),
.A2(n_178),
.B1(n_131),
.B2(n_148),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_126),
.B(n_108),
.Y(n_166)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_166),
.Y(n_182)
);

INVxp67_ASAP7_75t_L g168 ( 
.A(n_145),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_168),
.B(n_169),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_SL g169 ( 
.A(n_146),
.B(n_17),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_170),
.B(n_171),
.C(n_132),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_125),
.B(n_109),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_172),
.B(n_174),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_132),
.B(n_109),
.Y(n_173)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_173),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_127),
.Y(n_174)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_131),
.Y(n_176)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_176),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_127),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_177),
.B(n_73),
.Y(n_200)
);

CKINVDCx16_ASAP7_75t_R g179 ( 
.A(n_166),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_179),
.B(n_152),
.Y(n_214)
);

INVxp67_ASAP7_75t_L g180 ( 
.A(n_162),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_180),
.B(n_178),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_175),
.A2(n_134),
.B1(n_130),
.B2(n_129),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_183),
.A2(n_187),
.B1(n_155),
.B2(n_152),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_184),
.B(n_185),
.C(n_186),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_171),
.B(n_150),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_170),
.B(n_128),
.C(n_139),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_160),
.A2(n_137),
.B1(n_141),
.B2(n_126),
.Y(n_187)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_190),
.Y(n_212)
);

INVx5_ASAP7_75t_L g193 ( 
.A(n_176),
.Y(n_193)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_193),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_159),
.B(n_141),
.C(n_149),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_194),
.B(n_203),
.C(n_186),
.Y(n_221)
);

AOI21xp5_ASAP7_75t_L g197 ( 
.A1(n_160),
.A2(n_109),
.B(n_62),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_L g211 ( 
.A1(n_197),
.A2(n_161),
.B(n_177),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_163),
.A2(n_121),
.B1(n_18),
.B2(n_25),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_199),
.A2(n_153),
.B1(n_161),
.B2(n_174),
.Y(n_208)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_200),
.Y(n_213)
);

OA21x2_ASAP7_75t_L g201 ( 
.A1(n_157),
.A2(n_121),
.B(n_50),
.Y(n_201)
);

OA21x2_ASAP7_75t_L g227 ( 
.A1(n_201),
.A2(n_50),
.B(n_47),
.Y(n_227)
);

HB1xp67_ASAP7_75t_L g202 ( 
.A(n_153),
.Y(n_202)
);

CKINVDCx16_ASAP7_75t_R g209 ( 
.A(n_202),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_173),
.B(n_147),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_156),
.B(n_147),
.Y(n_204)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_204),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_156),
.B(n_0),
.Y(n_205)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_205),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_200),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_207),
.B(n_219),
.Y(n_241)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_208),
.Y(n_231)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_210),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_211),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_214),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_196),
.B(n_154),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_215),
.B(n_222),
.Y(n_243)
);

AND2x2_ASAP7_75t_L g216 ( 
.A(n_191),
.B(n_172),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_216),
.A2(n_187),
.B1(n_180),
.B2(n_195),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_181),
.A2(n_167),
.B1(n_155),
.B2(n_158),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_218),
.A2(n_224),
.B1(n_189),
.B2(n_198),
.Y(n_236)
);

INVxp67_ASAP7_75t_L g219 ( 
.A(n_193),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_220),
.B(n_221),
.C(n_194),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_196),
.B(n_154),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_192),
.A2(n_164),
.B1(n_151),
.B2(n_169),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_205),
.B(n_0),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_225),
.B(n_227),
.Y(n_247)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_195),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_228),
.A2(n_192),
.B1(n_197),
.B2(n_199),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_217),
.B(n_185),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_229),
.B(n_232),
.C(n_237),
.Y(n_254)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_230),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_217),
.B(n_184),
.Y(n_232)
);

AND2x2_ASAP7_75t_L g250 ( 
.A(n_236),
.B(n_216),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_221),
.B(n_189),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_238),
.B(n_239),
.C(n_245),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_211),
.B(n_203),
.Y(n_239)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_240),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_210),
.A2(n_201),
.B1(n_183),
.B2(n_182),
.Y(n_242)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_242),
.Y(n_263)
);

XOR2x2_ASAP7_75t_SL g244 ( 
.A(n_223),
.B(n_201),
.Y(n_244)
);

A2O1A1O1Ixp25_ASAP7_75t_L g255 ( 
.A1(n_244),
.A2(n_216),
.B(n_227),
.C(n_218),
.D(n_223),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_213),
.B(n_204),
.C(n_188),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_L g246 ( 
.A1(n_212),
.A2(n_104),
.B1(n_82),
.B2(n_67),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_246),
.B(n_227),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_220),
.A2(n_104),
.B1(n_82),
.B2(n_67),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_248),
.A2(n_219),
.B1(n_206),
.B2(n_226),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_213),
.B(n_104),
.C(n_60),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_249),
.B(n_18),
.C(n_25),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_250),
.A2(n_256),
.B1(n_266),
.B2(n_234),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_238),
.B(n_224),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_251),
.B(n_260),
.Y(n_279)
);

INVxp67_ASAP7_75t_L g252 ( 
.A(n_248),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_252),
.B(n_257),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_235),
.B(n_209),
.Y(n_253)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_253),
.Y(n_269)
);

NAND3xp33_ASAP7_75t_SL g277 ( 
.A(n_255),
.B(n_259),
.C(n_249),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_242),
.B(n_206),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_258),
.B(n_264),
.Y(n_273)
);

OAI31xp33_ASAP7_75t_SL g259 ( 
.A1(n_244),
.A2(n_226),
.A3(n_225),
.B(n_18),
.Y(n_259)
);

BUFx24_ASAP7_75t_SL g264 ( 
.A(n_232),
.Y(n_264)
);

INVxp67_ASAP7_75t_SL g265 ( 
.A(n_241),
.Y(n_265)
);

CKINVDCx14_ASAP7_75t_R g275 ( 
.A(n_265),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_233),
.A2(n_25),
.B1(n_21),
.B2(n_27),
.Y(n_266)
);

CKINVDCx14_ASAP7_75t_R g280 ( 
.A(n_267),
.Y(n_280)
);

OAI221xp5_ASAP7_75t_L g268 ( 
.A1(n_265),
.A2(n_230),
.B1(n_247),
.B2(n_243),
.C(n_239),
.Y(n_268)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_268),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_261),
.B(n_245),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_271),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_L g286 ( 
.A1(n_272),
.A2(n_283),
.B1(n_254),
.B2(n_27),
.Y(n_286)
);

INVx1_ASAP7_75t_SL g274 ( 
.A(n_259),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_274),
.B(n_1),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_263),
.A2(n_231),
.B1(n_237),
.B2(n_236),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_276),
.B(n_278),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_277),
.B(n_2),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_262),
.A2(n_229),
.B1(n_11),
.B2(n_12),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_279),
.B(n_27),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_L g281 ( 
.A1(n_252),
.A2(n_52),
.B1(n_25),
.B2(n_21),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_SL g289 ( 
.A(n_281),
.B(n_1),
.Y(n_289)
);

OA21x2_ASAP7_75t_SL g282 ( 
.A1(n_250),
.A2(n_21),
.B(n_18),
.Y(n_282)
);

AOI221xp5_ASAP7_75t_L g292 ( 
.A1(n_282),
.A2(n_27),
.B1(n_16),
.B2(n_4),
.C(n_5),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_255),
.A2(n_21),
.B1(n_18),
.B2(n_27),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_275),
.A2(n_280),
.B1(n_269),
.B2(n_272),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_284),
.B(n_287),
.C(n_295),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_286),
.A2(n_294),
.B1(n_3),
.B2(n_5),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_279),
.B(n_1),
.C(n_2),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_289),
.B(n_283),
.Y(n_298)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_291),
.Y(n_301)
);

OR2x2_ASAP7_75t_L g300 ( 
.A(n_292),
.B(n_2),
.Y(n_300)
);

XOR2xp5_ASAP7_75t_L g304 ( 
.A(n_293),
.B(n_287),
.Y(n_304)
);

OAI21xp5_ASAP7_75t_SL g295 ( 
.A1(n_270),
.A2(n_2),
.B(n_3),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_273),
.B(n_274),
.Y(n_296)
);

OAI21xp5_ASAP7_75t_L g302 ( 
.A1(n_296),
.A2(n_16),
.B(n_5),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_298),
.B(n_299),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_288),
.A2(n_276),
.B1(n_3),
.B2(n_4),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_300),
.B(n_303),
.Y(n_311)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_302),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_293),
.B(n_3),
.Y(n_303)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_304),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_305),
.B(n_306),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_290),
.B(n_6),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_284),
.B(n_6),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_307),
.B(n_7),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_SL g309 ( 
.A1(n_297),
.A2(n_285),
.B1(n_295),
.B2(n_9),
.Y(n_309)
);

XOR2xp5_ASAP7_75t_L g319 ( 
.A(n_309),
.B(n_7),
.Y(n_319)
);

AOI21xp5_ASAP7_75t_L g317 ( 
.A1(n_313),
.A2(n_300),
.B(n_8),
.Y(n_317)
);

INVx1_ASAP7_75t_SL g314 ( 
.A(n_307),
.Y(n_314)
);

OAI21xp5_ASAP7_75t_L g316 ( 
.A1(n_314),
.A2(n_301),
.B(n_306),
.Y(n_316)
);

XOR2xp5_ASAP7_75t_L g321 ( 
.A(n_316),
.B(n_318),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_317),
.B(n_319),
.Y(n_320)
);

OAI21xp5_ASAP7_75t_L g318 ( 
.A1(n_315),
.A2(n_7),
.B(n_8),
.Y(n_318)
);

AND2x2_ASAP7_75t_L g322 ( 
.A(n_321),
.B(n_312),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_322),
.B(n_308),
.C(n_311),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_323),
.B(n_320),
.C(n_310),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_324),
.B(n_310),
.Y(n_325)
);

MAJx2_ASAP7_75t_L g326 ( 
.A(n_325),
.B(n_8),
.C(n_9),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_326),
.B(n_9),
.C(n_10),
.Y(n_327)
);

AOI22xp5_ASAP7_75t_L g328 ( 
.A1(n_327),
.A2(n_9),
.B1(n_10),
.B2(n_310),
.Y(n_328)
);


endmodule