module fake_jpeg_8555_n_48 (n_3, n_2, n_1, n_0, n_4, n_5, n_48);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_48;

wire n_13;
wire n_21;
wire n_33;
wire n_45;
wire n_23;
wire n_10;
wire n_27;
wire n_6;
wire n_22;
wire n_47;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_31;
wire n_25;
wire n_29;
wire n_37;
wire n_43;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

CKINVDCx20_ASAP7_75t_R g6 ( 
.A(n_0),
.Y(n_6)
);

BUFx6f_ASAP7_75t_L g7 ( 
.A(n_3),
.Y(n_7)
);

INVx4_ASAP7_75t_L g8 ( 
.A(n_5),
.Y(n_8)
);

NOR2xp33_ASAP7_75t_L g9 ( 
.A(n_2),
.B(n_1),
.Y(n_9)
);

INVx1_ASAP7_75t_L g10 ( 
.A(n_1),
.Y(n_10)
);

INVx2_ASAP7_75t_L g11 ( 
.A(n_2),
.Y(n_11)
);

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_0),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_1),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_SL g14 ( 
.A(n_3),
.B(n_2),
.Y(n_14)
);

AND2x4_ASAP7_75t_SL g15 ( 
.A(n_11),
.B(n_0),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_15),
.B(n_16),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_SL g16 ( 
.A(n_14),
.B(n_3),
.Y(n_16)
);

AOI22xp33_ASAP7_75t_L g17 ( 
.A1(n_11),
.A2(n_4),
.B1(n_5),
.B2(n_8),
.Y(n_17)
);

OAI22xp5_ASAP7_75t_L g27 ( 
.A1(n_17),
.A2(n_18),
.B1(n_23),
.B2(n_7),
.Y(n_27)
);

AOI22xp33_ASAP7_75t_SL g18 ( 
.A1(n_8),
.A2(n_4),
.B1(n_5),
.B2(n_10),
.Y(n_18)
);

INVx13_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_19),
.Y(n_24)
);

OAI22xp33_ASAP7_75t_SL g20 ( 
.A1(n_6),
.A2(n_4),
.B1(n_7),
.B2(n_10),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g28 ( 
.A1(n_20),
.A2(n_12),
.B1(n_13),
.B2(n_15),
.Y(n_28)
);

OR2x2_ASAP7_75t_SL g21 ( 
.A(n_14),
.B(n_7),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_21),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_9),
.B(n_6),
.Y(n_22)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_22),
.Y(n_25)
);

AOI22xp5_ASAP7_75t_SL g23 ( 
.A1(n_7),
.A2(n_13),
.B1(n_12),
.B2(n_9),
.Y(n_23)
);

AOI22xp33_ASAP7_75t_SL g31 ( 
.A1(n_27),
.A2(n_15),
.B1(n_21),
.B2(n_19),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_L g30 ( 
.A1(n_28),
.A2(n_17),
.B1(n_23),
.B2(n_15),
.Y(n_30)
);

XOR2xp5_ASAP7_75t_L g36 ( 
.A(n_30),
.B(n_32),
.Y(n_36)
);

CKINVDCx14_ASAP7_75t_R g35 ( 
.A(n_31),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_L g32 ( 
.A1(n_29),
.A2(n_15),
.B1(n_21),
.B2(n_19),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_28),
.Y(n_33)
);

MAJIxp5_ASAP7_75t_L g37 ( 
.A(n_33),
.B(n_29),
.C(n_24),
.Y(n_37)
);

XNOR2xp5_ASAP7_75t_SL g34 ( 
.A(n_32),
.B(n_26),
.Y(n_34)
);

MAJIxp5_ASAP7_75t_L g38 ( 
.A(n_34),
.B(n_37),
.C(n_26),
.Y(n_38)
);

XNOR2xp5_ASAP7_75t_L g42 ( 
.A(n_38),
.B(n_39),
.Y(n_42)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_36),
.Y(n_39)
);

OAI221xp5_ASAP7_75t_L g40 ( 
.A1(n_35),
.A2(n_33),
.B1(n_30),
.B2(n_25),
.C(n_24),
.Y(n_40)
);

XNOR2xp5_ASAP7_75t_L g44 ( 
.A(n_40),
.B(n_20),
.Y(n_44)
);

XOR2xp5_ASAP7_75t_L g41 ( 
.A(n_35),
.B(n_16),
.Y(n_41)
);

MAJIxp5_ASAP7_75t_L g43 ( 
.A(n_41),
.B(n_25),
.C(n_22),
.Y(n_43)
);

OAI211xp5_ASAP7_75t_L g46 ( 
.A1(n_43),
.A2(n_41),
.B(n_12),
.C(n_13),
.Y(n_46)
);

CKINVDCx14_ASAP7_75t_R g45 ( 
.A(n_44),
.Y(n_45)
);

AOI21xp5_ASAP7_75t_L g47 ( 
.A1(n_46),
.A2(n_43),
.B(n_42),
.Y(n_47)
);

XOR2xp5_ASAP7_75t_L g48 ( 
.A(n_47),
.B(n_45),
.Y(n_48)
);


endmodule