module real_aes_18116_n_103 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_103);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_103;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_800;
wire n_618;
wire n_778;
wire n_522;
wire n_838;
wire n_485;
wire n_822;
wire n_846;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_841;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_555;
wire n_421;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_815;
wire n_564;
wire n_519;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_816;
wire n_292;
wire n_539;
wire n_400;
wire n_626;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_559;
wire n_466;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_840;
wire n_570;
wire n_675;
wire n_530;
wire n_835;
wire n_104;
wire n_535;
wire n_732;
wire n_834;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_781;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_812;
wire n_817;
wire n_443;
wire n_565;
wire n_782;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_417;
wire n_449;
wire n_363;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_505;
wire n_527;
wire n_434;
wire n_502;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_552;
wire n_402;
wire n_617;
wire n_733;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_807;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_832;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_848;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_756;
wire n_735;
wire n_728;
wire n_713;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_785;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_845;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_847;
wire n_779;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_765;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_831;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_789;
wire n_268;
wire n_544;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_839;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_836;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_837;
wire n_474;
wire n_829;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_729;
wire n_687;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_802;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_842;
wire n_259;
wire n_143;
wire n_849;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
AND2x4_ASAP7_75t_L g845 ( .A(n_0), .B(n_846), .Y(n_845) );
AOI22xp5_ASAP7_75t_L g497 ( .A1(n_1), .A2(n_3), .B1(n_171), .B2(n_498), .Y(n_497) );
OAI22x1_ASAP7_75t_R g107 ( .A1(n_2), .A2(n_44), .B1(n_108), .B2(n_109), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_2), .Y(n_108) );
AOI22xp33_ASAP7_75t_L g150 ( .A1(n_4), .A2(n_42), .B1(n_128), .B2(n_151), .Y(n_150) );
AOI22xp33_ASAP7_75t_L g472 ( .A1(n_5), .A2(n_25), .B1(n_151), .B2(n_227), .Y(n_472) );
AOI22xp5_ASAP7_75t_L g205 ( .A1(n_6), .A2(n_16), .B1(n_170), .B2(n_206), .Y(n_205) );
AOI22xp33_ASAP7_75t_L g508 ( .A1(n_7), .A2(n_61), .B1(n_188), .B2(n_229), .Y(n_508) );
AOI22xp5_ASAP7_75t_L g514 ( .A1(n_8), .A2(n_17), .B1(n_127), .B2(n_128), .Y(n_514) );
INVx1_ASAP7_75t_L g846 ( .A(n_9), .Y(n_846) );
CKINVDCx5p33_ASAP7_75t_R g568 ( .A(n_10), .Y(n_568) );
CKINVDCx5p33_ASAP7_75t_R g126 ( .A(n_11), .Y(n_126) );
AOI22xp5_ASAP7_75t_L g186 ( .A1(n_12), .A2(n_18), .B1(n_187), .B2(n_190), .Y(n_186) );
OR2x2_ASAP7_75t_L g799 ( .A(n_13), .B(n_39), .Y(n_799) );
BUFx2_ASAP7_75t_L g840 ( .A(n_13), .Y(n_840) );
BUFx6f_ASAP7_75t_L g129 ( .A(n_14), .Y(n_129) );
CKINVDCx5p33_ASAP7_75t_R g210 ( .A(n_15), .Y(n_210) );
INVx2_ASAP7_75t_L g816 ( .A(n_19), .Y(n_816) );
AOI22xp5_ASAP7_75t_L g169 ( .A1(n_20), .A2(n_101), .B1(n_170), .B2(n_171), .Y(n_169) );
AOI22xp33_ASAP7_75t_L g202 ( .A1(n_21), .A2(n_38), .B1(n_136), .B2(n_203), .Y(n_202) );
NAND2xp5_ASAP7_75t_SL g130 ( .A(n_22), .B(n_131), .Y(n_130) );
OAI21x1_ASAP7_75t_L g122 ( .A1(n_23), .A2(n_57), .B(n_123), .Y(n_122) );
CKINVDCx5p33_ASAP7_75t_R g477 ( .A(n_24), .Y(n_477) );
CKINVDCx5p33_ASAP7_75t_R g180 ( .A(n_26), .Y(n_180) );
NAND2xp5_ASAP7_75t_L g484 ( .A(n_27), .B(n_133), .Y(n_484) );
INVx4_ASAP7_75t_R g526 ( .A(n_28), .Y(n_526) );
AOI22xp33_ASAP7_75t_L g155 ( .A1(n_29), .A2(n_47), .B1(n_156), .B2(n_157), .Y(n_155) );
AOI22xp33_ASAP7_75t_L g265 ( .A1(n_30), .A2(n_54), .B1(n_157), .B2(n_170), .Y(n_265) );
CKINVDCx5p33_ASAP7_75t_R g233 ( .A(n_31), .Y(n_233) );
NAND2xp5_ASAP7_75t_L g135 ( .A(n_32), .B(n_136), .Y(n_135) );
CKINVDCx5p33_ASAP7_75t_R g219 ( .A(n_33), .Y(n_219) );
NAND2xp5_ASAP7_75t_SL g491 ( .A(n_34), .B(n_151), .Y(n_491) );
INVx1_ASAP7_75t_L g500 ( .A(n_35), .Y(n_500) );
A2O1A1Ixp33_ASAP7_75t_SL g566 ( .A1(n_36), .A2(n_128), .B(n_132), .C(n_567), .Y(n_566) );
AOI22xp33_ASAP7_75t_L g473 ( .A1(n_37), .A2(n_55), .B1(n_128), .B2(n_157), .Y(n_473) );
HB1xp67_ASAP7_75t_L g839 ( .A(n_39), .Y(n_839) );
AOI22xp5_ASAP7_75t_L g225 ( .A1(n_40), .A2(n_88), .B1(n_128), .B2(n_226), .Y(n_225) );
AOI22xp33_ASAP7_75t_L g191 ( .A1(n_41), .A2(n_46), .B1(n_127), .B2(n_128), .Y(n_191) );
CKINVDCx5p33_ASAP7_75t_R g564 ( .A(n_43), .Y(n_564) );
CKINVDCx5p33_ASAP7_75t_R g109 ( .A(n_44), .Y(n_109) );
AOI22xp33_ASAP7_75t_L g173 ( .A1(n_45), .A2(n_60), .B1(n_170), .B2(n_174), .Y(n_173) );
INVx1_ASAP7_75t_L g488 ( .A(n_48), .Y(n_488) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_49), .B(n_128), .Y(n_490) );
CKINVDCx5p33_ASAP7_75t_R g547 ( .A(n_50), .Y(n_547) );
INVx2_ASAP7_75t_L g794 ( .A(n_51), .Y(n_794) );
CKINVDCx5p33_ASAP7_75t_R g825 ( .A(n_52), .Y(n_825) );
BUFx3_ASAP7_75t_L g797 ( .A(n_53), .Y(n_797) );
INVx1_ASAP7_75t_L g812 ( .A(n_53), .Y(n_812) );
AOI22xp33_ASAP7_75t_L g515 ( .A1(n_56), .A2(n_89), .B1(n_128), .B2(n_157), .Y(n_515) );
CKINVDCx5p33_ASAP7_75t_R g527 ( .A(n_58), .Y(n_527) );
OAI22xp5_ASAP7_75t_L g105 ( .A1(n_59), .A2(n_106), .B1(n_788), .B2(n_789), .Y(n_105) );
INVx1_ASAP7_75t_L g788 ( .A(n_59), .Y(n_788) );
AOI22xp33_ASAP7_75t_L g264 ( .A1(n_62), .A2(n_76), .B1(n_156), .B2(n_174), .Y(n_264) );
CKINVDCx5p33_ASAP7_75t_R g517 ( .A(n_63), .Y(n_517) );
AOI22xp33_ASAP7_75t_L g217 ( .A1(n_64), .A2(n_79), .B1(n_127), .B2(n_128), .Y(n_217) );
AOI22xp5_ASAP7_75t_L g216 ( .A1(n_65), .A2(n_99), .B1(n_170), .B2(n_190), .Y(n_216) );
INVx1_ASAP7_75t_L g123 ( .A(n_66), .Y(n_123) );
AND2x4_ASAP7_75t_L g142 ( .A(n_67), .B(n_143), .Y(n_142) );
AOI22xp5_ASAP7_75t_L g814 ( .A1(n_68), .A2(n_815), .B1(n_816), .B2(n_817), .Y(n_814) );
CKINVDCx5p33_ASAP7_75t_R g817 ( .A(n_68), .Y(n_817) );
AOI22xp33_ASAP7_75t_L g496 ( .A1(n_69), .A2(n_92), .B1(n_156), .B2(n_157), .Y(n_496) );
AO22x1_ASAP7_75t_L g505 ( .A1(n_70), .A2(n_77), .B1(n_203), .B2(n_506), .Y(n_505) );
INVx1_ASAP7_75t_L g143 ( .A(n_71), .Y(n_143) );
AND2x2_ASAP7_75t_L g569 ( .A(n_72), .B(n_145), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_73), .B(n_229), .Y(n_553) );
CKINVDCx5p33_ASAP7_75t_R g562 ( .A(n_74), .Y(n_562) );
AOI22xp5_ASAP7_75t_L g103 ( .A1(n_75), .A2(n_104), .B1(n_834), .B2(n_847), .Y(n_103) );
CKINVDCx16_ASAP7_75t_R g818 ( .A(n_78), .Y(n_818) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_80), .B(n_151), .Y(n_548) );
INVx2_ASAP7_75t_L g133 ( .A(n_81), .Y(n_133) );
NAND2xp5_ASAP7_75t_L g481 ( .A(n_82), .B(n_145), .Y(n_481) );
CKINVDCx5p33_ASAP7_75t_R g523 ( .A(n_83), .Y(n_523) );
AOI22xp33_ASAP7_75t_L g228 ( .A1(n_84), .A2(n_100), .B1(n_157), .B2(n_229), .Y(n_228) );
CKINVDCx5p33_ASAP7_75t_R g267 ( .A(n_85), .Y(n_267) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_86), .B(n_178), .Y(n_509) );
CKINVDCx5p33_ASAP7_75t_R g160 ( .A(n_87), .Y(n_160) );
AOI21xp5_ASAP7_75t_L g826 ( .A1(n_90), .A2(n_823), .B(n_827), .Y(n_826) );
NAND2xp5_ASAP7_75t_SL g144 ( .A(n_91), .B(n_145), .Y(n_144) );
CKINVDCx5p33_ASAP7_75t_R g197 ( .A(n_93), .Y(n_197) );
NAND2xp5_ASAP7_75t_SL g544 ( .A(n_94), .B(n_145), .Y(n_544) );
INVx1_ASAP7_75t_L g460 ( .A(n_95), .Y(n_460) );
NOR2xp33_ASAP7_75t_L g810 ( .A(n_95), .B(n_811), .Y(n_810) );
NAND2xp33_ASAP7_75t_L g138 ( .A(n_96), .B(n_131), .Y(n_138) );
A2O1A1Ixp33_ASAP7_75t_L g521 ( .A1(n_97), .A2(n_193), .B(n_229), .C(n_522), .Y(n_521) );
AND2x2_ASAP7_75t_L g528 ( .A(n_98), .B(n_529), .Y(n_528) );
NAND2xp33_ASAP7_75t_L g552 ( .A(n_102), .B(n_137), .Y(n_552) );
AO21x2_ASAP7_75t_L g104 ( .A1(n_105), .A2(n_790), .B(n_800), .Y(n_104) );
INVx2_ASAP7_75t_L g789 ( .A(n_106), .Y(n_789) );
XNOR2x1_ASAP7_75t_L g106 ( .A(n_107), .B(n_110), .Y(n_106) );
AOI22x1_ASAP7_75t_L g110 ( .A1(n_111), .A2(n_457), .B1(n_461), .B2(n_785), .Y(n_110) );
XNOR2x1_ASAP7_75t_SL g813 ( .A(n_111), .B(n_814), .Y(n_813) );
NAND2x1p5_ASAP7_75t_L g111 ( .A(n_112), .B(n_401), .Y(n_111) );
NOR3x1_ASAP7_75t_L g112 ( .A(n_113), .B(n_319), .C(n_356), .Y(n_112) );
NAND4xp75_ASAP7_75t_L g113 ( .A(n_114), .B(n_239), .C(n_273), .D(n_303), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
OAI32xp33_ASAP7_75t_L g115 ( .A1(n_116), .A2(n_161), .A3(n_211), .B1(n_220), .B2(n_234), .Y(n_115) );
OR2x2_ASAP7_75t_L g220 ( .A(n_116), .B(n_221), .Y(n_220) );
INVx1_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
OAI21xp5_ASAP7_75t_L g430 ( .A1(n_117), .A2(n_431), .B(n_433), .Y(n_430) );
AND2x2_ASAP7_75t_L g117 ( .A(n_118), .B(n_146), .Y(n_117) );
NAND2xp5_ASAP7_75t_L g271 ( .A(n_118), .B(n_272), .Y(n_271) );
AND2x4_ASAP7_75t_L g302 ( .A(n_118), .B(n_248), .Y(n_302) );
AND2x2_ASAP7_75t_L g397 ( .A(n_118), .B(n_213), .Y(n_397) );
INVx2_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
BUFx2_ASAP7_75t_L g246 ( .A(n_119), .Y(n_246) );
OAI21x1_ASAP7_75t_L g119 ( .A1(n_120), .A2(n_124), .B(n_144), .Y(n_119) );
OAI21x1_ASAP7_75t_L g279 ( .A1(n_120), .A2(n_124), .B(n_144), .Y(n_279) );
INVx2_ASAP7_75t_SL g120 ( .A(n_121), .Y(n_120) );
INVx4_ASAP7_75t_L g145 ( .A(n_121), .Y(n_145) );
NOR2xp33_ASAP7_75t_L g159 ( .A(n_121), .B(n_160), .Y(n_159) );
BUFx3_ASAP7_75t_L g208 ( .A(n_121), .Y(n_208) );
NOR2xp33_ASAP7_75t_L g209 ( .A(n_121), .B(n_210), .Y(n_209) );
NOR2xp33_ASAP7_75t_L g218 ( .A(n_121), .B(n_219), .Y(n_218) );
AND2x2_ASAP7_75t_L g492 ( .A(n_121), .B(n_475), .Y(n_492) );
BUFx6f_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
INVx2_ASAP7_75t_L g178 ( .A(n_122), .Y(n_178) );
OAI21x1_ASAP7_75t_L g124 ( .A1(n_125), .A2(n_134), .B(n_140), .Y(n_124) );
O2A1O1Ixp5_ASAP7_75t_L g125 ( .A1(n_126), .A2(n_127), .B(n_130), .C(n_132), .Y(n_125) );
O2A1O1Ixp33_ASAP7_75t_L g546 ( .A1(n_127), .A2(n_547), .B(n_548), .C(n_549), .Y(n_546) );
INVx4_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
INVx1_ASAP7_75t_L g174 ( .A(n_128), .Y(n_174) );
INVx1_ASAP7_75t_L g190 ( .A(n_128), .Y(n_190) );
INVx3_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
BUFx6f_ASAP7_75t_L g131 ( .A(n_129), .Y(n_131) );
BUFx6f_ASAP7_75t_L g137 ( .A(n_129), .Y(n_137) );
BUFx6f_ASAP7_75t_L g151 ( .A(n_129), .Y(n_151) );
BUFx6f_ASAP7_75t_L g157 ( .A(n_129), .Y(n_157) );
INVx1_ASAP7_75t_L g172 ( .A(n_129), .Y(n_172) );
INVx1_ASAP7_75t_L g189 ( .A(n_129), .Y(n_189) );
INVx1_ASAP7_75t_L g204 ( .A(n_129), .Y(n_204) );
INVx1_ASAP7_75t_L g207 ( .A(n_129), .Y(n_207) );
INVx2_ASAP7_75t_L g227 ( .A(n_129), .Y(n_227) );
INVx1_ASAP7_75t_L g229 ( .A(n_129), .Y(n_229) );
INVx3_ASAP7_75t_L g170 ( .A(n_131), .Y(n_170) );
INVxp67_ASAP7_75t_SL g506 ( .A(n_131), .Y(n_506) );
INVx6_ASAP7_75t_L g139 ( .A(n_132), .Y(n_139) );
A2O1A1Ixp33_ASAP7_75t_L g504 ( .A1(n_132), .A2(n_505), .B(n_507), .C(n_510), .Y(n_504) );
AOI21xp5_ASAP7_75t_L g551 ( .A1(n_132), .A2(n_552), .B(n_553), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g578 ( .A(n_132), .B(n_505), .Y(n_578) );
BUFx8_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
INVx2_ASAP7_75t_L g154 ( .A(n_133), .Y(n_154) );
INVx1_ASAP7_75t_L g193 ( .A(n_133), .Y(n_193) );
INVx1_ASAP7_75t_L g487 ( .A(n_133), .Y(n_487) );
AOI21xp5_ASAP7_75t_L g134 ( .A1(n_135), .A2(n_138), .B(n_139), .Y(n_134) );
INVx1_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
INVx2_ASAP7_75t_L g156 ( .A(n_137), .Y(n_156) );
OAI22xp33_ASAP7_75t_L g525 ( .A1(n_137), .A2(n_207), .B1(n_526), .B2(n_527), .Y(n_525) );
OAI22xp5_ASAP7_75t_L g149 ( .A1(n_139), .A2(n_150), .B1(n_152), .B2(n_155), .Y(n_149) );
OAI22xp5_ASAP7_75t_L g168 ( .A1(n_139), .A2(n_152), .B1(n_169), .B2(n_173), .Y(n_168) );
OAI22xp5_ASAP7_75t_L g185 ( .A1(n_139), .A2(n_186), .B1(n_191), .B2(n_192), .Y(n_185) );
OAI22xp5_ASAP7_75t_L g201 ( .A1(n_139), .A2(n_152), .B1(n_202), .B2(n_205), .Y(n_201) );
OAI22xp5_ASAP7_75t_L g215 ( .A1(n_139), .A2(n_192), .B1(n_216), .B2(n_217), .Y(n_215) );
OAI22xp5_ASAP7_75t_L g224 ( .A1(n_139), .A2(n_225), .B1(n_228), .B2(n_230), .Y(n_224) );
OAI22xp5_ASAP7_75t_L g263 ( .A1(n_139), .A2(n_152), .B1(n_264), .B2(n_265), .Y(n_263) );
OAI22xp5_ASAP7_75t_L g471 ( .A1(n_139), .A2(n_472), .B1(n_473), .B2(n_474), .Y(n_471) );
OAI22xp5_ASAP7_75t_L g495 ( .A1(n_139), .A2(n_230), .B1(n_496), .B2(n_497), .Y(n_495) );
OAI22x1_ASAP7_75t_L g513 ( .A1(n_139), .A2(n_230), .B1(n_514), .B2(n_515), .Y(n_513) );
INVx2_ASAP7_75t_SL g140 ( .A(n_141), .Y(n_140) );
INVx2_ASAP7_75t_SL g231 ( .A(n_141), .Y(n_231) );
INVx1_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
BUFx10_ASAP7_75t_L g148 ( .A(n_142), .Y(n_148) );
BUFx10_ASAP7_75t_L g475 ( .A(n_142), .Y(n_475) );
INVx1_ASAP7_75t_L g511 ( .A(n_142), .Y(n_511) );
INVx2_ASAP7_75t_L g158 ( .A(n_145), .Y(n_158) );
NOR2x1_ASAP7_75t_L g554 ( .A(n_145), .B(n_555), .Y(n_554) );
INVx2_ASAP7_75t_L g270 ( .A(n_146), .Y(n_270) );
NAND2xp5_ASAP7_75t_L g278 ( .A(n_146), .B(n_279), .Y(n_278) );
INVx2_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
HB1xp67_ASAP7_75t_L g257 ( .A(n_147), .Y(n_257) );
INVx1_ASAP7_75t_L g301 ( .A(n_147), .Y(n_301) );
AND2x2_ASAP7_75t_L g345 ( .A(n_147), .B(n_279), .Y(n_345) );
OR2x2_ASAP7_75t_L g399 ( .A(n_147), .B(n_223), .Y(n_399) );
AO31x2_ASAP7_75t_L g147 ( .A1(n_148), .A2(n_149), .A3(n_158), .B(n_159), .Y(n_147) );
INVx2_ASAP7_75t_L g167 ( .A(n_148), .Y(n_167) );
AO31x2_ASAP7_75t_L g184 ( .A1(n_148), .A2(n_185), .A3(n_194), .B(n_196), .Y(n_184) );
AO31x2_ASAP7_75t_L g200 ( .A1(n_148), .A2(n_201), .A3(n_208), .B(n_209), .Y(n_200) );
AO31x2_ASAP7_75t_L g512 ( .A1(n_148), .A2(n_181), .A3(n_513), .B(n_516), .Y(n_512) );
NOR2xp33_ASAP7_75t_L g561 ( .A(n_151), .B(n_562), .Y(n_561) );
INVx2_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
INVx2_ASAP7_75t_L g474 ( .A(n_153), .Y(n_474) );
BUFx3_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
INVx2_ASAP7_75t_L g550 ( .A(n_154), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g485 ( .A(n_157), .B(n_486), .Y(n_485) );
INVx2_ASAP7_75t_L g498 ( .A(n_157), .Y(n_498) );
AO31x2_ASAP7_75t_L g470 ( .A1(n_158), .A2(n_471), .A3(n_475), .B(n_476), .Y(n_470) );
INVx1_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
AOI22xp33_ASAP7_75t_L g416 ( .A1(n_162), .A2(n_325), .B1(n_417), .B2(n_419), .Y(n_416) );
AND2x2_ASAP7_75t_L g162 ( .A(n_163), .B(n_182), .Y(n_162) );
INVx4_ASAP7_75t_L g242 ( .A(n_163), .Y(n_242) );
AOI22xp5_ASAP7_75t_L g253 ( .A1(n_163), .A2(n_222), .B1(n_254), .B2(n_256), .Y(n_253) );
OR2x2_ASAP7_75t_L g259 ( .A(n_163), .B(n_260), .Y(n_259) );
AND2x2_ASAP7_75t_L g378 ( .A(n_163), .B(n_277), .Y(n_378) );
INVx3_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
AND2x2_ASAP7_75t_L g298 ( .A(n_164), .B(n_183), .Y(n_298) );
AND2x2_ASAP7_75t_L g389 ( .A(n_164), .B(n_261), .Y(n_389) );
AND2x2_ASAP7_75t_L g444 ( .A(n_164), .B(n_200), .Y(n_444) );
INVx2_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
INVx2_ASAP7_75t_L g238 ( .A(n_165), .Y(n_238) );
AND2x4_ASAP7_75t_L g365 ( .A(n_165), .B(n_261), .Y(n_365) );
AO31x2_ASAP7_75t_L g165 ( .A1(n_166), .A2(n_168), .A3(n_175), .B(n_179), .Y(n_165) );
AO31x2_ASAP7_75t_L g214 ( .A1(n_166), .A2(n_194), .A3(n_215), .B(n_218), .Y(n_214) );
INVx1_ASAP7_75t_L g166 ( .A(n_167), .Y(n_166) );
AOI21xp5_ASAP7_75t_L g520 ( .A1(n_167), .A2(n_521), .B(n_524), .Y(n_520) );
INVx2_ASAP7_75t_L g171 ( .A(n_172), .Y(n_171) );
NOR2xp33_ASAP7_75t_L g563 ( .A(n_172), .B(n_564), .Y(n_563) );
AO31x2_ASAP7_75t_L g262 ( .A1(n_175), .A2(n_231), .A3(n_263), .B(n_266), .Y(n_262) );
AO21x2_ASAP7_75t_L g519 ( .A1(n_175), .A2(n_520), .B(n_528), .Y(n_519) );
INVx2_ASAP7_75t_L g175 ( .A(n_176), .Y(n_175) );
INVx2_ASAP7_75t_L g176 ( .A(n_177), .Y(n_176) );
NOR2xp33_ASAP7_75t_SL g196 ( .A(n_177), .B(n_197), .Y(n_196) );
NOR2xp33_ASAP7_75t_L g232 ( .A(n_177), .B(n_233), .Y(n_232) );
INVx2_ASAP7_75t_L g177 ( .A(n_178), .Y(n_177) );
INVx2_ASAP7_75t_L g181 ( .A(n_178), .Y(n_181) );
INVx2_ASAP7_75t_L g195 ( .A(n_178), .Y(n_195) );
OAI21xp33_ASAP7_75t_L g510 ( .A1(n_178), .A2(n_509), .B(n_511), .Y(n_510) );
NOR2xp33_ASAP7_75t_L g179 ( .A(n_180), .B(n_181), .Y(n_179) );
NOR2xp33_ASAP7_75t_L g266 ( .A(n_181), .B(n_267), .Y(n_266) );
NAND2x1_ASAP7_75t_L g241 ( .A(n_182), .B(n_242), .Y(n_241) );
NAND2xp5_ASAP7_75t_SL g348 ( .A(n_182), .B(n_349), .Y(n_348) );
AND2x4_ASAP7_75t_L g182 ( .A(n_183), .B(n_198), .Y(n_182) );
INVx2_ASAP7_75t_L g236 ( .A(n_183), .Y(n_236) );
NAND2xp5_ASAP7_75t_L g260 ( .A(n_183), .B(n_261), .Y(n_260) );
INVx1_ASAP7_75t_L g284 ( .A(n_183), .Y(n_284) );
NAND2xp5_ASAP7_75t_L g311 ( .A(n_183), .B(n_286), .Y(n_311) );
AND2x2_ASAP7_75t_L g314 ( .A(n_183), .B(n_315), .Y(n_314) );
INVx1_ASAP7_75t_L g374 ( .A(n_183), .Y(n_374) );
INVx4_ASAP7_75t_SL g183 ( .A(n_184), .Y(n_183) );
NAND2xp5_ASAP7_75t_L g252 ( .A(n_184), .B(n_199), .Y(n_252) );
BUFx2_ASAP7_75t_L g290 ( .A(n_184), .Y(n_290) );
AND2x2_ASAP7_75t_L g339 ( .A(n_184), .B(n_200), .Y(n_339) );
AND2x2_ASAP7_75t_L g381 ( .A(n_184), .B(n_262), .Y(n_381) );
NAND2xp5_ASAP7_75t_L g413 ( .A(n_184), .B(n_414), .Y(n_413) );
INVx1_ASAP7_75t_L g187 ( .A(n_188), .Y(n_187) );
INVx2_ASAP7_75t_L g188 ( .A(n_189), .Y(n_188) );
NOR2xp33_ASAP7_75t_L g522 ( .A(n_189), .B(n_523), .Y(n_522) );
INVx1_ASAP7_75t_SL g192 ( .A(n_193), .Y(n_192) );
INVx1_ASAP7_75t_L g230 ( .A(n_193), .Y(n_230) );
AO31x2_ASAP7_75t_L g494 ( .A1(n_194), .A2(n_231), .A3(n_495), .B(n_499), .Y(n_494) );
AOI21x1_ASAP7_75t_L g558 ( .A1(n_194), .A2(n_559), .B(n_569), .Y(n_558) );
BUFx2_ASAP7_75t_L g194 ( .A(n_195), .Y(n_194) );
NOR2xp33_ASAP7_75t_L g476 ( .A(n_195), .B(n_477), .Y(n_476) );
NOR2xp33_ASAP7_75t_L g499 ( .A(n_195), .B(n_500), .Y(n_499) );
NOR2xp33_ASAP7_75t_L g516 ( .A(n_195), .B(n_517), .Y(n_516) );
INVx2_ASAP7_75t_L g529 ( .A(n_195), .Y(n_529) );
INVx1_ASAP7_75t_L g198 ( .A(n_199), .Y(n_198) );
INVx1_ASAP7_75t_L g199 ( .A(n_200), .Y(n_199) );
NAND2xp5_ASAP7_75t_L g285 ( .A(n_200), .B(n_286), .Y(n_285) );
OR2x2_ASAP7_75t_L g292 ( .A(n_200), .B(n_262), .Y(n_292) );
INVx1_ASAP7_75t_L g315 ( .A(n_200), .Y(n_315) );
INVx2_ASAP7_75t_L g335 ( .A(n_200), .Y(n_335) );
HB1xp67_ASAP7_75t_L g380 ( .A(n_200), .Y(n_380) );
OAI21xp33_ASAP7_75t_SL g483 ( .A1(n_203), .A2(n_484), .B(n_485), .Y(n_483) );
INVx1_ASAP7_75t_L g203 ( .A(n_204), .Y(n_203) );
INVx1_ASAP7_75t_L g206 ( .A(n_207), .Y(n_206) );
AO31x2_ASAP7_75t_L g223 ( .A1(n_208), .A2(n_224), .A3(n_231), .B(n_232), .Y(n_223) );
INVx1_ASAP7_75t_L g211 ( .A(n_212), .Y(n_211) );
AND2x2_ASAP7_75t_L g299 ( .A(n_212), .B(n_300), .Y(n_299) );
NOR2x1p5_ASAP7_75t_L g405 ( .A(n_212), .B(n_399), .Y(n_405) );
INVx2_ASAP7_75t_L g212 ( .A(n_213), .Y(n_212) );
AND2x4_ASAP7_75t_L g222 ( .A(n_213), .B(n_223), .Y(n_222) );
INVx3_ASAP7_75t_L g255 ( .A(n_213), .Y(n_255) );
NAND2xp5_ASAP7_75t_L g269 ( .A(n_213), .B(n_270), .Y(n_269) );
NAND2xp5_ASAP7_75t_L g330 ( .A(n_213), .B(n_331), .Y(n_330) );
INVx3_ASAP7_75t_L g213 ( .A(n_214), .Y(n_213) );
AND2x2_ASAP7_75t_L g247 ( .A(n_214), .B(n_248), .Y(n_247) );
AND2x2_ASAP7_75t_L g305 ( .A(n_214), .B(n_223), .Y(n_305) );
BUFx2_ASAP7_75t_L g418 ( .A(n_214), .Y(n_418) );
NAND2xp5_ASAP7_75t_L g243 ( .A(n_220), .B(n_244), .Y(n_243) );
INVx1_ASAP7_75t_L g456 ( .A(n_220), .Y(n_456) );
INVx2_ASAP7_75t_SL g221 ( .A(n_222), .Y(n_221) );
INVx1_ASAP7_75t_L g392 ( .A(n_222), .Y(n_392) );
AND2x4_ASAP7_75t_L g415 ( .A(n_222), .B(n_345), .Y(n_415) );
AND2x2_ASAP7_75t_L g439 ( .A(n_222), .B(n_440), .Y(n_439) );
INVx2_ASAP7_75t_L g248 ( .A(n_223), .Y(n_248) );
BUFx2_ASAP7_75t_L g272 ( .A(n_223), .Y(n_272) );
INVx1_ASAP7_75t_L g328 ( .A(n_223), .Y(n_328) );
OR2x2_ASAP7_75t_L g450 ( .A(n_223), .B(n_307), .Y(n_450) );
INVx2_ASAP7_75t_SL g226 ( .A(n_227), .Y(n_226) );
NOR2xp33_ASAP7_75t_L g567 ( .A(n_227), .B(n_568), .Y(n_567) );
NAND2xp5_ASAP7_75t_SL g524 ( .A(n_230), .B(n_525), .Y(n_524) );
HB1xp67_ASAP7_75t_L g234 ( .A(n_235), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g235 ( .A(n_236), .B(n_237), .Y(n_235) );
INVx2_ASAP7_75t_L g296 ( .A(n_236), .Y(n_296) );
HB1xp67_ASAP7_75t_L g313 ( .A(n_237), .Y(n_313) );
INVx1_ASAP7_75t_L g317 ( .A(n_237), .Y(n_317) );
INVx1_ASAP7_75t_L g237 ( .A(n_238), .Y(n_237) );
INVx2_ASAP7_75t_L g258 ( .A(n_238), .Y(n_258) );
OR2x2_ASAP7_75t_L g295 ( .A(n_238), .B(n_287), .Y(n_295) );
AOI21xp5_ASAP7_75t_L g239 ( .A1(n_240), .A2(n_243), .B(n_249), .Y(n_239) );
INVx2_ASAP7_75t_L g240 ( .A(n_241), .Y(n_240) );
OAI22xp5_ASAP7_75t_L g337 ( .A1(n_244), .A2(n_338), .B1(n_340), .B2(n_343), .Y(n_337) );
INVx1_ASAP7_75t_L g244 ( .A(n_245), .Y(n_244) );
AND2x2_ASAP7_75t_L g245 ( .A(n_246), .B(n_247), .Y(n_245) );
OR2x2_ASAP7_75t_L g383 ( .A(n_246), .B(n_384), .Y(n_383) );
INVx1_ASAP7_75t_L g391 ( .A(n_246), .Y(n_391) );
AND2x2_ASAP7_75t_L g404 ( .A(n_246), .B(n_405), .Y(n_404) );
AND2x2_ASAP7_75t_L g366 ( .A(n_247), .B(n_345), .Y(n_366) );
OAI22xp5_ASAP7_75t_L g249 ( .A1(n_250), .A2(n_253), .B1(n_259), .B2(n_268), .Y(n_249) );
INVx1_ASAP7_75t_L g250 ( .A(n_251), .Y(n_250) );
INVx1_ASAP7_75t_L g251 ( .A(n_252), .Y(n_251) );
INVx1_ASAP7_75t_L g318 ( .A(n_252), .Y(n_318) );
INVx1_ASAP7_75t_L g254 ( .A(n_255), .Y(n_254) );
AND2x4_ASAP7_75t_L g276 ( .A(n_255), .B(n_277), .Y(n_276) );
AND2x2_ASAP7_75t_L g344 ( .A(n_255), .B(n_345), .Y(n_344) );
INVx2_ASAP7_75t_L g353 ( .A(n_255), .Y(n_353) );
NAND2xp5_ASAP7_75t_L g369 ( .A(n_255), .B(n_370), .Y(n_369) );
NAND2xp5_ASAP7_75t_L g424 ( .A(n_256), .B(n_425), .Y(n_424) );
AND2x2_ASAP7_75t_L g256 ( .A(n_257), .B(n_258), .Y(n_256) );
AND2x2_ASAP7_75t_L g341 ( .A(n_258), .B(n_342), .Y(n_341) );
INVx3_ASAP7_75t_L g355 ( .A(n_258), .Y(n_355) );
INVx2_ASAP7_75t_L g261 ( .A(n_262), .Y(n_261) );
INVx2_ASAP7_75t_L g287 ( .A(n_262), .Y(n_287) );
AND2x4_ASAP7_75t_L g334 ( .A(n_262), .B(n_335), .Y(n_334) );
HB1xp67_ASAP7_75t_L g350 ( .A(n_262), .Y(n_350) );
INVx1_ASAP7_75t_L g414 ( .A(n_262), .Y(n_414) );
OR2x2_ASAP7_75t_L g268 ( .A(n_269), .B(n_271), .Y(n_268) );
AND2x4_ASAP7_75t_L g306 ( .A(n_270), .B(n_307), .Y(n_306) );
INVx1_ASAP7_75t_L g323 ( .A(n_270), .Y(n_323) );
INVx1_ASAP7_75t_L g281 ( .A(n_272), .Y(n_281) );
AOI22xp5_ASAP7_75t_L g273 ( .A1(n_274), .A2(n_282), .B1(n_293), .B2(n_299), .Y(n_273) );
INVx1_ASAP7_75t_L g274 ( .A(n_275), .Y(n_274) );
NAND2x1p5_ASAP7_75t_L g275 ( .A(n_276), .B(n_280), .Y(n_275) );
INVx1_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
INVxp67_ASAP7_75t_SL g331 ( .A(n_278), .Y(n_331) );
INVx1_ASAP7_75t_L g307 ( .A(n_279), .Y(n_307) );
INVx1_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
NAND2xp5_ASAP7_75t_SL g282 ( .A(n_283), .B(n_288), .Y(n_282) );
OR2x2_ASAP7_75t_L g283 ( .A(n_284), .B(n_285), .Y(n_283) );
NAND2xp5_ASAP7_75t_L g333 ( .A(n_284), .B(n_334), .Y(n_333) );
INVx1_ASAP7_75t_L g436 ( .A(n_285), .Y(n_436) );
INVx1_ASAP7_75t_L g455 ( .A(n_285), .Y(n_455) );
INVx1_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
INVx1_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
NAND2x1_ASAP7_75t_L g432 ( .A(n_289), .B(n_355), .Y(n_432) );
AND2x4_ASAP7_75t_L g289 ( .A(n_290), .B(n_291), .Y(n_289) );
INVx1_ASAP7_75t_L g448 ( .A(n_290), .Y(n_448) );
INVx2_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
NAND2xp5_ASAP7_75t_L g293 ( .A(n_294), .B(n_297), .Y(n_293) );
INVx2_ASAP7_75t_L g386 ( .A(n_294), .Y(n_386) );
OR2x2_ASAP7_75t_L g294 ( .A(n_295), .B(n_296), .Y(n_294) );
INVx2_ASAP7_75t_L g375 ( .A(n_295), .Y(n_375) );
AND2x4_ASAP7_75t_L g377 ( .A(n_296), .B(n_334), .Y(n_377) );
INVx1_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
AOI22xp5_ASAP7_75t_L g445 ( .A1(n_300), .A2(n_446), .B1(n_449), .B2(n_451), .Y(n_445) );
AND2x4_ASAP7_75t_L g300 ( .A(n_301), .B(n_302), .Y(n_300) );
INVx2_ASAP7_75t_L g370 ( .A(n_301), .Y(n_370) );
INVx1_ASAP7_75t_L g324 ( .A(n_302), .Y(n_324) );
AND2x4_ASAP7_75t_L g417 ( .A(n_302), .B(n_418), .Y(n_417) );
AND2x2_ASAP7_75t_L g425 ( .A(n_302), .B(n_426), .Y(n_425) );
NAND2xp5_ASAP7_75t_L g303 ( .A(n_304), .B(n_308), .Y(n_303) );
AND2x4_ASAP7_75t_SL g304 ( .A(n_305), .B(n_306), .Y(n_304) );
INVx1_ASAP7_75t_SL g368 ( .A(n_305), .Y(n_368) );
INVx2_ASAP7_75t_L g384 ( .A(n_305), .Y(n_384) );
INVx1_ASAP7_75t_L g411 ( .A(n_306), .Y(n_411) );
AND2x2_ASAP7_75t_L g442 ( .A(n_306), .B(n_353), .Y(n_442) );
NAND3xp33_ASAP7_75t_L g308 ( .A(n_309), .B(n_312), .C(n_316), .Y(n_308) );
INVx1_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
INVx1_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
NAND2xp5_ASAP7_75t_L g312 ( .A(n_313), .B(n_314), .Y(n_312) );
NAND2xp5_ASAP7_75t_L g338 ( .A(n_313), .B(n_339), .Y(n_338) );
AND2x2_ASAP7_75t_L g354 ( .A(n_314), .B(n_355), .Y(n_354) );
NAND2xp5_ASAP7_75t_L g422 ( .A(n_314), .B(n_389), .Y(n_422) );
INVx1_ASAP7_75t_L g342 ( .A(n_315), .Y(n_342) );
NAND2xp5_ASAP7_75t_L g316 ( .A(n_317), .B(n_318), .Y(n_316) );
NAND2xp5_ASAP7_75t_L g407 ( .A(n_317), .B(n_381), .Y(n_407) );
INVx1_ASAP7_75t_L g362 ( .A(n_318), .Y(n_362) );
NAND3xp33_ASAP7_75t_L g319 ( .A(n_320), .B(n_336), .C(n_346), .Y(n_319) );
OAI21xp5_ASAP7_75t_L g320 ( .A1(n_321), .A2(n_325), .B(n_332), .Y(n_320) );
INVxp67_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
OR2x2_ASAP7_75t_L g322 ( .A(n_323), .B(n_324), .Y(n_322) );
INVx1_ASAP7_75t_L g440 ( .A(n_323), .Y(n_440) );
AND2x4_ASAP7_75t_L g325 ( .A(n_326), .B(n_329), .Y(n_325) );
INVx1_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
AOI32xp33_ASAP7_75t_L g376 ( .A1(n_327), .A2(n_377), .A3(n_378), .B1(n_379), .B2(n_382), .Y(n_376) );
NOR2xp33_ASAP7_75t_L g410 ( .A(n_327), .B(n_411), .Y(n_410) );
BUFx2_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
INVx1_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
INVx1_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
INVx2_ASAP7_75t_L g360 ( .A(n_334), .Y(n_360) );
NAND2x1p5_ASAP7_75t_L g395 ( .A(n_334), .B(n_355), .Y(n_395) );
INVx1_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
NAND2xp5_ASAP7_75t_L g388 ( .A(n_339), .B(n_389), .Y(n_388) );
AND2x2_ASAP7_75t_L g400 ( .A(n_339), .B(n_349), .Y(n_400) );
INVx1_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
INVx1_ASAP7_75t_L g428 ( .A(n_342), .Y(n_428) );
INVx1_ASAP7_75t_SL g343 ( .A(n_344), .Y(n_343) );
AOI22xp33_ASAP7_75t_SL g346 ( .A1(n_344), .A2(n_347), .B1(n_351), .B2(n_354), .Y(n_346) );
NAND2xp5_ASAP7_75t_L g352 ( .A(n_345), .B(n_353), .Y(n_352) );
AOI22xp5_ASAP7_75t_L g441 ( .A1(n_347), .A2(n_405), .B1(n_442), .B2(n_443), .Y(n_441) );
INVx1_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
AND2x2_ASAP7_75t_L g443 ( .A(n_349), .B(n_444), .Y(n_443) );
INVx1_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
AOI22xp33_ASAP7_75t_L g393 ( .A1(n_351), .A2(n_394), .B1(n_396), .B2(n_400), .Y(n_393) );
INVx2_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
INVx2_ASAP7_75t_L g435 ( .A(n_355), .Y(n_435) );
NAND4xp25_ASAP7_75t_L g356 ( .A(n_357), .B(n_376), .C(n_385), .D(n_393), .Y(n_356) );
O2A1O1Ixp5_ASAP7_75t_L g357 ( .A1(n_358), .A2(n_363), .B(n_366), .C(n_367), .Y(n_357) );
NOR2x1_ASAP7_75t_L g358 ( .A(n_359), .B(n_361), .Y(n_358) );
INVx1_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
INVx1_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
INVx2_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
INVx3_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
AND2x4_ASAP7_75t_L g421 ( .A(n_365), .B(n_380), .Y(n_421) );
NAND2xp5_ASAP7_75t_L g447 ( .A(n_365), .B(n_448), .Y(n_447) );
AOI21xp5_ASAP7_75t_L g367 ( .A1(n_368), .A2(n_369), .B(n_371), .Y(n_367) );
INVx1_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
AOI22xp5_ASAP7_75t_L g409 ( .A1(n_372), .A2(n_410), .B1(n_412), .B2(n_415), .Y(n_409) );
AND2x4_ASAP7_75t_L g372 ( .A(n_373), .B(n_375), .Y(n_372) );
INVx1_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
OAI21xp5_ASAP7_75t_L g438 ( .A1(n_377), .A2(n_382), .B(n_439), .Y(n_438) );
AND2x4_ASAP7_75t_L g379 ( .A(n_380), .B(n_381), .Y(n_379) );
INVx1_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
OAI21xp33_ASAP7_75t_L g385 ( .A1(n_386), .A2(n_387), .B(n_390), .Y(n_385) );
INVx2_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
NOR2xp33_ASAP7_75t_R g390 ( .A(n_391), .B(n_392), .Y(n_390) );
INVx2_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
AND2x2_ASAP7_75t_L g396 ( .A(n_397), .B(n_398), .Y(n_396) );
INVx1_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
AOI22xp5_ASAP7_75t_L g453 ( .A1(n_400), .A2(n_417), .B1(n_454), .B2(n_456), .Y(n_453) );
NOR3x1_ASAP7_75t_L g401 ( .A(n_402), .B(n_423), .C(n_437), .Y(n_401) );
NAND2xp5_ASAP7_75t_L g402 ( .A(n_403), .B(n_416), .Y(n_402) );
AOI21xp33_ASAP7_75t_L g403 ( .A1(n_404), .A2(n_406), .B(n_408), .Y(n_403) );
INVx1_ASAP7_75t_L g429 ( .A(n_404), .Y(n_429) );
INVx2_ASAP7_75t_SL g406 ( .A(n_407), .Y(n_406) );
INVxp67_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
INVx1_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
INVx1_ASAP7_75t_L g452 ( .A(n_414), .Y(n_452) );
INVx1_ASAP7_75t_L g426 ( .A(n_418), .Y(n_426) );
NAND2xp5_ASAP7_75t_L g419 ( .A(n_420), .B(n_422), .Y(n_419) );
OAI221xp5_ASAP7_75t_L g423 ( .A1(n_420), .A2(n_424), .B1(n_427), .B2(n_429), .C(n_430), .Y(n_423) );
INVx1_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
INVx1_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
INVx1_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
INVx2_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
NAND2xp5_ASAP7_75t_L g434 ( .A(n_435), .B(n_436), .Y(n_434) );
NAND4xp25_ASAP7_75t_SL g437 ( .A(n_438), .B(n_441), .C(n_445), .D(n_453), .Y(n_437) );
AND2x2_ASAP7_75t_L g451 ( .A(n_444), .B(n_452), .Y(n_451) );
INVxp67_ASAP7_75t_SL g446 ( .A(n_447), .Y(n_446) );
INVxp67_ASAP7_75t_SL g449 ( .A(n_450), .Y(n_449) );
HB1xp67_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
INVx1_ASAP7_75t_SL g457 ( .A(n_458), .Y(n_457) );
HB1xp67_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
CKINVDCx5p33_ASAP7_75t_R g787 ( .A(n_459), .Y(n_787) );
AND2x2_ASAP7_75t_L g832 ( .A(n_459), .B(n_833), .Y(n_832) );
INVx2_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
BUFx2_ASAP7_75t_L g844 ( .A(n_460), .Y(n_844) );
INVx2_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
AND2x4_ASAP7_75t_L g462 ( .A(n_463), .B(n_662), .Y(n_462) );
NOR2x1_ASAP7_75t_L g463 ( .A(n_464), .B(n_610), .Y(n_463) );
OAI211xp5_ASAP7_75t_L g464 ( .A1(n_465), .A2(n_501), .B(n_530), .C(n_595), .Y(n_464) );
HB1xp67_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
INVx1_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
OAI21xp5_ASAP7_75t_L g745 ( .A1(n_467), .A2(n_531), .B(n_746), .Y(n_745) );
AND2x4_ASAP7_75t_L g467 ( .A(n_468), .B(n_478), .Y(n_467) );
INVx2_ASAP7_75t_L g591 ( .A(n_468), .Y(n_591) );
NOR2xp33_ASAP7_75t_L g765 ( .A(n_468), .B(n_766), .Y(n_765) );
INVx2_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
AND2x2_ASAP7_75t_L g702 ( .A(n_469), .B(n_480), .Y(n_702) );
BUFx2_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
INVx2_ASAP7_75t_SL g570 ( .A(n_470), .Y(n_570) );
NAND2xp5_ASAP7_75t_L g607 ( .A(n_470), .B(n_494), .Y(n_607) );
AND2x2_ASAP7_75t_L g640 ( .A(n_470), .B(n_557), .Y(n_640) );
OR2x2_ASAP7_75t_L g645 ( .A(n_470), .B(n_494), .Y(n_645) );
AOI21xp5_ASAP7_75t_L g489 ( .A1(n_474), .A2(n_490), .B(n_491), .Y(n_489) );
OAI21x1_ASAP7_75t_L g507 ( .A1(n_474), .A2(n_508), .B(n_509), .Y(n_507) );
INVx1_ASAP7_75t_L g555 ( .A(n_475), .Y(n_555) );
INVx1_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
INVx1_ASAP7_75t_L g784 ( .A(n_479), .Y(n_784) );
OR2x2_ASAP7_75t_L g479 ( .A(n_480), .B(n_493), .Y(n_479) );
AND2x2_ASAP7_75t_L g585 ( .A(n_480), .B(n_494), .Y(n_585) );
INVx3_ASAP7_75t_L g593 ( .A(n_480), .Y(n_593) );
NAND2x1p5_ASAP7_75t_SL g625 ( .A(n_480), .B(n_609), .Y(n_625) );
INVx1_ASAP7_75t_L g643 ( .A(n_480), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g668 ( .A(n_480), .B(n_588), .Y(n_668) );
BUFx2_ASAP7_75t_L g754 ( .A(n_480), .Y(n_754) );
AND2x4_ASAP7_75t_L g480 ( .A(n_481), .B(n_482), .Y(n_480) );
OAI21xp5_ASAP7_75t_L g482 ( .A1(n_483), .A2(n_489), .B(n_492), .Y(n_482) );
NOR2xp33_ASAP7_75t_L g486 ( .A(n_487), .B(n_488), .Y(n_486) );
BUFx4f_ASAP7_75t_L g565 ( .A(n_487), .Y(n_565) );
INVx1_ASAP7_75t_L g493 ( .A(n_494), .Y(n_493) );
INVx1_ASAP7_75t_L g538 ( .A(n_494), .Y(n_538) );
INVx1_ASAP7_75t_L g594 ( .A(n_494), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g667 ( .A(n_494), .B(n_570), .Y(n_667) );
NOR2xp33_ASAP7_75t_L g703 ( .A(n_494), .B(n_557), .Y(n_703) );
OR2x2_ASAP7_75t_L g501 ( .A(n_502), .B(n_518), .Y(n_501) );
INVx1_ASAP7_75t_L g761 ( .A(n_502), .Y(n_761) );
NAND2xp5_ASAP7_75t_L g502 ( .A(n_503), .B(n_512), .Y(n_502) );
OR2x2_ASAP7_75t_L g533 ( .A(n_503), .B(n_534), .Y(n_533) );
INVx2_ASAP7_75t_L g598 ( .A(n_503), .Y(n_598) );
INVx1_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
INVx1_ASAP7_75t_L g577 ( .A(n_507), .Y(n_577) );
INVx1_ASAP7_75t_L g579 ( .A(n_510), .Y(n_579) );
AOI21xp5_ASAP7_75t_L g559 ( .A1(n_511), .A2(n_560), .B(n_566), .Y(n_559) );
INVx2_ASAP7_75t_L g534 ( .A(n_512), .Y(n_534) );
OR2x2_ASAP7_75t_L g599 ( .A(n_512), .B(n_519), .Y(n_599) );
AND2x2_ASAP7_75t_L g604 ( .A(n_512), .B(n_519), .Y(n_604) );
INVx2_ASAP7_75t_L g649 ( .A(n_512), .Y(n_649) );
AND2x2_ASAP7_75t_L g690 ( .A(n_512), .B(n_543), .Y(n_690) );
AND2x2_ASAP7_75t_L g724 ( .A(n_512), .B(n_621), .Y(n_724) );
INVx1_ASAP7_75t_L g535 ( .A(n_518), .Y(n_535) );
INVx1_ASAP7_75t_L g654 ( .A(n_518), .Y(n_654) );
INVx1_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
AND2x2_ASAP7_75t_L g574 ( .A(n_519), .B(n_575), .Y(n_574) );
AND2x4_ASAP7_75t_L g615 ( .A(n_519), .B(n_576), .Y(n_615) );
INVx2_ASAP7_75t_L g621 ( .A(n_519), .Y(n_621) );
AND2x2_ASAP7_75t_L g676 ( .A(n_519), .B(n_543), .Y(n_676) );
AND2x2_ASAP7_75t_L g733 ( .A(n_519), .B(n_542), .Y(n_733) );
AOI22xp5_ASAP7_75t_L g530 ( .A1(n_531), .A2(n_536), .B1(n_571), .B2(n_582), .Y(n_530) );
INVx3_ASAP7_75t_L g531 ( .A(n_532), .Y(n_531) );
OR2x2_ASAP7_75t_L g532 ( .A(n_533), .B(n_535), .Y(n_532) );
NAND3xp33_ASAP7_75t_SL g711 ( .A(n_533), .B(n_712), .C(n_714), .Y(n_711) );
INVx1_ASAP7_75t_L g630 ( .A(n_534), .Y(n_630) );
AND2x2_ASAP7_75t_L g680 ( .A(n_534), .B(n_542), .Y(n_680) );
INVx1_ASAP7_75t_L g780 ( .A(n_535), .Y(n_780) );
AND2x2_ASAP7_75t_L g536 ( .A(n_537), .B(n_539), .Y(n_536) );
NOR2xp33_ASAP7_75t_L g771 ( .A(n_537), .B(n_735), .Y(n_771) );
BUFx3_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
INVx1_ASAP7_75t_L g626 ( .A(n_538), .Y(n_626) );
INVx1_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
OR2x2_ASAP7_75t_L g540 ( .A(n_541), .B(n_556), .Y(n_540) );
INVx1_ASAP7_75t_L g614 ( .A(n_541), .Y(n_614) );
BUFx2_ASAP7_75t_L g541 ( .A(n_542), .Y(n_541) );
AND2x2_ASAP7_75t_L g694 ( .A(n_542), .B(n_575), .Y(n_694) );
AND2x2_ASAP7_75t_L g713 ( .A(n_542), .B(n_620), .Y(n_713) );
INVx2_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
INVx1_ASAP7_75t_L g581 ( .A(n_543), .Y(n_581) );
BUFx3_ASAP7_75t_L g619 ( .A(n_543), .Y(n_619) );
AND2x2_ASAP7_75t_L g648 ( .A(n_543), .B(n_649), .Y(n_648) );
NAND2x1p5_ASAP7_75t_L g543 ( .A(n_544), .B(n_545), .Y(n_543) );
OAI21x1_ASAP7_75t_L g545 ( .A1(n_546), .A2(n_551), .B(n_554), .Y(n_545) );
INVx2_ASAP7_75t_SL g549 ( .A(n_550), .Y(n_549) );
INVx2_ASAP7_75t_L g741 ( .A(n_556), .Y(n_741) );
OR2x2_ASAP7_75t_L g556 ( .A(n_557), .B(n_570), .Y(n_556) );
INVx2_ASAP7_75t_L g609 ( .A(n_557), .Y(n_609) );
INVx2_ASAP7_75t_L g557 ( .A(n_558), .Y(n_557) );
INVx1_ASAP7_75t_L g588 ( .A(n_558), .Y(n_588) );
OAI21xp5_ASAP7_75t_L g560 ( .A1(n_561), .A2(n_563), .B(n_565), .Y(n_560) );
INVx1_ASAP7_75t_L g589 ( .A(n_570), .Y(n_589) );
INVx3_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
OR2x6_ASAP7_75t_L g572 ( .A(n_573), .B(n_580), .Y(n_572) );
INVx2_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
AND2x2_ASAP7_75t_L g628 ( .A(n_574), .B(n_629), .Y(n_628) );
BUFx2_ASAP7_75t_L g758 ( .A(n_574), .Y(n_758) );
INVx1_ASAP7_75t_L g603 ( .A(n_575), .Y(n_603) );
AND2x2_ASAP7_75t_L g683 ( .A(n_575), .B(n_621), .Y(n_683) );
INVx2_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
AND2x2_ASAP7_75t_L g620 ( .A(n_576), .B(n_621), .Y(n_620) );
AOI21x1_ASAP7_75t_L g576 ( .A1(n_577), .A2(n_578), .B(n_579), .Y(n_576) );
INVx1_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
NOR2x1_ASAP7_75t_L g632 ( .A(n_581), .B(n_633), .Y(n_632) );
INVx2_ASAP7_75t_L g716 ( .A(n_581), .Y(n_716) );
NAND2xp5_ASAP7_75t_L g582 ( .A(n_583), .B(n_590), .Y(n_582) );
OAI22xp5_ASAP7_75t_L g623 ( .A1(n_583), .A2(n_624), .B1(n_627), .B2(n_631), .Y(n_623) );
INVx1_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
AOI22xp5_ASAP7_75t_L g641 ( .A1(n_584), .A2(n_604), .B1(n_636), .B2(n_642), .Y(n_641) );
AND2x2_ASAP7_75t_L g584 ( .A(n_585), .B(n_586), .Y(n_584) );
BUFx2_ASAP7_75t_SL g622 ( .A(n_585), .Y(n_622) );
AND2x4_ASAP7_75t_L g740 ( .A(n_585), .B(n_741), .Y(n_740) );
INVx1_ASAP7_75t_L g749 ( .A(n_585), .Y(n_749) );
INVx1_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
INVx1_ASAP7_75t_L g661 ( .A(n_587), .Y(n_661) );
OR2x2_ASAP7_75t_L g587 ( .A(n_588), .B(n_589), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g719 ( .A(n_588), .B(n_593), .Y(n_719) );
INVxp67_ASAP7_75t_L g748 ( .A(n_588), .Y(n_748) );
AND2x2_ASAP7_75t_L g753 ( .A(n_588), .B(n_619), .Y(n_753) );
OR2x2_ASAP7_75t_L g735 ( .A(n_589), .B(n_609), .Y(n_735) );
INVx1_ASAP7_75t_L g616 ( .A(n_590), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g590 ( .A(n_591), .B(n_592), .Y(n_590) );
NAND2xp5_ASAP7_75t_L g673 ( .A(n_591), .B(n_674), .Y(n_673) );
AND2x2_ASAP7_75t_L g655 ( .A(n_592), .B(n_640), .Y(n_655) );
AND2x4_ASAP7_75t_L g592 ( .A(n_593), .B(n_594), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g608 ( .A(n_593), .B(n_609), .Y(n_608) );
INVx2_ASAP7_75t_L g639 ( .A(n_593), .Y(n_639) );
OR2x2_ASAP7_75t_L g734 ( .A(n_593), .B(n_735), .Y(n_734) );
OAI21xp33_ASAP7_75t_L g595 ( .A1(n_596), .A2(n_600), .B(n_605), .Y(n_595) );
INVx1_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
INVx2_ASAP7_75t_L g658 ( .A(n_597), .Y(n_658) );
OR2x2_ASAP7_75t_L g597 ( .A(n_598), .B(n_599), .Y(n_597) );
AND2x2_ASAP7_75t_L g652 ( .A(n_598), .B(n_649), .Y(n_652) );
INVx2_ASAP7_75t_L g776 ( .A(n_598), .Y(n_776) );
INVx2_ASAP7_75t_SL g600 ( .A(n_601), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g601 ( .A(n_602), .B(n_604), .Y(n_601) );
AND2x2_ASAP7_75t_L g705 ( .A(n_602), .B(n_648), .Y(n_705) );
AND2x2_ASAP7_75t_L g730 ( .A(n_602), .B(n_676), .Y(n_730) );
INVx1_ASAP7_75t_L g602 ( .A(n_603), .Y(n_602) );
INVx2_ASAP7_75t_L g633 ( .A(n_603), .Y(n_633) );
AND2x2_ASAP7_75t_L g660 ( .A(n_604), .B(n_614), .Y(n_660) );
NAND2xp5_ASAP7_75t_L g672 ( .A(n_604), .B(n_659), .Y(n_672) );
INVx1_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
OR2x2_ASAP7_75t_L g606 ( .A(n_607), .B(n_608), .Y(n_606) );
INVx1_ASAP7_75t_L g757 ( .A(n_607), .Y(n_757) );
OR2x2_ASAP7_75t_L g773 ( .A(n_607), .B(n_668), .Y(n_773) );
INVx1_ASAP7_75t_L g697 ( .A(n_609), .Y(n_697) );
NAND3xp33_ASAP7_75t_L g610 ( .A(n_611), .B(n_634), .C(n_656), .Y(n_610) );
AOI221xp5_ASAP7_75t_L g611 ( .A1(n_612), .A2(n_616), .B1(n_617), .B2(n_622), .C(n_623), .Y(n_611) );
INVx1_ASAP7_75t_L g612 ( .A(n_613), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g613 ( .A(n_614), .B(n_615), .Y(n_613) );
AND2x2_ASAP7_75t_L g636 ( .A(n_615), .B(n_637), .Y(n_636) );
NAND2xp5_ASAP7_75t_L g764 ( .A(n_615), .B(n_680), .Y(n_764) );
AND2x2_ASAP7_75t_L g617 ( .A(n_618), .B(n_620), .Y(n_617) );
BUFx2_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
INVx3_ASAP7_75t_L g659 ( .A(n_619), .Y(n_659) );
AND3x1_ASAP7_75t_L g755 ( .A(n_619), .B(n_756), .C(n_757), .Y(n_755) );
AND2x2_ASAP7_75t_L g742 ( .A(n_620), .B(n_743), .Y(n_742) );
INVx2_ASAP7_75t_L g752 ( .A(n_620), .Y(n_752) );
INVxp67_ASAP7_75t_L g766 ( .A(n_622), .Y(n_766) );
OR2x2_ASAP7_75t_L g624 ( .A(n_625), .B(n_626), .Y(n_624) );
OR2x2_ASAP7_75t_L g721 ( .A(n_625), .B(n_645), .Y(n_721) );
INVx2_ASAP7_75t_L g756 ( .A(n_625), .Y(n_756) );
INVx1_ASAP7_75t_L g674 ( .A(n_626), .Y(n_674) );
INVx1_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
OAI21xp5_ASAP7_75t_L g675 ( .A1(n_628), .A2(n_676), .B(n_677), .Y(n_675) );
NAND2xp5_ASAP7_75t_L g775 ( .A(n_629), .B(n_776), .Y(n_775) );
INVx1_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
INVx1_ASAP7_75t_L g637 ( .A(n_630), .Y(n_637) );
OR2x2_ASAP7_75t_L g731 ( .A(n_630), .B(n_732), .Y(n_731) );
INVxp67_ASAP7_75t_SL g631 ( .A(n_632), .Y(n_631) );
INVx1_ASAP7_75t_L g691 ( .A(n_633), .Y(n_691) );
NAND2xp5_ASAP7_75t_L g770 ( .A(n_633), .B(n_690), .Y(n_770) );
AND3x1_ASAP7_75t_L g634 ( .A(n_635), .B(n_641), .C(n_646), .Y(n_634) );
NAND2xp5_ASAP7_75t_L g635 ( .A(n_636), .B(n_638), .Y(n_635) );
AND2x2_ASAP7_75t_L g685 ( .A(n_637), .B(n_676), .Y(n_685) );
AOI22xp5_ASAP7_75t_L g704 ( .A1(n_638), .A2(n_705), .B1(n_706), .B2(n_708), .Y(n_704) );
AND2x2_ASAP7_75t_L g638 ( .A(n_639), .B(n_640), .Y(n_638) );
OAI321xp33_ASAP7_75t_L g727 ( .A1(n_639), .A2(n_728), .A3(n_729), .B1(n_731), .B2(n_734), .C(n_736), .Y(n_727) );
AND2x2_ASAP7_75t_L g779 ( .A(n_639), .B(n_644), .Y(n_779) );
AND2x2_ASAP7_75t_L g677 ( .A(n_640), .B(n_643), .Y(n_677) );
INVx2_ASAP7_75t_L g686 ( .A(n_642), .Y(n_686) );
AND2x2_ASAP7_75t_L g695 ( .A(n_642), .B(n_696), .Y(n_695) );
AND2x4_ASAP7_75t_L g642 ( .A(n_643), .B(n_644), .Y(n_642) );
INVx2_ASAP7_75t_L g644 ( .A(n_645), .Y(n_644) );
OR2x2_ASAP7_75t_L g707 ( .A(n_645), .B(n_697), .Y(n_707) );
INVx2_ASAP7_75t_L g739 ( .A(n_645), .Y(n_739) );
OAI21xp33_ASAP7_75t_L g646 ( .A1(n_647), .A2(n_650), .B(n_655), .Y(n_646) );
HB1xp67_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
INVx1_ASAP7_75t_L g743 ( .A(n_649), .Y(n_743) );
NAND2xp5_ASAP7_75t_SL g650 ( .A(n_651), .B(n_653), .Y(n_650) );
INVx1_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
NAND2x1p5_ASAP7_75t_L g669 ( .A(n_652), .B(n_659), .Y(n_669) );
INVxp67_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
OAI21xp5_ASAP7_75t_L g656 ( .A1(n_657), .A2(n_660), .B(n_661), .Y(n_656) );
AND2x2_ASAP7_75t_L g657 ( .A(n_658), .B(n_659), .Y(n_657) );
NAND2xp5_ASAP7_75t_L g709 ( .A(n_659), .B(n_683), .Y(n_709) );
NAND2xp5_ASAP7_75t_L g723 ( .A(n_659), .B(n_724), .Y(n_723) );
AND2x2_ASAP7_75t_L g760 ( .A(n_659), .B(n_761), .Y(n_760) );
INVx1_ASAP7_75t_L g728 ( .A(n_661), .Y(n_728) );
NOR2xp67_ASAP7_75t_L g662 ( .A(n_663), .B(n_725), .Y(n_662) );
NAND3xp33_ASAP7_75t_L g663 ( .A(n_664), .B(n_687), .C(n_710), .Y(n_663) );
NOR2xp33_ASAP7_75t_L g664 ( .A(n_665), .B(n_678), .Y(n_664) );
OAI221xp5_ASAP7_75t_L g665 ( .A1(n_666), .A2(n_669), .B1(n_670), .B2(n_673), .C(n_675), .Y(n_665) );
OR2x2_ASAP7_75t_L g666 ( .A(n_667), .B(n_668), .Y(n_666) );
OR2x2_ASAP7_75t_L g718 ( .A(n_667), .B(n_719), .Y(n_718) );
INVx1_ASAP7_75t_L g670 ( .A(n_671), .Y(n_670) );
INVx1_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
AOI21xp33_ASAP7_75t_SL g678 ( .A1(n_679), .A2(n_684), .B(n_686), .Y(n_678) );
NAND2xp5_ASAP7_75t_L g679 ( .A(n_680), .B(n_681), .Y(n_679) );
INVx1_ASAP7_75t_L g681 ( .A(n_682), .Y(n_681) );
INVx2_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
AND2x2_ASAP7_75t_L g715 ( .A(n_683), .B(n_716), .Y(n_715) );
OAI21xp33_ASAP7_75t_SL g698 ( .A1(n_684), .A2(n_699), .B(n_704), .Y(n_698) );
INVx2_ASAP7_75t_SL g684 ( .A(n_685), .Y(n_684) );
O2A1O1Ixp33_ASAP7_75t_L g687 ( .A1(n_688), .A2(n_692), .B(n_695), .C(n_698), .Y(n_687) );
INVx2_ASAP7_75t_SL g688 ( .A(n_689), .Y(n_688) );
NAND2xp5_ASAP7_75t_L g763 ( .A(n_689), .B(n_764), .Y(n_763) );
NAND2x1_ASAP7_75t_L g689 ( .A(n_690), .B(n_691), .Y(n_689) );
INVx1_ASAP7_75t_L g692 ( .A(n_693), .Y(n_692) );
INVx1_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
INVx1_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
NAND2xp5_ASAP7_75t_L g738 ( .A(n_697), .B(n_739), .Y(n_738) );
INVxp67_ASAP7_75t_L g699 ( .A(n_700), .Y(n_699) );
NAND2xp5_ASAP7_75t_SL g759 ( .A(n_700), .B(n_760), .Y(n_759) );
INVx2_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
NAND2xp5_ASAP7_75t_L g701 ( .A(n_702), .B(n_703), .Y(n_701) );
INVx2_ASAP7_75t_L g706 ( .A(n_707), .Y(n_706) );
INVx1_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
AOI22xp5_ASAP7_75t_L g710 ( .A1(n_711), .A2(n_717), .B1(n_720), .B2(n_722), .Y(n_710) );
INVx1_ASAP7_75t_L g712 ( .A(n_713), .Y(n_712) );
INVx1_ASAP7_75t_L g714 ( .A(n_715), .Y(n_714) );
INVx1_ASAP7_75t_L g717 ( .A(n_718), .Y(n_717) );
HB1xp67_ASAP7_75t_L g782 ( .A(n_719), .Y(n_782) );
INVx1_ASAP7_75t_L g720 ( .A(n_721), .Y(n_720) );
INVx1_ASAP7_75t_L g722 ( .A(n_723), .Y(n_722) );
NAND3xp33_ASAP7_75t_L g725 ( .A(n_726), .B(n_762), .C(n_777), .Y(n_725) );
NOR2xp33_ASAP7_75t_L g726 ( .A(n_727), .B(n_744), .Y(n_726) );
INVx2_ASAP7_75t_L g729 ( .A(n_730), .Y(n_729) );
INVx2_ASAP7_75t_SL g732 ( .A(n_733), .Y(n_732) );
OAI21xp33_ASAP7_75t_L g736 ( .A1(n_737), .A2(n_740), .B(n_742), .Y(n_736) );
INVx1_ASAP7_75t_L g737 ( .A(n_738), .Y(n_737) );
NAND3xp33_ASAP7_75t_L g744 ( .A(n_745), .B(n_750), .C(n_759), .Y(n_744) );
INVx1_ASAP7_75t_L g746 ( .A(n_747), .Y(n_746) );
OR2x2_ASAP7_75t_L g747 ( .A(n_748), .B(n_749), .Y(n_747) );
AOI32xp33_ASAP7_75t_L g750 ( .A1(n_751), .A2(n_753), .A3(n_754), .B1(n_755), .B2(n_758), .Y(n_750) );
INVx3_ASAP7_75t_L g751 ( .A(n_752), .Y(n_751) );
AND2x2_ASAP7_75t_L g778 ( .A(n_753), .B(n_779), .Y(n_778) );
AOI21xp5_ASAP7_75t_L g762 ( .A1(n_763), .A2(n_765), .B(n_767), .Y(n_762) );
INVx1_ASAP7_75t_L g767 ( .A(n_768), .Y(n_767) );
AOI22x1_ASAP7_75t_L g768 ( .A1(n_769), .A2(n_771), .B1(n_772), .B2(n_774), .Y(n_768) );
INVx1_ASAP7_75t_L g769 ( .A(n_770), .Y(n_769) );
AOI21xp33_ASAP7_75t_L g781 ( .A1(n_770), .A2(n_782), .B(n_783), .Y(n_781) );
INVx2_ASAP7_75t_L g772 ( .A(n_773), .Y(n_772) );
INVx1_ASAP7_75t_L g774 ( .A(n_775), .Y(n_774) );
AOI21xp5_ASAP7_75t_L g777 ( .A1(n_778), .A2(n_780), .B(n_781), .Y(n_777) );
INVx1_ASAP7_75t_L g783 ( .A(n_784), .Y(n_783) );
INVx8_ASAP7_75t_L g785 ( .A(n_786), .Y(n_785) );
BUFx12f_ASAP7_75t_L g786 ( .A(n_787), .Y(n_786) );
INVx2_ASAP7_75t_L g790 ( .A(n_791), .Y(n_790) );
INVx5_ASAP7_75t_L g791 ( .A(n_792), .Y(n_791) );
AND2x6_ASAP7_75t_SL g792 ( .A(n_793), .B(n_795), .Y(n_792) );
INVx1_ASAP7_75t_L g793 ( .A(n_794), .Y(n_793) );
INVx3_ASAP7_75t_L g804 ( .A(n_794), .Y(n_804) );
NOR2xp33_ASAP7_75t_L g830 ( .A(n_794), .B(n_831), .Y(n_830) );
NAND2xp5_ASAP7_75t_L g795 ( .A(n_796), .B(n_798), .Y(n_795) );
INVx1_ASAP7_75t_L g796 ( .A(n_797), .Y(n_796) );
NOR2x1_ASAP7_75t_L g833 ( .A(n_797), .B(n_799), .Y(n_833) );
AND2x6_ASAP7_75t_SL g809 ( .A(n_798), .B(n_810), .Y(n_809) );
INVx1_ASAP7_75t_L g798 ( .A(n_799), .Y(n_798) );
OAI21x1_ASAP7_75t_SL g800 ( .A1(n_801), .A2(n_805), .B(n_826), .Y(n_800) );
INVx1_ASAP7_75t_SL g801 ( .A(n_802), .Y(n_801) );
CKINVDCx11_ASAP7_75t_R g802 ( .A(n_803), .Y(n_802) );
BUFx6f_ASAP7_75t_L g803 ( .A(n_804), .Y(n_803) );
AOI21xp5_ASAP7_75t_L g805 ( .A1(n_806), .A2(n_818), .B(n_819), .Y(n_805) );
AND2x2_ASAP7_75t_L g806 ( .A(n_807), .B(n_813), .Y(n_806) );
BUFx12f_ASAP7_75t_L g807 ( .A(n_808), .Y(n_807) );
INVx4_ASAP7_75t_L g808 ( .A(n_809), .Y(n_808) );
INVx3_ASAP7_75t_L g821 ( .A(n_809), .Y(n_821) );
INVx1_ASAP7_75t_L g811 ( .A(n_812), .Y(n_811) );
HB1xp67_ASAP7_75t_L g842 ( .A(n_812), .Y(n_842) );
OAI31xp33_ASAP7_75t_SL g819 ( .A1(n_813), .A2(n_818), .A3(n_820), .B(n_822), .Y(n_819) );
CKINVDCx5p33_ASAP7_75t_R g815 ( .A(n_816), .Y(n_815) );
INVx2_ASAP7_75t_L g820 ( .A(n_821), .Y(n_820) );
BUFx2_ASAP7_75t_SL g824 ( .A(n_821), .Y(n_824) );
INVxp67_ASAP7_75t_L g822 ( .A(n_823), .Y(n_822) );
NOR2xp33_ASAP7_75t_L g823 ( .A(n_824), .B(n_825), .Y(n_823) );
INVx1_ASAP7_75t_L g827 ( .A(n_828), .Y(n_827) );
INVx2_ASAP7_75t_L g828 ( .A(n_829), .Y(n_828) );
BUFx10_ASAP7_75t_L g829 ( .A(n_830), .Y(n_829) );
INVx1_ASAP7_75t_L g831 ( .A(n_832), .Y(n_831) );
INVx1_ASAP7_75t_SL g834 ( .A(n_835), .Y(n_834) );
INVx2_ASAP7_75t_L g835 ( .A(n_836), .Y(n_835) );
AND2x4_ASAP7_75t_L g836 ( .A(n_837), .B(n_841), .Y(n_836) );
AND2x4_ASAP7_75t_L g849 ( .A(n_837), .B(n_841), .Y(n_849) );
INVx1_ASAP7_75t_L g837 ( .A(n_838), .Y(n_837) );
NAND2xp5_ASAP7_75t_L g838 ( .A(n_839), .B(n_840), .Y(n_838) );
NOR2x1p5_ASAP7_75t_L g841 ( .A(n_842), .B(n_843), .Y(n_841) );
NAND2xp5_ASAP7_75t_L g843 ( .A(n_844), .B(n_845), .Y(n_843) );
INVx3_ASAP7_75t_L g847 ( .A(n_848), .Y(n_847) );
BUFx6f_ASAP7_75t_SL g848 ( .A(n_849), .Y(n_848) );
endmodule