module fake_jpeg_435_n_88 (n_13, n_21, n_1, n_10, n_23, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_9, n_5, n_11, n_17, n_25, n_2, n_12, n_8, n_15, n_7, n_88);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_88;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_57;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_44;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_12),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_21),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_9),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_23),
.Y(n_30)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_25),
.Y(n_31)
);

HB1xp67_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_11),
.Y(n_33)
);

INVx5_ASAP7_75t_L g34 ( 
.A(n_31),
.Y(n_34)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_34),
.Y(n_48)
);

INVx13_ASAP7_75t_L g35 ( 
.A(n_26),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_35),
.B(n_36),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_32),
.Y(n_36)
);

INVx2_ASAP7_75t_SL g37 ( 
.A(n_29),
.Y(n_37)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_37),
.Y(n_47)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_31),
.Y(n_38)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_38),
.Y(n_44)
);

INVx11_ASAP7_75t_L g39 ( 
.A(n_33),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_39),
.B(n_27),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_37),
.B(n_30),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_40),
.B(n_43),
.Y(n_51)
);

O2A1O1Ixp33_ASAP7_75t_L g42 ( 
.A1(n_38),
.A2(n_30),
.B(n_29),
.C(n_28),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_42),
.A2(n_0),
.B1(n_3),
.B2(n_4),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_34),
.B(n_28),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_35),
.B(n_27),
.Y(n_45)
);

CKINVDCx14_ASAP7_75t_R g52 ( 
.A(n_45),
.Y(n_52)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_46),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_L g50 ( 
.A1(n_47),
.A2(n_39),
.B1(n_1),
.B2(n_2),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_L g63 ( 
.A1(n_50),
.A2(n_54),
.B1(n_5),
.B2(n_6),
.Y(n_63)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_48),
.Y(n_53)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_53),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_44),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_54)
);

BUFx2_ASAP7_75t_L g55 ( 
.A(n_48),
.Y(n_55)
);

HB1xp67_ASAP7_75t_L g67 ( 
.A(n_55),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_41),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_56),
.B(n_4),
.Y(n_61)
);

INVxp67_ASAP7_75t_L g64 ( 
.A(n_57),
.Y(n_64)
);

XNOR2xp5_ASAP7_75t_L g59 ( 
.A(n_51),
.B(n_42),
.Y(n_59)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_59),
.B(n_60),
.C(n_62),
.Y(n_71)
);

XNOR2xp5_ASAP7_75t_L g60 ( 
.A(n_49),
.B(n_3),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_61),
.B(n_66),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_52),
.B(n_17),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_62),
.B(n_63),
.Y(n_74)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_55),
.Y(n_65)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_65),
.Y(n_73)
);

OR2x2_ASAP7_75t_L g66 ( 
.A(n_57),
.B(n_5),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_64),
.A2(n_50),
.B1(n_53),
.B2(n_13),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_69),
.A2(n_75),
.B1(n_74),
.B2(n_72),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_67),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_70),
.B(n_72),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_R g79 ( 
.A(n_71),
.B(n_16),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g72 ( 
.A(n_58),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_64),
.A2(n_7),
.B1(n_10),
.B2(n_15),
.Y(n_75)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_73),
.Y(n_76)
);

INVxp33_ASAP7_75t_L g82 ( 
.A(n_76),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_68),
.B(n_24),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_77),
.B(n_78),
.Y(n_81)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_82),
.Y(n_83)
);

AOI31xp67_ASAP7_75t_SL g84 ( 
.A1(n_83),
.A2(n_80),
.A3(n_81),
.B(n_77),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_84),
.B(n_79),
.C(n_19),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_85),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_SL g87 ( 
.A1(n_86),
.A2(n_18),
.B(n_20),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_87),
.B(n_22),
.Y(n_88)
);


endmodule