module real_jpeg_12331_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_54;
wire n_37;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_68;
wire n_83;
wire n_78;
wire n_64;
wire n_47;
wire n_22;
wire n_87;
wire n_40;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_13;
wire n_93;
wire n_95;
wire n_65;
wire n_33;
wire n_76;
wire n_67;
wire n_79;
wire n_66;
wire n_28;
wire n_44;
wire n_62;
wire n_45;
wire n_42;
wire n_18;
wire n_77;
wire n_39;
wire n_94;
wire n_26;
wire n_19;
wire n_17;
wire n_21;
wire n_50;
wire n_69;
wire n_31;
wire n_72;
wire n_100;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_30;
wire n_15;
wire n_57;
wire n_43;
wire n_84;
wire n_82;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_24;
wire n_92;
wire n_97;
wire n_75;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_25;
wire n_53;
wire n_36;
wire n_81;
wire n_85;
wire n_101;
wire n_96;
wire n_89;
wire n_16;

BUFx2_ASAP7_75t_L g44 ( 
.A(n_0),
.Y(n_44)
);

BUFx4f_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

OAI22xp5_ASAP7_75t_L g33 ( 
.A1(n_3),
.A2(n_20),
.B1(n_23),
.B2(n_34),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_3),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_L g84 ( 
.A1(n_3),
.A2(n_29),
.B1(n_31),
.B2(n_34),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_4),
.A2(n_29),
.B1(n_31),
.B2(n_49),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_4),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_5),
.Y(n_55)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_6),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_7),
.B(n_37),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_7),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_7),
.A2(n_20),
.B1(n_23),
.B2(n_56),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_7),
.A2(n_42),
.B1(n_61),
.B2(n_91),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g19 ( 
.A1(n_8),
.A2(n_20),
.B1(n_22),
.B2(n_23),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_8),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_8),
.A2(n_22),
.B1(n_55),
.B2(n_58),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_8),
.A2(n_22),
.B1(n_29),
.B2(n_31),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g62 ( 
.A1(n_9),
.A2(n_29),
.B1(n_31),
.B2(n_63),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_9),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g45 ( 
.A1(n_10),
.A2(n_29),
.B1(n_31),
.B2(n_46),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_10),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_10),
.A2(n_20),
.B1(n_23),
.B2(n_46),
.Y(n_66)
);

INVx11_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

XOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_72),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_71),
.Y(n_13)
);

INVxp67_ASAP7_75t_L g14 ( 
.A(n_15),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_50),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_16),
.B(n_50),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_35),
.C(n_41),
.Y(n_16)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_17),
.A2(n_18),
.B1(n_35),
.B2(n_36),
.Y(n_100)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

AOI22xp5_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_24),
.B1(n_32),
.B2(n_33),
.Y(n_18)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_19),
.A2(n_24),
.B1(n_32),
.B2(n_79),
.Y(n_78)
);

INVx6_ASAP7_75t_SL g23 ( 
.A(n_20),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_L g25 ( 
.A1(n_20),
.A2(n_23),
.B1(n_26),
.B2(n_27),
.Y(n_25)
);

OA22x2_ASAP7_75t_SL g38 ( 
.A1(n_20),
.A2(n_23),
.B1(n_39),
.B2(n_40),
.Y(n_38)
);

NOR3xp33_ASAP7_75t_L g57 ( 
.A(n_20),
.B(n_40),
.C(n_58),
.Y(n_57)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

O2A1O1Ixp33_ASAP7_75t_SL g52 ( 
.A1(n_23),
.A2(n_39),
.B(n_53),
.C(n_57),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_23),
.B(n_77),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_24),
.A2(n_32),
.B1(n_33),
.B2(n_66),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_28),
.Y(n_24)
);

INVx13_ASAP7_75t_L g27 ( 
.A(n_26),
.Y(n_27)
);

OA22x2_ASAP7_75t_L g28 ( 
.A1(n_26),
.A2(n_27),
.B1(n_29),
.B2(n_31),
.Y(n_28)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_27),
.B(n_31),
.C(n_56),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_28),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_28),
.B(n_56),
.Y(n_94)
);

CKINVDCx6p67_ASAP7_75t_R g31 ( 
.A(n_29),
.Y(n_31)
);

INVx5_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_31),
.B(n_44),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_31),
.B(n_89),
.Y(n_88)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_37),
.A2(n_54),
.B1(n_68),
.B2(n_70),
.Y(n_67)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

AND2x2_ASAP7_75t_L g68 ( 
.A(n_38),
.B(n_69),
.Y(n_68)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_39),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_39),
.A2(n_40),
.B1(n_55),
.B2(n_58),
.Y(n_69)
);

XNOR2xp5_ASAP7_75t_L g99 ( 
.A(n_41),
.B(n_100),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_L g41 ( 
.A1(n_42),
.A2(n_45),
.B(n_47),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_42),
.A2(n_61),
.B1(n_84),
.B2(n_91),
.Y(n_93)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

AOI21xp5_ASAP7_75t_L g59 ( 
.A1(n_43),
.A2(n_48),
.B(n_60),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_43),
.A2(n_44),
.B1(n_83),
.B2(n_85),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_44),
.B(n_48),
.Y(n_47)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_44),
.Y(n_61)
);

CKINVDCx16_ASAP7_75t_R g85 ( 
.A(n_45),
.Y(n_85)
);

XOR2xp5_ASAP7_75t_L g50 ( 
.A(n_51),
.B(n_64),
.Y(n_50)
);

XNOR2xp5_ASAP7_75t_SL g51 ( 
.A(n_52),
.B(n_59),
.Y(n_51)
);

CKINVDCx5p33_ASAP7_75t_R g53 ( 
.A(n_54),
.Y(n_53)
);

HAxp5_ASAP7_75t_SL g54 ( 
.A(n_55),
.B(n_56),
.CON(n_54),
.SN(n_54)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_55),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_56),
.B(n_61),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_61),
.B(n_62),
.Y(n_60)
);

XOR2xp5_ASAP7_75t_L g64 ( 
.A(n_65),
.B(n_67),
.Y(n_64)
);

OAI21xp5_ASAP7_75t_L g72 ( 
.A1(n_73),
.A2(n_97),
.B(n_101),
.Y(n_72)
);

AOI21xp5_ASAP7_75t_L g73 ( 
.A1(n_74),
.A2(n_86),
.B(n_96),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_75),
.B(n_82),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_75),
.B(n_82),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_76),
.A2(n_78),
.B1(n_80),
.B2(n_81),
.Y(n_75)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_76),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_78),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_78),
.B(n_80),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

OAI21xp5_ASAP7_75t_L g86 ( 
.A1(n_87),
.A2(n_92),
.B(n_95),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_90),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_93),
.B(n_94),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_93),
.B(n_94),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_99),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_98),
.B(n_99),
.Y(n_101)
);


endmodule