module real_jpeg_12857_n_18 (n_17, n_8, n_0, n_2, n_297, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_18);

input n_17;
input n_8;
input n_0;
input n_2;
input n_297;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_18;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_201;
wire n_114;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_249;
wire n_166;
wire n_176;
wire n_215;
wire n_221;
wire n_292;
wire n_286;
wire n_288;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_280;
wire n_64;
wire n_177;
wire n_291;
wire n_236;
wire n_271;
wire n_47;
wire n_281;
wire n_131;
wire n_163;
wire n_276;
wire n_22;
wire n_287;
wire n_237;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_243;
wire n_255;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_293;
wire n_275;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_188;
wire n_139;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_290;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_172;
wire n_211;
wire n_160;
wire n_45;
wire n_285;
wire n_112;
wire n_42;
wire n_268;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_294;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_203;
wire n_198;
wire n_100;
wire n_192;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_110;
wire n_195;
wire n_61;
wire n_205;
wire n_258;
wire n_289;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_278;
wire n_130;
wire n_144;
wire n_241;
wire n_103;
wire n_259;
wire n_225;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_284;
wire n_226;
wire n_277;
wire n_125;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_240;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_97;
wire n_187;
wire n_75;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_279;
wire n_167;
wire n_295;
wire n_202;
wire n_128;
wire n_179;
wire n_216;
wire n_133;
wire n_213;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_181;
wire n_283;
wire n_101;
wire n_256;
wire n_274;
wire n_182;
wire n_269;
wire n_96;
wire n_253;
wire n_273;
wire n_89;

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

BUFx16f_ASAP7_75t_L g49 ( 
.A(n_1),
.Y(n_49)
);

BUFx12_ASAP7_75t_L g67 ( 
.A(n_2),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_3),
.A2(n_65),
.B1(n_66),
.B2(n_69),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_3),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_3),
.A2(n_43),
.B1(n_44),
.B2(n_69),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_SL g167 ( 
.A1(n_3),
.A2(n_60),
.B1(n_63),
.B2(n_69),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_3),
.A2(n_29),
.B1(n_35),
.B2(n_69),
.Y(n_197)
);

AOI22xp33_ASAP7_75t_L g34 ( 
.A1(n_4),
.A2(n_29),
.B1(n_35),
.B2(n_36),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_4),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_4),
.A2(n_36),
.B1(n_43),
.B2(n_44),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_L g288 ( 
.A1(n_4),
.A2(n_36),
.B1(n_60),
.B2(n_63),
.Y(n_288)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_5),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_6),
.A2(n_60),
.B1(n_63),
.B2(n_80),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_6),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_6),
.A2(n_43),
.B1(n_44),
.B2(n_80),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_6),
.A2(n_65),
.B1(n_66),
.B2(n_80),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_6),
.A2(n_29),
.B1(n_35),
.B2(n_80),
.Y(n_142)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_7),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_L g42 ( 
.A1(n_8),
.A2(n_43),
.B1(n_44),
.B2(n_46),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_8),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_8),
.A2(n_46),
.B1(n_60),
.B2(n_63),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_8),
.A2(n_29),
.B1(n_35),
.B2(n_46),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_SL g281 ( 
.A1(n_8),
.A2(n_46),
.B1(n_65),
.B2(n_66),
.Y(n_281)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_9),
.A2(n_60),
.B1(n_63),
.B2(n_135),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_9),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_L g164 ( 
.A1(n_9),
.A2(n_65),
.B1(n_66),
.B2(n_135),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_9),
.A2(n_43),
.B1(n_44),
.B2(n_135),
.Y(n_188)
);

OAI22xp33_ASAP7_75t_SL g209 ( 
.A1(n_9),
.A2(n_29),
.B1(n_35),
.B2(n_135),
.Y(n_209)
);

BUFx12_ASAP7_75t_L g76 ( 
.A(n_10),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_11),
.B(n_140),
.Y(n_139)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_11),
.Y(n_153)
);

AOI21xp33_ASAP7_75t_L g161 ( 
.A1(n_11),
.A2(n_65),
.B(n_162),
.Y(n_161)
);

OAI22xp33_ASAP7_75t_L g187 ( 
.A1(n_11),
.A2(n_43),
.B1(n_44),
.B2(n_153),
.Y(n_187)
);

O2A1O1Ixp33_ASAP7_75t_L g189 ( 
.A1(n_11),
.A2(n_43),
.B(n_49),
.C(n_190),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_11),
.B(n_110),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_11),
.B(n_32),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_11),
.B(n_54),
.Y(n_214)
);

A2O1A1Ixp33_ASAP7_75t_L g223 ( 
.A1(n_11),
.A2(n_63),
.B(n_74),
.C(n_224),
.Y(n_223)
);

BUFx8_ASAP7_75t_L g62 ( 
.A(n_12),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g37 ( 
.A1(n_13),
.A2(n_29),
.B1(n_35),
.B2(n_38),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_13),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_13),
.A2(n_38),
.B1(n_43),
.B2(n_44),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g52 ( 
.A1(n_14),
.A2(n_43),
.B1(n_44),
.B2(n_53),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_14),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_14),
.A2(n_29),
.B1(n_35),
.B2(n_53),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_14),
.A2(n_53),
.B1(n_60),
.B2(n_63),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_15),
.A2(n_65),
.B1(n_66),
.B2(n_71),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_15),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_15),
.A2(n_60),
.B1(n_63),
.B2(n_71),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_15),
.A2(n_43),
.B1(n_44),
.B2(n_71),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_15),
.A2(n_29),
.B1(n_35),
.B2(n_71),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_16),
.A2(n_65),
.B1(n_66),
.B2(n_103),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_16),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_16),
.A2(n_60),
.B1(n_63),
.B2(n_103),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_16),
.A2(n_43),
.B1(n_44),
.B2(n_103),
.Y(n_195)
);

OAI22xp33_ASAP7_75t_SL g202 ( 
.A1(n_16),
.A2(n_29),
.B1(n_35),
.B2(n_103),
.Y(n_202)
);

INVx11_ASAP7_75t_L g30 ( 
.A(n_17),
.Y(n_30)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

OAI22xp5_ASAP7_75t_SL g19 ( 
.A1(n_20),
.A2(n_272),
.B1(n_294),
.B2(n_295),
.Y(n_19)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_20),
.Y(n_294)
);

OAI21xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_125),
.B(n_271),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_104),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_22),
.B(n_104),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_82),
.C(n_88),
.Y(n_22)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_23),
.B(n_82),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_25),
.B1(n_55),
.B2(n_56),
.Y(n_23)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_24),
.B(n_57),
.C(n_72),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_25),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_39),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_26),
.A2(n_27),
.B1(n_39),
.B2(n_40),
.Y(n_257)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g27 ( 
.A1(n_28),
.A2(n_32),
.B1(n_33),
.B2(n_37),
.Y(n_27)
);

OAI21xp5_ASAP7_75t_SL g84 ( 
.A1(n_28),
.A2(n_32),
.B(n_37),
.Y(n_84)
);

CKINVDCx16_ASAP7_75t_R g92 ( 
.A(n_28),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_28),
.A2(n_32),
.B1(n_142),
.B2(n_143),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_28),
.A2(n_32),
.B1(n_142),
.B2(n_156),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_28),
.A2(n_32),
.B1(n_94),
.B2(n_143),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_28),
.A2(n_32),
.B1(n_156),
.B2(n_197),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_28),
.A2(n_32),
.B1(n_153),
.B2(n_209),
.Y(n_208)
);

AOI22xp33_ASAP7_75t_L g213 ( 
.A1(n_28),
.A2(n_32),
.B1(n_202),
.B2(n_209),
.Y(n_213)
);

AND2x2_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_31),
.Y(n_28)
);

INVx3_ASAP7_75t_SL g35 ( 
.A(n_29),
.Y(n_35)
);

OA22x2_ASAP7_75t_L g51 ( 
.A1(n_29),
.A2(n_35),
.B1(n_49),
.B2(n_50),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_29),
.B(n_211),
.Y(n_210)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_31),
.A2(n_34),
.B1(n_92),
.B2(n_93),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_31),
.A2(n_92),
.B1(n_201),
.B2(n_203),
.Y(n_200)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVxp67_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

OAI21xp33_ASAP7_75t_L g190 ( 
.A1(n_35),
.A2(n_50),
.B(n_153),
.Y(n_190)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g40 ( 
.A1(n_41),
.A2(n_47),
.B1(n_52),
.B2(n_54),
.Y(n_40)
);

INVxp67_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_42),
.A2(n_51),
.B1(n_96),
.B2(n_98),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_43),
.A2(n_44),
.B1(n_49),
.B2(n_50),
.Y(n_48)
);

OA22x2_ASAP7_75t_L g78 ( 
.A1(n_43),
.A2(n_44),
.B1(n_76),
.B2(n_77),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_43),
.B(n_77),
.Y(n_154)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

OAI32xp33_ASAP7_75t_L g151 ( 
.A1(n_44),
.A2(n_63),
.A3(n_76),
.B1(n_152),
.B2(n_154),
.Y(n_151)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_47),
.A2(n_52),
.B1(n_54),
.B2(n_86),
.Y(n_85)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_47),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_47),
.A2(n_54),
.B1(n_86),
.B2(n_112),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_47),
.A2(n_54),
.B1(n_145),
.B2(n_147),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_47),
.A2(n_54),
.B1(n_97),
.B2(n_147),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_47),
.A2(n_54),
.B1(n_187),
.B2(n_188),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_47),
.A2(n_54),
.B1(n_188),
.B2(n_195),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_L g284 ( 
.A1(n_47),
.A2(n_54),
.B(n_112),
.Y(n_284)
);

AND2x2_ASAP7_75t_L g47 ( 
.A(n_48),
.B(n_51),
.Y(n_47)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_49),
.Y(n_50)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_51),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_51),
.A2(n_98),
.B1(n_146),
.B2(n_226),
.Y(n_225)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

XOR2xp5_ASAP7_75t_L g56 ( 
.A(n_57),
.B(n_72),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_58),
.A2(n_59),
.B1(n_68),
.B2(n_70),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_58),
.A2(n_59),
.B1(n_68),
.B2(n_102),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_58),
.A2(n_59),
.B1(n_70),
.B2(n_121),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_58),
.A2(n_59),
.B1(n_161),
.B2(n_164),
.Y(n_160)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_58),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_L g280 ( 
.A1(n_58),
.A2(n_59),
.B1(n_121),
.B2(n_281),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_59),
.B(n_64),
.Y(n_58)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_59),
.Y(n_140)
);

OA22x2_ASAP7_75t_L g59 ( 
.A1(n_60),
.A2(n_61),
.B1(n_62),
.B2(n_63),
.Y(n_59)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_60),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_60),
.A2(n_63),
.B1(n_76),
.B2(n_77),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_60),
.B(n_153),
.Y(n_152)
);

OAI32xp33_ASAP7_75t_L g176 ( 
.A1(n_60),
.A2(n_62),
.A3(n_65),
.B1(n_163),
.B2(n_177),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_61),
.A2(n_62),
.B1(n_65),
.B2(n_66),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_61),
.B(n_63),
.Y(n_177)
);

INVx11_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_66),
.B(n_153),
.Y(n_163)
);

BUFx16f_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_73),
.A2(n_78),
.B1(n_79),
.B2(n_81),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_73),
.A2(n_78),
.B1(n_79),
.B2(n_100),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_73),
.A2(n_78),
.B1(n_137),
.B2(n_167),
.Y(n_166)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_74),
.A2(n_108),
.B1(n_109),
.B2(n_110),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_74),
.A2(n_110),
.B1(n_133),
.B2(n_136),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_74),
.A2(n_110),
.B1(n_246),
.B2(n_247),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_74),
.A2(n_109),
.B1(n_110),
.B2(n_287),
.Y(n_286)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_75),
.B(n_78),
.Y(n_74)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_76),
.Y(n_77)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_78),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_L g222 ( 
.A1(n_78),
.A2(n_134),
.B(n_223),
.Y(n_222)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_81),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_83),
.A2(n_84),
.B1(n_85),
.B2(n_87),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_83),
.B(n_87),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_83),
.A2(n_84),
.B1(n_119),
.B2(n_120),
.Y(n_118)
);

CKINVDCx16_ASAP7_75t_R g83 ( 
.A(n_84),
.Y(n_83)
);

OAI21xp5_ASAP7_75t_L g276 ( 
.A1(n_84),
.A2(n_120),
.B(n_122),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_85),
.Y(n_87)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_88),
.B(n_269),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_99),
.C(n_101),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_89),
.A2(n_90),
.B1(n_259),
.B2(n_260),
.Y(n_258)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_95),
.Y(n_90)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_91),
.B(n_95),
.Y(n_242)
);

CKINVDCx16_ASAP7_75t_R g93 ( 
.A(n_94),
.Y(n_93)
);

CKINVDCx16_ASAP7_75t_R g96 ( 
.A(n_97),
.Y(n_96)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_99),
.B(n_101),
.Y(n_260)
);

INVxp67_ASAP7_75t_L g247 ( 
.A(n_100),
.Y(n_247)
);

INVxp67_ASAP7_75t_L g251 ( 
.A(n_102),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_124),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_106),
.A2(n_114),
.B1(n_115),
.B2(n_123),
.Y(n_105)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_106),
.Y(n_123)
);

OAI21xp33_ASAP7_75t_L g106 ( 
.A1(n_107),
.A2(n_111),
.B(n_113),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_107),
.B(n_111),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_113),
.A2(n_278),
.B1(n_290),
.B2(n_291),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_113),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_114),
.B(n_123),
.C(n_124),
.Y(n_292)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_116),
.A2(n_117),
.B1(n_118),
.B2(n_122),
.Y(n_115)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_116),
.Y(n_122)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

CKINVDCx14_ASAP7_75t_R g119 ( 
.A(n_120),
.Y(n_119)
);

AOI21xp5_ASAP7_75t_L g125 ( 
.A1(n_126),
.A2(n_266),
.B(n_270),
.Y(n_125)
);

OAI221xp5_ASAP7_75t_L g126 ( 
.A1(n_127),
.A2(n_253),
.B1(n_264),
.B2(n_265),
.C(n_297),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_128),
.B(n_237),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_L g128 ( 
.A1(n_129),
.A2(n_180),
.B(n_236),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_157),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_130),
.B(n_157),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_144),
.C(n_148),
.Y(n_130)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_131),
.B(n_233),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_SL g131 ( 
.A(n_132),
.B(n_138),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_132),
.B(n_139),
.C(n_141),
.Y(n_178)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_141),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_140),
.A2(n_249),
.B1(n_250),
.B2(n_251),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_L g233 ( 
.A1(n_144),
.A2(n_148),
.B1(n_149),
.B2(n_234),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_144),
.Y(n_234)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_155),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_150),
.A2(n_151),
.B1(n_155),
.B2(n_228),
.Y(n_227)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

CKINVDCx16_ASAP7_75t_R g224 ( 
.A(n_152),
.Y(n_224)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_155),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_158),
.A2(n_159),
.B1(n_171),
.B2(n_179),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_158),
.B(n_172),
.C(n_178),
.Y(n_238)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_165),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_160),
.B(n_166),
.C(n_170),
.Y(n_241)
);

CKINVDCx16_ASAP7_75t_R g162 ( 
.A(n_163),
.Y(n_162)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_164),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_166),
.A2(n_168),
.B1(n_169),
.B2(n_170),
.Y(n_165)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_166),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g246 ( 
.A(n_167),
.Y(n_246)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_168),
.Y(n_170)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_171),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_SL g171 ( 
.A(n_172),
.B(n_178),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_173),
.A2(n_174),
.B1(n_175),
.B2(n_176),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_173),
.B(n_176),
.Y(n_252)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

AOI21xp5_ASAP7_75t_L g180 ( 
.A1(n_181),
.A2(n_230),
.B(n_235),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_SL g181 ( 
.A1(n_182),
.A2(n_218),
.B(n_229),
.Y(n_181)
);

AOI21xp5_ASAP7_75t_L g182 ( 
.A1(n_183),
.A2(n_198),
.B(n_217),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_191),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_SL g217 ( 
.A(n_184),
.B(n_191),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_185),
.B(n_189),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_185),
.A2(n_186),
.B1(n_189),
.B2(n_205),
.Y(n_204)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_189),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_196),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_194),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_193),
.B(n_194),
.C(n_196),
.Y(n_219)
);

INVxp67_ASAP7_75t_L g226 ( 
.A(n_195),
.Y(n_226)
);

INVxp67_ASAP7_75t_L g203 ( 
.A(n_197),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_SL g198 ( 
.A1(n_199),
.A2(n_206),
.B(n_216),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_204),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_200),
.B(n_204),
.Y(n_216)
);

INVxp67_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

AOI21xp5_ASAP7_75t_L g206 ( 
.A1(n_207),
.A2(n_212),
.B(n_215),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_SL g207 ( 
.A(n_208),
.B(n_210),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_214),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_SL g215 ( 
.A(n_213),
.B(n_214),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_220),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_219),
.B(n_220),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_227),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_225),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_222),
.B(n_225),
.C(n_227),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_232),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_SL g235 ( 
.A(n_231),
.B(n_232),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_238),
.B(n_239),
.Y(n_237)
);

OR2x2_ASAP7_75t_L g264 ( 
.A(n_238),
.B(n_239),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_243),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_242),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_241),
.B(n_242),
.C(n_243),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_252),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_248),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_245),
.B(n_248),
.C(n_252),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_255),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_254),
.B(n_255),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_263),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_257),
.A2(n_258),
.B1(n_261),
.B2(n_262),
.Y(n_256)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_257),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_257),
.B(n_262),
.C(n_263),
.Y(n_267)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_258),
.Y(n_262)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_267),
.B(n_268),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_267),
.B(n_268),
.Y(n_270)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_272),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_273),
.B(n_293),
.Y(n_272)
);

INVxp67_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_SL g274 ( 
.A(n_275),
.B(n_292),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_275),
.B(n_292),
.Y(n_293)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_276),
.B(n_277),
.Y(n_275)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_278),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_279),
.A2(n_280),
.B1(n_282),
.B2(n_283),
.Y(n_278)
);

CKINVDCx14_ASAP7_75t_R g279 ( 
.A(n_280),
.Y(n_279)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_284),
.A2(n_285),
.B1(n_286),
.B2(n_289),
.Y(n_283)
);

CKINVDCx16_ASAP7_75t_R g289 ( 
.A(n_284),
.Y(n_289)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

CKINVDCx14_ASAP7_75t_R g287 ( 
.A(n_288),
.Y(n_287)
);


endmodule