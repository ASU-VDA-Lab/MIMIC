module fake_jpeg_27813_n_65 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_65);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_65;

wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_23;
wire n_27;
wire n_55;
wire n_64;
wire n_22;
wire n_47;
wire n_51;
wire n_40;
wire n_20;
wire n_59;
wire n_48;
wire n_35;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_44;
wire n_24;
wire n_38;
wire n_26;
wire n_28;
wire n_36;
wire n_62;
wire n_25;
wire n_31;
wire n_56;
wire n_43;
wire n_37;
wire n_29;
wire n_50;
wire n_32;

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

AOI21xp33_ASAP7_75t_L g21 ( 
.A1(n_7),
.A2(n_12),
.B(n_11),
.Y(n_21)
);

INVx8_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_3),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_17),
.Y(n_26)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_19),
.Y(n_32)
);

BUFx10_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

BUFx4f_ASAP7_75t_SL g35 ( 
.A(n_6),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_6),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_15),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_22),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_38),
.B(n_40),
.Y(n_55)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_32),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_39),
.A2(n_44),
.B1(n_45),
.B2(n_47),
.Y(n_54)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_24),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_27),
.Y(n_41)
);

CKINVDCx16_ASAP7_75t_R g56 ( 
.A(n_41),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g42 ( 
.A1(n_21),
.A2(n_13),
.B1(n_16),
.B2(n_18),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_42),
.A2(n_43),
.B1(n_46),
.B2(n_48),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g43 ( 
.A1(n_25),
.A2(n_5),
.B1(n_1),
.B2(n_2),
.Y(n_43)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_20),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_37),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_L g46 ( 
.A1(n_30),
.A2(n_5),
.B1(n_34),
.B2(n_31),
.Y(n_46)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_33),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g49 ( 
.A(n_36),
.B(n_23),
.Y(n_49)
);

CKINVDCx12_ASAP7_75t_R g50 ( 
.A(n_26),
.Y(n_50)
);

HB1xp67_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_26),
.A2(n_23),
.B1(n_33),
.B2(n_29),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_55),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_57),
.A2(n_58),
.B1(n_53),
.B2(n_49),
.Y(n_59)
);

AOI21xp5_ASAP7_75t_L g58 ( 
.A1(n_53),
.A2(n_28),
.B(n_52),
.Y(n_58)
);

OAI321xp33_ASAP7_75t_L g60 ( 
.A1(n_59),
.A2(n_52),
.A3(n_46),
.B1(n_43),
.B2(n_50),
.C(n_54),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_60),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_61),
.Y(n_62)
);

OAI221xp5_ASAP7_75t_L g63 ( 
.A1(n_62),
.A2(n_41),
.B1(n_51),
.B2(n_56),
.C(n_59),
.Y(n_63)
);

INVxp67_ASAP7_75t_L g64 ( 
.A(n_63),
.Y(n_64)
);

XNOR2xp5_ASAP7_75t_L g65 ( 
.A(n_64),
.B(n_51),
.Y(n_65)
);


endmodule