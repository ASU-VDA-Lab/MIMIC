module real_jpeg_17287_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_425;
wire n_50;
wire n_409;
wire n_186;
wire n_137;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_366;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_432;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_368;
wire n_100;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

AOI21xp5_ASAP7_75t_L g18 ( 
.A1(n_0),
.A2(n_19),
.B(n_440),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g440 ( 
.A(n_0),
.B(n_441),
.Y(n_440)
);

AOI22xp5_ASAP7_75t_SL g41 ( 
.A1(n_1),
.A2(n_14),
.B1(n_42),
.B2(n_43),
.Y(n_41)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_1),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_1),
.B(n_140),
.Y(n_139)
);

AND2x2_ASAP7_75t_SL g156 ( 
.A(n_1),
.B(n_157),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_1),
.B(n_310),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_1),
.B(n_329),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_SL g353 ( 
.A(n_1),
.B(n_354),
.Y(n_353)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_2),
.Y(n_60)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_2),
.Y(n_133)
);

BUFx3_ASAP7_75t_L g158 ( 
.A(n_2),
.Y(n_158)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_2),
.Y(n_436)
);

AND2x2_ASAP7_75t_L g36 ( 
.A(n_3),
.B(n_37),
.Y(n_36)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_3),
.B(n_81),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_3),
.B(n_111),
.Y(n_110)
);

AND2x2_ASAP7_75t_L g120 ( 
.A(n_3),
.B(n_121),
.Y(n_120)
);

AND2x2_ASAP7_75t_L g135 ( 
.A(n_3),
.B(n_136),
.Y(n_135)
);

AND2x2_ASAP7_75t_L g194 ( 
.A(n_3),
.B(n_195),
.Y(n_194)
);

AND2x2_ASAP7_75t_L g428 ( 
.A(n_3),
.B(n_429),
.Y(n_428)
);

AND2x2_ASAP7_75t_SL g56 ( 
.A(n_4),
.B(n_57),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_4),
.B(n_70),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_4),
.B(n_107),
.Y(n_106)
);

AND2x2_ASAP7_75t_SL g159 ( 
.A(n_4),
.B(n_160),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_4),
.B(n_191),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_4),
.B(n_261),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_4),
.B(n_267),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_4),
.B(n_154),
.Y(n_326)
);

BUFx5_ASAP7_75t_L g68 ( 
.A(n_5),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_5),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_5),
.Y(n_166)
);

BUFx5_ASAP7_75t_L g264 ( 
.A(n_5),
.Y(n_264)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_5),
.Y(n_312)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_6),
.B(n_74),
.Y(n_73)
);

NAND2x1p5_ASAP7_75t_L g94 ( 
.A(n_6),
.B(n_70),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g124 ( 
.A(n_6),
.B(n_125),
.Y(n_124)
);

AND2x2_ASAP7_75t_SL g129 ( 
.A(n_6),
.B(n_130),
.Y(n_129)
);

AND2x2_ASAP7_75t_L g163 ( 
.A(n_6),
.B(n_164),
.Y(n_163)
);

AND2x2_ASAP7_75t_L g201 ( 
.A(n_6),
.B(n_202),
.Y(n_201)
);

AND2x2_ASAP7_75t_L g206 ( 
.A(n_6),
.B(n_207),
.Y(n_206)
);

AND2x2_ASAP7_75t_L g413 ( 
.A(n_6),
.B(n_414),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_7),
.B(n_77),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g242 ( 
.A(n_7),
.B(n_243),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_7),
.B(n_248),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_7),
.B(n_307),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_7),
.B(n_341),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_SL g361 ( 
.A(n_7),
.B(n_362),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_SL g367 ( 
.A(n_7),
.B(n_368),
.Y(n_367)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_8),
.Y(n_38)
);

BUFx5_ASAP7_75t_L g125 ( 
.A(n_8),
.Y(n_125)
);

BUFx5_ASAP7_75t_L g154 ( 
.A(n_8),
.Y(n_154)
);

AND2x2_ASAP7_75t_L g50 ( 
.A(n_9),
.B(n_51),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_9),
.B(n_68),
.Y(n_67)
);

AND2x2_ASAP7_75t_L g102 ( 
.A(n_9),
.B(n_103),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_9),
.B(n_153),
.Y(n_152)
);

AND2x2_ASAP7_75t_L g216 ( 
.A(n_9),
.B(n_217),
.Y(n_216)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_9),
.Y(n_423)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_10),
.Y(n_75)
);

BUFx3_ASAP7_75t_L g104 ( 
.A(n_10),
.Y(n_104)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_10),
.Y(n_138)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_10),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g241 ( 
.A(n_10),
.Y(n_241)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_11),
.Y(n_441)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_12),
.Y(n_64)
);

INVx6_ASAP7_75t_L g109 ( 
.A(n_12),
.Y(n_109)
);

BUFx5_ASAP7_75t_L g142 ( 
.A(n_12),
.Y(n_142)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_12),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g28 ( 
.A(n_13),
.B(n_29),
.Y(n_28)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_13),
.B(n_62),
.Y(n_61)
);

AND2x2_ASAP7_75t_L g236 ( 
.A(n_13),
.B(n_237),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_13),
.B(n_251),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_13),
.B(n_302),
.Y(n_301)
);

AND2x2_ASAP7_75t_L g343 ( 
.A(n_13),
.B(n_164),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_13),
.B(n_352),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_SL g370 ( 
.A(n_13),
.B(n_354),
.Y(n_370)
);

AND2x2_ASAP7_75t_L g32 ( 
.A(n_14),
.B(n_33),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_14),
.B(n_93),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g218 ( 
.A(n_14),
.B(n_160),
.Y(n_218)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_14),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g432 ( 
.A(n_14),
.B(n_433),
.Y(n_432)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_15),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_15),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_16),
.Y(n_55)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_16),
.Y(n_123)
);

BUFx4f_ASAP7_75t_L g209 ( 
.A(n_16),
.Y(n_209)
);

BUFx8_ASAP7_75t_L g29 ( 
.A(n_17),
.Y(n_29)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_17),
.Y(n_79)
);

BUFx5_ASAP7_75t_L g414 ( 
.A(n_17),
.Y(n_414)
);

XOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_397),
.Y(n_19)
);

OAI21xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_222),
.B(n_395),
.Y(n_20)
);

INVxp67_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_175),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g396 ( 
.A(n_23),
.B(n_175),
.Y(n_396)
);

MAJIxp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_99),
.C(n_145),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_SL g390 ( 
.A1(n_24),
.A2(n_25),
.B1(n_100),
.B2(n_391),
.Y(n_390)
);

INVx1_ASAP7_75t_SL g24 ( 
.A(n_25),
.Y(n_24)
);

XNOR2xp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_65),
.Y(n_25)
);

INVxp33_ASAP7_75t_SL g177 ( 
.A(n_26),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_40),
.C(n_48),
.Y(n_26)
);

XNOR2xp5_ASAP7_75t_L g384 ( 
.A(n_27),
.B(n_385),
.Y(n_384)
);

XNOR2xp5_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_30),
.Y(n_27)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_28),
.B(n_32),
.C(n_36),
.Y(n_88)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_29),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g30 ( 
.A1(n_31),
.A2(n_32),
.B1(n_36),
.B2(n_39),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_35),
.Y(n_268)
);

INVx1_ASAP7_75t_SL g39 ( 
.A(n_36),
.Y(n_39)
);

AND2x2_ASAP7_75t_L g256 ( 
.A(n_36),
.B(n_206),
.Y(n_256)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_37),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g289 ( 
.A(n_37),
.Y(n_289)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_39),
.B(n_206),
.Y(n_258)
);

AOI22xp33_ASAP7_75t_SL g385 ( 
.A1(n_40),
.A2(n_41),
.B1(n_48),
.B2(n_49),
.Y(n_385)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

AOI21xp5_ASAP7_75t_L g280 ( 
.A1(n_41),
.A2(n_281),
.B(n_286),
.Y(n_280)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g244 ( 
.A(n_46),
.Y(n_244)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

BUFx5_ASAP7_75t_L g195 ( 
.A(n_47),
.Y(n_195)
);

BUFx6f_ASAP7_75t_L g285 ( 
.A(n_47),
.Y(n_285)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

MAJIxp5_ASAP7_75t_L g49 ( 
.A(n_50),
.B(n_56),
.C(n_61),
.Y(n_49)
);

XNOR2xp5_ASAP7_75t_L g148 ( 
.A(n_50),
.B(n_61),
.Y(n_148)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx4_ASAP7_75t_L g330 ( 
.A(n_55),
.Y(n_330)
);

BUFx6f_ASAP7_75t_L g352 ( 
.A(n_55),
.Y(n_352)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_56),
.B(n_148),
.Y(n_147)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_60),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g217 ( 
.A(n_60),
.Y(n_217)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx2_ASAP7_75t_L g430 ( 
.A(n_64),
.Y(n_430)
);

AOI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_66),
.A2(n_87),
.B1(n_97),
.B2(n_98),
.Y(n_65)
);

INVxp67_ASAP7_75t_SL g97 ( 
.A(n_66),
.Y(n_97)
);

HB1xp67_ASAP7_75t_L g178 ( 
.A(n_66),
.Y(n_178)
);

A2O1A1Ixp33_ASAP7_75t_L g66 ( 
.A1(n_67),
.A2(n_69),
.B(n_72),
.C(n_84),
.Y(n_66)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_67),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_67),
.A2(n_69),
.B1(n_85),
.B2(n_86),
.Y(n_174)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_69),
.Y(n_86)
);

INVx6_ASAP7_75t_L g424 ( 
.A(n_70),
.Y(n_424)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx3_ASAP7_75t_L g254 ( 
.A(n_71),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g173 ( 
.A(n_72),
.B(n_174),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_73),
.B(n_76),
.C(n_80),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_73),
.A2(n_80),
.B1(n_292),
.B2(n_293),
.Y(n_291)
);

INVx1_ASAP7_75t_SL g292 ( 
.A(n_73),
.Y(n_292)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_76),
.B(n_291),
.Y(n_290)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g192 ( 
.A(n_79),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_80),
.B(n_214),
.Y(n_213)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_80),
.Y(n_293)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx6_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_83),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_86),
.Y(n_84)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_87),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_88),
.A2(n_89),
.B1(n_90),
.B2(n_96),
.Y(n_87)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_88),
.Y(n_96)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_91),
.A2(n_92),
.B1(n_94),
.B2(n_95),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_91),
.B(n_95),
.C(n_96),
.Y(n_186)
);

INVx1_ASAP7_75t_SL g91 ( 
.A(n_92),
.Y(n_91)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_94),
.Y(n_95)
);

HB1xp67_ASAP7_75t_L g179 ( 
.A(n_98),
.Y(n_179)
);

HB1xp67_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_100),
.Y(n_391)
);

XNOR2x1_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_113),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_101),
.B(n_127),
.C(n_143),
.Y(n_183)
);

XNOR2x2_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_105),
.Y(n_101)
);

MAJx2_ASAP7_75t_L g196 ( 
.A(n_102),
.B(n_106),
.C(n_110),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

XNOR2xp5_ASAP7_75t_SL g105 ( 
.A(n_106),
.B(n_110),
.Y(n_105)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx4_ASAP7_75t_L g248 ( 
.A(n_109),
.Y(n_248)
);

HB1xp67_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_112),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_114),
.A2(n_127),
.B1(n_143),
.B2(n_144),
.Y(n_113)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_114),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_118),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_115),
.B(n_119),
.C(n_126),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_117),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_116),
.B(n_240),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_116),
.B(n_282),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_119),
.A2(n_120),
.B1(n_124),
.B2(n_126),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_119),
.A2(n_120),
.B1(n_151),
.B2(n_152),
.Y(n_234)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_120),
.B(n_151),
.Y(n_150)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_124),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_124),
.A2(n_126),
.B1(n_206),
.B2(n_210),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g332 ( 
.A(n_124),
.B(n_266),
.Y(n_332)
);

INVx2_ASAP7_75t_L g355 ( 
.A(n_125),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_126),
.B(n_266),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g415 ( 
.A(n_126),
.B(n_201),
.C(n_206),
.Y(n_415)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_127),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_134),
.C(n_139),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_128),
.A2(n_129),
.B1(n_139),
.B2(n_171),
.Y(n_170)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_134),
.A2(n_135),
.B1(n_169),
.B2(n_170),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_SL g431 ( 
.A1(n_134),
.A2(n_135),
.B1(n_432),
.B2(n_437),
.Y(n_431)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

BUFx3_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx2_ASAP7_75t_L g342 ( 
.A(n_138),
.Y(n_342)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_139),
.Y(n_171)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g389 ( 
.A(n_145),
.B(n_390),
.Y(n_389)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_167),
.C(n_172),
.Y(n_145)
);

XOR2xp5_ASAP7_75t_L g381 ( 
.A(n_146),
.B(n_382),
.Y(n_381)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_149),
.C(n_155),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_SL g272 ( 
.A(n_147),
.B(n_273),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_149),
.A2(n_150),
.B1(n_155),
.B2(n_274),
.Y(n_273)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

BUFx12f_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_155),
.Y(n_274)
);

MAJx2_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_159),
.C(n_163),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_156),
.A2(n_163),
.B1(n_231),
.B2(n_232),
.Y(n_230)
);

CKINVDCx14_ASAP7_75t_R g231 ( 
.A(n_156),
.Y(n_231)
);

BUFx3_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_SL g229 ( 
.A(n_159),
.B(n_230),
.Y(n_229)
);

INVx6_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

INVx1_ASAP7_75t_SL g232 ( 
.A(n_163),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g421 ( 
.A1(n_163),
.A2(n_206),
.B1(n_210),
.B2(n_232),
.Y(n_421)
);

INVx4_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

INVx8_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g382 ( 
.A(n_168),
.B(n_173),
.Y(n_382)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_180),
.Y(n_175)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_176),
.Y(n_401)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_178),
.C(n_179),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_181),
.A2(n_199),
.B1(n_220),
.B2(n_221),
.Y(n_180)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_181),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_182),
.A2(n_183),
.B1(n_184),
.B2(n_198),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g403 ( 
.A(n_182),
.B(n_185),
.C(n_404),
.Y(n_403)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_184),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_185),
.A2(n_186),
.B1(n_187),
.B2(n_197),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_187),
.Y(n_197)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_187),
.Y(n_404)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_188),
.B(n_196),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_189),
.A2(n_190),
.B1(n_193),
.B2(n_194),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

MAJx2_ASAP7_75t_L g410 ( 
.A(n_190),
.B(n_193),
.C(n_196),
.Y(n_410)
);

INVx4_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

INVx2_ASAP7_75t_SL g193 ( 
.A(n_194),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g412 ( 
.A(n_194),
.B(n_413),
.Y(n_412)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_199),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g400 ( 
.A(n_199),
.B(n_220),
.C(n_401),
.Y(n_400)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_211),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g408 ( 
.A(n_200),
.B(n_212),
.C(n_213),
.Y(n_408)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_205),
.Y(n_200)
);

INVx3_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

BUFx3_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_206),
.Y(n_210)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_213),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_215),
.A2(n_216),
.B1(n_218),
.B2(n_219),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g426 ( 
.A(n_215),
.B(n_219),
.C(n_293),
.Y(n_426)
);

CKINVDCx16_ASAP7_75t_R g215 ( 
.A(n_216),
.Y(n_215)
);

INVx5_ASAP7_75t_L g308 ( 
.A(n_217),
.Y(n_308)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_218),
.Y(n_219)
);

AOI21xp5_ASAP7_75t_L g222 ( 
.A1(n_223),
.A2(n_377),
.B(n_392),
.Y(n_222)
);

HB1xp67_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_L g224 ( 
.A1(n_225),
.A2(n_294),
.B(n_376),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_269),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g376 ( 
.A(n_226),
.B(n_269),
.Y(n_376)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_245),
.C(n_257),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_227),
.A2(n_228),
.B1(n_316),
.B2(n_317),
.Y(n_315)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_SL g228 ( 
.A(n_229),
.B(n_233),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_229),
.B(n_234),
.C(n_235),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_235),
.Y(n_233)
);

MAJx2_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_239),
.C(n_242),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_236),
.B(n_242),
.Y(n_314)
);

INVx3_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_239),
.B(n_314),
.Y(n_313)
);

INVx4_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

INVx4_ASAP7_75t_L g305 ( 
.A(n_241),
.Y(n_305)
);

INVx4_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_SL g317 ( 
.A(n_245),
.B(n_257),
.Y(n_317)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_256),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_247),
.A2(n_249),
.B1(n_250),
.B2(n_255),
.Y(n_246)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_247),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_249),
.B(n_255),
.C(n_256),
.Y(n_278)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_259),
.C(n_265),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_258),
.A2(n_259),
.B1(n_260),
.B2(n_299),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_258),
.Y(n_299)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

BUFx2_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

INVx2_ASAP7_75t_L g364 ( 
.A(n_263),
.Y(n_364)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_SL g297 ( 
.A(n_265),
.B(n_298),
.Y(n_297)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_267),
.Y(n_369)
);

INVx5_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_270),
.B(n_277),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_271),
.A2(n_272),
.B1(n_275),
.B2(n_276),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g379 ( 
.A(n_271),
.B(n_276),
.C(n_277),
.Y(n_379)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_SL g277 ( 
.A(n_278),
.B(n_279),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g386 ( 
.A(n_278),
.B(n_280),
.C(n_290),
.Y(n_386)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_280),
.B(n_290),
.Y(n_279)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_287),
.B(n_288),
.Y(n_286)
);

INVx2_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

AOI21x1_ASAP7_75t_SL g294 ( 
.A1(n_295),
.A2(n_318),
.B(n_375),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_296),
.B(n_315),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_SL g375 ( 
.A(n_296),
.B(n_315),
.Y(n_375)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_297),
.B(n_300),
.C(n_313),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g333 ( 
.A(n_297),
.B(n_334),
.Y(n_333)
);

XNOR2xp5_ASAP7_75t_L g334 ( 
.A(n_300),
.B(n_313),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_301),
.B(n_306),
.C(n_309),
.Y(n_300)
);

XOR2xp5_ASAP7_75t_L g322 ( 
.A(n_301),
.B(n_323),
.Y(n_322)
);

INVx1_ASAP7_75t_SL g302 ( 
.A(n_303),
.Y(n_302)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g323 ( 
.A(n_306),
.B(n_309),
.Y(n_323)
);

INVx5_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

INVx4_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

BUFx3_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

OAI21x1_ASAP7_75t_L g318 ( 
.A1(n_319),
.A2(n_335),
.B(n_374),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_320),
.B(n_333),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_SL g374 ( 
.A(n_320),
.B(n_333),
.Y(n_374)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_321),
.B(n_324),
.C(n_331),
.Y(n_320)
);

AOI22xp33_ASAP7_75t_SL g344 ( 
.A1(n_321),
.A2(n_322),
.B1(n_345),
.B2(n_347),
.Y(n_344)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_L g345 ( 
.A1(n_324),
.A2(n_331),
.B1(n_332),
.B2(n_346),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_324),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_325),
.B(n_327),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_SL g338 ( 
.A1(n_325),
.A2(n_326),
.B1(n_327),
.B2(n_328),
.Y(n_338)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_332),
.Y(n_331)
);

AOI21xp5_ASAP7_75t_L g335 ( 
.A1(n_336),
.A2(n_348),
.B(n_373),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_337),
.B(n_344),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_SL g373 ( 
.A(n_337),
.B(n_344),
.Y(n_373)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_338),
.B(n_339),
.C(n_343),
.Y(n_337)
);

XOR2xp5_ASAP7_75t_L g356 ( 
.A(n_338),
.B(n_357),
.Y(n_356)
);

OAI22xp5_ASAP7_75t_SL g357 ( 
.A1(n_339),
.A2(n_340),
.B1(n_343),
.B2(n_358),
.Y(n_357)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_340),
.Y(n_339)
);

HB1xp67_ASAP7_75t_L g341 ( 
.A(n_342),
.Y(n_341)
);

CKINVDCx16_ASAP7_75t_R g358 ( 
.A(n_343),
.Y(n_358)
);

INVxp67_ASAP7_75t_SL g347 ( 
.A(n_345),
.Y(n_347)
);

OAI21xp5_ASAP7_75t_SL g348 ( 
.A1(n_349),
.A2(n_359),
.B(n_372),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_350),
.B(n_356),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_SL g372 ( 
.A(n_350),
.B(n_356),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_L g350 ( 
.A(n_351),
.B(n_353),
.Y(n_350)
);

XNOR2xp5_ASAP7_75t_L g365 ( 
.A(n_351),
.B(n_353),
.Y(n_365)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_355),
.Y(n_354)
);

AOI21xp5_ASAP7_75t_L g359 ( 
.A1(n_360),
.A2(n_366),
.B(n_371),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_361),
.B(n_365),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_SL g371 ( 
.A(n_361),
.B(n_365),
.Y(n_371)
);

INVx2_ASAP7_75t_L g362 ( 
.A(n_363),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_364),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_L g366 ( 
.A(n_367),
.B(n_370),
.Y(n_366)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_369),
.Y(n_368)
);

NOR2x1_ASAP7_75t_L g377 ( 
.A(n_378),
.B(n_387),
.Y(n_377)
);

NOR2x1_ASAP7_75t_L g378 ( 
.A(n_379),
.B(n_380),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_379),
.B(n_380),
.Y(n_393)
);

XNOR2xp5_ASAP7_75t_L g380 ( 
.A(n_381),
.B(n_383),
.Y(n_380)
);

MAJIxp5_ASAP7_75t_L g388 ( 
.A(n_381),
.B(n_384),
.C(n_386),
.Y(n_388)
);

XNOR2xp5_ASAP7_75t_L g383 ( 
.A(n_384),
.B(n_386),
.Y(n_383)
);

OAI21x1_ASAP7_75t_SL g392 ( 
.A1(n_387),
.A2(n_393),
.B(n_394),
.Y(n_392)
);

AND2x2_ASAP7_75t_L g387 ( 
.A(n_388),
.B(n_389),
.Y(n_387)
);

OR2x2_ASAP7_75t_L g394 ( 
.A(n_388),
.B(n_389),
.Y(n_394)
);

INVxp67_ASAP7_75t_SL g395 ( 
.A(n_396),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_L g397 ( 
.A(n_398),
.B(n_438),
.Y(n_397)
);

HB1xp67_ASAP7_75t_L g398 ( 
.A(n_399),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_L g399 ( 
.A(n_400),
.B(n_402),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_400),
.B(n_402),
.Y(n_439)
);

XNOR2xp5_ASAP7_75t_L g402 ( 
.A(n_403),
.B(n_405),
.Y(n_402)
);

XNOR2xp5_ASAP7_75t_L g405 ( 
.A(n_406),
.B(n_419),
.Y(n_405)
);

AOI22xp5_ASAP7_75t_L g406 ( 
.A1(n_407),
.A2(n_408),
.B1(n_409),
.B2(n_418),
.Y(n_406)
);

INVx1_ASAP7_75t_SL g407 ( 
.A(n_408),
.Y(n_407)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_409),
.Y(n_418)
);

XNOR2xp5_ASAP7_75t_SL g409 ( 
.A(n_410),
.B(n_411),
.Y(n_409)
);

AO22x1_ASAP7_75t_SL g411 ( 
.A1(n_412),
.A2(n_415),
.B1(n_416),
.B2(n_417),
.Y(n_411)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_412),
.Y(n_416)
);

INVx1_ASAP7_75t_SL g417 ( 
.A(n_415),
.Y(n_417)
);

XOR2xp5_ASAP7_75t_L g419 ( 
.A(n_420),
.B(n_425),
.Y(n_419)
);

XNOR2xp5_ASAP7_75t_SL g420 ( 
.A(n_421),
.B(n_422),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_L g422 ( 
.A(n_423),
.B(n_424),
.Y(n_422)
);

XNOR2xp5_ASAP7_75t_L g425 ( 
.A(n_426),
.B(n_427),
.Y(n_425)
);

XNOR2xp5_ASAP7_75t_L g427 ( 
.A(n_428),
.B(n_431),
.Y(n_427)
);

INVx1_ASAP7_75t_SL g429 ( 
.A(n_430),
.Y(n_429)
);

INVx1_ASAP7_75t_SL g437 ( 
.A(n_432),
.Y(n_437)
);

BUFx2_ASAP7_75t_L g433 ( 
.A(n_434),
.Y(n_433)
);

INVx3_ASAP7_75t_L g434 ( 
.A(n_435),
.Y(n_434)
);

BUFx6f_ASAP7_75t_L g435 ( 
.A(n_436),
.Y(n_435)
);

INVxp33_ASAP7_75t_L g438 ( 
.A(n_439),
.Y(n_438)
);


endmodule