module real_jpeg_22515_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_323, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_323;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_215;
wire n_176;
wire n_312;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

OAI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_0),
.A2(n_26),
.B1(n_35),
.B2(n_95),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_0),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_L g149 ( 
.A1(n_0),
.A2(n_47),
.B1(n_50),
.B2(n_95),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_0),
.A2(n_64),
.B1(n_65),
.B2(n_95),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_L g203 ( 
.A1(n_0),
.A2(n_32),
.B1(n_33),
.B2(n_95),
.Y(n_203)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_1),
.A2(n_26),
.B1(n_35),
.B2(n_132),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_1),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_SL g165 ( 
.A1(n_1),
.A2(n_64),
.B1(n_65),
.B2(n_132),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_L g199 ( 
.A1(n_1),
.A2(n_47),
.B1(n_50),
.B2(n_132),
.Y(n_199)
);

AOI22xp33_ASAP7_75t_SL g256 ( 
.A1(n_1),
.A2(n_32),
.B1(n_33),
.B2(n_132),
.Y(n_256)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_2),
.A2(n_32),
.B1(n_33),
.B2(n_56),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_2),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_2),
.A2(n_47),
.B1(n_50),
.B2(n_56),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_2),
.A2(n_56),
.B1(n_64),
.B2(n_65),
.Y(n_124)
);

A2O1A1O1Ixp25_ASAP7_75t_L g146 ( 
.A1(n_3),
.A2(n_50),
.B(n_60),
.C(n_147),
.D(n_148),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_3),
.B(n_50),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_3),
.B(n_46),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_3),
.Y(n_182)
);

OAI21xp33_ASAP7_75t_L g187 ( 
.A1(n_3),
.A2(n_83),
.B(n_166),
.Y(n_187)
);

A2O1A1O1Ixp25_ASAP7_75t_L g200 ( 
.A1(n_3),
.A2(n_32),
.B(n_43),
.C(n_201),
.D(n_202),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_3),
.B(n_32),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_3),
.B(n_134),
.Y(n_227)
);

AOI21xp33_ASAP7_75t_L g243 ( 
.A1(n_3),
.A2(n_31),
.B(n_33),
.Y(n_243)
);

OAI22xp33_ASAP7_75t_SL g259 ( 
.A1(n_3),
.A2(n_26),
.B1(n_35),
.B2(n_182),
.Y(n_259)
);

AOI22xp33_ASAP7_75t_SL g34 ( 
.A1(n_4),
.A2(n_26),
.B1(n_35),
.B2(n_36),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_4),
.Y(n_36)
);

OAI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_4),
.A2(n_32),
.B1(n_33),
.B2(n_36),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_L g212 ( 
.A1(n_4),
.A2(n_36),
.B1(n_64),
.B2(n_65),
.Y(n_212)
);

AOI22xp33_ASAP7_75t_L g253 ( 
.A1(n_4),
.A2(n_36),
.B1(n_47),
.B2(n_50),
.Y(n_253)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_5),
.A2(n_47),
.B1(n_50),
.B2(n_69),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_5),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_5),
.A2(n_64),
.B1(n_65),
.B2(n_69),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_5),
.A2(n_32),
.B1(n_33),
.B2(n_69),
.Y(n_106)
);

BUFx16f_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

INVx8_ASAP7_75t_L g84 ( 
.A(n_7),
.Y(n_84)
);

INVx6_ASAP7_75t_L g87 ( 
.A(n_7),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_7),
.B(n_167),
.Y(n_166)
);

BUFx12_ASAP7_75t_L g64 ( 
.A(n_8),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_9),
.A2(n_47),
.B1(n_50),
.B2(n_161),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_9),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_SL g173 ( 
.A1(n_9),
.A2(n_64),
.B1(n_65),
.B2(n_161),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_SL g221 ( 
.A1(n_9),
.A2(n_32),
.B1(n_33),
.B2(n_161),
.Y(n_221)
);

AOI22xp33_ASAP7_75t_SL g268 ( 
.A1(n_9),
.A2(n_26),
.B1(n_35),
.B2(n_161),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_10),
.A2(n_32),
.B1(n_33),
.B2(n_53),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_10),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_L g90 ( 
.A1(n_10),
.A2(n_47),
.B1(n_50),
.B2(n_53),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_10),
.A2(n_26),
.B1(n_35),
.B2(n_53),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g246 ( 
.A1(n_10),
.A2(n_53),
.B1(n_64),
.B2(n_65),
.Y(n_246)
);

BUFx12_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_SL g37 ( 
.A1(n_12),
.A2(n_26),
.B1(n_35),
.B2(n_38),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_12),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_12),
.A2(n_32),
.B1(n_33),
.B2(n_38),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_12),
.A2(n_38),
.B1(n_47),
.B2(n_50),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g226 ( 
.A1(n_12),
.A2(n_38),
.B1(n_64),
.B2(n_65),
.Y(n_226)
);

INVx13_ASAP7_75t_L g44 ( 
.A(n_13),
.Y(n_44)
);

INVx13_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

INVx11_ASAP7_75t_L g61 ( 
.A(n_15),
.Y(n_61)
);

INVx11_ASAP7_75t_SL g48 ( 
.A(n_16),
.Y(n_48)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_111),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_110),
.Y(n_18)
);

INVxp67_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_97),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_21),
.B(n_97),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_71),
.C(n_79),
.Y(n_21)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_22),
.A2(n_71),
.B1(n_72),
.B2(n_137),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_22),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_24),
.B1(n_39),
.B2(n_40),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_23),
.A2(n_24),
.B1(n_99),
.B2(n_100),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_24),
.Y(n_23)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_24),
.B(n_57),
.C(n_70),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g24 ( 
.A1(n_25),
.A2(n_30),
.B1(n_34),
.B2(n_37),
.Y(n_24)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_25),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_25),
.A2(n_30),
.B1(n_37),
.B2(n_102),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_SL g130 ( 
.A1(n_25),
.A2(n_131),
.B(n_133),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_25),
.A2(n_30),
.B1(n_131),
.B2(n_268),
.Y(n_288)
);

A2O1A1Ixp33_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_28),
.B(n_29),
.C(n_30),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_26),
.B(n_28),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_26),
.Y(n_35)
);

A2O1A1Ixp33_ASAP7_75t_L g242 ( 
.A1(n_26),
.A2(n_28),
.B(n_182),
.C(n_243),
.Y(n_242)
);

BUFx2_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g30 ( 
.A1(n_28),
.A2(n_31),
.B1(n_32),
.B2(n_33),
.Y(n_30)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_28),
.Y(n_31)
);

OAI21xp5_ASAP7_75t_L g92 ( 
.A1(n_30),
.A2(n_34),
.B(n_93),
.Y(n_92)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_30),
.Y(n_134)
);

OAI21xp33_ASAP7_75t_L g267 ( 
.A1(n_30),
.A2(n_93),
.B(n_268),
.Y(n_267)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

O2A1O1Ixp33_ASAP7_75t_SL g43 ( 
.A1(n_33),
.A2(n_44),
.B(n_45),
.C(n_46),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_33),
.B(n_44),
.Y(n_45)
);

CKINVDCx14_ASAP7_75t_R g39 ( 
.A(n_40),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g40 ( 
.A1(n_41),
.A2(n_57),
.B1(n_58),
.B2(n_70),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_41),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g41 ( 
.A1(n_42),
.A2(n_51),
.B1(n_54),
.B2(n_55),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_42),
.A2(n_54),
.B1(n_55),
.B2(n_106),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_42),
.A2(n_54),
.B1(n_221),
.B2(n_256),
.Y(n_255)
);

OAI21xp5_ASAP7_75t_L g270 ( 
.A1(n_42),
.A2(n_256),
.B(n_271),
.Y(n_270)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_43),
.A2(n_46),
.B1(n_52),
.B2(n_74),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_43),
.A2(n_46),
.B1(n_74),
.B2(n_128),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_43),
.B(n_223),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_L g46 ( 
.A1(n_44),
.A2(n_47),
.B1(n_49),
.B2(n_50),
.Y(n_46)
);

INVx11_ASAP7_75t_L g49 ( 
.A(n_44),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_45),
.Y(n_209)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_46),
.Y(n_54)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_47),
.Y(n_50)
);

O2A1O1Ixp33_ASAP7_75t_L g60 ( 
.A1(n_47),
.A2(n_61),
.B(n_62),
.C(n_63),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_47),
.B(n_61),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_47),
.B(n_49),
.Y(n_208)
);

INVx11_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_50),
.A2(n_201),
.B1(n_208),
.B2(n_209),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_52),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_54),
.B(n_203),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_L g220 ( 
.A1(n_54),
.A2(n_221),
.B(n_222),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_L g285 ( 
.A1(n_54),
.A2(n_222),
.B(n_286),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_57),
.A2(n_58),
.B1(n_105),
.B2(n_107),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_58),
.Y(n_57)
);

AOI21xp5_ASAP7_75t_SL g58 ( 
.A1(n_59),
.A2(n_67),
.B(n_68),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_59),
.A2(n_67),
.B1(n_77),
.B2(n_90),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_59),
.A2(n_67),
.B1(n_90),
.B2(n_126),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_59),
.A2(n_67),
.B1(n_160),
.B2(n_199),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_SL g233 ( 
.A1(n_59),
.A2(n_199),
.B(n_234),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_L g276 ( 
.A1(n_59),
.A2(n_67),
.B1(n_126),
.B2(n_253),
.Y(n_276)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_60),
.A2(n_63),
.B1(n_76),
.B2(n_78),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_60),
.B(n_163),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_61),
.A2(n_64),
.B1(n_65),
.B2(n_66),
.Y(n_63)
);

CKINVDCx9p33_ASAP7_75t_R g66 ( 
.A(n_61),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g152 ( 
.A(n_61),
.B(n_65),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_62),
.A2(n_64),
.B1(n_152),
.B2(n_153),
.Y(n_151)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_63),
.Y(n_67)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_64),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_64),
.B(n_84),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g188 ( 
.A(n_65),
.B(n_189),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_67),
.B(n_149),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_L g159 ( 
.A1(n_67),
.A2(n_160),
.B(n_162),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_SL g181 ( 
.A(n_67),
.B(n_182),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_L g252 ( 
.A1(n_67),
.A2(n_162),
.B(n_253),
.Y(n_252)
);

INVxp67_ASAP7_75t_L g78 ( 
.A(n_68),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_72),
.Y(n_71)
);

OAI21xp5_ASAP7_75t_L g119 ( 
.A1(n_72),
.A2(n_73),
.B(n_75),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_73),
.B(n_75),
.Y(n_72)
);

INVxp67_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

XNOR2xp5_ASAP7_75t_L g135 ( 
.A(n_79),
.B(n_136),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_L g79 ( 
.A1(n_80),
.A2(n_91),
.B(n_92),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_80),
.A2(n_81),
.B1(n_115),
.B2(n_117),
.Y(n_114)
);

CKINVDCx16_ASAP7_75t_R g80 ( 
.A(n_81),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_82),
.B(n_89),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_82),
.Y(n_91)
);

AOI22x1_ASAP7_75t_SL g115 ( 
.A1(n_82),
.A2(n_91),
.B1(n_92),
.B2(n_116),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g302 ( 
.A1(n_82),
.A2(n_89),
.B1(n_91),
.B2(n_303),
.Y(n_302)
);

AOI21xp5_ASAP7_75t_L g82 ( 
.A1(n_83),
.A2(n_85),
.B(n_88),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_83),
.A2(n_84),
.B1(n_88),
.B2(n_124),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_SL g164 ( 
.A1(n_83),
.A2(n_165),
.B(n_166),
.Y(n_164)
);

INVxp67_ASAP7_75t_L g174 ( 
.A(n_83),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_83),
.B(n_168),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_83),
.A2(n_84),
.B1(n_212),
.B2(n_226),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_83),
.A2(n_87),
.B1(n_226),
.B2(n_246),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_L g275 ( 
.A1(n_83),
.A2(n_85),
.B1(n_124),
.B2(n_246),
.Y(n_275)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_84),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_L g183 ( 
.A1(n_84),
.A2(n_173),
.B(n_184),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_84),
.B(n_182),
.Y(n_189)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

AOI21xp5_ASAP7_75t_L g210 ( 
.A1(n_86),
.A2(n_185),
.B(n_211),
.Y(n_210)
);

INVx5_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_89),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_92),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_96),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_94),
.B(n_134),
.Y(n_133)
);

AOI21xp5_ASAP7_75t_L g258 ( 
.A1(n_96),
.A2(n_259),
.B(n_260),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_109),
.Y(n_97)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_101),
.A2(n_103),
.B1(n_104),
.B2(n_108),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_101),
.Y(n_108)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_105),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_L g111 ( 
.A1(n_112),
.A2(n_138),
.B(n_321),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_135),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g321 ( 
.A(n_113),
.B(n_135),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_118),
.C(n_120),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g307 ( 
.A1(n_114),
.A2(n_118),
.B1(n_119),
.B2(n_308),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_114),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_115),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_119),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_SL g305 ( 
.A1(n_120),
.A2(n_121),
.B1(n_306),
.B2(n_307),
.Y(n_305)
);

CKINVDCx14_ASAP7_75t_R g120 ( 
.A(n_121),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_127),
.C(n_129),
.Y(n_121)
);

XOR2xp5_ASAP7_75t_L g299 ( 
.A(n_122),
.B(n_300),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_125),
.Y(n_122)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_123),
.B(n_125),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_L g300 ( 
.A1(n_127),
.A2(n_129),
.B1(n_130),
.B2(n_301),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_127),
.Y(n_301)
);

CKINVDCx16_ASAP7_75t_R g286 ( 
.A(n_128),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_130),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_133),
.Y(n_260)
);

AOI321xp33_ASAP7_75t_L g138 ( 
.A1(n_139),
.A2(n_296),
.A3(n_309),
.B1(n_315),
.B2(n_320),
.C(n_323),
.Y(n_138)
);

NOR3xp33_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_262),
.C(n_292),
.Y(n_139)
);

AOI21xp5_ASAP7_75t_L g140 ( 
.A1(n_141),
.A2(n_236),
.B(n_261),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_SL g141 ( 
.A1(n_142),
.A2(n_215),
.B(n_235),
.Y(n_141)
);

AOI21xp5_ASAP7_75t_L g142 ( 
.A1(n_143),
.A2(n_193),
.B(n_214),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_SL g143 ( 
.A1(n_144),
.A2(n_169),
.B(n_192),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_154),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_145),
.B(n_154),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_SL g145 ( 
.A(n_146),
.B(n_150),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_146),
.A2(n_150),
.B1(n_151),
.B2(n_178),
.Y(n_177)
);

CKINVDCx14_ASAP7_75t_R g178 ( 
.A(n_146),
.Y(n_178)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_147),
.Y(n_153)
);

INVxp67_ASAP7_75t_L g234 ( 
.A(n_148),
.Y(n_234)
);

INVxp67_ASAP7_75t_L g163 ( 
.A(n_149),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_151),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_164),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_156),
.A2(n_157),
.B1(n_158),
.B2(n_159),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_156),
.B(n_159),
.C(n_164),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_157),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_159),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_165),
.Y(n_175)
);

CKINVDCx16_ASAP7_75t_R g167 ( 
.A(n_168),
.Y(n_167)
);

AOI21xp5_ASAP7_75t_L g169 ( 
.A1(n_170),
.A2(n_179),
.B(n_191),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_177),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_SL g191 ( 
.A(n_171),
.B(n_177),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_172),
.A2(n_174),
.B1(n_175),
.B2(n_176),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_173),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_SL g179 ( 
.A1(n_180),
.A2(n_186),
.B(n_190),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_183),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_181),
.B(n_183),
.Y(n_190)
);

INVxp67_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_187),
.B(n_188),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_195),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_SL g214 ( 
.A(n_194),
.B(n_195),
.Y(n_214)
);

AOI22xp33_ASAP7_75t_SL g195 ( 
.A1(n_196),
.A2(n_197),
.B1(n_206),
.B2(n_213),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_198),
.A2(n_200),
.B1(n_204),
.B2(n_205),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_198),
.Y(n_205)
);

CKINVDCx16_ASAP7_75t_R g204 ( 
.A(n_200),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_200),
.B(n_205),
.C(n_213),
.Y(n_216)
);

INVxp67_ASAP7_75t_L g271 ( 
.A(n_202),
.Y(n_271)
);

INVxp67_ASAP7_75t_L g223 ( 
.A(n_203),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_206),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_210),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_207),
.B(n_210),
.Y(n_232)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_217),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_216),
.B(n_217),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_231),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_218),
.B(n_232),
.C(n_233),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_219),
.A2(n_220),
.B1(n_224),
.B2(n_230),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_219),
.B(n_227),
.C(n_228),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_220),
.Y(n_219)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_224),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_225),
.A2(n_227),
.B1(n_228),
.B2(n_229),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_225),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_227),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_233),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_238),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_SL g261 ( 
.A(n_237),
.B(n_238),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_250),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_L g239 ( 
.A1(n_240),
.A2(n_247),
.B1(n_248),
.B2(n_249),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_240),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_240),
.B(n_249),
.C(n_250),
.Y(n_293)
);

AOI22x1_ASAP7_75t_SL g240 ( 
.A1(n_241),
.A2(n_242),
.B1(n_244),
.B2(n_245),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_241),
.B(n_245),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_242),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_245),
.Y(n_244)
);

CKINVDCx14_ASAP7_75t_R g249 ( 
.A(n_247),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_258),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_252),
.A2(n_254),
.B1(n_255),
.B2(n_257),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_252),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_254),
.B(n_257),
.C(n_258),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_255),
.Y(n_254)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

AOI21xp33_ASAP7_75t_L g316 ( 
.A1(n_263),
.A2(n_317),
.B(n_318),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_264),
.B(n_278),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_264),
.B(n_278),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_274),
.C(n_277),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_265),
.B(n_295),
.Y(n_294)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_266),
.B(n_273),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_267),
.A2(n_269),
.B1(n_270),
.B2(n_272),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_267),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_269),
.B(n_272),
.C(n_273),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_270),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_274),
.B(n_277),
.Y(n_295)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_275),
.B(n_276),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_275),
.B(n_276),
.Y(n_283)
);

AOI22xp33_ASAP7_75t_SL g278 ( 
.A1(n_279),
.A2(n_280),
.B1(n_290),
.B2(n_291),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_281),
.B(n_282),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_281),
.B(n_282),
.C(n_291),
.Y(n_311)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_283),
.B(n_284),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_283),
.B(n_287),
.C(n_289),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_285),
.A2(n_287),
.B1(n_288),
.B2(n_289),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_285),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_288),
.Y(n_287)
);

CKINVDCx16_ASAP7_75t_R g291 ( 
.A(n_290),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_293),
.B(n_294),
.Y(n_292)
);

AND2x2_ASAP7_75t_L g317 ( 
.A(n_293),
.B(n_294),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_297),
.B(n_305),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_SL g320 ( 
.A(n_297),
.B(n_305),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_298),
.B(n_302),
.C(n_304),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_SL g313 ( 
.A1(n_298),
.A2(n_299),
.B1(n_302),
.B2(n_314),
.Y(n_313)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

CKINVDCx16_ASAP7_75t_R g314 ( 
.A(n_302),
.Y(n_314)
);

XOR2xp5_ASAP7_75t_L g312 ( 
.A(n_304),
.B(n_313),
.Y(n_312)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

OAI21xp5_ASAP7_75t_SL g315 ( 
.A1(n_310),
.A2(n_316),
.B(n_319),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_311),
.B(n_312),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_SL g319 ( 
.A(n_311),
.B(n_312),
.Y(n_319)
);


endmodule