module fake_netlist_5_2438_n_1648 (n_137, n_91, n_82, n_122, n_142, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_60, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_125, n_35, n_128, n_73, n_17, n_92, n_19, n_120, n_135, n_30, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_29, n_79, n_131, n_47, n_25, n_53, n_8, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_109, n_112, n_85, n_95, n_119, n_59, n_26, n_133, n_55, n_99, n_2, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_12, n_67, n_121, n_36, n_76, n_87, n_27, n_64, n_77, n_102, n_106, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_134, n_32, n_41, n_104, n_103, n_56, n_51, n_63, n_97, n_141, n_11, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_1648);

input n_137;
input n_91;
input n_82;
input n_122;
input n_142;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_60;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_125;
input n_35;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_120;
input n_135;
input n_30;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_29;
input n_79;
input n_131;
input n_47;
input n_25;
input n_53;
input n_8;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_109;
input n_112;
input n_85;
input n_95;
input n_119;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_27;
input n_64;
input n_77;
input n_102;
input n_106;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_134;
input n_32;
input n_41;
input n_104;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_11;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_1648;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1166;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1150;
wire n_226;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_155;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1021;
wire n_551;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_1545;
wire n_864;
wire n_173;
wire n_859;
wire n_951;
wire n_1264;
wire n_447;
wire n_247;
wire n_1494;
wire n_292;
wire n_625;
wire n_854;
wire n_1462;
wire n_1580;
wire n_674;
wire n_417;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_1607;
wire n_1563;
wire n_606;
wire n_275;
wire n_877;
wire n_755;
wire n_1118;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1359;
wire n_530;
wire n_150;
wire n_1107;
wire n_556;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_929;
wire n_1124;
wire n_902;
wire n_1576;
wire n_191;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1257;
wire n_171;
wire n_1182;
wire n_579;
wire n_1261;
wire n_938;
wire n_1098;
wire n_320;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_406;
wire n_519;
wire n_1016;
wire n_1243;
wire n_546;
wire n_1280;
wire n_281;
wire n_240;
wire n_291;
wire n_231;
wire n_257;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_317;
wire n_1236;
wire n_1633;
wire n_569;
wire n_227;
wire n_920;
wire n_1289;
wire n_1517;
wire n_335;
wire n_370;
wire n_976;
wire n_343;
wire n_1449;
wire n_308;
wire n_1566;
wire n_297;
wire n_156;
wire n_1078;
wire n_775;
wire n_219;
wire n_157;
wire n_600;
wire n_1484;
wire n_1374;
wire n_1328;
wire n_223;
wire n_264;
wire n_1598;
wire n_955;
wire n_163;
wire n_339;
wire n_1146;
wire n_882;
wire n_183;
wire n_243;
wire n_1036;
wire n_1097;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_215;
wire n_350;
wire n_196;
wire n_798;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_580;
wire n_290;
wire n_1040;
wire n_578;
wire n_926;
wire n_344;
wire n_1218;
wire n_422;
wire n_475;
wire n_777;
wire n_1070;
wire n_1547;
wire n_1030;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_663;
wire n_845;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_680;
wire n_1473;
wire n_1587;
wire n_395;
wire n_164;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_214;
wire n_675;
wire n_888;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1384;
wire n_1556;
wire n_184;
wire n_446;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_468;
wire n_213;
wire n_342;
wire n_464;
wire n_363;
wire n_1582;
wire n_197;
wire n_1069;
wire n_1075;
wire n_1450;
wire n_1322;
wire n_1471;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1599;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_907;
wire n_1447;
wire n_1377;
wire n_190;
wire n_989;
wire n_1039;
wire n_228;
wire n_283;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_310;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1248;
wire n_230;
wire n_1331;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_476;
wire n_1527;
wire n_534;
wire n_884;
wire n_345;
wire n_944;
wire n_1623;
wire n_1565;
wire n_182;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_857;
wire n_832;
wire n_207;
wire n_561;
wire n_1319;
wire n_1387;
wire n_1532;
wire n_1027;
wire n_971;
wire n_1156;
wire n_326;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1538;
wire n_1199;
wire n_352;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_887;
wire n_154;
wire n_300;
wire n_809;
wire n_931;
wire n_870;
wire n_599;
wire n_1481;
wire n_434;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1629;
wire n_1293;
wire n_965;
wire n_935;
wire n_1175;
wire n_817;
wire n_360;
wire n_1479;
wire n_759;
wire n_806;
wire n_1477;
wire n_324;
wire n_1635;
wire n_1571;
wire n_187;
wire n_1189;
wire n_1259;
wire n_706;
wire n_746;
wire n_747;
wire n_784;
wire n_1244;
wire n_431;
wire n_1194;
wire n_615;
wire n_851;
wire n_843;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_776;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1647;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_284;
wire n_1128;
wire n_744;
wire n_629;
wire n_590;
wire n_1308;
wire n_254;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_526;
wire n_293;
wire n_372;
wire n_677;
wire n_244;
wire n_1333;
wire n_1121;
wire n_368;
wire n_314;
wire n_433;
wire n_604;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_498;
wire n_1468;
wire n_1559;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_252;
wire n_624;
wire n_1380;
wire n_1617;
wire n_295;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_610;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_448;
wire n_259;
wire n_758;
wire n_999;
wire n_1158;
wire n_1509;
wire n_563;
wire n_1145;
wire n_878;
wire n_524;
wire n_204;
wire n_394;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_331;
wire n_906;
wire n_1163;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_658;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_152;
wire n_940;
wire n_1445;
wire n_1492;
wire n_592;
wire n_1169;
wire n_1596;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1269;
wire n_1095;
wire n_1614;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_1431;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1640;
wire n_1009;
wire n_1148;
wire n_742;
wire n_750;
wire n_995;
wire n_454;
wire n_1609;
wire n_374;
wire n_185;
wire n_396;
wire n_1383;
wire n_1073;
wire n_255;
wire n_662;
wire n_459;
wire n_218;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1574;
wire n_473;
wire n_1309;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_1548;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_168;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_208;
wire n_743;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_1240;
wire n_829;
wire n_1612;
wire n_1416;
wire n_361;
wire n_700;
wire n_1237;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1568;
wire n_1006;
wire n_329;
wire n_274;
wire n_1270;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_309;
wire n_512;
wire n_1591;
wire n_322;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1349;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_224;
wire n_1562;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_239;
wire n_630;
wire n_504;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_1304;
wire n_1324;
wire n_987;
wire n_261;
wire n_174;
wire n_1455;
wire n_767;
wire n_993;
wire n_1407;
wire n_1551;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_729;
wire n_1131;
wire n_1084;
wire n_970;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_340;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_1645;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_233;
wire n_572;
wire n_366;
wire n_815;
wire n_327;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_426;
wire n_1438;
wire n_1082;
wire n_589;
wire n_716;
wire n_1630;
wire n_562;
wire n_1436;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_531;
wire n_890;
wire n_764;
wire n_1056;
wire n_1424;
wire n_162;
wire n_960;
wire n_222;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_634;
wire n_199;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_1519;
wire n_256;
wire n_950;
wire n_1553;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1060;
wire n_1141;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_912;
wire n_968;
wire n_315;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_1608;
wire n_983;
wire n_280;
wire n_1305;
wire n_873;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_1644;
wire n_690;
wire n_583;
wire n_302;
wire n_1343;
wire n_1203;
wire n_1631;
wire n_821;
wire n_321;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1288;
wire n_385;
wire n_212;
wire n_507;
wire n_1560;
wire n_1605;
wire n_330;
wire n_1228;
wire n_972;
wire n_692;
wire n_820;
wire n_1200;
wire n_1301;
wire n_1363;
wire n_1185;
wire n_991;
wire n_828;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_945;
wire n_492;
wire n_153;
wire n_1504;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_286;
wire n_1643;
wire n_883;
wire n_470;
wire n_325;
wire n_449;
wire n_1594;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_856;
wire n_918;
wire n_942;
wire n_189;
wire n_1147;
wire n_1557;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_195;
wire n_356;
wire n_894;
wire n_1636;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1470;
wire n_1096;
wire n_234;
wire n_1575;
wire n_833;
wire n_1646;
wire n_225;
wire n_1307;
wire n_988;
wire n_814;
wire n_192;
wire n_1549;
wire n_1201;
wire n_1114;
wire n_655;
wire n_1616;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_387;
wire n_1149;
wire n_398;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_211;
wire n_1219;
wire n_1204;
wire n_178;
wire n_1035;
wire n_287;
wire n_555;
wire n_783;
wire n_1188;
wire n_661;
wire n_849;
wire n_336;
wire n_681;
wire n_584;
wire n_1638;
wire n_430;
wire n_510;
wire n_216;
wire n_311;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_445;
wire n_749;
wire n_1134;
wire n_1358;
wire n_717;
wire n_165;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_249;
wire n_304;
wire n_1338;
wire n_577;
wire n_1522;
wire n_1637;
wire n_1419;
wire n_338;
wire n_149;
wire n_693;
wire n_1506;
wire n_836;
wire n_990;
wire n_1389;
wire n_975;
wire n_1256;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_151;
wire n_306;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1164;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_1572;
wire n_876;
wire n_1516;
wire n_1190;
wire n_601;
wire n_917;
wire n_966;
wire n_253;
wire n_1116;
wire n_1212;
wire n_1541;
wire n_206;
wire n_172;
wire n_217;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_818;
wire n_861;
wire n_1183;
wire n_899;
wire n_1253;
wire n_210;
wire n_774;
wire n_1628;
wire n_1335;
wire n_1514;
wire n_1059;
wire n_1345;
wire n_176;
wire n_1133;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_1168;
wire n_707;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_1584;
wire n_665;
wire n_1440;
wire n_177;
wire n_421;
wire n_1356;
wire n_910;
wire n_768;
wire n_1475;
wire n_1302;
wire n_205;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_179;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_735;
wire n_232;
wire n_1109;
wire n_895;
wire n_1310;
wire n_202;
wire n_427;
wire n_1399;
wire n_1543;
wire n_791;
wire n_732;
wire n_1533;
wire n_193;
wire n_808;
wire n_797;
wire n_1025;
wire n_500;
wire n_1067;
wire n_435;
wire n_159;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_594;
wire n_200;
wire n_1291;
wire n_1297;
wire n_1155;
wire n_1418;
wire n_1524;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_985;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1352;
wire n_626;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_305;
wire n_676;
wire n_294;
wire n_318;
wire n_653;
wire n_642;
wire n_1602;
wire n_194;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_268;
wire n_664;
wire n_503;
wire n_235;
wire n_1372;
wire n_605;
wire n_1273;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_581;
wire n_382;
wire n_554;
wire n_1625;
wire n_898;
wire n_1013;
wire n_1452;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_198;
wire n_714;
wire n_909;
wire n_1497;
wire n_1530;
wire n_997;
wire n_932;
wire n_612;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_508;
wire n_506;
wire n_1320;
wire n_737;
wire n_986;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1281;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_209;
wire n_1564;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1376;
wire n_941;
wire n_981;
wire n_1569;
wire n_867;
wire n_186;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_518;
wire n_505;
wire n_282;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1620;
wire n_381;
wire n_220;
wire n_390;
wire n_1330;
wire n_481;
wire n_1554;
wire n_769;
wire n_1046;
wire n_271;
wire n_934;
wire n_1618;
wire n_826;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_167;
wire n_428;
wire n_379;
wire n_1341;
wire n_570;
wire n_1641;
wire n_1361;
wire n_853;
wire n_377;
wire n_751;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_158;
wire n_704;
wire n_787;
wire n_961;
wire n_771;
wire n_276;
wire n_1225;
wire n_1520;
wire n_169;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_181;
wire n_1411;
wire n_221;
wire n_622;
wire n_1577;
wire n_1087;
wire n_386;
wire n_994;
wire n_848;
wire n_1550;
wire n_1498;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_591;
wire n_1536;
wire n_1344;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_432;
wire n_839;
wire n_1210;
wire n_1364;
wire n_328;
wire n_1250;
wire n_369;
wire n_871;
wire n_598;
wire n_685;
wire n_608;
wire n_928;
wire n_1367;
wire n_1460;
wire n_772;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_402;
wire n_413;
wire n_1086;
wire n_796;
wire n_1619;
wire n_236;
wire n_1502;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_903;
wire n_1525;
wire n_740;
wire n_203;
wire n_384;
wire n_1404;
wire n_1315;
wire n_277;
wire n_1061;
wire n_333;
wire n_1298;
wire n_462;
wire n_1193;
wire n_1255;
wire n_258;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_188;
wire n_844;
wire n_201;
wire n_471;
wire n_852;
wire n_1487;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_465;
wire n_362;
wire n_1321;
wire n_170;
wire n_161;
wire n_273;
wire n_585;
wire n_270;
wire n_616;
wire n_745;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_641;
wire n_730;
wire n_1325;
wire n_1595;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_180;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1540;
wire n_229;
wire n_437;
wire n_1642;
wire n_403;
wire n_453;
wire n_1130;
wire n_720;
wire n_1526;
wire n_863;
wire n_805;
wire n_1604;
wire n_1275;
wire n_712;
wire n_246;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_269;
wire n_285;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_1621;
wire n_251;
wire n_160;
wire n_566;
wire n_565;
wire n_1448;
wire n_1507;
wire n_1398;
wire n_597;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_651;
wire n_1340;
wire n_334;
wire n_811;
wire n_1558;
wire n_807;
wire n_835;
wire n_175;
wire n_666;
wire n_262;
wire n_1433;
wire n_1254;
wire n_1026;
wire n_1234;
wire n_319;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_242;
wire n_1018;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_166;
wire n_1180;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;
wire n_278;

CKINVDCx5p33_ASAP7_75t_R g149 ( 
.A(n_31),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_40),
.Y(n_150)
);

CKINVDCx5p33_ASAP7_75t_R g151 ( 
.A(n_132),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_109),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_82),
.Y(n_153)
);

CKINVDCx5p33_ASAP7_75t_R g154 ( 
.A(n_125),
.Y(n_154)
);

CKINVDCx5p33_ASAP7_75t_R g155 ( 
.A(n_50),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_8),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_52),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_89),
.Y(n_158)
);

CKINVDCx5p33_ASAP7_75t_R g159 ( 
.A(n_85),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_114),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_138),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_15),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_77),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_23),
.Y(n_164)
);

BUFx3_ASAP7_75t_L g165 ( 
.A(n_15),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_51),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_30),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_134),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_127),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_111),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_93),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_60),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_3),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_136),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_63),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_43),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_86),
.Y(n_177)
);

INVx1_ASAP7_75t_SL g178 ( 
.A(n_98),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_27),
.Y(n_179)
);

INVx1_ASAP7_75t_SL g180 ( 
.A(n_49),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_102),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_145),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_28),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_135),
.Y(n_184)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_96),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_90),
.Y(n_186)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_83),
.Y(n_187)
);

INVx1_ASAP7_75t_SL g188 ( 
.A(n_110),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_43),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_21),
.Y(n_190)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_8),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_24),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_67),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_16),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_46),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_33),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_37),
.Y(n_197)
);

INVx1_ASAP7_75t_SL g198 ( 
.A(n_4),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_87),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_28),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_65),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_42),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_24),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_66),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_142),
.Y(n_205)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_41),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_101),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_55),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_144),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_25),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_0),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_53),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_36),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_92),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_54),
.Y(n_215)
);

BUFx10_ASAP7_75t_L g216 ( 
.A(n_81),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_105),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_57),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_9),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_115),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_103),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_70),
.Y(n_222)
);

BUFx6f_ASAP7_75t_L g223 ( 
.A(n_30),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_147),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_100),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_130),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_16),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_47),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_35),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_124),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_97),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_141),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_40),
.Y(n_233)
);

INVx1_ASAP7_75t_SL g234 ( 
.A(n_64),
.Y(n_234)
);

INVx2_ASAP7_75t_SL g235 ( 
.A(n_0),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_38),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_5),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_76),
.Y(n_238)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_47),
.Y(n_239)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_94),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_37),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_88),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_10),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_1),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_22),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_17),
.Y(n_246)
);

BUFx6f_ASAP7_75t_L g247 ( 
.A(n_72),
.Y(n_247)
);

BUFx2_ASAP7_75t_SL g248 ( 
.A(n_113),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_35),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_123),
.Y(n_250)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_42),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_122),
.Y(n_252)
);

INVx1_ASAP7_75t_SL g253 ( 
.A(n_117),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_128),
.Y(n_254)
);

BUFx6f_ASAP7_75t_L g255 ( 
.A(n_91),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_74),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_139),
.Y(n_257)
);

HB1xp67_ASAP7_75t_L g258 ( 
.A(n_56),
.Y(n_258)
);

INVx1_ASAP7_75t_SL g259 ( 
.A(n_112),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_5),
.Y(n_260)
);

INVx2_ASAP7_75t_SL g261 ( 
.A(n_131),
.Y(n_261)
);

INVx2_ASAP7_75t_SL g262 ( 
.A(n_19),
.Y(n_262)
);

BUFx3_ASAP7_75t_L g263 ( 
.A(n_34),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_1),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_99),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_6),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_119),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_12),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_11),
.Y(n_269)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_68),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_29),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_25),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_2),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_120),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_3),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_18),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_148),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_7),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_69),
.Y(n_279)
);

INVx2_ASAP7_75t_SL g280 ( 
.A(n_2),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_19),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_48),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_143),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_4),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_18),
.Y(n_285)
);

BUFx3_ASAP7_75t_L g286 ( 
.A(n_12),
.Y(n_286)
);

BUFx3_ASAP7_75t_L g287 ( 
.A(n_31),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_58),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_121),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_118),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_10),
.Y(n_291)
);

INVx1_ASAP7_75t_SL g292 ( 
.A(n_13),
.Y(n_292)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_17),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_9),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_61),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_6),
.Y(n_296)
);

CKINVDCx16_ASAP7_75t_R g297 ( 
.A(n_32),
.Y(n_297)
);

INVx1_ASAP7_75t_SL g298 ( 
.A(n_21),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_73),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_29),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_11),
.Y(n_301)
);

BUFx10_ASAP7_75t_L g302 ( 
.A(n_133),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_129),
.Y(n_303)
);

INVx2_ASAP7_75t_SL g304 ( 
.A(n_95),
.Y(n_304)
);

HB1xp67_ASAP7_75t_L g305 ( 
.A(n_297),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_150),
.Y(n_306)
);

INVxp67_ASAP7_75t_L g307 ( 
.A(n_156),
.Y(n_307)
);

INVxp67_ASAP7_75t_SL g308 ( 
.A(n_258),
.Y(n_308)
);

INVxp67_ASAP7_75t_SL g309 ( 
.A(n_150),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_152),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_157),
.Y(n_311)
);

HB1xp67_ASAP7_75t_L g312 ( 
.A(n_149),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_163),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_150),
.Y(n_314)
);

INVxp67_ASAP7_75t_SL g315 ( 
.A(n_150),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_150),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_223),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_199),
.Y(n_318)
);

HB1xp67_ASAP7_75t_L g319 ( 
.A(n_149),
.Y(n_319)
);

HB1xp67_ASAP7_75t_L g320 ( 
.A(n_167),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_223),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_223),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_201),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_223),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_223),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_174),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_184),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_191),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_191),
.Y(n_329)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_247),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_215),
.Y(n_331)
);

INVxp67_ASAP7_75t_SL g332 ( 
.A(n_165),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_204),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_207),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_208),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_214),
.Y(n_336)
);

INVxp67_ASAP7_75t_SL g337 ( 
.A(n_165),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_206),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_206),
.Y(n_339)
);

HB1xp67_ASAP7_75t_L g340 ( 
.A(n_167),
.Y(n_340)
);

CKINVDCx20_ASAP7_75t_R g341 ( 
.A(n_283),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_239),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_239),
.Y(n_343)
);

INVxp67_ASAP7_75t_L g344 ( 
.A(n_162),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_251),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_251),
.Y(n_346)
);

INVxp33_ASAP7_75t_SL g347 ( 
.A(n_179),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_293),
.Y(n_348)
);

INVxp67_ASAP7_75t_SL g349 ( 
.A(n_263),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_293),
.Y(n_350)
);

CKINVDCx14_ASAP7_75t_R g351 ( 
.A(n_216),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_263),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_286),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_286),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_218),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_287),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_287),
.Y(n_357)
);

HB1xp67_ASAP7_75t_L g358 ( 
.A(n_179),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_176),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_192),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_195),
.Y(n_361)
);

HB1xp67_ASAP7_75t_L g362 ( 
.A(n_268),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_228),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_229),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_243),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_244),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_246),
.Y(n_367)
);

BUFx6f_ASAP7_75t_L g368 ( 
.A(n_247),
.Y(n_368)
);

INVx2_ASAP7_75t_L g369 ( 
.A(n_247),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_249),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_220),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_266),
.Y(n_372)
);

INVx2_ASAP7_75t_L g373 ( 
.A(n_247),
.Y(n_373)
);

INVxp67_ASAP7_75t_L g374 ( 
.A(n_269),
.Y(n_374)
);

INVxp67_ASAP7_75t_SL g375 ( 
.A(n_153),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_273),
.Y(n_376)
);

CKINVDCx20_ASAP7_75t_R g377 ( 
.A(n_222),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_284),
.Y(n_378)
);

INVxp33_ASAP7_75t_SL g379 ( 
.A(n_268),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_291),
.Y(n_380)
);

AND2x4_ASAP7_75t_L g381 ( 
.A(n_309),
.B(n_261),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_R g382 ( 
.A(n_351),
.B(n_224),
.Y(n_382)
);

BUFx6f_ASAP7_75t_L g383 ( 
.A(n_368),
.Y(n_383)
);

NAND2xp33_ASAP7_75t_L g384 ( 
.A(n_318),
.B(n_271),
.Y(n_384)
);

HB1xp67_ASAP7_75t_L g385 ( 
.A(n_305),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_306),
.Y(n_386)
);

AND2x4_ASAP7_75t_L g387 ( 
.A(n_315),
.B(n_261),
.Y(n_387)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_330),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_306),
.Y(n_389)
);

BUFx3_ASAP7_75t_L g390 ( 
.A(n_314),
.Y(n_390)
);

INVx2_ASAP7_75t_L g391 ( 
.A(n_330),
.Y(n_391)
);

AND2x2_ASAP7_75t_L g392 ( 
.A(n_332),
.B(n_235),
.Y(n_392)
);

INVx2_ASAP7_75t_L g393 ( 
.A(n_330),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_323),
.B(n_304),
.Y(n_394)
);

BUFx8_ASAP7_75t_L g395 ( 
.A(n_352),
.Y(n_395)
);

OAI22xp5_ASAP7_75t_SL g396 ( 
.A1(n_310),
.A2(n_164),
.B1(n_173),
.B2(n_190),
.Y(n_396)
);

INVx6_ASAP7_75t_L g397 ( 
.A(n_368),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_SL g398 ( 
.A(n_347),
.B(n_216),
.Y(n_398)
);

INVx2_ASAP7_75t_L g399 ( 
.A(n_369),
.Y(n_399)
);

OA21x2_ASAP7_75t_L g400 ( 
.A1(n_369),
.A2(n_187),
.B(n_185),
.Y(n_400)
);

AND2x2_ASAP7_75t_L g401 ( 
.A(n_337),
.B(n_235),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_333),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_314),
.Y(n_403)
);

BUFx6f_ASAP7_75t_L g404 ( 
.A(n_368),
.Y(n_404)
);

CKINVDCx8_ASAP7_75t_R g405 ( 
.A(n_334),
.Y(n_405)
);

INVx2_ASAP7_75t_L g406 ( 
.A(n_369),
.Y(n_406)
);

BUFx6f_ASAP7_75t_L g407 ( 
.A(n_368),
.Y(n_407)
);

NOR2xp33_ASAP7_75t_L g408 ( 
.A(n_335),
.B(n_304),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_336),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_355),
.B(n_185),
.Y(n_410)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_373),
.Y(n_411)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_373),
.Y(n_412)
);

BUFx6f_ASAP7_75t_L g413 ( 
.A(n_368),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_371),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_SL g415 ( 
.A(n_379),
.B(n_216),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_349),
.B(n_187),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_375),
.B(n_308),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_377),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_SL g419 ( 
.A(n_312),
.B(n_302),
.Y(n_419)
);

INVx2_ASAP7_75t_L g420 ( 
.A(n_373),
.Y(n_420)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_368),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_311),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_316),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_316),
.Y(n_424)
);

NOR2xp33_ASAP7_75t_L g425 ( 
.A(n_319),
.B(n_320),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_317),
.Y(n_426)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_317),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_321),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_SL g429 ( 
.A(n_340),
.B(n_302),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_321),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_322),
.Y(n_431)
);

BUFx2_ASAP7_75t_L g432 ( 
.A(n_358),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_322),
.Y(n_433)
);

HB1xp67_ASAP7_75t_L g434 ( 
.A(n_362),
.Y(n_434)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_324),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_324),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_325),
.Y(n_437)
);

BUFx8_ASAP7_75t_L g438 ( 
.A(n_352),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_325),
.Y(n_439)
);

HB1xp67_ASAP7_75t_L g440 ( 
.A(n_353),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_359),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_313),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_353),
.B(n_240),
.Y(n_443)
);

INVx4_ASAP7_75t_L g444 ( 
.A(n_328),
.Y(n_444)
);

INVx2_ASAP7_75t_L g445 ( 
.A(n_328),
.Y(n_445)
);

AND2x6_ASAP7_75t_L g446 ( 
.A(n_329),
.B(n_247),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_359),
.Y(n_447)
);

BUFx6f_ASAP7_75t_L g448 ( 
.A(n_329),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_360),
.Y(n_449)
);

CKINVDCx16_ASAP7_75t_R g450 ( 
.A(n_326),
.Y(n_450)
);

CKINVDCx20_ASAP7_75t_R g451 ( 
.A(n_327),
.Y(n_451)
);

NOR2xp33_ASAP7_75t_L g452 ( 
.A(n_394),
.B(n_354),
.Y(n_452)
);

INVx2_ASAP7_75t_L g453 ( 
.A(n_427),
.Y(n_453)
);

INVx2_ASAP7_75t_L g454 ( 
.A(n_427),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_390),
.Y(n_455)
);

AOI22xp33_ASAP7_75t_L g456 ( 
.A1(n_381),
.A2(n_280),
.B1(n_262),
.B2(n_300),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_SL g457 ( 
.A(n_382),
.B(n_302),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_381),
.B(n_178),
.Y(n_458)
);

INVx3_ASAP7_75t_L g459 ( 
.A(n_383),
.Y(n_459)
);

INVx3_ASAP7_75t_L g460 ( 
.A(n_383),
.Y(n_460)
);

INVx3_ASAP7_75t_L g461 ( 
.A(n_383),
.Y(n_461)
);

BUFx10_ASAP7_75t_L g462 ( 
.A(n_402),
.Y(n_462)
);

NOR2x1p5_ASAP7_75t_L g463 ( 
.A(n_409),
.B(n_271),
.Y(n_463)
);

INVx2_ASAP7_75t_L g464 ( 
.A(n_427),
.Y(n_464)
);

BUFx6f_ASAP7_75t_SL g465 ( 
.A(n_381),
.Y(n_465)
);

BUFx3_ASAP7_75t_L g466 ( 
.A(n_390),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_390),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_386),
.Y(n_468)
);

INVx4_ASAP7_75t_L g469 ( 
.A(n_383),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_SL g470 ( 
.A(n_405),
.B(n_151),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_386),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_389),
.Y(n_472)
);

NOR2x1p5_ASAP7_75t_L g473 ( 
.A(n_414),
.B(n_272),
.Y(n_473)
);

INVx2_ASAP7_75t_L g474 ( 
.A(n_435),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_381),
.B(n_180),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_387),
.B(n_188),
.Y(n_476)
);

INVx2_ASAP7_75t_L g477 ( 
.A(n_435),
.Y(n_477)
);

INVx2_ASAP7_75t_SL g478 ( 
.A(n_392),
.Y(n_478)
);

INVx2_ASAP7_75t_L g479 ( 
.A(n_435),
.Y(n_479)
);

BUFx2_ASAP7_75t_L g480 ( 
.A(n_385),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_389),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_403),
.Y(n_482)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_448),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_403),
.Y(n_484)
);

INVxp33_ASAP7_75t_L g485 ( 
.A(n_425),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_423),
.Y(n_486)
);

OAI22xp33_ASAP7_75t_L g487 ( 
.A1(n_417),
.A2(n_292),
.B1(n_198),
.B2(n_298),
.Y(n_487)
);

OAI22xp33_ASAP7_75t_SL g488 ( 
.A1(n_410),
.A2(n_280),
.B1(n_262),
.B2(n_374),
.Y(n_488)
);

NOR3xp33_ASAP7_75t_L g489 ( 
.A(n_396),
.B(n_344),
.C(n_307),
.Y(n_489)
);

INVx3_ASAP7_75t_L g490 ( 
.A(n_383),
.Y(n_490)
);

INVx4_ASAP7_75t_L g491 ( 
.A(n_383),
.Y(n_491)
);

INVxp67_ASAP7_75t_L g492 ( 
.A(n_432),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_387),
.B(n_234),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_SL g494 ( 
.A(n_405),
.B(n_151),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_SL g495 ( 
.A(n_408),
.B(n_154),
.Y(n_495)
);

BUFx8_ASAP7_75t_SL g496 ( 
.A(n_451),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_SL g497 ( 
.A(n_398),
.B(n_415),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_387),
.B(n_253),
.Y(n_498)
);

INVx3_ASAP7_75t_L g499 ( 
.A(n_404),
.Y(n_499)
);

OR2x6_ASAP7_75t_L g500 ( 
.A(n_419),
.B(n_248),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_SL g501 ( 
.A(n_429),
.B(n_154),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_440),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_441),
.Y(n_503)
);

INVx2_ASAP7_75t_L g504 ( 
.A(n_448),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_441),
.Y(n_505)
);

AOI22xp33_ASAP7_75t_L g506 ( 
.A1(n_387),
.A2(n_301),
.B1(n_294),
.B2(n_270),
.Y(n_506)
);

OR2x6_ASAP7_75t_L g507 ( 
.A(n_432),
.B(n_354),
.Y(n_507)
);

AO22x2_ASAP7_75t_L g508 ( 
.A1(n_392),
.A2(n_270),
.B1(n_240),
.B2(n_401),
.Y(n_508)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_448),
.Y(n_509)
);

NAND2xp33_ASAP7_75t_L g510 ( 
.A(n_446),
.B(n_255),
.Y(n_510)
);

INVx5_ASAP7_75t_L g511 ( 
.A(n_446),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_423),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_L g513 ( 
.A(n_401),
.B(n_259),
.Y(n_513)
);

HB1xp67_ASAP7_75t_L g514 ( 
.A(n_434),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_424),
.Y(n_515)
);

BUFx6f_ASAP7_75t_L g516 ( 
.A(n_404),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_424),
.Y(n_517)
);

INVx2_ASAP7_75t_L g518 ( 
.A(n_448),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_SL g519 ( 
.A(n_395),
.B(n_438),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_426),
.Y(n_520)
);

INVx4_ASAP7_75t_L g521 ( 
.A(n_404),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_426),
.Y(n_522)
);

INVx2_ASAP7_75t_L g523 ( 
.A(n_448),
.Y(n_523)
);

INVxp33_ASAP7_75t_L g524 ( 
.A(n_396),
.Y(n_524)
);

BUFx6f_ASAP7_75t_L g525 ( 
.A(n_404),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_428),
.Y(n_526)
);

INVx2_ASAP7_75t_L g527 ( 
.A(n_448),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_416),
.B(n_225),
.Y(n_528)
);

INVx8_ASAP7_75t_L g529 ( 
.A(n_446),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_428),
.Y(n_530)
);

INVx1_ASAP7_75t_SL g531 ( 
.A(n_418),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_430),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_430),
.Y(n_533)
);

BUFx6f_ASAP7_75t_SL g534 ( 
.A(n_447),
.Y(n_534)
);

OR2x6_ASAP7_75t_L g535 ( 
.A(n_443),
.B(n_356),
.Y(n_535)
);

INVx2_ASAP7_75t_L g536 ( 
.A(n_431),
.Y(n_536)
);

HB1xp67_ASAP7_75t_L g537 ( 
.A(n_422),
.Y(n_537)
);

INVx2_ASAP7_75t_L g538 ( 
.A(n_431),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_433),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_433),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_436),
.Y(n_541)
);

INVx2_ASAP7_75t_SL g542 ( 
.A(n_395),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_SL g543 ( 
.A(n_395),
.B(n_155),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_SL g544 ( 
.A(n_395),
.B(n_155),
.Y(n_544)
);

INVx2_ASAP7_75t_L g545 ( 
.A(n_436),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_437),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_437),
.Y(n_547)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_439),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_439),
.Y(n_549)
);

NOR2xp33_ASAP7_75t_R g550 ( 
.A(n_442),
.B(n_331),
.Y(n_550)
);

INVx3_ASAP7_75t_L g551 ( 
.A(n_404),
.Y(n_551)
);

INVx2_ASAP7_75t_L g552 ( 
.A(n_388),
.Y(n_552)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_388),
.Y(n_553)
);

AND2x2_ASAP7_75t_L g554 ( 
.A(n_449),
.B(n_356),
.Y(n_554)
);

INVx2_ASAP7_75t_L g555 ( 
.A(n_388),
.Y(n_555)
);

CKINVDCx5p33_ASAP7_75t_R g556 ( 
.A(n_450),
.Y(n_556)
);

INVx2_ASAP7_75t_SL g557 ( 
.A(n_438),
.Y(n_557)
);

NAND2xp33_ASAP7_75t_L g558 ( 
.A(n_446),
.B(n_255),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_L g559 ( 
.A(n_444),
.B(n_230),
.Y(n_559)
);

INVx2_ASAP7_75t_L g560 ( 
.A(n_391),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_444),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_444),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_444),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_391),
.Y(n_564)
);

INVx2_ASAP7_75t_L g565 ( 
.A(n_391),
.Y(n_565)
);

NOR2xp33_ASAP7_75t_L g566 ( 
.A(n_384),
.B(n_357),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_L g567 ( 
.A(n_421),
.B(n_231),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_393),
.Y(n_568)
);

INVx4_ASAP7_75t_L g569 ( 
.A(n_404),
.Y(n_569)
);

OR2x6_ASAP7_75t_L g570 ( 
.A(n_445),
.B(n_357),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_393),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_399),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_399),
.Y(n_573)
);

OR2x2_ASAP7_75t_L g574 ( 
.A(n_450),
.B(n_360),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_399),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_406),
.Y(n_576)
);

NOR2xp33_ASAP7_75t_L g577 ( 
.A(n_438),
.B(n_341),
.Y(n_577)
);

BUFx3_ASAP7_75t_L g578 ( 
.A(n_400),
.Y(n_578)
);

NOR2xp33_ASAP7_75t_R g579 ( 
.A(n_438),
.B(n_232),
.Y(n_579)
);

AOI22xp33_ASAP7_75t_L g580 ( 
.A1(n_400),
.A2(n_255),
.B1(n_378),
.B2(n_376),
.Y(n_580)
);

BUFx3_ASAP7_75t_L g581 ( 
.A(n_400),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_406),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_406),
.Y(n_583)
);

BUFx6f_ASAP7_75t_L g584 ( 
.A(n_407),
.Y(n_584)
);

INVx3_ASAP7_75t_L g585 ( 
.A(n_407),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_445),
.Y(n_586)
);

INVx3_ASAP7_75t_L g587 ( 
.A(n_407),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_SL g588 ( 
.A(n_445),
.B(n_159),
.Y(n_588)
);

INVx2_ASAP7_75t_L g589 ( 
.A(n_411),
.Y(n_589)
);

INVx3_ASAP7_75t_L g590 ( 
.A(n_407),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_411),
.Y(n_591)
);

OAI22x1_ASAP7_75t_L g592 ( 
.A1(n_400),
.A2(n_285),
.B1(n_296),
.B2(n_281),
.Y(n_592)
);

INVx2_ASAP7_75t_L g593 ( 
.A(n_412),
.Y(n_593)
);

AND2x2_ASAP7_75t_L g594 ( 
.A(n_412),
.B(n_338),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_412),
.Y(n_595)
);

INVx2_ASAP7_75t_L g596 ( 
.A(n_420),
.Y(n_596)
);

INVx3_ASAP7_75t_L g597 ( 
.A(n_407),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_L g598 ( 
.A(n_421),
.B(n_238),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_455),
.Y(n_599)
);

NAND2xp33_ASAP7_75t_L g600 ( 
.A(n_478),
.B(n_242),
.Y(n_600)
);

BUFx6f_ASAP7_75t_SL g601 ( 
.A(n_462),
.Y(n_601)
);

NOR2xp33_ASAP7_75t_L g602 ( 
.A(n_485),
.B(n_159),
.Y(n_602)
);

BUFx5_ASAP7_75t_L g603 ( 
.A(n_578),
.Y(n_603)
);

OR2x6_ASAP7_75t_L g604 ( 
.A(n_519),
.B(n_361),
.Y(n_604)
);

INVx2_ASAP7_75t_L g605 ( 
.A(n_552),
.Y(n_605)
);

INVx2_ASAP7_75t_L g606 ( 
.A(n_552),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_455),
.Y(n_607)
);

NOR2x1p5_ASAP7_75t_L g608 ( 
.A(n_574),
.B(n_272),
.Y(n_608)
);

AO22x2_ASAP7_75t_L g609 ( 
.A1(n_497),
.A2(n_205),
.B1(n_160),
.B2(n_161),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_L g610 ( 
.A(n_452),
.B(n_421),
.Y(n_610)
);

OR2x2_ASAP7_75t_L g611 ( 
.A(n_574),
.B(n_361),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_467),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_L g613 ( 
.A(n_561),
.B(n_158),
.Y(n_613)
);

NOR2xp33_ASAP7_75t_L g614 ( 
.A(n_502),
.B(n_168),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_SL g615 ( 
.A(n_513),
.B(n_168),
.Y(n_615)
);

INVx2_ASAP7_75t_L g616 ( 
.A(n_553),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_L g617 ( 
.A(n_561),
.B(n_166),
.Y(n_617)
);

NOR2xp67_ASAP7_75t_L g618 ( 
.A(n_542),
.B(n_557),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_L g619 ( 
.A(n_562),
.B(n_171),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_SL g620 ( 
.A(n_566),
.B(n_458),
.Y(n_620)
);

INVx2_ASAP7_75t_SL g621 ( 
.A(n_507),
.Y(n_621)
);

NOR3xp33_ASAP7_75t_L g622 ( 
.A(n_487),
.B(n_226),
.C(n_221),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_562),
.B(n_181),
.Y(n_623)
);

BUFx6f_ASAP7_75t_SL g624 ( 
.A(n_462),
.Y(n_624)
);

A2O1A1Ixp33_ASAP7_75t_L g625 ( 
.A1(n_563),
.A2(n_252),
.B(n_182),
.C(n_250),
.Y(n_625)
);

BUFx3_ASAP7_75t_L g626 ( 
.A(n_496),
.Y(n_626)
);

INVx2_ASAP7_75t_SL g627 ( 
.A(n_507),
.Y(n_627)
);

INVx2_ASAP7_75t_L g628 ( 
.A(n_553),
.Y(n_628)
);

NOR2xp33_ASAP7_75t_L g629 ( 
.A(n_475),
.B(n_169),
.Y(n_629)
);

OR2x2_ASAP7_75t_L g630 ( 
.A(n_492),
.B(n_363),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_L g631 ( 
.A(n_563),
.B(n_186),
.Y(n_631)
);

OAI22xp5_ASAP7_75t_SL g632 ( 
.A1(n_524),
.A2(n_245),
.B1(n_282),
.B2(n_202),
.Y(n_632)
);

NOR2xp33_ASAP7_75t_L g633 ( 
.A(n_476),
.B(n_169),
.Y(n_633)
);

NOR2xp33_ASAP7_75t_L g634 ( 
.A(n_493),
.B(n_170),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_L g635 ( 
.A(n_498),
.B(n_193),
.Y(n_635)
);

INVx2_ASAP7_75t_L g636 ( 
.A(n_555),
.Y(n_636)
);

INVx2_ASAP7_75t_L g637 ( 
.A(n_555),
.Y(n_637)
);

OAI22xp33_ASAP7_75t_L g638 ( 
.A1(n_500),
.A2(n_276),
.B1(n_275),
.B2(n_278),
.Y(n_638)
);

NOR2xp33_ASAP7_75t_L g639 ( 
.A(n_528),
.B(n_170),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_L g640 ( 
.A(n_503),
.B(n_209),
.Y(n_640)
);

INVx2_ASAP7_75t_L g641 ( 
.A(n_560),
.Y(n_641)
);

OAI22xp5_ASAP7_75t_L g642 ( 
.A1(n_465),
.A2(n_217),
.B1(n_212),
.B2(n_277),
.Y(n_642)
);

NOR2xp33_ASAP7_75t_L g643 ( 
.A(n_495),
.B(n_172),
.Y(n_643)
);

OR2x2_ASAP7_75t_L g644 ( 
.A(n_507),
.B(n_363),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_L g645 ( 
.A(n_505),
.B(n_420),
.Y(n_645)
);

O2A1O1Ixp5_ASAP7_75t_L g646 ( 
.A1(n_468),
.A2(n_420),
.B(n_370),
.C(n_364),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_554),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_554),
.Y(n_648)
);

BUFx6f_ASAP7_75t_L g649 ( 
.A(n_466),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_L g650 ( 
.A(n_468),
.B(n_407),
.Y(n_650)
);

NOR2xp33_ASAP7_75t_L g651 ( 
.A(n_535),
.B(n_175),
.Y(n_651)
);

AND2x2_ASAP7_75t_L g652 ( 
.A(n_507),
.B(n_364),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_471),
.Y(n_653)
);

AOI22xp33_ASAP7_75t_L g654 ( 
.A1(n_592),
.A2(n_255),
.B1(n_296),
.B2(n_285),
.Y(n_654)
);

INVx2_ASAP7_75t_SL g655 ( 
.A(n_480),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_471),
.B(n_413),
.Y(n_656)
);

INVxp67_ASAP7_75t_L g657 ( 
.A(n_514),
.Y(n_657)
);

CKINVDCx5p33_ASAP7_75t_R g658 ( 
.A(n_550),
.Y(n_658)
);

NAND3xp33_ASAP7_75t_L g659 ( 
.A(n_456),
.B(n_506),
.C(n_489),
.Y(n_659)
);

INVx2_ASAP7_75t_L g660 ( 
.A(n_560),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_SL g661 ( 
.A(n_578),
.B(n_255),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_472),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_SL g663 ( 
.A(n_579),
.B(n_175),
.Y(n_663)
);

AND2x2_ASAP7_75t_L g664 ( 
.A(n_480),
.B(n_365),
.Y(n_664)
);

CKINVDCx5p33_ASAP7_75t_R g665 ( 
.A(n_462),
.Y(n_665)
);

NOR2xp33_ASAP7_75t_L g666 ( 
.A(n_535),
.B(n_177),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_SL g667 ( 
.A(n_488),
.B(n_177),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_472),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_481),
.B(n_413),
.Y(n_669)
);

O2A1O1Ixp33_ASAP7_75t_L g670 ( 
.A1(n_481),
.A2(n_365),
.B(n_380),
.C(n_378),
.Y(n_670)
);

NOR2xp33_ASAP7_75t_L g671 ( 
.A(n_535),
.B(n_265),
.Y(n_671)
);

INVx2_ASAP7_75t_SL g672 ( 
.A(n_463),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_482),
.B(n_413),
.Y(n_673)
);

INVx2_ASAP7_75t_L g674 ( 
.A(n_565),
.Y(n_674)
);

INVx3_ASAP7_75t_L g675 ( 
.A(n_466),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_SL g676 ( 
.A(n_470),
.B(n_265),
.Y(n_676)
);

AND2x2_ASAP7_75t_SL g677 ( 
.A(n_510),
.B(n_366),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_L g678 ( 
.A(n_482),
.B(n_413),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_484),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_SL g680 ( 
.A(n_581),
.B(n_254),
.Y(n_680)
);

OR2x2_ASAP7_75t_L g681 ( 
.A(n_494),
.B(n_366),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_SL g682 ( 
.A(n_559),
.B(n_543),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_484),
.B(n_413),
.Y(n_683)
);

AOI22xp5_ASAP7_75t_L g684 ( 
.A1(n_465),
.A2(n_256),
.B1(n_257),
.B2(n_295),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_486),
.Y(n_685)
);

BUFx6f_ASAP7_75t_L g686 ( 
.A(n_581),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_486),
.Y(n_687)
);

OAI22xp5_ASAP7_75t_L g688 ( 
.A1(n_465),
.A2(n_279),
.B1(n_267),
.B2(n_274),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_SL g689 ( 
.A(n_544),
.B(n_267),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_512),
.B(n_413),
.Y(n_690)
);

NAND2xp33_ASAP7_75t_L g691 ( 
.A(n_592),
.B(n_580),
.Y(n_691)
);

AND2x6_ASAP7_75t_L g692 ( 
.A(n_483),
.B(n_367),
.Y(n_692)
);

NAND2xp33_ASAP7_75t_L g693 ( 
.A(n_508),
.B(n_274),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_512),
.Y(n_694)
);

AO22x2_ASAP7_75t_L g695 ( 
.A1(n_501),
.A2(n_380),
.B1(n_376),
.B2(n_372),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_SL g696 ( 
.A(n_457),
.B(n_279),
.Y(n_696)
);

OAI22xp5_ASAP7_75t_SL g697 ( 
.A1(n_556),
.A2(n_281),
.B1(n_278),
.B2(n_276),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_SL g698 ( 
.A(n_515),
.B(n_288),
.Y(n_698)
);

AOI221xp5_ASAP7_75t_L g699 ( 
.A1(n_508),
.A2(n_275),
.B1(n_211),
.B2(n_210),
.C(n_203),
.Y(n_699)
);

BUFx2_ASAP7_75t_L g700 ( 
.A(n_556),
.Y(n_700)
);

AO22x2_ASAP7_75t_L g701 ( 
.A1(n_508),
.A2(n_372),
.B1(n_370),
.B2(n_367),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_L g702 ( 
.A(n_515),
.B(n_446),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_L g703 ( 
.A(n_517),
.B(n_446),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_L g704 ( 
.A(n_517),
.B(n_446),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_520),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_520),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_522),
.B(n_446),
.Y(n_707)
);

AOI22xp33_ASAP7_75t_L g708 ( 
.A1(n_508),
.A2(n_264),
.B1(n_189),
.B2(n_194),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_522),
.B(n_288),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_L g710 ( 
.A(n_526),
.B(n_289),
.Y(n_710)
);

AOI22xp5_ASAP7_75t_L g711 ( 
.A1(n_535),
.A2(n_289),
.B1(n_290),
.B2(n_295),
.Y(n_711)
);

AND2x2_ASAP7_75t_L g712 ( 
.A(n_473),
.B(n_338),
.Y(n_712)
);

AND2x4_ASAP7_75t_L g713 ( 
.A(n_570),
.B(n_339),
.Y(n_713)
);

INVxp67_ASAP7_75t_L g714 ( 
.A(n_588),
.Y(n_714)
);

INVx2_ASAP7_75t_L g715 ( 
.A(n_589),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_526),
.Y(n_716)
);

NAND2xp33_ASAP7_75t_L g717 ( 
.A(n_529),
.B(n_290),
.Y(n_717)
);

AOI22xp5_ASAP7_75t_SL g718 ( 
.A1(n_531),
.A2(n_183),
.B1(n_196),
.B2(n_197),
.Y(n_718)
);

NOR2xp33_ASAP7_75t_L g719 ( 
.A(n_500),
.B(n_299),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_530),
.B(n_299),
.Y(n_720)
);

AOI21x1_ASAP7_75t_L g721 ( 
.A1(n_567),
.A2(n_345),
.B(n_350),
.Y(n_721)
);

NOR3xp33_ASAP7_75t_L g722 ( 
.A(n_577),
.B(n_303),
.C(n_213),
.Y(n_722)
);

BUFx6f_ASAP7_75t_SL g723 ( 
.A(n_500),
.Y(n_723)
);

OAI22x1_ASAP7_75t_SL g724 ( 
.A1(n_500),
.A2(n_200),
.B1(n_219),
.B2(n_227),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_530),
.Y(n_725)
);

AND2x2_ASAP7_75t_SL g726 ( 
.A(n_510),
.B(n_339),
.Y(n_726)
);

INVx2_ASAP7_75t_L g727 ( 
.A(n_593),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_532),
.Y(n_728)
);

INVx3_ASAP7_75t_L g729 ( 
.A(n_570),
.Y(n_729)
);

HB1xp67_ASAP7_75t_L g730 ( 
.A(n_570),
.Y(n_730)
);

INVxp67_ASAP7_75t_L g731 ( 
.A(n_570),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_533),
.B(n_397),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_L g733 ( 
.A(n_533),
.B(n_397),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_L g734 ( 
.A(n_539),
.B(n_540),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_SL g735 ( 
.A(n_539),
.B(n_233),
.Y(n_735)
);

BUFx5_ASAP7_75t_L g736 ( 
.A(n_564),
.Y(n_736)
);

INVx2_ASAP7_75t_L g737 ( 
.A(n_595),
.Y(n_737)
);

AOI22xp5_ASAP7_75t_L g738 ( 
.A1(n_534),
.A2(n_236),
.B1(n_237),
.B2(n_241),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_SL g739 ( 
.A(n_540),
.B(n_260),
.Y(n_739)
);

BUFx2_ASAP7_75t_L g740 ( 
.A(n_537),
.Y(n_740)
);

INVx2_ASAP7_75t_L g741 ( 
.A(n_595),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_SL g742 ( 
.A(n_541),
.B(n_342),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_L g743 ( 
.A(n_541),
.B(n_546),
.Y(n_743)
);

NOR3xp33_ASAP7_75t_L g744 ( 
.A(n_546),
.B(n_342),
.C(n_343),
.Y(n_744)
);

CKINVDCx20_ASAP7_75t_R g745 ( 
.A(n_598),
.Y(n_745)
);

INVx2_ASAP7_75t_SL g746 ( 
.A(n_594),
.Y(n_746)
);

AOI22xp5_ASAP7_75t_L g747 ( 
.A1(n_534),
.A2(n_350),
.B1(n_348),
.B2(n_346),
.Y(n_747)
);

INVx2_ASAP7_75t_SL g748 ( 
.A(n_594),
.Y(n_748)
);

NOR2xp33_ASAP7_75t_L g749 ( 
.A(n_547),
.B(n_7),
.Y(n_749)
);

OAI221xp5_ASAP7_75t_L g750 ( 
.A1(n_547),
.A2(n_549),
.B1(n_536),
.B2(n_545),
.C(n_548),
.Y(n_750)
);

INVx2_ASAP7_75t_SL g751 ( 
.A(n_549),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_536),
.Y(n_752)
);

AND2x2_ASAP7_75t_L g753 ( 
.A(n_538),
.B(n_343),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_SL g754 ( 
.A(n_538),
.B(n_345),
.Y(n_754)
);

NOR2xp33_ASAP7_75t_SL g755 ( 
.A(n_534),
.B(n_348),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_SL g756 ( 
.A(n_545),
.B(n_346),
.Y(n_756)
);

INVx2_ASAP7_75t_L g757 ( 
.A(n_596),
.Y(n_757)
);

A2O1A1Ixp33_ASAP7_75t_L g758 ( 
.A1(n_548),
.A2(n_13),
.B(n_14),
.C(n_20),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_586),
.Y(n_759)
);

INVx2_ASAP7_75t_L g760 ( 
.A(n_752),
.Y(n_760)
);

INVx5_ASAP7_75t_L g761 ( 
.A(n_686),
.Y(n_761)
);

BUFx12f_ASAP7_75t_L g762 ( 
.A(n_655),
.Y(n_762)
);

AOI22xp33_ASAP7_75t_L g763 ( 
.A1(n_691),
.A2(n_518),
.B1(n_523),
.B2(n_509),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_599),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_L g765 ( 
.A(n_686),
.B(n_483),
.Y(n_765)
);

O2A1O1Ixp33_ASAP7_75t_L g766 ( 
.A1(n_693),
.A2(n_661),
.B(n_620),
.C(n_749),
.Y(n_766)
);

NOR3xp33_ASAP7_75t_SL g767 ( 
.A(n_638),
.B(n_591),
.C(n_583),
.Y(n_767)
);

INVx2_ASAP7_75t_L g768 ( 
.A(n_607),
.Y(n_768)
);

INVxp67_ASAP7_75t_SL g769 ( 
.A(n_686),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_L g770 ( 
.A(n_686),
.B(n_504),
.Y(n_770)
);

INVx2_ASAP7_75t_L g771 ( 
.A(n_612),
.Y(n_771)
);

NOR2xp33_ASAP7_75t_L g772 ( 
.A(n_602),
.B(n_469),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_653),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_L g774 ( 
.A(n_603),
.B(n_504),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_662),
.Y(n_775)
);

OAI22xp5_ASAP7_75t_L g776 ( 
.A1(n_654),
.A2(n_477),
.B1(n_479),
.B2(n_474),
.Y(n_776)
);

INVx3_ASAP7_75t_L g777 ( 
.A(n_649),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_L g778 ( 
.A(n_603),
.B(n_509),
.Y(n_778)
);

CKINVDCx5p33_ASAP7_75t_R g779 ( 
.A(n_658),
.Y(n_779)
);

INVx6_ASAP7_75t_L g780 ( 
.A(n_626),
.Y(n_780)
);

AOI22xp33_ASAP7_75t_L g781 ( 
.A1(n_654),
.A2(n_527),
.B1(n_518),
.B2(n_523),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_L g782 ( 
.A(n_603),
.B(n_527),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_668),
.Y(n_783)
);

NAND2xp33_ASAP7_75t_SL g784 ( 
.A(n_723),
.B(n_516),
.Y(n_784)
);

BUFx6f_ASAP7_75t_L g785 ( 
.A(n_649),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_L g786 ( 
.A(n_603),
.B(n_453),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_L g787 ( 
.A(n_603),
.B(n_453),
.Y(n_787)
);

INVx2_ASAP7_75t_SL g788 ( 
.A(n_664),
.Y(n_788)
);

AOI22xp5_ASAP7_75t_L g789 ( 
.A1(n_639),
.A2(n_597),
.B1(n_459),
.B2(n_460),
.Y(n_789)
);

NAND2x1p5_ASAP7_75t_L g790 ( 
.A(n_729),
.B(n_511),
.Y(n_790)
);

INVx2_ASAP7_75t_L g791 ( 
.A(n_605),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_746),
.B(n_459),
.Y(n_792)
);

AND2x4_ASAP7_75t_L g793 ( 
.A(n_647),
.B(n_459),
.Y(n_793)
);

AOI22xp5_ASAP7_75t_L g794 ( 
.A1(n_639),
.A2(n_597),
.B1(n_460),
.B2(n_461),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_679),
.Y(n_795)
);

AND2x4_ASAP7_75t_L g796 ( 
.A(n_648),
.B(n_460),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_748),
.B(n_461),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_685),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_SL g799 ( 
.A(n_755),
.B(n_511),
.Y(n_799)
);

INVx2_ASAP7_75t_L g800 ( 
.A(n_606),
.Y(n_800)
);

HB1xp67_ASAP7_75t_L g801 ( 
.A(n_657),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_687),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_694),
.Y(n_803)
);

INVx2_ASAP7_75t_L g804 ( 
.A(n_616),
.Y(n_804)
);

INVx2_ASAP7_75t_L g805 ( 
.A(n_628),
.Y(n_805)
);

NOR2xp33_ASAP7_75t_R g806 ( 
.A(n_665),
.B(n_745),
.Y(n_806)
);

BUFx6f_ASAP7_75t_L g807 ( 
.A(n_649),
.Y(n_807)
);

INVx2_ASAP7_75t_L g808 ( 
.A(n_636),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_SL g809 ( 
.A(n_603),
.B(n_511),
.Y(n_809)
);

CKINVDCx5p33_ASAP7_75t_R g810 ( 
.A(n_601),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_705),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_SL g812 ( 
.A(n_649),
.B(n_511),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_SL g813 ( 
.A(n_751),
.B(n_516),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_L g814 ( 
.A(n_734),
.B(n_454),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_706),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_716),
.Y(n_816)
);

AND2x4_ASAP7_75t_L g817 ( 
.A(n_713),
.B(n_461),
.Y(n_817)
);

BUFx2_ASAP7_75t_L g818 ( 
.A(n_740),
.Y(n_818)
);

NOR2xp33_ASAP7_75t_L g819 ( 
.A(n_602),
.B(n_469),
.Y(n_819)
);

NOR2xp33_ASAP7_75t_L g820 ( 
.A(n_657),
.B(n_469),
.Y(n_820)
);

BUFx3_ASAP7_75t_L g821 ( 
.A(n_700),
.Y(n_821)
);

NOR2xp33_ASAP7_75t_L g822 ( 
.A(n_714),
.B(n_491),
.Y(n_822)
);

INVx2_ASAP7_75t_L g823 ( 
.A(n_637),
.Y(n_823)
);

OAI21xp33_ASAP7_75t_L g824 ( 
.A1(n_614),
.A2(n_558),
.B(n_464),
.Y(n_824)
);

BUFx6f_ASAP7_75t_L g825 ( 
.A(n_729),
.Y(n_825)
);

BUFx2_ASAP7_75t_L g826 ( 
.A(n_652),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_L g827 ( 
.A(n_743),
.B(n_454),
.Y(n_827)
);

INVx1_ASAP7_75t_SL g828 ( 
.A(n_611),
.Y(n_828)
);

HB1xp67_ASAP7_75t_L g829 ( 
.A(n_644),
.Y(n_829)
);

OR2x6_ASAP7_75t_L g830 ( 
.A(n_621),
.B(n_627),
.Y(n_830)
);

INVx2_ASAP7_75t_L g831 ( 
.A(n_641),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_SL g832 ( 
.A(n_629),
.B(n_516),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_725),
.B(n_464),
.Y(n_833)
);

OAI21xp5_ASAP7_75t_L g834 ( 
.A1(n_661),
.A2(n_479),
.B(n_477),
.Y(n_834)
);

NOR2xp67_ASAP7_75t_L g835 ( 
.A(n_714),
.B(n_474),
.Y(n_835)
);

BUFx3_ASAP7_75t_L g836 ( 
.A(n_672),
.Y(n_836)
);

AND2x4_ASAP7_75t_L g837 ( 
.A(n_713),
.B(n_490),
.Y(n_837)
);

HB1xp67_ASAP7_75t_L g838 ( 
.A(n_730),
.Y(n_838)
);

AND2x6_ASAP7_75t_L g839 ( 
.A(n_712),
.B(n_490),
.Y(n_839)
);

INVx2_ASAP7_75t_L g840 ( 
.A(n_660),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_728),
.Y(n_841)
);

OAI22xp5_ASAP7_75t_L g842 ( 
.A1(n_708),
.A2(n_571),
.B1(n_591),
.B2(n_568),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_610),
.B(n_499),
.Y(n_843)
);

BUFx4f_ASAP7_75t_SL g844 ( 
.A(n_663),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_753),
.Y(n_845)
);

BUFx2_ASAP7_75t_L g846 ( 
.A(n_695),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_L g847 ( 
.A(n_675),
.B(n_499),
.Y(n_847)
);

AND2x4_ASAP7_75t_L g848 ( 
.A(n_730),
.B(n_551),
.Y(n_848)
);

INVx2_ASAP7_75t_SL g849 ( 
.A(n_630),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_759),
.Y(n_850)
);

NAND2x1p5_ASAP7_75t_L g851 ( 
.A(n_675),
.B(n_491),
.Y(n_851)
);

INVx4_ASAP7_75t_L g852 ( 
.A(n_692),
.Y(n_852)
);

BUFx6f_ASAP7_75t_L g853 ( 
.A(n_692),
.Y(n_853)
);

INVx1_ASAP7_75t_SL g854 ( 
.A(n_681),
.Y(n_854)
);

BUFx2_ASAP7_75t_L g855 ( 
.A(n_695),
.Y(n_855)
);

INVx4_ASAP7_75t_L g856 ( 
.A(n_692),
.Y(n_856)
);

INVx1_ASAP7_75t_SL g857 ( 
.A(n_709),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_650),
.Y(n_858)
);

INVx2_ASAP7_75t_SL g859 ( 
.A(n_608),
.Y(n_859)
);

AOI22xp5_ASAP7_75t_L g860 ( 
.A1(n_629),
.A2(n_551),
.B1(n_590),
.B2(n_587),
.Y(n_860)
);

INVxp67_ASAP7_75t_L g861 ( 
.A(n_614),
.Y(n_861)
);

NOR2xp33_ASAP7_75t_L g862 ( 
.A(n_651),
.B(n_491),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_656),
.Y(n_863)
);

INVx3_ASAP7_75t_L g864 ( 
.A(n_692),
.Y(n_864)
);

INVx2_ASAP7_75t_L g865 ( 
.A(n_674),
.Y(n_865)
);

OR2x2_ASAP7_75t_L g866 ( 
.A(n_615),
.B(n_14),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_633),
.B(n_551),
.Y(n_867)
);

INVxp67_ASAP7_75t_SL g868 ( 
.A(n_736),
.Y(n_868)
);

INVx2_ASAP7_75t_SL g869 ( 
.A(n_735),
.Y(n_869)
);

BUFx6f_ASAP7_75t_SL g870 ( 
.A(n_604),
.Y(n_870)
);

OR2x6_ASAP7_75t_L g871 ( 
.A(n_604),
.B(n_529),
.Y(n_871)
);

AOI22xp33_ASAP7_75t_L g872 ( 
.A1(n_622),
.A2(n_529),
.B1(n_572),
.B2(n_564),
.Y(n_872)
);

INVx3_ASAP7_75t_L g873 ( 
.A(n_692),
.Y(n_873)
);

NOR2xp33_ASAP7_75t_L g874 ( 
.A(n_651),
.B(n_521),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_SL g875 ( 
.A(n_633),
.B(n_516),
.Y(n_875)
);

AOI22xp33_ASAP7_75t_L g876 ( 
.A1(n_622),
.A2(n_529),
.B1(n_572),
.B2(n_568),
.Y(n_876)
);

BUFx6f_ASAP7_75t_L g877 ( 
.A(n_677),
.Y(n_877)
);

NOR2xp33_ASAP7_75t_L g878 ( 
.A(n_666),
.B(n_521),
.Y(n_878)
);

HB1xp67_ASAP7_75t_L g879 ( 
.A(n_731),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_L g880 ( 
.A(n_635),
.B(n_613),
.Y(n_880)
);

NOR2xp33_ASAP7_75t_SL g881 ( 
.A(n_601),
.B(n_569),
.Y(n_881)
);

INVx2_ASAP7_75t_SL g882 ( 
.A(n_739),
.Y(n_882)
);

AOI22xp5_ASAP7_75t_L g883 ( 
.A1(n_634),
.A2(n_590),
.B1(n_587),
.B2(n_585),
.Y(n_883)
);

AOI22xp5_ASAP7_75t_L g884 ( 
.A1(n_634),
.A2(n_590),
.B1(n_587),
.B2(n_585),
.Y(n_884)
);

AND2x2_ASAP7_75t_L g885 ( 
.A(n_666),
.B(n_596),
.Y(n_885)
);

NAND3xp33_ASAP7_75t_SL g886 ( 
.A(n_722),
.B(n_571),
.C(n_573),
.Y(n_886)
);

AOI22xp5_ASAP7_75t_L g887 ( 
.A1(n_680),
.A2(n_585),
.B1(n_521),
.B2(n_569),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_SL g888 ( 
.A(n_643),
.B(n_516),
.Y(n_888)
);

BUFx2_ASAP7_75t_L g889 ( 
.A(n_695),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_669),
.Y(n_890)
);

NAND3xp33_ASAP7_75t_SL g891 ( 
.A(n_722),
.B(n_573),
.C(n_575),
.Y(n_891)
);

INVx4_ASAP7_75t_L g892 ( 
.A(n_624),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_673),
.Y(n_893)
);

NOR2xp33_ASAP7_75t_L g894 ( 
.A(n_671),
.B(n_569),
.Y(n_894)
);

AND2x4_ASAP7_75t_L g895 ( 
.A(n_731),
.B(n_584),
.Y(n_895)
);

AND2x6_ASAP7_75t_L g896 ( 
.A(n_749),
.B(n_584),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_678),
.Y(n_897)
);

AND2x4_ASAP7_75t_L g898 ( 
.A(n_618),
.B(n_584),
.Y(n_898)
);

BUFx4f_ASAP7_75t_L g899 ( 
.A(n_604),
.Y(n_899)
);

AND2x4_ASAP7_75t_L g900 ( 
.A(n_747),
.B(n_584),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_683),
.Y(n_901)
);

INVx4_ASAP7_75t_L g902 ( 
.A(n_624),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_SL g903 ( 
.A(n_638),
.B(n_525),
.Y(n_903)
);

OAI22xp5_ASAP7_75t_L g904 ( 
.A1(n_708),
.A2(n_582),
.B1(n_576),
.B2(n_575),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_L g905 ( 
.A(n_710),
.B(n_525),
.Y(n_905)
);

INVx2_ASAP7_75t_SL g906 ( 
.A(n_609),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_690),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_754),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_754),
.Y(n_909)
);

INVxp67_ASAP7_75t_L g910 ( 
.A(n_667),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_756),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_SL g912 ( 
.A(n_659),
.B(n_719),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_L g913 ( 
.A(n_720),
.B(n_525),
.Y(n_913)
);

BUFx6f_ASAP7_75t_L g914 ( 
.A(n_677),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_L g915 ( 
.A(n_609),
.B(n_525),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_756),
.Y(n_916)
);

AOI22xp33_ASAP7_75t_L g917 ( 
.A1(n_609),
.A2(n_558),
.B1(n_525),
.B2(n_397),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_SL g918 ( 
.A(n_719),
.B(n_75),
.Y(n_918)
);

NOR2xp33_ASAP7_75t_R g919 ( 
.A(n_600),
.B(n_78),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_645),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_L g921 ( 
.A(n_640),
.B(n_397),
.Y(n_921)
);

NOR3xp33_ASAP7_75t_SL g922 ( 
.A(n_632),
.B(n_20),
.C(n_22),
.Y(n_922)
);

NAND2x1p5_ASAP7_75t_L g923 ( 
.A(n_742),
.B(n_79),
.Y(n_923)
);

A2O1A1Ixp33_ASAP7_75t_L g924 ( 
.A1(n_699),
.A2(n_23),
.B(n_26),
.C(n_27),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_715),
.Y(n_925)
);

OAI21xp5_ASAP7_75t_L g926 ( 
.A1(n_646),
.A2(n_397),
.B(n_84),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_L g927 ( 
.A(n_617),
.B(n_80),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_L g928 ( 
.A(n_619),
.B(n_71),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_L g929 ( 
.A(n_623),
.B(n_59),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_631),
.B(n_736),
.Y(n_930)
);

AOI22xp33_ASAP7_75t_L g931 ( 
.A1(n_701),
.A2(n_26),
.B1(n_32),
.B2(n_33),
.Y(n_931)
);

INVx2_ASAP7_75t_SL g932 ( 
.A(n_698),
.Y(n_932)
);

INVx1_ASAP7_75t_L g933 ( 
.A(n_727),
.Y(n_933)
);

NAND3xp33_ASAP7_75t_SL g934 ( 
.A(n_711),
.B(n_34),
.C(n_36),
.Y(n_934)
);

NOR2xp33_ASAP7_75t_L g935 ( 
.A(n_676),
.B(n_38),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_737),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_L g937 ( 
.A(n_736),
.B(n_106),
.Y(n_937)
);

AOI222xp33_ASAP7_75t_L g938 ( 
.A1(n_861),
.A2(n_724),
.B1(n_697),
.B2(n_723),
.C1(n_689),
.C2(n_696),
.Y(n_938)
);

AOI21xp5_ASAP7_75t_L g939 ( 
.A1(n_930),
.A2(n_717),
.B(n_750),
.Y(n_939)
);

AOI21xp5_ASAP7_75t_L g940 ( 
.A1(n_930),
.A2(n_704),
.B(n_703),
.Y(n_940)
);

O2A1O1Ixp33_ASAP7_75t_L g941 ( 
.A1(n_912),
.A2(n_758),
.B(n_625),
.C(n_642),
.Y(n_941)
);

AOI21xp5_ASAP7_75t_L g942 ( 
.A1(n_761),
.A2(n_707),
.B(n_702),
.Y(n_942)
);

AO21x1_ASAP7_75t_L g943 ( 
.A1(n_766),
.A2(n_733),
.B(n_732),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_L g944 ( 
.A(n_857),
.B(n_701),
.Y(n_944)
);

AOI21xp5_ASAP7_75t_L g945 ( 
.A1(n_761),
.A2(n_726),
.B(n_757),
.Y(n_945)
);

O2A1O1Ixp33_ASAP7_75t_L g946 ( 
.A1(n_924),
.A2(n_670),
.B(n_688),
.C(n_744),
.Y(n_946)
);

O2A1O1Ixp33_ASAP7_75t_SL g947 ( 
.A1(n_918),
.A2(n_684),
.B(n_741),
.C(n_738),
.Y(n_947)
);

O2A1O1Ixp5_ASAP7_75t_L g948 ( 
.A1(n_772),
.A2(n_721),
.B(n_646),
.C(n_736),
.Y(n_948)
);

INVx2_ASAP7_75t_SL g949 ( 
.A(n_818),
.Y(n_949)
);

OAI22xp5_ASAP7_75t_SL g950 ( 
.A1(n_844),
.A2(n_726),
.B1(n_718),
.B2(n_44),
.Y(n_950)
);

AOI21xp5_ASAP7_75t_L g951 ( 
.A1(n_761),
.A2(n_736),
.B(n_670),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_773),
.Y(n_952)
);

INVx2_ASAP7_75t_L g953 ( 
.A(n_768),
.Y(n_953)
);

NAND3xp33_ASAP7_75t_SL g954 ( 
.A(n_857),
.B(n_744),
.C(n_41),
.Y(n_954)
);

NOR2xp33_ASAP7_75t_L g955 ( 
.A(n_828),
.B(n_736),
.Y(n_955)
);

AOI22xp5_ASAP7_75t_L g956 ( 
.A1(n_826),
.A2(n_107),
.B1(n_140),
.B2(n_137),
.Y(n_956)
);

INVx1_ASAP7_75t_SL g957 ( 
.A(n_828),
.Y(n_957)
);

INVx3_ASAP7_75t_L g958 ( 
.A(n_785),
.Y(n_958)
);

BUFx2_ASAP7_75t_L g959 ( 
.A(n_821),
.Y(n_959)
);

NOR2xp67_ASAP7_75t_L g960 ( 
.A(n_779),
.B(n_788),
.Y(n_960)
);

AND2x4_ASAP7_75t_L g961 ( 
.A(n_830),
.B(n_62),
.Y(n_961)
);

AND2x2_ASAP7_75t_L g962 ( 
.A(n_854),
.B(n_39),
.Y(n_962)
);

NOR2xp33_ASAP7_75t_R g963 ( 
.A(n_784),
.B(n_104),
.Y(n_963)
);

INVx3_ASAP7_75t_L g964 ( 
.A(n_785),
.Y(n_964)
);

INVx2_ASAP7_75t_L g965 ( 
.A(n_771),
.Y(n_965)
);

OAI22xp5_ASAP7_75t_L g966 ( 
.A1(n_877),
.A2(n_914),
.B1(n_846),
.B2(n_855),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_L g967 ( 
.A(n_880),
.B(n_44),
.Y(n_967)
);

CKINVDCx6p67_ASAP7_75t_R g968 ( 
.A(n_762),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_L g969 ( 
.A(n_920),
.B(n_45),
.Y(n_969)
);

A2O1A1Ixp33_ASAP7_75t_L g970 ( 
.A1(n_935),
.A2(n_45),
.B(n_46),
.C(n_48),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_L g971 ( 
.A(n_845),
.B(n_108),
.Y(n_971)
);

OAI22x1_ASAP7_75t_L g972 ( 
.A1(n_889),
.A2(n_116),
.B1(n_126),
.B2(n_146),
.Y(n_972)
);

BUFx12f_ASAP7_75t_L g973 ( 
.A(n_892),
.Y(n_973)
);

BUFx6f_ASAP7_75t_L g974 ( 
.A(n_785),
.Y(n_974)
);

AND2x2_ASAP7_75t_L g975 ( 
.A(n_854),
.B(n_829),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_L g976 ( 
.A(n_885),
.B(n_819),
.Y(n_976)
);

AOI21xp5_ASAP7_75t_L g977 ( 
.A1(n_786),
.A2(n_787),
.B(n_868),
.Y(n_977)
);

NOR2xp33_ASAP7_75t_L g978 ( 
.A(n_801),
.B(n_849),
.Y(n_978)
);

NAND3xp33_ASAP7_75t_SL g979 ( 
.A(n_806),
.B(n_922),
.C(n_866),
.Y(n_979)
);

AOI21xp5_ASAP7_75t_L g980 ( 
.A1(n_787),
.A2(n_778),
.B(n_774),
.Y(n_980)
);

OAI21x1_ASAP7_75t_L g981 ( 
.A1(n_774),
.A2(n_782),
.B(n_778),
.Y(n_981)
);

INVx1_ASAP7_75t_SL g982 ( 
.A(n_838),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_SL g983 ( 
.A(n_877),
.B(n_914),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_SL g984 ( 
.A(n_877),
.B(n_914),
.Y(n_984)
);

OAI22xp5_ASAP7_75t_L g985 ( 
.A1(n_931),
.A2(n_906),
.B1(n_899),
.B2(n_767),
.Y(n_985)
);

NOR2xp33_ASAP7_75t_L g986 ( 
.A(n_879),
.B(n_910),
.Y(n_986)
);

OAI22xp5_ASAP7_75t_SL g987 ( 
.A1(n_810),
.A2(n_859),
.B1(n_932),
.B2(n_869),
.Y(n_987)
);

INVx2_ASAP7_75t_L g988 ( 
.A(n_760),
.Y(n_988)
);

AOI21xp5_ASAP7_75t_L g989 ( 
.A1(n_782),
.A2(n_913),
.B(n_905),
.Y(n_989)
);

O2A1O1Ixp33_ASAP7_75t_SL g990 ( 
.A1(n_937),
.A2(n_903),
.B(n_928),
.C(n_927),
.Y(n_990)
);

NOR2xp33_ASAP7_75t_L g991 ( 
.A(n_882),
.B(n_820),
.Y(n_991)
);

INVx2_ASAP7_75t_L g992 ( 
.A(n_791),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_775),
.Y(n_993)
);

O2A1O1Ixp5_ASAP7_75t_L g994 ( 
.A1(n_888),
.A2(n_832),
.B(n_875),
.C(n_894),
.Y(n_994)
);

AOI21xp5_ASAP7_75t_L g995 ( 
.A1(n_814),
.A2(n_827),
.B(n_765),
.Y(n_995)
);

OAI22xp5_ASAP7_75t_L g996 ( 
.A1(n_899),
.A2(n_803),
.B1(n_811),
.B2(n_841),
.Y(n_996)
);

NOR2xp33_ASAP7_75t_L g997 ( 
.A(n_783),
.B(n_795),
.Y(n_997)
);

OR2x6_ASAP7_75t_L g998 ( 
.A(n_780),
.B(n_892),
.Y(n_998)
);

OAI22xp5_ASAP7_75t_L g999 ( 
.A1(n_798),
.A2(n_815),
.B1(n_802),
.B2(n_816),
.Y(n_999)
);

INVx1_ASAP7_75t_L g1000 ( 
.A(n_764),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_L g1001 ( 
.A(n_862),
.B(n_874),
.Y(n_1001)
);

CKINVDCx5p33_ASAP7_75t_R g1002 ( 
.A(n_780),
.Y(n_1002)
);

AOI21xp5_ASAP7_75t_L g1003 ( 
.A1(n_765),
.A2(n_770),
.B(n_843),
.Y(n_1003)
);

OR2x2_ASAP7_75t_L g1004 ( 
.A(n_850),
.B(n_836),
.Y(n_1004)
);

BUFx3_ASAP7_75t_L g1005 ( 
.A(n_830),
.Y(n_1005)
);

INVx2_ASAP7_75t_L g1006 ( 
.A(n_800),
.Y(n_1006)
);

BUFx6f_ASAP7_75t_L g1007 ( 
.A(n_807),
.Y(n_1007)
);

NOR2xp33_ASAP7_75t_R g1008 ( 
.A(n_881),
.B(n_886),
.Y(n_1008)
);

OAI21xp33_ASAP7_75t_L g1009 ( 
.A1(n_934),
.A2(n_878),
.B(n_830),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_L g1010 ( 
.A(n_822),
.B(n_835),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_SL g1011 ( 
.A(n_825),
.B(n_881),
.Y(n_1011)
);

AOI21xp5_ASAP7_75t_L g1012 ( 
.A1(n_843),
.A2(n_867),
.B(n_809),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_L g1013 ( 
.A(n_858),
.B(n_863),
.Y(n_1013)
);

A2O1A1Ixp33_ASAP7_75t_L g1014 ( 
.A1(n_908),
.A2(n_911),
.B(n_909),
.C(n_916),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_833),
.Y(n_1015)
);

OAI21x1_ASAP7_75t_L g1016 ( 
.A1(n_834),
.A2(n_763),
.B(n_847),
.Y(n_1016)
);

INVx5_ASAP7_75t_L g1017 ( 
.A(n_853),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_SL g1018 ( 
.A(n_825),
.B(n_807),
.Y(n_1018)
);

NOR2xp67_ASAP7_75t_L g1019 ( 
.A(n_902),
.B(n_891),
.Y(n_1019)
);

AOI22xp33_ASAP7_75t_L g1020 ( 
.A1(n_793),
.A2(n_796),
.B1(n_837),
.B2(n_817),
.Y(n_1020)
);

INVx2_ASAP7_75t_SL g1021 ( 
.A(n_848),
.Y(n_1021)
);

INVx1_ASAP7_75t_L g1022 ( 
.A(n_833),
.Y(n_1022)
);

AOI22xp5_ASAP7_75t_L g1023 ( 
.A1(n_817),
.A2(n_837),
.B1(n_848),
.B2(n_895),
.Y(n_1023)
);

INVx4_ASAP7_75t_L g1024 ( 
.A(n_807),
.Y(n_1024)
);

INVx1_ASAP7_75t_L g1025 ( 
.A(n_925),
.Y(n_1025)
);

INVx2_ASAP7_75t_SL g1026 ( 
.A(n_825),
.Y(n_1026)
);

OAI21xp5_ASAP7_75t_L g1027 ( 
.A1(n_926),
.A2(n_834),
.B(n_776),
.Y(n_1027)
);

INVx1_ASAP7_75t_L g1028 ( 
.A(n_933),
.Y(n_1028)
);

INVx2_ASAP7_75t_L g1029 ( 
.A(n_804),
.Y(n_1029)
);

CKINVDCx5p33_ASAP7_75t_R g1030 ( 
.A(n_902),
.Y(n_1030)
);

INVx2_ASAP7_75t_L g1031 ( 
.A(n_805),
.Y(n_1031)
);

INVx1_ASAP7_75t_L g1032 ( 
.A(n_936),
.Y(n_1032)
);

NAND2xp5_ASAP7_75t_L g1033 ( 
.A(n_890),
.B(n_893),
.Y(n_1033)
);

INVx4_ASAP7_75t_L g1034 ( 
.A(n_777),
.Y(n_1034)
);

INVx2_ASAP7_75t_L g1035 ( 
.A(n_808),
.Y(n_1035)
);

OAI22xp5_ASAP7_75t_L g1036 ( 
.A1(n_871),
.A2(n_926),
.B1(n_915),
.B2(n_900),
.Y(n_1036)
);

INVx5_ASAP7_75t_L g1037 ( 
.A(n_853),
.Y(n_1037)
);

CKINVDCx20_ASAP7_75t_R g1038 ( 
.A(n_919),
.Y(n_1038)
);

BUFx2_ASAP7_75t_L g1039 ( 
.A(n_895),
.Y(n_1039)
);

NAND2xp5_ASAP7_75t_L g1040 ( 
.A(n_897),
.B(n_907),
.Y(n_1040)
);

NAND2xp5_ASAP7_75t_SL g1041 ( 
.A(n_793),
.B(n_796),
.Y(n_1041)
);

NOR2xp33_ASAP7_75t_R g1042 ( 
.A(n_777),
.B(n_864),
.Y(n_1042)
);

INVx1_ASAP7_75t_L g1043 ( 
.A(n_823),
.Y(n_1043)
);

INVx1_ASAP7_75t_SL g1044 ( 
.A(n_792),
.Y(n_1044)
);

INVx4_ASAP7_75t_L g1045 ( 
.A(n_839),
.Y(n_1045)
);

OAI22xp5_ASAP7_75t_L g1046 ( 
.A1(n_871),
.A2(n_900),
.B1(n_937),
.B2(n_781),
.Y(n_1046)
);

INVx3_ASAP7_75t_L g1047 ( 
.A(n_853),
.Y(n_1047)
);

O2A1O1Ixp33_ASAP7_75t_L g1048 ( 
.A1(n_842),
.A2(n_904),
.B(n_776),
.C(n_824),
.Y(n_1048)
);

INVx2_ASAP7_75t_L g1049 ( 
.A(n_831),
.Y(n_1049)
);

O2A1O1Ixp33_ASAP7_75t_L g1050 ( 
.A1(n_842),
.A2(n_904),
.B(n_901),
.C(n_797),
.Y(n_1050)
);

BUFx6f_ASAP7_75t_L g1051 ( 
.A(n_839),
.Y(n_1051)
);

INVx1_ASAP7_75t_L g1052 ( 
.A(n_840),
.Y(n_1052)
);

OAI22xp5_ASAP7_75t_L g1053 ( 
.A1(n_917),
.A2(n_769),
.B1(n_876),
.B2(n_872),
.Y(n_1053)
);

AOI21xp5_ASAP7_75t_L g1054 ( 
.A1(n_851),
.A2(n_929),
.B(n_927),
.Y(n_1054)
);

NOR2xp33_ASAP7_75t_L g1055 ( 
.A(n_870),
.B(n_865),
.Y(n_1055)
);

BUFx6f_ASAP7_75t_L g1056 ( 
.A(n_839),
.Y(n_1056)
);

A2O1A1Ixp33_ASAP7_75t_L g1057 ( 
.A1(n_864),
.A2(n_873),
.B(n_789),
.C(n_794),
.Y(n_1057)
);

A2O1A1Ixp33_ASAP7_75t_L g1058 ( 
.A1(n_873),
.A2(n_860),
.B(n_884),
.C(n_883),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_813),
.Y(n_1059)
);

NAND2xp5_ASAP7_75t_SL g1060 ( 
.A(n_898),
.B(n_852),
.Y(n_1060)
);

BUFx2_ASAP7_75t_L g1061 ( 
.A(n_923),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_SL g1062 ( 
.A(n_852),
.B(n_856),
.Y(n_1062)
);

INVx4_ASAP7_75t_L g1063 ( 
.A(n_856),
.Y(n_1063)
);

BUFx6f_ASAP7_75t_L g1064 ( 
.A(n_923),
.Y(n_1064)
);

AOI21xp5_ASAP7_75t_L g1065 ( 
.A1(n_812),
.A2(n_921),
.B(n_887),
.Y(n_1065)
);

INVx1_ASAP7_75t_L g1066 ( 
.A(n_790),
.Y(n_1066)
);

HAxp5_ASAP7_75t_L g1067 ( 
.A(n_896),
.B(n_799),
.CON(n_1067),
.SN(n_1067)
);

INVx2_ASAP7_75t_L g1068 ( 
.A(n_896),
.Y(n_1068)
);

OAI21xp33_ASAP7_75t_L g1069 ( 
.A1(n_828),
.A2(n_485),
.B(n_602),
.Y(n_1069)
);

INVx2_ASAP7_75t_L g1070 ( 
.A(n_768),
.Y(n_1070)
);

INVx2_ASAP7_75t_L g1071 ( 
.A(n_768),
.Y(n_1071)
);

INVx2_ASAP7_75t_L g1072 ( 
.A(n_768),
.Y(n_1072)
);

O2A1O1Ixp5_ASAP7_75t_L g1073 ( 
.A1(n_772),
.A2(n_682),
.B(n_819),
.C(n_912),
.Y(n_1073)
);

NOR2xp33_ASAP7_75t_L g1074 ( 
.A(n_861),
.B(n_485),
.Y(n_1074)
);

A2O1A1Ixp33_ASAP7_75t_L g1075 ( 
.A1(n_1048),
.A2(n_1001),
.B(n_1073),
.C(n_941),
.Y(n_1075)
);

AOI21xp5_ASAP7_75t_L g1076 ( 
.A1(n_1054),
.A2(n_990),
.B(n_989),
.Y(n_1076)
);

AO31x2_ASAP7_75t_L g1077 ( 
.A1(n_943),
.A2(n_1036),
.A3(n_1046),
.B(n_1058),
.Y(n_1077)
);

OAI21x1_ASAP7_75t_L g1078 ( 
.A1(n_981),
.A2(n_1003),
.B(n_980),
.Y(n_1078)
);

OAI21x1_ASAP7_75t_L g1079 ( 
.A1(n_977),
.A2(n_1016),
.B(n_940),
.Y(n_1079)
);

OR2x2_ASAP7_75t_L g1080 ( 
.A(n_957),
.B(n_944),
.Y(n_1080)
);

AOI21xp5_ASAP7_75t_L g1081 ( 
.A1(n_939),
.A2(n_976),
.B(n_1027),
.Y(n_1081)
);

AOI21xp5_ASAP7_75t_L g1082 ( 
.A1(n_1027),
.A2(n_1012),
.B(n_1010),
.Y(n_1082)
);

INVx2_ASAP7_75t_L g1083 ( 
.A(n_993),
.Y(n_1083)
);

BUFx6f_ASAP7_75t_L g1084 ( 
.A(n_974),
.Y(n_1084)
);

INVx3_ASAP7_75t_L g1085 ( 
.A(n_1051),
.Y(n_1085)
);

AOI21xp5_ASAP7_75t_L g1086 ( 
.A1(n_1065),
.A2(n_1050),
.B(n_1046),
.Y(n_1086)
);

INVxp67_ASAP7_75t_L g1087 ( 
.A(n_978),
.Y(n_1087)
);

INVx1_ASAP7_75t_SL g1088 ( 
.A(n_957),
.Y(n_1088)
);

AOI21xp5_ASAP7_75t_L g1089 ( 
.A1(n_1033),
.A2(n_945),
.B(n_1013),
.Y(n_1089)
);

INVx1_ASAP7_75t_L g1090 ( 
.A(n_1000),
.Y(n_1090)
);

OAI21x1_ASAP7_75t_L g1091 ( 
.A1(n_942),
.A2(n_951),
.B(n_948),
.Y(n_1091)
);

AOI21xp5_ASAP7_75t_L g1092 ( 
.A1(n_1040),
.A2(n_1036),
.B(n_1053),
.Y(n_1092)
);

OAI22xp5_ASAP7_75t_L g1093 ( 
.A1(n_1015),
.A2(n_1022),
.B1(n_997),
.B2(n_967),
.Y(n_1093)
);

CKINVDCx5p33_ASAP7_75t_R g1094 ( 
.A(n_959),
.Y(n_1094)
);

AND2x2_ASAP7_75t_L g1095 ( 
.A(n_975),
.B(n_1074),
.Y(n_1095)
);

NAND2xp5_ASAP7_75t_L g1096 ( 
.A(n_1044),
.B(n_955),
.Y(n_1096)
);

AND3x4_ASAP7_75t_L g1097 ( 
.A(n_960),
.B(n_1019),
.C(n_1005),
.Y(n_1097)
);

AOI22xp5_ASAP7_75t_L g1098 ( 
.A1(n_979),
.A2(n_1069),
.B1(n_950),
.B2(n_938),
.Y(n_1098)
);

AOI21xp5_ASAP7_75t_L g1099 ( 
.A1(n_1053),
.A2(n_1060),
.B(n_1062),
.Y(n_1099)
);

AOI21x1_ASAP7_75t_L g1100 ( 
.A1(n_1061),
.A2(n_1011),
.B(n_996),
.Y(n_1100)
);

NAND2xp5_ASAP7_75t_L g1101 ( 
.A(n_1044),
.B(n_969),
.Y(n_1101)
);

NAND2xp5_ASAP7_75t_L g1102 ( 
.A(n_1014),
.B(n_985),
.Y(n_1102)
);

AOI21x1_ASAP7_75t_SL g1103 ( 
.A1(n_961),
.A2(n_971),
.B(n_962),
.Y(n_1103)
);

AOI221x1_ASAP7_75t_L g1104 ( 
.A1(n_1009),
.A2(n_985),
.B1(n_970),
.B2(n_966),
.C(n_996),
.Y(n_1104)
);

INVx1_ASAP7_75t_SL g1105 ( 
.A(n_982),
.Y(n_1105)
);

OAI21xp33_ASAP7_75t_L g1106 ( 
.A1(n_986),
.A2(n_954),
.B(n_938),
.Y(n_1106)
);

AOI21x1_ASAP7_75t_L g1107 ( 
.A1(n_983),
.A2(n_984),
.B(n_999),
.Y(n_1107)
);

OAI21x1_ASAP7_75t_L g1108 ( 
.A1(n_1059),
.A2(n_1047),
.B(n_1066),
.Y(n_1108)
);

AND2x2_ASAP7_75t_L g1109 ( 
.A(n_1021),
.B(n_1039),
.Y(n_1109)
);

AOI221xp5_ASAP7_75t_L g1110 ( 
.A1(n_946),
.A2(n_1055),
.B1(n_1008),
.B2(n_982),
.C(n_947),
.Y(n_1110)
);

OAI22xp5_ASAP7_75t_L g1111 ( 
.A1(n_966),
.A2(n_1023),
.B1(n_1032),
.B2(n_1028),
.Y(n_1111)
);

BUFx2_ASAP7_75t_L g1112 ( 
.A(n_949),
.Y(n_1112)
);

NAND2xp5_ASAP7_75t_L g1113 ( 
.A(n_953),
.B(n_1072),
.Y(n_1113)
);

AOI221x1_ASAP7_75t_L g1114 ( 
.A1(n_972),
.A2(n_1064),
.B1(n_1025),
.B2(n_987),
.C(n_961),
.Y(n_1114)
);

AOI21x1_ASAP7_75t_L g1115 ( 
.A1(n_1018),
.A2(n_1052),
.B(n_1043),
.Y(n_1115)
);

OAI21x1_ASAP7_75t_L g1116 ( 
.A1(n_1047),
.A2(n_988),
.B(n_958),
.Y(n_1116)
);

INVxp67_ASAP7_75t_L g1117 ( 
.A(n_1004),
.Y(n_1117)
);

NAND2xp5_ASAP7_75t_SL g1118 ( 
.A(n_1020),
.B(n_1071),
.Y(n_1118)
);

INVx4_ASAP7_75t_L g1119 ( 
.A(n_998),
.Y(n_1119)
);

AOI21xp5_ASAP7_75t_L g1120 ( 
.A1(n_1041),
.A2(n_1045),
.B(n_1064),
.Y(n_1120)
);

OAI21xp33_ASAP7_75t_L g1121 ( 
.A1(n_965),
.A2(n_1070),
.B(n_956),
.Y(n_1121)
);

OAI21x1_ASAP7_75t_L g1122 ( 
.A1(n_958),
.A2(n_964),
.B(n_1049),
.Y(n_1122)
);

NAND2xp5_ASAP7_75t_L g1123 ( 
.A(n_992),
.B(n_1029),
.Y(n_1123)
);

NAND2xp5_ASAP7_75t_SL g1124 ( 
.A(n_1030),
.B(n_1035),
.Y(n_1124)
);

AND2x2_ASAP7_75t_L g1125 ( 
.A(n_1006),
.B(n_1031),
.Y(n_1125)
);

NAND2xp5_ASAP7_75t_L g1126 ( 
.A(n_964),
.B(n_1034),
.Y(n_1126)
);

A2O1A1Ixp33_ASAP7_75t_L g1127 ( 
.A1(n_1026),
.A2(n_1056),
.B(n_1051),
.C(n_1067),
.Y(n_1127)
);

AO31x2_ASAP7_75t_L g1128 ( 
.A1(n_1034),
.A2(n_1063),
.A3(n_1024),
.B(n_1042),
.Y(n_1128)
);

BUFx6f_ASAP7_75t_L g1129 ( 
.A(n_1007),
.Y(n_1129)
);

XNOR2xp5_ASAP7_75t_L g1130 ( 
.A(n_998),
.B(n_968),
.Y(n_1130)
);

BUFx6f_ASAP7_75t_L g1131 ( 
.A(n_1007),
.Y(n_1131)
);

INVx1_ASAP7_75t_L g1132 ( 
.A(n_1017),
.Y(n_1132)
);

OAI21x1_ASAP7_75t_L g1133 ( 
.A1(n_1017),
.A2(n_1037),
.B(n_1051),
.Y(n_1133)
);

OAI21xp5_ASAP7_75t_L g1134 ( 
.A1(n_1037),
.A2(n_998),
.B(n_963),
.Y(n_1134)
);

NAND2xp5_ASAP7_75t_L g1135 ( 
.A(n_1037),
.B(n_1056),
.Y(n_1135)
);

AOI21xp5_ASAP7_75t_L g1136 ( 
.A1(n_1056),
.A2(n_1054),
.B(n_990),
.Y(n_1136)
);

AO21x1_ASAP7_75t_L g1137 ( 
.A1(n_973),
.A2(n_1001),
.B(n_1048),
.Y(n_1137)
);

O2A1O1Ixp33_ASAP7_75t_SL g1138 ( 
.A1(n_1057),
.A2(n_918),
.B(n_1014),
.C(n_924),
.Y(n_1138)
);

AND2x2_ASAP7_75t_L g1139 ( 
.A(n_975),
.B(n_826),
.Y(n_1139)
);

BUFx3_ASAP7_75t_L g1140 ( 
.A(n_1002),
.Y(n_1140)
);

OAI21xp5_ASAP7_75t_L g1141 ( 
.A1(n_1048),
.A2(n_1073),
.B(n_995),
.Y(n_1141)
);

NAND2xp5_ASAP7_75t_L g1142 ( 
.A(n_1015),
.B(n_1022),
.Y(n_1142)
);

AND2x4_ASAP7_75t_L g1143 ( 
.A(n_1021),
.B(n_1005),
.Y(n_1143)
);

NAND2xp5_ASAP7_75t_L g1144 ( 
.A(n_1015),
.B(n_1022),
.Y(n_1144)
);

NOR2xp33_ASAP7_75t_L g1145 ( 
.A(n_1074),
.B(n_485),
.Y(n_1145)
);

NAND2xp5_ASAP7_75t_L g1146 ( 
.A(n_1015),
.B(n_1022),
.Y(n_1146)
);

OAI21x1_ASAP7_75t_L g1147 ( 
.A1(n_981),
.A2(n_1003),
.B(n_980),
.Y(n_1147)
);

NOR2xp67_ASAP7_75t_L g1148 ( 
.A(n_1002),
.B(n_779),
.Y(n_1148)
);

AOI21xp5_ASAP7_75t_L g1149 ( 
.A1(n_1054),
.A2(n_990),
.B(n_1001),
.Y(n_1149)
);

OR2x2_ASAP7_75t_L g1150 ( 
.A(n_957),
.B(n_828),
.Y(n_1150)
);

AOI22xp5_ASAP7_75t_L g1151 ( 
.A1(n_1074),
.A2(n_310),
.B1(n_313),
.B2(n_311),
.Y(n_1151)
);

BUFx2_ASAP7_75t_L g1152 ( 
.A(n_959),
.Y(n_1152)
);

AOI21xp33_ASAP7_75t_L g1153 ( 
.A1(n_1001),
.A2(n_1048),
.B(n_912),
.Y(n_1153)
);

NOR2xp33_ASAP7_75t_L g1154 ( 
.A(n_1074),
.B(n_485),
.Y(n_1154)
);

HB1xp67_ASAP7_75t_L g1155 ( 
.A(n_957),
.Y(n_1155)
);

OAI21xp5_ASAP7_75t_L g1156 ( 
.A1(n_1048),
.A2(n_1073),
.B(n_995),
.Y(n_1156)
);

INVx2_ASAP7_75t_L g1157 ( 
.A(n_952),
.Y(n_1157)
);

AOI21xp5_ASAP7_75t_L g1158 ( 
.A1(n_1054),
.A2(n_990),
.B(n_1001),
.Y(n_1158)
);

NOR2xp33_ASAP7_75t_R g1159 ( 
.A(n_1002),
.B(n_422),
.Y(n_1159)
);

AOI21xp5_ASAP7_75t_L g1160 ( 
.A1(n_1054),
.A2(n_990),
.B(n_1001),
.Y(n_1160)
);

O2A1O1Ixp5_ASAP7_75t_L g1161 ( 
.A1(n_1001),
.A2(n_1073),
.B(n_1027),
.C(n_912),
.Y(n_1161)
);

INVx2_ASAP7_75t_SL g1162 ( 
.A(n_1002),
.Y(n_1162)
);

NOR2xp33_ASAP7_75t_L g1163 ( 
.A(n_1074),
.B(n_485),
.Y(n_1163)
);

NAND2x1_ASAP7_75t_L g1164 ( 
.A(n_1063),
.B(n_1045),
.Y(n_1164)
);

NAND2xp5_ASAP7_75t_L g1165 ( 
.A(n_1015),
.B(n_1022),
.Y(n_1165)
);

AOI21xp5_ASAP7_75t_L g1166 ( 
.A1(n_1054),
.A2(n_990),
.B(n_1001),
.Y(n_1166)
);

NAND2xp5_ASAP7_75t_L g1167 ( 
.A(n_1015),
.B(n_1022),
.Y(n_1167)
);

NAND2xp5_ASAP7_75t_L g1168 ( 
.A(n_1015),
.B(n_1022),
.Y(n_1168)
);

INVxp67_ASAP7_75t_L g1169 ( 
.A(n_978),
.Y(n_1169)
);

INVx1_ASAP7_75t_L g1170 ( 
.A(n_952),
.Y(n_1170)
);

OAI21xp5_ASAP7_75t_L g1171 ( 
.A1(n_1048),
.A2(n_1073),
.B(n_995),
.Y(n_1171)
);

NAND2xp5_ASAP7_75t_L g1172 ( 
.A(n_1015),
.B(n_1022),
.Y(n_1172)
);

AND2x2_ASAP7_75t_L g1173 ( 
.A(n_975),
.B(n_826),
.Y(n_1173)
);

OAI21x1_ASAP7_75t_L g1174 ( 
.A1(n_981),
.A2(n_1003),
.B(n_980),
.Y(n_1174)
);

INVx1_ASAP7_75t_L g1175 ( 
.A(n_952),
.Y(n_1175)
);

AOI21xp5_ASAP7_75t_L g1176 ( 
.A1(n_1054),
.A2(n_990),
.B(n_1001),
.Y(n_1176)
);

NAND2xp5_ASAP7_75t_L g1177 ( 
.A(n_1015),
.B(n_1022),
.Y(n_1177)
);

AND2x2_ASAP7_75t_L g1178 ( 
.A(n_975),
.B(n_826),
.Y(n_1178)
);

NAND2xp5_ASAP7_75t_L g1179 ( 
.A(n_976),
.B(n_991),
.Y(n_1179)
);

AOI21xp5_ASAP7_75t_L g1180 ( 
.A1(n_1054),
.A2(n_990),
.B(n_1001),
.Y(n_1180)
);

INVx3_ASAP7_75t_L g1181 ( 
.A(n_1051),
.Y(n_1181)
);

NAND2xp5_ASAP7_75t_L g1182 ( 
.A(n_1015),
.B(n_1022),
.Y(n_1182)
);

AOI21xp5_ASAP7_75t_L g1183 ( 
.A1(n_1054),
.A2(n_990),
.B(n_1001),
.Y(n_1183)
);

OAI21x1_ASAP7_75t_L g1184 ( 
.A1(n_981),
.A2(n_1003),
.B(n_980),
.Y(n_1184)
);

BUFx2_ASAP7_75t_L g1185 ( 
.A(n_959),
.Y(n_1185)
);

OAI21x1_ASAP7_75t_L g1186 ( 
.A1(n_981),
.A2(n_1003),
.B(n_980),
.Y(n_1186)
);

CKINVDCx20_ASAP7_75t_R g1187 ( 
.A(n_1002),
.Y(n_1187)
);

NOR2xp33_ASAP7_75t_L g1188 ( 
.A(n_1074),
.B(n_485),
.Y(n_1188)
);

NAND2xp5_ASAP7_75t_L g1189 ( 
.A(n_1015),
.B(n_1022),
.Y(n_1189)
);

A2O1A1Ixp33_ASAP7_75t_L g1190 ( 
.A1(n_1048),
.A2(n_1001),
.B(n_643),
.C(n_766),
.Y(n_1190)
);

INVx3_ASAP7_75t_L g1191 ( 
.A(n_1051),
.Y(n_1191)
);

OAI21xp5_ASAP7_75t_L g1192 ( 
.A1(n_1048),
.A2(n_1073),
.B(n_995),
.Y(n_1192)
);

OAI21x1_ASAP7_75t_L g1193 ( 
.A1(n_981),
.A2(n_1003),
.B(n_980),
.Y(n_1193)
);

AO31x2_ASAP7_75t_L g1194 ( 
.A1(n_943),
.A2(n_1036),
.A3(n_1046),
.B(n_1058),
.Y(n_1194)
);

A2O1A1Ixp33_ASAP7_75t_L g1195 ( 
.A1(n_1048),
.A2(n_1001),
.B(n_643),
.C(n_766),
.Y(n_1195)
);

NAND2xp5_ASAP7_75t_L g1196 ( 
.A(n_1015),
.B(n_1022),
.Y(n_1196)
);

AOI21xp5_ASAP7_75t_L g1197 ( 
.A1(n_1054),
.A2(n_990),
.B(n_1001),
.Y(n_1197)
);

INVx1_ASAP7_75t_L g1198 ( 
.A(n_952),
.Y(n_1198)
);

OA21x2_ASAP7_75t_L g1199 ( 
.A1(n_1027),
.A2(n_948),
.B(n_994),
.Y(n_1199)
);

INVx1_ASAP7_75t_L g1200 ( 
.A(n_952),
.Y(n_1200)
);

OAI21x1_ASAP7_75t_L g1201 ( 
.A1(n_1136),
.A2(n_1147),
.B(n_1078),
.Y(n_1201)
);

INVx1_ASAP7_75t_L g1202 ( 
.A(n_1083),
.Y(n_1202)
);

CKINVDCx5p33_ASAP7_75t_R g1203 ( 
.A(n_1159),
.Y(n_1203)
);

INVx1_ASAP7_75t_L g1204 ( 
.A(n_1157),
.Y(n_1204)
);

OR2x2_ASAP7_75t_L g1205 ( 
.A(n_1080),
.B(n_1150),
.Y(n_1205)
);

NAND2xp5_ASAP7_75t_L g1206 ( 
.A(n_1179),
.B(n_1095),
.Y(n_1206)
);

OAI21xp5_ASAP7_75t_L g1207 ( 
.A1(n_1190),
.A2(n_1195),
.B(n_1075),
.Y(n_1207)
);

BUFx4f_ASAP7_75t_SL g1208 ( 
.A(n_1187),
.Y(n_1208)
);

NAND2xp5_ASAP7_75t_L g1209 ( 
.A(n_1145),
.B(n_1154),
.Y(n_1209)
);

INVx1_ASAP7_75t_L g1210 ( 
.A(n_1090),
.Y(n_1210)
);

NAND2xp5_ASAP7_75t_L g1211 ( 
.A(n_1163),
.B(n_1188),
.Y(n_1211)
);

INVxp67_ASAP7_75t_L g1212 ( 
.A(n_1155),
.Y(n_1212)
);

INVx2_ASAP7_75t_SL g1213 ( 
.A(n_1140),
.Y(n_1213)
);

NAND2x1p5_ASAP7_75t_L g1214 ( 
.A(n_1119),
.B(n_1164),
.Y(n_1214)
);

AND2x2_ASAP7_75t_L g1215 ( 
.A(n_1139),
.B(n_1173),
.Y(n_1215)
);

OAI21x1_ASAP7_75t_L g1216 ( 
.A1(n_1174),
.A2(n_1184),
.B(n_1186),
.Y(n_1216)
);

BUFx12f_ASAP7_75t_L g1217 ( 
.A(n_1094),
.Y(n_1217)
);

OAI21x1_ASAP7_75t_L g1218 ( 
.A1(n_1193),
.A2(n_1079),
.B(n_1091),
.Y(n_1218)
);

NOR2xp67_ASAP7_75t_L g1219 ( 
.A(n_1087),
.B(n_1169),
.Y(n_1219)
);

AND2x2_ASAP7_75t_L g1220 ( 
.A(n_1178),
.B(n_1109),
.Y(n_1220)
);

INVx3_ASAP7_75t_L g1221 ( 
.A(n_1133),
.Y(n_1221)
);

AO31x2_ASAP7_75t_L g1222 ( 
.A1(n_1076),
.A2(n_1176),
.A3(n_1183),
.B(n_1149),
.Y(n_1222)
);

AOI22xp33_ASAP7_75t_L g1223 ( 
.A1(n_1106),
.A2(n_1098),
.B1(n_1153),
.B2(n_1110),
.Y(n_1223)
);

INVx1_ASAP7_75t_L g1224 ( 
.A(n_1170),
.Y(n_1224)
);

NAND2xp5_ASAP7_75t_L g1225 ( 
.A(n_1101),
.B(n_1096),
.Y(n_1225)
);

NAND2xp5_ASAP7_75t_L g1226 ( 
.A(n_1096),
.B(n_1142),
.Y(n_1226)
);

NAND2x1p5_ASAP7_75t_L g1227 ( 
.A(n_1119),
.B(n_1088),
.Y(n_1227)
);

HB1xp67_ASAP7_75t_L g1228 ( 
.A(n_1088),
.Y(n_1228)
);

AOI22xp33_ASAP7_75t_L g1229 ( 
.A1(n_1153),
.A2(n_1102),
.B1(n_1137),
.B2(n_1092),
.Y(n_1229)
);

INVx1_ASAP7_75t_L g1230 ( 
.A(n_1175),
.Y(n_1230)
);

OAI21xp5_ASAP7_75t_SL g1231 ( 
.A1(n_1151),
.A2(n_1104),
.B(n_1114),
.Y(n_1231)
);

INVx1_ASAP7_75t_L g1232 ( 
.A(n_1198),
.Y(n_1232)
);

AOI22xp33_ASAP7_75t_L g1233 ( 
.A1(n_1102),
.A2(n_1086),
.B1(n_1141),
.B2(n_1171),
.Y(n_1233)
);

AOI22xp33_ASAP7_75t_L g1234 ( 
.A1(n_1141),
.A2(n_1156),
.B1(n_1192),
.B2(n_1171),
.Y(n_1234)
);

AO21x2_ASAP7_75t_L g1235 ( 
.A1(n_1158),
.A2(n_1180),
.B(n_1166),
.Y(n_1235)
);

INVx1_ASAP7_75t_L g1236 ( 
.A(n_1200),
.Y(n_1236)
);

INVx2_ASAP7_75t_SL g1237 ( 
.A(n_1162),
.Y(n_1237)
);

AO21x2_ASAP7_75t_L g1238 ( 
.A1(n_1160),
.A2(n_1197),
.B(n_1192),
.Y(n_1238)
);

OA21x2_ASAP7_75t_L g1239 ( 
.A1(n_1156),
.A2(n_1081),
.B(n_1082),
.Y(n_1239)
);

BUFx3_ASAP7_75t_L g1240 ( 
.A(n_1152),
.Y(n_1240)
);

OAI21x1_ASAP7_75t_L g1241 ( 
.A1(n_1103),
.A2(n_1099),
.B(n_1089),
.Y(n_1241)
);

OAI22xp5_ASAP7_75t_L g1242 ( 
.A1(n_1142),
.A2(n_1165),
.B1(n_1196),
.B2(n_1167),
.Y(n_1242)
);

OAI21x1_ASAP7_75t_L g1243 ( 
.A1(n_1122),
.A2(n_1116),
.B(n_1115),
.Y(n_1243)
);

NAND2xp5_ASAP7_75t_L g1244 ( 
.A(n_1144),
.B(n_1146),
.Y(n_1244)
);

OA21x2_ASAP7_75t_L g1245 ( 
.A1(n_1161),
.A2(n_1093),
.B(n_1107),
.Y(n_1245)
);

OAI21x1_ASAP7_75t_L g1246 ( 
.A1(n_1100),
.A2(n_1199),
.B(n_1108),
.Y(n_1246)
);

INVx2_ASAP7_75t_L g1247 ( 
.A(n_1144),
.Y(n_1247)
);

INVx1_ASAP7_75t_L g1248 ( 
.A(n_1113),
.Y(n_1248)
);

NAND3xp33_ASAP7_75t_L g1249 ( 
.A(n_1093),
.B(n_1111),
.C(n_1118),
.Y(n_1249)
);

OAI22xp33_ASAP7_75t_L g1250 ( 
.A1(n_1146),
.A2(n_1196),
.B1(n_1182),
.B2(n_1168),
.Y(n_1250)
);

AOI22xp33_ASAP7_75t_SL g1251 ( 
.A1(n_1134),
.A2(n_1111),
.B1(n_1105),
.B2(n_1185),
.Y(n_1251)
);

INVx1_ASAP7_75t_L g1252 ( 
.A(n_1113),
.Y(n_1252)
);

INVx2_ASAP7_75t_L g1253 ( 
.A(n_1165),
.Y(n_1253)
);

AND2x4_ASAP7_75t_L g1254 ( 
.A(n_1127),
.B(n_1181),
.Y(n_1254)
);

INVx1_ASAP7_75t_L g1255 ( 
.A(n_1123),
.Y(n_1255)
);

BUFx3_ASAP7_75t_L g1256 ( 
.A(n_1112),
.Y(n_1256)
);

INVx2_ASAP7_75t_L g1257 ( 
.A(n_1167),
.Y(n_1257)
);

OA21x2_ASAP7_75t_L g1258 ( 
.A1(n_1168),
.A2(n_1189),
.B(n_1182),
.Y(n_1258)
);

INVx3_ASAP7_75t_L g1259 ( 
.A(n_1085),
.Y(n_1259)
);

OR2x2_ASAP7_75t_L g1260 ( 
.A(n_1105),
.B(n_1117),
.Y(n_1260)
);

AND2x2_ASAP7_75t_L g1261 ( 
.A(n_1125),
.B(n_1143),
.Y(n_1261)
);

AND2x4_ASAP7_75t_L g1262 ( 
.A(n_1085),
.B(n_1191),
.Y(n_1262)
);

NAND2xp5_ASAP7_75t_L g1263 ( 
.A(n_1172),
.B(n_1177),
.Y(n_1263)
);

OAI21x1_ASAP7_75t_L g1264 ( 
.A1(n_1134),
.A2(n_1126),
.B(n_1135),
.Y(n_1264)
);

OAI21x1_ASAP7_75t_L g1265 ( 
.A1(n_1126),
.A2(n_1135),
.B(n_1123),
.Y(n_1265)
);

NAND2xp5_ASAP7_75t_SL g1266 ( 
.A(n_1121),
.B(n_1124),
.Y(n_1266)
);

OAI21x1_ASAP7_75t_L g1267 ( 
.A1(n_1181),
.A2(n_1191),
.B(n_1132),
.Y(n_1267)
);

OAI22xp5_ASAP7_75t_L g1268 ( 
.A1(n_1097),
.A2(n_1143),
.B1(n_1130),
.B2(n_1148),
.Y(n_1268)
);

INVx3_ASAP7_75t_L g1269 ( 
.A(n_1128),
.Y(n_1269)
);

OAI21xp5_ASAP7_75t_L g1270 ( 
.A1(n_1138),
.A2(n_1077),
.B(n_1194),
.Y(n_1270)
);

BUFx4f_ASAP7_75t_L g1271 ( 
.A(n_1084),
.Y(n_1271)
);

AO21x2_ASAP7_75t_L g1272 ( 
.A1(n_1077),
.A2(n_1194),
.B(n_1128),
.Y(n_1272)
);

OR2x6_ASAP7_75t_L g1273 ( 
.A(n_1129),
.B(n_1131),
.Y(n_1273)
);

AND2x2_ASAP7_75t_L g1274 ( 
.A(n_1131),
.B(n_1095),
.Y(n_1274)
);

NAND2xp5_ASAP7_75t_L g1275 ( 
.A(n_1179),
.B(n_1095),
.Y(n_1275)
);

OAI21xp5_ASAP7_75t_L g1276 ( 
.A1(n_1190),
.A2(n_1195),
.B(n_1073),
.Y(n_1276)
);

CKINVDCx5p33_ASAP7_75t_R g1277 ( 
.A(n_1159),
.Y(n_1277)
);

NAND3xp33_ASAP7_75t_L g1278 ( 
.A(n_1098),
.B(n_1106),
.C(n_722),
.Y(n_1278)
);

OR3x4_ASAP7_75t_SL g1279 ( 
.A(n_1106),
.B(n_308),
.C(n_375),
.Y(n_1279)
);

NAND2xp5_ASAP7_75t_L g1280 ( 
.A(n_1179),
.B(n_1095),
.Y(n_1280)
);

BUFx2_ASAP7_75t_L g1281 ( 
.A(n_1094),
.Y(n_1281)
);

A2O1A1Ixp33_ASAP7_75t_L g1282 ( 
.A1(n_1190),
.A2(n_1048),
.B(n_1195),
.C(n_1106),
.Y(n_1282)
);

OAI221xp5_ASAP7_75t_L g1283 ( 
.A1(n_1106),
.A2(n_1098),
.B1(n_497),
.B2(n_415),
.C(n_398),
.Y(n_1283)
);

NOR2xp33_ASAP7_75t_L g1284 ( 
.A(n_1106),
.B(n_1145),
.Y(n_1284)
);

AOI221xp5_ASAP7_75t_L g1285 ( 
.A1(n_1106),
.A2(n_487),
.B1(n_638),
.B2(n_485),
.C(n_861),
.Y(n_1285)
);

INVx2_ASAP7_75t_L g1286 ( 
.A(n_1083),
.Y(n_1286)
);

OAI21x1_ASAP7_75t_L g1287 ( 
.A1(n_1136),
.A2(n_1193),
.B(n_1147),
.Y(n_1287)
);

OAI21x1_ASAP7_75t_SL g1288 ( 
.A1(n_1137),
.A2(n_1100),
.B(n_1107),
.Y(n_1288)
);

INVx1_ASAP7_75t_L g1289 ( 
.A(n_1083),
.Y(n_1289)
);

AOI22xp33_ASAP7_75t_L g1290 ( 
.A1(n_1106),
.A2(n_934),
.B1(n_1098),
.B2(n_912),
.Y(n_1290)
);

OAI21xp5_ASAP7_75t_L g1291 ( 
.A1(n_1190),
.A2(n_1195),
.B(n_1073),
.Y(n_1291)
);

OAI21xp5_ASAP7_75t_L g1292 ( 
.A1(n_1190),
.A2(n_1195),
.B(n_1073),
.Y(n_1292)
);

INVx1_ASAP7_75t_SL g1293 ( 
.A(n_1150),
.Y(n_1293)
);

BUFx3_ASAP7_75t_L g1294 ( 
.A(n_1187),
.Y(n_1294)
);

OR2x6_ASAP7_75t_L g1295 ( 
.A(n_1134),
.B(n_1120),
.Y(n_1295)
);

OAI21x1_ASAP7_75t_L g1296 ( 
.A1(n_1136),
.A2(n_1079),
.B(n_1078),
.Y(n_1296)
);

INVx1_ASAP7_75t_L g1297 ( 
.A(n_1083),
.Y(n_1297)
);

OAI21x1_ASAP7_75t_L g1298 ( 
.A1(n_1136),
.A2(n_1079),
.B(n_1078),
.Y(n_1298)
);

OAI22xp5_ASAP7_75t_L g1299 ( 
.A1(n_1098),
.A2(n_1038),
.B1(n_1001),
.B2(n_861),
.Y(n_1299)
);

INVx2_ASAP7_75t_L g1300 ( 
.A(n_1083),
.Y(n_1300)
);

BUFx6f_ASAP7_75t_L g1301 ( 
.A(n_1084),
.Y(n_1301)
);

OAI21x1_ASAP7_75t_L g1302 ( 
.A1(n_1136),
.A2(n_1193),
.B(n_1147),
.Y(n_1302)
);

OR2x6_ASAP7_75t_L g1303 ( 
.A(n_1134),
.B(n_1120),
.Y(n_1303)
);

AOI21xp5_ASAP7_75t_L g1304 ( 
.A1(n_1076),
.A2(n_1158),
.B(n_1149),
.Y(n_1304)
);

INVx2_ASAP7_75t_L g1305 ( 
.A(n_1083),
.Y(n_1305)
);

NAND3xp33_ASAP7_75t_SL g1306 ( 
.A(n_1106),
.B(n_1098),
.C(n_938),
.Y(n_1306)
);

AO21x2_ASAP7_75t_L g1307 ( 
.A1(n_1076),
.A2(n_1158),
.B(n_1149),
.Y(n_1307)
);

OAI21x1_ASAP7_75t_L g1308 ( 
.A1(n_1136),
.A2(n_1193),
.B(n_1147),
.Y(n_1308)
);

INVx2_ASAP7_75t_L g1309 ( 
.A(n_1083),
.Y(n_1309)
);

AO21x2_ASAP7_75t_L g1310 ( 
.A1(n_1076),
.A2(n_1158),
.B(n_1149),
.Y(n_1310)
);

AOI21xp5_ASAP7_75t_SL g1311 ( 
.A1(n_1190),
.A2(n_1195),
.B(n_1075),
.Y(n_1311)
);

A2O1A1Ixp33_ASAP7_75t_L g1312 ( 
.A1(n_1190),
.A2(n_1048),
.B(n_1195),
.C(n_1106),
.Y(n_1312)
);

OAI21x1_ASAP7_75t_L g1313 ( 
.A1(n_1136),
.A2(n_1193),
.B(n_1147),
.Y(n_1313)
);

OA21x2_ASAP7_75t_L g1314 ( 
.A1(n_1149),
.A2(n_1160),
.B(n_1158),
.Y(n_1314)
);

O2A1O1Ixp33_ASAP7_75t_SL g1315 ( 
.A1(n_1190),
.A2(n_1195),
.B(n_970),
.C(n_924),
.Y(n_1315)
);

INVx2_ASAP7_75t_SL g1316 ( 
.A(n_1140),
.Y(n_1316)
);

OAI21x1_ASAP7_75t_L g1317 ( 
.A1(n_1136),
.A2(n_1193),
.B(n_1147),
.Y(n_1317)
);

AND2x6_ASAP7_75t_L g1318 ( 
.A(n_1102),
.B(n_1068),
.Y(n_1318)
);

AOI221x1_ASAP7_75t_SL g1319 ( 
.A1(n_1284),
.A2(n_1278),
.B1(n_1299),
.B2(n_1306),
.C(n_1219),
.Y(n_1319)
);

OR2x2_ASAP7_75t_L g1320 ( 
.A(n_1205),
.B(n_1293),
.Y(n_1320)
);

OAI22xp5_ASAP7_75t_L g1321 ( 
.A1(n_1223),
.A2(n_1290),
.B1(n_1284),
.B2(n_1283),
.Y(n_1321)
);

OAI211xp5_ASAP7_75t_L g1322 ( 
.A1(n_1285),
.A2(n_1223),
.B(n_1290),
.C(n_1231),
.Y(n_1322)
);

NAND2xp5_ASAP7_75t_L g1323 ( 
.A(n_1225),
.B(n_1226),
.Y(n_1323)
);

AND2x2_ASAP7_75t_L g1324 ( 
.A(n_1274),
.B(n_1220),
.Y(n_1324)
);

OAI22xp5_ASAP7_75t_L g1325 ( 
.A1(n_1251),
.A2(n_1209),
.B1(n_1211),
.B2(n_1282),
.Y(n_1325)
);

HB1xp67_ASAP7_75t_L g1326 ( 
.A(n_1272),
.Y(n_1326)
);

NAND2xp5_ASAP7_75t_L g1327 ( 
.A(n_1206),
.B(n_1275),
.Y(n_1327)
);

AND2x2_ASAP7_75t_L g1328 ( 
.A(n_1215),
.B(n_1261),
.Y(n_1328)
);

OAI22xp5_ASAP7_75t_L g1329 ( 
.A1(n_1282),
.A2(n_1312),
.B1(n_1234),
.B2(n_1229),
.Y(n_1329)
);

OR2x2_ASAP7_75t_L g1330 ( 
.A(n_1280),
.B(n_1228),
.Y(n_1330)
);

OAI22xp5_ASAP7_75t_L g1331 ( 
.A1(n_1312),
.A2(n_1234),
.B1(n_1229),
.B2(n_1244),
.Y(n_1331)
);

NOR2xp67_ASAP7_75t_L g1332 ( 
.A(n_1203),
.B(n_1277),
.Y(n_1332)
);

AOI21xp5_ASAP7_75t_L g1333 ( 
.A1(n_1304),
.A2(n_1238),
.B(n_1311),
.Y(n_1333)
);

O2A1O1Ixp33_ASAP7_75t_L g1334 ( 
.A1(n_1315),
.A2(n_1207),
.B(n_1292),
.C(n_1276),
.Y(n_1334)
);

INVxp67_ASAP7_75t_L g1335 ( 
.A(n_1260),
.Y(n_1335)
);

O2A1O1Ixp5_ASAP7_75t_SL g1336 ( 
.A1(n_1266),
.A2(n_1269),
.B(n_1291),
.C(n_1270),
.Y(n_1336)
);

NAND2xp5_ASAP7_75t_L g1337 ( 
.A(n_1263),
.B(n_1247),
.Y(n_1337)
);

A2O1A1Ixp33_ASAP7_75t_L g1338 ( 
.A1(n_1249),
.A2(n_1233),
.B(n_1242),
.C(n_1279),
.Y(n_1338)
);

NOR2xp33_ASAP7_75t_L g1339 ( 
.A(n_1266),
.B(n_1250),
.Y(n_1339)
);

AND2x4_ASAP7_75t_L g1340 ( 
.A(n_1295),
.B(n_1303),
.Y(n_1340)
);

OAI22xp5_ASAP7_75t_L g1341 ( 
.A1(n_1233),
.A2(n_1240),
.B1(n_1256),
.B2(n_1268),
.Y(n_1341)
);

AND2x2_ASAP7_75t_L g1342 ( 
.A(n_1286),
.B(n_1300),
.Y(n_1342)
);

NAND2xp5_ASAP7_75t_L g1343 ( 
.A(n_1247),
.B(n_1253),
.Y(n_1343)
);

NOR2xp67_ASAP7_75t_L g1344 ( 
.A(n_1203),
.B(n_1277),
.Y(n_1344)
);

OAI22xp5_ASAP7_75t_L g1345 ( 
.A1(n_1240),
.A2(n_1256),
.B1(n_1254),
.B2(n_1212),
.Y(n_1345)
);

O2A1O1Ixp33_ASAP7_75t_L g1346 ( 
.A1(n_1315),
.A2(n_1288),
.B(n_1295),
.C(n_1303),
.Y(n_1346)
);

OAI22xp5_ASAP7_75t_L g1347 ( 
.A1(n_1254),
.A2(n_1227),
.B1(n_1237),
.B2(n_1295),
.Y(n_1347)
);

OAI22xp5_ASAP7_75t_L g1348 ( 
.A1(n_1227),
.A2(n_1303),
.B1(n_1253),
.B2(n_1257),
.Y(n_1348)
);

OA21x2_ASAP7_75t_L g1349 ( 
.A1(n_1241),
.A2(n_1246),
.B(n_1218),
.Y(n_1349)
);

O2A1O1Ixp33_ASAP7_75t_L g1350 ( 
.A1(n_1210),
.A2(n_1232),
.B(n_1224),
.C(n_1230),
.Y(n_1350)
);

O2A1O1Ixp33_ASAP7_75t_L g1351 ( 
.A1(n_1236),
.A2(n_1297),
.B(n_1202),
.C(n_1204),
.Y(n_1351)
);

AND2x2_ASAP7_75t_L g1352 ( 
.A(n_1305),
.B(n_1309),
.Y(n_1352)
);

HB1xp67_ASAP7_75t_L g1353 ( 
.A(n_1238),
.Y(n_1353)
);

OR2x2_ASAP7_75t_L g1354 ( 
.A(n_1309),
.B(n_1289),
.Y(n_1354)
);

OA21x2_ASAP7_75t_L g1355 ( 
.A1(n_1246),
.A2(n_1218),
.B(n_1317),
.Y(n_1355)
);

INVxp67_ASAP7_75t_L g1356 ( 
.A(n_1281),
.Y(n_1356)
);

OAI22xp5_ASAP7_75t_L g1357 ( 
.A1(n_1258),
.A2(n_1316),
.B1(n_1213),
.B2(n_1255),
.Y(n_1357)
);

OA21x2_ASAP7_75t_L g1358 ( 
.A1(n_1201),
.A2(n_1308),
.B(n_1302),
.Y(n_1358)
);

OAI22xp5_ASAP7_75t_L g1359 ( 
.A1(n_1258),
.A2(n_1248),
.B1(n_1252),
.B2(n_1271),
.Y(n_1359)
);

HB1xp67_ASAP7_75t_L g1360 ( 
.A(n_1269),
.Y(n_1360)
);

INVx1_ASAP7_75t_SL g1361 ( 
.A(n_1208),
.Y(n_1361)
);

OAI22xp5_ASAP7_75t_L g1362 ( 
.A1(n_1271),
.A2(n_1214),
.B1(n_1217),
.B2(n_1262),
.Y(n_1362)
);

OAI22xp5_ASAP7_75t_L g1363 ( 
.A1(n_1214),
.A2(n_1217),
.B1(n_1259),
.B2(n_1294),
.Y(n_1363)
);

AND2x2_ASAP7_75t_L g1364 ( 
.A(n_1264),
.B(n_1265),
.Y(n_1364)
);

AOI21xp5_ASAP7_75t_L g1365 ( 
.A1(n_1307),
.A2(n_1310),
.B(n_1235),
.Y(n_1365)
);

A2O1A1Ixp33_ASAP7_75t_L g1366 ( 
.A1(n_1222),
.A2(n_1314),
.B(n_1307),
.C(n_1310),
.Y(n_1366)
);

AOI21xp5_ASAP7_75t_SL g1367 ( 
.A1(n_1314),
.A2(n_1239),
.B(n_1245),
.Y(n_1367)
);

O2A1O1Ixp33_ASAP7_75t_L g1368 ( 
.A1(n_1239),
.A2(n_1294),
.B(n_1245),
.C(n_1273),
.Y(n_1368)
);

HB1xp67_ASAP7_75t_L g1369 ( 
.A(n_1222),
.Y(n_1369)
);

INVx1_ASAP7_75t_L g1370 ( 
.A(n_1267),
.Y(n_1370)
);

AND2x4_ASAP7_75t_L g1371 ( 
.A(n_1267),
.B(n_1221),
.Y(n_1371)
);

NAND2xp5_ASAP7_75t_L g1372 ( 
.A(n_1318),
.B(n_1301),
.Y(n_1372)
);

HB1xp67_ASAP7_75t_L g1373 ( 
.A(n_1243),
.Y(n_1373)
);

HB1xp67_ASAP7_75t_L g1374 ( 
.A(n_1243),
.Y(n_1374)
);

AND2x4_ASAP7_75t_L g1375 ( 
.A(n_1296),
.B(n_1298),
.Y(n_1375)
);

OR2x6_ASAP7_75t_L g1376 ( 
.A(n_1313),
.B(n_1287),
.Y(n_1376)
);

INVx2_ASAP7_75t_L g1377 ( 
.A(n_1313),
.Y(n_1377)
);

AND2x2_ASAP7_75t_L g1378 ( 
.A(n_1216),
.B(n_1272),
.Y(n_1378)
);

AOI21xp5_ASAP7_75t_L g1379 ( 
.A1(n_1304),
.A2(n_1001),
.B(n_1238),
.Y(n_1379)
);

OAI22x1_ASAP7_75t_L g1380 ( 
.A1(n_1278),
.A2(n_1098),
.B1(n_1249),
.B2(n_1284),
.Y(n_1380)
);

O2A1O1Ixp5_ASAP7_75t_L g1381 ( 
.A1(n_1207),
.A2(n_1291),
.B(n_1292),
.C(n_1276),
.Y(n_1381)
);

AND2x4_ASAP7_75t_L g1382 ( 
.A(n_1295),
.B(n_1303),
.Y(n_1382)
);

NAND2xp5_ASAP7_75t_L g1383 ( 
.A(n_1225),
.B(n_1226),
.Y(n_1383)
);

BUFx3_ASAP7_75t_L g1384 ( 
.A(n_1281),
.Y(n_1384)
);

OAI22xp5_ASAP7_75t_L g1385 ( 
.A1(n_1223),
.A2(n_1098),
.B1(n_1290),
.B2(n_1278),
.Y(n_1385)
);

NAND2xp5_ASAP7_75t_L g1386 ( 
.A(n_1225),
.B(n_1226),
.Y(n_1386)
);

INVx3_ASAP7_75t_L g1387 ( 
.A(n_1371),
.Y(n_1387)
);

AO21x2_ASAP7_75t_L g1388 ( 
.A1(n_1365),
.A2(n_1333),
.B(n_1366),
.Y(n_1388)
);

HB1xp67_ASAP7_75t_L g1389 ( 
.A(n_1326),
.Y(n_1389)
);

AOI21xp5_ASAP7_75t_L g1390 ( 
.A1(n_1334),
.A2(n_1379),
.B(n_1381),
.Y(n_1390)
);

BUFx6f_ASAP7_75t_L g1391 ( 
.A(n_1340),
.Y(n_1391)
);

AND2x4_ASAP7_75t_L g1392 ( 
.A(n_1371),
.B(n_1340),
.Y(n_1392)
);

AOI21xp5_ASAP7_75t_L g1393 ( 
.A1(n_1329),
.A2(n_1366),
.B(n_1367),
.Y(n_1393)
);

HB1xp67_ASAP7_75t_L g1394 ( 
.A(n_1326),
.Y(n_1394)
);

BUFx3_ASAP7_75t_L g1395 ( 
.A(n_1340),
.Y(n_1395)
);

INVx2_ASAP7_75t_L g1396 ( 
.A(n_1370),
.Y(n_1396)
);

NOR2x1_ASAP7_75t_R g1397 ( 
.A(n_1384),
.B(n_1382),
.Y(n_1397)
);

AOI22xp33_ASAP7_75t_L g1398 ( 
.A1(n_1385),
.A2(n_1321),
.B1(n_1380),
.B2(n_1325),
.Y(n_1398)
);

INVx1_ASAP7_75t_SL g1399 ( 
.A(n_1330),
.Y(n_1399)
);

AND2x2_ASAP7_75t_L g1400 ( 
.A(n_1364),
.B(n_1378),
.Y(n_1400)
);

AO21x2_ASAP7_75t_L g1401 ( 
.A1(n_1338),
.A2(n_1368),
.B(n_1377),
.Y(n_1401)
);

NAND2xp5_ASAP7_75t_L g1402 ( 
.A(n_1339),
.B(n_1331),
.Y(n_1402)
);

OAI221xp5_ASAP7_75t_L g1403 ( 
.A1(n_1322),
.A2(n_1319),
.B1(n_1339),
.B2(n_1346),
.C(n_1341),
.Y(n_1403)
);

BUFx3_ASAP7_75t_L g1404 ( 
.A(n_1382),
.Y(n_1404)
);

OR2x2_ASAP7_75t_L g1405 ( 
.A(n_1353),
.B(n_1369),
.Y(n_1405)
);

HB1xp67_ASAP7_75t_L g1406 ( 
.A(n_1357),
.Y(n_1406)
);

AND2x2_ASAP7_75t_L g1407 ( 
.A(n_1378),
.B(n_1369),
.Y(n_1407)
);

INVx1_ASAP7_75t_L g1408 ( 
.A(n_1350),
.Y(n_1408)
);

INVx2_ASAP7_75t_L g1409 ( 
.A(n_1349),
.Y(n_1409)
);

OA21x2_ASAP7_75t_L g1410 ( 
.A1(n_1373),
.A2(n_1374),
.B(n_1375),
.Y(n_1410)
);

INVx1_ASAP7_75t_L g1411 ( 
.A(n_1360),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_1343),
.Y(n_1412)
);

INVx1_ASAP7_75t_L g1413 ( 
.A(n_1354),
.Y(n_1413)
);

OR2x6_ASAP7_75t_L g1414 ( 
.A(n_1376),
.B(n_1348),
.Y(n_1414)
);

INVx1_ASAP7_75t_L g1415 ( 
.A(n_1342),
.Y(n_1415)
);

AND2x4_ASAP7_75t_L g1416 ( 
.A(n_1376),
.B(n_1372),
.Y(n_1416)
);

OR2x6_ASAP7_75t_L g1417 ( 
.A(n_1376),
.B(n_1347),
.Y(n_1417)
);

BUFx2_ASAP7_75t_L g1418 ( 
.A(n_1410),
.Y(n_1418)
);

AND2x2_ASAP7_75t_L g1419 ( 
.A(n_1400),
.B(n_1355),
.Y(n_1419)
);

INVx1_ASAP7_75t_SL g1420 ( 
.A(n_1399),
.Y(n_1420)
);

INVx1_ASAP7_75t_L g1421 ( 
.A(n_1396),
.Y(n_1421)
);

AND2x4_ASAP7_75t_L g1422 ( 
.A(n_1387),
.B(n_1352),
.Y(n_1422)
);

NOR2xp33_ASAP7_75t_L g1423 ( 
.A(n_1402),
.B(n_1345),
.Y(n_1423)
);

HB1xp67_ASAP7_75t_L g1424 ( 
.A(n_1389),
.Y(n_1424)
);

NAND2xp5_ASAP7_75t_L g1425 ( 
.A(n_1412),
.B(n_1359),
.Y(n_1425)
);

INVx2_ASAP7_75t_L g1426 ( 
.A(n_1409),
.Y(n_1426)
);

HB1xp67_ASAP7_75t_L g1427 ( 
.A(n_1389),
.Y(n_1427)
);

NAND2xp5_ASAP7_75t_L g1428 ( 
.A(n_1412),
.B(n_1335),
.Y(n_1428)
);

NAND2xp5_ASAP7_75t_L g1429 ( 
.A(n_1413),
.B(n_1336),
.Y(n_1429)
);

HB1xp67_ASAP7_75t_L g1430 ( 
.A(n_1394),
.Y(n_1430)
);

AND2x2_ASAP7_75t_L g1431 ( 
.A(n_1407),
.B(n_1358),
.Y(n_1431)
);

AND2x2_ASAP7_75t_L g1432 ( 
.A(n_1407),
.B(n_1358),
.Y(n_1432)
);

AO21x2_ASAP7_75t_L g1433 ( 
.A1(n_1393),
.A2(n_1351),
.B(n_1337),
.Y(n_1433)
);

INVx2_ASAP7_75t_SL g1434 ( 
.A(n_1392),
.Y(n_1434)
);

BUFx2_ASAP7_75t_L g1435 ( 
.A(n_1410),
.Y(n_1435)
);

INVxp67_ASAP7_75t_L g1436 ( 
.A(n_1406),
.Y(n_1436)
);

OAI221xp5_ASAP7_75t_L g1437 ( 
.A1(n_1423),
.A2(n_1398),
.B1(n_1402),
.B2(n_1403),
.C(n_1393),
.Y(n_1437)
);

OAI31xp33_ASAP7_75t_L g1438 ( 
.A1(n_1423),
.A2(n_1398),
.A3(n_1403),
.B(n_1408),
.Y(n_1438)
);

OAI31xp33_ASAP7_75t_SL g1439 ( 
.A1(n_1420),
.A2(n_1363),
.A3(n_1408),
.B(n_1362),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_1421),
.Y(n_1440)
);

NAND2xp5_ASAP7_75t_L g1441 ( 
.A(n_1436),
.B(n_1420),
.Y(n_1441)
);

INVx1_ASAP7_75t_L g1442 ( 
.A(n_1421),
.Y(n_1442)
);

AND2x4_ASAP7_75t_SL g1443 ( 
.A(n_1422),
.B(n_1391),
.Y(n_1443)
);

INVx1_ASAP7_75t_L g1444 ( 
.A(n_1421),
.Y(n_1444)
);

NAND2xp5_ASAP7_75t_L g1445 ( 
.A(n_1436),
.B(n_1406),
.Y(n_1445)
);

AOI22xp33_ASAP7_75t_L g1446 ( 
.A1(n_1433),
.A2(n_1380),
.B1(n_1391),
.B2(n_1395),
.Y(n_1446)
);

OAI21xp5_ASAP7_75t_L g1447 ( 
.A1(n_1425),
.A2(n_1390),
.B(n_1323),
.Y(n_1447)
);

AND2x2_ASAP7_75t_SL g1448 ( 
.A(n_1418),
.B(n_1391),
.Y(n_1448)
);

HB1xp67_ASAP7_75t_L g1449 ( 
.A(n_1424),
.Y(n_1449)
);

OAI33xp33_ASAP7_75t_L g1450 ( 
.A1(n_1429),
.A2(n_1413),
.A3(n_1411),
.B1(n_1405),
.B2(n_1327),
.B3(n_1383),
.Y(n_1450)
);

NOR2xp33_ASAP7_75t_R g1451 ( 
.A(n_1428),
.B(n_1384),
.Y(n_1451)
);

NAND2xp5_ASAP7_75t_L g1452 ( 
.A(n_1425),
.B(n_1411),
.Y(n_1452)
);

AND2x2_ASAP7_75t_L g1453 ( 
.A(n_1434),
.B(n_1392),
.Y(n_1453)
);

AOI22xp33_ASAP7_75t_L g1454 ( 
.A1(n_1433),
.A2(n_1391),
.B1(n_1395),
.B2(n_1404),
.Y(n_1454)
);

NAND3xp33_ASAP7_75t_L g1455 ( 
.A(n_1429),
.B(n_1390),
.C(n_1386),
.Y(n_1455)
);

AOI22xp5_ASAP7_75t_L g1456 ( 
.A1(n_1433),
.A2(n_1356),
.B1(n_1328),
.B2(n_1324),
.Y(n_1456)
);

AND2x2_ASAP7_75t_L g1457 ( 
.A(n_1434),
.B(n_1392),
.Y(n_1457)
);

BUFx3_ASAP7_75t_L g1458 ( 
.A(n_1427),
.Y(n_1458)
);

NAND2xp5_ASAP7_75t_L g1459 ( 
.A(n_1433),
.B(n_1427),
.Y(n_1459)
);

OAI211xp5_ASAP7_75t_SL g1460 ( 
.A1(n_1428),
.A2(n_1320),
.B(n_1361),
.C(n_1415),
.Y(n_1460)
);

HB1xp67_ASAP7_75t_L g1461 ( 
.A(n_1430),
.Y(n_1461)
);

AND2x2_ASAP7_75t_L g1462 ( 
.A(n_1419),
.B(n_1407),
.Y(n_1462)
);

AND2x2_ASAP7_75t_L g1463 ( 
.A(n_1419),
.B(n_1416),
.Y(n_1463)
);

BUFx6f_ASAP7_75t_L g1464 ( 
.A(n_1448),
.Y(n_1464)
);

NAND3xp33_ASAP7_75t_L g1465 ( 
.A(n_1438),
.B(n_1437),
.C(n_1455),
.Y(n_1465)
);

INVx1_ASAP7_75t_L g1466 ( 
.A(n_1440),
.Y(n_1466)
);

AND2x2_ASAP7_75t_L g1467 ( 
.A(n_1448),
.B(n_1431),
.Y(n_1467)
);

NAND2xp5_ASAP7_75t_SL g1468 ( 
.A(n_1451),
.B(n_1447),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_1440),
.Y(n_1469)
);

CKINVDCx16_ASAP7_75t_R g1470 ( 
.A(n_1456),
.Y(n_1470)
);

INVx1_ASAP7_75t_L g1471 ( 
.A(n_1442),
.Y(n_1471)
);

OA21x2_ASAP7_75t_L g1472 ( 
.A1(n_1459),
.A2(n_1418),
.B(n_1435),
.Y(n_1472)
);

INVx1_ASAP7_75t_L g1473 ( 
.A(n_1444),
.Y(n_1473)
);

AOI21xp5_ASAP7_75t_SL g1474 ( 
.A1(n_1447),
.A2(n_1397),
.B(n_1401),
.Y(n_1474)
);

AND2x2_ASAP7_75t_L g1475 ( 
.A(n_1448),
.B(n_1431),
.Y(n_1475)
);

AND2x2_ASAP7_75t_L g1476 ( 
.A(n_1462),
.B(n_1431),
.Y(n_1476)
);

AND2x2_ASAP7_75t_L g1477 ( 
.A(n_1463),
.B(n_1432),
.Y(n_1477)
);

HB1xp67_ASAP7_75t_L g1478 ( 
.A(n_1449),
.Y(n_1478)
);

AOI21x1_ASAP7_75t_L g1479 ( 
.A1(n_1455),
.A2(n_1435),
.B(n_1426),
.Y(n_1479)
);

INVx1_ASAP7_75t_SL g1480 ( 
.A(n_1458),
.Y(n_1480)
);

HB1xp67_ASAP7_75t_L g1481 ( 
.A(n_1461),
.Y(n_1481)
);

INVxp67_ASAP7_75t_SL g1482 ( 
.A(n_1445),
.Y(n_1482)
);

AND2x2_ASAP7_75t_L g1483 ( 
.A(n_1464),
.B(n_1463),
.Y(n_1483)
);

NOR2xp33_ASAP7_75t_L g1484 ( 
.A(n_1465),
.B(n_1460),
.Y(n_1484)
);

OR2x2_ASAP7_75t_L g1485 ( 
.A(n_1482),
.B(n_1445),
.Y(n_1485)
);

AND2x4_ASAP7_75t_L g1486 ( 
.A(n_1464),
.B(n_1443),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_1466),
.Y(n_1487)
);

AND2x2_ASAP7_75t_SL g1488 ( 
.A(n_1470),
.B(n_1439),
.Y(n_1488)
);

AND2x2_ASAP7_75t_L g1489 ( 
.A(n_1464),
.B(n_1453),
.Y(n_1489)
);

INVx1_ASAP7_75t_L g1490 ( 
.A(n_1466),
.Y(n_1490)
);

INVx1_ASAP7_75t_L g1491 ( 
.A(n_1466),
.Y(n_1491)
);

INVx1_ASAP7_75t_L g1492 ( 
.A(n_1469),
.Y(n_1492)
);

INVx1_ASAP7_75t_L g1493 ( 
.A(n_1469),
.Y(n_1493)
);

INVx1_ASAP7_75t_L g1494 ( 
.A(n_1469),
.Y(n_1494)
);

INVx2_ASAP7_75t_SL g1495 ( 
.A(n_1464),
.Y(n_1495)
);

INVx1_ASAP7_75t_SL g1496 ( 
.A(n_1468),
.Y(n_1496)
);

INVx1_ASAP7_75t_L g1497 ( 
.A(n_1471),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_1471),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_1471),
.Y(n_1499)
);

NAND2xp5_ASAP7_75t_L g1500 ( 
.A(n_1465),
.B(n_1452),
.Y(n_1500)
);

NAND2xp5_ASAP7_75t_L g1501 ( 
.A(n_1468),
.B(n_1456),
.Y(n_1501)
);

NAND2xp5_ASAP7_75t_SL g1502 ( 
.A(n_1470),
.B(n_1439),
.Y(n_1502)
);

AND2x2_ASAP7_75t_L g1503 ( 
.A(n_1464),
.B(n_1453),
.Y(n_1503)
);

AND2x2_ASAP7_75t_L g1504 ( 
.A(n_1464),
.B(n_1457),
.Y(n_1504)
);

NAND3x1_ASAP7_75t_L g1505 ( 
.A(n_1479),
.B(n_1438),
.C(n_1441),
.Y(n_1505)
);

AND2x2_ASAP7_75t_L g1506 ( 
.A(n_1464),
.B(n_1457),
.Y(n_1506)
);

AND2x4_ASAP7_75t_L g1507 ( 
.A(n_1464),
.B(n_1443),
.Y(n_1507)
);

HB1xp67_ASAP7_75t_L g1508 ( 
.A(n_1478),
.Y(n_1508)
);

NAND2xp5_ASAP7_75t_L g1509 ( 
.A(n_1470),
.B(n_1441),
.Y(n_1509)
);

INVx1_ASAP7_75t_SL g1510 ( 
.A(n_1480),
.Y(n_1510)
);

OR2x2_ASAP7_75t_L g1511 ( 
.A(n_1478),
.B(n_1458),
.Y(n_1511)
);

INVx1_ASAP7_75t_SL g1512 ( 
.A(n_1480),
.Y(n_1512)
);

NAND3xp33_ASAP7_75t_L g1513 ( 
.A(n_1474),
.B(n_1446),
.C(n_1454),
.Y(n_1513)
);

AND2x2_ASAP7_75t_L g1514 ( 
.A(n_1464),
.B(n_1467),
.Y(n_1514)
);

OR2x2_ASAP7_75t_L g1515 ( 
.A(n_1481),
.B(n_1458),
.Y(n_1515)
);

AOI21xp33_ASAP7_75t_SL g1516 ( 
.A1(n_1488),
.A2(n_1502),
.B(n_1484),
.Y(n_1516)
);

AND2x2_ASAP7_75t_L g1517 ( 
.A(n_1514),
.B(n_1467),
.Y(n_1517)
);

AND2x2_ASAP7_75t_L g1518 ( 
.A(n_1514),
.B(n_1467),
.Y(n_1518)
);

OAI22xp5_ASAP7_75t_L g1519 ( 
.A1(n_1488),
.A2(n_1475),
.B1(n_1417),
.B2(n_1414),
.Y(n_1519)
);

NOR2xp33_ASAP7_75t_SL g1520 ( 
.A(n_1496),
.B(n_1450),
.Y(n_1520)
);

INVx2_ASAP7_75t_SL g1521 ( 
.A(n_1486),
.Y(n_1521)
);

INVx2_ASAP7_75t_L g1522 ( 
.A(n_1495),
.Y(n_1522)
);

OR2x2_ASAP7_75t_L g1523 ( 
.A(n_1508),
.B(n_1481),
.Y(n_1523)
);

NAND2xp5_ASAP7_75t_L g1524 ( 
.A(n_1500),
.B(n_1477),
.Y(n_1524)
);

AND2x2_ASAP7_75t_L g1525 ( 
.A(n_1486),
.B(n_1475),
.Y(n_1525)
);

BUFx2_ASAP7_75t_L g1526 ( 
.A(n_1505),
.Y(n_1526)
);

AND2x4_ASAP7_75t_L g1527 ( 
.A(n_1486),
.B(n_1475),
.Y(n_1527)
);

INVxp67_ASAP7_75t_SL g1528 ( 
.A(n_1505),
.Y(n_1528)
);

INVx2_ASAP7_75t_L g1529 ( 
.A(n_1495),
.Y(n_1529)
);

OR2x2_ASAP7_75t_L g1530 ( 
.A(n_1485),
.B(n_1473),
.Y(n_1530)
);

AND2x2_ASAP7_75t_L g1531 ( 
.A(n_1507),
.B(n_1477),
.Y(n_1531)
);

INVx1_ASAP7_75t_L g1532 ( 
.A(n_1499),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_1499),
.Y(n_1533)
);

NAND2xp5_ASAP7_75t_L g1534 ( 
.A(n_1510),
.B(n_1477),
.Y(n_1534)
);

BUFx2_ASAP7_75t_L g1535 ( 
.A(n_1507),
.Y(n_1535)
);

NAND2xp5_ASAP7_75t_L g1536 ( 
.A(n_1512),
.B(n_1501),
.Y(n_1536)
);

AND2x2_ASAP7_75t_SL g1537 ( 
.A(n_1502),
.B(n_1472),
.Y(n_1537)
);

NAND2xp5_ASAP7_75t_L g1538 ( 
.A(n_1509),
.B(n_1476),
.Y(n_1538)
);

INVx1_ASAP7_75t_L g1539 ( 
.A(n_1487),
.Y(n_1539)
);

AND2x2_ASAP7_75t_L g1540 ( 
.A(n_1507),
.B(n_1483),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_1490),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_1491),
.Y(n_1542)
);

INVx1_ASAP7_75t_L g1543 ( 
.A(n_1492),
.Y(n_1543)
);

NAND2xp5_ASAP7_75t_L g1544 ( 
.A(n_1485),
.B(n_1483),
.Y(n_1544)
);

INVx1_ASAP7_75t_L g1545 ( 
.A(n_1493),
.Y(n_1545)
);

INVx1_ASAP7_75t_L g1546 ( 
.A(n_1494),
.Y(n_1546)
);

INVx1_ASAP7_75t_L g1547 ( 
.A(n_1497),
.Y(n_1547)
);

AND2x2_ASAP7_75t_L g1548 ( 
.A(n_1489),
.B(n_1476),
.Y(n_1548)
);

OR2x2_ASAP7_75t_L g1549 ( 
.A(n_1511),
.B(n_1515),
.Y(n_1549)
);

INVx1_ASAP7_75t_L g1550 ( 
.A(n_1498),
.Y(n_1550)
);

AND2x4_ASAP7_75t_L g1551 ( 
.A(n_1527),
.B(n_1489),
.Y(n_1551)
);

INVx1_ASAP7_75t_L g1552 ( 
.A(n_1532),
.Y(n_1552)
);

INVx2_ASAP7_75t_SL g1553 ( 
.A(n_1527),
.Y(n_1553)
);

NAND2xp5_ASAP7_75t_L g1554 ( 
.A(n_1516),
.B(n_1503),
.Y(n_1554)
);

CKINVDCx16_ASAP7_75t_R g1555 ( 
.A(n_1526),
.Y(n_1555)
);

INVx1_ASAP7_75t_L g1556 ( 
.A(n_1532),
.Y(n_1556)
);

NAND2xp5_ASAP7_75t_L g1557 ( 
.A(n_1528),
.B(n_1503),
.Y(n_1557)
);

INVx2_ASAP7_75t_L g1558 ( 
.A(n_1537),
.Y(n_1558)
);

NAND2xp5_ASAP7_75t_L g1559 ( 
.A(n_1535),
.B(n_1504),
.Y(n_1559)
);

INVx2_ASAP7_75t_SL g1560 ( 
.A(n_1527),
.Y(n_1560)
);

AND2x2_ASAP7_75t_L g1561 ( 
.A(n_1540),
.B(n_1504),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1533),
.Y(n_1562)
);

AND2x2_ASAP7_75t_L g1563 ( 
.A(n_1540),
.B(n_1506),
.Y(n_1563)
);

AOI22xp33_ASAP7_75t_L g1564 ( 
.A1(n_1526),
.A2(n_1513),
.B1(n_1506),
.B2(n_1388),
.Y(n_1564)
);

INVx1_ASAP7_75t_L g1565 ( 
.A(n_1533),
.Y(n_1565)
);

OR2x6_ASAP7_75t_L g1566 ( 
.A(n_1521),
.B(n_1479),
.Y(n_1566)
);

INVx1_ASAP7_75t_L g1567 ( 
.A(n_1523),
.Y(n_1567)
);

INVx1_ASAP7_75t_SL g1568 ( 
.A(n_1535),
.Y(n_1568)
);

INVx2_ASAP7_75t_L g1569 ( 
.A(n_1537),
.Y(n_1569)
);

INVx2_ASAP7_75t_L g1570 ( 
.A(n_1517),
.Y(n_1570)
);

AND2x4_ASAP7_75t_L g1571 ( 
.A(n_1525),
.B(n_1521),
.Y(n_1571)
);

BUFx2_ASAP7_75t_L g1572 ( 
.A(n_1523),
.Y(n_1572)
);

HB1xp67_ASAP7_75t_L g1573 ( 
.A(n_1549),
.Y(n_1573)
);

INVx2_ASAP7_75t_L g1574 ( 
.A(n_1517),
.Y(n_1574)
);

INVx4_ASAP7_75t_L g1575 ( 
.A(n_1549),
.Y(n_1575)
);

INVx1_ASAP7_75t_L g1576 ( 
.A(n_1573),
.Y(n_1576)
);

NAND4xp25_ASAP7_75t_L g1577 ( 
.A(n_1554),
.B(n_1536),
.C(n_1520),
.D(n_1544),
.Y(n_1577)
);

AOI221xp5_ASAP7_75t_L g1578 ( 
.A1(n_1555),
.A2(n_1519),
.B1(n_1524),
.B2(n_1550),
.C(n_1539),
.Y(n_1578)
);

OAI33xp33_ASAP7_75t_L g1579 ( 
.A1(n_1557),
.A2(n_1567),
.A3(n_1559),
.B1(n_1558),
.B2(n_1569),
.B3(n_1556),
.Y(n_1579)
);

INVx2_ASAP7_75t_L g1580 ( 
.A(n_1575),
.Y(n_1580)
);

AND2x2_ASAP7_75t_L g1581 ( 
.A(n_1561),
.B(n_1525),
.Y(n_1581)
);

NAND2xp5_ASAP7_75t_L g1582 ( 
.A(n_1555),
.B(n_1541),
.Y(n_1582)
);

CKINVDCx20_ASAP7_75t_R g1583 ( 
.A(n_1561),
.Y(n_1583)
);

INVx2_ASAP7_75t_SL g1584 ( 
.A(n_1571),
.Y(n_1584)
);

INVx1_ASAP7_75t_L g1585 ( 
.A(n_1572),
.Y(n_1585)
);

INVx1_ASAP7_75t_L g1586 ( 
.A(n_1572),
.Y(n_1586)
);

AOI221xp5_ASAP7_75t_L g1587 ( 
.A1(n_1564),
.A2(n_1542),
.B1(n_1547),
.B2(n_1546),
.C(n_1543),
.Y(n_1587)
);

INVx1_ASAP7_75t_L g1588 ( 
.A(n_1575),
.Y(n_1588)
);

INVx1_ASAP7_75t_L g1589 ( 
.A(n_1575),
.Y(n_1589)
);

AOI221xp5_ASAP7_75t_L g1590 ( 
.A1(n_1568),
.A2(n_1542),
.B1(n_1547),
.B2(n_1546),
.C(n_1543),
.Y(n_1590)
);

INVx1_ASAP7_75t_L g1591 ( 
.A(n_1575),
.Y(n_1591)
);

AND2x4_ASAP7_75t_L g1592 ( 
.A(n_1553),
.B(n_1531),
.Y(n_1592)
);

INVx2_ASAP7_75t_L g1593 ( 
.A(n_1571),
.Y(n_1593)
);

INVx2_ASAP7_75t_L g1594 ( 
.A(n_1571),
.Y(n_1594)
);

BUFx2_ASAP7_75t_L g1595 ( 
.A(n_1583),
.Y(n_1595)
);

AND2x2_ASAP7_75t_L g1596 ( 
.A(n_1581),
.B(n_1571),
.Y(n_1596)
);

NAND2xp5_ASAP7_75t_L g1597 ( 
.A(n_1584),
.B(n_1568),
.Y(n_1597)
);

NOR2xp33_ASAP7_75t_L g1598 ( 
.A(n_1585),
.B(n_1586),
.Y(n_1598)
);

NAND2xp5_ASAP7_75t_L g1599 ( 
.A(n_1593),
.B(n_1553),
.Y(n_1599)
);

INVx1_ASAP7_75t_L g1600 ( 
.A(n_1576),
.Y(n_1600)
);

NAND2xp5_ASAP7_75t_SL g1601 ( 
.A(n_1578),
.B(n_1551),
.Y(n_1601)
);

AND2x2_ASAP7_75t_L g1602 ( 
.A(n_1592),
.B(n_1560),
.Y(n_1602)
);

INVx1_ASAP7_75t_L g1603 ( 
.A(n_1588),
.Y(n_1603)
);

HB1xp67_ASAP7_75t_L g1604 ( 
.A(n_1589),
.Y(n_1604)
);

NOR2x1_ASAP7_75t_L g1605 ( 
.A(n_1591),
.B(n_1567),
.Y(n_1605)
);

O2A1O1Ixp5_ASAP7_75t_SL g1606 ( 
.A1(n_1604),
.A2(n_1562),
.B(n_1556),
.C(n_1552),
.Y(n_1606)
);

CKINVDCx20_ASAP7_75t_R g1607 ( 
.A(n_1595),
.Y(n_1607)
);

OAI21xp33_ASAP7_75t_L g1608 ( 
.A1(n_1596),
.A2(n_1577),
.B(n_1560),
.Y(n_1608)
);

AOI21xp5_ASAP7_75t_L g1609 ( 
.A1(n_1601),
.A2(n_1587),
.B(n_1578),
.Y(n_1609)
);

NOR3xp33_ASAP7_75t_L g1610 ( 
.A(n_1597),
.B(n_1579),
.C(n_1582),
.Y(n_1610)
);

AOI22xp5_ASAP7_75t_L g1611 ( 
.A1(n_1602),
.A2(n_1592),
.B1(n_1551),
.B2(n_1587),
.Y(n_1611)
);

AOI222xp33_ASAP7_75t_L g1612 ( 
.A1(n_1598),
.A2(n_1590),
.B1(n_1582),
.B2(n_1558),
.C1(n_1569),
.C2(n_1580),
.Y(n_1612)
);

OAI221xp5_ASAP7_75t_L g1613 ( 
.A1(n_1598),
.A2(n_1590),
.B1(n_1558),
.B2(n_1569),
.C(n_1594),
.Y(n_1613)
);

AOI22xp5_ASAP7_75t_L g1614 ( 
.A1(n_1600),
.A2(n_1551),
.B1(n_1563),
.B2(n_1574),
.Y(n_1614)
);

AOI211xp5_ASAP7_75t_L g1615 ( 
.A1(n_1599),
.A2(n_1574),
.B(n_1570),
.C(n_1551),
.Y(n_1615)
);

OAI21xp5_ASAP7_75t_L g1616 ( 
.A1(n_1609),
.A2(n_1605),
.B(n_1603),
.Y(n_1616)
);

AOI22xp33_ASAP7_75t_L g1617 ( 
.A1(n_1610),
.A2(n_1563),
.B1(n_1574),
.B2(n_1570),
.Y(n_1617)
);

INVxp67_ASAP7_75t_L g1618 ( 
.A(n_1613),
.Y(n_1618)
);

INVx1_ASAP7_75t_L g1619 ( 
.A(n_1614),
.Y(n_1619)
);

OAI31xp33_ASAP7_75t_L g1620 ( 
.A1(n_1608),
.A2(n_1612),
.A3(n_1604),
.B(n_1570),
.Y(n_1620)
);

NAND2xp5_ASAP7_75t_L g1621 ( 
.A(n_1617),
.B(n_1611),
.Y(n_1621)
);

OR2x2_ASAP7_75t_L g1622 ( 
.A(n_1619),
.B(n_1538),
.Y(n_1622)
);

NAND2xp5_ASAP7_75t_L g1623 ( 
.A(n_1620),
.B(n_1607),
.Y(n_1623)
);

HB1xp67_ASAP7_75t_L g1624 ( 
.A(n_1616),
.Y(n_1624)
);

INVx1_ASAP7_75t_L g1625 ( 
.A(n_1619),
.Y(n_1625)
);

NOR2xp67_ASAP7_75t_L g1626 ( 
.A(n_1618),
.B(n_1552),
.Y(n_1626)
);

AND2x2_ASAP7_75t_L g1627 ( 
.A(n_1625),
.B(n_1615),
.Y(n_1627)
);

HB1xp67_ASAP7_75t_L g1628 ( 
.A(n_1626),
.Y(n_1628)
);

INVx1_ASAP7_75t_L g1629 ( 
.A(n_1622),
.Y(n_1629)
);

OAI22xp5_ASAP7_75t_L g1630 ( 
.A1(n_1624),
.A2(n_1566),
.B1(n_1565),
.B2(n_1562),
.Y(n_1630)
);

XOR2x2_ASAP7_75t_L g1631 ( 
.A(n_1623),
.B(n_1332),
.Y(n_1631)
);

AND3x2_ASAP7_75t_L g1632 ( 
.A(n_1628),
.B(n_1621),
.C(n_1606),
.Y(n_1632)
);

NAND2xp5_ASAP7_75t_L g1633 ( 
.A(n_1627),
.B(n_1518),
.Y(n_1633)
);

INVx1_ASAP7_75t_SL g1634 ( 
.A(n_1629),
.Y(n_1634)
);

NAND2xp5_ASAP7_75t_SL g1635 ( 
.A(n_1634),
.B(n_1630),
.Y(n_1635)
);

AOI221xp5_ASAP7_75t_L g1636 ( 
.A1(n_1635),
.A2(n_1633),
.B1(n_1630),
.B2(n_1632),
.C(n_1565),
.Y(n_1636)
);

INVx2_ASAP7_75t_L g1637 ( 
.A(n_1636),
.Y(n_1637)
);

AND3x2_ASAP7_75t_L g1638 ( 
.A(n_1636),
.B(n_1631),
.C(n_1529),
.Y(n_1638)
);

OAI211xp5_ASAP7_75t_SL g1639 ( 
.A1(n_1637),
.A2(n_1529),
.B(n_1522),
.C(n_1541),
.Y(n_1639)
);

NAND2xp5_ASAP7_75t_L g1640 ( 
.A(n_1638),
.B(n_1522),
.Y(n_1640)
);

INVx2_ASAP7_75t_L g1641 ( 
.A(n_1640),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_1639),
.Y(n_1642)
);

INVx1_ASAP7_75t_SL g1643 ( 
.A(n_1642),
.Y(n_1643)
);

NAND2xp5_ASAP7_75t_SL g1644 ( 
.A(n_1643),
.B(n_1641),
.Y(n_1644)
);

AOI22xp33_ASAP7_75t_SL g1645 ( 
.A1(n_1644),
.A2(n_1566),
.B1(n_1545),
.B2(n_1518),
.Y(n_1645)
);

OAI21x1_ASAP7_75t_SL g1646 ( 
.A1(n_1645),
.A2(n_1545),
.B(n_1534),
.Y(n_1646)
);

AOI22xp5_ASAP7_75t_L g1647 ( 
.A1(n_1646),
.A2(n_1566),
.B1(n_1531),
.B2(n_1344),
.Y(n_1647)
);

AOI211xp5_ASAP7_75t_L g1648 ( 
.A1(n_1647),
.A2(n_1530),
.B(n_1548),
.C(n_1515),
.Y(n_1648)
);


endmodule