module fake_jpeg_19463_n_333 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_333);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_333;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_12),
.Y(n_20)
);

BUFx12_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

INVx5_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

BUFx6f_ASAP7_75t_SL g25 ( 
.A(n_12),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_15),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_14),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

INVx11_ASAP7_75t_SL g32 ( 
.A(n_5),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

CKINVDCx12_ASAP7_75t_R g35 ( 
.A(n_1),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_11),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_7),
.Y(n_37)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_8),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_35),
.B(n_15),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_39),
.B(n_43),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_23),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g69 ( 
.A(n_40),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_23),
.Y(n_41)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_23),
.Y(n_42)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_42),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g43 ( 
.A(n_20),
.B(n_14),
.Y(n_43)
);

INVx11_ASAP7_75t_L g44 ( 
.A(n_32),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_23),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_45),
.Y(n_62)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_23),
.Y(n_46)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_46),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_L g47 ( 
.A1(n_30),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_47),
.A2(n_33),
.B1(n_37),
.B2(n_17),
.Y(n_60)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_19),
.Y(n_48)
);

INVx6_ASAP7_75t_L g92 ( 
.A(n_48),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_19),
.Y(n_49)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_49),
.Y(n_64)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

INVx11_ASAP7_75t_L g65 ( 
.A(n_50),
.Y(n_65)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_24),
.Y(n_51)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_51),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_21),
.B(n_13),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_52),
.B(n_21),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_43),
.B(n_20),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_53),
.B(n_57),
.Y(n_102)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_50),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_55),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_43),
.B(n_29),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_51),
.A2(n_30),
.B1(n_33),
.B2(n_38),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_58),
.A2(n_73),
.B1(n_91),
.B2(n_3),
.Y(n_121)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_46),
.Y(n_59)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_59),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_60),
.A2(n_63),
.B1(n_74),
.B2(n_77),
.Y(n_117)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_50),
.Y(n_61)
);

CKINVDCx16_ASAP7_75t_R g128 ( 
.A(n_61),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_48),
.A2(n_38),
.B1(n_34),
.B2(n_24),
.Y(n_63)
);

HAxp5_ASAP7_75t_SL g66 ( 
.A(n_50),
.B(n_32),
.CON(n_66),
.SN(n_66)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_66),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_67),
.B(n_71),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_52),
.B(n_28),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_68),
.B(n_80),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_39),
.B(n_28),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_50),
.B(n_36),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_72),
.B(n_75),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_51),
.A2(n_38),
.B1(n_34),
.B2(n_24),
.Y(n_73)
);

OAI22xp33_ASAP7_75t_L g74 ( 
.A1(n_48),
.A2(n_34),
.B1(n_25),
.B2(n_27),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_50),
.B(n_36),
.Y(n_75)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_46),
.Y(n_76)
);

INVx5_ASAP7_75t_L g115 ( 
.A(n_76),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_51),
.A2(n_29),
.B1(n_16),
.B2(n_37),
.Y(n_77)
);

INVx5_ASAP7_75t_L g78 ( 
.A(n_45),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_78),
.B(n_81),
.Y(n_120)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_45),
.Y(n_79)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_79),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_47),
.B(n_16),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_41),
.B(n_18),
.Y(n_81)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_40),
.Y(n_82)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_82),
.Y(n_122)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_45),
.Y(n_83)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_83),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_L g85 ( 
.A1(n_44),
.A2(n_18),
.B1(n_26),
.B2(n_17),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_L g105 ( 
.A1(n_85),
.A2(n_93),
.B1(n_27),
.B2(n_22),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_41),
.B(n_26),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_86),
.Y(n_130)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_40),
.Y(n_87)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_87),
.Y(n_131)
);

INVx11_ASAP7_75t_L g88 ( 
.A(n_40),
.Y(n_88)
);

INVx1_ASAP7_75t_SL g118 ( 
.A(n_88),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_40),
.B(n_21),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_89),
.B(n_96),
.Y(n_132)
);

INVx5_ASAP7_75t_L g91 ( 
.A(n_40),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_L g93 ( 
.A1(n_44),
.A2(n_25),
.B1(n_49),
.B2(n_21),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_42),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_94),
.B(n_97),
.Y(n_111)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_42),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_95),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_49),
.B(n_31),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_49),
.B(n_31),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_43),
.B(n_21),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_98),
.B(n_100),
.C(n_7),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_43),
.B(n_25),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_99),
.A2(n_13),
.B1(n_11),
.B2(n_10),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_43),
.B(n_22),
.Y(n_100)
);

OA22x2_ASAP7_75t_L g101 ( 
.A1(n_92),
.A2(n_27),
.B1(n_19),
.B2(n_31),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_101),
.A2(n_124),
.B1(n_64),
.B2(n_83),
.Y(n_135)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_105),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_L g106 ( 
.A1(n_97),
.A2(n_22),
.B1(n_1),
.B2(n_2),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_106),
.A2(n_108),
.B1(n_119),
.B2(n_123),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_80),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_65),
.A2(n_66),
.B1(n_70),
.B2(n_88),
.Y(n_109)
);

CKINVDCx14_ASAP7_75t_R g161 ( 
.A(n_109),
.Y(n_161)
);

AND2x2_ASAP7_75t_L g151 ( 
.A(n_113),
.B(n_56),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_65),
.A2(n_13),
.B1(n_11),
.B2(n_4),
.Y(n_116)
);

CKINVDCx16_ASAP7_75t_R g141 ( 
.A(n_116),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_96),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_119)
);

CKINVDCx16_ASAP7_75t_R g157 ( 
.A(n_121),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_60),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_123)
);

OAI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_92),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_70),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_SL g168 ( 
.A(n_125),
.B(n_9),
.C(n_69),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_129),
.B(n_9),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_130),
.B(n_72),
.Y(n_134)
);

CKINVDCx14_ASAP7_75t_R g190 ( 
.A(n_134),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_135),
.A2(n_147),
.B1(n_149),
.B2(n_101),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_132),
.B(n_112),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_136),
.B(n_137),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_132),
.B(n_99),
.Y(n_137)
);

INVx1_ASAP7_75t_SL g138 ( 
.A(n_110),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_138),
.B(n_144),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_112),
.B(n_77),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_139),
.B(n_145),
.Y(n_182)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_110),
.Y(n_140)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_140),
.Y(n_170)
);

BUFx2_ASAP7_75t_L g142 ( 
.A(n_127),
.Y(n_142)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_142),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_130),
.B(n_71),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_111),
.B(n_67),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_107),
.B(n_68),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_146),
.B(n_155),
.Y(n_180)
);

O2A1O1Ixp33_ASAP7_75t_L g147 ( 
.A1(n_114),
.A2(n_79),
.B(n_89),
.C(n_59),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_111),
.B(n_63),
.C(n_94),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_148),
.B(n_152),
.C(n_161),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_117),
.A2(n_121),
.B1(n_123),
.B2(n_105),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_108),
.B(n_56),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_150),
.B(n_152),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_151),
.A2(n_113),
.B1(n_124),
.B2(n_91),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_119),
.B(n_64),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_126),
.Y(n_153)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_153),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_102),
.B(n_76),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_154),
.B(n_165),
.Y(n_189)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_126),
.Y(n_156)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_156),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_107),
.B(n_55),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_159),
.B(n_163),
.Y(n_186)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_103),
.Y(n_160)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_160),
.Y(n_191)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_103),
.Y(n_162)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_162),
.Y(n_200)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_127),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_122),
.Y(n_164)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_164),
.Y(n_204)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_122),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_SL g166 ( 
.A(n_104),
.B(n_90),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_166),
.B(n_169),
.Y(n_193)
);

INVx3_ASAP7_75t_L g167 ( 
.A(n_115),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_SL g195 ( 
.A1(n_167),
.A2(n_168),
.B1(n_118),
.B2(n_87),
.Y(n_195)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_131),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_136),
.B(n_129),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_171),
.B(n_173),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_157),
.A2(n_143),
.B1(n_117),
.B2(n_149),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_172),
.A2(n_176),
.B1(n_184),
.B2(n_194),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_SL g173 ( 
.A(n_137),
.B(n_104),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_174),
.B(n_198),
.C(n_69),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_164),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_175),
.B(n_196),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_143),
.A2(n_101),
.B1(n_120),
.B2(n_106),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g177 ( 
.A(n_166),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g232 ( 
.A(n_177),
.Y(n_232)
);

INVxp67_ASAP7_75t_L g178 ( 
.A(n_148),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_178),
.B(n_202),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_L g217 ( 
.A1(n_181),
.A2(n_147),
.B(n_168),
.Y(n_217)
);

AOI22xp33_ASAP7_75t_L g184 ( 
.A1(n_157),
.A2(n_101),
.B1(n_120),
.B2(n_74),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_192),
.A2(n_158),
.B1(n_141),
.B2(n_135),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_139),
.A2(n_101),
.B1(n_90),
.B2(n_78),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_SL g230 ( 
.A1(n_195),
.A2(n_118),
.B(n_133),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_165),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_150),
.B(n_102),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_197),
.B(n_160),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_145),
.B(n_69),
.C(n_131),
.Y(n_198)
);

BUFx24_ASAP7_75t_SL g201 ( 
.A(n_151),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_201),
.B(n_151),
.Y(n_210)
);

INVxp67_ASAP7_75t_L g202 ( 
.A(n_155),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_169),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_203),
.B(n_196),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_158),
.A2(n_84),
.B1(n_54),
.B2(n_95),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_205),
.A2(n_138),
.B1(n_141),
.B2(n_140),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_207),
.B(n_213),
.Y(n_236)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_204),
.Y(n_209)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_209),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_210),
.B(n_215),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_190),
.B(n_167),
.Y(n_211)
);

CKINVDCx14_ASAP7_75t_R g242 ( 
.A(n_211),
.Y(n_242)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_204),
.Y(n_212)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_212),
.Y(n_248)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_179),
.Y(n_214)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_214),
.Y(n_253)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_170),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_188),
.B(n_115),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_216),
.B(n_218),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_L g235 ( 
.A1(n_217),
.A2(n_228),
.B(n_230),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_220),
.B(n_221),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_182),
.B(n_162),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_182),
.B(n_185),
.Y(n_222)
);

CKINVDCx16_ASAP7_75t_R g250 ( 
.A(n_222),
.Y(n_250)
);

AOI21xp5_ASAP7_75t_L g223 ( 
.A1(n_192),
.A2(n_156),
.B(n_153),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_SL g251 ( 
.A1(n_223),
.A2(n_230),
.B(n_203),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_185),
.B(n_115),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_SL g237 ( 
.A(n_224),
.B(n_229),
.Y(n_237)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_179),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_225),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_226),
.B(n_233),
.Y(n_256)
);

AOI21x1_ASAP7_75t_SL g228 ( 
.A1(n_170),
.A2(n_69),
.B(n_118),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_193),
.B(n_189),
.Y(n_229)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_183),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_231),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_173),
.B(n_61),
.Y(n_233)
);

AOI21xp5_ASAP7_75t_L g271 ( 
.A1(n_235),
.A2(n_240),
.B(n_251),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_206),
.B(n_199),
.C(n_174),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_238),
.B(n_249),
.C(n_256),
.Y(n_257)
);

OAI21xp5_ASAP7_75t_L g240 ( 
.A1(n_217),
.A2(n_181),
.B(n_193),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_223),
.A2(n_172),
.B1(n_199),
.B2(n_197),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_243),
.A2(n_207),
.B1(n_221),
.B2(n_224),
.Y(n_262)
);

AOI322xp5_ASAP7_75t_SL g246 ( 
.A1(n_232),
.A2(n_180),
.A3(n_188),
.B1(n_171),
.B2(n_205),
.C1(n_189),
.C2(n_198),
.Y(n_246)
);

NOR3xp33_ASAP7_75t_L g258 ( 
.A(n_246),
.B(n_240),
.C(n_235),
.Y(n_258)
);

HB1xp67_ASAP7_75t_L g247 ( 
.A(n_220),
.Y(n_247)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_247),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_206),
.B(n_187),
.C(n_183),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_233),
.B(n_186),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_252),
.B(n_255),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_226),
.B(n_176),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_257),
.B(n_259),
.C(n_264),
.Y(n_276)
);

AOI321xp33_ASAP7_75t_L g284 ( 
.A1(n_258),
.A2(n_237),
.A3(n_234),
.B1(n_242),
.B2(n_191),
.C(n_200),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_256),
.B(n_208),
.C(n_222),
.Y(n_259)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_245),
.Y(n_261)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_261),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_262),
.A2(n_244),
.B1(n_248),
.B2(n_237),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_236),
.A2(n_227),
.B1(n_218),
.B2(n_219),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_263),
.A2(n_225),
.B1(n_214),
.B2(n_163),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_238),
.B(n_208),
.C(n_227),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_250),
.B(n_229),
.Y(n_265)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_265),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_L g266 ( 
.A1(n_236),
.A2(n_219),
.B1(n_175),
.B2(n_215),
.Y(n_266)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_266),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_252),
.B(n_213),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_267),
.B(n_269),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_SL g268 ( 
.A(n_234),
.B(n_187),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_268),
.B(n_274),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_SL g269 ( 
.A(n_249),
.B(n_194),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_255),
.B(n_231),
.C(n_209),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_272),
.B(n_241),
.C(n_250),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_243),
.B(n_212),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_273),
.B(n_244),
.Y(n_288)
);

A2O1A1Ixp33_ASAP7_75t_L g274 ( 
.A1(n_251),
.A2(n_200),
.B(n_191),
.C(n_228),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_245),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_SL g277 ( 
.A(n_275),
.B(n_254),
.Y(n_277)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_277),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_278),
.B(n_289),
.C(n_270),
.Y(n_292)
);

AOI21xp5_ASAP7_75t_L g279 ( 
.A1(n_274),
.A2(n_241),
.B(n_254),
.Y(n_279)
);

OAI21xp5_ASAP7_75t_SL g304 ( 
.A1(n_279),
.A2(n_290),
.B(n_128),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_281),
.B(n_291),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_284),
.B(n_142),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_264),
.A2(n_248),
.B1(n_239),
.B2(n_253),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_287),
.A2(n_260),
.B1(n_271),
.B2(n_263),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_SL g295 ( 
.A(n_288),
.B(n_267),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_257),
.B(n_272),
.C(n_270),
.Y(n_289)
);

OAI21xp5_ASAP7_75t_SL g290 ( 
.A1(n_271),
.A2(n_239),
.B(n_253),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_292),
.B(n_297),
.C(n_303),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_276),
.B(n_259),
.C(n_269),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_294),
.B(n_295),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_296),
.B(n_301),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_276),
.B(n_273),
.C(n_262),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_282),
.B(n_142),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_SL g313 ( 
.A(n_298),
.B(n_299),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_SL g299 ( 
.A(n_283),
.B(n_9),
.Y(n_299)
);

AOI21xp5_ASAP7_75t_L g307 ( 
.A1(n_300),
.A2(n_291),
.B(n_281),
.Y(n_307)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_279),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_289),
.B(n_127),
.C(n_128),
.Y(n_303)
);

AO21x1_ASAP7_75t_L g308 ( 
.A1(n_304),
.A2(n_278),
.B(n_288),
.Y(n_308)
);

AOI21xp5_ASAP7_75t_SL g305 ( 
.A1(n_293),
.A2(n_286),
.B(n_284),
.Y(n_305)
);

OAI21xp5_ASAP7_75t_L g315 ( 
.A1(n_305),
.A2(n_314),
.B(n_303),
.Y(n_315)
);

OAI21xp5_ASAP7_75t_SL g306 ( 
.A1(n_302),
.A2(n_287),
.B(n_280),
.Y(n_306)
);

OAI21xp5_ASAP7_75t_SL g318 ( 
.A1(n_306),
.A2(n_84),
.B(n_54),
.Y(n_318)
);

XOR2xp5_ASAP7_75t_L g320 ( 
.A(n_307),
.B(n_62),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_308),
.B(n_310),
.Y(n_321)
);

INVxp67_ASAP7_75t_L g310 ( 
.A(n_296),
.Y(n_310)
);

AOI21xp5_ASAP7_75t_SL g314 ( 
.A1(n_297),
.A2(n_285),
.B(n_82),
.Y(n_314)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_315),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_313),
.B(n_294),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_L g326 ( 
.A(n_316),
.B(n_318),
.Y(n_326)
);

OAI21xp33_ASAP7_75t_L g317 ( 
.A1(n_312),
.A2(n_285),
.B(n_292),
.Y(n_317)
);

OAI21xp5_ASAP7_75t_L g323 ( 
.A1(n_317),
.A2(n_322),
.B(n_310),
.Y(n_323)
);

INVxp33_ASAP7_75t_SL g319 ( 
.A(n_309),
.Y(n_319)
);

INVxp67_ASAP7_75t_L g324 ( 
.A(n_319),
.Y(n_324)
);

INVxp67_ASAP7_75t_L g327 ( 
.A(n_320),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_SL g322 ( 
.A(n_311),
.B(n_9),
.Y(n_322)
);

XNOR2xp5_ASAP7_75t_L g328 ( 
.A(n_323),
.B(n_321),
.Y(n_328)
);

AO21x1_ASAP7_75t_L g331 ( 
.A1(n_328),
.A2(n_329),
.B(n_330),
.Y(n_331)
);

XNOR2xp5_ASAP7_75t_L g329 ( 
.A(n_326),
.B(n_308),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g330 ( 
.A(n_325),
.Y(n_330)
);

A2O1A1Ixp33_ASAP7_75t_L g332 ( 
.A1(n_331),
.A2(n_324),
.B(n_319),
.C(n_327),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_SL g333 ( 
.A(n_332),
.B(n_62),
.Y(n_333)
);


endmodule