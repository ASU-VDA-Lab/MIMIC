module fake_jpeg_2755_n_554 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_554);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_554;

wire n_529;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_417;
wire n_362;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_349;
wire n_21;
wire n_288;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx8_ASAP7_75t_L g19 ( 
.A(n_18),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_16),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_17),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_18),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_13),
.Y(n_24)
);

INVx8_ASAP7_75t_L g25 ( 
.A(n_18),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_13),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_6),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_8),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_4),
.Y(n_31)
);

INVx11_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

BUFx24_ASAP7_75t_L g34 ( 
.A(n_9),
.Y(n_34)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_0),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_14),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_3),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_1),
.Y(n_38)
);

AOI21xp5_ASAP7_75t_L g39 ( 
.A1(n_15),
.A2(n_2),
.B(n_14),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_14),
.Y(n_40)
);

BUFx3_ASAP7_75t_SL g41 ( 
.A(n_1),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_11),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_13),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_6),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_8),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_7),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_8),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_8),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_16),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_0),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_12),
.Y(n_51)
);

BUFx5_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

INVx4_ASAP7_75t_L g138 ( 
.A(n_52),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_53),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_23),
.B(n_16),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_54),
.B(n_59),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_55),
.Y(n_149)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_33),
.Y(n_56)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_56),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_57),
.Y(n_121)
);

INVx11_ASAP7_75t_L g58 ( 
.A(n_44),
.Y(n_58)
);

INVx11_ASAP7_75t_L g117 ( 
.A(n_58),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_23),
.B(n_17),
.Y(n_59)
);

NAND2xp33_ASAP7_75t_SL g60 ( 
.A(n_39),
.B(n_30),
.Y(n_60)
);

OR2x2_ASAP7_75t_L g126 ( 
.A(n_60),
.B(n_86),
.Y(n_126)
);

INVx11_ASAP7_75t_L g61 ( 
.A(n_44),
.Y(n_61)
);

INVx11_ASAP7_75t_L g167 ( 
.A(n_61),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_40),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_62),
.Y(n_125)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_30),
.Y(n_63)
);

INVx4_ASAP7_75t_SL g123 ( 
.A(n_63),
.Y(n_123)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_19),
.Y(n_64)
);

BUFx4f_ASAP7_75t_SL g131 ( 
.A(n_64),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_21),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_65),
.Y(n_148)
);

INVx11_ASAP7_75t_L g66 ( 
.A(n_44),
.Y(n_66)
);

INVx4_ASAP7_75t_L g139 ( 
.A(n_66),
.Y(n_139)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_30),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g105 ( 
.A(n_67),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_20),
.B(n_17),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_68),
.B(n_71),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_21),
.Y(n_69)
);

INVx6_ASAP7_75t_L g115 ( 
.A(n_69),
.Y(n_115)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_32),
.Y(n_70)
);

INVx2_ASAP7_75t_SL g151 ( 
.A(n_70),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_20),
.B(n_15),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_29),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_72),
.B(n_85),
.Y(n_142)
);

INVx8_ASAP7_75t_L g73 ( 
.A(n_44),
.Y(n_73)
);

INVx5_ASAP7_75t_L g113 ( 
.A(n_73),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_21),
.Y(n_74)
);

BUFx12f_ASAP7_75t_L g116 ( 
.A(n_74),
.Y(n_116)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_33),
.Y(n_75)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_75),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_42),
.Y(n_76)
);

BUFx12f_ASAP7_75t_L g158 ( 
.A(n_76),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_42),
.B(n_0),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_77),
.B(n_101),
.Y(n_136)
);

INVx11_ASAP7_75t_L g78 ( 
.A(n_44),
.Y(n_78)
);

BUFx24_ASAP7_75t_L g150 ( 
.A(n_78),
.Y(n_150)
);

BUFx5_ASAP7_75t_L g79 ( 
.A(n_41),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_79),
.Y(n_120)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_42),
.Y(n_80)
);

INVx5_ASAP7_75t_L g128 ( 
.A(n_80),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_35),
.Y(n_81)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_81),
.Y(n_122)
);

INVx3_ASAP7_75t_SL g82 ( 
.A(n_41),
.Y(n_82)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_82),
.Y(n_132)
);

INVx8_ASAP7_75t_L g83 ( 
.A(n_36),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g141 ( 
.A(n_83),
.B(n_84),
.Y(n_141)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_36),
.Y(n_84)
);

AOI21xp33_ASAP7_75t_L g85 ( 
.A1(n_39),
.A2(n_15),
.B(n_1),
.Y(n_85)
);

NAND2x1_ASAP7_75t_L g86 ( 
.A(n_36),
.B(n_0),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_35),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_87),
.Y(n_110)
);

INVx11_ASAP7_75t_L g88 ( 
.A(n_34),
.Y(n_88)
);

CKINVDCx16_ASAP7_75t_R g161 ( 
.A(n_88),
.Y(n_161)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_29),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_89),
.B(n_95),
.Y(n_144)
);

INVx13_ASAP7_75t_L g90 ( 
.A(n_41),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_90),
.Y(n_156)
);

INVx5_ASAP7_75t_L g91 ( 
.A(n_19),
.Y(n_91)
);

NAND2xp33_ASAP7_75t_SL g108 ( 
.A(n_91),
.B(n_99),
.Y(n_108)
);

BUFx12f_ASAP7_75t_L g92 ( 
.A(n_19),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g159 ( 
.A(n_92),
.B(n_94),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_35),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_93),
.Y(n_157)
);

BUFx12f_ASAP7_75t_L g94 ( 
.A(n_25),
.Y(n_94)
);

CKINVDCx16_ASAP7_75t_R g95 ( 
.A(n_41),
.Y(n_95)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_36),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g163 ( 
.A(n_96),
.B(n_100),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_36),
.B(n_1),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_97),
.B(n_98),
.Y(n_146)
);

CKINVDCx14_ASAP7_75t_R g98 ( 
.A(n_41),
.Y(n_98)
);

BUFx3_ASAP7_75t_L g99 ( 
.A(n_41),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_49),
.Y(n_100)
);

INVx6_ASAP7_75t_L g101 ( 
.A(n_49),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_49),
.B(n_2),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_102),
.B(n_2),
.Y(n_137)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_32),
.Y(n_103)
);

OR2x2_ASAP7_75t_L g154 ( 
.A(n_103),
.B(n_104),
.Y(n_154)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_49),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_L g107 ( 
.A1(n_77),
.A2(n_27),
.B1(n_50),
.B2(n_46),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_107),
.A2(n_134),
.B1(n_162),
.B2(n_4),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_102),
.B(n_51),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_109),
.B(n_112),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_86),
.B(n_51),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_60),
.B(n_48),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_114),
.B(n_127),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_63),
.A2(n_32),
.B1(n_48),
.B2(n_47),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g179 ( 
.A1(n_119),
.A2(n_135),
.B1(n_152),
.B2(n_34),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_56),
.B(n_75),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_65),
.A2(n_47),
.B1(n_25),
.B2(n_50),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_129),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_104),
.A2(n_96),
.B1(n_91),
.B2(n_67),
.Y(n_130)
);

AND2x2_ASAP7_75t_L g196 ( 
.A(n_130),
.B(n_155),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_82),
.B(n_49),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_133),
.B(n_160),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_L g134 ( 
.A1(n_69),
.A2(n_24),
.B1(n_45),
.B2(n_43),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_88),
.A2(n_25),
.B1(n_46),
.B2(n_24),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_137),
.B(n_10),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_81),
.A2(n_45),
.B1(n_43),
.B2(n_38),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_140),
.A2(n_143),
.B1(n_103),
.B2(n_57),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_87),
.A2(n_38),
.B1(n_37),
.B2(n_26),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_83),
.B(n_37),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_SL g224 ( 
.A(n_147),
.B(n_153),
.Y(n_224)
);

AOI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_58),
.A2(n_31),
.B1(n_28),
.B2(n_27),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_84),
.B(n_31),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_70),
.A2(n_28),
.B1(n_26),
.B2(n_22),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_93),
.B(n_76),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_L g162 ( 
.A1(n_74),
.A2(n_34),
.B1(n_22),
.B2(n_4),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_101),
.B(n_2),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_164),
.B(n_165),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_64),
.B(n_3),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_64),
.B(n_4),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_166),
.B(n_131),
.Y(n_220)
);

INVx4_ASAP7_75t_L g168 ( 
.A(n_113),
.Y(n_168)
);

INVx3_ASAP7_75t_L g261 ( 
.A(n_168),
.Y(n_261)
);

INVx4_ASAP7_75t_L g170 ( 
.A(n_113),
.Y(n_170)
);

INVx3_ASAP7_75t_L g262 ( 
.A(n_170),
.Y(n_262)
);

INVx4_ASAP7_75t_L g171 ( 
.A(n_117),
.Y(n_171)
);

INVx1_ASAP7_75t_SL g258 ( 
.A(n_171),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_L g245 ( 
.A1(n_172),
.A2(n_178),
.B1(n_193),
.B2(n_202),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_144),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_173),
.B(n_174),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_141),
.Y(n_174)
);

BUFx3_ASAP7_75t_L g175 ( 
.A(n_120),
.Y(n_175)
);

BUFx3_ASAP7_75t_L g231 ( 
.A(n_175),
.Y(n_231)
);

AOI22xp33_ASAP7_75t_L g178 ( 
.A1(n_114),
.A2(n_55),
.B1(n_62),
.B2(n_53),
.Y(n_178)
);

INVxp67_ASAP7_75t_L g254 ( 
.A(n_179),
.Y(n_254)
);

CKINVDCx14_ASAP7_75t_R g180 ( 
.A(n_159),
.Y(n_180)
);

CKINVDCx14_ASAP7_75t_R g230 ( 
.A(n_180),
.Y(n_230)
);

AOI22xp33_ASAP7_75t_SL g181 ( 
.A1(n_140),
.A2(n_94),
.B1(n_92),
.B2(n_61),
.Y(n_181)
);

INVxp67_ASAP7_75t_L g265 ( 
.A(n_181),
.Y(n_265)
);

INVx6_ASAP7_75t_L g182 ( 
.A(n_148),
.Y(n_182)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_182),
.Y(n_249)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_123),
.Y(n_183)
);

HB1xp67_ASAP7_75t_L g256 ( 
.A(n_183),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_109),
.B(n_99),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_184),
.B(n_188),
.Y(n_234)
);

AO22x1_ASAP7_75t_SL g185 ( 
.A1(n_126),
.A2(n_90),
.B1(n_94),
.B2(n_92),
.Y(n_185)
);

A2O1A1Ixp33_ASAP7_75t_SL g241 ( 
.A1(n_185),
.A2(n_219),
.B(n_150),
.C(n_128),
.Y(n_241)
);

INVxp67_ASAP7_75t_L g186 ( 
.A(n_159),
.Y(n_186)
);

BUFx3_ASAP7_75t_L g247 ( 
.A(n_186),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_136),
.B(n_127),
.Y(n_188)
);

INVx5_ASAP7_75t_L g189 ( 
.A(n_105),
.Y(n_189)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_189),
.Y(n_253)
);

BUFx3_ASAP7_75t_L g190 ( 
.A(n_120),
.Y(n_190)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_190),
.Y(n_267)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_106),
.Y(n_191)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_191),
.Y(n_233)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_106),
.Y(n_192)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_192),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_126),
.A2(n_100),
.B1(n_73),
.B2(n_80),
.Y(n_193)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_118),
.Y(n_194)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_194),
.Y(n_246)
);

A2O1A1Ixp33_ASAP7_75t_L g195 ( 
.A1(n_142),
.A2(n_34),
.B(n_52),
.C(n_79),
.Y(n_195)
);

AND2x2_ASAP7_75t_L g238 ( 
.A(n_195),
.B(n_198),
.Y(n_238)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_123),
.Y(n_197)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_197),
.Y(n_248)
);

OAI32xp33_ASAP7_75t_L g198 ( 
.A1(n_112),
.A2(n_78),
.A3(n_66),
.B1(n_22),
.B2(n_34),
.Y(n_198)
);

AND2x2_ASAP7_75t_L g255 ( 
.A(n_199),
.B(n_212),
.Y(n_255)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_118),
.Y(n_200)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_200),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_201),
.A2(n_148),
.B1(n_121),
.B2(n_125),
.Y(n_232)
);

AOI22xp33_ASAP7_75t_L g202 ( 
.A1(n_110),
.A2(n_5),
.B1(n_7),
.B2(n_9),
.Y(n_202)
);

AOI22xp33_ASAP7_75t_L g203 ( 
.A1(n_110),
.A2(n_5),
.B1(n_7),
.B2(n_9),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_203),
.A2(n_204),
.B1(n_209),
.B2(n_211),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_146),
.A2(n_160),
.B1(n_129),
.B2(n_155),
.Y(n_204)
);

INVx3_ASAP7_75t_L g205 ( 
.A(n_105),
.Y(n_205)
);

INVxp67_ASAP7_75t_L g278 ( 
.A(n_205),
.Y(n_278)
);

INVx4_ASAP7_75t_L g206 ( 
.A(n_117),
.Y(n_206)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_206),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_130),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_207),
.A2(n_201),
.B1(n_196),
.B2(n_195),
.Y(n_283)
);

INVx5_ASAP7_75t_L g208 ( 
.A(n_116),
.Y(n_208)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_208),
.Y(n_264)
);

AOI22xp33_ASAP7_75t_L g209 ( 
.A1(n_157),
.A2(n_12),
.B1(n_10),
.B2(n_11),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_210),
.B(n_214),
.Y(n_257)
);

AOI22xp33_ASAP7_75t_L g211 ( 
.A1(n_157),
.A2(n_12),
.B1(n_10),
.B2(n_11),
.Y(n_211)
);

AND2x2_ASAP7_75t_L g212 ( 
.A(n_133),
.B(n_12),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_123),
.Y(n_213)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_213),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_141),
.Y(n_214)
);

INVx3_ASAP7_75t_SL g215 ( 
.A(n_141),
.Y(n_215)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_215),
.Y(n_275)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_122),
.Y(n_216)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_216),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_156),
.B(n_111),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_217),
.B(n_218),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_156),
.B(n_143),
.Y(n_218)
);

AO22x1_ASAP7_75t_SL g219 ( 
.A1(n_108),
.A2(n_163),
.B1(n_159),
.B2(n_132),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_220),
.B(n_223),
.Y(n_269)
);

AND2x2_ASAP7_75t_L g221 ( 
.A(n_154),
.B(n_132),
.Y(n_221)
);

AND2x2_ASAP7_75t_L g259 ( 
.A(n_221),
.B(n_228),
.Y(n_259)
);

BUFx2_ASAP7_75t_L g222 ( 
.A(n_138),
.Y(n_222)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_222),
.Y(n_281)
);

INVxp67_ASAP7_75t_L g223 ( 
.A(n_154),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_124),
.B(n_163),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_225),
.B(n_226),
.Y(n_270)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_122),
.Y(n_226)
);

AOI22xp33_ASAP7_75t_SL g227 ( 
.A1(n_151),
.A2(n_108),
.B1(n_138),
.B2(n_163),
.Y(n_227)
);

AOI22xp33_ASAP7_75t_SL g239 ( 
.A1(n_227),
.A2(n_116),
.B1(n_158),
.B2(n_167),
.Y(n_239)
);

A2O1A1Ixp33_ASAP7_75t_L g228 ( 
.A1(n_161),
.A2(n_131),
.B(n_150),
.C(n_151),
.Y(n_228)
);

CKINVDCx16_ASAP7_75t_R g229 ( 
.A(n_131),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_229),
.B(n_158),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_232),
.A2(n_242),
.B1(n_260),
.B2(n_274),
.Y(n_291)
);

AOI32xp33_ASAP7_75t_L g236 ( 
.A1(n_176),
.A2(n_139),
.A3(n_150),
.B1(n_128),
.B2(n_151),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_236),
.B(n_277),
.Y(n_287)
);

INVxp67_ASAP7_75t_L g325 ( 
.A(n_239),
.Y(n_325)
);

AND2x2_ASAP7_75t_L g332 ( 
.A(n_241),
.B(n_222),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_176),
.A2(n_115),
.B1(n_148),
.B2(n_145),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_188),
.B(n_115),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_243),
.B(n_273),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_217),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_244),
.Y(n_295)
);

NAND2xp33_ASAP7_75t_SL g252 ( 
.A(n_221),
.B(n_139),
.Y(n_252)
);

INVx1_ASAP7_75t_SL g311 ( 
.A(n_252),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_L g260 ( 
.A1(n_218),
.A2(n_149),
.B1(n_145),
.B2(n_125),
.Y(n_260)
);

AOI21xp5_ASAP7_75t_L g266 ( 
.A1(n_223),
.A2(n_150),
.B(n_167),
.Y(n_266)
);

AOI21xp5_ASAP7_75t_L g326 ( 
.A1(n_266),
.A2(n_236),
.B(n_259),
.Y(n_326)
);

INVxp67_ASAP7_75t_SL g319 ( 
.A(n_271),
.Y(n_319)
);

AOI22xp33_ASAP7_75t_L g272 ( 
.A1(n_215),
.A2(n_149),
.B1(n_121),
.B2(n_125),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_SL g312 ( 
.A1(n_272),
.A2(n_193),
.B1(n_186),
.B2(n_182),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_177),
.B(n_121),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_L g274 ( 
.A1(n_172),
.A2(n_116),
.B1(n_158),
.B2(n_169),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_177),
.B(n_116),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_276),
.B(n_185),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_224),
.B(n_158),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_187),
.B(n_184),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_280),
.B(n_282),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_169),
.B(n_212),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_283),
.A2(n_228),
.B1(n_207),
.B2(n_219),
.Y(n_316)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_248),
.Y(n_284)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_284),
.Y(n_334)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_248),
.Y(n_285)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_285),
.Y(n_343)
);

OA21x2_ASAP7_75t_L g286 ( 
.A1(n_238),
.A2(n_196),
.B(n_185),
.Y(n_286)
);

AND2x2_ASAP7_75t_L g342 ( 
.A(n_286),
.B(n_308),
.Y(n_342)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_234),
.B(n_221),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g345 ( 
.A(n_289),
.B(n_320),
.Y(n_345)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_268),
.Y(n_290)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_290),
.Y(n_347)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_268),
.Y(n_292)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_292),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_244),
.B(n_235),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_SL g355 ( 
.A(n_294),
.B(n_299),
.Y(n_355)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_233),
.Y(n_296)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_296),
.Y(n_374)
);

AO21x2_ASAP7_75t_L g297 ( 
.A1(n_241),
.A2(n_232),
.B(n_245),
.Y(n_297)
);

INVx1_ASAP7_75t_SL g336 ( 
.A(n_297),
.Y(n_336)
);

INVx8_ASAP7_75t_L g298 ( 
.A(n_278),
.Y(n_298)
);

INVx2_ASAP7_75t_L g359 ( 
.A(n_298),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_240),
.B(n_269),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_270),
.B(n_212),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_SL g346 ( 
.A(n_300),
.B(n_307),
.Y(n_346)
);

OAI21xp5_ASAP7_75t_L g301 ( 
.A1(n_259),
.A2(n_196),
.B(n_198),
.Y(n_301)
);

OAI21xp5_ASAP7_75t_SL g353 ( 
.A1(n_301),
.A2(n_326),
.B(n_332),
.Y(n_353)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_256),
.Y(n_302)
);

INVx13_ASAP7_75t_L g363 ( 
.A(n_302),
.Y(n_363)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_249),
.Y(n_303)
);

INVx2_ASAP7_75t_L g362 ( 
.A(n_303),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_304),
.B(n_314),
.Y(n_335)
);

BUFx12_ASAP7_75t_L g305 ( 
.A(n_278),
.Y(n_305)
);

INVxp67_ASAP7_75t_L g356 ( 
.A(n_305),
.Y(n_356)
);

BUFx3_ASAP7_75t_L g306 ( 
.A(n_231),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_306),
.B(n_329),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_257),
.B(n_194),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_233),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_267),
.B(n_200),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_SL g351 ( 
.A(n_309),
.B(n_318),
.Y(n_351)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_237),
.Y(n_310)
);

AND2x2_ASAP7_75t_L g368 ( 
.A(n_310),
.B(n_312),
.Y(n_368)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_237),
.Y(n_313)
);

INVxp67_ASAP7_75t_L g357 ( 
.A(n_313),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_234),
.B(n_219),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_238),
.A2(n_283),
.B1(n_235),
.B2(n_255),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_L g341 ( 
.A1(n_315),
.A2(n_316),
.B1(n_327),
.B2(n_255),
.Y(n_341)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_246),
.Y(n_317)
);

INVxp67_ASAP7_75t_L g360 ( 
.A(n_317),
.Y(n_360)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_246),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_243),
.B(n_191),
.C(n_192),
.Y(n_320)
);

CKINVDCx16_ASAP7_75t_R g321 ( 
.A(n_266),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_SL g370 ( 
.A(n_321),
.B(n_322),
.Y(n_370)
);

CKINVDCx16_ASAP7_75t_R g322 ( 
.A(n_259),
.Y(n_322)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_249),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_323),
.B(n_251),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_267),
.B(n_190),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_SL g375 ( 
.A(n_324),
.B(n_328),
.Y(n_375)
);

OAI22xp5_ASAP7_75t_SL g327 ( 
.A1(n_238),
.A2(n_216),
.B1(n_168),
.B2(n_170),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_231),
.B(n_247),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_247),
.B(n_175),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_SL g330 ( 
.A(n_255),
.B(n_205),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g358 ( 
.A(n_330),
.B(n_331),
.Y(n_358)
);

INVx3_ASAP7_75t_L g331 ( 
.A(n_261),
.Y(n_331)
);

AND2x2_ASAP7_75t_L g333 ( 
.A(n_252),
.B(n_171),
.Y(n_333)
);

OAI21xp5_ASAP7_75t_L g339 ( 
.A1(n_333),
.A2(n_326),
.B(n_230),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_295),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_337),
.B(n_340),
.Y(n_380)
);

AND2x2_ASAP7_75t_L g379 ( 
.A(n_339),
.B(n_341),
.Y(n_379)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_295),
.Y(n_340)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_344),
.Y(n_399)
);

AOI22xp5_ASAP7_75t_L g348 ( 
.A1(n_297),
.A2(n_250),
.B1(n_254),
.B2(n_273),
.Y(n_348)
);

AOI22xp5_ASAP7_75t_L g383 ( 
.A1(n_348),
.A2(n_371),
.B1(n_332),
.B2(n_297),
.Y(n_383)
);

XNOR2xp5_ASAP7_75t_L g349 ( 
.A(n_289),
.B(n_276),
.Y(n_349)
);

MAJIxp5_ASAP7_75t_L g378 ( 
.A(n_349),
.B(n_365),
.C(n_367),
.Y(n_378)
);

CKINVDCx20_ASAP7_75t_R g350 ( 
.A(n_302),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g405 ( 
.A(n_350),
.B(n_361),
.Y(n_405)
);

AO22x1_ASAP7_75t_SL g354 ( 
.A1(n_332),
.A2(n_241),
.B1(n_242),
.B2(n_275),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_354),
.B(n_369),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_L g361 ( 
.A(n_319),
.B(n_261),
.Y(n_361)
);

CKINVDCx20_ASAP7_75t_R g364 ( 
.A(n_284),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g407 ( 
.A(n_364),
.B(n_372),
.Y(n_407)
);

XOR2xp5_ASAP7_75t_L g365 ( 
.A(n_315),
.B(n_275),
.Y(n_365)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_285),
.Y(n_366)
);

AND2x2_ASAP7_75t_L g403 ( 
.A(n_366),
.B(n_323),
.Y(n_403)
);

XOR2xp5_ASAP7_75t_L g367 ( 
.A(n_314),
.B(n_293),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_293),
.B(n_241),
.Y(n_369)
);

AOI22xp5_ASAP7_75t_L g371 ( 
.A1(n_297),
.A2(n_254),
.B1(n_241),
.B2(n_265),
.Y(n_371)
);

CKINVDCx20_ASAP7_75t_R g372 ( 
.A(n_290),
.Y(n_372)
);

XOR2xp5_ASAP7_75t_L g373 ( 
.A(n_288),
.B(n_251),
.Y(n_373)
);

MAJIxp5_ASAP7_75t_L g394 ( 
.A(n_373),
.B(n_292),
.C(n_317),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_320),
.B(n_279),
.Y(n_376)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_376),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_304),
.B(n_279),
.Y(n_377)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_377),
.Y(n_413)
);

XOR2xp5_ASAP7_75t_L g381 ( 
.A(n_345),
.B(n_287),
.Y(n_381)
);

MAJIxp5_ASAP7_75t_L g434 ( 
.A(n_381),
.B(n_389),
.C(n_395),
.Y(n_434)
);

INVxp67_ASAP7_75t_L g382 ( 
.A(n_338),
.Y(n_382)
);

INVx2_ASAP7_75t_L g422 ( 
.A(n_382),
.Y(n_422)
);

AOI22xp5_ASAP7_75t_L g421 ( 
.A1(n_383),
.A2(n_391),
.B1(n_398),
.B2(n_411),
.Y(n_421)
);

AOI322xp5_ASAP7_75t_L g384 ( 
.A1(n_335),
.A2(n_301),
.A3(n_297),
.B1(n_311),
.B2(n_316),
.C1(n_286),
.C2(n_330),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_SL g417 ( 
.A(n_384),
.B(n_393),
.Y(n_417)
);

XNOR2xp5_ASAP7_75t_L g385 ( 
.A(n_345),
.B(n_286),
.Y(n_385)
);

XOR2xp5_ASAP7_75t_L g423 ( 
.A(n_385),
.B(n_387),
.Y(n_423)
);

AOI22xp5_ASAP7_75t_SL g386 ( 
.A1(n_370),
.A2(n_336),
.B1(n_325),
.B2(n_342),
.Y(n_386)
);

OAI21xp5_ASAP7_75t_SL g418 ( 
.A1(n_386),
.A2(n_390),
.B(n_392),
.Y(n_418)
);

XNOR2xp5_ASAP7_75t_L g387 ( 
.A(n_349),
.B(n_311),
.Y(n_387)
);

INVxp67_ASAP7_75t_L g388 ( 
.A(n_358),
.Y(n_388)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_388),
.Y(n_419)
);

XOR2xp5_ASAP7_75t_L g389 ( 
.A(n_373),
.B(n_333),
.Y(n_389)
);

AOI21xp5_ASAP7_75t_L g390 ( 
.A1(n_353),
.A2(n_325),
.B(n_265),
.Y(n_390)
);

AOI22xp5_ASAP7_75t_L g391 ( 
.A1(n_336),
.A2(n_291),
.B1(n_327),
.B2(n_312),
.Y(n_391)
);

OAI21xp5_ASAP7_75t_SL g392 ( 
.A1(n_353),
.A2(n_333),
.B(n_291),
.Y(n_392)
);

CKINVDCx20_ASAP7_75t_R g393 ( 
.A(n_357),
.Y(n_393)
);

XOR2xp5_ASAP7_75t_L g425 ( 
.A(n_394),
.B(n_397),
.Y(n_425)
);

MAJIxp5_ASAP7_75t_L g395 ( 
.A(n_365),
.B(n_313),
.C(n_310),
.Y(n_395)
);

OAI21xp5_ASAP7_75t_SL g396 ( 
.A1(n_339),
.A2(n_331),
.B(n_296),
.Y(n_396)
);

CKINVDCx14_ASAP7_75t_R g437 ( 
.A(n_396),
.Y(n_437)
);

XNOR2xp5_ASAP7_75t_L g397 ( 
.A(n_367),
.B(n_318),
.Y(n_397)
);

AOI22xp5_ASAP7_75t_L g398 ( 
.A1(n_348),
.A2(n_341),
.B1(n_371),
.B2(n_368),
.Y(n_398)
);

AOI22xp5_ASAP7_75t_SL g400 ( 
.A1(n_342),
.A2(n_308),
.B1(n_306),
.B2(n_253),
.Y(n_400)
);

INVxp67_ASAP7_75t_L g430 ( 
.A(n_400),
.Y(n_430)
);

CKINVDCx16_ASAP7_75t_R g401 ( 
.A(n_375),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_SL g442 ( 
.A(n_401),
.B(n_406),
.Y(n_442)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_403),
.Y(n_420)
);

OAI21xp5_ASAP7_75t_L g404 ( 
.A1(n_342),
.A2(n_298),
.B(n_253),
.Y(n_404)
);

INVxp67_ASAP7_75t_L g436 ( 
.A(n_404),
.Y(n_436)
);

OAI21xp5_ASAP7_75t_SL g406 ( 
.A1(n_340),
.A2(n_262),
.B(n_189),
.Y(n_406)
);

NOR2xp33_ASAP7_75t_L g409 ( 
.A(n_355),
.B(n_262),
.Y(n_409)
);

OAI221xp5_ASAP7_75t_L g416 ( 
.A1(n_409),
.A2(n_356),
.B1(n_351),
.B2(n_359),
.C(n_366),
.Y(n_416)
);

XOR2x2_ASAP7_75t_SL g410 ( 
.A(n_335),
.B(n_305),
.Y(n_410)
);

XNOR2xp5_ASAP7_75t_L g426 ( 
.A(n_410),
.B(n_414),
.Y(n_426)
);

AOI22xp5_ASAP7_75t_L g411 ( 
.A1(n_368),
.A2(n_303),
.B1(n_263),
.B2(n_258),
.Y(n_411)
);

OAI21xp5_ASAP7_75t_SL g412 ( 
.A1(n_369),
.A2(n_264),
.B(n_258),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_L g424 ( 
.A(n_412),
.B(n_360),
.Y(n_424)
);

MAJIxp5_ASAP7_75t_L g414 ( 
.A(n_376),
.B(n_264),
.C(n_263),
.Y(n_414)
);

XNOR2xp5_ASAP7_75t_SL g415 ( 
.A(n_381),
.B(n_346),
.Y(n_415)
);

XOR2xp5_ASAP7_75t_L g450 ( 
.A(n_415),
.B(n_429),
.Y(n_450)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_416),
.Y(n_448)
);

AOI22xp33_ASAP7_75t_SL g457 ( 
.A1(n_424),
.A2(n_379),
.B1(n_347),
.B2(n_334),
.Y(n_457)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_380),
.Y(n_427)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_427),
.Y(n_461)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_407),
.Y(n_428)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_428),
.Y(n_462)
);

XNOR2xp5_ASAP7_75t_L g429 ( 
.A(n_378),
.B(n_377),
.Y(n_429)
);

XNOR2xp5_ASAP7_75t_SL g431 ( 
.A(n_385),
.B(n_368),
.Y(n_431)
);

XOR2xp5_ASAP7_75t_L g454 ( 
.A(n_431),
.B(n_445),
.Y(n_454)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_403),
.Y(n_432)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_432),
.Y(n_473)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_405),
.Y(n_433)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_433),
.Y(n_463)
);

AOI22xp5_ASAP7_75t_L g435 ( 
.A1(n_383),
.A2(n_354),
.B1(n_360),
.B2(n_357),
.Y(n_435)
);

OAI22xp5_ASAP7_75t_SL g472 ( 
.A1(n_435),
.A2(n_444),
.B1(n_343),
.B2(n_334),
.Y(n_472)
);

CKINVDCx20_ASAP7_75t_R g438 ( 
.A(n_403),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_SL g456 ( 
.A(n_438),
.B(n_439),
.Y(n_456)
);

CKINVDCx20_ASAP7_75t_R g439 ( 
.A(n_388),
.Y(n_439)
);

CKINVDCx16_ASAP7_75t_R g440 ( 
.A(n_404),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_L g471 ( 
.A(n_440),
.B(n_443),
.Y(n_471)
);

NOR2xp33_ASAP7_75t_L g441 ( 
.A(n_382),
.B(n_356),
.Y(n_441)
);

NOR2xp33_ASAP7_75t_SL g460 ( 
.A(n_441),
.B(n_379),
.Y(n_460)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_399),
.Y(n_443)
);

AOI22xp5_ASAP7_75t_L g444 ( 
.A1(n_398),
.A2(n_354),
.B1(n_347),
.B2(n_352),
.Y(n_444)
);

XNOR2xp5_ASAP7_75t_L g445 ( 
.A(n_378),
.B(n_352),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_413),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_446),
.B(n_343),
.Y(n_449)
);

OA21x2_ASAP7_75t_SL g447 ( 
.A1(n_428),
.A2(n_402),
.B(n_390),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_447),
.B(n_455),
.Y(n_487)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_449),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_432),
.B(n_414),
.Y(n_451)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_451),
.Y(n_479)
);

MAJIxp5_ASAP7_75t_L g452 ( 
.A(n_445),
.B(n_395),
.C(n_394),
.Y(n_452)
);

MAJIxp5_ASAP7_75t_L g493 ( 
.A(n_452),
.B(n_459),
.C(n_465),
.Y(n_493)
);

XNOR2xp5_ASAP7_75t_L g453 ( 
.A(n_425),
.B(n_389),
.Y(n_453)
);

XNOR2xp5_ASAP7_75t_L g477 ( 
.A(n_453),
.B(n_464),
.Y(n_477)
);

CKINVDCx20_ASAP7_75t_R g455 ( 
.A(n_442),
.Y(n_455)
);

INVxp67_ASAP7_75t_L g476 ( 
.A(n_457),
.Y(n_476)
);

AOI21xp5_ASAP7_75t_L g458 ( 
.A1(n_437),
.A2(n_379),
.B(n_396),
.Y(n_458)
);

HB1xp67_ASAP7_75t_L g494 ( 
.A(n_458),
.Y(n_494)
);

MAJIxp5_ASAP7_75t_L g459 ( 
.A(n_434),
.B(n_397),
.C(n_387),
.Y(n_459)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_460),
.Y(n_483)
);

XNOR2xp5_ASAP7_75t_L g464 ( 
.A(n_425),
.B(n_410),
.Y(n_464)
);

MAJIxp5_ASAP7_75t_L g465 ( 
.A(n_434),
.B(n_392),
.C(n_412),
.Y(n_465)
);

MAJIxp5_ASAP7_75t_L g466 ( 
.A(n_429),
.B(n_423),
.C(n_426),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_SL g478 ( 
.A(n_466),
.B(n_468),
.Y(n_478)
);

AOI22xp5_ASAP7_75t_L g467 ( 
.A1(n_421),
.A2(n_408),
.B1(n_391),
.B2(n_386),
.Y(n_467)
);

OAI22xp5_ASAP7_75t_SL g482 ( 
.A1(n_467),
.A2(n_421),
.B1(n_435),
.B2(n_444),
.Y(n_482)
);

MAJIxp5_ASAP7_75t_L g468 ( 
.A(n_423),
.B(n_408),
.C(n_400),
.Y(n_468)
);

XOR2xp5_ASAP7_75t_L g469 ( 
.A(n_426),
.B(n_411),
.Y(n_469)
);

XOR2xp5_ASAP7_75t_L g486 ( 
.A(n_469),
.B(n_418),
.Y(n_486)
);

XNOR2xp5_ASAP7_75t_L g470 ( 
.A(n_415),
.B(n_406),
.Y(n_470)
);

XNOR2xp5_ASAP7_75t_L g485 ( 
.A(n_470),
.B(n_431),
.Y(n_485)
);

AOI22xp5_ASAP7_75t_L g484 ( 
.A1(n_472),
.A2(n_420),
.B1(n_446),
.B2(n_436),
.Y(n_484)
);

NAND4xp25_ASAP7_75t_L g474 ( 
.A(n_448),
.B(n_417),
.C(n_430),
.D(n_436),
.Y(n_474)
);

NOR2xp33_ASAP7_75t_L g497 ( 
.A(n_474),
.B(n_485),
.Y(n_497)
);

CKINVDCx16_ASAP7_75t_R g480 ( 
.A(n_471),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_SL g504 ( 
.A(n_480),
.B(n_463),
.Y(n_504)
);

XNOR2xp5_ASAP7_75t_SL g481 ( 
.A(n_464),
.B(n_454),
.Y(n_481)
);

INVxp67_ASAP7_75t_L g499 ( 
.A(n_481),
.Y(n_499)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_482),
.Y(n_507)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_484),
.Y(n_512)
);

MAJIxp5_ASAP7_75t_L g511 ( 
.A(n_486),
.B(n_496),
.C(n_450),
.Y(n_511)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_462),
.Y(n_488)
);

NOR2xp33_ASAP7_75t_L g505 ( 
.A(n_488),
.B(n_495),
.Y(n_505)
);

OAI22xp5_ASAP7_75t_SL g489 ( 
.A1(n_467),
.A2(n_473),
.B1(n_458),
.B2(n_430),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_489),
.B(n_456),
.Y(n_500)
);

XNOR2xp5_ASAP7_75t_SL g490 ( 
.A(n_454),
.B(n_418),
.Y(n_490)
);

NAND3xp33_ASAP7_75t_L g513 ( 
.A(n_490),
.B(n_491),
.C(n_344),
.Y(n_513)
);

NOR2xp33_ASAP7_75t_L g491 ( 
.A(n_463),
.B(n_419),
.Y(n_491)
);

AOI22xp33_ASAP7_75t_SL g492 ( 
.A1(n_472),
.A2(n_422),
.B1(n_359),
.B2(n_374),
.Y(n_492)
);

OAI22xp5_ASAP7_75t_L g498 ( 
.A1(n_492),
.A2(n_451),
.B1(n_468),
.B2(n_374),
.Y(n_498)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_449),
.Y(n_495)
);

XOR2xp5_ASAP7_75t_L g496 ( 
.A(n_453),
.B(n_422),
.Y(n_496)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_498),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_500),
.Y(n_527)
);

AOI21xp5_ASAP7_75t_L g501 ( 
.A1(n_494),
.A2(n_470),
.B(n_465),
.Y(n_501)
);

AOI21xp33_ASAP7_75t_L g524 ( 
.A1(n_501),
.A2(n_363),
.B(n_362),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_479),
.B(n_483),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_502),
.B(n_503),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_475),
.B(n_461),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_504),
.B(n_506),
.Y(n_517)
);

NOR2xp33_ASAP7_75t_L g506 ( 
.A(n_487),
.B(n_452),
.Y(n_506)
);

CKINVDCx20_ASAP7_75t_R g508 ( 
.A(n_484),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_508),
.B(n_510),
.Y(n_525)
);

OAI22xp5_ASAP7_75t_SL g509 ( 
.A1(n_476),
.A2(n_469),
.B1(n_450),
.B2(n_466),
.Y(n_509)
);

AOI22xp5_ASAP7_75t_SL g528 ( 
.A1(n_509),
.A2(n_499),
.B1(n_497),
.B2(n_512),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_SL g510 ( 
.A(n_493),
.B(n_459),
.Y(n_510)
);

XOR2xp5_ASAP7_75t_L g523 ( 
.A(n_511),
.B(n_363),
.Y(n_523)
);

NOR2xp33_ASAP7_75t_L g516 ( 
.A(n_513),
.B(n_490),
.Y(n_516)
);

NOR2xp33_ASAP7_75t_L g514 ( 
.A(n_476),
.B(n_362),
.Y(n_514)
);

NOR2xp33_ASAP7_75t_SL g515 ( 
.A(n_514),
.B(n_489),
.Y(n_515)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_515),
.Y(n_535)
);

AOI31xp33_ASAP7_75t_L g538 ( 
.A1(n_516),
.A2(n_503),
.A3(n_509),
.B(n_499),
.Y(n_538)
);

OAI22xp5_ASAP7_75t_SL g518 ( 
.A1(n_507),
.A2(n_482),
.B1(n_478),
.B2(n_486),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_518),
.B(n_519),
.Y(n_532)
);

MAJIxp5_ASAP7_75t_L g519 ( 
.A(n_511),
.B(n_493),
.C(n_496),
.Y(n_519)
);

OAI22xp5_ASAP7_75t_SL g521 ( 
.A1(n_507),
.A2(n_485),
.B1(n_481),
.B2(n_477),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_L g536 ( 
.A(n_521),
.B(n_522),
.Y(n_536)
);

XNOR2xp5_ASAP7_75t_L g522 ( 
.A(n_500),
.B(n_477),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_523),
.B(n_524),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_528),
.B(n_501),
.Y(n_529)
);

MAJx2_ASAP7_75t_L g543 ( 
.A(n_529),
.B(n_518),
.C(n_523),
.Y(n_543)
);

NOR2xp33_ASAP7_75t_L g530 ( 
.A(n_522),
.B(n_502),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_L g541 ( 
.A(n_530),
.B(n_531),
.Y(n_541)
);

MAJIxp5_ASAP7_75t_L g531 ( 
.A(n_519),
.B(n_512),
.C(n_508),
.Y(n_531)
);

CKINVDCx20_ASAP7_75t_R g533 ( 
.A(n_520),
.Y(n_533)
);

NOR2xp33_ASAP7_75t_L g539 ( 
.A(n_533),
.B(n_527),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_L g534 ( 
.A(n_520),
.B(n_505),
.Y(n_534)
);

AOI21xp33_ASAP7_75t_L g544 ( 
.A1(n_534),
.A2(n_521),
.B(n_305),
.Y(n_544)
);

OAI21xp5_ASAP7_75t_L g540 ( 
.A1(n_538),
.A2(n_525),
.B(n_528),
.Y(n_540)
);

NOR2xp33_ASAP7_75t_SL g545 ( 
.A(n_539),
.B(n_542),
.Y(n_545)
);

AOI21xp5_ASAP7_75t_L g548 ( 
.A1(n_540),
.A2(n_544),
.B(n_534),
.Y(n_548)
);

MAJIxp5_ASAP7_75t_L g542 ( 
.A(n_532),
.B(n_517),
.C(n_526),
.Y(n_542)
);

OAI21xp5_ASAP7_75t_L g546 ( 
.A1(n_543),
.A2(n_537),
.B(n_529),
.Y(n_546)
);

HB1xp67_ASAP7_75t_L g550 ( 
.A(n_546),
.Y(n_550)
);

NOR2xp33_ASAP7_75t_SL g547 ( 
.A(n_541),
.B(n_535),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_L g549 ( 
.A(n_547),
.B(n_548),
.Y(n_549)
);

OAI321xp33_ASAP7_75t_L g551 ( 
.A1(n_549),
.A2(n_545),
.A3(n_536),
.B1(n_531),
.B2(n_543),
.C(n_281),
.Y(n_551)
);

AOI21xp5_ASAP7_75t_L g553 ( 
.A1(n_551),
.A2(n_552),
.B(n_206),
.Y(n_553)
);

AOI21xp5_ASAP7_75t_L g552 ( 
.A1(n_550),
.A2(n_305),
.B(n_281),
.Y(n_552)
);

XNOR2xp5_ASAP7_75t_L g554 ( 
.A(n_553),
.B(n_208),
.Y(n_554)
);


endmodule