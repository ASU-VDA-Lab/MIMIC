module fake_netlist_1_6618_n_33 (n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_8, n_0, n_33);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_8;
input n_0;
output n_33;
wire n_20;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_30;
wire n_18;
wire n_32;
wire n_12;
wire n_17;
wire n_14;
wire n_10;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_27;
INVx1_ASAP7_75t_L g10 ( .A(n_8), .Y(n_10) );
INVx1_ASAP7_75t_L g11 ( .A(n_8), .Y(n_11) );
INVx3_ASAP7_75t_L g12 ( .A(n_9), .Y(n_12) );
INVx1_ASAP7_75t_L g13 ( .A(n_5), .Y(n_13) );
CKINVDCx20_ASAP7_75t_R g14 ( .A(n_5), .Y(n_14) );
CKINVDCx5p33_ASAP7_75t_R g15 ( .A(n_4), .Y(n_15) );
NAND2xp5_ASAP7_75t_L g16 ( .A(n_12), .B(n_0), .Y(n_16) );
OAI22xp5_ASAP7_75t_L g17 ( .A1(n_10), .A2(n_0), .B1(n_1), .B2(n_2), .Y(n_17) );
INVx2_ASAP7_75t_SL g18 ( .A(n_12), .Y(n_18) );
INVx2_ASAP7_75t_SL g19 ( .A(n_12), .Y(n_19) );
INVx2_ASAP7_75t_SL g20 ( .A(n_18), .Y(n_20) );
NAND2xp5_ASAP7_75t_L g21 ( .A(n_18), .B(n_12), .Y(n_21) );
INVxp67_ASAP7_75t_L g22 ( .A(n_21), .Y(n_22) );
NOR2xp33_ASAP7_75t_L g23 ( .A(n_20), .B(n_16), .Y(n_23) );
AND2x2_ASAP7_75t_L g24 ( .A(n_21), .B(n_19), .Y(n_24) );
AOI22xp33_ASAP7_75t_SL g25 ( .A1(n_22), .A2(n_14), .B1(n_17), .B2(n_15), .Y(n_25) );
NAND2xp5_ASAP7_75t_L g26 ( .A(n_22), .B(n_20), .Y(n_26) );
OAI211xp5_ASAP7_75t_L g27 ( .A1(n_25), .A2(n_23), .B(n_14), .C(n_11), .Y(n_27) );
AOI221xp5_ASAP7_75t_L g28 ( .A1(n_26), .A2(n_24), .B1(n_10), .B2(n_11), .C(n_13), .Y(n_28) );
INVx1_ASAP7_75t_L g29 ( .A(n_28), .Y(n_29) );
CKINVDCx5p33_ASAP7_75t_R g30 ( .A(n_27), .Y(n_30) );
BUFx2_ASAP7_75t_L g31 ( .A(n_28), .Y(n_31) );
XNOR2xp5_ASAP7_75t_L g32 ( .A(n_31), .B(n_1), .Y(n_32) );
AOI322xp5_ASAP7_75t_L g33 ( .A1(n_32), .A2(n_3), .A3(n_6), .B1(n_7), .B2(n_29), .C1(n_30), .C2(n_14), .Y(n_33) );
endmodule