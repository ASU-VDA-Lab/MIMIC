module real_aes_7756_n_103 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_103);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_103;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_555;
wire n_421;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_376;
wire n_571;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_744;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_746;
wire n_178;
wire n_409;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_449;
wire n_754;
wire n_417;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_434;
wire n_502;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_756;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_735;
wire n_713;
wire n_728;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_749;
wire n_358;
wire n_275;
wire n_214;
wire n_385;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_637;
wire n_526;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_420;
wire n_349;
wire n_336;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_753;
wire n_741;
wire n_283;
wire n_252;
wire n_314;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_424;
wire n_225;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
INVx1_ASAP7_75t_L g113 ( .A(n_0), .Y(n_113) );
INVx1_ASAP7_75t_L g497 ( .A(n_1), .Y(n_497) );
INVx1_ASAP7_75t_L g211 ( .A(n_2), .Y(n_211) );
AOI22xp5_ASAP7_75t_L g754 ( .A1(n_3), .A2(n_80), .B1(n_755), .B2(n_756), .Y(n_754) );
CKINVDCx20_ASAP7_75t_R g756 ( .A(n_3), .Y(n_756) );
AOI22xp33_ASAP7_75t_L g523 ( .A1(n_4), .A2(n_40), .B1(n_167), .B2(n_513), .Y(n_523) );
AOI21xp33_ASAP7_75t_L g191 ( .A1(n_5), .A2(n_148), .B(n_192), .Y(n_191) );
NAND2xp5_ASAP7_75t_L g488 ( .A(n_6), .B(n_141), .Y(n_488) );
AND2x6_ASAP7_75t_L g153 ( .A(n_7), .B(n_154), .Y(n_153) );
AOI21xp5_ASAP7_75t_L g249 ( .A1(n_8), .A2(n_250), .B(n_251), .Y(n_249) );
NOR2xp33_ASAP7_75t_L g114 ( .A(n_9), .B(n_41), .Y(n_114) );
INVx1_ASAP7_75t_L g198 ( .A(n_10), .Y(n_198) );
NAND2xp5_ASAP7_75t_L g241 ( .A(n_11), .B(n_242), .Y(n_241) );
INVx1_ASAP7_75t_L g146 ( .A(n_12), .Y(n_146) );
INVx1_ASAP7_75t_L g492 ( .A(n_13), .Y(n_492) );
INVx1_ASAP7_75t_L g256 ( .A(n_14), .Y(n_256) );
NAND2xp5_ASAP7_75t_L g508 ( .A(n_15), .B(n_179), .Y(n_508) );
CKINVDCx20_ASAP7_75t_R g123 ( .A(n_16), .Y(n_123) );
NAND2xp5_ASAP7_75t_L g469 ( .A(n_17), .B(n_142), .Y(n_469) );
AO32x2_ASAP7_75t_L g521 ( .A1(n_18), .A2(n_141), .A3(n_176), .B1(n_475), .B2(n_522), .Y(n_521) );
NAND2xp5_ASAP7_75t_SL g511 ( .A(n_19), .B(n_167), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g267 ( .A(n_20), .B(n_162), .Y(n_267) );
NAND2xp5_ASAP7_75t_L g499 ( .A(n_21), .B(n_142), .Y(n_499) );
AOI22xp33_ASAP7_75t_L g524 ( .A1(n_22), .A2(n_53), .B1(n_167), .B2(n_513), .Y(n_524) );
NAND2xp5_ASAP7_75t_SL g222 ( .A(n_23), .B(n_148), .Y(n_222) );
AOI22xp33_ASAP7_75t_SL g519 ( .A1(n_24), .A2(n_77), .B1(n_167), .B2(n_179), .Y(n_519) );
NAND2xp5_ASAP7_75t_SL g534 ( .A(n_25), .B(n_167), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g169 ( .A(n_26), .B(n_170), .Y(n_169) );
A2O1A1Ixp33_ASAP7_75t_L g253 ( .A1(n_27), .A2(n_254), .B(n_255), .C(n_257), .Y(n_253) );
BUFx6f_ASAP7_75t_L g152 ( .A(n_28), .Y(n_152) );
NAND2xp5_ASAP7_75t_L g557 ( .A(n_29), .B(n_200), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g213 ( .A(n_30), .B(n_196), .Y(n_213) );
AOI222xp33_ASAP7_75t_SL g124 ( .A1(n_31), .A2(n_125), .B1(n_131), .B2(n_739), .C1(n_740), .C2(n_745), .Y(n_124) );
OAI22xp5_ASAP7_75t_L g126 ( .A1(n_32), .A2(n_44), .B1(n_127), .B2(n_128), .Y(n_126) );
CKINVDCx20_ASAP7_75t_R g127 ( .A(n_32), .Y(n_127) );
INVx1_ASAP7_75t_L g185 ( .A(n_33), .Y(n_185) );
AOI22xp33_ASAP7_75t_L g103 ( .A1(n_34), .A2(n_104), .B1(n_115), .B2(n_760), .Y(n_103) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_35), .B(n_200), .Y(n_536) );
INVx2_ASAP7_75t_L g151 ( .A(n_36), .Y(n_151) );
NAND2xp5_ASAP7_75t_SL g552 ( .A(n_37), .B(n_167), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_38), .B(n_200), .Y(n_514) );
A2O1A1Ixp33_ASAP7_75t_L g223 ( .A1(n_39), .A2(n_153), .B(n_157), .C(n_224), .Y(n_223) );
INVx1_ASAP7_75t_L g183 ( .A(n_42), .Y(n_183) );
NAND2xp5_ASAP7_75t_SL g266 ( .A(n_43), .B(n_196), .Y(n_266) );
CKINVDCx14_ASAP7_75t_R g128 ( .A(n_44), .Y(n_128) );
NAND2xp5_ASAP7_75t_SL g482 ( .A(n_45), .B(n_167), .Y(n_482) );
OAI22xp5_ASAP7_75t_SL g125 ( .A1(n_46), .A2(n_126), .B1(n_129), .B2(n_130), .Y(n_125) );
CKINVDCx20_ASAP7_75t_R g130 ( .A(n_46), .Y(n_130) );
AOI22xp33_ASAP7_75t_L g518 ( .A1(n_47), .A2(n_88), .B1(n_229), .B2(n_513), .Y(n_518) );
NAND2xp5_ASAP7_75t_SL g485 ( .A(n_48), .B(n_167), .Y(n_485) );
NAND2xp5_ASAP7_75t_L g493 ( .A(n_49), .B(n_167), .Y(n_493) );
CKINVDCx16_ASAP7_75t_R g186 ( .A(n_50), .Y(n_186) );
NAND2xp5_ASAP7_75t_L g486 ( .A(n_51), .B(n_487), .Y(n_486) );
NAND2xp5_ASAP7_75t_L g244 ( .A(n_52), .B(n_148), .Y(n_244) );
AOI22xp33_ASAP7_75t_SL g474 ( .A1(n_54), .A2(n_63), .B1(n_167), .B2(n_179), .Y(n_474) );
AOI22xp5_ASAP7_75t_L g178 ( .A1(n_55), .A2(n_157), .B1(n_179), .B2(n_181), .Y(n_178) );
CKINVDCx20_ASAP7_75t_R g232 ( .A(n_56), .Y(n_232) );
NAND2xp5_ASAP7_75t_SL g507 ( .A(n_57), .B(n_167), .Y(n_507) );
CKINVDCx16_ASAP7_75t_R g208 ( .A(n_58), .Y(n_208) );
NAND2xp5_ASAP7_75t_SL g556 ( .A(n_59), .B(n_167), .Y(n_556) );
A2O1A1Ixp33_ASAP7_75t_L g194 ( .A1(n_60), .A2(n_166), .B(n_195), .C(n_197), .Y(n_194) );
CKINVDCx20_ASAP7_75t_R g270 ( .A(n_61), .Y(n_270) );
INVx1_ASAP7_75t_L g193 ( .A(n_62), .Y(n_193) );
INVx1_ASAP7_75t_L g154 ( .A(n_64), .Y(n_154) );
NAND2xp5_ASAP7_75t_L g498 ( .A(n_65), .B(n_167), .Y(n_498) );
INVx1_ASAP7_75t_L g145 ( .A(n_66), .Y(n_145) );
CKINVDCx20_ASAP7_75t_R g119 ( .A(n_67), .Y(n_119) );
AO32x2_ASAP7_75t_L g516 ( .A1(n_68), .A2(n_141), .A3(n_236), .B1(n_475), .B2(n_517), .Y(n_516) );
INVx1_ASAP7_75t_L g555 ( .A(n_69), .Y(n_555) );
INVx1_ASAP7_75t_L g531 ( .A(n_70), .Y(n_531) );
A2O1A1Ixp33_ASAP7_75t_SL g161 ( .A1(n_71), .A2(n_162), .B(n_163), .C(n_166), .Y(n_161) );
INVxp67_ASAP7_75t_L g164 ( .A(n_72), .Y(n_164) );
NAND2xp5_ASAP7_75t_SL g532 ( .A(n_73), .B(n_179), .Y(n_532) );
INVx1_ASAP7_75t_L g107 ( .A(n_74), .Y(n_107) );
CKINVDCx20_ASAP7_75t_R g189 ( .A(n_75), .Y(n_189) );
INVx1_ASAP7_75t_L g263 ( .A(n_76), .Y(n_263) );
A2O1A1Ixp33_ASAP7_75t_L g264 ( .A1(n_78), .A2(n_153), .B(n_157), .C(n_265), .Y(n_264) );
NAND2xp5_ASAP7_75t_L g512 ( .A(n_79), .B(n_513), .Y(n_512) );
CKINVDCx20_ASAP7_75t_R g755 ( .A(n_80), .Y(n_755) );
NAND2xp5_ASAP7_75t_SL g535 ( .A(n_81), .B(n_179), .Y(n_535) );
NAND2xp5_ASAP7_75t_SL g225 ( .A(n_82), .B(n_212), .Y(n_225) );
INVx2_ASAP7_75t_L g143 ( .A(n_83), .Y(n_143) );
NAND2xp5_ASAP7_75t_L g226 ( .A(n_84), .B(n_162), .Y(n_226) );
NAND2xp5_ASAP7_75t_L g483 ( .A(n_85), .B(n_179), .Y(n_483) );
A2O1A1Ixp33_ASAP7_75t_L g209 ( .A1(n_86), .A2(n_153), .B(n_157), .C(n_210), .Y(n_209) );
INVx2_ASAP7_75t_L g110 ( .A(n_87), .Y(n_110) );
OR2x2_ASAP7_75t_L g122 ( .A(n_87), .B(n_111), .Y(n_122) );
OR2x2_ASAP7_75t_L g460 ( .A(n_87), .B(n_112), .Y(n_460) );
AOI22xp33_ASAP7_75t_L g472 ( .A1(n_89), .A2(n_102), .B1(n_179), .B2(n_180), .Y(n_472) );
NAND2xp5_ASAP7_75t_L g199 ( .A(n_90), .B(n_200), .Y(n_199) );
CKINVDCx20_ASAP7_75t_R g216 ( .A(n_91), .Y(n_216) );
A2O1A1Ixp33_ASAP7_75t_L g238 ( .A1(n_92), .A2(n_153), .B(n_157), .C(n_239), .Y(n_238) );
CKINVDCx20_ASAP7_75t_R g246 ( .A(n_93), .Y(n_246) );
INVx1_ASAP7_75t_L g160 ( .A(n_94), .Y(n_160) );
CKINVDCx16_ASAP7_75t_R g252 ( .A(n_95), .Y(n_252) );
NAND2xp5_ASAP7_75t_SL g240 ( .A(n_96), .B(n_212), .Y(n_240) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_97), .B(n_179), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g258 ( .A(n_98), .B(n_141), .Y(n_258) );
NAND2xp5_ASAP7_75t_L g106 ( .A(n_99), .B(n_107), .Y(n_106) );
AOI21xp5_ASAP7_75t_L g147 ( .A1(n_100), .A2(n_148), .B(n_155), .Y(n_147) );
OAI22xp5_ASAP7_75t_SL g752 ( .A1(n_101), .A2(n_753), .B1(n_754), .B2(n_757), .Y(n_752) );
CKINVDCx20_ASAP7_75t_R g757 ( .A(n_101), .Y(n_757) );
INVx1_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
INVx1_ASAP7_75t_L g761 ( .A(n_105), .Y(n_761) );
OR2x2_ASAP7_75t_L g105 ( .A(n_106), .B(n_108), .Y(n_105) );
INVx3_ASAP7_75t_SL g108 ( .A(n_109), .Y(n_108) );
INVx2_ASAP7_75t_L g746 ( .A(n_109), .Y(n_746) );
NOR2x2_ASAP7_75t_L g109 ( .A(n_110), .B(n_111), .Y(n_109) );
OR2x2_ASAP7_75t_L g461 ( .A(n_110), .B(n_112), .Y(n_461) );
INVx2_ASAP7_75t_L g111 ( .A(n_112), .Y(n_111) );
AND2x2_ASAP7_75t_L g112 ( .A(n_113), .B(n_114), .Y(n_112) );
AOI22x1_ASAP7_75t_L g115 ( .A1(n_116), .A2(n_124), .B1(n_747), .B2(n_749), .Y(n_115) );
NOR2xp33_ASAP7_75t_L g116 ( .A(n_117), .B(n_120), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
BUFx2_ASAP7_75t_L g748 ( .A(n_118), .Y(n_748) );
INVx2_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
AOI21xp5_ASAP7_75t_L g749 ( .A1(n_120), .A2(n_750), .B(n_758), .Y(n_749) );
NOR2xp33_ASAP7_75t_SL g120 ( .A(n_121), .B(n_123), .Y(n_120) );
HB1xp67_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
INVx1_ASAP7_75t_SL g759 ( .A(n_122), .Y(n_759) );
CKINVDCx14_ASAP7_75t_R g739 ( .A(n_125), .Y(n_739) );
INVx1_ASAP7_75t_L g129 ( .A(n_126), .Y(n_129) );
OAI22x1_ASAP7_75t_SL g131 ( .A1(n_132), .A2(n_458), .B1(n_461), .B2(n_462), .Y(n_131) );
OAI22xp5_ASAP7_75t_L g750 ( .A1(n_132), .A2(n_133), .B1(n_751), .B2(n_752), .Y(n_750) );
INVx1_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
OAI22xp5_ASAP7_75t_L g740 ( .A1(n_133), .A2(n_741), .B1(n_742), .B2(n_744), .Y(n_740) );
AND2x2_ASAP7_75t_SL g133 ( .A(n_134), .B(n_395), .Y(n_133) );
NOR4xp25_ASAP7_75t_L g134 ( .A(n_135), .B(n_325), .C(n_356), .D(n_375), .Y(n_134) );
NAND4xp25_ASAP7_75t_L g135 ( .A(n_136), .B(n_283), .C(n_298), .D(n_316), .Y(n_135) );
AOI222xp33_ASAP7_75t_L g136 ( .A1(n_137), .A2(n_218), .B1(n_259), .B2(n_271), .C1(n_276), .C2(n_278), .Y(n_136) );
NAND2xp5_ASAP7_75t_L g137 ( .A(n_138), .B(n_201), .Y(n_137) );
INVx1_ASAP7_75t_L g339 ( .A(n_138), .Y(n_339) );
NAND2xp5_ASAP7_75t_L g138 ( .A(n_139), .B(n_172), .Y(n_138) );
AND2x2_ASAP7_75t_L g202 ( .A(n_139), .B(n_190), .Y(n_202) );
NAND2xp5_ASAP7_75t_L g368 ( .A(n_139), .B(n_205), .Y(n_368) );
INVx3_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
OR2x2_ASAP7_75t_L g275 ( .A(n_140), .B(n_174), .Y(n_275) );
AND2x2_ASAP7_75t_L g284 ( .A(n_140), .B(n_285), .Y(n_284) );
INVx1_ASAP7_75t_L g310 ( .A(n_140), .Y(n_310) );
AND2x2_ASAP7_75t_L g331 ( .A(n_140), .B(n_174), .Y(n_331) );
BUFx2_ASAP7_75t_L g354 ( .A(n_140), .Y(n_354) );
AND2x2_ASAP7_75t_L g378 ( .A(n_140), .B(n_175), .Y(n_378) );
AND2x2_ASAP7_75t_L g442 ( .A(n_140), .B(n_190), .Y(n_442) );
OA21x2_ASAP7_75t_L g140 ( .A1(n_141), .A2(n_147), .B(n_169), .Y(n_140) );
INVx4_ASAP7_75t_L g171 ( .A(n_141), .Y(n_171) );
OA21x2_ASAP7_75t_L g479 ( .A1(n_141), .A2(n_480), .B(n_488), .Y(n_479) );
BUFx6f_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
INVx1_ASAP7_75t_L g176 ( .A(n_142), .Y(n_176) );
AND2x2_ASAP7_75t_L g142 ( .A(n_143), .B(n_144), .Y(n_142) );
AND2x2_ASAP7_75t_SL g200 ( .A(n_143), .B(n_144), .Y(n_200) );
NAND2xp5_ASAP7_75t_L g144 ( .A(n_145), .B(n_146), .Y(n_144) );
BUFx2_ASAP7_75t_L g250 ( .A(n_148), .Y(n_250) );
AND2x4_ASAP7_75t_L g148 ( .A(n_149), .B(n_153), .Y(n_148) );
NAND2x1p5_ASAP7_75t_L g187 ( .A(n_149), .B(n_153), .Y(n_187) );
AND2x2_ASAP7_75t_L g149 ( .A(n_150), .B(n_152), .Y(n_149) );
INVx1_ASAP7_75t_L g487 ( .A(n_150), .Y(n_487) );
INVx1_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
INVx2_ASAP7_75t_L g158 ( .A(n_151), .Y(n_158) );
INVx1_ASAP7_75t_L g180 ( .A(n_151), .Y(n_180) );
INVx1_ASAP7_75t_L g159 ( .A(n_152), .Y(n_159) );
INVx1_ASAP7_75t_L g162 ( .A(n_152), .Y(n_162) );
INVx3_ASAP7_75t_L g165 ( .A(n_152), .Y(n_165) );
BUFx6f_ASAP7_75t_L g182 ( .A(n_152), .Y(n_182) );
BUFx6f_ASAP7_75t_L g196 ( .A(n_152), .Y(n_196) );
INVx4_ASAP7_75t_SL g168 ( .A(n_153), .Y(n_168) );
BUFx3_ASAP7_75t_L g475 ( .A(n_153), .Y(n_475) );
OAI21xp5_ASAP7_75t_L g480 ( .A1(n_153), .A2(n_481), .B(n_484), .Y(n_480) );
OAI21xp5_ASAP7_75t_L g490 ( .A1(n_153), .A2(n_491), .B(n_495), .Y(n_490) );
OAI21xp5_ASAP7_75t_L g505 ( .A1(n_153), .A2(n_506), .B(n_510), .Y(n_505) );
OAI21xp5_ASAP7_75t_L g529 ( .A1(n_153), .A2(n_530), .B(n_533), .Y(n_529) );
O2A1O1Ixp33_ASAP7_75t_L g155 ( .A1(n_156), .A2(n_160), .B(n_161), .C(n_168), .Y(n_155) );
O2A1O1Ixp33_ASAP7_75t_L g192 ( .A1(n_156), .A2(n_168), .B(n_193), .C(n_194), .Y(n_192) );
O2A1O1Ixp33_ASAP7_75t_L g251 ( .A1(n_156), .A2(n_168), .B(n_252), .C(n_253), .Y(n_251) );
INVx5_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
AND2x6_ASAP7_75t_L g157 ( .A(n_158), .B(n_159), .Y(n_157) );
BUFx6f_ASAP7_75t_L g167 ( .A(n_158), .Y(n_167) );
BUFx3_ASAP7_75t_L g229 ( .A(n_158), .Y(n_229) );
INVx1_ASAP7_75t_L g513 ( .A(n_158), .Y(n_513) );
INVx1_ASAP7_75t_L g509 ( .A(n_162), .Y(n_509) );
NOR2xp33_ASAP7_75t_L g163 ( .A(n_164), .B(n_165), .Y(n_163) );
NOR2xp33_ASAP7_75t_L g197 ( .A(n_165), .B(n_198), .Y(n_197) );
INVx5_ASAP7_75t_L g212 ( .A(n_165), .Y(n_212) );
OAI22xp5_ASAP7_75t_SL g517 ( .A1(n_165), .A2(n_196), .B1(n_518), .B2(n_519), .Y(n_517) );
O2A1O1Ixp5_ASAP7_75t_SL g530 ( .A1(n_166), .A2(n_212), .B(n_531), .C(n_532), .Y(n_530) );
INVx3_ASAP7_75t_L g166 ( .A(n_167), .Y(n_166) );
HB1xp67_ASAP7_75t_L g243 ( .A(n_167), .Y(n_243) );
OAI22xp33_ASAP7_75t_L g177 ( .A1(n_168), .A2(n_178), .B1(n_186), .B2(n_187), .Y(n_177) );
OA21x2_ASAP7_75t_L g190 ( .A1(n_170), .A2(n_191), .B(n_199), .Y(n_190) );
INVx3_ASAP7_75t_L g170 ( .A(n_171), .Y(n_170) );
NOR2xp33_ASAP7_75t_SL g231 ( .A(n_171), .B(n_232), .Y(n_231) );
NAND3xp33_ASAP7_75t_L g470 ( .A(n_171), .B(n_471), .C(n_475), .Y(n_470) );
AO21x1_ASAP7_75t_L g563 ( .A1(n_171), .A2(n_471), .B(n_564), .Y(n_563) );
AND2x2_ASAP7_75t_L g343 ( .A(n_172), .B(n_274), .Y(n_343) );
INVx1_ASAP7_75t_L g172 ( .A(n_173), .Y(n_172) );
NOR2xp33_ASAP7_75t_L g367 ( .A(n_173), .B(n_368), .Y(n_367) );
OR2x2_ASAP7_75t_L g173 ( .A(n_174), .B(n_190), .Y(n_173) );
OR2x2_ASAP7_75t_L g303 ( .A(n_174), .B(n_206), .Y(n_303) );
AND2x2_ASAP7_75t_L g315 ( .A(n_174), .B(n_274), .Y(n_315) );
BUFx2_ASAP7_75t_L g447 ( .A(n_174), .Y(n_447) );
INVx3_ASAP7_75t_L g174 ( .A(n_175), .Y(n_174) );
OR2x2_ASAP7_75t_L g204 ( .A(n_175), .B(n_205), .Y(n_204) );
AND2x2_ASAP7_75t_L g297 ( .A(n_175), .B(n_206), .Y(n_297) );
AND2x2_ASAP7_75t_L g350 ( .A(n_175), .B(n_190), .Y(n_350) );
HB1xp67_ASAP7_75t_L g386 ( .A(n_175), .Y(n_386) );
AO21x2_ASAP7_75t_L g175 ( .A1(n_176), .A2(n_177), .B(n_188), .Y(n_175) );
NOR2xp33_ASAP7_75t_L g188 ( .A(n_176), .B(n_189), .Y(n_188) );
AO21x2_ASAP7_75t_L g206 ( .A1(n_176), .A2(n_207), .B(n_215), .Y(n_206) );
INVx2_ASAP7_75t_L g230 ( .A(n_176), .Y(n_230) );
INVx2_ASAP7_75t_L g214 ( .A(n_179), .Y(n_214) );
INVx3_ASAP7_75t_L g179 ( .A(n_180), .Y(n_179) );
OAI22xp5_ASAP7_75t_SL g181 ( .A1(n_182), .A2(n_183), .B1(n_184), .B2(n_185), .Y(n_181) );
INVx2_ASAP7_75t_L g184 ( .A(n_182), .Y(n_184) );
INVx4_ASAP7_75t_L g254 ( .A(n_182), .Y(n_254) );
OAI21xp5_ASAP7_75t_L g207 ( .A1(n_187), .A2(n_208), .B(n_209), .Y(n_207) );
OAI21xp5_ASAP7_75t_L g262 ( .A1(n_187), .A2(n_263), .B(n_264), .Y(n_262) );
AND2x2_ASAP7_75t_L g273 ( .A(n_190), .B(n_274), .Y(n_273) );
INVx1_ASAP7_75t_SL g285 ( .A(n_190), .Y(n_285) );
INVx2_ASAP7_75t_L g296 ( .A(n_190), .Y(n_296) );
BUFx2_ASAP7_75t_L g320 ( .A(n_190), .Y(n_320) );
AND2x2_ASAP7_75t_SL g377 ( .A(n_190), .B(n_378), .Y(n_377) );
AOI21xp5_ASAP7_75t_L g510 ( .A1(n_195), .A2(n_511), .B(n_512), .Y(n_510) );
O2A1O1Ixp5_ASAP7_75t_L g554 ( .A1(n_195), .A2(n_496), .B(n_555), .C(n_556), .Y(n_554) );
INVx2_ASAP7_75t_L g195 ( .A(n_196), .Y(n_195) );
INVx4_ASAP7_75t_L g242 ( .A(n_196), .Y(n_242) );
OAI22xp5_ASAP7_75t_L g471 ( .A1(n_196), .A2(n_472), .B1(n_473), .B2(n_474), .Y(n_471) );
OAI22xp5_ASAP7_75t_L g522 ( .A1(n_196), .A2(n_473), .B1(n_523), .B2(n_524), .Y(n_522) );
INVx1_ASAP7_75t_L g217 ( .A(n_200), .Y(n_217) );
INVx2_ASAP7_75t_L g236 ( .A(n_200), .Y(n_236) );
OA21x2_ASAP7_75t_L g248 ( .A1(n_200), .A2(n_249), .B(n_258), .Y(n_248) );
OA21x2_ASAP7_75t_L g504 ( .A1(n_200), .A2(n_505), .B(n_514), .Y(n_504) );
OA21x2_ASAP7_75t_L g528 ( .A1(n_200), .A2(n_529), .B(n_536), .Y(n_528) );
NAND2xp5_ASAP7_75t_L g201 ( .A(n_202), .B(n_203), .Y(n_201) );
AOI332xp33_ASAP7_75t_L g298 ( .A1(n_202), .A2(n_299), .A3(n_303), .B1(n_304), .B2(n_308), .B3(n_311), .C1(n_312), .C2(n_314), .Y(n_298) );
NAND2x1_ASAP7_75t_L g383 ( .A(n_202), .B(n_274), .Y(n_383) );
NAND2xp5_ASAP7_75t_L g434 ( .A(n_202), .B(n_288), .Y(n_434) );
A2O1A1Ixp33_ASAP7_75t_SL g316 ( .A1(n_203), .A2(n_317), .B(n_320), .C(n_321), .Y(n_316) );
AND2x2_ASAP7_75t_L g455 ( .A(n_203), .B(n_296), .Y(n_455) );
INVx3_ASAP7_75t_SL g203 ( .A(n_204), .Y(n_203) );
OR2x2_ASAP7_75t_L g352 ( .A(n_204), .B(n_353), .Y(n_352) );
OR2x2_ASAP7_75t_L g357 ( .A(n_204), .B(n_354), .Y(n_357) );
INVx1_ASAP7_75t_L g288 ( .A(n_205), .Y(n_288) );
AND2x2_ASAP7_75t_L g391 ( .A(n_205), .B(n_350), .Y(n_391) );
AND2x2_ASAP7_75t_L g392 ( .A(n_205), .B(n_331), .Y(n_392) );
NAND2xp5_ASAP7_75t_L g401 ( .A(n_205), .B(n_402), .Y(n_401) );
NAND2xp5_ASAP7_75t_L g417 ( .A(n_205), .B(n_309), .Y(n_417) );
INVx3_ASAP7_75t_L g205 ( .A(n_206), .Y(n_205) );
INVx3_ASAP7_75t_L g274 ( .A(n_206), .Y(n_274) );
O2A1O1Ixp33_ASAP7_75t_L g210 ( .A1(n_211), .A2(n_212), .B(n_213), .C(n_214), .Y(n_210) );
INVx2_ASAP7_75t_L g473 ( .A(n_212), .Y(n_473) );
AOI21xp5_ASAP7_75t_L g481 ( .A1(n_212), .A2(n_482), .B(n_483), .Y(n_481) );
AOI21xp5_ASAP7_75t_L g551 ( .A1(n_212), .A2(n_552), .B(n_553), .Y(n_551) );
O2A1O1Ixp33_ASAP7_75t_L g491 ( .A1(n_214), .A2(n_492), .B(n_493), .C(n_494), .Y(n_491) );
NOR2xp33_ASAP7_75t_L g215 ( .A(n_216), .B(n_217), .Y(n_215) );
NOR2xp33_ASAP7_75t_L g245 ( .A(n_217), .B(n_246), .Y(n_245) );
NOR2xp33_ASAP7_75t_L g269 ( .A(n_217), .B(n_270), .Y(n_269) );
OAI31xp33_ASAP7_75t_L g456 ( .A1(n_218), .A2(n_377), .A3(n_384), .B(n_457), .Y(n_456) );
AND2x2_ASAP7_75t_L g218 ( .A(n_219), .B(n_233), .Y(n_218) );
AND2x2_ASAP7_75t_L g259 ( .A(n_219), .B(n_260), .Y(n_259) );
NAND2x1_ASAP7_75t_SL g279 ( .A(n_219), .B(n_280), .Y(n_279) );
HB1xp67_ASAP7_75t_L g366 ( .A(n_219), .Y(n_366) );
AND2x2_ASAP7_75t_L g371 ( .A(n_219), .B(n_282), .Y(n_371) );
INVx3_ASAP7_75t_L g219 ( .A(n_220), .Y(n_219) );
A2O1A1Ixp33_ASAP7_75t_L g283 ( .A1(n_220), .A2(n_284), .B(n_286), .C(n_289), .Y(n_283) );
OR2x2_ASAP7_75t_L g300 ( .A(n_220), .B(n_301), .Y(n_300) );
INVx1_ASAP7_75t_L g313 ( .A(n_220), .Y(n_313) );
AND2x2_ASAP7_75t_L g319 ( .A(n_220), .B(n_261), .Y(n_319) );
INVx2_ASAP7_75t_L g337 ( .A(n_220), .Y(n_337) );
AND2x2_ASAP7_75t_L g348 ( .A(n_220), .B(n_302), .Y(n_348) );
AND2x2_ASAP7_75t_L g380 ( .A(n_220), .B(n_338), .Y(n_380) );
AND2x2_ASAP7_75t_L g384 ( .A(n_220), .B(n_307), .Y(n_384) );
NAND2xp5_ASAP7_75t_L g389 ( .A(n_220), .B(n_233), .Y(n_389) );
AND2x2_ASAP7_75t_L g423 ( .A(n_220), .B(n_424), .Y(n_423) );
NOR2xp33_ASAP7_75t_L g457 ( .A(n_220), .B(n_326), .Y(n_457) );
OR2x6_ASAP7_75t_L g220 ( .A(n_221), .B(n_231), .Y(n_220) );
AOI21xp5_ASAP7_75t_SL g221 ( .A1(n_222), .A2(n_223), .B(n_230), .Y(n_221) );
AOI21xp5_ASAP7_75t_L g224 ( .A1(n_225), .A2(n_226), .B(n_227), .Y(n_224) );
AOI21xp5_ASAP7_75t_L g265 ( .A1(n_227), .A2(n_266), .B(n_267), .Y(n_265) );
INVx2_ASAP7_75t_L g227 ( .A(n_228), .Y(n_227) );
INVx2_ASAP7_75t_L g228 ( .A(n_229), .Y(n_228) );
INVx1_ASAP7_75t_L g257 ( .A(n_229), .Y(n_257) );
INVx1_ASAP7_75t_L g268 ( .A(n_230), .Y(n_268) );
OA21x2_ASAP7_75t_L g489 ( .A1(n_230), .A2(n_490), .B(n_499), .Y(n_489) );
OA21x2_ASAP7_75t_L g549 ( .A1(n_230), .A2(n_550), .B(n_557), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g287 ( .A(n_233), .B(n_288), .Y(n_287) );
INVx1_ASAP7_75t_L g365 ( .A(n_233), .Y(n_365) );
AND2x2_ASAP7_75t_L g427 ( .A(n_233), .B(n_348), .Y(n_427) );
AND2x2_ASAP7_75t_L g233 ( .A(n_234), .B(n_247), .Y(n_233) );
OR2x2_ASAP7_75t_L g281 ( .A(n_234), .B(n_282), .Y(n_281) );
AND2x2_ASAP7_75t_L g291 ( .A(n_234), .B(n_292), .Y(n_291) );
NAND2xp5_ASAP7_75t_L g301 ( .A(n_234), .B(n_302), .Y(n_301) );
INVx1_ASAP7_75t_L g399 ( .A(n_234), .Y(n_399) );
AND2x2_ASAP7_75t_L g416 ( .A(n_234), .B(n_261), .Y(n_416) );
INVx2_ASAP7_75t_L g234 ( .A(n_235), .Y(n_234) );
AND2x2_ASAP7_75t_L g307 ( .A(n_235), .B(n_247), .Y(n_307) );
AND2x2_ASAP7_75t_L g336 ( .A(n_235), .B(n_337), .Y(n_336) );
INVx1_ASAP7_75t_L g347 ( .A(n_235), .Y(n_347) );
NAND2xp5_ASAP7_75t_L g438 ( .A(n_235), .B(n_302), .Y(n_438) );
AO21x2_ASAP7_75t_L g235 ( .A1(n_236), .A2(n_237), .B(n_245), .Y(n_235) );
NAND2xp5_ASAP7_75t_L g237 ( .A(n_238), .B(n_244), .Y(n_237) );
AOI21xp5_ASAP7_75t_L g239 ( .A1(n_240), .A2(n_241), .B(n_243), .Y(n_239) );
INVx1_ASAP7_75t_L g247 ( .A(n_248), .Y(n_247) );
AND2x2_ASAP7_75t_L g260 ( .A(n_248), .B(n_261), .Y(n_260) );
INVx2_ASAP7_75t_L g282 ( .A(n_248), .Y(n_282) );
AND2x2_ASAP7_75t_L g338 ( .A(n_248), .B(n_302), .Y(n_338) );
NOR2xp33_ASAP7_75t_L g255 ( .A(n_254), .B(n_256), .Y(n_255) );
INVx1_ASAP7_75t_L g494 ( .A(n_254), .Y(n_494) );
AOI21xp5_ASAP7_75t_L g533 ( .A1(n_254), .A2(n_534), .B(n_535), .Y(n_533) );
INVx1_ASAP7_75t_L g440 ( .A(n_259), .Y(n_440) );
INVx1_ASAP7_75t_L g444 ( .A(n_260), .Y(n_444) );
INVx2_ASAP7_75t_L g302 ( .A(n_261), .Y(n_302) );
AO21x2_ASAP7_75t_L g261 ( .A1(n_262), .A2(n_268), .B(n_269), .Y(n_261) );
NOR2xp33_ASAP7_75t_L g271 ( .A(n_272), .B(n_275), .Y(n_271) );
INVx1_ASAP7_75t_SL g272 ( .A(n_273), .Y(n_272) );
NAND2xp5_ASAP7_75t_L g418 ( .A(n_273), .B(n_419), .Y(n_418) );
NAND2xp5_ASAP7_75t_L g436 ( .A(n_273), .B(n_378), .Y(n_436) );
OR2x2_ASAP7_75t_L g277 ( .A(n_274), .B(n_275), .Y(n_277) );
INVx1_ASAP7_75t_SL g329 ( .A(n_274), .Y(n_329) );
INVx1_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
INVx1_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
AOI221xp5_ASAP7_75t_L g332 ( .A1(n_280), .A2(n_333), .B1(n_335), .B2(n_339), .C(n_340), .Y(n_332) );
INVx2_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
OR2x2_ASAP7_75t_L g360 ( .A(n_281), .B(n_324), .Y(n_360) );
INVx2_ASAP7_75t_L g292 ( .A(n_282), .Y(n_292) );
INVx1_ASAP7_75t_L g318 ( .A(n_282), .Y(n_318) );
NAND2xp5_ASAP7_75t_L g326 ( .A(n_282), .B(n_302), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g412 ( .A(n_282), .B(n_305), .Y(n_412) );
INVx1_ASAP7_75t_L g420 ( .A(n_282), .Y(n_420) );
NAND2xp5_ASAP7_75t_L g334 ( .A(n_284), .B(n_288), .Y(n_334) );
AND2x4_ASAP7_75t_L g309 ( .A(n_285), .B(n_310), .Y(n_309) );
INVx1_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
AND2x2_ASAP7_75t_L g422 ( .A(n_288), .B(n_378), .Y(n_422) );
NOR2xp33_ASAP7_75t_L g289 ( .A(n_290), .B(n_293), .Y(n_289) );
INVx1_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
NAND2xp5_ASAP7_75t_L g322 ( .A(n_291), .B(n_323), .Y(n_322) );
INVxp67_ASAP7_75t_L g430 ( .A(n_292), .Y(n_430) );
INVxp67_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
AND2x2_ASAP7_75t_L g294 ( .A(n_295), .B(n_297), .Y(n_294) );
INVx1_ASAP7_75t_SL g295 ( .A(n_296), .Y(n_295) );
AND2x2_ASAP7_75t_L g330 ( .A(n_296), .B(n_331), .Y(n_330) );
AND2x2_ASAP7_75t_L g402 ( .A(n_296), .B(n_378), .Y(n_402) );
NAND2xp5_ASAP7_75t_L g408 ( .A(n_296), .B(n_315), .Y(n_408) );
AOI322xp5_ASAP7_75t_L g362 ( .A1(n_297), .A2(n_331), .A3(n_338), .B1(n_363), .B2(n_366), .C1(n_367), .C2(n_369), .Y(n_362) );
NAND2xp5_ASAP7_75t_L g405 ( .A(n_297), .B(n_406), .Y(n_405) );
INVx1_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
OR2x2_ASAP7_75t_L g428 ( .A(n_300), .B(n_429), .Y(n_428) );
INVx1_ASAP7_75t_L g374 ( .A(n_301), .Y(n_374) );
INVx2_ASAP7_75t_L g305 ( .A(n_302), .Y(n_305) );
INVx1_ASAP7_75t_L g364 ( .A(n_302), .Y(n_364) );
CKINVDCx16_ASAP7_75t_R g311 ( .A(n_303), .Y(n_311) );
NOR2xp33_ASAP7_75t_L g304 ( .A(n_305), .B(n_306), .Y(n_304) );
AND2x2_ASAP7_75t_L g400 ( .A(n_305), .B(n_313), .Y(n_400) );
INVx1_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
AND2x2_ASAP7_75t_L g312 ( .A(n_307), .B(n_313), .Y(n_312) );
AND2x2_ASAP7_75t_L g355 ( .A(n_307), .B(n_348), .Y(n_355) );
AND2x2_ASAP7_75t_L g359 ( .A(n_307), .B(n_319), .Y(n_359) );
OAI21xp33_ASAP7_75t_SL g369 ( .A1(n_308), .A2(n_370), .B(n_372), .Y(n_369) );
OAI22xp33_ASAP7_75t_L g439 ( .A1(n_308), .A2(n_440), .B1(n_441), .B2(n_443), .Y(n_439) );
INVx3_ASAP7_75t_SL g308 ( .A(n_309), .Y(n_308) );
AND2x2_ASAP7_75t_L g314 ( .A(n_309), .B(n_315), .Y(n_314) );
NAND2xp5_ASAP7_75t_L g341 ( .A(n_309), .B(n_329), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g448 ( .A(n_311), .B(n_449), .Y(n_448) );
AND2x2_ASAP7_75t_L g317 ( .A(n_318), .B(n_319), .Y(n_317) );
INVx1_ASAP7_75t_L g451 ( .A(n_318), .Y(n_451) );
INVx4_ASAP7_75t_L g324 ( .A(n_319), .Y(n_324) );
NAND2xp5_ASAP7_75t_L g394 ( .A(n_319), .B(n_346), .Y(n_394) );
INVx1_ASAP7_75t_SL g406 ( .A(n_320), .Y(n_406) );
INVx1_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
INVx1_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
NOR2xp67_ASAP7_75t_L g419 ( .A(n_324), .B(n_420), .Y(n_419) );
OAI211xp5_ASAP7_75t_SL g325 ( .A1(n_326), .A2(n_327), .B(n_332), .C(n_349), .Y(n_325) );
OAI221xp5_ASAP7_75t_SL g445 ( .A1(n_327), .A2(n_365), .B1(n_444), .B2(n_446), .C(n_448), .Y(n_445) );
INVx1_ASAP7_75t_SL g327 ( .A(n_328), .Y(n_327) );
AND2x2_ASAP7_75t_L g328 ( .A(n_329), .B(n_330), .Y(n_328) );
NAND2xp5_ASAP7_75t_L g441 ( .A(n_329), .B(n_442), .Y(n_441) );
OAI31xp33_ASAP7_75t_L g421 ( .A1(n_330), .A2(n_407), .A3(n_422), .B(n_423), .Y(n_421) );
INVx1_ASAP7_75t_L g361 ( .A(n_331), .Y(n_361) );
INVx1_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
AND2x2_ASAP7_75t_L g335 ( .A(n_336), .B(n_338), .Y(n_335) );
INVx1_ASAP7_75t_L g411 ( .A(n_336), .Y(n_411) );
AND2x2_ASAP7_75t_L g424 ( .A(n_338), .B(n_347), .Y(n_424) );
AOI21xp33_ASAP7_75t_L g340 ( .A1(n_341), .A2(n_342), .B(n_344), .Y(n_340) );
INVx1_ASAP7_75t_SL g342 ( .A(n_343), .Y(n_342) );
INVxp67_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
AND2x2_ASAP7_75t_L g345 ( .A(n_346), .B(n_348), .Y(n_345) );
INVx1_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
NAND2xp5_ASAP7_75t_L g450 ( .A(n_348), .B(n_451), .Y(n_450) );
OAI21xp33_ASAP7_75t_L g349 ( .A1(n_350), .A2(n_351), .B(n_355), .Y(n_349) );
INVx1_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
INVx1_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
OAI221xp5_ASAP7_75t_SL g356 ( .A1(n_357), .A2(n_358), .B1(n_360), .B2(n_361), .C(n_362), .Y(n_356) );
A2O1A1Ixp33_ASAP7_75t_L g425 ( .A1(n_357), .A2(n_426), .B(n_428), .C(n_431), .Y(n_425) );
CKINVDCx16_ASAP7_75t_R g358 ( .A(n_359), .Y(n_358) );
NAND2xp5_ASAP7_75t_SL g409 ( .A(n_360), .B(n_410), .Y(n_409) );
NOR2xp33_ASAP7_75t_L g363 ( .A(n_364), .B(n_365), .Y(n_363) );
INVx1_ASAP7_75t_L g387 ( .A(n_368), .Y(n_387) );
INVx1_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
AND2x2_ASAP7_75t_L g373 ( .A(n_371), .B(n_374), .Y(n_373) );
AND2x2_ASAP7_75t_L g415 ( .A(n_371), .B(n_416), .Y(n_415) );
INVx2_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
OAI211xp5_ASAP7_75t_L g375 ( .A1(n_376), .A2(n_379), .B(n_381), .C(n_390), .Y(n_375) );
INVx1_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
OAI221xp5_ASAP7_75t_L g452 ( .A1(n_379), .A2(n_389), .B1(n_453), .B2(n_454), .C(n_456), .Y(n_452) );
INVx1_ASAP7_75t_SL g379 ( .A(n_380), .Y(n_379) );
AOI22xp5_ASAP7_75t_L g381 ( .A1(n_382), .A2(n_384), .B1(n_385), .B2(n_388), .Y(n_381) );
INVx1_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
AND2x2_ASAP7_75t_L g385 ( .A(n_386), .B(n_387), .Y(n_385) );
INVx1_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
OAI21xp5_ASAP7_75t_SL g390 ( .A1(n_391), .A2(n_392), .B(n_393), .Y(n_390) );
INVx1_ASAP7_75t_SL g453 ( .A(n_392), .Y(n_453) );
INVxp67_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
NOR4xp25_ASAP7_75t_L g395 ( .A(n_396), .B(n_425), .C(n_445), .D(n_452), .Y(n_395) );
OAI211xp5_ASAP7_75t_L g396 ( .A1(n_397), .A2(n_401), .B(n_403), .C(n_421), .Y(n_396) );
NAND2xp5_ASAP7_75t_L g397 ( .A(n_398), .B(n_400), .Y(n_397) );
INVxp67_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
O2A1O1Ixp33_ASAP7_75t_L g403 ( .A1(n_404), .A2(n_407), .B(n_409), .C(n_413), .Y(n_403) );
INVx1_ASAP7_75t_SL g404 ( .A(n_405), .Y(n_404) );
INVx1_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
INVx1_ASAP7_75t_SL g432 ( .A(n_410), .Y(n_432) );
OR2x2_ASAP7_75t_L g410 ( .A(n_411), .B(n_412), .Y(n_410) );
OR2x2_ASAP7_75t_L g443 ( .A(n_411), .B(n_444), .Y(n_443) );
OAI21xp33_ASAP7_75t_L g413 ( .A1(n_414), .A2(n_417), .B(n_418), .Y(n_413) );
INVx1_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
INVx1_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
HB1xp67_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
AOI221xp5_ASAP7_75t_L g431 ( .A1(n_432), .A2(n_433), .B1(n_435), .B2(n_437), .C(n_439), .Y(n_431) );
INVx1_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
INVx1_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
INVxp67_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
NAND2xp5_ASAP7_75t_L g446 ( .A(n_442), .B(n_447), .Y(n_446) );
INVx1_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
INVx1_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
INVx2_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
INVx2_ASAP7_75t_L g741 ( .A(n_459), .Y(n_741) );
INVx1_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
INVx1_ASAP7_75t_L g743 ( .A(n_461), .Y(n_743) );
INVx1_ASAP7_75t_L g744 ( .A(n_462), .Y(n_744) );
INVx2_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
AND2x2_ASAP7_75t_SL g463 ( .A(n_464), .B(n_673), .Y(n_463) );
NOR5xp2_ASAP7_75t_L g464 ( .A(n_465), .B(n_586), .C(n_632), .D(n_645), .E(n_657), .Y(n_464) );
OAI211xp5_ASAP7_75t_L g465 ( .A1(n_466), .A2(n_500), .B(n_540), .C(n_567), .Y(n_465) );
INVx1_ASAP7_75t_SL g668 ( .A(n_466), .Y(n_668) );
OR2x2_ASAP7_75t_L g466 ( .A(n_467), .B(n_476), .Y(n_466) );
AND2x2_ASAP7_75t_L g592 ( .A(n_467), .B(n_477), .Y(n_592) );
AND2x2_ASAP7_75t_L g620 ( .A(n_467), .B(n_566), .Y(n_620) );
AND2x2_ASAP7_75t_L g628 ( .A(n_467), .B(n_571), .Y(n_628) );
INVx3_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
AND2x2_ASAP7_75t_L g558 ( .A(n_468), .B(n_478), .Y(n_558) );
INVx2_ASAP7_75t_L g570 ( .A(n_468), .Y(n_570) );
AND2x2_ASAP7_75t_L g695 ( .A(n_468), .B(n_637), .Y(n_695) );
OR2x2_ASAP7_75t_L g697 ( .A(n_468), .B(n_698), .Y(n_697) );
AND2x4_ASAP7_75t_L g468 ( .A(n_469), .B(n_470), .Y(n_468) );
INVx1_ASAP7_75t_L g564 ( .A(n_469), .Y(n_564) );
AOI21xp5_ASAP7_75t_L g484 ( .A1(n_473), .A2(n_485), .B(n_486), .Y(n_484) );
O2A1O1Ixp33_ASAP7_75t_L g495 ( .A1(n_473), .A2(n_496), .B(n_497), .C(n_498), .Y(n_495) );
OAI21xp5_ASAP7_75t_L g550 ( .A1(n_475), .A2(n_551), .B(n_554), .Y(n_550) );
INVx2_ASAP7_75t_SL g476 ( .A(n_477), .Y(n_476) );
AND2x2_ASAP7_75t_L g608 ( .A(n_477), .B(n_580), .Y(n_608) );
NOR2xp33_ASAP7_75t_L g636 ( .A(n_477), .B(n_637), .Y(n_636) );
AND2x2_ASAP7_75t_L g722 ( .A(n_477), .B(n_562), .Y(n_722) );
AND2x2_ASAP7_75t_L g477 ( .A(n_478), .B(n_489), .Y(n_477) );
AND2x2_ASAP7_75t_L g565 ( .A(n_478), .B(n_566), .Y(n_565) );
INVx2_ASAP7_75t_L g612 ( .A(n_478), .Y(n_612) );
AND2x2_ASAP7_75t_L g637 ( .A(n_478), .B(n_549), .Y(n_637) );
NAND2xp5_ASAP7_75t_L g707 ( .A(n_478), .B(n_670), .Y(n_707) );
INVx3_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
AND2x2_ASAP7_75t_L g571 ( .A(n_479), .B(n_549), .Y(n_571) );
AND2x2_ASAP7_75t_L g585 ( .A(n_479), .B(n_548), .Y(n_585) );
AND2x2_ASAP7_75t_L g602 ( .A(n_479), .B(n_489), .Y(n_602) );
AND2x2_ASAP7_75t_L g659 ( .A(n_479), .B(n_660), .Y(n_659) );
NAND2xp5_ASAP7_75t_L g672 ( .A(n_479), .B(n_566), .Y(n_672) );
AND2x2_ASAP7_75t_L g724 ( .A(n_479), .B(n_649), .Y(n_724) );
INVx2_ASAP7_75t_L g496 ( .A(n_487), .Y(n_496) );
AND2x2_ASAP7_75t_L g547 ( .A(n_489), .B(n_548), .Y(n_547) );
INVx2_ASAP7_75t_L g566 ( .A(n_489), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g643 ( .A(n_489), .B(n_549), .Y(n_643) );
AOI21xp5_ASAP7_75t_L g500 ( .A1(n_501), .A2(n_525), .B(n_537), .Y(n_500) );
INVx1_ASAP7_75t_SL g656 ( .A(n_501), .Y(n_656) );
AND2x4_ASAP7_75t_L g501 ( .A(n_502), .B(n_515), .Y(n_501) );
BUFx3_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
AND2x2_ASAP7_75t_SL g544 ( .A(n_503), .B(n_545), .Y(n_544) );
INVx1_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
INVx2_ASAP7_75t_L g539 ( .A(n_504), .Y(n_539) );
INVx1_ASAP7_75t_L g576 ( .A(n_504), .Y(n_576) );
AND2x2_ASAP7_75t_L g597 ( .A(n_504), .B(n_520), .Y(n_597) );
AND2x2_ASAP7_75t_L g631 ( .A(n_504), .B(n_521), .Y(n_631) );
OR2x2_ASAP7_75t_L g650 ( .A(n_504), .B(n_527), .Y(n_650) );
HB1xp67_ASAP7_75t_L g664 ( .A(n_504), .Y(n_664) );
AND2x2_ASAP7_75t_L g677 ( .A(n_504), .B(n_678), .Y(n_677) );
AOI21xp5_ASAP7_75t_L g506 ( .A1(n_507), .A2(n_508), .B(n_509), .Y(n_506) );
AOI22xp5_ASAP7_75t_L g598 ( .A1(n_515), .A2(n_599), .B1(n_600), .B2(n_609), .Y(n_598) );
AND2x2_ASAP7_75t_L g682 ( .A(n_515), .B(n_683), .Y(n_682) );
AND2x2_ASAP7_75t_L g515 ( .A(n_516), .B(n_520), .Y(n_515) );
INVx1_ASAP7_75t_L g543 ( .A(n_516), .Y(n_543) );
BUFx6f_ASAP7_75t_L g580 ( .A(n_516), .Y(n_580) );
INVx1_ASAP7_75t_L g591 ( .A(n_516), .Y(n_591) );
AND2x2_ASAP7_75t_L g606 ( .A(n_516), .B(n_521), .Y(n_606) );
OR2x2_ASAP7_75t_L g560 ( .A(n_520), .B(n_545), .Y(n_560) );
AND2x2_ASAP7_75t_L g590 ( .A(n_520), .B(n_591), .Y(n_590) );
NOR2xp67_ASAP7_75t_L g678 ( .A(n_520), .B(n_679), .Y(n_678) );
INVx2_ASAP7_75t_L g520 ( .A(n_521), .Y(n_520) );
AND2x2_ASAP7_75t_L g538 ( .A(n_521), .B(n_539), .Y(n_538) );
BUFx2_ASAP7_75t_L g647 ( .A(n_521), .Y(n_647) );
NAND2xp5_ASAP7_75t_L g662 ( .A(n_525), .B(n_663), .Y(n_662) );
BUFx2_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
AND2x2_ASAP7_75t_L g625 ( .A(n_526), .B(n_591), .Y(n_625) );
INVx2_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
AND2x2_ASAP7_75t_L g537 ( .A(n_527), .B(n_538), .Y(n_537) );
INVx1_ASAP7_75t_L g596 ( .A(n_527), .Y(n_596) );
INVx2_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
INVx2_ASAP7_75t_L g545 ( .A(n_528), .Y(n_545) );
OR2x2_ASAP7_75t_L g575 ( .A(n_528), .B(n_576), .Y(n_575) );
HB1xp67_ASAP7_75t_L g630 ( .A(n_528), .Y(n_630) );
AOI32xp33_ASAP7_75t_L g667 ( .A1(n_537), .A2(n_597), .A3(n_668), .B1(n_669), .B2(n_671), .Y(n_667) );
AND2x2_ASAP7_75t_L g593 ( .A(n_538), .B(n_594), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g691 ( .A(n_538), .B(n_692), .Y(n_691) );
NAND2xp5_ASAP7_75t_L g711 ( .A(n_538), .B(n_625), .Y(n_711) );
INVx1_ASAP7_75t_L g716 ( .A(n_538), .Y(n_716) );
AOI22xp5_ASAP7_75t_L g540 ( .A1(n_541), .A2(n_546), .B1(n_559), .B2(n_561), .Y(n_540) );
AND2x2_ASAP7_75t_L g541 ( .A(n_542), .B(n_544), .Y(n_541) );
AND2x2_ASAP7_75t_L g646 ( .A(n_542), .B(n_647), .Y(n_646) );
HB1xp67_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g690 ( .A(n_543), .B(n_545), .Y(n_690) );
AOI22xp5_ASAP7_75t_L g567 ( .A1(n_544), .A2(n_568), .B1(n_572), .B2(n_582), .Y(n_567) );
AND2x2_ASAP7_75t_L g589 ( .A(n_544), .B(n_590), .Y(n_589) );
A2O1A1Ixp33_ASAP7_75t_L g640 ( .A1(n_544), .A2(n_558), .B(n_606), .C(n_641), .Y(n_640) );
OAI332xp33_ASAP7_75t_L g645 ( .A1(n_544), .A2(n_646), .A3(n_648), .B1(n_650), .B2(n_651), .B3(n_653), .C1(n_654), .C2(n_656), .Y(n_645) );
INVx2_ASAP7_75t_L g686 ( .A(n_544), .Y(n_686) );
HB1xp67_ASAP7_75t_L g604 ( .A(n_545), .Y(n_604) );
INVx1_ASAP7_75t_L g679 ( .A(n_545), .Y(n_679) );
AND2x2_ASAP7_75t_L g733 ( .A(n_545), .B(n_597), .Y(n_733) );
AND2x2_ASAP7_75t_L g546 ( .A(n_547), .B(n_558), .Y(n_546) );
AND2x2_ASAP7_75t_L g613 ( .A(n_548), .B(n_563), .Y(n_613) );
INVx2_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
AND2x2_ASAP7_75t_L g562 ( .A(n_549), .B(n_563), .Y(n_562) );
OR2x2_ASAP7_75t_L g661 ( .A(n_549), .B(n_563), .Y(n_661) );
INVx1_ASAP7_75t_L g670 ( .A(n_549), .Y(n_670) );
INVx1_ASAP7_75t_L g644 ( .A(n_558), .Y(n_644) );
INVxp67_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
OR2x2_ASAP7_75t_L g728 ( .A(n_560), .B(n_580), .Y(n_728) );
INVx1_ASAP7_75t_SL g639 ( .A(n_561), .Y(n_639) );
AND2x2_ASAP7_75t_L g561 ( .A(n_562), .B(n_565), .Y(n_561) );
AND2x2_ASAP7_75t_L g666 ( .A(n_562), .B(n_624), .Y(n_666) );
INVx1_ASAP7_75t_L g685 ( .A(n_562), .Y(n_685) );
NAND2xp5_ASAP7_75t_SL g687 ( .A(n_562), .B(n_652), .Y(n_687) );
INVx1_ASAP7_75t_L g584 ( .A(n_563), .Y(n_584) );
AND2x2_ASAP7_75t_L g588 ( .A(n_565), .B(n_569), .Y(n_588) );
AND2x2_ASAP7_75t_L g655 ( .A(n_565), .B(n_613), .Y(n_655) );
INVx2_ASAP7_75t_L g698 ( .A(n_565), .Y(n_698) );
INVx2_ASAP7_75t_L g581 ( .A(n_566), .Y(n_581) );
AND2x2_ASAP7_75t_L g583 ( .A(n_566), .B(n_584), .Y(n_583) );
AND2x2_ASAP7_75t_L g568 ( .A(n_569), .B(n_571), .Y(n_568) );
INVx1_ASAP7_75t_L g599 ( .A(n_569), .Y(n_599) );
INVx2_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
NOR2xp33_ASAP7_75t_L g649 ( .A(n_570), .B(n_643), .Y(n_649) );
OR2x2_ASAP7_75t_L g713 ( .A(n_570), .B(n_672), .Y(n_713) );
INVx1_ASAP7_75t_L g737 ( .A(n_570), .Y(n_737) );
INVx1_ASAP7_75t_L g693 ( .A(n_571), .Y(n_693) );
AND2x2_ASAP7_75t_L g738 ( .A(n_571), .B(n_581), .Y(n_738) );
INVx1_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g573 ( .A(n_574), .B(n_577), .Y(n_573) );
INVx2_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
OAI22xp5_ASAP7_75t_L g600 ( .A1(n_575), .A2(n_601), .B1(n_603), .B2(n_607), .Y(n_600) );
INVx1_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
OAI322xp33_ASAP7_75t_SL g684 ( .A1(n_578), .A2(n_685), .A3(n_686), .B1(n_687), .B2(n_688), .C1(n_691), .C2(n_693), .Y(n_684) );
OR2x2_ASAP7_75t_L g578 ( .A(n_579), .B(n_581), .Y(n_578) );
AND2x2_ASAP7_75t_L g681 ( .A(n_579), .B(n_597), .Y(n_681) );
OR2x2_ASAP7_75t_L g715 ( .A(n_579), .B(n_716), .Y(n_715) );
OR2x2_ASAP7_75t_L g718 ( .A(n_579), .B(n_650), .Y(n_718) );
INVx2_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
AND2x2_ASAP7_75t_L g663 ( .A(n_580), .B(n_664), .Y(n_663) );
OR2x2_ASAP7_75t_L g719 ( .A(n_580), .B(n_650), .Y(n_719) );
INVx3_ASAP7_75t_L g652 ( .A(n_581), .Y(n_652) );
AND2x2_ASAP7_75t_L g582 ( .A(n_583), .B(n_585), .Y(n_582) );
INVx1_ASAP7_75t_L g708 ( .A(n_583), .Y(n_708) );
AOI222xp33_ASAP7_75t_L g587 ( .A1(n_585), .A2(n_588), .B1(n_589), .B2(n_592), .C1(n_593), .C2(n_595), .Y(n_587) );
INVx1_ASAP7_75t_L g618 ( .A(n_585), .Y(n_618) );
NAND3xp33_ASAP7_75t_SL g586 ( .A(n_587), .B(n_598), .C(n_615), .Y(n_586) );
AND2x2_ASAP7_75t_L g703 ( .A(n_590), .B(n_604), .Y(n_703) );
BUFx2_ASAP7_75t_L g594 ( .A(n_591), .Y(n_594) );
INVx1_ASAP7_75t_L g635 ( .A(n_591), .Y(n_635) );
AOI221xp5_ASAP7_75t_L g680 ( .A1(n_592), .A2(n_628), .B1(n_681), .B2(n_682), .C(n_684), .Y(n_680) );
NAND2xp5_ASAP7_75t_L g676 ( .A(n_594), .B(n_677), .Y(n_676) );
AND2x2_ASAP7_75t_L g595 ( .A(n_596), .B(n_597), .Y(n_595) );
HB1xp67_ASAP7_75t_L g621 ( .A(n_597), .Y(n_621) );
AND2x2_ASAP7_75t_L g634 ( .A(n_597), .B(n_635), .Y(n_634) );
INVx1_ASAP7_75t_SL g601 ( .A(n_602), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g614 ( .A(n_602), .B(n_613), .Y(n_614) );
OR2x2_ASAP7_75t_L g603 ( .A(n_604), .B(n_605), .Y(n_603) );
OAI21xp33_ASAP7_75t_L g609 ( .A1(n_604), .A2(n_610), .B(n_614), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g633 ( .A(n_604), .B(n_634), .Y(n_633) );
INVx1_ASAP7_75t_SL g605 ( .A(n_606), .Y(n_605) );
AND2x2_ASAP7_75t_L g701 ( .A(n_606), .B(n_683), .Y(n_701) );
INVx1_ASAP7_75t_L g607 ( .A(n_608), .Y(n_607) );
INVx1_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
AND2x2_ASAP7_75t_L g611 ( .A(n_612), .B(n_613), .Y(n_611) );
INVx1_ASAP7_75t_L g624 ( .A(n_612), .Y(n_624) );
NAND2xp5_ASAP7_75t_L g623 ( .A(n_613), .B(n_624), .Y(n_623) );
INVx2_ASAP7_75t_L g730 ( .A(n_613), .Y(n_730) );
AOI221xp5_ASAP7_75t_L g615 ( .A1(n_616), .A2(n_621), .B1(n_622), .B2(n_625), .C(n_626), .Y(n_615) );
INVx2_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
NAND2xp5_ASAP7_75t_SL g705 ( .A(n_617), .B(n_706), .Y(n_705) );
OR2x2_ASAP7_75t_L g617 ( .A(n_618), .B(n_619), .Y(n_617) );
INVx1_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
INVx1_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
AND2x2_ASAP7_75t_L g726 ( .A(n_625), .B(n_631), .Y(n_726) );
INVxp67_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
NAND2xp5_ASAP7_75t_L g627 ( .A(n_628), .B(n_629), .Y(n_627) );
OAI31xp33_ASAP7_75t_SL g694 ( .A1(n_629), .A2(n_668), .A3(n_695), .B(n_696), .Y(n_694) );
AND2x2_ASAP7_75t_L g629 ( .A(n_630), .B(n_631), .Y(n_629) );
INVx1_ASAP7_75t_L g683 ( .A(n_630), .Y(n_683) );
NAND2xp5_ASAP7_75t_SL g734 ( .A(n_631), .B(n_635), .Y(n_734) );
OAI221xp5_ASAP7_75t_SL g632 ( .A1(n_633), .A2(n_636), .B1(n_638), .B2(n_639), .C(n_640), .Y(n_632) );
INVx1_ASAP7_75t_L g638 ( .A(n_634), .Y(n_638) );
NAND2xp5_ASAP7_75t_L g651 ( .A(n_637), .B(n_652), .Y(n_651) );
INVx1_ASAP7_75t_L g641 ( .A(n_642), .Y(n_641) );
OR2x2_ASAP7_75t_L g642 ( .A(n_643), .B(n_644), .Y(n_642) );
INVx1_ASAP7_75t_L g653 ( .A(n_646), .Y(n_653) );
INVx2_ASAP7_75t_L g689 ( .A(n_647), .Y(n_689) );
INVx1_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
OR2x2_ASAP7_75t_L g675 ( .A(n_652), .B(n_661), .Y(n_675) );
A2O1A1Ixp33_ASAP7_75t_L g725 ( .A1(n_652), .A2(n_669), .B(n_726), .C(n_727), .Y(n_725) );
OAI221xp5_ASAP7_75t_SL g657 ( .A1(n_653), .A2(n_658), .B1(n_662), .B2(n_665), .C(n_667), .Y(n_657) );
INVx1_ASAP7_75t_SL g654 ( .A(n_655), .Y(n_654) );
A2O1A1Ixp33_ASAP7_75t_L g720 ( .A1(n_656), .A2(n_721), .B(n_723), .C(n_725), .Y(n_720) );
INVx1_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
AOI221xp5_ASAP7_75t_L g709 ( .A1(n_659), .A2(n_710), .B1(n_712), .B2(n_714), .C(n_717), .Y(n_709) );
INVx1_ASAP7_75t_SL g660 ( .A(n_661), .Y(n_660) );
INVx1_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
INVx1_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
INVx1_ASAP7_75t_SL g671 ( .A(n_672), .Y(n_671) );
NOR4xp25_ASAP7_75t_L g673 ( .A(n_674), .B(n_699), .C(n_720), .D(n_731), .Y(n_673) );
OAI211xp5_ASAP7_75t_SL g674 ( .A1(n_675), .A2(n_676), .B(n_680), .C(n_694), .Y(n_674) );
INVx1_ASAP7_75t_SL g729 ( .A(n_681), .Y(n_729) );
OR2x2_ASAP7_75t_L g688 ( .A(n_689), .B(n_690), .Y(n_688) );
INVx1_ASAP7_75t_SL g692 ( .A(n_690), .Y(n_692) );
INVx1_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
OAI22xp5_ASAP7_75t_L g717 ( .A1(n_697), .A2(n_706), .B1(n_718), .B2(n_719), .Y(n_717) );
A2O1A1Ixp33_ASAP7_75t_L g699 ( .A1(n_700), .A2(n_702), .B(n_704), .C(n_709), .Y(n_699) );
INVx1_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
AOI31xp33_ASAP7_75t_L g731 ( .A1(n_702), .A2(n_732), .A3(n_734), .B(n_735), .Y(n_731) );
INVx1_ASAP7_75t_L g702 ( .A(n_703), .Y(n_702) );
INVxp67_ASAP7_75t_L g704 ( .A(n_705), .Y(n_704) );
OR2x2_ASAP7_75t_L g706 ( .A(n_707), .B(n_708), .Y(n_706) );
INVx1_ASAP7_75t_L g710 ( .A(n_711), .Y(n_710) );
INVx1_ASAP7_75t_SL g712 ( .A(n_713), .Y(n_712) );
INVx1_ASAP7_75t_L g714 ( .A(n_715), .Y(n_714) );
INVx1_ASAP7_75t_L g721 ( .A(n_722), .Y(n_721) );
INVx1_ASAP7_75t_SL g723 ( .A(n_724), .Y(n_723) );
AOI21xp5_ASAP7_75t_L g727 ( .A1(n_728), .A2(n_729), .B(n_730), .Y(n_727) );
INVx1_ASAP7_75t_L g732 ( .A(n_733), .Y(n_732) );
NAND2xp5_ASAP7_75t_L g735 ( .A(n_736), .B(n_738), .Y(n_735) );
INVx1_ASAP7_75t_L g736 ( .A(n_737), .Y(n_736) );
INVx2_ASAP7_75t_L g742 ( .A(n_743), .Y(n_742) );
INVx2_ASAP7_75t_L g745 ( .A(n_746), .Y(n_745) );
INVx1_ASAP7_75t_SL g747 ( .A(n_748), .Y(n_747) );
CKINVDCx20_ASAP7_75t_R g751 ( .A(n_752), .Y(n_751) );
CKINVDCx20_ASAP7_75t_R g753 ( .A(n_754), .Y(n_753) );
INVx1_ASAP7_75t_SL g758 ( .A(n_759), .Y(n_758) );
INVx1_ASAP7_75t_L g760 ( .A(n_761), .Y(n_760) );
endmodule