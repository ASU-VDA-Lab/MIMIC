module real_aes_754_n_104 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_104);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_104;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_800;
wire n_778;
wire n_522;
wire n_485;
wire n_822;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_503;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_571;
wire n_376;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_453;
wire n_374;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_816;
wire n_292;
wire n_539;
wire n_400;
wire n_626;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_578;
wire n_528;
wire n_372;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_732;
wire n_834;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_781;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_812;
wire n_782;
wire n_443;
wire n_565;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_449;
wire n_417;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_733;
wire n_552;
wire n_402;
wire n_602;
wire n_617;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_807;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_832;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_569;
wire n_303;
wire n_563;
wire n_785;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_810;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_831;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_456;
wire n_359;
wire n_717;
wire n_312;
wire n_266;
wire n_183;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_521;
wire n_140;
wire n_418;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_829;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_710;
wire n_650;
wire n_105;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_802;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_554;
wire n_475;
wire n_264;
wire n_798;
wire n_237;
wire n_797;
wire n_668;
NAND2xp5_ASAP7_75t_SL g543 ( .A(n_0), .B(n_520), .Y(n_543) );
AOI21xp5_ASAP7_75t_L g587 ( .A1(n_1), .A2(n_523), .B(n_588), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g113 ( .A(n_2), .B(n_114), .Y(n_113) );
NAND2xp5_ASAP7_75t_SL g526 ( .A(n_3), .B(n_230), .Y(n_526) );
INVx1_ASAP7_75t_L g162 ( .A(n_4), .Y(n_162) );
XNOR2xp5_ASAP7_75t_L g131 ( .A(n_5), .B(n_132), .Y(n_131) );
NAND2xp5_ASAP7_75t_SL g218 ( .A(n_6), .B(n_219), .Y(n_218) );
NAND2xp5_ASAP7_75t_L g596 ( .A(n_7), .B(n_230), .Y(n_596) );
INVx1_ASAP7_75t_L g194 ( .A(n_8), .Y(n_194) );
CKINVDCx16_ASAP7_75t_R g114 ( .A(n_9), .Y(n_114) );
XNOR2xp5_ASAP7_75t_L g132 ( .A(n_10), .B(n_133), .Y(n_132) );
CKINVDCx5p33_ASAP7_75t_R g209 ( .A(n_11), .Y(n_209) );
NAND2xp33_ASAP7_75t_L g581 ( .A(n_12), .B(n_227), .Y(n_581) );
INVx2_ASAP7_75t_L g154 ( .A(n_13), .Y(n_154) );
AOI221x1_ASAP7_75t_L g530 ( .A1(n_14), .A2(n_26), .B1(n_520), .B2(n_523), .C(n_531), .Y(n_530) );
NOR3xp33_ASAP7_75t_L g112 ( .A(n_15), .B(n_113), .C(n_115), .Y(n_112) );
CKINVDCx16_ASAP7_75t_R g126 ( .A(n_15), .Y(n_126) );
NAND2xp5_ASAP7_75t_SL g577 ( .A(n_16), .B(n_520), .Y(n_577) );
INVx1_ASAP7_75t_L g228 ( .A(n_17), .Y(n_228) );
AO21x2_ASAP7_75t_L g575 ( .A1(n_18), .A2(n_191), .B(n_576), .Y(n_575) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_19), .B(n_185), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g570 ( .A(n_20), .B(n_230), .Y(n_570) );
AO21x1_ASAP7_75t_L g519 ( .A1(n_21), .A2(n_520), .B(n_521), .Y(n_519) );
INVx1_ASAP7_75t_L g110 ( .A(n_22), .Y(n_110) );
INVx1_ASAP7_75t_L g225 ( .A(n_23), .Y(n_225) );
INVx1_ASAP7_75t_SL g279 ( .A(n_24), .Y(n_279) );
NAND2xp5_ASAP7_75t_SL g241 ( .A(n_25), .B(n_177), .Y(n_241) );
AOI33xp33_ASAP7_75t_L g265 ( .A1(n_27), .A2(n_56), .A3(n_159), .B1(n_170), .B2(n_266), .B3(n_267), .Y(n_265) );
NAND2x1_ASAP7_75t_L g541 ( .A(n_28), .B(n_230), .Y(n_541) );
AOI22xp5_ASAP7_75t_SL g823 ( .A1(n_29), .A2(n_824), .B1(n_827), .B2(n_828), .Y(n_823) );
CKINVDCx20_ASAP7_75t_R g828 ( .A(n_29), .Y(n_828) );
NAND2x1_ASAP7_75t_L g595 ( .A(n_30), .B(n_227), .Y(n_595) );
INVx1_ASAP7_75t_L g202 ( .A(n_31), .Y(n_202) );
OA21x2_ASAP7_75t_L g153 ( .A1(n_32), .A2(n_89), .B(n_154), .Y(n_153) );
OR2x2_ASAP7_75t_L g187 ( .A(n_32), .B(n_89), .Y(n_187) );
NAND2xp5_ASAP7_75t_L g276 ( .A(n_33), .B(n_157), .Y(n_276) );
NAND2xp5_ASAP7_75t_L g590 ( .A(n_34), .B(n_227), .Y(n_590) );
NAND2xp5_ASAP7_75t_L g580 ( .A(n_35), .B(n_230), .Y(n_580) );
AOI22xp5_ASAP7_75t_L g824 ( .A1(n_36), .A2(n_67), .B1(n_825), .B2(n_826), .Y(n_824) );
CKINVDCx20_ASAP7_75t_R g826 ( .A(n_36), .Y(n_826) );
NAND2xp5_ASAP7_75t_L g525 ( .A(n_37), .B(n_227), .Y(n_525) );
AOI21xp5_ASAP7_75t_L g549 ( .A1(n_38), .A2(n_523), .B(n_550), .Y(n_549) );
AND2x2_ASAP7_75t_L g164 ( .A(n_39), .B(n_165), .Y(n_164) );
INVx1_ASAP7_75t_L g169 ( .A(n_39), .Y(n_169) );
AND2x2_ASAP7_75t_L g183 ( .A(n_39), .B(n_162), .Y(n_183) );
INVxp67_ASAP7_75t_L g115 ( .A(n_40), .Y(n_115) );
OR2x6_ASAP7_75t_L g128 ( .A(n_40), .B(n_109), .Y(n_128) );
CKINVDCx20_ASAP7_75t_R g205 ( .A(n_41), .Y(n_205) );
NAND2xp5_ASAP7_75t_SL g553 ( .A(n_42), .B(n_520), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g156 ( .A(n_43), .B(n_157), .Y(n_156) );
AOI22xp5_ASAP7_75t_L g234 ( .A1(n_44), .A2(n_152), .B1(n_219), .B2(n_235), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g242 ( .A(n_45), .B(n_243), .Y(n_242) );
NAND2xp5_ASAP7_75t_L g280 ( .A(n_46), .B(n_177), .Y(n_280) );
AOI22xp5_ASAP7_75t_L g133 ( .A1(n_47), .A2(n_98), .B1(n_134), .B2(n_135), .Y(n_133) );
CKINVDCx20_ASAP7_75t_R g135 ( .A(n_47), .Y(n_135) );
CKINVDCx20_ASAP7_75t_R g574 ( .A(n_48), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g551 ( .A(n_49), .B(n_227), .Y(n_551) );
NAND2xp5_ASAP7_75t_SL g196 ( .A(n_50), .B(n_191), .Y(n_196) );
NAND2xp5_ASAP7_75t_L g195 ( .A(n_51), .B(n_177), .Y(n_195) );
AOI21xp5_ASAP7_75t_L g593 ( .A1(n_52), .A2(n_523), .B(n_594), .Y(n_593) );
CKINVDCx5p33_ASAP7_75t_R g238 ( .A(n_53), .Y(n_238) );
CKINVDCx20_ASAP7_75t_R g833 ( .A(n_54), .Y(n_833) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_55), .B(n_227), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g176 ( .A(n_57), .B(n_177), .Y(n_176) );
INVx1_ASAP7_75t_L g160 ( .A(n_58), .Y(n_160) );
INVx1_ASAP7_75t_L g179 ( .A(n_58), .Y(n_179) );
AND2x2_ASAP7_75t_L g184 ( .A(n_59), .B(n_185), .Y(n_184) );
AOI221xp5_ASAP7_75t_L g192 ( .A1(n_60), .A2(n_78), .B1(n_157), .B2(n_167), .C(n_193), .Y(n_192) );
NAND2xp5_ASAP7_75t_L g253 ( .A(n_61), .B(n_157), .Y(n_253) );
NAND2xp5_ASAP7_75t_L g122 ( .A(n_62), .B(n_123), .Y(n_122) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_63), .B(n_230), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g211 ( .A(n_64), .B(n_152), .Y(n_211) );
AOI21xp5_ASAP7_75t_SL g249 ( .A1(n_65), .A2(n_167), .B(n_250), .Y(n_249) );
AOI21xp5_ASAP7_75t_L g539 ( .A1(n_66), .A2(n_523), .B(n_540), .Y(n_539) );
CKINVDCx20_ASAP7_75t_R g825 ( .A(n_67), .Y(n_825) );
INVx1_ASAP7_75t_L g222 ( .A(n_68), .Y(n_222) );
AO21x1_ASAP7_75t_L g522 ( .A1(n_69), .A2(n_523), .B(n_524), .Y(n_522) );
NAND2xp5_ASAP7_75t_SL g586 ( .A(n_70), .B(n_520), .Y(n_586) );
INVx1_ASAP7_75t_L g174 ( .A(n_71), .Y(n_174) );
NAND2xp5_ASAP7_75t_SL g597 ( .A(n_72), .B(n_520), .Y(n_597) );
AOI21xp5_ASAP7_75t_L g166 ( .A1(n_73), .A2(n_167), .B(n_173), .Y(n_166) );
AND2x2_ASAP7_75t_L g554 ( .A(n_74), .B(n_186), .Y(n_554) );
INVx1_ASAP7_75t_L g165 ( .A(n_75), .Y(n_165) );
INVx1_ASAP7_75t_L g181 ( .A(n_75), .Y(n_181) );
AND2x2_ASAP7_75t_L g598 ( .A(n_76), .B(n_151), .Y(n_598) );
NAND2xp5_ASAP7_75t_L g268 ( .A(n_77), .B(n_157), .Y(n_268) );
AND2x2_ASAP7_75t_L g281 ( .A(n_79), .B(n_151), .Y(n_281) );
CKINVDCx20_ASAP7_75t_R g829 ( .A(n_79), .Y(n_829) );
INVx1_ASAP7_75t_L g223 ( .A(n_80), .Y(n_223) );
AOI21xp5_ASAP7_75t_L g277 ( .A1(n_81), .A2(n_167), .B(n_278), .Y(n_277) );
A2O1A1Ixp33_ASAP7_75t_L g239 ( .A1(n_82), .A2(n_167), .B(n_240), .C(n_244), .Y(n_239) );
INVx1_ASAP7_75t_L g111 ( .A(n_83), .Y(n_111) );
NAND2xp5_ASAP7_75t_SL g572 ( .A(n_84), .B(n_520), .Y(n_572) );
AND2x2_ASAP7_75t_SL g247 ( .A(n_85), .B(n_151), .Y(n_247) );
AND2x2_ASAP7_75t_L g584 ( .A(n_86), .B(n_151), .Y(n_584) );
AOI22xp5_ASAP7_75t_L g262 ( .A1(n_87), .A2(n_167), .B1(n_263), .B2(n_264), .Y(n_262) );
AND2x2_ASAP7_75t_L g521 ( .A(n_88), .B(n_219), .Y(n_521) );
AND2x2_ASAP7_75t_L g544 ( .A(n_90), .B(n_151), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g571 ( .A(n_91), .B(n_227), .Y(n_571) );
INVx1_ASAP7_75t_L g251 ( .A(n_92), .Y(n_251) );
CKINVDCx20_ASAP7_75t_R g811 ( .A(n_93), .Y(n_811) );
NAND2xp5_ASAP7_75t_L g552 ( .A(n_94), .B(n_230), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_95), .B(n_227), .Y(n_532) );
AOI21xp5_ASAP7_75t_L g568 ( .A1(n_96), .A2(n_523), .B(n_569), .Y(n_568) );
AND2x2_ASAP7_75t_L g269 ( .A(n_97), .B(n_151), .Y(n_269) );
CKINVDCx20_ASAP7_75t_R g134 ( .A(n_98), .Y(n_134) );
NAND2xp5_ASAP7_75t_L g589 ( .A(n_99), .B(n_230), .Y(n_589) );
A2O1A1Ixp33_ASAP7_75t_L g199 ( .A1(n_100), .A2(n_200), .B(n_201), .C(n_204), .Y(n_199) );
BUFx2_ASAP7_75t_L g121 ( .A(n_101), .Y(n_121) );
AOI21xp5_ASAP7_75t_L g578 ( .A1(n_102), .A2(n_523), .B(n_579), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g252 ( .A(n_103), .B(n_177), .Y(n_252) );
AOI21xp33_ASAP7_75t_SL g104 ( .A1(n_105), .A2(n_116), .B(n_832), .Y(n_104) );
CKINVDCx5p33_ASAP7_75t_R g105 ( .A(n_106), .Y(n_105) );
CKINVDCx20_ASAP7_75t_R g834 ( .A(n_106), .Y(n_834) );
INVx2_ASAP7_75t_SL g106 ( .A(n_107), .Y(n_106) );
AND2x2_ASAP7_75t_SL g107 ( .A(n_108), .B(n_112), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
NAND2xp5_ASAP7_75t_L g109 ( .A(n_110), .B(n_111), .Y(n_109) );
OA22x2_ASAP7_75t_L g116 ( .A1(n_117), .A2(n_129), .B1(n_814), .B2(n_816), .Y(n_116) );
NAND2xp5_ASAP7_75t_L g117 ( .A(n_118), .B(n_122), .Y(n_117) );
CKINVDCx11_ASAP7_75t_R g118 ( .A(n_119), .Y(n_118) );
CKINVDCx20_ASAP7_75t_R g119 ( .A(n_120), .Y(n_119) );
HB1xp67_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
CKINVDCx20_ASAP7_75t_R g815 ( .A(n_121), .Y(n_815) );
CKINVDCx20_ASAP7_75t_R g830 ( .A(n_122), .Y(n_830) );
INVx1_ASAP7_75t_SL g123 ( .A(n_124), .Y(n_123) );
BUFx2_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
BUFx3_ASAP7_75t_L g821 ( .A(n_125), .Y(n_821) );
NAND2xp5_ASAP7_75t_L g125 ( .A(n_126), .B(n_127), .Y(n_125) );
CKINVDCx16_ASAP7_75t_R g138 ( .A(n_126), .Y(n_138) );
OR2x2_ASAP7_75t_L g813 ( .A(n_126), .B(n_128), .Y(n_813) );
OAI22xp5_ASAP7_75t_SL g129 ( .A1(n_127), .A2(n_130), .B1(n_811), .B2(n_812), .Y(n_129) );
CKINVDCx5p33_ASAP7_75t_R g127 ( .A(n_128), .Y(n_127) );
XNOR2xp5_ASAP7_75t_L g130 ( .A(n_131), .B(n_136), .Y(n_130) );
OAI22xp5_ASAP7_75t_L g136 ( .A1(n_137), .A2(n_138), .B1(n_139), .B2(n_511), .Y(n_136) );
CKINVDCx5p33_ASAP7_75t_R g137 ( .A(n_138), .Y(n_137) );
INVx2_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
NAND4xp75_ASAP7_75t_L g140 ( .A(n_141), .B(n_383), .C(n_428), .D(n_497), .Y(n_140) );
INVx1_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
NAND2x1_ASAP7_75t_L g142 ( .A(n_143), .B(n_343), .Y(n_142) );
NOR3xp33_ASAP7_75t_L g143 ( .A(n_144), .B(n_299), .C(n_324), .Y(n_143) );
OAI222xp33_ASAP7_75t_L g144 ( .A1(n_145), .A2(n_213), .B1(n_254), .B2(n_270), .C1(n_286), .C2(n_293), .Y(n_144) );
INVxp67_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
AND2x2_ASAP7_75t_L g146 ( .A(n_147), .B(n_188), .Y(n_146) );
AND2x2_ASAP7_75t_L g508 ( .A(n_147), .B(n_322), .Y(n_508) );
INVx1_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
HB1xp67_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
NAND2xp5_ASAP7_75t_L g259 ( .A(n_149), .B(n_260), .Y(n_259) );
NAND2xp5_ASAP7_75t_L g298 ( .A(n_149), .B(n_197), .Y(n_298) );
INVx3_ASAP7_75t_L g313 ( .A(n_149), .Y(n_313) );
AND2x2_ASAP7_75t_L g446 ( .A(n_149), .B(n_447), .Y(n_446) );
AO21x2_ASAP7_75t_L g149 ( .A1(n_150), .A2(n_155), .B(n_184), .Y(n_149) );
OAI22xp5_ASAP7_75t_L g198 ( .A1(n_150), .A2(n_151), .B1(n_199), .B2(n_205), .Y(n_198) );
AO21x2_ASAP7_75t_L g331 ( .A1(n_150), .A2(n_155), .B(n_184), .Y(n_331) );
AO21x2_ASAP7_75t_L g537 ( .A1(n_150), .A2(n_538), .B(n_544), .Y(n_537) );
AO21x2_ASAP7_75t_L g547 ( .A1(n_150), .A2(n_548), .B(n_554), .Y(n_547) );
AO21x2_ASAP7_75t_L g559 ( .A1(n_150), .A2(n_538), .B(n_544), .Y(n_559) );
AO21x2_ASAP7_75t_L g561 ( .A1(n_150), .A2(n_548), .B(n_554), .Y(n_561) );
INVx3_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
INVx4_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
NAND2xp5_ASAP7_75t_L g207 ( .A(n_152), .B(n_208), .Y(n_207) );
INVx3_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
BUFx4f_ASAP7_75t_L g191 ( .A(n_153), .Y(n_191) );
AND2x2_ASAP7_75t_SL g186 ( .A(n_154), .B(n_187), .Y(n_186) );
AND2x4_ASAP7_75t_L g219 ( .A(n_154), .B(n_187), .Y(n_219) );
NAND2xp5_ASAP7_75t_L g155 ( .A(n_156), .B(n_166), .Y(n_155) );
INVx1_ASAP7_75t_L g212 ( .A(n_157), .Y(n_212) );
AND2x4_ASAP7_75t_L g157 ( .A(n_158), .B(n_163), .Y(n_157) );
INVx1_ASAP7_75t_L g236 ( .A(n_158), .Y(n_236) );
AND2x2_ASAP7_75t_L g158 ( .A(n_159), .B(n_161), .Y(n_158) );
OR2x6_ASAP7_75t_L g175 ( .A(n_159), .B(n_171), .Y(n_175) );
INVxp33_ASAP7_75t_L g266 ( .A(n_159), .Y(n_266) );
INVx2_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
AND2x2_ASAP7_75t_L g172 ( .A(n_160), .B(n_162), .Y(n_172) );
AND2x4_ASAP7_75t_L g230 ( .A(n_160), .B(n_180), .Y(n_230) );
HB1xp67_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
INVx1_ASAP7_75t_L g237 ( .A(n_163), .Y(n_237) );
BUFx3_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
AND2x6_ASAP7_75t_L g523 ( .A(n_164), .B(n_172), .Y(n_523) );
INVx2_ASAP7_75t_L g171 ( .A(n_165), .Y(n_171) );
AND2x6_ASAP7_75t_L g227 ( .A(n_165), .B(n_178), .Y(n_227) );
INVxp67_ASAP7_75t_L g210 ( .A(n_167), .Y(n_210) );
AND2x4_ASAP7_75t_L g167 ( .A(n_168), .B(n_172), .Y(n_167) );
NOR2x1p5_ASAP7_75t_L g168 ( .A(n_169), .B(n_170), .Y(n_168) );
INVx1_ASAP7_75t_L g267 ( .A(n_170), .Y(n_267) );
INVx3_ASAP7_75t_L g170 ( .A(n_171), .Y(n_170) );
O2A1O1Ixp33_ASAP7_75t_L g173 ( .A1(n_174), .A2(n_175), .B(n_176), .C(n_182), .Y(n_173) );
O2A1O1Ixp33_ASAP7_75t_SL g193 ( .A1(n_175), .A2(n_182), .B(n_194), .C(n_195), .Y(n_193) );
INVxp67_ASAP7_75t_L g200 ( .A(n_175), .Y(n_200) );
OAI22xp5_ASAP7_75t_L g221 ( .A1(n_175), .A2(n_203), .B1(n_222), .B2(n_223), .Y(n_221) );
INVx2_ASAP7_75t_L g243 ( .A(n_175), .Y(n_243) );
O2A1O1Ixp33_ASAP7_75t_L g250 ( .A1(n_175), .A2(n_182), .B(n_251), .C(n_252), .Y(n_250) );
O2A1O1Ixp33_ASAP7_75t_SL g278 ( .A1(n_175), .A2(n_182), .B(n_279), .C(n_280), .Y(n_278) );
INVx1_ASAP7_75t_L g203 ( .A(n_177), .Y(n_203) );
AND2x4_ASAP7_75t_L g520 ( .A(n_177), .B(n_183), .Y(n_520) );
AND2x4_ASAP7_75t_L g177 ( .A(n_178), .B(n_180), .Y(n_177) );
INVx2_ASAP7_75t_L g178 ( .A(n_179), .Y(n_178) );
INVx2_ASAP7_75t_L g180 ( .A(n_181), .Y(n_180) );
NOR2xp33_ASAP7_75t_L g231 ( .A(n_182), .B(n_219), .Y(n_231) );
AOI21xp5_ASAP7_75t_L g240 ( .A1(n_182), .A2(n_241), .B(n_242), .Y(n_240) );
INVx1_ASAP7_75t_L g263 ( .A(n_182), .Y(n_263) );
AOI21xp5_ASAP7_75t_L g524 ( .A1(n_182), .A2(n_525), .B(n_526), .Y(n_524) );
AOI21xp5_ASAP7_75t_L g531 ( .A1(n_182), .A2(n_532), .B(n_533), .Y(n_531) );
AOI21xp5_ASAP7_75t_L g540 ( .A1(n_182), .A2(n_541), .B(n_542), .Y(n_540) );
AOI21xp5_ASAP7_75t_L g550 ( .A1(n_182), .A2(n_551), .B(n_552), .Y(n_550) );
AOI21xp5_ASAP7_75t_L g569 ( .A1(n_182), .A2(n_570), .B(n_571), .Y(n_569) );
AOI21xp5_ASAP7_75t_L g579 ( .A1(n_182), .A2(n_580), .B(n_581), .Y(n_579) );
AOI21xp5_ASAP7_75t_L g588 ( .A1(n_182), .A2(n_589), .B(n_590), .Y(n_588) );
AOI21xp5_ASAP7_75t_L g594 ( .A1(n_182), .A2(n_595), .B(n_596), .Y(n_594) );
INVx5_ASAP7_75t_L g182 ( .A(n_183), .Y(n_182) );
HB1xp67_ASAP7_75t_L g204 ( .A(n_183), .Y(n_204) );
CKINVDCx5p33_ASAP7_75t_R g274 ( .A(n_185), .Y(n_274) );
OA21x2_ASAP7_75t_L g529 ( .A1(n_185), .A2(n_530), .B(n_534), .Y(n_529) );
OA21x2_ASAP7_75t_L g557 ( .A1(n_185), .A2(n_530), .B(n_534), .Y(n_557) );
AOI21xp5_ASAP7_75t_L g585 ( .A1(n_185), .A2(n_586), .B(n_587), .Y(n_585) );
BUFx6f_ASAP7_75t_L g185 ( .A(n_186), .Y(n_185) );
AND2x2_ASAP7_75t_L g376 ( .A(n_188), .B(n_329), .Y(n_376) );
AND2x2_ASAP7_75t_L g378 ( .A(n_188), .B(n_379), .Y(n_378) );
INVx3_ASAP7_75t_L g413 ( .A(n_188), .Y(n_413) );
AND2x4_ASAP7_75t_L g188 ( .A(n_189), .B(n_197), .Y(n_188) );
INVx2_ASAP7_75t_L g189 ( .A(n_190), .Y(n_189) );
INVxp67_ASAP7_75t_L g296 ( .A(n_190), .Y(n_296) );
INVx1_ASAP7_75t_L g315 ( .A(n_190), .Y(n_315) );
AND2x4_ASAP7_75t_L g322 ( .A(n_190), .B(n_323), .Y(n_322) );
NAND2xp5_ASAP7_75t_L g338 ( .A(n_190), .B(n_260), .Y(n_338) );
HB1xp67_ASAP7_75t_L g447 ( .A(n_190), .Y(n_447) );
INVx1_ASAP7_75t_L g457 ( .A(n_190), .Y(n_457) );
OA21x2_ASAP7_75t_L g190 ( .A1(n_191), .A2(n_192), .B(n_196), .Y(n_190) );
INVx2_ASAP7_75t_SL g244 ( .A(n_191), .Y(n_244) );
INVx1_ASAP7_75t_L g257 ( .A(n_197), .Y(n_257) );
INVx2_ASAP7_75t_L g310 ( .A(n_197), .Y(n_310) );
INVx1_ASAP7_75t_L g391 ( .A(n_197), .Y(n_391) );
OR2x2_ASAP7_75t_L g197 ( .A(n_198), .B(n_206), .Y(n_197) );
NOR2xp33_ASAP7_75t_L g201 ( .A(n_202), .B(n_203), .Y(n_201) );
OAI22xp5_ASAP7_75t_L g206 ( .A1(n_207), .A2(n_210), .B1(n_211), .B2(n_212), .Y(n_206) );
INVx1_ASAP7_75t_L g208 ( .A(n_209), .Y(n_208) );
INVx1_ASAP7_75t_L g213 ( .A(n_214), .Y(n_213) );
AND2x2_ASAP7_75t_SL g214 ( .A(n_215), .B(n_245), .Y(n_214) );
NAND2xp5_ASAP7_75t_L g366 ( .A(n_215), .B(n_272), .Y(n_366) );
INVx2_ASAP7_75t_L g387 ( .A(n_215), .Y(n_387) );
AND2x2_ASAP7_75t_L g395 ( .A(n_215), .B(n_396), .Y(n_395) );
AND2x2_ASAP7_75t_L g215 ( .A(n_216), .B(n_232), .Y(n_215) );
AND2x4_ASAP7_75t_L g285 ( .A(n_216), .B(n_233), .Y(n_285) );
INVx1_ASAP7_75t_L g292 ( .A(n_216), .Y(n_292) );
AND2x2_ASAP7_75t_L g468 ( .A(n_216), .B(n_273), .Y(n_468) );
INVx3_ASAP7_75t_L g216 ( .A(n_217), .Y(n_216) );
AND2x2_ASAP7_75t_L g306 ( .A(n_217), .B(n_233), .Y(n_306) );
INVx2_ASAP7_75t_L g342 ( .A(n_217), .Y(n_342) );
AND2x2_ASAP7_75t_L g421 ( .A(n_217), .B(n_273), .Y(n_421) );
NOR2x1_ASAP7_75t_SL g464 ( .A(n_217), .B(n_246), .Y(n_464) );
AND2x4_ASAP7_75t_L g217 ( .A(n_218), .B(n_220), .Y(n_217) );
AOI21xp5_ASAP7_75t_L g248 ( .A1(n_219), .A2(n_249), .B(n_253), .Y(n_248) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_219), .B(n_528), .Y(n_527) );
INVx1_ASAP7_75t_SL g566 ( .A(n_219), .Y(n_566) );
AOI21xp5_ASAP7_75t_L g576 ( .A1(n_219), .A2(n_577), .B(n_578), .Y(n_576) );
OAI21xp5_ASAP7_75t_L g220 ( .A1(n_221), .A2(n_224), .B(n_231), .Y(n_220) );
OAI22xp5_ASAP7_75t_L g224 ( .A1(n_225), .A2(n_226), .B1(n_228), .B2(n_229), .Y(n_224) );
INVxp67_ASAP7_75t_L g226 ( .A(n_227), .Y(n_226) );
INVxp67_ASAP7_75t_L g229 ( .A(n_230), .Y(n_229) );
INVx1_ASAP7_75t_L g304 ( .A(n_232), .Y(n_304) );
INVx2_ASAP7_75t_L g232 ( .A(n_233), .Y(n_232) );
AND2x2_ASAP7_75t_L g318 ( .A(n_233), .B(n_246), .Y(n_318) );
INVx1_ASAP7_75t_L g334 ( .A(n_233), .Y(n_334) );
HB1xp67_ASAP7_75t_L g442 ( .A(n_233), .Y(n_442) );
AND2x2_ASAP7_75t_L g233 ( .A(n_234), .B(n_239), .Y(n_233) );
NOR3xp33_ASAP7_75t_L g235 ( .A(n_236), .B(n_237), .C(n_238), .Y(n_235) );
AO21x2_ASAP7_75t_L g260 ( .A1(n_244), .A2(n_261), .B(n_269), .Y(n_260) );
AO21x2_ASAP7_75t_L g311 ( .A1(n_244), .A2(n_261), .B(n_269), .Y(n_311) );
AND2x2_ASAP7_75t_L g305 ( .A(n_245), .B(n_306), .Y(n_305) );
OR2x6_ASAP7_75t_L g386 ( .A(n_245), .B(n_387), .Y(n_386) );
AND2x2_ASAP7_75t_L g424 ( .A(n_245), .B(n_421), .Y(n_424) );
BUFx6f_ASAP7_75t_L g245 ( .A(n_246), .Y(n_245) );
INVx4_ASAP7_75t_L g283 ( .A(n_246), .Y(n_283) );
NAND2xp5_ASAP7_75t_SL g291 ( .A(n_246), .B(n_292), .Y(n_291) );
INVx2_ASAP7_75t_L g353 ( .A(n_246), .Y(n_353) );
OR2x2_ASAP7_75t_L g359 ( .A(n_246), .B(n_273), .Y(n_359) );
AND2x4_ASAP7_75t_L g373 ( .A(n_246), .B(n_334), .Y(n_373) );
AND2x2_ASAP7_75t_L g374 ( .A(n_246), .B(n_342), .Y(n_374) );
OR2x6_ASAP7_75t_L g246 ( .A(n_247), .B(n_248), .Y(n_246) );
INVx1_ASAP7_75t_L g254 ( .A(n_255), .Y(n_254) );
AND2x2_ASAP7_75t_L g255 ( .A(n_256), .B(n_258), .Y(n_255) );
INVx1_ASAP7_75t_SL g256 ( .A(n_257), .Y(n_256) );
AND2x2_ASAP7_75t_L g418 ( .A(n_257), .B(n_337), .Y(n_418) );
BUFx2_ASAP7_75t_L g470 ( .A(n_257), .Y(n_470) );
INVx1_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
OR2x2_ASAP7_75t_L g501 ( .A(n_259), .B(n_413), .Y(n_501) );
INVx2_ASAP7_75t_L g295 ( .A(n_260), .Y(n_295) );
NAND2xp5_ASAP7_75t_SL g261 ( .A(n_262), .B(n_268), .Y(n_261) );
INVx1_ASAP7_75t_L g264 ( .A(n_265), .Y(n_264) );
NAND2xp5_ASAP7_75t_L g270 ( .A(n_271), .B(n_282), .Y(n_270) );
AND2x2_ASAP7_75t_L g317 ( .A(n_271), .B(n_318), .Y(n_317) );
HB1xp67_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
AND2x4_ASAP7_75t_SL g302 ( .A(n_272), .B(n_292), .Y(n_302) );
INVx1_ASAP7_75t_L g272 ( .A(n_273), .Y(n_272) );
INVx2_ASAP7_75t_L g290 ( .A(n_273), .Y(n_290) );
HB1xp67_ASAP7_75t_L g396 ( .A(n_273), .Y(n_396) );
HB1xp67_ASAP7_75t_L g463 ( .A(n_273), .Y(n_463) );
INVx1_ASAP7_75t_L g503 ( .A(n_273), .Y(n_503) );
AO21x2_ASAP7_75t_L g273 ( .A1(n_274), .A2(n_275), .B(n_281), .Y(n_273) );
AO21x2_ASAP7_75t_L g591 ( .A1(n_274), .A2(n_592), .B(n_598), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g275 ( .A(n_276), .B(n_277), .Y(n_275) );
BUFx2_ASAP7_75t_L g417 ( .A(n_282), .Y(n_417) );
NOR2x1_ASAP7_75t_L g282 ( .A(n_283), .B(n_284), .Y(n_282) );
AND2x4_ASAP7_75t_L g333 ( .A(n_283), .B(n_334), .Y(n_333) );
NOR2xp67_ASAP7_75t_SL g365 ( .A(n_283), .B(n_366), .Y(n_365) );
AND2x2_ASAP7_75t_L g438 ( .A(n_283), .B(n_421), .Y(n_438) );
AND2x4_ASAP7_75t_SL g441 ( .A(n_283), .B(n_442), .Y(n_441) );
OR2x2_ASAP7_75t_L g490 ( .A(n_283), .B(n_491), .Y(n_490) );
INVx2_ASAP7_75t_L g357 ( .A(n_284), .Y(n_357) );
INVx4_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
AND2x2_ASAP7_75t_L g352 ( .A(n_285), .B(n_353), .Y(n_352) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_285), .B(n_350), .Y(n_370) );
NAND2xp5_ASAP7_75t_L g409 ( .A(n_285), .B(n_410), .Y(n_409) );
NOR2xp33_ASAP7_75t_L g473 ( .A(n_285), .B(n_474), .Y(n_473) );
INVx1_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
NOR2x1_ASAP7_75t_L g287 ( .A(n_288), .B(n_291), .Y(n_287) );
INVx1_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
OR2x2_ASAP7_75t_L g435 ( .A(n_289), .B(n_436), .Y(n_435) );
HB1xp67_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
INVx2_ASAP7_75t_L g351 ( .A(n_290), .Y(n_351) );
NAND2x1p5_ASAP7_75t_L g293 ( .A(n_294), .B(n_297), .Y(n_293) );
AND2x2_ASAP7_75t_L g469 ( .A(n_294), .B(n_470), .Y(n_469) );
AND2x2_ASAP7_75t_L g477 ( .A(n_294), .B(n_406), .Y(n_477) );
AND2x2_ASAP7_75t_L g294 ( .A(n_295), .B(n_296), .Y(n_294) );
AND2x2_ASAP7_75t_L g346 ( .A(n_295), .B(n_331), .Y(n_346) );
AND2x4_ASAP7_75t_L g379 ( .A(n_295), .B(n_313), .Y(n_379) );
INVx1_ASAP7_75t_L g496 ( .A(n_295), .Y(n_496) );
AND2x2_ASAP7_75t_L g382 ( .A(n_297), .B(n_322), .Y(n_382) );
INVx2_ASAP7_75t_SL g297 ( .A(n_298), .Y(n_297) );
OR2x2_ASAP7_75t_L g403 ( .A(n_298), .B(n_338), .Y(n_403) );
OAI22xp5_ASAP7_75t_L g299 ( .A1(n_300), .A2(n_307), .B1(n_316), .B2(n_319), .Y(n_299) );
AOI21xp5_ASAP7_75t_L g300 ( .A1(n_301), .A2(n_303), .B(n_305), .Y(n_300) );
OAI22xp5_ASAP7_75t_SL g482 ( .A1(n_301), .A2(n_370), .B1(n_478), .B2(n_483), .Y(n_482) );
INVx1_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
NAND2xp5_ASAP7_75t_L g332 ( .A(n_302), .B(n_333), .Y(n_332) );
AND2x4_ASAP7_75t_L g371 ( .A(n_302), .B(n_303), .Y(n_371) );
AND2x2_ASAP7_75t_SL g401 ( .A(n_302), .B(n_373), .Y(n_401) );
AOI211xp5_ASAP7_75t_SL g489 ( .A1(n_302), .A2(n_490), .B(n_492), .C(n_493), .Y(n_489) );
AND2x2_ASAP7_75t_SL g420 ( .A(n_303), .B(n_421), .Y(n_420) );
NAND2xp5_ASAP7_75t_L g475 ( .A(n_303), .B(n_349), .Y(n_475) );
INVx2_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
INVx1_ASAP7_75t_L g380 ( .A(n_305), .Y(n_380) );
INVx2_ASAP7_75t_L g436 ( .A(n_306), .Y(n_436) );
AND2x2_ASAP7_75t_L g510 ( .A(n_306), .B(n_503), .Y(n_510) );
OAI21xp5_ASAP7_75t_L g458 ( .A1(n_307), .A2(n_459), .B(n_465), .Y(n_458) );
OR2x2_ASAP7_75t_L g307 ( .A(n_308), .B(n_312), .Y(n_307) );
INVx1_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
AND2x4_ASAP7_75t_L g445 ( .A(n_309), .B(n_446), .Y(n_445) );
AND2x2_ASAP7_75t_L g455 ( .A(n_309), .B(n_456), .Y(n_455) );
AND2x2_ASAP7_75t_L g309 ( .A(n_310), .B(n_311), .Y(n_309) );
AND2x2_ASAP7_75t_L g362 ( .A(n_310), .B(n_315), .Y(n_362) );
NOR2xp67_ASAP7_75t_L g364 ( .A(n_310), .B(n_331), .Y(n_364) );
AND2x2_ASAP7_75t_L g406 ( .A(n_310), .B(n_331), .Y(n_406) );
INVx2_ASAP7_75t_L g323 ( .A(n_311), .Y(n_323) );
AND2x4_ASAP7_75t_L g329 ( .A(n_311), .B(n_330), .Y(n_329) );
NAND2x1p5_ASAP7_75t_L g312 ( .A(n_313), .B(n_314), .Y(n_312) );
INVx3_ASAP7_75t_L g321 ( .A(n_313), .Y(n_321) );
INVx3_ASAP7_75t_L g327 ( .A(n_314), .Y(n_327) );
BUFx3_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
INVx1_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
OAI21xp5_ASAP7_75t_L g504 ( .A1(n_318), .A2(n_424), .B(n_500), .Y(n_504) );
INVx1_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
AND2x2_ASAP7_75t_L g320 ( .A(n_321), .B(n_322), .Y(n_320) );
INVx1_ASAP7_75t_L g336 ( .A(n_321), .Y(n_336) );
NAND2xp5_ASAP7_75t_L g361 ( .A(n_321), .B(n_362), .Y(n_361) );
NAND2xp5_ASAP7_75t_L g411 ( .A(n_321), .B(n_396), .Y(n_411) );
OR2x2_ASAP7_75t_L g426 ( .A(n_321), .B(n_427), .Y(n_426) );
AND2x2_ASAP7_75t_L g433 ( .A(n_321), .B(n_337), .Y(n_433) );
AND2x2_ASAP7_75t_L g389 ( .A(n_322), .B(n_390), .Y(n_389) );
AND2x2_ASAP7_75t_L g405 ( .A(n_322), .B(n_406), .Y(n_405) );
AND2x2_ASAP7_75t_L g422 ( .A(n_322), .B(n_391), .Y(n_422) );
OAI22xp33_ASAP7_75t_L g324 ( .A1(n_325), .A2(n_332), .B1(n_335), .B2(n_339), .Y(n_324) );
NAND2xp5_ASAP7_75t_L g325 ( .A(n_326), .B(n_328), .Y(n_325) );
INVx1_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
NOR2xp67_ASAP7_75t_L g399 ( .A(n_327), .B(n_328), .Y(n_399) );
NOR2xp67_ASAP7_75t_SL g437 ( .A(n_327), .B(n_345), .Y(n_437) );
INVxp67_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
INVx2_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
NOR2x1_ASAP7_75t_L g456 ( .A(n_331), .B(n_457), .Y(n_456) );
AND2x2_ASAP7_75t_L g340 ( .A(n_333), .B(n_341), .Y(n_340) );
AND2x2_ASAP7_75t_L g404 ( .A(n_333), .B(n_350), .Y(n_404) );
NAND2xp5_ASAP7_75t_L g467 ( .A(n_333), .B(n_468), .Y(n_467) );
NAND2xp5_ASAP7_75t_L g335 ( .A(n_336), .B(n_337), .Y(n_335) );
INVx2_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
INVx1_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
AND2x2_ASAP7_75t_L g507 ( .A(n_341), .B(n_373), .Y(n_507) );
INVx1_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
NOR2x1_ASAP7_75t_L g452 ( .A(n_342), .B(n_453), .Y(n_452) );
NOR2xp67_ASAP7_75t_SL g343 ( .A(n_344), .B(n_367), .Y(n_343) );
OAI211xp5_ASAP7_75t_L g344 ( .A1(n_345), .A2(n_347), .B(n_354), .C(n_363), .Y(n_344) );
A2O1A1Ixp33_ASAP7_75t_L g407 ( .A1(n_345), .A2(n_398), .B(n_408), .C(n_412), .Y(n_407) );
INVx1_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
AND2x2_ASAP7_75t_L g487 ( .A(n_346), .B(n_488), .Y(n_487) );
INVx2_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
AND2x2_ASAP7_75t_L g348 ( .A(n_349), .B(n_352), .Y(n_348) );
INVx1_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
AND2x2_ASAP7_75t_L g398 ( .A(n_350), .B(n_374), .Y(n_398) );
AND2x2_ASAP7_75t_L g485 ( .A(n_350), .B(n_464), .Y(n_485) );
INVx3_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
INVx1_ASAP7_75t_L g453 ( .A(n_353), .Y(n_453) );
NAND2xp5_ASAP7_75t_L g354 ( .A(n_355), .B(n_360), .Y(n_354) );
INVx1_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
NAND2x1_ASAP7_75t_L g356 ( .A(n_357), .B(n_358), .Y(n_356) );
NAND2xp5_ASAP7_75t_L g381 ( .A(n_357), .B(n_382), .Y(n_381) );
INVx2_ASAP7_75t_SL g358 ( .A(n_359), .Y(n_358) );
INVx1_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
INVx2_ASAP7_75t_L g427 ( .A(n_362), .Y(n_427) );
NAND2xp33_ASAP7_75t_SL g363 ( .A(n_364), .B(n_365), .Y(n_363) );
OAI221xp5_ASAP7_75t_L g367 ( .A1(n_368), .A2(n_375), .B1(n_377), .B2(n_380), .C(n_381), .Y(n_367) );
NOR4xp25_ASAP7_75t_L g368 ( .A(n_369), .B(n_371), .C(n_372), .D(n_374), .Y(n_368) );
INVx1_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
HB1xp67_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
AND2x2_ASAP7_75t_L g486 ( .A(n_373), .B(n_449), .Y(n_486) );
INVx2_ASAP7_75t_L g492 ( .A(n_373), .Y(n_492) );
INVx2_ASAP7_75t_SL g375 ( .A(n_376), .Y(n_375) );
NAND2xp5_ASAP7_75t_L g439 ( .A(n_376), .B(n_440), .Y(n_439) );
INVx2_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
AND2x2_ASAP7_75t_L g479 ( .A(n_379), .B(n_480), .Y(n_479) );
INVx2_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
NAND4xp75_ASAP7_75t_L g384 ( .A(n_385), .B(n_407), .C(n_414), .D(n_423), .Y(n_384) );
OA211x2_ASAP7_75t_L g385 ( .A1(n_386), .A2(n_388), .B(n_392), .C(n_400), .Y(n_385) );
NAND2xp5_ASAP7_75t_L g434 ( .A(n_386), .B(n_435), .Y(n_434) );
INVx3_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
INVx1_ASAP7_75t_L g480 ( .A(n_390), .Y(n_480) );
INVx2_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
INVx1_ASAP7_75t_L g488 ( .A(n_391), .Y(n_488) );
NAND2xp5_ASAP7_75t_SL g392 ( .A(n_393), .B(n_399), .Y(n_392) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_394), .B(n_397), .Y(n_393) );
INVx2_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
BUFx2_ASAP7_75t_L g449 ( .A(n_396), .Y(n_449) );
INVx1_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
AOI22xp33_ASAP7_75t_L g400 ( .A1(n_401), .A2(n_402), .B1(n_404), .B2(n_405), .Y(n_400) );
INVx1_ASAP7_75t_SL g402 ( .A(n_403), .Y(n_402) );
OAI21xp5_ASAP7_75t_L g509 ( .A1(n_404), .A2(n_455), .B(n_510), .Y(n_509) );
INVx1_ASAP7_75t_SL g483 ( .A(n_405), .Y(n_483) );
NAND2x1p5_ASAP7_75t_L g495 ( .A(n_406), .B(n_496), .Y(n_495) );
INVxp67_ASAP7_75t_SL g408 ( .A(n_409), .Y(n_408) );
INVx1_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
INVx1_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
NOR2x1_ASAP7_75t_L g414 ( .A(n_415), .B(n_419), .Y(n_414) );
INVx1_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
NAND2xp5_ASAP7_75t_L g416 ( .A(n_417), .B(n_418), .Y(n_416) );
INVxp67_ASAP7_75t_L g481 ( .A(n_417), .Y(n_481) );
AND2x2_ASAP7_75t_L g419 ( .A(n_420), .B(n_422), .Y(n_419) );
AND2x2_ASAP7_75t_SL g440 ( .A(n_421), .B(n_441), .Y(n_440) );
AOI22xp5_ASAP7_75t_L g506 ( .A1(n_422), .A2(n_485), .B1(n_507), .B2(n_508), .Y(n_506) );
NAND2xp5_ASAP7_75t_L g423 ( .A(n_424), .B(n_425), .Y(n_423) );
INVx1_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
INVx2_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
NAND3x1_ASAP7_75t_L g429 ( .A(n_430), .B(n_471), .C(n_484), .Y(n_429) );
NOR3x1_ASAP7_75t_L g430 ( .A(n_431), .B(n_443), .C(n_458), .Y(n_430) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_432), .B(n_439), .Y(n_431) );
AOI22xp5_ASAP7_75t_L g432 ( .A1(n_433), .A2(n_434), .B1(n_437), .B2(n_438), .Y(n_432) );
OAI22xp5_ASAP7_75t_L g443 ( .A1(n_444), .A2(n_448), .B1(n_450), .B2(n_454), .Y(n_443) );
INVx1_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
INVx1_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
INVxp67_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
HB1xp67_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
AND2x2_ASAP7_75t_L g502 ( .A(n_452), .B(n_503), .Y(n_502) );
INVx1_ASAP7_75t_SL g454 ( .A(n_455), .Y(n_454) );
INVx1_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
AND2x2_ASAP7_75t_L g460 ( .A(n_461), .B(n_464), .Y(n_460) );
INVx1_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
INVx1_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
NAND2xp5_ASAP7_75t_L g465 ( .A(n_466), .B(n_469), .Y(n_465) );
INVxp67_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
INVx1_ASAP7_75t_SL g491 ( .A(n_468), .Y(n_491) );
OAI21xp5_ASAP7_75t_SL g499 ( .A1(n_469), .A2(n_500), .B(n_502), .Y(n_499) );
NOR2x1_ASAP7_75t_L g471 ( .A(n_472), .B(n_482), .Y(n_471) );
OAI22xp5_ASAP7_75t_L g472 ( .A1(n_473), .A2(n_476), .B1(n_478), .B2(n_481), .Y(n_472) );
INVxp67_ASAP7_75t_SL g474 ( .A(n_475), .Y(n_474) );
INVx1_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
INVx1_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
O2A1O1Ixp5_ASAP7_75t_L g484 ( .A1(n_485), .A2(n_486), .B(n_487), .C(n_489), .Y(n_484) );
INVx1_ASAP7_75t_L g493 ( .A(n_494), .Y(n_493) );
INVx1_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
NOR2x1_ASAP7_75t_SL g497 ( .A(n_498), .B(n_505), .Y(n_497) );
NAND2xp5_ASAP7_75t_L g498 ( .A(n_499), .B(n_504), .Y(n_498) );
INVx1_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
NAND2xp5_ASAP7_75t_SL g505 ( .A(n_506), .B(n_509), .Y(n_505) );
XOR2x1_ASAP7_75t_SL g822 ( .A(n_511), .B(n_823), .Y(n_822) );
AND2x4_ASAP7_75t_L g511 ( .A(n_512), .B(n_710), .Y(n_511) );
NOR3xp33_ASAP7_75t_L g512 ( .A(n_513), .B(n_647), .C(n_670), .Y(n_512) );
NAND3xp33_ASAP7_75t_SL g513 ( .A(n_514), .B(n_599), .C(n_616), .Y(n_513) );
OAI31xp33_ASAP7_75t_SL g514 ( .A1(n_515), .A2(n_535), .A3(n_555), .B(n_562), .Y(n_514) );
NAND2xp5_ASAP7_75t_L g673 ( .A(n_515), .B(n_674), .Y(n_673) );
INVx1_ASAP7_75t_SL g515 ( .A(n_516), .Y(n_515) );
OR2x2_ASAP7_75t_L g516 ( .A(n_517), .B(n_529), .Y(n_516) );
AND2x4_ASAP7_75t_L g602 ( .A(n_517), .B(n_529), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g631 ( .A(n_517), .B(n_546), .Y(n_631) );
AND2x4_ASAP7_75t_L g633 ( .A(n_517), .B(n_627), .Y(n_633) );
AND2x2_ASAP7_75t_L g764 ( .A(n_517), .B(n_559), .Y(n_764) );
INVx2_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
INVx2_ASAP7_75t_L g609 ( .A(n_518), .Y(n_609) );
OAI21x1_ASAP7_75t_SL g518 ( .A1(n_519), .A2(n_522), .B(n_527), .Y(n_518) );
INVx1_ASAP7_75t_L g528 ( .A(n_521), .Y(n_528) );
AND2x2_ASAP7_75t_L g545 ( .A(n_529), .B(n_546), .Y(n_545) );
AND2x2_ASAP7_75t_SL g700 ( .A(n_529), .B(n_608), .Y(n_700) );
AND2x2_ASAP7_75t_L g706 ( .A(n_529), .B(n_547), .Y(n_706) );
AND2x2_ASAP7_75t_L g795 ( .A(n_529), .B(n_796), .Y(n_795) );
INVx1_ASAP7_75t_SL g777 ( .A(n_535), .Y(n_777) );
AND2x2_ASAP7_75t_L g535 ( .A(n_536), .B(n_545), .Y(n_535) );
BUFx2_ASAP7_75t_L g606 ( .A(n_536), .Y(n_606) );
AND2x2_ASAP7_75t_L g640 ( .A(n_536), .B(n_546), .Y(n_640) );
AND2x2_ASAP7_75t_L g689 ( .A(n_536), .B(n_547), .Y(n_689) );
INVx2_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
AND2x2_ASAP7_75t_L g646 ( .A(n_537), .B(n_547), .Y(n_646) );
INVxp67_ASAP7_75t_L g658 ( .A(n_537), .Y(n_658) );
BUFx3_ASAP7_75t_L g703 ( .A(n_537), .Y(n_703) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_539), .B(n_543), .Y(n_538) );
OAI31xp33_ASAP7_75t_L g599 ( .A1(n_545), .A2(n_600), .A3(n_605), .B(n_610), .Y(n_599) );
AND2x2_ASAP7_75t_L g607 ( .A(n_546), .B(n_608), .Y(n_607) );
INVx2_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
AND2x2_ASAP7_75t_L g626 ( .A(n_547), .B(n_627), .Y(n_626) );
NAND2xp5_ASAP7_75t_SL g548 ( .A(n_549), .B(n_553), .Y(n_548) );
AOI322xp5_ASAP7_75t_L g800 ( .A1(n_555), .A2(n_675), .A3(n_704), .B1(n_709), .B2(n_801), .C1(n_804), .C2(n_805), .Y(n_800) );
AND2x2_ASAP7_75t_L g555 ( .A(n_556), .B(n_558), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g651 ( .A(n_556), .B(n_646), .Y(n_651) );
NAND2x1_ASAP7_75t_L g688 ( .A(n_556), .B(n_689), .Y(n_688) );
AND2x4_ASAP7_75t_L g732 ( .A(n_556), .B(n_636), .Y(n_732) );
INVx1_ASAP7_75t_SL g746 ( .A(n_556), .Y(n_746) );
INVx2_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
INVx2_ASAP7_75t_L g627 ( .A(n_557), .Y(n_627) );
HB1xp67_ASAP7_75t_L g770 ( .A(n_557), .Y(n_770) );
AND2x2_ASAP7_75t_L g699 ( .A(n_558), .B(n_700), .Y(n_699) );
NAND2xp5_ASAP7_75t_L g745 ( .A(n_558), .B(n_746), .Y(n_745) );
AND2x4_ASAP7_75t_SL g558 ( .A(n_559), .B(n_560), .Y(n_558) );
BUFx2_ASAP7_75t_L g604 ( .A(n_559), .Y(n_604) );
INVx1_ASAP7_75t_L g796 ( .A(n_559), .Y(n_796) );
OR2x2_ASAP7_75t_L g663 ( .A(n_560), .B(n_608), .Y(n_663) );
NAND2xp5_ASAP7_75t_SL g697 ( .A(n_560), .B(n_633), .Y(n_697) );
INVx2_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
AND2x4_ASAP7_75t_L g636 ( .A(n_561), .B(n_608), .Y(n_636) );
AND2x2_ASAP7_75t_L g562 ( .A(n_563), .B(n_582), .Y(n_562) );
INVxp67_ASAP7_75t_SL g563 ( .A(n_564), .Y(n_563) );
INVx1_ASAP7_75t_L g692 ( .A(n_564), .Y(n_692) );
OR2x2_ASAP7_75t_L g719 ( .A(n_564), .B(n_720), .Y(n_719) );
NAND2xp5_ASAP7_75t_L g564 ( .A(n_565), .B(n_575), .Y(n_564) );
NOR2x1_ASAP7_75t_SL g613 ( .A(n_565), .B(n_583), .Y(n_613) );
AND2x2_ASAP7_75t_L g620 ( .A(n_565), .B(n_621), .Y(n_620) );
AND2x2_ASAP7_75t_L g792 ( .A(n_565), .B(n_654), .Y(n_792) );
AO21x2_ASAP7_75t_L g565 ( .A1(n_566), .A2(n_567), .B(n_573), .Y(n_565) );
NOR2xp33_ASAP7_75t_L g573 ( .A(n_566), .B(n_574), .Y(n_573) );
AO21x2_ASAP7_75t_L g669 ( .A1(n_566), .A2(n_567), .B(n_573), .Y(n_669) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_568), .B(n_572), .Y(n_567) );
OR2x2_ASAP7_75t_L g614 ( .A(n_575), .B(n_615), .Y(n_614) );
BUFx3_ASAP7_75t_L g623 ( .A(n_575), .Y(n_623) );
INVx2_ASAP7_75t_L g654 ( .A(n_575), .Y(n_654) );
INVx1_ASAP7_75t_L g695 ( .A(n_575), .Y(n_695) );
AND2x2_ASAP7_75t_L g726 ( .A(n_575), .B(n_583), .Y(n_726) );
AND2x2_ASAP7_75t_L g757 ( .A(n_575), .B(n_684), .Y(n_757) );
AND2x2_ASAP7_75t_L g653 ( .A(n_582), .B(n_654), .Y(n_653) );
NAND2xp5_ASAP7_75t_L g665 ( .A(n_582), .B(n_666), .Y(n_665) );
AND2x2_ASAP7_75t_SL g756 ( .A(n_582), .B(n_757), .Y(n_756) );
AND2x2_ASAP7_75t_L g761 ( .A(n_582), .B(n_623), .Y(n_761) );
AND2x2_ASAP7_75t_L g582 ( .A(n_583), .B(n_591), .Y(n_582) );
INVx5_ASAP7_75t_L g621 ( .A(n_583), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g693 ( .A(n_583), .B(n_615), .Y(n_693) );
BUFx2_ASAP7_75t_L g753 ( .A(n_583), .Y(n_753) );
OR2x6_ASAP7_75t_L g583 ( .A(n_584), .B(n_585), .Y(n_583) );
INVx4_ASAP7_75t_L g615 ( .A(n_591), .Y(n_615) );
AND2x2_ASAP7_75t_L g738 ( .A(n_591), .B(n_621), .Y(n_738) );
NAND2xp5_ASAP7_75t_L g592 ( .A(n_593), .B(n_597), .Y(n_592) );
INVx1_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
OAI221xp5_ASAP7_75t_L g727 ( .A1(n_601), .A2(n_728), .B1(n_731), .B2(n_733), .C(n_734), .Y(n_727) );
NAND2xp5_ASAP7_75t_SL g601 ( .A(n_602), .B(n_603), .Y(n_601) );
AND2x2_ASAP7_75t_L g749 ( .A(n_602), .B(n_640), .Y(n_749) );
INVx1_ASAP7_75t_SL g775 ( .A(n_602), .Y(n_775) );
AND2x2_ASAP7_75t_L g760 ( .A(n_603), .B(n_732), .Y(n_760) );
INVx2_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
NOR2xp33_ASAP7_75t_L g705 ( .A(n_604), .B(n_706), .Y(n_705) );
AND2x2_ASAP7_75t_L g605 ( .A(n_606), .B(n_607), .Y(n_605) );
AND2x2_ASAP7_75t_L g629 ( .A(n_606), .B(n_630), .Y(n_629) );
AND2x2_ASAP7_75t_L g635 ( .A(n_606), .B(n_636), .Y(n_635) );
INVx1_ASAP7_75t_L g659 ( .A(n_607), .Y(n_659) );
AND2x2_ASAP7_75t_L g717 ( .A(n_607), .B(n_645), .Y(n_717) );
INVx2_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
BUFx2_ASAP7_75t_L g642 ( .A(n_609), .Y(n_642) );
INVx1_ASAP7_75t_SL g610 ( .A(n_611), .Y(n_610) );
OR2x2_ASAP7_75t_L g611 ( .A(n_612), .B(n_614), .Y(n_611) );
INVx1_ASAP7_75t_L g612 ( .A(n_613), .Y(n_612) );
INVx2_ASAP7_75t_L g638 ( .A(n_614), .Y(n_638) );
OR2x2_ASAP7_75t_L g806 ( .A(n_614), .B(n_807), .Y(n_806) );
INVx2_ASAP7_75t_L g622 ( .A(n_615), .Y(n_622) );
AND2x4_ASAP7_75t_L g678 ( .A(n_615), .B(n_679), .Y(n_678) );
NAND2xp5_ASAP7_75t_L g682 ( .A(n_615), .B(n_683), .Y(n_682) );
NAND2x1p5_ASAP7_75t_L g720 ( .A(n_615), .B(n_621), .Y(n_720) );
AND2x2_ASAP7_75t_L g780 ( .A(n_615), .B(n_683), .Y(n_780) );
AOI22xp33_ASAP7_75t_L g616 ( .A1(n_617), .A2(n_624), .B1(n_637), .B2(n_639), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g698 ( .A(n_617), .B(n_699), .Y(n_698) );
INVx1_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
INVx2_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
AND3x2_ASAP7_75t_L g619 ( .A(n_620), .B(n_622), .C(n_623), .Y(n_619) );
AND2x4_ASAP7_75t_L g637 ( .A(n_620), .B(n_638), .Y(n_637) );
INVx4_ASAP7_75t_L g677 ( .A(n_621), .Y(n_677) );
AND2x2_ASAP7_75t_SL g810 ( .A(n_621), .B(n_678), .Y(n_810) );
NAND2xp5_ASAP7_75t_L g785 ( .A(n_622), .B(n_786), .Y(n_785) );
INVx2_ASAP7_75t_L g722 ( .A(n_623), .Y(n_722) );
AOI322xp5_ASAP7_75t_L g787 ( .A1(n_623), .A2(n_752), .A3(n_788), .B1(n_790), .B2(n_793), .C1(n_797), .C2(n_798), .Y(n_787) );
NAND4xp25_ASAP7_75t_SL g624 ( .A(n_625), .B(n_628), .C(n_632), .D(n_634), .Y(n_624) );
INVx1_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
AND2x2_ASAP7_75t_SL g754 ( .A(n_626), .B(n_642), .Y(n_754) );
BUFx2_ASAP7_75t_L g645 ( .A(n_627), .Y(n_645) );
INVx1_ASAP7_75t_SL g628 ( .A(n_629), .Y(n_628) );
AND2x2_ASAP7_75t_L g769 ( .A(n_630), .B(n_770), .Y(n_769) );
INVx1_ASAP7_75t_L g630 ( .A(n_631), .Y(n_630) );
OR2x2_ASAP7_75t_L g783 ( .A(n_631), .B(n_658), .Y(n_783) );
INVx1_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
AND2x2_ASAP7_75t_L g649 ( .A(n_633), .B(n_650), .Y(n_649) );
OAI211xp5_ASAP7_75t_L g701 ( .A1(n_633), .A2(n_702), .B(n_704), .C(n_707), .Y(n_701) );
NAND2xp5_ASAP7_75t_L g759 ( .A(n_633), .B(n_640), .Y(n_759) );
INVx1_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
AOI22xp5_ASAP7_75t_L g716 ( .A1(n_635), .A2(n_717), .B1(n_718), .B2(n_721), .Y(n_716) );
AOI22xp5_ASAP7_75t_L g671 ( .A1(n_636), .A2(n_672), .B1(n_676), .B2(n_680), .Y(n_671) );
NAND2xp5_ASAP7_75t_L g724 ( .A(n_636), .B(n_725), .Y(n_724) );
NAND2xp5_ASAP7_75t_L g772 ( .A(n_636), .B(n_773), .Y(n_772) );
NAND2xp5_ASAP7_75t_L g794 ( .A(n_636), .B(n_795), .Y(n_794) );
INVx2_ASAP7_75t_L g803 ( .A(n_636), .Y(n_803) );
INVx1_ASAP7_75t_L g742 ( .A(n_637), .Y(n_742) );
OAI21xp33_ASAP7_75t_SL g639 ( .A1(n_640), .A2(n_641), .B(n_643), .Y(n_639) );
INVx1_ASAP7_75t_L g650 ( .A(n_640), .Y(n_650) );
NAND2xp5_ASAP7_75t_L g799 ( .A(n_640), .B(n_645), .Y(n_799) );
INVx1_ASAP7_75t_L g641 ( .A(n_642), .Y(n_641) );
AND2x2_ASAP7_75t_L g735 ( .A(n_642), .B(n_646), .Y(n_735) );
NAND2xp5_ASAP7_75t_L g643 ( .A(n_644), .B(n_646), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g661 ( .A(n_644), .B(n_662), .Y(n_661) );
INVx1_ASAP7_75t_L g644 ( .A(n_645), .Y(n_644) );
OR2x2_ASAP7_75t_L g802 ( .A(n_645), .B(n_803), .Y(n_802) );
INVx1_ASAP7_75t_L g776 ( .A(n_646), .Y(n_776) );
A2O1A1Ixp33_ASAP7_75t_L g647 ( .A1(n_648), .A2(n_651), .B(n_652), .C(n_655), .Y(n_647) );
INVxp67_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
OAI22xp33_ASAP7_75t_SL g762 ( .A1(n_650), .A2(n_681), .B1(n_728), .B2(n_763), .Y(n_762) );
INVx1_ASAP7_75t_SL g652 ( .A(n_653), .Y(n_652) );
NAND2xp5_ASAP7_75t_L g685 ( .A(n_654), .B(n_677), .Y(n_685) );
OR2x2_ASAP7_75t_L g714 ( .A(n_654), .B(n_715), .Y(n_714) );
OAI21xp5_ASAP7_75t_SL g655 ( .A1(n_656), .A2(n_660), .B(n_664), .Y(n_655) );
INVx1_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
OR2x2_ASAP7_75t_L g657 ( .A(n_658), .B(n_659), .Y(n_657) );
INVx1_ASAP7_75t_L g675 ( .A(n_658), .Y(n_675) );
INVx1_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
OAI211xp5_ASAP7_75t_SL g713 ( .A1(n_661), .A2(n_714), .B(n_716), .C(n_724), .Y(n_713) );
INVx1_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
INVx1_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
NOR2xp67_ASAP7_75t_SL g747 ( .A(n_666), .B(n_693), .Y(n_747) );
INVx1_ASAP7_75t_L g750 ( .A(n_666), .Y(n_750) );
INVx2_ASAP7_75t_L g666 ( .A(n_667), .Y(n_666) );
INVx2_ASAP7_75t_L g667 ( .A(n_668), .Y(n_667) );
NAND2xp5_ASAP7_75t_L g807 ( .A(n_668), .B(n_677), .Y(n_807) );
INVx1_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
INVx1_ASAP7_75t_L g679 ( .A(n_669), .Y(n_679) );
INVx2_ASAP7_75t_L g684 ( .A(n_669), .Y(n_684) );
NAND4xp25_ASAP7_75t_L g670 ( .A(n_671), .B(n_686), .C(n_698), .D(n_701), .Y(n_670) );
INVx1_ASAP7_75t_L g672 ( .A(n_673), .Y(n_672) );
OAI22xp33_ASAP7_75t_L g805 ( .A1(n_674), .A2(n_806), .B1(n_808), .B2(n_809), .Y(n_805) );
INVx1_ASAP7_75t_L g674 ( .A(n_675), .Y(n_674) );
AND2x2_ASAP7_75t_L g676 ( .A(n_677), .B(n_678), .Y(n_676) );
AND2x4_ASAP7_75t_L g773 ( .A(n_677), .B(n_703), .Y(n_773) );
AND2x2_ASAP7_75t_L g694 ( .A(n_678), .B(n_695), .Y(n_694) );
INVx2_ASAP7_75t_L g715 ( .A(n_678), .Y(n_715) );
AND2x2_ASAP7_75t_L g725 ( .A(n_678), .B(n_726), .Y(n_725) );
INVx1_ASAP7_75t_L g680 ( .A(n_681), .Y(n_680) );
OR2x2_ASAP7_75t_L g681 ( .A(n_682), .B(n_685), .Y(n_681) );
INVx1_ASAP7_75t_L g683 ( .A(n_684), .Y(n_683) );
HB1xp67_ASAP7_75t_L g739 ( .A(n_684), .Y(n_739) );
INVx1_ASAP7_75t_L g729 ( .A(n_685), .Y(n_729) );
AOI32xp33_ASAP7_75t_L g686 ( .A1(n_687), .A2(n_690), .A3(n_693), .B1(n_694), .B2(n_696), .Y(n_686) );
OAI21xp33_ASAP7_75t_L g734 ( .A1(n_687), .A2(n_735), .B(n_736), .Y(n_734) );
INVx2_ASAP7_75t_L g687 ( .A(n_688), .Y(n_687) );
AOI221xp5_ASAP7_75t_L g766 ( .A1(n_690), .A2(n_767), .B1(n_769), .B2(n_771), .C(n_774), .Y(n_766) );
INVx1_ASAP7_75t_SL g690 ( .A(n_691), .Y(n_690) );
INVx1_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
AND2x2_ASAP7_75t_L g751 ( .A(n_692), .B(n_752), .Y(n_751) );
INVx1_ASAP7_75t_L g709 ( .A(n_693), .Y(n_709) );
AOI22xp5_ASAP7_75t_L g781 ( .A1(n_694), .A2(n_732), .B1(n_782), .B2(n_784), .Y(n_781) );
INVx1_ASAP7_75t_L g708 ( .A(n_695), .Y(n_708) );
AND2x2_ASAP7_75t_L g786 ( .A(n_695), .B(n_739), .Y(n_786) );
INVx1_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
NAND2xp5_ASAP7_75t_SL g789 ( .A(n_702), .B(n_754), .Y(n_789) );
INVx1_ASAP7_75t_L g808 ( .A(n_702), .Y(n_808) );
INVx1_ASAP7_75t_SL g702 ( .A(n_703), .Y(n_702) );
INVx1_ASAP7_75t_L g704 ( .A(n_705), .Y(n_704) );
AND2x2_ASAP7_75t_L g707 ( .A(n_708), .B(n_709), .Y(n_707) );
NOR2xp67_ASAP7_75t_L g710 ( .A(n_711), .B(n_765), .Y(n_710) );
NAND2xp5_ASAP7_75t_L g711 ( .A(n_712), .B(n_755), .Y(n_711) );
NOR3xp33_ASAP7_75t_SL g712 ( .A(n_713), .B(n_727), .C(n_740), .Y(n_712) );
INVx1_ASAP7_75t_L g730 ( .A(n_715), .Y(n_730) );
INVx1_ASAP7_75t_SL g741 ( .A(n_717), .Y(n_741) );
INVx2_ASAP7_75t_L g718 ( .A(n_719), .Y(n_718) );
INVx2_ASAP7_75t_L g723 ( .A(n_720), .Y(n_723) );
INVx2_ASAP7_75t_L g733 ( .A(n_721), .Y(n_733) );
AND2x2_ASAP7_75t_L g721 ( .A(n_722), .B(n_723), .Y(n_721) );
AND2x4_ASAP7_75t_L g779 ( .A(n_722), .B(n_780), .Y(n_779) );
AND2x4_ASAP7_75t_L g797 ( .A(n_726), .B(n_780), .Y(n_797) );
NAND2xp5_ASAP7_75t_SL g728 ( .A(n_729), .B(n_730), .Y(n_728) );
INVx1_ASAP7_75t_SL g731 ( .A(n_732), .Y(n_731) );
NOR2xp33_ASAP7_75t_L g736 ( .A(n_737), .B(n_739), .Y(n_736) );
AOI32xp33_ASAP7_75t_L g748 ( .A1(n_737), .A2(n_749), .A3(n_750), .B1(n_751), .B2(n_754), .Y(n_748) );
NOR2xp33_ASAP7_75t_SL g767 ( .A(n_737), .B(n_768), .Y(n_767) );
INVx2_ASAP7_75t_SL g737 ( .A(n_738), .Y(n_737) );
INVx1_ASAP7_75t_L g768 ( .A(n_739), .Y(n_768) );
OAI211xp5_ASAP7_75t_SL g740 ( .A1(n_741), .A2(n_742), .B(n_743), .C(n_748), .Y(n_740) );
NAND2xp5_ASAP7_75t_L g743 ( .A(n_744), .B(n_747), .Y(n_743) );
INVx1_ASAP7_75t_L g744 ( .A(n_745), .Y(n_744) );
AND2x2_ASAP7_75t_L g804 ( .A(n_752), .B(n_792), .Y(n_804) );
INVx2_ASAP7_75t_L g752 ( .A(n_753), .Y(n_752) );
NAND2xp5_ASAP7_75t_L g791 ( .A(n_753), .B(n_792), .Y(n_791) );
AOI221xp5_ASAP7_75t_L g755 ( .A1(n_756), .A2(n_758), .B1(n_760), .B2(n_761), .C(n_762), .Y(n_755) );
INVx1_ASAP7_75t_SL g758 ( .A(n_759), .Y(n_758) );
CKINVDCx16_ASAP7_75t_R g763 ( .A(n_764), .Y(n_763) );
NAND4xp25_ASAP7_75t_L g765 ( .A(n_766), .B(n_781), .C(n_787), .D(n_800), .Y(n_765) );
INVxp33_ASAP7_75t_L g771 ( .A(n_772), .Y(n_771) );
O2A1O1Ixp33_ASAP7_75t_L g774 ( .A1(n_775), .A2(n_776), .B(n_777), .C(n_778), .Y(n_774) );
INVx2_ASAP7_75t_L g778 ( .A(n_779), .Y(n_778) );
INVx1_ASAP7_75t_L g782 ( .A(n_783), .Y(n_782) );
INVx1_ASAP7_75t_SL g784 ( .A(n_785), .Y(n_784) );
INVx1_ASAP7_75t_L g788 ( .A(n_789), .Y(n_788) );
INVx1_ASAP7_75t_L g790 ( .A(n_791), .Y(n_790) );
INVx1_ASAP7_75t_SL g793 ( .A(n_794), .Y(n_793) );
INVx1_ASAP7_75t_L g798 ( .A(n_799), .Y(n_798) );
INVx2_ASAP7_75t_L g801 ( .A(n_802), .Y(n_801) );
INVx3_ASAP7_75t_SL g809 ( .A(n_810), .Y(n_809) );
BUFx2_ASAP7_75t_L g812 ( .A(n_813), .Y(n_812) );
CKINVDCx5p33_ASAP7_75t_R g814 ( .A(n_815), .Y(n_814) );
NAND2xp5_ASAP7_75t_L g816 ( .A(n_817), .B(n_831), .Y(n_816) );
AOI31xp33_ASAP7_75t_L g817 ( .A1(n_818), .A2(n_822), .A3(n_829), .B(n_830), .Y(n_817) );
INVx1_ASAP7_75t_L g818 ( .A(n_819), .Y(n_818) );
OR3x1_ASAP7_75t_L g831 ( .A(n_819), .B(n_822), .C(n_829), .Y(n_831) );
INVx1_ASAP7_75t_L g819 ( .A(n_820), .Y(n_819) );
HB1xp67_ASAP7_75t_L g820 ( .A(n_821), .Y(n_820) );
INVx1_ASAP7_75t_L g827 ( .A(n_824), .Y(n_827) );
NOR2xp33_ASAP7_75t_L g832 ( .A(n_833), .B(n_834), .Y(n_832) );
endmodule