module fake_jpeg_2327_n_329 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_329);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_329;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_0),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_3),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

BUFx10_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

INVx3_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

INVx4_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_10),
.Y(n_24)
);

BUFx8_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_2),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_11),
.Y(n_28)
);

BUFx10_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

INVx2_ASAP7_75t_SL g31 ( 
.A(n_10),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_6),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_2),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_1),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_22),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_19),
.Y(n_37)
);

INVx2_ASAP7_75t_SL g89 ( 
.A(n_37),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_22),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_38),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g39 ( 
.A(n_24),
.B(n_7),
.Y(n_39)
);

OR2x2_ASAP7_75t_L g57 ( 
.A(n_39),
.B(n_31),
.Y(n_57)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_40),
.Y(n_63)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_30),
.Y(n_41)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_41),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_22),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_42),
.Y(n_97)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_25),
.Y(n_43)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_43),
.Y(n_55)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_19),
.Y(n_44)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_44),
.Y(n_71)
);

AND2x2_ASAP7_75t_L g45 ( 
.A(n_30),
.B(n_0),
.Y(n_45)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_45),
.B(n_31),
.Y(n_58)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_25),
.Y(n_46)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_46),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_18),
.B(n_0),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_47),
.B(n_51),
.Y(n_54)
);

BUFx5_ASAP7_75t_L g48 ( 
.A(n_25),
.Y(n_48)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_48),
.Y(n_53)
);

INVx2_ASAP7_75t_SL g49 ( 
.A(n_25),
.Y(n_49)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_49),
.Y(n_96)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_25),
.Y(n_50)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_50),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_18),
.B(n_1),
.Y(n_51)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_36),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_56),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_57),
.B(n_59),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_58),
.B(n_78),
.Y(n_106)
);

NOR2xp67_ASAP7_75t_L g59 ( 
.A(n_39),
.B(n_23),
.Y(n_59)
);

INVx11_ASAP7_75t_L g60 ( 
.A(n_43),
.Y(n_60)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_60),
.Y(n_113)
);

NOR2x1_ASAP7_75t_L g61 ( 
.A(n_47),
.B(n_23),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_61),
.B(n_64),
.Y(n_127)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_37),
.Y(n_62)
);

INVx1_ASAP7_75t_SL g105 ( 
.A(n_62),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_51),
.B(n_32),
.Y(n_64)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_36),
.Y(n_65)
);

BUFx2_ASAP7_75t_L g129 ( 
.A(n_65),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_45),
.A2(n_18),
.B1(n_21),
.B2(n_20),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_66),
.A2(n_72),
.B1(n_75),
.B2(n_81),
.Y(n_117)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_38),
.Y(n_67)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_67),
.Y(n_102)
);

OAI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_40),
.A2(n_41),
.B1(n_38),
.B2(n_42),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_68),
.A2(n_82),
.B1(n_34),
.B2(n_33),
.Y(n_120)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_44),
.Y(n_70)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_70),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_45),
.A2(n_19),
.B1(n_20),
.B2(n_21),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_43),
.B(n_28),
.Y(n_73)
);

CKINVDCx16_ASAP7_75t_R g124 ( 
.A(n_73),
.Y(n_124)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_49),
.Y(n_74)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_74),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_43),
.A2(n_49),
.B1(n_50),
.B2(n_46),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_50),
.B(n_28),
.Y(n_76)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_76),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_42),
.B(n_24),
.Y(n_78)
);

BUFx12_ASAP7_75t_L g80 ( 
.A(n_48),
.Y(n_80)
);

INVx13_ASAP7_75t_L g125 ( 
.A(n_80),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_47),
.A2(n_20),
.B1(n_21),
.B2(n_35),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_47),
.A2(n_20),
.B1(n_21),
.B2(n_35),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_43),
.A2(n_31),
.B1(n_35),
.B2(n_26),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_83),
.A2(n_99),
.B1(n_100),
.B2(n_101),
.Y(n_111)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_40),
.Y(n_84)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_84),
.Y(n_126)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_50),
.Y(n_85)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_85),
.Y(n_115)
);

INVx5_ASAP7_75t_L g86 ( 
.A(n_43),
.Y(n_86)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_86),
.Y(n_119)
);

INVx13_ASAP7_75t_L g87 ( 
.A(n_49),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_87),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_39),
.B(n_32),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_88),
.B(n_93),
.Y(n_121)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_50),
.Y(n_91)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_91),
.Y(n_130)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_45),
.B(n_31),
.Y(n_92)
);

XNOR2xp5_ASAP7_75t_L g108 ( 
.A(n_92),
.B(n_98),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_39),
.B(n_33),
.Y(n_93)
);

CKINVDCx12_ASAP7_75t_R g94 ( 
.A(n_43),
.Y(n_94)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_94),
.Y(n_131)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_40),
.Y(n_95)
);

INVx6_ASAP7_75t_L g133 ( 
.A(n_95),
.Y(n_133)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_45),
.B(n_34),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_47),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_43),
.A2(n_22),
.B1(n_26),
.B2(n_16),
.Y(n_100)
);

BUFx12f_ASAP7_75t_L g101 ( 
.A(n_37),
.Y(n_101)
);

AO22x1_ASAP7_75t_SL g104 ( 
.A1(n_58),
.A2(n_26),
.B1(n_16),
.B2(n_17),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_104),
.B(n_114),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_L g112 ( 
.A1(n_68),
.A2(n_27),
.B1(n_14),
.B2(n_15),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_112),
.A2(n_120),
.B1(n_123),
.B2(n_128),
.Y(n_153)
);

AO22x1_ASAP7_75t_SL g114 ( 
.A1(n_92),
.A2(n_26),
.B1(n_16),
.B2(n_17),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_96),
.A2(n_98),
.B1(n_15),
.B2(n_14),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g137 ( 
.A(n_118),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_96),
.A2(n_27),
.B1(n_17),
.B2(n_29),
.Y(n_123)
);

OAI22xp33_ASAP7_75t_L g128 ( 
.A1(n_100),
.A2(n_17),
.B1(n_29),
.B2(n_4),
.Y(n_128)
);

AO22x2_ASAP7_75t_L g132 ( 
.A1(n_83),
.A2(n_17),
.B1(n_29),
.B2(n_4),
.Y(n_132)
);

HB1xp67_ASAP7_75t_L g158 ( 
.A(n_132),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_106),
.B(n_54),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_135),
.B(n_114),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_124),
.B(n_61),
.Y(n_136)
);

CKINVDCx14_ASAP7_75t_R g179 ( 
.A(n_136),
.Y(n_179)
);

INVx8_ASAP7_75t_L g138 ( 
.A(n_110),
.Y(n_138)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_138),
.Y(n_176)
);

INVx4_ASAP7_75t_L g139 ( 
.A(n_115),
.Y(n_139)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_139),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_SL g140 ( 
.A1(n_111),
.A2(n_57),
.B(n_75),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_SL g184 ( 
.A1(n_140),
.A2(n_132),
.B(n_105),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_107),
.B(n_63),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_141),
.B(n_154),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_120),
.A2(n_69),
.B1(n_56),
.B2(n_65),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_142),
.A2(n_97),
.B1(n_79),
.B2(n_52),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g143 ( 
.A(n_108),
.B(n_89),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_143),
.B(n_149),
.Y(n_194)
);

AND2x2_ASAP7_75t_L g144 ( 
.A(n_122),
.B(n_77),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_SL g175 ( 
.A(n_144),
.B(n_145),
.Y(n_175)
);

AND2x2_ASAP7_75t_L g145 ( 
.A(n_108),
.B(n_90),
.Y(n_145)
);

INVx2_ASAP7_75t_SL g146 ( 
.A(n_129),
.Y(n_146)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_146),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g147 ( 
.A(n_102),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g178 ( 
.A(n_147),
.Y(n_178)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_103),
.Y(n_148)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_148),
.Y(n_187)
);

CKINVDCx16_ASAP7_75t_R g149 ( 
.A(n_125),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_126),
.Y(n_150)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_150),
.Y(n_195)
);

FAx1_ASAP7_75t_SL g151 ( 
.A(n_106),
.B(n_87),
.CI(n_89),
.CON(n_151),
.SN(n_151)
);

OAI32xp33_ASAP7_75t_L g182 ( 
.A1(n_151),
.A2(n_132),
.A3(n_105),
.B1(n_113),
.B2(n_128),
.Y(n_182)
);

INVxp33_ASAP7_75t_L g152 ( 
.A(n_131),
.Y(n_152)
);

INVxp67_ASAP7_75t_L g192 ( 
.A(n_152),
.Y(n_192)
);

AND2x2_ASAP7_75t_L g154 ( 
.A(n_104),
.B(n_55),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_102),
.Y(n_155)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_155),
.Y(n_197)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_133),
.Y(n_156)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_156),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_109),
.B(n_127),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_157),
.B(n_160),
.Y(n_173)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_126),
.Y(n_159)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_159),
.Y(n_204)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_133),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_129),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_161),
.B(n_162),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_121),
.B(n_71),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_113),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_163),
.B(n_165),
.Y(n_186)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_115),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_SL g190 ( 
.A1(n_164),
.A2(n_166),
.B1(n_168),
.B2(n_101),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_121),
.B(n_97),
.Y(n_165)
);

INVx4_ASAP7_75t_L g166 ( 
.A(n_116),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_116),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_167),
.B(n_169),
.Y(n_201)
);

INVx4_ASAP7_75t_L g168 ( 
.A(n_125),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_130),
.B(n_62),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g170 ( 
.A(n_119),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_170),
.Y(n_189)
);

AO21x1_ASAP7_75t_L g171 ( 
.A1(n_134),
.A2(n_114),
.B(n_104),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_SL g220 ( 
.A1(n_171),
.A2(n_184),
.B(n_185),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_174),
.B(n_181),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_135),
.B(n_117),
.Y(n_181)
);

AND2x2_ASAP7_75t_L g222 ( 
.A(n_182),
.B(n_188),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_143),
.B(n_67),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_183),
.B(n_206),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_137),
.A2(n_132),
.B1(n_53),
.B2(n_80),
.Y(n_185)
);

INVxp67_ASAP7_75t_L g227 ( 
.A(n_190),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_134),
.A2(n_79),
.B1(n_52),
.B2(n_62),
.Y(n_191)
);

AOI22xp33_ASAP7_75t_SL g224 ( 
.A1(n_191),
.A2(n_146),
.B1(n_164),
.B2(n_166),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_170),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_193),
.B(n_203),
.Y(n_215)
);

AOI21xp5_ASAP7_75t_L g196 ( 
.A1(n_140),
.A2(n_101),
.B(n_17),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_L g223 ( 
.A1(n_196),
.A2(n_205),
.B(n_153),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_158),
.A2(n_29),
.B1(n_8),
.B2(n_9),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_200),
.A2(n_142),
.B1(n_174),
.B2(n_186),
.Y(n_213)
);

OR2x4_ASAP7_75t_L g202 ( 
.A(n_151),
.B(n_29),
.Y(n_202)
);

OR2x2_ASAP7_75t_L g232 ( 
.A(n_202),
.B(n_156),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_144),
.Y(n_203)
);

AOI21xp5_ASAP7_75t_L g205 ( 
.A1(n_137),
.A2(n_29),
.B(n_2),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_151),
.B(n_1),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_145),
.B(n_1),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_207),
.B(n_168),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_208),
.B(n_214),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_192),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_209),
.B(n_211),
.Y(n_236)
);

AND2x6_ASAP7_75t_L g210 ( 
.A(n_202),
.B(n_154),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_210),
.B(n_212),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_179),
.B(n_152),
.Y(n_211)
);

AND2x6_ASAP7_75t_L g212 ( 
.A(n_181),
.B(n_196),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_213),
.A2(n_233),
.B1(n_234),
.B2(n_180),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_SL g214 ( 
.A(n_173),
.B(n_139),
.Y(n_214)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_187),
.Y(n_216)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_216),
.Y(n_238)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_187),
.Y(n_217)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_217),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_192),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_218),
.B(n_225),
.Y(n_242)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_195),
.Y(n_221)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_221),
.Y(n_241)
);

INVx1_ASAP7_75t_SL g247 ( 
.A(n_223),
.Y(n_247)
);

INVxp67_ASAP7_75t_L g244 ( 
.A(n_224),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_201),
.Y(n_225)
);

AND2x6_ASAP7_75t_L g226 ( 
.A(n_184),
.B(n_12),
.Y(n_226)
);

INVxp67_ASAP7_75t_L g249 ( 
.A(n_226),
.Y(n_249)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_195),
.Y(n_228)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_228),
.Y(n_248)
);

NAND3xp33_ASAP7_75t_L g229 ( 
.A(n_203),
.B(n_12),
.C(n_5),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_229),
.Y(n_243)
);

INVxp67_ASAP7_75t_L g230 ( 
.A(n_199),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_230),
.Y(n_245)
);

AOI21xp5_ASAP7_75t_L g253 ( 
.A1(n_232),
.A2(n_205),
.B(n_175),
.Y(n_253)
);

CKINVDCx16_ASAP7_75t_R g233 ( 
.A(n_177),
.Y(n_233)
);

INVx2_ASAP7_75t_SL g234 ( 
.A(n_198),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_SL g235 ( 
.A(n_172),
.B(n_10),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_235),
.B(n_206),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_219),
.B(n_194),
.C(n_183),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_237),
.B(n_251),
.C(n_254),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g269 ( 
.A(n_246),
.B(n_217),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_L g264 ( 
.A1(n_250),
.A2(n_255),
.B1(n_218),
.B2(n_215),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_219),
.B(n_220),
.C(n_231),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_231),
.B(n_175),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_252),
.B(n_258),
.Y(n_263)
);

INVx1_ASAP7_75t_SL g265 ( 
.A(n_253),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_220),
.B(n_207),
.C(n_204),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_222),
.A2(n_223),
.B1(n_232),
.B2(n_213),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_222),
.B(n_204),
.C(n_185),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_257),
.B(n_258),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_222),
.B(n_182),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_245),
.B(n_209),
.Y(n_259)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_259),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_242),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_SL g287 ( 
.A(n_260),
.B(n_261),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_236),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_264),
.A2(n_272),
.B1(n_274),
.B2(n_275),
.Y(n_277)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_248),
.Y(n_266)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_266),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_252),
.B(n_225),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_SL g288 ( 
.A(n_267),
.B(n_269),
.Y(n_288)
);

INVxp67_ASAP7_75t_L g268 ( 
.A(n_239),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_L g284 ( 
.A1(n_268),
.A2(n_271),
.B1(n_273),
.B2(n_250),
.Y(n_284)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_270),
.B(n_276),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_246),
.B(n_199),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_238),
.Y(n_272)
);

CKINVDCx14_ASAP7_75t_R g273 ( 
.A(n_256),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_255),
.A2(n_212),
.B1(n_210),
.B2(n_226),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_247),
.A2(n_227),
.B1(n_171),
.B2(n_216),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g276 ( 
.A(n_251),
.B(n_221),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_262),
.B(n_254),
.C(n_249),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_SL g292 ( 
.A(n_279),
.B(n_285),
.Y(n_292)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_270),
.B(n_262),
.Y(n_281)
);

XOR2xp5_ASAP7_75t_L g291 ( 
.A(n_281),
.B(n_283),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_SL g283 ( 
.A(n_263),
.B(n_237),
.Y(n_283)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_284),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_268),
.B(n_249),
.C(n_247),
.Y(n_285)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_276),
.B(n_257),
.Y(n_286)
);

XOR2xp5_ASAP7_75t_L g296 ( 
.A(n_286),
.B(n_272),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_263),
.B(n_253),
.C(n_241),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_289),
.B(n_290),
.C(n_240),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_259),
.B(n_265),
.C(n_275),
.Y(n_290)
);

OAI21xp5_ASAP7_75t_L g294 ( 
.A1(n_290),
.A2(n_265),
.B(n_274),
.Y(n_294)
);

XOR2xp5_ASAP7_75t_L g305 ( 
.A(n_294),
.B(n_296),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_281),
.B(n_266),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g304 ( 
.A(n_295),
.B(n_298),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_288),
.B(n_243),
.Y(n_297)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_297),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_278),
.B(n_286),
.C(n_283),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_SL g307 ( 
.A(n_299),
.B(n_278),
.Y(n_307)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_287),
.Y(n_300)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_300),
.Y(n_306)
);

OAI21xp5_ASAP7_75t_L g301 ( 
.A1(n_280),
.A2(n_244),
.B(n_227),
.Y(n_301)
);

XOR2xp5_ASAP7_75t_L g309 ( 
.A(n_301),
.B(n_200),
.Y(n_309)
);

AOI21xp5_ASAP7_75t_L g302 ( 
.A1(n_289),
.A2(n_244),
.B(n_230),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_302),
.B(n_180),
.C(n_178),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_307),
.B(n_310),
.Y(n_313)
);

A2O1A1O1Ixp25_ASAP7_75t_L g308 ( 
.A1(n_294),
.A2(n_277),
.B(n_282),
.C(n_228),
.D(n_189),
.Y(n_308)
);

AOI21xp5_ASAP7_75t_L g318 ( 
.A1(n_308),
.A2(n_189),
.B(n_193),
.Y(n_318)
);

XOR2xp5_ASAP7_75t_L g316 ( 
.A(n_309),
.B(n_305),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_L g311 ( 
.A(n_296),
.B(n_295),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_311),
.B(n_299),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_SL g312 ( 
.A1(n_308),
.A2(n_293),
.B1(n_292),
.B2(n_301),
.Y(n_312)
);

INVxp67_ASAP7_75t_L g321 ( 
.A(n_312),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_306),
.A2(n_298),
.B1(n_234),
.B2(n_188),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g319 ( 
.A1(n_314),
.A2(n_316),
.B1(n_309),
.B2(n_305),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_315),
.B(n_318),
.Y(n_320)
);

OAI21xp5_ASAP7_75t_SL g317 ( 
.A1(n_303),
.A2(n_291),
.B(n_234),
.Y(n_317)
);

OAI21xp5_ASAP7_75t_L g322 ( 
.A1(n_317),
.A2(n_304),
.B(n_291),
.Y(n_322)
);

OAI21xp5_ASAP7_75t_L g323 ( 
.A1(n_319),
.A2(n_322),
.B(n_320),
.Y(n_323)
);

OAI21xp33_ASAP7_75t_SL g325 ( 
.A1(n_323),
.A2(n_324),
.B(n_176),
.Y(n_325)
);

AOI22xp33_ASAP7_75t_SL g324 ( 
.A1(n_321),
.A2(n_312),
.B1(n_313),
.B2(n_316),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_325),
.B(n_176),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_326),
.B(n_198),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_327),
.B(n_197),
.Y(n_328)
);

XNOR2xp5_ASAP7_75t_L g329 ( 
.A(n_328),
.B(n_197),
.Y(n_329)
);


endmodule