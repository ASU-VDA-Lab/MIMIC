module fake_aes_9759_n_39 (n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_39);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_39;
wire n_20;
wire n_38;
wire n_36;
wire n_37;
wire n_34;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_30;
wire n_33;
wire n_18;
wire n_32;
wire n_35;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_27;
XOR2xp5_ASAP7_75t_L g11 ( .A(n_3), .B(n_7), .Y(n_11) );
CKINVDCx5p33_ASAP7_75t_R g12 ( .A(n_2), .Y(n_12) );
AOI22xp5_ASAP7_75t_L g13 ( .A1(n_10), .A2(n_2), .B1(n_1), .B2(n_0), .Y(n_13) );
AND2x2_ASAP7_75t_L g14 ( .A(n_6), .B(n_5), .Y(n_14) );
INVx1_ASAP7_75t_L g15 ( .A(n_1), .Y(n_15) );
NOR2xp33_ASAP7_75t_L g16 ( .A(n_9), .B(n_8), .Y(n_16) );
INVx2_ASAP7_75t_L g17 ( .A(n_15), .Y(n_17) );
CKINVDCx5p33_ASAP7_75t_R g18 ( .A(n_12), .Y(n_18) );
INVx3_ASAP7_75t_L g19 ( .A(n_12), .Y(n_19) );
AOI22xp5_ASAP7_75t_L g20 ( .A1(n_13), .A2(n_0), .B1(n_3), .B2(n_4), .Y(n_20) );
OAI21x1_ASAP7_75t_L g21 ( .A1(n_17), .A2(n_14), .B(n_16), .Y(n_21) );
AND2x4_ASAP7_75t_L g22 ( .A(n_19), .B(n_14), .Y(n_22) );
INVx2_ASAP7_75t_L g23 ( .A(n_17), .Y(n_23) );
INVx3_ASAP7_75t_L g24 ( .A(n_23), .Y(n_24) );
INVx1_ASAP7_75t_L g25 ( .A(n_23), .Y(n_25) );
AND2x2_ASAP7_75t_L g26 ( .A(n_25), .B(n_18), .Y(n_26) );
AOI211xp5_ASAP7_75t_L g27 ( .A1(n_25), .A2(n_20), .B(n_19), .C(n_22), .Y(n_27) );
NAND2xp5_ASAP7_75t_L g28 ( .A(n_27), .B(n_22), .Y(n_28) );
INVx1_ASAP7_75t_L g29 ( .A(n_26), .Y(n_29) );
OR2x2_ASAP7_75t_L g30 ( .A(n_29), .B(n_22), .Y(n_30) );
AOI22xp5_ASAP7_75t_L g31 ( .A1(n_28), .A2(n_11), .B1(n_22), .B2(n_24), .Y(n_31) );
AOI21xp5_ASAP7_75t_SL g32 ( .A1(n_28), .A2(n_23), .B(n_21), .Y(n_32) );
NOR2xp33_ASAP7_75t_L g33 ( .A(n_31), .B(n_21), .Y(n_33) );
HB1xp67_ASAP7_75t_L g34 ( .A(n_30), .Y(n_34) );
NAND3xp33_ASAP7_75t_SL g35 ( .A(n_32), .B(n_4), .C(n_24), .Y(n_35) );
BUFx3_ASAP7_75t_L g36 ( .A(n_34), .Y(n_36) );
NAND2xp5_ASAP7_75t_L g37 ( .A(n_33), .B(n_24), .Y(n_37) );
INVx2_ASAP7_75t_L g38 ( .A(n_36), .Y(n_38) );
OAI22xp33_ASAP7_75t_L g39 ( .A1(n_38), .A2(n_37), .B1(n_35), .B2(n_24), .Y(n_39) );
endmodule