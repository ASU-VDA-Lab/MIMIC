module fake_jpeg_1322_n_378 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_378);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_378;

wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

INVx6_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

BUFx10_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

BUFx12_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_5),
.Y(n_21)
);

CKINVDCx16_ASAP7_75t_R g22 ( 
.A(n_12),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_9),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_7),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_10),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_3),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_5),
.Y(n_32)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_5),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_7),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_2),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_2),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_4),
.Y(n_39)
);

INVx1_ASAP7_75t_SL g40 ( 
.A(n_1),
.Y(n_40)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_11),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_9),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_3),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_11),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_14),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_15),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_46),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_22),
.B(n_14),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_47),
.B(n_63),
.Y(n_109)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_20),
.Y(n_48)
);

INVx4_ASAP7_75t_SL g110 ( 
.A(n_48),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_15),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_49),
.Y(n_114)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_41),
.Y(n_50)
);

INVx2_ASAP7_75t_SL g143 ( 
.A(n_50),
.Y(n_143)
);

OR2x2_ASAP7_75t_L g51 ( 
.A(n_25),
.B(n_13),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_51),
.B(n_64),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_15),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_52),
.Y(n_142)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_27),
.Y(n_53)
);

HB1xp67_ASAP7_75t_L g136 ( 
.A(n_53),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_16),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_54),
.Y(n_146)
);

INVx11_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

INVx11_ASAP7_75t_L g116 ( 
.A(n_55),
.Y(n_116)
);

INVx11_ASAP7_75t_L g56 ( 
.A(n_36),
.Y(n_56)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_56),
.Y(n_106)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_36),
.Y(n_57)
);

INVx5_ASAP7_75t_L g117 ( 
.A(n_57),
.Y(n_117)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_20),
.Y(n_58)
);

INVx5_ASAP7_75t_L g118 ( 
.A(n_58),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_16),
.Y(n_59)
);

INVx6_ASAP7_75t_L g152 ( 
.A(n_59),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_16),
.Y(n_60)
);

BUFx12f_ASAP7_75t_L g137 ( 
.A(n_60),
.Y(n_137)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_33),
.Y(n_61)
);

INVx4_ASAP7_75t_L g129 ( 
.A(n_61),
.Y(n_129)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_44),
.Y(n_62)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_62),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_40),
.B(n_42),
.Y(n_63)
);

OR2x2_ASAP7_75t_L g64 ( 
.A(n_25),
.B(n_13),
.Y(n_64)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_33),
.Y(n_65)
);

INVx4_ASAP7_75t_L g132 ( 
.A(n_65),
.Y(n_132)
);

INVx6_ASAP7_75t_SL g66 ( 
.A(n_18),
.Y(n_66)
);

INVx5_ASAP7_75t_SL g122 ( 
.A(n_66),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_19),
.Y(n_67)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_67),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_19),
.Y(n_68)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_68),
.Y(n_123)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_35),
.Y(n_69)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_69),
.Y(n_99)
);

BUFx5_ASAP7_75t_L g70 ( 
.A(n_35),
.Y(n_70)
);

BUFx5_ASAP7_75t_L g126 ( 
.A(n_70),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_19),
.Y(n_71)
);

INVx4_ASAP7_75t_L g145 ( 
.A(n_71),
.Y(n_145)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_27),
.Y(n_72)
);

HB1xp67_ASAP7_75t_L g148 ( 
.A(n_72),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_17),
.Y(n_73)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_73),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_17),
.Y(n_74)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_74),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_36),
.Y(n_75)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_75),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_37),
.Y(n_76)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_76),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_37),
.Y(n_77)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_77),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_40),
.B(n_9),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g150 ( 
.A(n_78),
.B(n_89),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_37),
.Y(n_79)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_79),
.Y(n_121)
);

INVx5_ASAP7_75t_L g80 ( 
.A(n_31),
.Y(n_80)
);

BUFx5_ASAP7_75t_L g139 ( 
.A(n_80),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_37),
.Y(n_81)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_81),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_38),
.Y(n_82)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_82),
.Y(n_138)
);

BUFx4f_ASAP7_75t_SL g83 ( 
.A(n_20),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_83),
.B(n_88),
.Y(n_128)
);

BUFx3_ASAP7_75t_L g84 ( 
.A(n_31),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g151 ( 
.A(n_84),
.B(n_92),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_38),
.Y(n_85)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_85),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_26),
.B(n_23),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_86),
.B(n_93),
.Y(n_101)
);

INVx11_ASAP7_75t_L g87 ( 
.A(n_18),
.Y(n_87)
);

AOI21xp33_ASAP7_75t_L g124 ( 
.A1(n_87),
.A2(n_90),
.B(n_20),
.Y(n_124)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_44),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_23),
.B(n_13),
.Y(n_89)
);

INVx11_ASAP7_75t_L g90 ( 
.A(n_18),
.Y(n_90)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_45),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_91),
.B(n_96),
.Y(n_131)
);

INVx8_ASAP7_75t_L g92 ( 
.A(n_18),
.Y(n_92)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_45),
.Y(n_93)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_41),
.Y(n_94)
);

OR2x2_ASAP7_75t_L g111 ( 
.A(n_94),
.B(n_95),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_29),
.B(n_0),
.Y(n_95)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_26),
.Y(n_96)
);

INVx6_ASAP7_75t_L g97 ( 
.A(n_28),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_97),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_89),
.B(n_42),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_103),
.B(n_113),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_63),
.A2(n_28),
.B1(n_29),
.B2(n_34),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_104),
.A2(n_107),
.B1(n_130),
.B2(n_141),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_78),
.A2(n_43),
.B1(n_39),
.B2(n_34),
.Y(n_105)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_105),
.B(n_5),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_95),
.A2(n_43),
.B1(n_39),
.B2(n_32),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_82),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_112),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_47),
.B(n_32),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_51),
.B(n_24),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_115),
.B(n_85),
.Y(n_163)
);

AOI21xp5_ASAP7_75t_L g158 ( 
.A1(n_124),
.A2(n_58),
.B(n_3),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_64),
.A2(n_30),
.B1(n_24),
.B2(n_21),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_83),
.B(n_30),
.Y(n_134)
);

CKINVDCx14_ASAP7_75t_R g156 ( 
.A(n_134),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_L g141 ( 
.A1(n_73),
.A2(n_21),
.B1(n_1),
.B2(n_2),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_74),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_144),
.A2(n_7),
.B1(n_105),
.B2(n_152),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_48),
.B(n_8),
.Y(n_149)
);

CKINVDCx14_ASAP7_75t_R g183 ( 
.A(n_149),
.Y(n_183)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_138),
.Y(n_154)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_154),
.Y(n_200)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_147),
.Y(n_155)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_155),
.Y(n_194)
);

AOI22xp33_ASAP7_75t_SL g157 ( 
.A1(n_102),
.A2(n_92),
.B1(n_57),
.B2(n_79),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g197 ( 
.A(n_157),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_SL g212 ( 
.A1(n_158),
.A2(n_118),
.B(n_122),
.Y(n_212)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_120),
.Y(n_159)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_159),
.Y(n_198)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_131),
.Y(n_160)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_160),
.Y(n_201)
);

AOI22xp33_ASAP7_75t_L g162 ( 
.A1(n_108),
.A2(n_54),
.B1(n_71),
.B2(n_68),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_162),
.A2(n_164),
.B1(n_137),
.B2(n_110),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_163),
.B(n_173),
.Y(n_214)
);

AOI22xp33_ASAP7_75t_L g164 ( 
.A1(n_108),
.A2(n_49),
.B1(n_52),
.B2(n_59),
.Y(n_164)
);

AOI32xp33_ASAP7_75t_L g165 ( 
.A1(n_98),
.A2(n_81),
.A3(n_77),
.B1(n_76),
.B2(n_75),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_165),
.B(n_174),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_111),
.A2(n_67),
.B1(n_60),
.B2(n_46),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_166),
.A2(n_181),
.B1(n_187),
.B2(n_188),
.Y(n_195)
);

O2A1O1Ixp33_ASAP7_75t_SL g167 ( 
.A1(n_141),
.A2(n_8),
.B(n_3),
.C(n_4),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_L g213 ( 
.A1(n_167),
.A2(n_168),
.B(n_148),
.Y(n_213)
);

AOI21xp5_ASAP7_75t_L g168 ( 
.A1(n_111),
.A2(n_0),
.B(n_4),
.Y(n_168)
);

INVx3_ASAP7_75t_L g169 ( 
.A(n_117),
.Y(n_169)
);

INVx4_ASAP7_75t_SL g192 ( 
.A(n_169),
.Y(n_192)
);

BUFx4f_ASAP7_75t_L g170 ( 
.A(n_145),
.Y(n_170)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_170),
.Y(n_207)
);

INVx3_ASAP7_75t_L g171 ( 
.A(n_117),
.Y(n_171)
);

INVx4_ASAP7_75t_L g196 ( 
.A(n_171),
.Y(n_196)
);

INVx3_ASAP7_75t_L g172 ( 
.A(n_129),
.Y(n_172)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_172),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_128),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_SL g176 ( 
.A1(n_151),
.A2(n_143),
.B1(n_132),
.B2(n_129),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g199 ( 
.A(n_176),
.Y(n_199)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_121),
.Y(n_177)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_177),
.Y(n_205)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_135),
.Y(n_178)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_178),
.Y(n_217)
);

INVx3_ASAP7_75t_L g179 ( 
.A(n_132),
.Y(n_179)
);

INVx5_ASAP7_75t_L g216 ( 
.A(n_179),
.Y(n_216)
);

INVx3_ASAP7_75t_L g180 ( 
.A(n_137),
.Y(n_180)
);

INVxp67_ASAP7_75t_L g206 ( 
.A(n_180),
.Y(n_206)
);

AOI22xp33_ASAP7_75t_L g181 ( 
.A1(n_123),
.A2(n_107),
.B1(n_101),
.B2(n_104),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_127),
.Y(n_182)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_182),
.Y(n_219)
);

OAI22xp33_ASAP7_75t_L g184 ( 
.A1(n_123),
.A2(n_6),
.B1(n_7),
.B2(n_152),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_184),
.A2(n_122),
.B1(n_114),
.B2(n_142),
.Y(n_193)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_119),
.Y(n_185)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_185),
.Y(n_220)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_125),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_186),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_150),
.B(n_6),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_109),
.A2(n_99),
.B1(n_100),
.B2(n_146),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_189),
.A2(n_190),
.B1(n_191),
.B2(n_116),
.Y(n_211)
);

AOI22xp33_ASAP7_75t_L g190 ( 
.A1(n_145),
.A2(n_143),
.B1(n_146),
.B2(n_100),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_133),
.B(n_140),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g241 ( 
.A1(n_193),
.A2(n_170),
.B1(n_178),
.B2(n_154),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_158),
.A2(n_114),
.B1(n_142),
.B2(n_151),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_202),
.A2(n_169),
.B1(n_171),
.B2(n_118),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_156),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_203),
.B(n_204),
.Y(n_229)
);

CKINVDCx16_ASAP7_75t_R g204 ( 
.A(n_168),
.Y(n_204)
);

INVx8_ASAP7_75t_L g209 ( 
.A(n_170),
.Y(n_209)
);

INVx3_ASAP7_75t_L g243 ( 
.A(n_209),
.Y(n_243)
);

INVxp67_ASAP7_75t_L g233 ( 
.A(n_211),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_SL g245 ( 
.A1(n_212),
.A2(n_179),
.B(n_180),
.Y(n_245)
);

CKINVDCx16_ASAP7_75t_R g228 ( 
.A(n_213),
.Y(n_228)
);

O2A1O1Ixp33_ASAP7_75t_L g218 ( 
.A1(n_175),
.A2(n_136),
.B(n_110),
.C(n_116),
.Y(n_218)
);

AOI21xp5_ASAP7_75t_L g244 ( 
.A1(n_218),
.A2(n_184),
.B(n_172),
.Y(n_244)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_221),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_214),
.B(n_183),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_222),
.B(n_224),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_215),
.A2(n_195),
.B1(n_213),
.B2(n_166),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_223),
.A2(n_241),
.B1(n_193),
.B2(n_197),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_198),
.B(n_161),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_198),
.B(n_163),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_225),
.B(n_231),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_212),
.B(n_159),
.C(n_191),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_226),
.B(n_234),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_216),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_230),
.B(n_235),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_194),
.B(n_174),
.Y(n_231)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_192),
.Y(n_232)
);

INVx2_ASAP7_75t_SL g254 ( 
.A(n_232),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_202),
.B(n_182),
.C(n_153),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_216),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_194),
.B(n_187),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_236),
.B(n_238),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_237),
.A2(n_199),
.B1(n_192),
.B2(n_196),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_217),
.B(n_161),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_219),
.B(n_155),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_239),
.B(n_242),
.Y(n_265)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_192),
.Y(n_240)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_240),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_201),
.B(n_205),
.Y(n_242)
);

OAI21xp5_ASAP7_75t_SL g266 ( 
.A1(n_244),
.A2(n_245),
.B(n_206),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_247),
.A2(n_253),
.B1(n_260),
.B2(n_244),
.Y(n_269)
);

CKINVDCx16_ASAP7_75t_R g248 ( 
.A(n_242),
.Y(n_248)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_248),
.Y(n_270)
);

A2O1A1Ixp33_ASAP7_75t_SL g249 ( 
.A1(n_228),
.A2(n_197),
.B(n_218),
.C(n_167),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_249),
.B(n_257),
.Y(n_273)
);

INVxp67_ASAP7_75t_L g252 ( 
.A(n_229),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_252),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_223),
.A2(n_199),
.B1(n_217),
.B2(n_205),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_256),
.A2(n_267),
.B1(n_227),
.B2(n_240),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_241),
.Y(n_257)
);

INVxp67_ASAP7_75t_L g258 ( 
.A(n_229),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_258),
.Y(n_281)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_239),
.Y(n_259)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_259),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_228),
.A2(n_219),
.B1(n_210),
.B2(n_185),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_222),
.B(n_201),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_262),
.B(n_224),
.Y(n_274)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_232),
.Y(n_264)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_264),
.Y(n_287)
);

OAI21xp5_ASAP7_75t_SL g271 ( 
.A1(n_266),
.A2(n_245),
.B(n_237),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_233),
.A2(n_196),
.B1(n_210),
.B2(n_220),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_246),
.B(n_226),
.C(n_234),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_268),
.B(n_277),
.C(n_279),
.Y(n_303)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_269),
.Y(n_290)
);

OAI21xp5_ASAP7_75t_L g293 ( 
.A1(n_271),
.A2(n_286),
.B(n_249),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_SL g272 ( 
.A(n_246),
.B(n_226),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g295 ( 
.A(n_272),
.B(n_282),
.Y(n_295)
);

OAI211xp5_ASAP7_75t_L g299 ( 
.A1(n_274),
.A2(n_262),
.B(n_265),
.C(n_259),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_248),
.B(n_225),
.Y(n_275)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_275),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_276),
.A2(n_283),
.B1(n_257),
.B2(n_270),
.Y(n_289)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_246),
.B(n_234),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_256),
.A2(n_227),
.B1(n_238),
.B2(n_236),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_278),
.A2(n_275),
.B1(n_284),
.B2(n_269),
.Y(n_301)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_261),
.B(n_231),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_261),
.B(n_220),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_L g283 ( 
.A1(n_247),
.A2(n_235),
.B1(n_230),
.B2(n_243),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_250),
.B(n_243),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_285),
.B(n_255),
.Y(n_296)
);

NOR2x1_ASAP7_75t_L g286 ( 
.A(n_263),
.B(n_200),
.Y(n_286)
);

AND2x6_ASAP7_75t_L g288 ( 
.A(n_272),
.B(n_273),
.Y(n_288)
);

OAI21xp5_ASAP7_75t_SL g312 ( 
.A1(n_288),
.A2(n_299),
.B(n_305),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g319 ( 
.A1(n_289),
.A2(n_301),
.B1(n_302),
.B2(n_276),
.Y(n_319)
);

FAx1_ASAP7_75t_SL g291 ( 
.A(n_268),
.B(n_250),
.CI(n_263),
.CON(n_291),
.SN(n_291)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_291),
.B(n_293),
.Y(n_316)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_287),
.Y(n_294)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_294),
.Y(n_310)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_296),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_280),
.B(n_264),
.Y(n_297)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_297),
.Y(n_318)
);

CKINVDCx16_ASAP7_75t_R g298 ( 
.A(n_285),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_298),
.B(n_306),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_280),
.B(n_265),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_SL g314 ( 
.A(n_300),
.B(n_304),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_273),
.A2(n_266),
.B1(n_249),
.B2(n_267),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_281),
.B(n_208),
.Y(n_304)
);

AOI21xp5_ASAP7_75t_L g305 ( 
.A1(n_271),
.A2(n_253),
.B(n_255),
.Y(n_305)
);

INVxp67_ASAP7_75t_L g306 ( 
.A(n_287),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_303),
.B(n_272),
.C(n_277),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_307),
.B(n_311),
.C(n_321),
.Y(n_331)
);

XOR2xp5_ASAP7_75t_L g309 ( 
.A(n_303),
.B(n_279),
.Y(n_309)
);

XOR2xp5_ASAP7_75t_L g325 ( 
.A(n_309),
.B(n_313),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_295),
.B(n_284),
.C(n_282),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_295),
.B(n_278),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_301),
.B(n_274),
.Y(n_315)
);

XOR2xp5_ASAP7_75t_L g333 ( 
.A(n_315),
.B(n_320),
.Y(n_333)
);

OAI22xp5_ASAP7_75t_SL g324 ( 
.A1(n_319),
.A2(n_290),
.B1(n_289),
.B2(n_298),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_292),
.B(n_270),
.Y(n_320)
);

XOR2xp5_ASAP7_75t_L g321 ( 
.A(n_292),
.B(n_286),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_297),
.B(n_281),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_322),
.B(n_286),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_308),
.B(n_306),
.Y(n_323)
);

OAI22xp5_ASAP7_75t_L g336 ( 
.A1(n_323),
.A2(n_329),
.B1(n_330),
.B2(n_334),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_L g339 ( 
.A1(n_324),
.A2(n_326),
.B1(n_327),
.B2(n_316),
.Y(n_339)
);

OAI22xp5_ASAP7_75t_SL g326 ( 
.A1(n_319),
.A2(n_290),
.B1(n_293),
.B2(n_305),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_SL g327 ( 
.A1(n_317),
.A2(n_296),
.B1(n_291),
.B2(n_288),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_SL g328 ( 
.A(n_312),
.B(n_251),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_SL g337 ( 
.A(n_328),
.B(n_332),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_320),
.B(n_294),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_SL g332 ( 
.A(n_309),
.B(n_251),
.Y(n_332)
);

AOI21xp5_ASAP7_75t_SL g334 ( 
.A1(n_321),
.A2(n_302),
.B(n_291),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_307),
.B(n_283),
.C(n_260),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_SL g343 ( 
.A(n_335),
.B(n_254),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_331),
.B(n_313),
.C(n_311),
.Y(n_338)
);

OR2x2_ASAP7_75t_L g350 ( 
.A(n_338),
.B(n_340),
.Y(n_350)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_339),
.Y(n_349)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_331),
.B(n_315),
.C(n_318),
.Y(n_340)
);

OAI22xp5_ASAP7_75t_SL g341 ( 
.A1(n_334),
.A2(n_314),
.B1(n_310),
.B2(n_249),
.Y(n_341)
);

HB1xp67_ASAP7_75t_L g348 ( 
.A(n_341),
.Y(n_348)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_325),
.B(n_254),
.C(n_243),
.Y(n_342)
);

OR2x2_ASAP7_75t_L g351 ( 
.A(n_342),
.B(n_343),
.Y(n_351)
);

OAI22xp5_ASAP7_75t_SL g344 ( 
.A1(n_323),
.A2(n_249),
.B1(n_254),
.B2(n_206),
.Y(n_344)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_344),
.Y(n_355)
);

NOR2x1_ASAP7_75t_SL g345 ( 
.A(n_327),
.B(n_249),
.Y(n_345)
);

AOI21xp5_ASAP7_75t_SL g353 ( 
.A1(n_345),
.A2(n_335),
.B(n_326),
.Y(n_353)
);

XOR2xp5_ASAP7_75t_L g346 ( 
.A(n_325),
.B(n_254),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_346),
.B(n_330),
.C(n_333),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_L g347 ( 
.A(n_336),
.B(n_340),
.Y(n_347)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_347),
.Y(n_356)
);

XNOR2xp5_ASAP7_75t_L g363 ( 
.A(n_352),
.B(n_207),
.Y(n_363)
);

OAI21xp5_ASAP7_75t_L g362 ( 
.A1(n_353),
.A2(n_346),
.B(n_208),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_337),
.B(n_324),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_SL g358 ( 
.A(n_354),
.B(n_341),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_350),
.B(n_339),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_357),
.B(n_358),
.Y(n_368)
);

AND2x2_ASAP7_75t_L g359 ( 
.A(n_351),
.B(n_338),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_R g365 ( 
.A(n_359),
.B(n_348),
.Y(n_365)
);

INVxp67_ASAP7_75t_L g360 ( 
.A(n_347),
.Y(n_360)
);

OAI22xp5_ASAP7_75t_SL g369 ( 
.A1(n_360),
.A2(n_362),
.B1(n_207),
.B2(n_186),
.Y(n_369)
);

OAI22xp5_ASAP7_75t_SL g361 ( 
.A1(n_349),
.A2(n_344),
.B1(n_333),
.B2(n_342),
.Y(n_361)
);

INVxp67_ASAP7_75t_L g366 ( 
.A(n_361),
.Y(n_366)
);

MAJx2_ASAP7_75t_L g364 ( 
.A(n_363),
.B(n_359),
.C(n_360),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_364),
.B(n_365),
.Y(n_371)
);

AOI21xp5_ASAP7_75t_SL g367 ( 
.A1(n_356),
.A2(n_355),
.B(n_200),
.Y(n_367)
);

AOI21xp5_ASAP7_75t_L g373 ( 
.A1(n_367),
.A2(n_209),
.B(n_126),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_369),
.B(n_106),
.Y(n_372)
);

MAJIxp5_ASAP7_75t_L g370 ( 
.A(n_366),
.B(n_106),
.C(n_137),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_370),
.B(n_372),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_SL g374 ( 
.A(n_373),
.B(n_368),
.Y(n_374)
);

MAJIxp5_ASAP7_75t_L g376 ( 
.A(n_374),
.B(n_371),
.C(n_139),
.Y(n_376)
);

MAJIxp5_ASAP7_75t_L g377 ( 
.A(n_376),
.B(n_375),
.C(n_126),
.Y(n_377)
);

XOR2xp5_ASAP7_75t_L g378 ( 
.A(n_377),
.B(n_139),
.Y(n_378)
);


endmodule