module fake_jpeg_2826_n_242 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_242);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_242;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_182;
wire n_19;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_140;
wire n_82;
wire n_128;
wire n_100;
wire n_96;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_6),
.Y(n_17)
);

INVx11_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

BUFx2_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_6),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

BUFx16f_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_0),
.Y(n_35)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_11),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_16),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_12),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_27),
.B(n_0),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_39),
.B(n_41),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_19),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_40),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_37),
.B(n_15),
.Y(n_41)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_28),
.Y(n_42)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_42),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_28),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_43),
.B(n_55),
.Y(n_98)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_20),
.Y(n_44)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_44),
.Y(n_64)
);

BUFx16f_ASAP7_75t_L g45 ( 
.A(n_28),
.Y(n_45)
);

BUFx4f_ASAP7_75t_SL g96 ( 
.A(n_45),
.Y(n_96)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_18),
.Y(n_46)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_46),
.Y(n_66)
);

INVx11_ASAP7_75t_L g47 ( 
.A(n_28),
.Y(n_47)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_47),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_19),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_48),
.Y(n_69)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_27),
.Y(n_49)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_49),
.Y(n_86)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_22),
.Y(n_50)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_50),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_34),
.B(n_0),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_51),
.B(n_57),
.Y(n_76)
);

INVx11_ASAP7_75t_L g52 ( 
.A(n_18),
.Y(n_52)
);

INVx5_ASAP7_75t_SL g88 ( 
.A(n_52),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g53 ( 
.A(n_37),
.B(n_15),
.Y(n_53)
);

OR2x2_ASAP7_75t_L g81 ( 
.A(n_53),
.B(n_38),
.Y(n_81)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_22),
.Y(n_54)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_54),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_22),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_34),
.Y(n_56)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_56),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_32),
.Y(n_57)
);

OR2x2_ASAP7_75t_L g58 ( 
.A(n_26),
.B(n_1),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_58),
.B(n_23),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_19),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_59),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_26),
.B(n_12),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_60),
.B(n_61),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_30),
.B(n_1),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_24),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_62),
.Y(n_78)
);

BUFx24_ASAP7_75t_L g63 ( 
.A(n_18),
.Y(n_63)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_63),
.Y(n_95)
);

CKINVDCx12_ASAP7_75t_R g65 ( 
.A(n_45),
.Y(n_65)
);

CKINVDCx14_ASAP7_75t_R g111 ( 
.A(n_65),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_51),
.A2(n_33),
.B1(n_25),
.B2(n_31),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_68),
.A2(n_72),
.B1(n_85),
.B2(n_97),
.Y(n_109)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_45),
.Y(n_70)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_70),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_71),
.B(n_81),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_55),
.A2(n_47),
.B1(n_57),
.B2(n_43),
.Y(n_72)
);

INVx6_ASAP7_75t_SL g77 ( 
.A(n_42),
.Y(n_77)
);

CKINVDCx16_ASAP7_75t_R g123 ( 
.A(n_77),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_40),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_82),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_39),
.B(n_38),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_83),
.B(n_20),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_58),
.A2(n_33),
.B1(n_25),
.B2(n_32),
.Y(n_85)
);

AND2x2_ASAP7_75t_SL g87 ( 
.A(n_56),
.B(n_31),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_87),
.B(n_63),
.C(n_36),
.Y(n_124)
);

OAI21xp33_ASAP7_75t_L g89 ( 
.A1(n_44),
.A2(n_21),
.B(n_35),
.Y(n_89)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_89),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_49),
.A2(n_31),
.B1(n_25),
.B2(n_33),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_92),
.A2(n_24),
.B1(n_54),
.B2(n_50),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_53),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_93),
.B(n_99),
.Y(n_100)
);

INVx6_ASAP7_75t_L g94 ( 
.A(n_48),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_94),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_59),
.A2(n_32),
.B1(n_24),
.B2(n_17),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_62),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_79),
.B(n_30),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_101),
.B(n_110),
.Y(n_131)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_64),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_102),
.B(n_106),
.Y(n_136)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_90),
.Y(n_105)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_105),
.Y(n_152)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_98),
.Y(n_106)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_75),
.Y(n_107)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_107),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_81),
.B(n_21),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_71),
.A2(n_23),
.B1(n_17),
.B2(n_35),
.Y(n_114)
);

CKINVDCx14_ASAP7_75t_R g142 ( 
.A(n_114),
.Y(n_142)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_86),
.Y(n_115)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_115),
.Y(n_132)
);

INVx8_ASAP7_75t_L g116 ( 
.A(n_67),
.Y(n_116)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_116),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_67),
.Y(n_117)
);

INVx8_ASAP7_75t_L g143 ( 
.A(n_117),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_SL g139 ( 
.A(n_118),
.B(n_126),
.Y(n_139)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_80),
.Y(n_119)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_119),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_120),
.A2(n_78),
.B1(n_69),
.B2(n_74),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_95),
.A2(n_29),
.B1(n_46),
.B2(n_52),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_121),
.B(n_88),
.Y(n_137)
);

OAI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_76),
.A2(n_29),
.B1(n_63),
.B2(n_36),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_L g135 ( 
.A1(n_122),
.A2(n_95),
.B1(n_96),
.B2(n_91),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_124),
.B(n_87),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_89),
.B(n_1),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_125),
.B(n_113),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_73),
.B(n_2),
.Y(n_126)
);

BUFx3_ASAP7_75t_L g127 ( 
.A(n_75),
.Y(n_127)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_127),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_69),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_128),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_SL g160 ( 
.A(n_130),
.B(n_147),
.Y(n_160)
);

INVxp33_ASAP7_75t_L g169 ( 
.A(n_135),
.Y(n_169)
);

CKINVDCx16_ASAP7_75t_R g175 ( 
.A(n_137),
.Y(n_175)
);

NAND3xp33_ASAP7_75t_L g172 ( 
.A(n_138),
.B(n_145),
.C(n_131),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_140),
.A2(n_150),
.B1(n_104),
.B2(n_117),
.Y(n_162)
);

OAI32xp33_ASAP7_75t_L g144 ( 
.A1(n_113),
.A2(n_84),
.A3(n_72),
.B1(n_88),
.B2(n_63),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_144),
.B(n_145),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_125),
.B(n_94),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_112),
.B(n_70),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_100),
.B(n_96),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_148),
.B(n_127),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_118),
.B(n_82),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_149),
.B(n_151),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_109),
.A2(n_78),
.B1(n_74),
.B2(n_66),
.Y(n_150)
);

AO22x1_ASAP7_75t_L g151 ( 
.A1(n_120),
.A2(n_91),
.B1(n_66),
.B2(n_96),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_124),
.B(n_2),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_153),
.B(n_2),
.Y(n_171)
);

NOR3xp33_ASAP7_75t_SL g154 ( 
.A(n_139),
.B(n_123),
.C(n_111),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_SL g187 ( 
.A(n_154),
.B(n_166),
.Y(n_187)
);

AOI21xp5_ASAP7_75t_L g156 ( 
.A1(n_130),
.A2(n_107),
.B(n_103),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_SL g191 ( 
.A1(n_156),
.A2(n_174),
.B(n_103),
.Y(n_191)
);

INVx13_ASAP7_75t_L g157 ( 
.A(n_141),
.Y(n_157)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_157),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_149),
.B(n_105),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_159),
.B(n_164),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_138),
.B(n_153),
.C(n_147),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_161),
.B(n_173),
.C(n_129),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_162),
.A2(n_172),
.B1(n_140),
.B2(n_146),
.Y(n_177)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_134),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_163),
.B(n_165),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_139),
.B(n_115),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_136),
.Y(n_165)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_134),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_167),
.B(n_168),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g168 ( 
.A(n_133),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_131),
.B(n_136),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_170),
.B(n_171),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_142),
.B(n_119),
.C(n_132),
.Y(n_173)
);

NOR4xp25_ASAP7_75t_L g174 ( 
.A(n_129),
.B(n_3),
.C(n_4),
.D(n_5),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_177),
.B(n_191),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_155),
.A2(n_150),
.B1(n_144),
.B2(n_151),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_178),
.A2(n_181),
.B1(n_188),
.B2(n_189),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g180 ( 
.A(n_161),
.B(n_132),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_180),
.B(n_182),
.C(n_183),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_155),
.A2(n_146),
.B1(n_133),
.B2(n_143),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_160),
.B(n_152),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_173),
.B(n_152),
.C(n_141),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_186),
.B(n_163),
.C(n_167),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_158),
.A2(n_143),
.B1(n_108),
.B2(n_116),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_158),
.A2(n_151),
.B1(n_143),
.B2(n_108),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_165),
.B(n_104),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_192),
.B(n_128),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_194),
.B(n_197),
.C(n_198),
.Y(n_213)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_185),
.Y(n_196)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_196),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_180),
.B(n_160),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_182),
.B(n_164),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_186),
.B(n_156),
.C(n_159),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_199),
.B(n_201),
.C(n_184),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_183),
.B(n_171),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_178),
.A2(n_175),
.B1(n_162),
.B2(n_169),
.Y(n_202)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_202),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_203),
.B(n_204),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_187),
.B(n_170),
.Y(n_204)
);

AO221x1_ASAP7_75t_L g205 ( 
.A1(n_189),
.A2(n_157),
.B1(n_154),
.B2(n_175),
.C(n_174),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_205),
.B(n_191),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_179),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_206),
.Y(n_212)
);

CKINVDCx16_ASAP7_75t_R g207 ( 
.A(n_200),
.Y(n_207)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_207),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_208),
.A2(n_195),
.B1(n_176),
.B2(n_190),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_209),
.B(n_193),
.Y(n_220)
);

INVx13_ASAP7_75t_L g211 ( 
.A(n_199),
.Y(n_211)
);

AOI21xp5_ASAP7_75t_L g223 ( 
.A1(n_211),
.A2(n_215),
.B(n_201),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_SL g215 ( 
.A1(n_202),
.A2(n_184),
.B(n_176),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_212),
.B(n_207),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_SL g228 ( 
.A(n_217),
.B(n_222),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_L g218 ( 
.A1(n_209),
.A2(n_194),
.B(n_198),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_218),
.B(n_219),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_220),
.B(n_223),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_SL g222 ( 
.A1(n_212),
.A2(n_197),
.B(n_193),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_216),
.A2(n_168),
.B1(n_157),
.B2(n_8),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_224),
.A2(n_214),
.B1(n_208),
.B2(n_216),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_219),
.B(n_213),
.C(n_209),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_225),
.B(n_227),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_221),
.B(n_210),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_229),
.B(n_215),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_232),
.A2(n_230),
.B1(n_213),
.B2(n_224),
.Y(n_235)
);

OAI21xp5_ASAP7_75t_SL g233 ( 
.A1(n_226),
.A2(n_228),
.B(n_225),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_SL g236 ( 
.A(n_233),
.B(n_229),
.Y(n_236)
);

OAI21x1_ASAP7_75t_L g234 ( 
.A1(n_230),
.A2(n_210),
.B(n_214),
.Y(n_234)
);

OAI21x1_ASAP7_75t_L g237 ( 
.A1(n_234),
.A2(n_211),
.B(n_168),
.Y(n_237)
);

MAJx2_ASAP7_75t_L g238 ( 
.A(n_235),
.B(n_237),
.C(n_232),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_L g239 ( 
.A1(n_236),
.A2(n_231),
.B1(n_211),
.B2(n_8),
.Y(n_239)
);

AOI21xp5_ASAP7_75t_SL g240 ( 
.A1(n_238),
.A2(n_239),
.B(n_4),
.Y(n_240)
);

AOI322xp5_ASAP7_75t_L g241 ( 
.A1(n_240),
.A2(n_4),
.A3(n_7),
.B1(n_8),
.B2(n_9),
.C1(n_212),
.C2(n_217),
.Y(n_241)
);

BUFx24_ASAP7_75t_SL g242 ( 
.A(n_241),
.Y(n_242)
);


endmodule