module fake_ariane_3242_n_2045 (n_83, n_8, n_56, n_60, n_170, n_190, n_160, n_64, n_179, n_180, n_119, n_124, n_167, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_176, n_149, n_34, n_158, n_172, n_69, n_95, n_175, n_92, n_143, n_183, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_181, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_174, n_100, n_17, n_50, n_187, n_132, n_62, n_147, n_51, n_166, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_159, n_107, n_189, n_72, n_105, n_128, n_44, n_30, n_82, n_178, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_188, n_185, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_148, n_164, n_52, n_157, n_184, n_177, n_135, n_73, n_77, n_171, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_182, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_191, n_151, n_136, n_192, n_28, n_80, n_146, n_194, n_97, n_154, n_142, n_161, n_14, n_163, n_88, n_186, n_141, n_68, n_116, n_104, n_145, n_78, n_193, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_2045);

input n_83;
input n_8;
input n_56;
input n_60;
input n_170;
input n_190;
input n_160;
input n_64;
input n_179;
input n_180;
input n_119;
input n_124;
input n_167;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_176;
input n_149;
input n_34;
input n_158;
input n_172;
input n_69;
input n_95;
input n_175;
input n_92;
input n_143;
input n_183;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_181;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_174;
input n_100;
input n_17;
input n_50;
input n_187;
input n_132;
input n_62;
input n_147;
input n_51;
input n_166;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_159;
input n_107;
input n_189;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_178;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_188;
input n_185;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_164;
input n_52;
input n_157;
input n_184;
input n_177;
input n_135;
input n_73;
input n_77;
input n_171;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_182;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_191;
input n_151;
input n_136;
input n_192;
input n_28;
input n_80;
input n_146;
input n_194;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_186;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_193;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_2045;

wire n_913;
wire n_1681;
wire n_1486;
wire n_1507;
wire n_1938;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_2030;
wire n_1169;
wire n_789;
wire n_850;
wire n_1916;
wire n_610;
wire n_245;
wire n_1713;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_2002;
wire n_1463;
wire n_1238;
wire n_2011;
wire n_1515;
wire n_817;
wire n_1837;
wire n_924;
wire n_781;
wire n_2013;
wire n_1566;
wire n_717;
wire n_2006;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_524;
wire n_1214;
wire n_634;
wire n_1839;
wire n_1246;
wire n_1138;
wire n_214;
wire n_2042;
wire n_1853;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_1999;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_232;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1835;
wire n_1457;
wire n_377;
wire n_1682;
wire n_1836;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_958;
wire n_945;
wire n_813;
wire n_419;
wire n_1985;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1909;
wire n_1184;
wire n_1961;
wire n_202;
wire n_1535;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1979;
wire n_1277;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_672;
wire n_740;
wire n_1283;
wire n_1974;
wire n_1736;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1888;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_242;
wire n_645;
wire n_1944;
wire n_331;
wire n_559;
wire n_495;
wire n_267;
wire n_1988;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_1936;
wire n_200;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1847;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1851;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_1900;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_1889;
wire n_587;
wire n_1977;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_206;
wire n_352;
wire n_899;
wire n_1703;
wire n_611;
wire n_1295;
wire n_1850;
wire n_238;
wire n_365;
wire n_2004;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_661;
wire n_1751;
wire n_300;
wire n_533;
wire n_1917;
wire n_1924;
wire n_438;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_1811;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_1840;
wire n_376;
wire n_512;
wire n_1597;
wire n_1771;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_237;
wire n_2043;
wire n_780;
wire n_1918;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1949;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_490;
wire n_209;
wire n_1461;
wire n_1391;
wire n_1947;
wire n_225;
wire n_1599;
wire n_1876;
wire n_1006;
wire n_1830;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_2038;
wire n_1838;
wire n_1594;
wire n_680;
wire n_1935;
wire n_287;
wire n_1716;
wire n_302;
wire n_1872;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_212;
wire n_444;
wire n_851;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_1819;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_1833;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_1884;
wire n_460;
wire n_1555;
wire n_1842;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_992;
wire n_966;
wire n_955;
wire n_1182;
wire n_794;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_1292;
wire n_1178;
wire n_1972;
wire n_2015;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_306;
wire n_203;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_437;
wire n_337;
wire n_274;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1787;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_1717;
wire n_1812;
wire n_824;
wire n_428;
wire n_892;
wire n_1880;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_1855;
wire n_990;
wire n_1623;
wire n_1903;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_1932;
wire n_1780;
wire n_1970;
wire n_1920;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1911;
wire n_1825;
wire n_1908;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1832;
wire n_1841;
wire n_1680;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_1731;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_1914;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_2019;
wire n_698;
wire n_1674;
wire n_2021;
wire n_2025;
wire n_1992;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_1913;
wire n_1058;
wire n_347;
wire n_1042;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_205;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_1728;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_2041;
wire n_1933;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_1817;
wire n_348;
wire n_552;
wire n_670;
wire n_1826;
wire n_379;
wire n_264;
wire n_441;
wire n_1951;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_1869;
wire n_1743;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_1943;
wire n_1802;
wire n_1163;
wire n_1795;
wire n_1384;
wire n_1868;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1879;
wire n_1886;
wire n_1648;
wire n_1413;
wire n_855;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_1901;
wire n_647;
wire n_2027;
wire n_1423;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_1939;
wire n_1906;
wire n_529;
wire n_1899;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1828;
wire n_1798;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_1105;
wire n_547;
wire n_439;
wire n_677;
wire n_604;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_2023;
wire n_1278;
wire n_707;
wire n_983;
wire n_727;
wire n_590;
wire n_699;
wire n_301;
wire n_1726;
wire n_1945;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_2031;
wire n_325;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_1963;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1693;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1823;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_2033;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_221;
wire n_321;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1863;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_1859;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_1883;
wire n_1969;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_845;
wire n_888;
wire n_1649;
wire n_1677;
wire n_1927;
wire n_1297;
wire n_551;
wire n_417;
wire n_1708;
wire n_343;
wire n_1222;
wire n_1844;
wire n_582;
wire n_1957;
wire n_1953;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_1919;
wire n_534;
wire n_1791;
wire n_1894;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_1898;
wire n_451;
wire n_745;
wire n_1741;
wire n_1572;
wire n_1907;
wire n_1793;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1975;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_769;
wire n_1797;
wire n_1753;
wire n_1990;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_1895;
wire n_982;
wire n_1800;
wire n_915;
wire n_215;
wire n_1075;
wire n_2008;
wire n_454;
wire n_298;
wire n_1331;
wire n_1890;
wire n_1529;
wire n_1227;
wire n_655;
wire n_1734;
wire n_1860;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_509;
wire n_1854;
wire n_666;
wire n_1747;
wire n_430;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_456;
wire n_1867;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_873;
wire n_1301;
wire n_1748;
wire n_1966;
wire n_1243;
wire n_1400;
wire n_342;
wire n_2035;
wire n_1466;
wire n_1513;
wire n_1527;
wire n_358;
wire n_1783;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1993;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1954;
wire n_1668;
wire n_1878;
wire n_1605;
wire n_1078;
wire n_266;
wire n_1897;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_2026;
wire n_1786;
wire n_480;
wire n_1327;
wire n_1475;
wire n_211;
wire n_642;
wire n_1804;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_1757;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_1632;
wire n_1769;
wire n_474;
wire n_1929;
wire n_1950;
wire n_805;
wire n_2032;
wire n_295;
wire n_1658;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1997;
wire n_1137;
wire n_1873;
wire n_1258;
wire n_197;
wire n_640;
wire n_463;
wire n_1476;
wire n_1524;
wire n_1733;
wire n_1856;
wire n_2016;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1874;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_1807;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_1784;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_283;
wire n_806;
wire n_1984;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_1824;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_1822;
wire n_682;
wire n_1616;
wire n_819;
wire n_1971;
wire n_586;
wire n_1324;
wire n_1429;
wire n_1778;
wire n_1776;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1759;
wire n_1829;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_2022;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_1815;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_198;
wire n_1864;
wire n_1887;
wire n_1208;
wire n_1987;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_1852;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1995;
wire n_1877;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_2001;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_1201;
wire n_1288;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_1367;
wire n_2044;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_420;
wire n_1291;
wire n_562;
wire n_2020;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1882;
wire n_1976;
wire n_1023;
wire n_1881;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_1958;
wire n_467;
wire n_1511;
wire n_1422;
wire n_1965;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_538;
wire n_1517;
wire n_2036;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_2003;
wire n_1307;
wire n_1128;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1921;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1955;
wire n_1773;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_1948;
wire n_810;
wire n_1290;
wire n_1959;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_1960;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_1968;
wire n_1885;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_1978;
wire n_414;
wire n_571;
wire n_1521;
wire n_1694;
wire n_1940;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_409;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_2007;
wire n_526;
wire n_1994;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1973;
wire n_1444;
wire n_1803;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_1739;
wire n_1814;
wire n_532;
wire n_1789;
wire n_763;
wire n_1986;
wire n_540;
wire n_216;
wire n_692;
wire n_1857;
wire n_984;
wire n_1687;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_1910;
wire n_1816;
wire n_1756;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_2018;
wire n_1772;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_2040;
wire n_493;
wire n_1311;
wire n_1956;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1962;
wire n_1335;
wire n_1715;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_1785;
wire n_792;
wire n_1262;
wire n_1942;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_2014;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1893;
wire n_1183;
wire n_1326;
wire n_1805;
wire n_981;
wire n_1110;
wire n_1758;
wire n_243;
wire n_1407;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_2010;
wire n_1054;
wire n_508;
wire n_1679;
wire n_1952;
wire n_1858;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_1834;
wire n_1011;
wire n_978;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_1536;
wire n_1471;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_1980;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_1998;
wire n_541;
wire n_499;
wire n_1775;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_2028;
wire n_919;
wire n_1663;
wire n_1625;
wire n_1926;
wire n_318;
wire n_1458;
wire n_244;
wire n_679;
wire n_1630;
wire n_220;
wire n_663;
wire n_1720;
wire n_443;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_1922;
wire n_1735;
wire n_1788;
wire n_391;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_1930;
wire n_765;
wire n_1809;
wire n_1843;
wire n_1904;
wire n_2000;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_857;
wire n_898;
wire n_363;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1937;
wire n_2012;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_2039;
wire n_1755;
wire n_1285;
wire n_733;
wire n_761;
wire n_731;
wire n_336;
wire n_1813;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1996;
wire n_1106;
wire n_2009;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_2024;
wire n_1348;
wire n_753;
wire n_1770;
wire n_701;
wire n_1003;
wire n_1125;
wire n_1710;
wire n_1865;
wire n_309;
wire n_1344;
wire n_1390;
wire n_401;
wire n_485;
wire n_1792;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_567;
wire n_240;
wire n_369;
wire n_1727;
wire n_1991;
wire n_1575;
wire n_1848;
wire n_1892;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_1902;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_2034;
wire n_1845;
wire n_1934;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1806;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_2005;
wire n_1696;
wire n_498;
wire n_1875;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1831;
wire n_1497;
wire n_1866;
wire n_459;
wire n_1136;
wire n_1782;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1941;
wire n_1316;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_1915;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_1781;
wire n_709;
wire n_809;
wire n_1686;
wire n_1964;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_1982;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_199;
wire n_217;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_308;
wire n_1223;
wire n_201;
wire n_1768;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1983;
wire n_1041;
wire n_993;
wire n_1862;
wire n_948;
wire n_2017;
wire n_922;
wire n_1004;
wire n_1810;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_1923;
wire n_1764;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_196;
wire n_1337;
wire n_774;
wire n_1946;
wire n_933;
wire n_1779;
wire n_596;
wire n_954;
wire n_1168;
wire n_1821;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_252;
wire n_664;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1896;
wire n_1732;
wire n_415;
wire n_1967;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1799;
wire n_1126;
wire n_2029;
wire n_195;
wire n_1846;
wire n_1912;
wire n_938;
wire n_1891;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_1928;
wire n_946;
wire n_757;
wire n_375;
wire n_1655;
wire n_1818;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_265;
wire n_1583;
wire n_1604;
wire n_208;
wire n_1631;
wire n_1702;
wire n_275;
wire n_1794;
wire n_1375;
wire n_204;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_1827;
wire n_866;
wire n_246;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_1871;
wire n_718;
wire n_329;
wire n_1434;
wire n_340;
wire n_1905;
wire n_1569;
wire n_289;
wire n_548;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_1870;
wire n_1925;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1861;
wire n_1228;
wire n_1931;
wire n_1244;
wire n_1796;
wire n_411;
wire n_484;
wire n_849;
wire n_1820;
wire n_357;
wire n_412;
wire n_1251;
wire n_1989;
wire n_447;
wire n_1421;
wire n_1762;
wire n_1233;
wire n_1808;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_1981;
wire n_2037;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_106),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_151),
.Y(n_196)
);

INVx1_ASAP7_75t_SL g197 ( 
.A(n_15),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_100),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_52),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_55),
.Y(n_200)
);

INVx1_ASAP7_75t_SL g201 ( 
.A(n_162),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_189),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_39),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_187),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_3),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_20),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_129),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_169),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_194),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_136),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_61),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_51),
.Y(n_212)
);

INVx2_ASAP7_75t_SL g213 ( 
.A(n_1),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_68),
.Y(n_214)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_130),
.Y(n_215)
);

INVx2_ASAP7_75t_SL g216 ( 
.A(n_8),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_57),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_29),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_48),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_51),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_105),
.Y(n_221)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_88),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_103),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_95),
.Y(n_224)
);

CKINVDCx14_ASAP7_75t_R g225 ( 
.A(n_86),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_44),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_58),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_74),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_147),
.Y(n_229)
);

INVx1_ASAP7_75t_SL g230 ( 
.A(n_145),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_76),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_92),
.Y(n_232)
);

INVx2_ASAP7_75t_SL g233 ( 
.A(n_24),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_188),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_178),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_159),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_30),
.Y(n_237)
);

BUFx3_ASAP7_75t_L g238 ( 
.A(n_53),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_141),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_112),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_191),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_37),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_185),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_80),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_34),
.Y(n_245)
);

BUFx10_ASAP7_75t_L g246 ( 
.A(n_23),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_78),
.Y(n_247)
);

BUFx10_ASAP7_75t_L g248 ( 
.A(n_168),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_146),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_98),
.Y(n_250)
);

BUFx6f_ASAP7_75t_L g251 ( 
.A(n_163),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_75),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_24),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_37),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_82),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_21),
.Y(n_256)
);

BUFx3_ASAP7_75t_L g257 ( 
.A(n_22),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_96),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_131),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_72),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_167),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_13),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_184),
.Y(n_263)
);

INVx1_ASAP7_75t_SL g264 ( 
.A(n_109),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_124),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_125),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_1),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_121),
.Y(n_268)
);

BUFx3_ASAP7_75t_L g269 ( 
.A(n_128),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_36),
.Y(n_270)
);

BUFx10_ASAP7_75t_L g271 ( 
.A(n_36),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_71),
.Y(n_272)
);

BUFx8_ASAP7_75t_SL g273 ( 
.A(n_31),
.Y(n_273)
);

INVx1_ASAP7_75t_SL g274 ( 
.A(n_79),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_165),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_74),
.Y(n_276)
);

BUFx10_ASAP7_75t_L g277 ( 
.A(n_85),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_70),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_148),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_160),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_157),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_16),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_83),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_154),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_75),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_2),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_39),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_52),
.Y(n_288)
);

CKINVDCx14_ASAP7_75t_R g289 ( 
.A(n_65),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_20),
.Y(n_290)
);

BUFx10_ASAP7_75t_L g291 ( 
.A(n_192),
.Y(n_291)
);

BUFx10_ASAP7_75t_L g292 ( 
.A(n_108),
.Y(n_292)
);

BUFx2_ASAP7_75t_L g293 ( 
.A(n_114),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_110),
.Y(n_294)
);

INVx1_ASAP7_75t_SL g295 ( 
.A(n_152),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_107),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_71),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_7),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_61),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_186),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_150),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_155),
.Y(n_302)
);

BUFx3_ASAP7_75t_L g303 ( 
.A(n_180),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_31),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_183),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_134),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_97),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_93),
.Y(n_308)
);

INVx2_ASAP7_75t_SL g309 ( 
.A(n_12),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_119),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_78),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_70),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_54),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_111),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_46),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_28),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_120),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_22),
.Y(n_318)
);

CKINVDCx14_ASAP7_75t_R g319 ( 
.A(n_84),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_135),
.Y(n_320)
);

BUFx6f_ASAP7_75t_L g321 ( 
.A(n_91),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_15),
.Y(n_322)
);

BUFx3_ASAP7_75t_L g323 ( 
.A(n_3),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_77),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_0),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_176),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_72),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_161),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_32),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g330 ( 
.A(n_122),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_174),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_144),
.Y(n_332)
);

BUFx3_ASAP7_75t_L g333 ( 
.A(n_153),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_99),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_132),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_41),
.Y(n_336)
);

BUFx10_ASAP7_75t_L g337 ( 
.A(n_21),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_65),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_9),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_127),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_149),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_182),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_177),
.Y(n_343)
);

BUFx8_ASAP7_75t_SL g344 ( 
.A(n_116),
.Y(n_344)
);

INVx2_ASAP7_75t_SL g345 ( 
.A(n_6),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_140),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_59),
.Y(n_347)
);

BUFx6f_ASAP7_75t_L g348 ( 
.A(n_62),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_19),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_17),
.Y(n_350)
);

INVx2_ASAP7_75t_L g351 ( 
.A(n_60),
.Y(n_351)
);

INVx1_ASAP7_75t_SL g352 ( 
.A(n_29),
.Y(n_352)
);

INVx2_ASAP7_75t_L g353 ( 
.A(n_133),
.Y(n_353)
);

BUFx3_ASAP7_75t_L g354 ( 
.A(n_8),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_172),
.Y(n_355)
);

INVx2_ASAP7_75t_SL g356 ( 
.A(n_181),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_104),
.Y(n_357)
);

INVx2_ASAP7_75t_L g358 ( 
.A(n_118),
.Y(n_358)
);

CKINVDCx16_ASAP7_75t_R g359 ( 
.A(n_90),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_58),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_23),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_35),
.Y(n_362)
);

INVx2_ASAP7_75t_SL g363 ( 
.A(n_32),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_190),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_50),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_101),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_94),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_171),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_47),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_102),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_59),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_53),
.Y(n_372)
);

BUFx3_ASAP7_75t_L g373 ( 
.A(n_7),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_139),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_64),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_13),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_16),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_156),
.Y(n_378)
);

INVx2_ASAP7_75t_L g379 ( 
.A(n_10),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_166),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_28),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_43),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_57),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_0),
.Y(n_384)
);

INVx1_ASAP7_75t_SL g385 ( 
.A(n_46),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_193),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_87),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_113),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_48),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_175),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_64),
.Y(n_391)
);

CKINVDCx20_ASAP7_75t_R g392 ( 
.A(n_170),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_68),
.Y(n_393)
);

BUFx3_ASAP7_75t_L g394 ( 
.A(n_12),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_89),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_196),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_196),
.Y(n_397)
);

INVx2_ASAP7_75t_L g398 ( 
.A(n_348),
.Y(n_398)
);

HB1xp67_ASAP7_75t_L g399 ( 
.A(n_289),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_273),
.Y(n_400)
);

INVx1_ASAP7_75t_SL g401 ( 
.A(n_214),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_198),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_198),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_207),
.Y(n_404)
);

INVxp67_ASAP7_75t_SL g405 ( 
.A(n_238),
.Y(n_405)
);

CKINVDCx20_ASAP7_75t_R g406 ( 
.A(n_224),
.Y(n_406)
);

INVxp67_ASAP7_75t_L g407 ( 
.A(n_199),
.Y(n_407)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_348),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_207),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_208),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_208),
.Y(n_411)
);

INVxp33_ASAP7_75t_SL g412 ( 
.A(n_200),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_234),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_234),
.Y(n_414)
);

BUFx3_ASAP7_75t_L g415 ( 
.A(n_293),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_344),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_305),
.Y(n_417)
);

CKINVDCx20_ASAP7_75t_R g418 ( 
.A(n_320),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_236),
.Y(n_419)
);

INVxp67_ASAP7_75t_SL g420 ( 
.A(n_257),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_330),
.Y(n_421)
);

BUFx6f_ASAP7_75t_L g422 ( 
.A(n_251),
.Y(n_422)
);

INVxp67_ASAP7_75t_SL g423 ( 
.A(n_257),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_236),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_240),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_240),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_241),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_241),
.Y(n_428)
);

CKINVDCx20_ASAP7_75t_R g429 ( 
.A(n_340),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_244),
.Y(n_430)
);

CKINVDCx20_ASAP7_75t_R g431 ( 
.A(n_392),
.Y(n_431)
);

CKINVDCx20_ASAP7_75t_R g432 ( 
.A(n_260),
.Y(n_432)
);

INVxp67_ASAP7_75t_L g433 ( 
.A(n_199),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_244),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_255),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_255),
.Y(n_436)
);

CKINVDCx20_ASAP7_75t_R g437 ( 
.A(n_293),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_266),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_203),
.Y(n_439)
);

HB1xp67_ASAP7_75t_L g440 ( 
.A(n_323),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_266),
.Y(n_441)
);

CKINVDCx16_ASAP7_75t_R g442 ( 
.A(n_359),
.Y(n_442)
);

INVxp67_ASAP7_75t_SL g443 ( 
.A(n_354),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_279),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_279),
.Y(n_445)
);

BUFx3_ASAP7_75t_L g446 ( 
.A(n_269),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_205),
.Y(n_447)
);

INVxp67_ASAP7_75t_SL g448 ( 
.A(n_354),
.Y(n_448)
);

INVx2_ASAP7_75t_L g449 ( 
.A(n_348),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_283),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_283),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_296),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_206),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_211),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_296),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_300),
.Y(n_456)
);

BUFx2_ASAP7_75t_SL g457 ( 
.A(n_248),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_300),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_219),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_301),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_301),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_306),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_237),
.Y(n_463)
);

INVxp33_ASAP7_75t_SL g464 ( 
.A(n_245),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_306),
.Y(n_465)
);

BUFx2_ASAP7_75t_L g466 ( 
.A(n_373),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_307),
.Y(n_467)
);

CKINVDCx5p33_ASAP7_75t_R g468 ( 
.A(n_247),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_307),
.Y(n_469)
);

CKINVDCx5p33_ASAP7_75t_R g470 ( 
.A(n_252),
.Y(n_470)
);

CKINVDCx5p33_ASAP7_75t_R g471 ( 
.A(n_253),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_308),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_308),
.Y(n_473)
);

CKINVDCx16_ASAP7_75t_R g474 ( 
.A(n_225),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_326),
.Y(n_475)
);

CKINVDCx20_ASAP7_75t_R g476 ( 
.A(n_319),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_326),
.Y(n_477)
);

CKINVDCx20_ASAP7_75t_R g478 ( 
.A(n_248),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_331),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_331),
.Y(n_480)
);

INVxp67_ASAP7_75t_L g481 ( 
.A(n_212),
.Y(n_481)
);

INVx2_ASAP7_75t_L g482 ( 
.A(n_348),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_346),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_346),
.Y(n_484)
);

INVxp67_ASAP7_75t_L g485 ( 
.A(n_212),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_355),
.Y(n_486)
);

INVxp33_ASAP7_75t_SL g487 ( 
.A(n_262),
.Y(n_487)
);

CKINVDCx16_ASAP7_75t_R g488 ( 
.A(n_246),
.Y(n_488)
);

CKINVDCx5p33_ASAP7_75t_R g489 ( 
.A(n_272),
.Y(n_489)
);

INVx2_ASAP7_75t_L g490 ( 
.A(n_348),
.Y(n_490)
);

INVxp67_ASAP7_75t_SL g491 ( 
.A(n_373),
.Y(n_491)
);

CKINVDCx16_ASAP7_75t_R g492 ( 
.A(n_246),
.Y(n_492)
);

CKINVDCx20_ASAP7_75t_R g493 ( 
.A(n_248),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_355),
.Y(n_494)
);

INVxp67_ASAP7_75t_SL g495 ( 
.A(n_394),
.Y(n_495)
);

BUFx2_ASAP7_75t_L g496 ( 
.A(n_394),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_357),
.Y(n_497)
);

CKINVDCx5p33_ASAP7_75t_R g498 ( 
.A(n_276),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_357),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_364),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_364),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_367),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_367),
.Y(n_503)
);

AND2x4_ASAP7_75t_L g504 ( 
.A(n_446),
.B(n_213),
.Y(n_504)
);

INVx2_ASAP7_75t_L g505 ( 
.A(n_398),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_SL g506 ( 
.A(n_474),
.B(n_248),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_398),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_408),
.Y(n_508)
);

AND2x4_ASAP7_75t_L g509 ( 
.A(n_446),
.B(n_213),
.Y(n_509)
);

CKINVDCx20_ASAP7_75t_R g510 ( 
.A(n_432),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_408),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_449),
.Y(n_512)
);

INVx2_ASAP7_75t_L g513 ( 
.A(n_449),
.Y(n_513)
);

BUFx6f_ASAP7_75t_L g514 ( 
.A(n_422),
.Y(n_514)
);

INVx3_ASAP7_75t_L g515 ( 
.A(n_482),
.Y(n_515)
);

AND2x2_ASAP7_75t_L g516 ( 
.A(n_466),
.B(n_246),
.Y(n_516)
);

NOR2xp33_ASAP7_75t_L g517 ( 
.A(n_457),
.B(n_370),
.Y(n_517)
);

CKINVDCx5p33_ASAP7_75t_R g518 ( 
.A(n_417),
.Y(n_518)
);

OAI22xp5_ASAP7_75t_SL g519 ( 
.A1(n_437),
.A2(n_197),
.B1(n_352),
.B2(n_274),
.Y(n_519)
);

CKINVDCx5p33_ASAP7_75t_R g520 ( 
.A(n_421),
.Y(n_520)
);

AND2x2_ASAP7_75t_L g521 ( 
.A(n_466),
.B(n_246),
.Y(n_521)
);

BUFx2_ASAP7_75t_L g522 ( 
.A(n_439),
.Y(n_522)
);

BUFx6f_ASAP7_75t_L g523 ( 
.A(n_422),
.Y(n_523)
);

INVx2_ASAP7_75t_L g524 ( 
.A(n_422),
.Y(n_524)
);

INVx3_ASAP7_75t_L g525 ( 
.A(n_482),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_457),
.B(n_370),
.Y(n_526)
);

CKINVDCx5p33_ASAP7_75t_R g527 ( 
.A(n_416),
.Y(n_527)
);

INVx2_ASAP7_75t_L g528 ( 
.A(n_490),
.Y(n_528)
);

AND2x2_ASAP7_75t_L g529 ( 
.A(n_496),
.B(n_271),
.Y(n_529)
);

HB1xp67_ASAP7_75t_L g530 ( 
.A(n_447),
.Y(n_530)
);

BUFx6f_ASAP7_75t_L g531 ( 
.A(n_422),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_490),
.Y(n_532)
);

BUFx6f_ASAP7_75t_L g533 ( 
.A(n_422),
.Y(n_533)
);

OAI22xp5_ASAP7_75t_SL g534 ( 
.A1(n_406),
.A2(n_385),
.B1(n_218),
.B2(n_220),
.Y(n_534)
);

AOI22xp5_ASAP7_75t_L g535 ( 
.A1(n_478),
.A2(n_233),
.B1(n_309),
.B2(n_216),
.Y(n_535)
);

AOI22xp5_ASAP7_75t_L g536 ( 
.A1(n_493),
.A2(n_233),
.B1(n_309),
.B2(n_216),
.Y(n_536)
);

BUFx2_ASAP7_75t_L g537 ( 
.A(n_453),
.Y(n_537)
);

BUFx8_ASAP7_75t_L g538 ( 
.A(n_496),
.Y(n_538)
);

AND2x2_ASAP7_75t_L g539 ( 
.A(n_405),
.B(n_420),
.Y(n_539)
);

CKINVDCx20_ASAP7_75t_R g540 ( 
.A(n_418),
.Y(n_540)
);

CKINVDCx16_ASAP7_75t_R g541 ( 
.A(n_488),
.Y(n_541)
);

INVxp67_ASAP7_75t_L g542 ( 
.A(n_399),
.Y(n_542)
);

HB1xp67_ASAP7_75t_L g543 ( 
.A(n_454),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_396),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_396),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_397),
.Y(n_546)
);

NOR2xp33_ASAP7_75t_L g547 ( 
.A(n_474),
.B(n_386),
.Y(n_547)
);

BUFx2_ASAP7_75t_L g548 ( 
.A(n_459),
.Y(n_548)
);

INVx2_ASAP7_75t_L g549 ( 
.A(n_397),
.Y(n_549)
);

INVx3_ASAP7_75t_L g550 ( 
.A(n_402),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_402),
.Y(n_551)
);

BUFx6f_ASAP7_75t_L g552 ( 
.A(n_403),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_403),
.Y(n_553)
);

HB1xp67_ASAP7_75t_L g554 ( 
.A(n_463),
.Y(n_554)
);

INVx2_ASAP7_75t_L g555 ( 
.A(n_404),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_L g556 ( 
.A(n_423),
.B(n_386),
.Y(n_556)
);

INVx2_ASAP7_75t_L g557 ( 
.A(n_404),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_SL g558 ( 
.A(n_442),
.B(n_277),
.Y(n_558)
);

INVx2_ASAP7_75t_L g559 ( 
.A(n_409),
.Y(n_559)
);

CKINVDCx16_ASAP7_75t_R g560 ( 
.A(n_492),
.Y(n_560)
);

INVx2_ASAP7_75t_L g561 ( 
.A(n_409),
.Y(n_561)
);

OAI22xp5_ASAP7_75t_SL g562 ( 
.A1(n_429),
.A2(n_217),
.B1(n_220),
.B2(n_218),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_410),
.Y(n_563)
);

CKINVDCx20_ASAP7_75t_R g564 ( 
.A(n_431),
.Y(n_564)
);

OAI22xp5_ASAP7_75t_SL g565 ( 
.A1(n_401),
.A2(n_217),
.B1(n_227),
.B2(n_226),
.Y(n_565)
);

OAI22xp5_ASAP7_75t_L g566 ( 
.A1(n_415),
.A2(n_363),
.B1(n_345),
.B2(n_286),
.Y(n_566)
);

AND2x4_ASAP7_75t_L g567 ( 
.A(n_410),
.B(n_345),
.Y(n_567)
);

BUFx6f_ASAP7_75t_L g568 ( 
.A(n_411),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_411),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_413),
.Y(n_570)
);

NOR2xp33_ASAP7_75t_L g571 ( 
.A(n_412),
.B(n_388),
.Y(n_571)
);

CKINVDCx5p33_ASAP7_75t_R g572 ( 
.A(n_400),
.Y(n_572)
);

NAND2xp33_ASAP7_75t_L g573 ( 
.A(n_468),
.B(n_363),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_413),
.Y(n_574)
);

INVx2_ASAP7_75t_SL g575 ( 
.A(n_470),
.Y(n_575)
);

CKINVDCx20_ASAP7_75t_R g576 ( 
.A(n_476),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_414),
.Y(n_577)
);

BUFx6f_ASAP7_75t_L g578 ( 
.A(n_414),
.Y(n_578)
);

AND2x2_ASAP7_75t_SL g579 ( 
.A(n_419),
.B(n_215),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_419),
.Y(n_580)
);

INVx2_ASAP7_75t_L g581 ( 
.A(n_424),
.Y(n_581)
);

AOI22xp5_ASAP7_75t_L g582 ( 
.A1(n_415),
.A2(n_278),
.B1(n_297),
.B2(n_288),
.Y(n_582)
);

BUFx3_ASAP7_75t_L g583 ( 
.A(n_424),
.Y(n_583)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_425),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_425),
.Y(n_585)
);

CKINVDCx5p33_ASAP7_75t_R g586 ( 
.A(n_471),
.Y(n_586)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_426),
.Y(n_587)
);

INVx2_ASAP7_75t_SL g588 ( 
.A(n_579),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_552),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_552),
.Y(n_590)
);

INVx2_ASAP7_75t_L g591 ( 
.A(n_505),
.Y(n_591)
);

INVx2_ASAP7_75t_L g592 ( 
.A(n_505),
.Y(n_592)
);

NOR2xp33_ASAP7_75t_L g593 ( 
.A(n_547),
.B(n_464),
.Y(n_593)
);

INVx2_ASAP7_75t_SL g594 ( 
.A(n_579),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_L g595 ( 
.A(n_517),
.B(n_426),
.Y(n_595)
);

INVx3_ASAP7_75t_L g596 ( 
.A(n_552),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_SL g597 ( 
.A(n_575),
.B(n_489),
.Y(n_597)
);

AOI22xp33_ASAP7_75t_SL g598 ( 
.A1(n_562),
.A2(n_487),
.B1(n_337),
.B2(n_271),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_552),
.Y(n_599)
);

INVx2_ASAP7_75t_L g600 ( 
.A(n_513),
.Y(n_600)
);

NOR2xp33_ASAP7_75t_L g601 ( 
.A(n_526),
.B(n_498),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_528),
.Y(n_602)
);

AND2x2_ASAP7_75t_L g603 ( 
.A(n_539),
.B(n_443),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_552),
.Y(n_604)
);

INVx2_ASAP7_75t_L g605 ( 
.A(n_528),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_552),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_L g607 ( 
.A(n_579),
.B(n_427),
.Y(n_607)
);

INVx8_ASAP7_75t_L g608 ( 
.A(n_539),
.Y(n_608)
);

INVx4_ASAP7_75t_L g609 ( 
.A(n_568),
.Y(n_609)
);

INVx3_ASAP7_75t_L g610 ( 
.A(n_568),
.Y(n_610)
);

INVx4_ASAP7_75t_L g611 ( 
.A(n_568),
.Y(n_611)
);

NOR2xp33_ASAP7_75t_L g612 ( 
.A(n_571),
.B(n_448),
.Y(n_612)
);

OAI22xp33_ASAP7_75t_L g613 ( 
.A1(n_582),
.A2(n_433),
.B1(n_481),
.B2(n_407),
.Y(n_613)
);

INVx2_ASAP7_75t_L g614 ( 
.A(n_568),
.Y(n_614)
);

INVx3_ASAP7_75t_L g615 ( 
.A(n_568),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_568),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_578),
.Y(n_617)
);

INVx2_ASAP7_75t_L g618 ( 
.A(n_578),
.Y(n_618)
);

BUFx6f_ASAP7_75t_L g619 ( 
.A(n_578),
.Y(n_619)
);

INVx3_ASAP7_75t_L g620 ( 
.A(n_578),
.Y(n_620)
);

INVx2_ASAP7_75t_L g621 ( 
.A(n_578),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_SL g622 ( 
.A(n_575),
.B(n_427),
.Y(n_622)
);

BUFx10_ASAP7_75t_L g623 ( 
.A(n_586),
.Y(n_623)
);

INVx2_ASAP7_75t_L g624 ( 
.A(n_578),
.Y(n_624)
);

INVx2_ASAP7_75t_L g625 ( 
.A(n_507),
.Y(n_625)
);

INVx2_ASAP7_75t_L g626 ( 
.A(n_507),
.Y(n_626)
);

NOR2xp33_ASAP7_75t_L g627 ( 
.A(n_542),
.B(n_491),
.Y(n_627)
);

OR2x6_ASAP7_75t_L g628 ( 
.A(n_562),
.B(n_428),
.Y(n_628)
);

INVx1_ASAP7_75t_SL g629 ( 
.A(n_510),
.Y(n_629)
);

BUFx2_ASAP7_75t_L g630 ( 
.A(n_522),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_L g631 ( 
.A(n_583),
.B(n_428),
.Y(n_631)
);

AOI22xp33_ASAP7_75t_L g632 ( 
.A1(n_565),
.A2(n_434),
.B1(n_435),
.B2(n_430),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_550),
.Y(n_633)
);

OAI21xp33_ASAP7_75t_SL g634 ( 
.A1(n_544),
.A2(n_434),
.B(n_430),
.Y(n_634)
);

INVx2_ASAP7_75t_SL g635 ( 
.A(n_516),
.Y(n_635)
);

INVx3_ASAP7_75t_L g636 ( 
.A(n_550),
.Y(n_636)
);

NOR2xp33_ASAP7_75t_L g637 ( 
.A(n_506),
.B(n_495),
.Y(n_637)
);

INVx2_ASAP7_75t_L g638 ( 
.A(n_549),
.Y(n_638)
);

INVxp33_ASAP7_75t_L g639 ( 
.A(n_522),
.Y(n_639)
);

INVx2_ASAP7_75t_L g640 ( 
.A(n_549),
.Y(n_640)
);

INVxp33_ASAP7_75t_L g641 ( 
.A(n_537),
.Y(n_641)
);

INVx2_ASAP7_75t_SL g642 ( 
.A(n_516),
.Y(n_642)
);

INVx2_ASAP7_75t_L g643 ( 
.A(n_549),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_550),
.Y(n_644)
);

OAI22xp33_ASAP7_75t_L g645 ( 
.A1(n_582),
.A2(n_485),
.B1(n_304),
.B2(n_311),
.Y(n_645)
);

INVx2_ASAP7_75t_L g646 ( 
.A(n_559),
.Y(n_646)
);

NAND2xp33_ASAP7_75t_L g647 ( 
.A(n_530),
.B(n_543),
.Y(n_647)
);

INVx2_ASAP7_75t_L g648 ( 
.A(n_559),
.Y(n_648)
);

INVx2_ASAP7_75t_L g649 ( 
.A(n_559),
.Y(n_649)
);

BUFx3_ASAP7_75t_L g650 ( 
.A(n_583),
.Y(n_650)
);

BUFx6f_ASAP7_75t_L g651 ( 
.A(n_514),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_550),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_587),
.Y(n_653)
);

INVx2_ASAP7_75t_L g654 ( 
.A(n_587),
.Y(n_654)
);

NAND2xp33_ASAP7_75t_L g655 ( 
.A(n_554),
.B(n_544),
.Y(n_655)
);

INVx2_ASAP7_75t_L g656 ( 
.A(n_587),
.Y(n_656)
);

AOI22xp5_ASAP7_75t_L g657 ( 
.A1(n_565),
.A2(n_298),
.B1(n_318),
.B2(n_316),
.Y(n_657)
);

INVx2_ASAP7_75t_L g658 ( 
.A(n_515),
.Y(n_658)
);

NOR2xp33_ASAP7_75t_L g659 ( 
.A(n_558),
.B(n_435),
.Y(n_659)
);

BUFx3_ASAP7_75t_L g660 ( 
.A(n_583),
.Y(n_660)
);

INVx2_ASAP7_75t_L g661 ( 
.A(n_515),
.Y(n_661)
);

INVx2_ASAP7_75t_L g662 ( 
.A(n_515),
.Y(n_662)
);

BUFx2_ASAP7_75t_L g663 ( 
.A(n_537),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_545),
.Y(n_664)
);

AOI22xp33_ASAP7_75t_L g665 ( 
.A1(n_567),
.A2(n_438),
.B1(n_441),
.B2(n_436),
.Y(n_665)
);

NOR2xp33_ASAP7_75t_L g666 ( 
.A(n_556),
.B(n_441),
.Y(n_666)
);

INVx3_ASAP7_75t_L g667 ( 
.A(n_514),
.Y(n_667)
);

BUFx3_ASAP7_75t_L g668 ( 
.A(n_545),
.Y(n_668)
);

INVx2_ASAP7_75t_L g669 ( 
.A(n_508),
.Y(n_669)
);

NAND3xp33_ASAP7_75t_L g670 ( 
.A(n_521),
.B(n_445),
.C(n_444),
.Y(n_670)
);

OAI22xp5_ASAP7_75t_SL g671 ( 
.A1(n_534),
.A2(n_327),
.B1(n_336),
.B2(n_322),
.Y(n_671)
);

INVx2_ASAP7_75t_L g672 ( 
.A(n_508),
.Y(n_672)
);

BUFx6f_ASAP7_75t_L g673 ( 
.A(n_514),
.Y(n_673)
);

OR2x6_ASAP7_75t_L g674 ( 
.A(n_567),
.B(n_444),
.Y(n_674)
);

OR2x2_ASAP7_75t_L g675 ( 
.A(n_541),
.B(n_440),
.Y(n_675)
);

NAND2xp33_ASAP7_75t_SL g676 ( 
.A(n_548),
.B(n_338),
.Y(n_676)
);

INVx2_ASAP7_75t_L g677 ( 
.A(n_511),
.Y(n_677)
);

INVx8_ASAP7_75t_L g678 ( 
.A(n_567),
.Y(n_678)
);

AND2x2_ASAP7_75t_L g679 ( 
.A(n_521),
.B(n_445),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_SL g680 ( 
.A(n_548),
.B(n_450),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_546),
.Y(n_681)
);

OR2x2_ASAP7_75t_L g682 ( 
.A(n_541),
.B(n_450),
.Y(n_682)
);

INVx3_ASAP7_75t_L g683 ( 
.A(n_514),
.Y(n_683)
);

HB1xp67_ASAP7_75t_L g684 ( 
.A(n_518),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_SL g685 ( 
.A(n_529),
.B(n_451),
.Y(n_685)
);

INVx2_ASAP7_75t_L g686 ( 
.A(n_515),
.Y(n_686)
);

INVx2_ASAP7_75t_L g687 ( 
.A(n_525),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_546),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_551),
.Y(n_689)
);

INVx2_ASAP7_75t_SL g690 ( 
.A(n_529),
.Y(n_690)
);

BUFx6f_ASAP7_75t_L g691 ( 
.A(n_514),
.Y(n_691)
);

AOI22xp5_ASAP7_75t_L g692 ( 
.A1(n_535),
.A2(n_347),
.B1(n_360),
.B2(n_339),
.Y(n_692)
);

INVx2_ASAP7_75t_L g693 ( 
.A(n_525),
.Y(n_693)
);

INVx2_ASAP7_75t_L g694 ( 
.A(n_525),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_551),
.B(n_451),
.Y(n_695)
);

AOI22xp33_ASAP7_75t_L g696 ( 
.A1(n_567),
.A2(n_455),
.B1(n_456),
.B2(n_452),
.Y(n_696)
);

INVx5_ASAP7_75t_L g697 ( 
.A(n_514),
.Y(n_697)
);

INVx2_ASAP7_75t_SL g698 ( 
.A(n_504),
.Y(n_698)
);

INVx5_ASAP7_75t_L g699 ( 
.A(n_523),
.Y(n_699)
);

BUFx6f_ASAP7_75t_L g700 ( 
.A(n_523),
.Y(n_700)
);

AND3x2_ASAP7_75t_L g701 ( 
.A(n_538),
.B(n_227),
.C(n_226),
.Y(n_701)
);

INVx5_ASAP7_75t_L g702 ( 
.A(n_523),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_L g703 ( 
.A(n_553),
.B(n_452),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_553),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_L g705 ( 
.A(n_563),
.B(n_455),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_L g706 ( 
.A(n_563),
.B(n_456),
.Y(n_706)
);

BUFx6f_ASAP7_75t_SL g707 ( 
.A(n_504),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_569),
.Y(n_708)
);

INVx3_ASAP7_75t_L g709 ( 
.A(n_523),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_569),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_570),
.Y(n_711)
);

INVx2_ASAP7_75t_L g712 ( 
.A(n_511),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_570),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_L g714 ( 
.A(n_574),
.B(n_458),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_574),
.Y(n_715)
);

NAND3xp33_ASAP7_75t_L g716 ( 
.A(n_566),
.B(n_503),
.C(n_460),
.Y(n_716)
);

INVx2_ASAP7_75t_L g717 ( 
.A(n_525),
.Y(n_717)
);

BUFx3_ASAP7_75t_L g718 ( 
.A(n_577),
.Y(n_718)
);

INVx3_ASAP7_75t_L g719 ( 
.A(n_523),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_SL g720 ( 
.A(n_504),
.B(n_458),
.Y(n_720)
);

INVx3_ASAP7_75t_L g721 ( 
.A(n_523),
.Y(n_721)
);

INVx2_ASAP7_75t_L g722 ( 
.A(n_524),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_577),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_SL g724 ( 
.A(n_504),
.B(n_509),
.Y(n_724)
);

INVx2_ASAP7_75t_L g725 ( 
.A(n_524),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_L g726 ( 
.A(n_580),
.B(n_460),
.Y(n_726)
);

NOR2xp33_ASAP7_75t_L g727 ( 
.A(n_573),
.B(n_461),
.Y(n_727)
);

INVx2_ASAP7_75t_L g728 ( 
.A(n_524),
.Y(n_728)
);

AND2x2_ASAP7_75t_L g729 ( 
.A(n_509),
.B(n_461),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_580),
.B(n_462),
.Y(n_730)
);

BUFx2_ASAP7_75t_L g731 ( 
.A(n_520),
.Y(n_731)
);

BUFx3_ASAP7_75t_L g732 ( 
.A(n_585),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_L g733 ( 
.A(n_585),
.B(n_462),
.Y(n_733)
);

INVx2_ASAP7_75t_L g734 ( 
.A(n_512),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_555),
.Y(n_735)
);

INVxp33_ASAP7_75t_L g736 ( 
.A(n_519),
.Y(n_736)
);

INVx4_ASAP7_75t_L g737 ( 
.A(n_531),
.Y(n_737)
);

INVx2_ASAP7_75t_L g738 ( 
.A(n_512),
.Y(n_738)
);

OR2x6_ASAP7_75t_L g739 ( 
.A(n_608),
.B(n_628),
.Y(n_739)
);

INVx2_ASAP7_75t_L g740 ( 
.A(n_591),
.Y(n_740)
);

INVx2_ASAP7_75t_L g741 ( 
.A(n_591),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_668),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_L g743 ( 
.A(n_612),
.B(n_509),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_SL g744 ( 
.A(n_588),
.B(n_555),
.Y(n_744)
);

AND2x4_ASAP7_75t_L g745 ( 
.A(n_674),
.B(n_509),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_SL g746 ( 
.A(n_588),
.B(n_557),
.Y(n_746)
);

NOR2xp33_ASAP7_75t_L g747 ( 
.A(n_593),
.B(n_535),
.Y(n_747)
);

INVx2_ASAP7_75t_L g748 ( 
.A(n_638),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_666),
.B(n_557),
.Y(n_749)
);

INVx4_ASAP7_75t_L g750 ( 
.A(n_678),
.Y(n_750)
);

INVx2_ASAP7_75t_L g751 ( 
.A(n_591),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_L g752 ( 
.A(n_595),
.B(n_561),
.Y(n_752)
);

INVx2_ASAP7_75t_SL g753 ( 
.A(n_682),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_SL g754 ( 
.A(n_594),
.B(n_561),
.Y(n_754)
);

INVx2_ASAP7_75t_L g755 ( 
.A(n_592),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_668),
.Y(n_756)
);

A2O1A1Ixp33_ASAP7_75t_L g757 ( 
.A1(n_634),
.A2(n_467),
.B(n_469),
.C(n_465),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_L g758 ( 
.A(n_601),
.B(n_581),
.Y(n_758)
);

NOR3xp33_ASAP7_75t_L g759 ( 
.A(n_630),
.B(n_663),
.C(n_731),
.Y(n_759)
);

NOR2xp33_ASAP7_75t_R g760 ( 
.A(n_623),
.B(n_527),
.Y(n_760)
);

NOR2xp33_ASAP7_75t_L g761 ( 
.A(n_635),
.B(n_536),
.Y(n_761)
);

INVxp67_ASAP7_75t_L g762 ( 
.A(n_663),
.Y(n_762)
);

BUFx6f_ASAP7_75t_L g763 ( 
.A(n_619),
.Y(n_763)
);

INVx2_ASAP7_75t_L g764 ( 
.A(n_592),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_668),
.Y(n_765)
);

AND2x2_ASAP7_75t_L g766 ( 
.A(n_639),
.B(n_560),
.Y(n_766)
);

NOR2xp33_ASAP7_75t_L g767 ( 
.A(n_635),
.B(n_536),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_718),
.Y(n_768)
);

AOI22xp5_ASAP7_75t_L g769 ( 
.A1(n_608),
.A2(n_584),
.B1(n_581),
.B2(n_388),
.Y(n_769)
);

NOR2xp33_ASAP7_75t_L g770 ( 
.A(n_642),
.B(n_584),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_727),
.B(n_465),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_L g772 ( 
.A(n_608),
.B(n_467),
.Y(n_772)
);

INVx2_ASAP7_75t_L g773 ( 
.A(n_638),
.Y(n_773)
);

AOI21xp5_ASAP7_75t_L g774 ( 
.A1(n_633),
.A2(n_472),
.B(n_469),
.Y(n_774)
);

BUFx3_ASAP7_75t_L g775 ( 
.A(n_623),
.Y(n_775)
);

BUFx8_ASAP7_75t_L g776 ( 
.A(n_731),
.Y(n_776)
);

NOR2xp33_ASAP7_75t_L g777 ( 
.A(n_642),
.B(n_362),
.Y(n_777)
);

BUFx6f_ASAP7_75t_L g778 ( 
.A(n_619),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_L g779 ( 
.A(n_679),
.B(n_473),
.Y(n_779)
);

O2A1O1Ixp33_ASAP7_75t_L g780 ( 
.A1(n_634),
.A2(n_231),
.B(n_242),
.C(n_228),
.Y(n_780)
);

INVx2_ASAP7_75t_L g781 ( 
.A(n_638),
.Y(n_781)
);

BUFx2_ASAP7_75t_L g782 ( 
.A(n_675),
.Y(n_782)
);

INVx4_ASAP7_75t_L g783 ( 
.A(n_678),
.Y(n_783)
);

AND2x6_ASAP7_75t_L g784 ( 
.A(n_607),
.B(n_215),
.Y(n_784)
);

AO22x2_ASAP7_75t_L g785 ( 
.A1(n_594),
.A2(n_534),
.B1(n_538),
.B2(n_519),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_718),
.Y(n_786)
);

NOR2xp33_ASAP7_75t_L g787 ( 
.A(n_690),
.B(n_365),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_SL g788 ( 
.A(n_636),
.B(n_572),
.Y(n_788)
);

INVx2_ASAP7_75t_SL g789 ( 
.A(n_682),
.Y(n_789)
);

NOR2xp67_ASAP7_75t_L g790 ( 
.A(n_684),
.B(n_475),
.Y(n_790)
);

AO22x2_ASAP7_75t_L g791 ( 
.A1(n_736),
.A2(n_538),
.B1(n_479),
.B2(n_480),
.Y(n_791)
);

NOR2x1p5_ASAP7_75t_L g792 ( 
.A(n_670),
.B(n_538),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_L g793 ( 
.A(n_659),
.B(n_477),
.Y(n_793)
);

BUFx6f_ASAP7_75t_L g794 ( 
.A(n_619),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_L g795 ( 
.A(n_698),
.B(n_477),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_SL g796 ( 
.A(n_636),
.B(n_479),
.Y(n_796)
);

OR2x2_ASAP7_75t_L g797 ( 
.A(n_629),
.B(n_540),
.Y(n_797)
);

OR2x6_ASAP7_75t_L g798 ( 
.A(n_628),
.B(n_678),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_L g799 ( 
.A(n_698),
.B(n_480),
.Y(n_799)
);

CKINVDCx5p33_ASAP7_75t_R g800 ( 
.A(n_623),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_SL g801 ( 
.A(n_636),
.B(n_483),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_L g802 ( 
.A(n_603),
.B(n_483),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_L g803 ( 
.A(n_603),
.B(n_729),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_L g804 ( 
.A(n_729),
.B(n_484),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_718),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_SL g806 ( 
.A(n_636),
.B(n_484),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_L g807 ( 
.A(n_674),
.B(n_486),
.Y(n_807)
);

AND2x2_ASAP7_75t_L g808 ( 
.A(n_641),
.B(n_576),
.Y(n_808)
);

INVx2_ASAP7_75t_L g809 ( 
.A(n_640),
.Y(n_809)
);

AOI22xp33_ASAP7_75t_L g810 ( 
.A1(n_628),
.A2(n_501),
.B1(n_497),
.B2(n_503),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_L g811 ( 
.A(n_674),
.B(n_494),
.Y(n_811)
);

INVx2_ASAP7_75t_L g812 ( 
.A(n_732),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_L g813 ( 
.A(n_674),
.B(n_497),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_L g814 ( 
.A(n_674),
.B(n_732),
.Y(n_814)
);

AO22x2_ASAP7_75t_L g815 ( 
.A1(n_671),
.A2(n_499),
.B1(n_500),
.B2(n_502),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_732),
.Y(n_816)
);

NOR2xp33_ASAP7_75t_L g817 ( 
.A(n_690),
.B(n_369),
.Y(n_817)
);

INVx2_ASAP7_75t_L g818 ( 
.A(n_640),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_664),
.Y(n_819)
);

NOR2xp33_ASAP7_75t_L g820 ( 
.A(n_637),
.B(n_371),
.Y(n_820)
);

OAI22xp5_ASAP7_75t_L g821 ( 
.A1(n_678),
.A2(n_372),
.B1(n_375),
.B2(n_376),
.Y(n_821)
);

AOI22xp5_ASAP7_75t_L g822 ( 
.A1(n_655),
.A2(n_356),
.B1(n_500),
.B2(n_502),
.Y(n_822)
);

INVx2_ASAP7_75t_SL g823 ( 
.A(n_623),
.Y(n_823)
);

OR2x2_ASAP7_75t_L g824 ( 
.A(n_628),
.B(n_564),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_L g825 ( 
.A(n_665),
.B(n_499),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_SL g826 ( 
.A(n_619),
.B(n_501),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_SL g827 ( 
.A(n_619),
.B(n_356),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_L g828 ( 
.A(n_696),
.B(n_201),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_SL g829 ( 
.A(n_619),
.B(n_268),
.Y(n_829)
);

HB1xp67_ASAP7_75t_L g830 ( 
.A(n_628),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_627),
.B(n_230),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_L g832 ( 
.A(n_685),
.B(n_264),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_681),
.B(n_295),
.Y(n_833)
);

INVx2_ASAP7_75t_L g834 ( 
.A(n_640),
.Y(n_834)
);

INVx2_ASAP7_75t_L g835 ( 
.A(n_643),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_SL g836 ( 
.A(n_644),
.B(n_341),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_681),
.Y(n_837)
);

OR2x6_ASAP7_75t_L g838 ( 
.A(n_671),
.B(n_351),
.Y(n_838)
);

NOR2xp33_ASAP7_75t_L g839 ( 
.A(n_680),
.B(n_381),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_L g840 ( 
.A(n_688),
.B(n_532),
.Y(n_840)
);

AND2x2_ASAP7_75t_L g841 ( 
.A(n_692),
.B(n_271),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_688),
.B(n_532),
.Y(n_842)
);

AND2x2_ASAP7_75t_L g843 ( 
.A(n_692),
.B(n_271),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_L g844 ( 
.A(n_689),
.B(n_351),
.Y(n_844)
);

OAI22xp5_ASAP7_75t_L g845 ( 
.A1(n_689),
.A2(n_383),
.B1(n_384),
.B2(n_393),
.Y(n_845)
);

OAI22xp5_ASAP7_75t_L g846 ( 
.A1(n_704),
.A2(n_389),
.B1(n_242),
.B2(n_391),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_L g847 ( 
.A(n_704),
.B(n_379),
.Y(n_847)
);

NOR2xp33_ASAP7_75t_L g848 ( 
.A(n_622),
.B(n_337),
.Y(n_848)
);

NAND2xp33_ASAP7_75t_L g849 ( 
.A(n_644),
.B(n_228),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_708),
.B(n_379),
.Y(n_850)
);

AND2x2_ASAP7_75t_L g851 ( 
.A(n_647),
.B(n_337),
.Y(n_851)
);

AND2x2_ASAP7_75t_L g852 ( 
.A(n_632),
.B(n_337),
.Y(n_852)
);

INVx2_ASAP7_75t_L g853 ( 
.A(n_600),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_708),
.B(n_231),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_L g855 ( 
.A(n_710),
.B(n_254),
.Y(n_855)
);

O2A1O1Ixp33_ASAP7_75t_L g856 ( 
.A1(n_710),
.A2(n_315),
.B(n_254),
.C(n_256),
.Y(n_856)
);

BUFx3_ASAP7_75t_L g857 ( 
.A(n_650),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_L g858 ( 
.A(n_711),
.B(n_256),
.Y(n_858)
);

AOI22xp33_ASAP7_75t_L g859 ( 
.A1(n_657),
.A2(n_598),
.B1(n_715),
.B2(n_713),
.Y(n_859)
);

NOR2xp33_ASAP7_75t_L g860 ( 
.A(n_724),
.B(n_342),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_L g861 ( 
.A(n_713),
.B(n_282),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_715),
.B(n_282),
.Y(n_862)
);

NOR2xp33_ASAP7_75t_L g863 ( 
.A(n_597),
.B(n_267),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_723),
.B(n_285),
.Y(n_864)
);

BUFx6f_ASAP7_75t_SL g865 ( 
.A(n_701),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_723),
.Y(n_866)
);

AOI22xp5_ASAP7_75t_L g867 ( 
.A1(n_707),
.A2(n_223),
.B1(n_239),
.B2(n_395),
.Y(n_867)
);

NAND3xp33_ASAP7_75t_L g868 ( 
.A(n_676),
.B(n_657),
.C(n_645),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_652),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_L g870 ( 
.A(n_631),
.B(n_285),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_652),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_SL g872 ( 
.A(n_650),
.B(n_222),
.Y(n_872)
);

NOR3xp33_ASAP7_75t_L g873 ( 
.A(n_613),
.B(n_270),
.C(n_287),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_L g874 ( 
.A(n_695),
.B(n_287),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_L g875 ( 
.A(n_703),
.B(n_705),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_SL g876 ( 
.A(n_650),
.B(n_222),
.Y(n_876)
);

INVx2_ASAP7_75t_L g877 ( 
.A(n_600),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_SL g878 ( 
.A(n_660),
.B(n_353),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_735),
.Y(n_879)
);

NOR2xp33_ASAP7_75t_L g880 ( 
.A(n_660),
.B(n_290),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_735),
.Y(n_881)
);

NAND3xp33_ASAP7_75t_L g882 ( 
.A(n_716),
.B(n_299),
.C(n_290),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_L g883 ( 
.A(n_706),
.B(n_299),
.Y(n_883)
);

BUFx3_ASAP7_75t_L g884 ( 
.A(n_660),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_L g885 ( 
.A(n_714),
.B(n_312),
.Y(n_885)
);

NOR2xp33_ASAP7_75t_L g886 ( 
.A(n_707),
.B(n_312),
.Y(n_886)
);

AND2x4_ASAP7_75t_L g887 ( 
.A(n_720),
.B(n_726),
.Y(n_887)
);

INVx2_ASAP7_75t_L g888 ( 
.A(n_602),
.Y(n_888)
);

NOR2xp33_ASAP7_75t_L g889 ( 
.A(n_707),
.B(n_313),
.Y(n_889)
);

NOR2xp33_ASAP7_75t_L g890 ( 
.A(n_707),
.B(n_313),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_L g891 ( 
.A(n_730),
.B(n_315),
.Y(n_891)
);

INVxp67_ASAP7_75t_L g892 ( 
.A(n_733),
.Y(n_892)
);

NOR2xp33_ASAP7_75t_L g893 ( 
.A(n_609),
.B(n_324),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_SL g894 ( 
.A(n_609),
.B(n_353),
.Y(n_894)
);

INVx2_ASAP7_75t_SL g895 ( 
.A(n_658),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_L g896 ( 
.A(n_653),
.B(n_324),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_819),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_L g898 ( 
.A(n_892),
.B(n_653),
.Y(n_898)
);

HB1xp67_ASAP7_75t_L g899 ( 
.A(n_762),
.Y(n_899)
);

BUFx3_ASAP7_75t_L g900 ( 
.A(n_776),
.Y(n_900)
);

CKINVDCx5p33_ASAP7_75t_R g901 ( 
.A(n_760),
.Y(n_901)
);

AND2x4_ASAP7_75t_L g902 ( 
.A(n_798),
.B(n_596),
.Y(n_902)
);

BUFx3_ASAP7_75t_L g903 ( 
.A(n_776),
.Y(n_903)
);

INVx3_ASAP7_75t_L g904 ( 
.A(n_750),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_SL g905 ( 
.A(n_750),
.B(n_609),
.Y(n_905)
);

INVx2_ASAP7_75t_L g906 ( 
.A(n_748),
.Y(n_906)
);

OAI21xp33_ASAP7_75t_SL g907 ( 
.A1(n_747),
.A2(n_611),
.B(n_609),
.Y(n_907)
);

INVxp67_ASAP7_75t_L g908 ( 
.A(n_782),
.Y(n_908)
);

AOI22xp33_ASAP7_75t_SL g909 ( 
.A1(n_747),
.A2(n_292),
.B1(n_277),
.B2(n_291),
.Y(n_909)
);

AOI22xp5_ASAP7_75t_L g910 ( 
.A1(n_820),
.A2(n_611),
.B1(n_615),
.B2(n_596),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_837),
.Y(n_911)
);

INVx2_ASAP7_75t_L g912 ( 
.A(n_748),
.Y(n_912)
);

INVx3_ASAP7_75t_L g913 ( 
.A(n_783),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_866),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_L g915 ( 
.A(n_820),
.B(n_646),
.Y(n_915)
);

NOR3xp33_ASAP7_75t_SL g916 ( 
.A(n_788),
.B(n_329),
.C(n_325),
.Y(n_916)
);

BUFx2_ASAP7_75t_L g917 ( 
.A(n_797),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_L g918 ( 
.A(n_771),
.B(n_646),
.Y(n_918)
);

NOR2xp33_ASAP7_75t_R g919 ( 
.A(n_800),
.B(n_596),
.Y(n_919)
);

AND2x4_ASAP7_75t_L g920 ( 
.A(n_798),
.B(n_596),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_L g921 ( 
.A(n_743),
.B(n_648),
.Y(n_921)
);

INVx2_ASAP7_75t_SL g922 ( 
.A(n_808),
.Y(n_922)
);

CKINVDCx5p33_ASAP7_75t_R g923 ( 
.A(n_760),
.Y(n_923)
);

INVx2_ASAP7_75t_SL g924 ( 
.A(n_766),
.Y(n_924)
);

BUFx8_ASAP7_75t_L g925 ( 
.A(n_865),
.Y(n_925)
);

INVxp67_ASAP7_75t_L g926 ( 
.A(n_753),
.Y(n_926)
);

BUFx6f_ASAP7_75t_L g927 ( 
.A(n_763),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_869),
.Y(n_928)
);

HB1xp67_ASAP7_75t_L g929 ( 
.A(n_745),
.Y(n_929)
);

BUFx6f_ASAP7_75t_L g930 ( 
.A(n_763),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_871),
.Y(n_931)
);

INVx2_ASAP7_75t_SL g932 ( 
.A(n_789),
.Y(n_932)
);

INVx3_ASAP7_75t_L g933 ( 
.A(n_783),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_879),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_L g935 ( 
.A(n_810),
.B(n_648),
.Y(n_935)
);

BUFx12f_ASAP7_75t_SL g936 ( 
.A(n_838),
.Y(n_936)
);

INVx4_ASAP7_75t_L g937 ( 
.A(n_798),
.Y(n_937)
);

BUFx3_ASAP7_75t_L g938 ( 
.A(n_775),
.Y(n_938)
);

AOI22xp5_ASAP7_75t_L g939 ( 
.A1(n_868),
.A2(n_859),
.B1(n_810),
.B2(n_767),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_L g940 ( 
.A(n_793),
.B(n_648),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_L g941 ( 
.A(n_802),
.B(n_649),
.Y(n_941)
);

CKINVDCx20_ASAP7_75t_R g942 ( 
.A(n_775),
.Y(n_942)
);

OR2x6_ASAP7_75t_L g943 ( 
.A(n_739),
.B(n_649),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_L g944 ( 
.A(n_803),
.B(n_649),
.Y(n_944)
);

OR2x2_ASAP7_75t_SL g945 ( 
.A(n_824),
.B(n_325),
.Y(n_945)
);

AOI22xp33_ASAP7_75t_L g946 ( 
.A1(n_852),
.A2(n_656),
.B1(n_654),
.B2(n_626),
.Y(n_946)
);

AND2x4_ASAP7_75t_L g947 ( 
.A(n_739),
.B(n_610),
.Y(n_947)
);

OR2x2_ASAP7_75t_L g948 ( 
.A(n_759),
.B(n_658),
.Y(n_948)
);

AND2x2_ASAP7_75t_SL g949 ( 
.A(n_830),
.B(n_358),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_881),
.Y(n_950)
);

AOI21x1_ASAP7_75t_L g951 ( 
.A1(n_744),
.A2(n_590),
.B(n_589),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_L g952 ( 
.A(n_831),
.B(n_654),
.Y(n_952)
);

INVx2_ASAP7_75t_L g953 ( 
.A(n_773),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_840),
.Y(n_954)
);

INVx3_ASAP7_75t_L g955 ( 
.A(n_857),
.Y(n_955)
);

INVx1_ASAP7_75t_L g956 ( 
.A(n_842),
.Y(n_956)
);

AND2x2_ASAP7_75t_L g957 ( 
.A(n_761),
.B(n_654),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_L g958 ( 
.A(n_770),
.B(n_804),
.Y(n_958)
);

AOI22xp33_ASAP7_75t_L g959 ( 
.A1(n_815),
.A2(n_656),
.B1(n_626),
.B2(n_625),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_SL g960 ( 
.A(n_814),
.B(n_610),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_807),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_L g962 ( 
.A(n_770),
.B(n_656),
.Y(n_962)
);

A2O1A1Ixp33_ASAP7_75t_L g963 ( 
.A1(n_780),
.A2(n_767),
.B(n_761),
.C(n_757),
.Y(n_963)
);

AOI22xp33_ASAP7_75t_L g964 ( 
.A1(n_815),
.A2(n_672),
.B1(n_625),
.B2(n_712),
.Y(n_964)
);

NOR2xp33_ASAP7_75t_L g965 ( 
.A(n_830),
.B(n_615),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_811),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_L g967 ( 
.A(n_875),
.B(n_669),
.Y(n_967)
);

NOR3xp33_ASAP7_75t_L g968 ( 
.A(n_790),
.B(n_350),
.C(n_349),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_L g969 ( 
.A(n_779),
.B(n_758),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_813),
.Y(n_970)
);

INVx2_ASAP7_75t_L g971 ( 
.A(n_773),
.Y(n_971)
);

BUFx8_ASAP7_75t_L g972 ( 
.A(n_865),
.Y(n_972)
);

CKINVDCx5p33_ASAP7_75t_R g973 ( 
.A(n_823),
.Y(n_973)
);

AOI22xp33_ASAP7_75t_L g974 ( 
.A1(n_815),
.A2(n_838),
.B1(n_843),
.B2(n_841),
.Y(n_974)
);

AND2x4_ASAP7_75t_L g975 ( 
.A(n_739),
.B(n_620),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_896),
.Y(n_976)
);

NOR2xp33_ASAP7_75t_R g977 ( 
.A(n_857),
.B(n_620),
.Y(n_977)
);

AND2x2_ASAP7_75t_L g978 ( 
.A(n_851),
.B(n_734),
.Y(n_978)
);

BUFx6f_ASAP7_75t_L g979 ( 
.A(n_763),
.Y(n_979)
);

INVx3_ASAP7_75t_L g980 ( 
.A(n_884),
.Y(n_980)
);

INVx1_ASAP7_75t_L g981 ( 
.A(n_844),
.Y(n_981)
);

OR2x6_ASAP7_75t_L g982 ( 
.A(n_745),
.B(n_734),
.Y(n_982)
);

OAI21xp5_ASAP7_75t_L g983 ( 
.A1(n_796),
.A2(n_590),
.B(n_589),
.Y(n_983)
);

BUFx6f_ASAP7_75t_L g984 ( 
.A(n_763),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_L g985 ( 
.A(n_749),
.B(n_669),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_SL g986 ( 
.A(n_778),
.B(n_614),
.Y(n_986)
);

NAND2xp5_ASAP7_75t_L g987 ( 
.A(n_887),
.B(n_672),
.Y(n_987)
);

INVx2_ASAP7_75t_L g988 ( 
.A(n_781),
.Y(n_988)
);

NOR2x2_ASAP7_75t_L g989 ( 
.A(n_838),
.B(n_658),
.Y(n_989)
);

AND2x4_ASAP7_75t_SL g990 ( 
.A(n_887),
.B(n_277),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_L g991 ( 
.A(n_772),
.B(n_677),
.Y(n_991)
);

AND2x2_ASAP7_75t_L g992 ( 
.A(n_777),
.B(n_787),
.Y(n_992)
);

BUFx4f_ASAP7_75t_L g993 ( 
.A(n_784),
.Y(n_993)
);

AND2x4_ASAP7_75t_L g994 ( 
.A(n_792),
.B(n_614),
.Y(n_994)
);

INVx2_ASAP7_75t_L g995 ( 
.A(n_781),
.Y(n_995)
);

INVx2_ASAP7_75t_L g996 ( 
.A(n_809),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_847),
.Y(n_997)
);

AND2x2_ASAP7_75t_L g998 ( 
.A(n_777),
.B(n_734),
.Y(n_998)
);

INVx8_ASAP7_75t_L g999 ( 
.A(n_784),
.Y(n_999)
);

AND2x4_ASAP7_75t_L g1000 ( 
.A(n_884),
.B(n_618),
.Y(n_1000)
);

INVx5_ASAP7_75t_L g1001 ( 
.A(n_778),
.Y(n_1001)
);

INVx1_ASAP7_75t_L g1002 ( 
.A(n_850),
.Y(n_1002)
);

INVx1_ASAP7_75t_L g1003 ( 
.A(n_854),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_855),
.Y(n_1004)
);

INVx1_ASAP7_75t_L g1005 ( 
.A(n_858),
.Y(n_1005)
);

INVx2_ASAP7_75t_SL g1006 ( 
.A(n_791),
.Y(n_1006)
);

NAND2xp5_ASAP7_75t_L g1007 ( 
.A(n_833),
.B(n_712),
.Y(n_1007)
);

INVx2_ASAP7_75t_L g1008 ( 
.A(n_809),
.Y(n_1008)
);

INVx1_ASAP7_75t_SL g1009 ( 
.A(n_886),
.Y(n_1009)
);

INVx1_ASAP7_75t_L g1010 ( 
.A(n_861),
.Y(n_1010)
);

CKINVDCx5p33_ASAP7_75t_R g1011 ( 
.A(n_821),
.Y(n_1011)
);

OR2x4_ASAP7_75t_L g1012 ( 
.A(n_787),
.B(n_350),
.Y(n_1012)
);

INVx2_ASAP7_75t_L g1013 ( 
.A(n_818),
.Y(n_1013)
);

NOR2xp33_ASAP7_75t_L g1014 ( 
.A(n_839),
.B(n_599),
.Y(n_1014)
);

BUFx6f_ASAP7_75t_L g1015 ( 
.A(n_794),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_L g1016 ( 
.A(n_880),
.B(n_738),
.Y(n_1016)
);

AOI221xp5_ASAP7_75t_SL g1017 ( 
.A1(n_757),
.A2(n_391),
.B1(n_361),
.B2(n_377),
.C(n_382),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_L g1018 ( 
.A(n_880),
.B(n_738),
.Y(n_1018)
);

AOI21xp33_ASAP7_75t_L g1019 ( 
.A1(n_839),
.A2(n_604),
.B(n_599),
.Y(n_1019)
);

INVx1_ASAP7_75t_L g1020 ( 
.A(n_862),
.Y(n_1020)
);

CKINVDCx5p33_ASAP7_75t_R g1021 ( 
.A(n_863),
.Y(n_1021)
);

NAND2xp5_ASAP7_75t_L g1022 ( 
.A(n_886),
.B(n_738),
.Y(n_1022)
);

CKINVDCx5p33_ASAP7_75t_R g1023 ( 
.A(n_863),
.Y(n_1023)
);

NOR2xp33_ASAP7_75t_L g1024 ( 
.A(n_889),
.B(n_604),
.Y(n_1024)
);

INVx3_ASAP7_75t_L g1025 ( 
.A(n_794),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_L g1026 ( 
.A(n_889),
.B(n_661),
.Y(n_1026)
);

AND2x4_ASAP7_75t_L g1027 ( 
.A(n_873),
.B(n_618),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_L g1028 ( 
.A(n_890),
.B(n_860),
.Y(n_1028)
);

INVx2_ASAP7_75t_SL g1029 ( 
.A(n_791),
.Y(n_1029)
);

BUFx2_ASAP7_75t_L g1030 ( 
.A(n_791),
.Y(n_1030)
);

NAND2xp5_ASAP7_75t_SL g1031 ( 
.A(n_812),
.B(n_769),
.Y(n_1031)
);

NOR2xp33_ASAP7_75t_R g1032 ( 
.A(n_742),
.B(n_667),
.Y(n_1032)
);

BUFx4f_ASAP7_75t_L g1033 ( 
.A(n_784),
.Y(n_1033)
);

INVx2_ASAP7_75t_L g1034 ( 
.A(n_834),
.Y(n_1034)
);

NAND2xp5_ASAP7_75t_L g1035 ( 
.A(n_890),
.B(n_860),
.Y(n_1035)
);

BUFx6f_ASAP7_75t_L g1036 ( 
.A(n_834),
.Y(n_1036)
);

AND2x4_ASAP7_75t_L g1037 ( 
.A(n_882),
.B(n_621),
.Y(n_1037)
);

NOR2xp33_ASAP7_75t_L g1038 ( 
.A(n_848),
.B(n_606),
.Y(n_1038)
);

INVx4_ASAP7_75t_L g1039 ( 
.A(n_756),
.Y(n_1039)
);

NOR2xp33_ASAP7_75t_L g1040 ( 
.A(n_848),
.B(n_606),
.Y(n_1040)
);

NOR2xp33_ASAP7_75t_L g1041 ( 
.A(n_752),
.B(n_616),
.Y(n_1041)
);

BUFx6f_ASAP7_75t_L g1042 ( 
.A(n_835),
.Y(n_1042)
);

NAND2xp5_ASAP7_75t_L g1043 ( 
.A(n_795),
.B(n_661),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_L g1044 ( 
.A(n_799),
.B(n_661),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_SL g1045 ( 
.A(n_765),
.B(n_621),
.Y(n_1045)
);

INVx1_ASAP7_75t_L g1046 ( 
.A(n_864),
.Y(n_1046)
);

AOI22xp33_ASAP7_75t_L g1047 ( 
.A1(n_785),
.A2(n_602),
.B1(n_605),
.B2(n_292),
.Y(n_1047)
);

AOI22xp33_ASAP7_75t_L g1048 ( 
.A1(n_785),
.A2(n_746),
.B1(n_754),
.B2(n_744),
.Y(n_1048)
);

OAI22xp5_ASAP7_75t_SL g1049 ( 
.A1(n_822),
.A2(n_361),
.B1(n_377),
.B2(n_382),
.Y(n_1049)
);

AND2x2_ASAP7_75t_L g1050 ( 
.A(n_817),
.B(n_662),
.Y(n_1050)
);

NAND2xp5_ASAP7_75t_L g1051 ( 
.A(n_817),
.B(n_662),
.Y(n_1051)
);

INVx2_ASAP7_75t_L g1052 ( 
.A(n_740),
.Y(n_1052)
);

NAND2xp5_ASAP7_75t_SL g1053 ( 
.A(n_768),
.B(n_621),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_796),
.Y(n_1054)
);

HB1xp67_ASAP7_75t_L g1055 ( 
.A(n_786),
.Y(n_1055)
);

AOI22xp5_ASAP7_75t_L g1056 ( 
.A1(n_893),
.A2(n_616),
.B1(n_617),
.B2(n_624),
.Y(n_1056)
);

CKINVDCx5p33_ASAP7_75t_R g1057 ( 
.A(n_845),
.Y(n_1057)
);

INVx2_ASAP7_75t_L g1058 ( 
.A(n_741),
.Y(n_1058)
);

HB1xp67_ASAP7_75t_L g1059 ( 
.A(n_805),
.Y(n_1059)
);

AND2x6_ASAP7_75t_SL g1060 ( 
.A(n_893),
.B(n_617),
.Y(n_1060)
);

BUFx3_ASAP7_75t_L g1061 ( 
.A(n_816),
.Y(n_1061)
);

BUFx10_ASAP7_75t_L g1062 ( 
.A(n_784),
.Y(n_1062)
);

BUFx6f_ASAP7_75t_L g1063 ( 
.A(n_895),
.Y(n_1063)
);

NOR3xp33_ASAP7_75t_SL g1064 ( 
.A(n_801),
.B(n_202),
.C(n_195),
.Y(n_1064)
);

AOI21x1_ASAP7_75t_L g1065 ( 
.A1(n_746),
.A2(n_624),
.B(n_722),
.Y(n_1065)
);

INVx1_ASAP7_75t_L g1066 ( 
.A(n_801),
.Y(n_1066)
);

INVxp67_ASAP7_75t_L g1067 ( 
.A(n_832),
.Y(n_1067)
);

AOI21xp5_ASAP7_75t_L g1068 ( 
.A1(n_806),
.A2(n_683),
.B(n_667),
.Y(n_1068)
);

INVx5_ASAP7_75t_L g1069 ( 
.A(n_784),
.Y(n_1069)
);

INVx3_ASAP7_75t_L g1070 ( 
.A(n_853),
.Y(n_1070)
);

INVx2_ASAP7_75t_L g1071 ( 
.A(n_751),
.Y(n_1071)
);

NOR2xp33_ASAP7_75t_L g1072 ( 
.A(n_1021),
.B(n_828),
.Y(n_1072)
);

AOI21xp5_ASAP7_75t_L g1073 ( 
.A1(n_958),
.A2(n_849),
.B(n_836),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_L g1074 ( 
.A(n_992),
.B(n_785),
.Y(n_1074)
);

NAND2x1p5_ASAP7_75t_L g1075 ( 
.A(n_937),
.B(n_1001),
.Y(n_1075)
);

AOI21xp5_ASAP7_75t_L g1076 ( 
.A1(n_969),
.A2(n_836),
.B(n_894),
.Y(n_1076)
);

INVx2_ASAP7_75t_L g1077 ( 
.A(n_906),
.Y(n_1077)
);

NAND2xp5_ASAP7_75t_SL g1078 ( 
.A(n_1023),
.B(n_867),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_SL g1079 ( 
.A(n_1028),
.B(n_825),
.Y(n_1079)
);

NAND2xp5_ASAP7_75t_L g1080 ( 
.A(n_939),
.B(n_754),
.Y(n_1080)
);

INVx2_ASAP7_75t_L g1081 ( 
.A(n_906),
.Y(n_1081)
);

NAND2xp5_ASAP7_75t_L g1082 ( 
.A(n_957),
.B(n_774),
.Y(n_1082)
);

AOI22xp33_ASAP7_75t_L g1083 ( 
.A1(n_949),
.A2(n_846),
.B1(n_877),
.B2(n_888),
.Y(n_1083)
);

AND2x4_ASAP7_75t_L g1084 ( 
.A(n_937),
.B(n_826),
.Y(n_1084)
);

AOI21xp5_ASAP7_75t_L g1085 ( 
.A1(n_967),
.A2(n_894),
.B(n_826),
.Y(n_1085)
);

NAND2x1p5_ASAP7_75t_L g1086 ( 
.A(n_1001),
.B(n_755),
.Y(n_1086)
);

BUFx6f_ASAP7_75t_L g1087 ( 
.A(n_927),
.Y(n_1087)
);

NOR3xp33_ASAP7_75t_SL g1088 ( 
.A(n_901),
.B(n_856),
.C(n_874),
.Y(n_1088)
);

AOI22xp33_ASAP7_75t_L g1089 ( 
.A1(n_949),
.A2(n_974),
.B1(n_1035),
.B2(n_1009),
.Y(n_1089)
);

OAI22xp5_ASAP7_75t_L g1090 ( 
.A1(n_963),
.A2(n_891),
.B1(n_885),
.B2(n_883),
.Y(n_1090)
);

INVx1_ASAP7_75t_L g1091 ( 
.A(n_897),
.Y(n_1091)
);

HB1xp67_ASAP7_75t_L g1092 ( 
.A(n_908),
.Y(n_1092)
);

AOI21xp5_ASAP7_75t_L g1093 ( 
.A1(n_915),
.A2(n_827),
.B(n_870),
.Y(n_1093)
);

A2O1A1Ixp33_ASAP7_75t_L g1094 ( 
.A1(n_963),
.A2(n_878),
.B(n_876),
.C(n_872),
.Y(n_1094)
);

OAI22xp5_ASAP7_75t_L g1095 ( 
.A1(n_974),
.A2(n_662),
.B1(n_693),
.B2(n_687),
.Y(n_1095)
);

NAND2x1p5_ASAP7_75t_L g1096 ( 
.A(n_1001),
.B(n_902),
.Y(n_1096)
);

INVx4_ASAP7_75t_L g1097 ( 
.A(n_1001),
.Y(n_1097)
);

O2A1O1Ixp33_ASAP7_75t_L g1098 ( 
.A1(n_899),
.A2(n_827),
.B(n_876),
.C(n_872),
.Y(n_1098)
);

A2O1A1Ixp33_ASAP7_75t_L g1099 ( 
.A1(n_1014),
.A2(n_878),
.B(n_829),
.C(n_694),
.Y(n_1099)
);

NAND2xp5_ASAP7_75t_SL g1100 ( 
.A(n_1057),
.B(n_737),
.Y(n_1100)
);

NAND2xp5_ASAP7_75t_L g1101 ( 
.A(n_954),
.B(n_764),
.Y(n_1101)
);

O2A1O1Ixp5_ASAP7_75t_SL g1102 ( 
.A1(n_986),
.A2(n_829),
.B(n_709),
.C(n_667),
.Y(n_1102)
);

NAND2xp5_ASAP7_75t_SL g1103 ( 
.A(n_1011),
.B(n_737),
.Y(n_1103)
);

INVx2_ASAP7_75t_L g1104 ( 
.A(n_912),
.Y(n_1104)
);

NOR2xp33_ASAP7_75t_L g1105 ( 
.A(n_917),
.B(n_737),
.Y(n_1105)
);

AOI22xp5_ASAP7_75t_L g1106 ( 
.A1(n_926),
.A2(n_686),
.B1(n_687),
.B2(n_693),
.Y(n_1106)
);

OAI22xp5_ASAP7_75t_L g1107 ( 
.A1(n_956),
.A2(n_693),
.B1(n_687),
.B2(n_686),
.Y(n_1107)
);

NOR2xp33_ASAP7_75t_L g1108 ( 
.A(n_899),
.B(n_667),
.Y(n_1108)
);

BUFx12f_ASAP7_75t_L g1109 ( 
.A(n_925),
.Y(n_1109)
);

BUFx6f_ASAP7_75t_L g1110 ( 
.A(n_927),
.Y(n_1110)
);

OAI22xp5_ASAP7_75t_L g1111 ( 
.A1(n_911),
.A2(n_717),
.B1(n_694),
.B2(n_709),
.Y(n_1111)
);

AND2x4_ASAP7_75t_L g1112 ( 
.A(n_929),
.B(n_694),
.Y(n_1112)
);

NAND3xp33_ASAP7_75t_SL g1113 ( 
.A(n_909),
.B(n_209),
.C(n_204),
.Y(n_1113)
);

OR2x6_ASAP7_75t_L g1114 ( 
.A(n_943),
.B(n_717),
.Y(n_1114)
);

NAND2xp5_ASAP7_75t_L g1115 ( 
.A(n_961),
.B(n_605),
.Y(n_1115)
);

OAI22xp5_ASAP7_75t_L g1116 ( 
.A1(n_914),
.A2(n_721),
.B1(n_719),
.B2(n_358),
.Y(n_1116)
);

O2A1O1Ixp33_ASAP7_75t_L g1117 ( 
.A1(n_916),
.A2(n_719),
.B(n_721),
.C(n_722),
.Y(n_1117)
);

NAND2xp5_ASAP7_75t_SL g1118 ( 
.A(n_932),
.B(n_651),
.Y(n_1118)
);

O2A1O1Ixp33_ASAP7_75t_L g1119 ( 
.A1(n_916),
.A2(n_721),
.B(n_725),
.C(n_722),
.Y(n_1119)
);

INVx1_ASAP7_75t_L g1120 ( 
.A(n_934),
.Y(n_1120)
);

INVx2_ASAP7_75t_L g1121 ( 
.A(n_912),
.Y(n_1121)
);

NAND2xp5_ASAP7_75t_SL g1122 ( 
.A(n_923),
.B(n_651),
.Y(n_1122)
);

AOI21xp5_ASAP7_75t_L g1123 ( 
.A1(n_962),
.A2(n_651),
.B(n_673),
.Y(n_1123)
);

AOI21xp5_ASAP7_75t_L g1124 ( 
.A1(n_921),
.A2(n_651),
.B(n_673),
.Y(n_1124)
);

AOI21xp5_ASAP7_75t_L g1125 ( 
.A1(n_1016),
.A2(n_651),
.B(n_673),
.Y(n_1125)
);

BUFx2_ASAP7_75t_L g1126 ( 
.A(n_942),
.Y(n_1126)
);

INVx3_ASAP7_75t_L g1127 ( 
.A(n_904),
.Y(n_1127)
);

XNOR2xp5_ASAP7_75t_L g1128 ( 
.A(n_900),
.B(n_725),
.Y(n_1128)
);

AOI21xp5_ASAP7_75t_L g1129 ( 
.A1(n_1018),
.A2(n_651),
.B(n_673),
.Y(n_1129)
);

INVx2_ASAP7_75t_L g1130 ( 
.A(n_953),
.Y(n_1130)
);

AOI21xp5_ASAP7_75t_L g1131 ( 
.A1(n_1041),
.A2(n_700),
.B(n_691),
.Y(n_1131)
);

AOI21xp5_ASAP7_75t_L g1132 ( 
.A1(n_1041),
.A2(n_700),
.B(n_691),
.Y(n_1132)
);

BUFx2_ASAP7_75t_L g1133 ( 
.A(n_936),
.Y(n_1133)
);

NOR2xp33_ASAP7_75t_L g1134 ( 
.A(n_929),
.B(n_728),
.Y(n_1134)
);

OAI22x1_ASAP7_75t_L g1135 ( 
.A1(n_1030),
.A2(n_922),
.B1(n_924),
.B2(n_994),
.Y(n_1135)
);

AOI22xp5_ASAP7_75t_L g1136 ( 
.A1(n_1024),
.A2(n_310),
.B1(n_221),
.B2(n_229),
.Y(n_1136)
);

AOI22xp5_ASAP7_75t_L g1137 ( 
.A1(n_1024),
.A2(n_314),
.B1(n_232),
.B2(n_235),
.Y(n_1137)
);

AOI21xp5_ASAP7_75t_L g1138 ( 
.A1(n_1051),
.A2(n_700),
.B(n_691),
.Y(n_1138)
);

NAND2xp5_ASAP7_75t_SL g1139 ( 
.A(n_977),
.B(n_673),
.Y(n_1139)
);

BUFx2_ASAP7_75t_L g1140 ( 
.A(n_982),
.Y(n_1140)
);

INVx2_ASAP7_75t_L g1141 ( 
.A(n_953),
.Y(n_1141)
);

BUFx2_ASAP7_75t_L g1142 ( 
.A(n_982),
.Y(n_1142)
);

AOI22xp33_ASAP7_75t_L g1143 ( 
.A1(n_1047),
.A2(n_291),
.B1(n_292),
.B2(n_303),
.Y(n_1143)
);

INVx3_ASAP7_75t_L g1144 ( 
.A(n_904),
.Y(n_1144)
);

AOI21xp5_ASAP7_75t_L g1145 ( 
.A1(n_918),
.A2(n_985),
.B(n_940),
.Y(n_1145)
);

OA22x2_ASAP7_75t_L g1146 ( 
.A1(n_990),
.A2(n_387),
.B1(n_284),
.B2(n_281),
.Y(n_1146)
);

NAND2xp5_ASAP7_75t_SL g1147 ( 
.A(n_977),
.B(n_673),
.Y(n_1147)
);

AOI21xp5_ASAP7_75t_L g1148 ( 
.A1(n_1014),
.A2(n_700),
.B(n_691),
.Y(n_1148)
);

NAND2xp5_ASAP7_75t_SL g1149 ( 
.A(n_919),
.B(n_691),
.Y(n_1149)
);

AOI21xp5_ASAP7_75t_L g1150 ( 
.A1(n_991),
.A2(n_700),
.B(n_691),
.Y(n_1150)
);

NOR2xp33_ASAP7_75t_L g1151 ( 
.A(n_1012),
.B(n_210),
.Y(n_1151)
);

AOI21x1_ASAP7_75t_L g1152 ( 
.A1(n_1065),
.A2(n_702),
.B(n_699),
.Y(n_1152)
);

OAI22xp5_ASAP7_75t_SL g1153 ( 
.A1(n_945),
.A2(n_280),
.B1(n_275),
.B2(n_265),
.Y(n_1153)
);

OAI22xp5_ASAP7_75t_L g1154 ( 
.A1(n_1012),
.A2(n_303),
.B1(n_333),
.B2(n_697),
.Y(n_1154)
);

INVx2_ASAP7_75t_L g1155 ( 
.A(n_971),
.Y(n_1155)
);

INVx2_ASAP7_75t_L g1156 ( 
.A(n_971),
.Y(n_1156)
);

OAI22x1_ASAP7_75t_L g1157 ( 
.A1(n_994),
.A2(n_258),
.B1(n_259),
.B2(n_250),
.Y(n_1157)
);

NAND2xp5_ASAP7_75t_L g1158 ( 
.A(n_966),
.B(n_697),
.Y(n_1158)
);

AOI21xp5_ASAP7_75t_L g1159 ( 
.A1(n_1038),
.A2(n_702),
.B(n_699),
.Y(n_1159)
);

AND2x4_ASAP7_75t_L g1160 ( 
.A(n_982),
.B(n_697),
.Y(n_1160)
);

AOI21x1_ASAP7_75t_L g1161 ( 
.A1(n_951),
.A2(n_699),
.B(n_697),
.Y(n_1161)
);

NAND2xp5_ASAP7_75t_L g1162 ( 
.A(n_970),
.B(n_697),
.Y(n_1162)
);

BUFx2_ASAP7_75t_L g1163 ( 
.A(n_919),
.Y(n_1163)
);

AOI21xp5_ASAP7_75t_L g1164 ( 
.A1(n_1040),
.A2(n_697),
.B(n_243),
.Y(n_1164)
);

NAND2xp5_ASAP7_75t_L g1165 ( 
.A(n_1003),
.B(n_333),
.Y(n_1165)
);

AOI21xp5_ASAP7_75t_L g1166 ( 
.A1(n_941),
.A2(n_334),
.B(n_261),
.Y(n_1166)
);

OR2x6_ASAP7_75t_SL g1167 ( 
.A(n_973),
.B(n_249),
.Y(n_1167)
);

AOI21xp5_ASAP7_75t_L g1168 ( 
.A1(n_1043),
.A2(n_1044),
.B(n_944),
.Y(n_1168)
);

OAI22xp5_ASAP7_75t_L g1169 ( 
.A1(n_1004),
.A2(n_335),
.B1(n_263),
.B2(n_294),
.Y(n_1169)
);

AND2x4_ASAP7_75t_L g1170 ( 
.A(n_943),
.B(n_2),
.Y(n_1170)
);

OR2x6_ASAP7_75t_L g1171 ( 
.A(n_943),
.B(n_251),
.Y(n_1171)
);

INVx2_ASAP7_75t_L g1172 ( 
.A(n_996),
.Y(n_1172)
);

AND2x2_ASAP7_75t_L g1173 ( 
.A(n_990),
.B(n_291),
.Y(n_1173)
);

BUFx6f_ASAP7_75t_L g1174 ( 
.A(n_927),
.Y(n_1174)
);

AOI21xp5_ASAP7_75t_L g1175 ( 
.A1(n_998),
.A2(n_366),
.B(n_302),
.Y(n_1175)
);

OAI22xp5_ASAP7_75t_L g1176 ( 
.A1(n_1005),
.A2(n_390),
.B1(n_380),
.B2(n_378),
.Y(n_1176)
);

NAND2xp5_ASAP7_75t_L g1177 ( 
.A(n_1010),
.B(n_4),
.Y(n_1177)
);

AOI21xp5_ASAP7_75t_L g1178 ( 
.A1(n_907),
.A2(n_332),
.B(n_317),
.Y(n_1178)
);

AOI22xp33_ASAP7_75t_SL g1179 ( 
.A1(n_1049),
.A2(n_291),
.B1(n_292),
.B2(n_343),
.Y(n_1179)
);

INVx1_ASAP7_75t_L g1180 ( 
.A(n_950),
.Y(n_1180)
);

CKINVDCx20_ASAP7_75t_R g1181 ( 
.A(n_925),
.Y(n_1181)
);

OAI22xp5_ASAP7_75t_L g1182 ( 
.A1(n_1020),
.A2(n_374),
.B1(n_368),
.B2(n_328),
.Y(n_1182)
);

NAND2xp5_ASAP7_75t_L g1183 ( 
.A(n_1046),
.B(n_4),
.Y(n_1183)
);

INVx2_ASAP7_75t_L g1184 ( 
.A(n_1008),
.Y(n_1184)
);

O2A1O1Ixp33_ASAP7_75t_SL g1185 ( 
.A1(n_905),
.A2(n_5),
.B(n_6),
.C(n_9),
.Y(n_1185)
);

BUFx3_ASAP7_75t_L g1186 ( 
.A(n_903),
.Y(n_1186)
);

NOR3xp33_ASAP7_75t_L g1187 ( 
.A(n_968),
.B(n_5),
.C(n_10),
.Y(n_1187)
);

NOR2xp33_ASAP7_75t_L g1188 ( 
.A(n_1067),
.B(n_11),
.Y(n_1188)
);

INVx3_ASAP7_75t_L g1189 ( 
.A(n_913),
.Y(n_1189)
);

CKINVDCx20_ASAP7_75t_R g1190 ( 
.A(n_972),
.Y(n_1190)
);

INVx1_ASAP7_75t_L g1191 ( 
.A(n_928),
.Y(n_1191)
);

AOI21xp5_ASAP7_75t_L g1192 ( 
.A1(n_1068),
.A2(n_321),
.B(n_251),
.Y(n_1192)
);

HB1xp67_ASAP7_75t_L g1193 ( 
.A(n_948),
.Y(n_1193)
);

NAND2xp5_ASAP7_75t_L g1194 ( 
.A(n_976),
.B(n_11),
.Y(n_1194)
);

A2O1A1Ixp33_ASAP7_75t_L g1195 ( 
.A1(n_965),
.A2(n_321),
.B(n_251),
.C(n_533),
.Y(n_1195)
);

BUFx2_ASAP7_75t_R g1196 ( 
.A(n_903),
.Y(n_1196)
);

INVx2_ASAP7_75t_SL g1197 ( 
.A(n_938),
.Y(n_1197)
);

AO22x1_ASAP7_75t_L g1198 ( 
.A1(n_968),
.A2(n_321),
.B1(n_251),
.B2(n_18),
.Y(n_1198)
);

INVx2_ASAP7_75t_L g1199 ( 
.A(n_1013),
.Y(n_1199)
);

AND2x4_ASAP7_75t_L g1200 ( 
.A(n_902),
.B(n_920),
.Y(n_1200)
);

O2A1O1Ixp33_ASAP7_75t_L g1201 ( 
.A1(n_1055),
.A2(n_14),
.B(n_19),
.C(n_25),
.Y(n_1201)
);

AND2x2_ASAP7_75t_L g1202 ( 
.A(n_978),
.B(n_25),
.Y(n_1202)
);

NOR2xp33_ASAP7_75t_L g1203 ( 
.A(n_898),
.B(n_26),
.Y(n_1203)
);

OAI21x1_ASAP7_75t_L g1204 ( 
.A1(n_983),
.A2(n_321),
.B(n_81),
.Y(n_1204)
);

O2A1O1Ixp33_ASAP7_75t_SL g1205 ( 
.A1(n_905),
.A2(n_26),
.B(n_27),
.C(n_30),
.Y(n_1205)
);

NOR2xp33_ASAP7_75t_L g1206 ( 
.A(n_1060),
.B(n_981),
.Y(n_1206)
);

AOI21xp5_ASAP7_75t_L g1207 ( 
.A1(n_1045),
.A2(n_1053),
.B(n_1022),
.Y(n_1207)
);

INVx4_ASAP7_75t_L g1208 ( 
.A(n_920),
.Y(n_1208)
);

NOR2x1_ASAP7_75t_L g1209 ( 
.A(n_955),
.B(n_321),
.Y(n_1209)
);

NAND2xp5_ASAP7_75t_L g1210 ( 
.A(n_997),
.B(n_27),
.Y(n_1210)
);

NAND2xp5_ASAP7_75t_SL g1211 ( 
.A(n_1063),
.B(n_533),
.Y(n_1211)
);

A2O1A1Ixp33_ASAP7_75t_L g1212 ( 
.A1(n_965),
.A2(n_533),
.B(n_531),
.C(n_35),
.Y(n_1212)
);

NAND2xp5_ASAP7_75t_SL g1213 ( 
.A(n_1063),
.B(n_1027),
.Y(n_1213)
);

BUFx6f_ASAP7_75t_L g1214 ( 
.A(n_927),
.Y(n_1214)
);

OAI21x1_ASAP7_75t_L g1215 ( 
.A1(n_1204),
.A2(n_1053),
.B(n_1045),
.Y(n_1215)
);

OAI21xp5_ASAP7_75t_SL g1216 ( 
.A1(n_1187),
.A2(n_1179),
.B(n_1201),
.Y(n_1216)
);

A2O1A1Ixp33_ASAP7_75t_L g1217 ( 
.A1(n_1203),
.A2(n_1002),
.B(n_1050),
.C(n_1007),
.Y(n_1217)
);

INVx2_ASAP7_75t_L g1218 ( 
.A(n_1077),
.Y(n_1218)
);

AOI21xp5_ASAP7_75t_L g1219 ( 
.A1(n_1145),
.A2(n_984),
.B(n_1015),
.Y(n_1219)
);

INVx1_ASAP7_75t_L g1220 ( 
.A(n_1091),
.Y(n_1220)
);

NAND2xp5_ASAP7_75t_L g1221 ( 
.A(n_1079),
.B(n_964),
.Y(n_1221)
);

NOR2xp33_ASAP7_75t_L g1222 ( 
.A(n_1072),
.B(n_947),
.Y(n_1222)
);

NOR2x1_ASAP7_75t_L g1223 ( 
.A(n_1163),
.B(n_955),
.Y(n_1223)
);

INVx2_ASAP7_75t_L g1224 ( 
.A(n_1081),
.Y(n_1224)
);

NAND2xp5_ASAP7_75t_L g1225 ( 
.A(n_1090),
.B(n_964),
.Y(n_1225)
);

AOI221x1_ASAP7_75t_L g1226 ( 
.A1(n_1090),
.A2(n_1154),
.B1(n_1212),
.B2(n_1074),
.C(n_1094),
.Y(n_1226)
);

CKINVDCx5p33_ASAP7_75t_R g1227 ( 
.A(n_1109),
.Y(n_1227)
);

INVx8_ASAP7_75t_L g1228 ( 
.A(n_1114),
.Y(n_1228)
);

NAND2xp5_ASAP7_75t_L g1229 ( 
.A(n_1080),
.B(n_959),
.Y(n_1229)
);

AOI21xp5_ASAP7_75t_L g1230 ( 
.A1(n_1148),
.A2(n_1015),
.B(n_984),
.Y(n_1230)
);

A2O1A1Ixp33_ASAP7_75t_L g1231 ( 
.A1(n_1073),
.A2(n_1019),
.B(n_1026),
.C(n_1064),
.Y(n_1231)
);

NOR2xp67_ASAP7_75t_L g1232 ( 
.A(n_1092),
.B(n_980),
.Y(n_1232)
);

AND2x4_ASAP7_75t_L g1233 ( 
.A(n_1200),
.B(n_947),
.Y(n_1233)
);

A2O1A1Ixp33_ASAP7_75t_L g1234 ( 
.A1(n_1206),
.A2(n_1064),
.B(n_1047),
.C(n_1027),
.Y(n_1234)
);

OAI22x1_ASAP7_75t_L g1235 ( 
.A1(n_1170),
.A2(n_1029),
.B1(n_1006),
.B2(n_989),
.Y(n_1235)
);

NAND2xp5_ASAP7_75t_L g1236 ( 
.A(n_1080),
.B(n_959),
.Y(n_1236)
);

INVx2_ASAP7_75t_L g1237 ( 
.A(n_1104),
.Y(n_1237)
);

NAND2xp5_ASAP7_75t_L g1238 ( 
.A(n_1089),
.B(n_935),
.Y(n_1238)
);

NAND2xp5_ASAP7_75t_L g1239 ( 
.A(n_1101),
.B(n_946),
.Y(n_1239)
);

AND2x6_ASAP7_75t_L g1240 ( 
.A(n_1170),
.B(n_975),
.Y(n_1240)
);

AOI21xp5_ASAP7_75t_L g1241 ( 
.A1(n_1168),
.A2(n_984),
.B(n_1015),
.Y(n_1241)
);

NOR2xp33_ASAP7_75t_L g1242 ( 
.A(n_1078),
.B(n_975),
.Y(n_1242)
);

OAI21x1_ASAP7_75t_L g1243 ( 
.A1(n_1152),
.A2(n_960),
.B(n_1034),
.Y(n_1243)
);

A2O1A1Ixp33_ASAP7_75t_L g1244 ( 
.A1(n_1188),
.A2(n_987),
.B(n_1017),
.C(n_1061),
.Y(n_1244)
);

OAI22xp5_ASAP7_75t_L g1245 ( 
.A1(n_1183),
.A2(n_931),
.B1(n_946),
.B2(n_1059),
.Y(n_1245)
);

AOI21xp5_ASAP7_75t_L g1246 ( 
.A1(n_1131),
.A2(n_1015),
.B(n_984),
.Y(n_1246)
);

BUFx6f_ASAP7_75t_L g1247 ( 
.A(n_1200),
.Y(n_1247)
);

INVx2_ASAP7_75t_L g1248 ( 
.A(n_1121),
.Y(n_1248)
);

AOI21xp5_ASAP7_75t_L g1249 ( 
.A1(n_1132),
.A2(n_930),
.B(n_979),
.Y(n_1249)
);

O2A1O1Ixp33_ASAP7_75t_SL g1250 ( 
.A1(n_1103),
.A2(n_913),
.B(n_933),
.C(n_1066),
.Y(n_1250)
);

NOR2xp33_ASAP7_75t_L g1251 ( 
.A(n_1208),
.B(n_1055),
.Y(n_1251)
);

OA21x2_ASAP7_75t_L g1252 ( 
.A1(n_1192),
.A2(n_1048),
.B(n_952),
.Y(n_1252)
);

AOI22xp33_ASAP7_75t_L g1253 ( 
.A1(n_1153),
.A2(n_1048),
.B1(n_1061),
.B2(n_1070),
.Y(n_1253)
);

O2A1O1Ixp33_ASAP7_75t_SL g1254 ( 
.A1(n_1100),
.A2(n_1149),
.B(n_1194),
.C(n_1122),
.Y(n_1254)
);

INVx1_ASAP7_75t_L g1255 ( 
.A(n_1120),
.Y(n_1255)
);

INVx2_ASAP7_75t_L g1256 ( 
.A(n_1130),
.Y(n_1256)
);

INVxp67_ASAP7_75t_SL g1257 ( 
.A(n_1193),
.Y(n_1257)
);

OR2x2_ASAP7_75t_L g1258 ( 
.A(n_1126),
.B(n_1059),
.Y(n_1258)
);

INVxp67_ASAP7_75t_SL g1259 ( 
.A(n_1134),
.Y(n_1259)
);

BUFx6f_ASAP7_75t_L g1260 ( 
.A(n_1096),
.Y(n_1260)
);

BUFx2_ASAP7_75t_L g1261 ( 
.A(n_1133),
.Y(n_1261)
);

OAI21x1_ASAP7_75t_L g1262 ( 
.A1(n_1123),
.A2(n_988),
.B(n_995),
.Y(n_1262)
);

INVxp67_ASAP7_75t_SL g1263 ( 
.A(n_1108),
.Y(n_1263)
);

OAI22x1_ASAP7_75t_L g1264 ( 
.A1(n_1173),
.A2(n_1151),
.B1(n_1128),
.B2(n_1142),
.Y(n_1264)
);

AOI21xp5_ASAP7_75t_L g1265 ( 
.A1(n_1125),
.A2(n_1129),
.B(n_1159),
.Y(n_1265)
);

OAI21x1_ASAP7_75t_L g1266 ( 
.A1(n_1102),
.A2(n_1025),
.B(n_1071),
.Y(n_1266)
);

OAI21xp5_ASAP7_75t_L g1267 ( 
.A1(n_1076),
.A2(n_1056),
.B(n_910),
.Y(n_1267)
);

INVx1_ASAP7_75t_L g1268 ( 
.A(n_1180),
.Y(n_1268)
);

BUFx2_ASAP7_75t_L g1269 ( 
.A(n_1186),
.Y(n_1269)
);

BUFx2_ASAP7_75t_L g1270 ( 
.A(n_1208),
.Y(n_1270)
);

AND2x4_ASAP7_75t_L g1271 ( 
.A(n_1140),
.B(n_980),
.Y(n_1271)
);

NAND2xp5_ASAP7_75t_L g1272 ( 
.A(n_1101),
.B(n_1082),
.Y(n_1272)
);

INVx1_ASAP7_75t_L g1273 ( 
.A(n_1191),
.Y(n_1273)
);

OAI21xp5_ASAP7_75t_L g1274 ( 
.A1(n_1082),
.A2(n_1031),
.B(n_1054),
.Y(n_1274)
);

AO31x2_ASAP7_75t_L g1275 ( 
.A1(n_1195),
.A2(n_1071),
.A3(n_1058),
.B(n_1052),
.Y(n_1275)
);

NOR2xp33_ASAP7_75t_R g1276 ( 
.A(n_1181),
.B(n_930),
.Y(n_1276)
);

INVx1_ASAP7_75t_L g1277 ( 
.A(n_1194),
.Y(n_1277)
);

AOI21xp5_ASAP7_75t_L g1278 ( 
.A1(n_1124),
.A2(n_979),
.B(n_930),
.Y(n_1278)
);

OAI22xp5_ASAP7_75t_L g1279 ( 
.A1(n_1177),
.A2(n_1210),
.B1(n_1088),
.B2(n_1202),
.Y(n_1279)
);

CKINVDCx20_ASAP7_75t_R g1280 ( 
.A(n_1190),
.Y(n_1280)
);

NAND2xp5_ASAP7_75t_L g1281 ( 
.A(n_1115),
.B(n_1036),
.Y(n_1281)
);

NAND3x1_ASAP7_75t_L g1282 ( 
.A(n_1210),
.B(n_1025),
.C(n_933),
.Y(n_1282)
);

INVx2_ASAP7_75t_L g1283 ( 
.A(n_1141),
.Y(n_1283)
);

OA21x2_ASAP7_75t_L g1284 ( 
.A1(n_1093),
.A2(n_1031),
.B(n_1058),
.Y(n_1284)
);

AOI21xp5_ASAP7_75t_L g1285 ( 
.A1(n_1150),
.A2(n_979),
.B(n_1033),
.Y(n_1285)
);

AO32x2_ASAP7_75t_L g1286 ( 
.A1(n_1154),
.A2(n_1039),
.A3(n_993),
.B1(n_1069),
.B2(n_1062),
.Y(n_1286)
);

INVx2_ASAP7_75t_L g1287 ( 
.A(n_1155),
.Y(n_1287)
);

INVx1_ASAP7_75t_L g1288 ( 
.A(n_1156),
.Y(n_1288)
);

AOI21xp5_ASAP7_75t_L g1289 ( 
.A1(n_1207),
.A2(n_999),
.B(n_1069),
.Y(n_1289)
);

OAI21x1_ASAP7_75t_L g1290 ( 
.A1(n_1161),
.A2(n_1052),
.B(n_1069),
.Y(n_1290)
);

NAND2xp5_ASAP7_75t_L g1291 ( 
.A(n_1115),
.B(n_1036),
.Y(n_1291)
);

NAND2xp5_ASAP7_75t_L g1292 ( 
.A(n_1213),
.B(n_1172),
.Y(n_1292)
);

NOR2xp33_ASAP7_75t_L g1293 ( 
.A(n_1105),
.B(n_1063),
.Y(n_1293)
);

NAND2xp5_ASAP7_75t_L g1294 ( 
.A(n_1184),
.B(n_1036),
.Y(n_1294)
);

BUFx6f_ASAP7_75t_L g1295 ( 
.A(n_1096),
.Y(n_1295)
);

AOI21xp5_ASAP7_75t_L g1296 ( 
.A1(n_1139),
.A2(n_999),
.B(n_1000),
.Y(n_1296)
);

BUFx2_ASAP7_75t_L g1297 ( 
.A(n_1197),
.Y(n_1297)
);

NAND2xp5_ASAP7_75t_L g1298 ( 
.A(n_1199),
.B(n_1042),
.Y(n_1298)
);

NAND2xp33_ASAP7_75t_R g1299 ( 
.A(n_1160),
.B(n_1032),
.Y(n_1299)
);

AOI221x1_ASAP7_75t_L g1300 ( 
.A1(n_1135),
.A2(n_1037),
.B1(n_1042),
.B2(n_1000),
.C(n_1063),
.Y(n_1300)
);

AO32x2_ASAP7_75t_L g1301 ( 
.A1(n_1095),
.A2(n_33),
.A3(n_34),
.B1(n_38),
.B2(n_40),
.Y(n_1301)
);

NAND2xp5_ASAP7_75t_L g1302 ( 
.A(n_1112),
.B(n_33),
.Y(n_1302)
);

AOI21xp5_ASAP7_75t_L g1303 ( 
.A1(n_1147),
.A2(n_533),
.B(n_531),
.Y(n_1303)
);

BUFx3_ASAP7_75t_L g1304 ( 
.A(n_1167),
.Y(n_1304)
);

NAND2xp5_ASAP7_75t_SL g1305 ( 
.A(n_1084),
.B(n_1160),
.Y(n_1305)
);

NAND2xp5_ASAP7_75t_SL g1306 ( 
.A(n_1084),
.B(n_533),
.Y(n_1306)
);

AO31x2_ASAP7_75t_L g1307 ( 
.A1(n_1107),
.A2(n_533),
.A3(n_531),
.B(n_115),
.Y(n_1307)
);

OAI21xp5_ASAP7_75t_L g1308 ( 
.A1(n_1085),
.A2(n_531),
.B(n_40),
.Y(n_1308)
);

INVxp67_ASAP7_75t_SL g1309 ( 
.A(n_1112),
.Y(n_1309)
);

AOI21xp33_ASAP7_75t_L g1310 ( 
.A1(n_1143),
.A2(n_38),
.B(n_41),
.Y(n_1310)
);

NAND2xp5_ASAP7_75t_SL g1311 ( 
.A(n_1127),
.B(n_42),
.Y(n_1311)
);

OR2x2_ASAP7_75t_L g1312 ( 
.A(n_1165),
.B(n_45),
.Y(n_1312)
);

AND2x4_ASAP7_75t_L g1313 ( 
.A(n_1114),
.B(n_179),
.Y(n_1313)
);

OAI21x1_ASAP7_75t_L g1314 ( 
.A1(n_1209),
.A2(n_1107),
.B(n_1111),
.Y(n_1314)
);

AOI21xp5_ASAP7_75t_L g1315 ( 
.A1(n_1111),
.A2(n_173),
.B(n_164),
.Y(n_1315)
);

NAND2xp5_ASAP7_75t_L g1316 ( 
.A(n_1127),
.B(n_45),
.Y(n_1316)
);

NAND2xp5_ASAP7_75t_SL g1317 ( 
.A(n_1144),
.B(n_47),
.Y(n_1317)
);

O2A1O1Ixp33_ASAP7_75t_SL g1318 ( 
.A1(n_1118),
.A2(n_49),
.B(n_50),
.C(n_54),
.Y(n_1318)
);

BUFx2_ASAP7_75t_R g1319 ( 
.A(n_1211),
.Y(n_1319)
);

NAND2xp5_ASAP7_75t_SL g1320 ( 
.A(n_1144),
.B(n_49),
.Y(n_1320)
);

NAND2xp5_ASAP7_75t_L g1321 ( 
.A(n_1189),
.B(n_1083),
.Y(n_1321)
);

AO31x2_ASAP7_75t_L g1322 ( 
.A1(n_1099),
.A2(n_1095),
.A3(n_1116),
.B(n_1162),
.Y(n_1322)
);

BUFx2_ASAP7_75t_SL g1323 ( 
.A(n_1097),
.Y(n_1323)
);

NAND2xp5_ASAP7_75t_SL g1324 ( 
.A(n_1189),
.B(n_55),
.Y(n_1324)
);

INVx1_ASAP7_75t_L g1325 ( 
.A(n_1106),
.Y(n_1325)
);

NOR2x1_ASAP7_75t_SL g1326 ( 
.A(n_1114),
.B(n_56),
.Y(n_1326)
);

INVx1_ASAP7_75t_L g1327 ( 
.A(n_1171),
.Y(n_1327)
);

AO22x2_ASAP7_75t_L g1328 ( 
.A1(n_1113),
.A2(n_56),
.B1(n_60),
.B2(n_62),
.Y(n_1328)
);

OAI21xp5_ASAP7_75t_L g1329 ( 
.A1(n_1116),
.A2(n_63),
.B(n_66),
.Y(n_1329)
);

INVx1_ASAP7_75t_SL g1330 ( 
.A(n_1087),
.Y(n_1330)
);

AOI21xp5_ASAP7_75t_L g1331 ( 
.A1(n_1164),
.A2(n_1162),
.B(n_1158),
.Y(n_1331)
);

BUFx2_ASAP7_75t_L g1332 ( 
.A(n_1087),
.Y(n_1332)
);

INVx1_ASAP7_75t_L g1333 ( 
.A(n_1171),
.Y(n_1333)
);

NAND2xp5_ASAP7_75t_L g1334 ( 
.A(n_1087),
.B(n_63),
.Y(n_1334)
);

AO32x2_ASAP7_75t_L g1335 ( 
.A1(n_1169),
.A2(n_66),
.A3(n_67),
.B1(n_69),
.B2(n_73),
.Y(n_1335)
);

NAND2xp5_ASAP7_75t_SL g1336 ( 
.A(n_1110),
.B(n_67),
.Y(n_1336)
);

BUFx3_ASAP7_75t_L g1337 ( 
.A(n_1075),
.Y(n_1337)
);

NAND2xp5_ASAP7_75t_L g1338 ( 
.A(n_1110),
.B(n_69),
.Y(n_1338)
);

NAND2xp5_ASAP7_75t_L g1339 ( 
.A(n_1110),
.B(n_73),
.Y(n_1339)
);

AOI21xp33_ASAP7_75t_L g1340 ( 
.A1(n_1098),
.A2(n_76),
.B(n_77),
.Y(n_1340)
);

AO21x1_ASAP7_75t_L g1341 ( 
.A1(n_1178),
.A2(n_79),
.B(n_117),
.Y(n_1341)
);

AOI21xp5_ASAP7_75t_L g1342 ( 
.A1(n_1117),
.A2(n_123),
.B(n_126),
.Y(n_1342)
);

AND2x2_ASAP7_75t_L g1343 ( 
.A(n_1146),
.B(n_158),
.Y(n_1343)
);

OAI21x1_ASAP7_75t_L g1344 ( 
.A1(n_1086),
.A2(n_137),
.B(n_138),
.Y(n_1344)
);

AOI21xp5_ASAP7_75t_L g1345 ( 
.A1(n_1119),
.A2(n_142),
.B(n_143),
.Y(n_1345)
);

AO31x2_ASAP7_75t_L g1346 ( 
.A1(n_1157),
.A2(n_1166),
.A3(n_1175),
.B(n_1176),
.Y(n_1346)
);

BUFx12f_ASAP7_75t_L g1347 ( 
.A(n_1174),
.Y(n_1347)
);

AOI21xp5_ASAP7_75t_L g1348 ( 
.A1(n_1171),
.A2(n_1214),
.B(n_1174),
.Y(n_1348)
);

INVx1_ASAP7_75t_L g1349 ( 
.A(n_1198),
.Y(n_1349)
);

INVx2_ASAP7_75t_L g1350 ( 
.A(n_1174),
.Y(n_1350)
);

INVx2_ASAP7_75t_L g1351 ( 
.A(n_1214),
.Y(n_1351)
);

AND2x6_ASAP7_75t_L g1352 ( 
.A(n_1214),
.B(n_1196),
.Y(n_1352)
);

AND2x2_ASAP7_75t_L g1353 ( 
.A(n_1146),
.B(n_1169),
.Y(n_1353)
);

AOI21x1_ASAP7_75t_L g1354 ( 
.A1(n_1176),
.A2(n_1182),
.B(n_1185),
.Y(n_1354)
);

NAND2xp5_ASAP7_75t_L g1355 ( 
.A(n_1182),
.B(n_1136),
.Y(n_1355)
);

AND2x2_ASAP7_75t_L g1356 ( 
.A(n_1137),
.B(n_1205),
.Y(n_1356)
);

O2A1O1Ixp5_ASAP7_75t_SL g1357 ( 
.A1(n_1118),
.A2(n_1090),
.B(n_1154),
.C(n_827),
.Y(n_1357)
);

O2A1O1Ixp5_ASAP7_75t_L g1358 ( 
.A1(n_1090),
.A2(n_747),
.B(n_593),
.C(n_992),
.Y(n_1358)
);

NAND2x1_ASAP7_75t_L g1359 ( 
.A(n_1097),
.B(n_1127),
.Y(n_1359)
);

AO31x2_ASAP7_75t_L g1360 ( 
.A1(n_1145),
.A2(n_1030),
.A3(n_1168),
.B(n_1094),
.Y(n_1360)
);

INVx3_ASAP7_75t_L g1361 ( 
.A(n_1097),
.Y(n_1361)
);

OAI21xp5_ASAP7_75t_SL g1362 ( 
.A1(n_1187),
.A2(n_747),
.B(n_974),
.Y(n_1362)
);

OAI21x1_ASAP7_75t_L g1363 ( 
.A1(n_1204),
.A2(n_1152),
.B(n_1138),
.Y(n_1363)
);

NAND2xp5_ASAP7_75t_L g1364 ( 
.A(n_1079),
.B(n_939),
.Y(n_1364)
);

NOR2xp33_ASAP7_75t_L g1365 ( 
.A(n_1362),
.B(n_1355),
.Y(n_1365)
);

NAND2xp5_ASAP7_75t_L g1366 ( 
.A(n_1259),
.B(n_1257),
.Y(n_1366)
);

OR2x6_ASAP7_75t_L g1367 ( 
.A(n_1228),
.B(n_1313),
.Y(n_1367)
);

O2A1O1Ixp5_ASAP7_75t_L g1368 ( 
.A1(n_1358),
.A2(n_1308),
.B(n_1329),
.C(n_1279),
.Y(n_1368)
);

OAI21xp5_ASAP7_75t_L g1369 ( 
.A1(n_1355),
.A2(n_1329),
.B(n_1362),
.Y(n_1369)
);

AND2x2_ASAP7_75t_L g1370 ( 
.A(n_1222),
.B(n_1353),
.Y(n_1370)
);

HB1xp67_ASAP7_75t_L g1371 ( 
.A(n_1360),
.Y(n_1371)
);

AND2x6_ASAP7_75t_L g1372 ( 
.A(n_1313),
.B(n_1225),
.Y(n_1372)
);

OAI22xp33_ASAP7_75t_L g1373 ( 
.A1(n_1225),
.A2(n_1216),
.B1(n_1364),
.B2(n_1226),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_1220),
.Y(n_1374)
);

AND2x2_ASAP7_75t_L g1375 ( 
.A(n_1233),
.B(n_1263),
.Y(n_1375)
);

INVx3_ASAP7_75t_L g1376 ( 
.A(n_1347),
.Y(n_1376)
);

OA21x2_ASAP7_75t_L g1377 ( 
.A1(n_1308),
.A2(n_1331),
.B(n_1243),
.Y(n_1377)
);

OAI21x1_ASAP7_75t_L g1378 ( 
.A1(n_1219),
.A2(n_1215),
.B(n_1241),
.Y(n_1378)
);

INVx1_ASAP7_75t_L g1379 ( 
.A(n_1255),
.Y(n_1379)
);

INVx2_ASAP7_75t_L g1380 ( 
.A(n_1224),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_1268),
.Y(n_1381)
);

OAI21x1_ASAP7_75t_L g1382 ( 
.A1(n_1278),
.A2(n_1249),
.B(n_1246),
.Y(n_1382)
);

INVx1_ASAP7_75t_L g1383 ( 
.A(n_1273),
.Y(n_1383)
);

NAND3xp33_ASAP7_75t_L g1384 ( 
.A(n_1279),
.B(n_1216),
.C(n_1234),
.Y(n_1384)
);

NOR2xp33_ASAP7_75t_L g1385 ( 
.A(n_1242),
.B(n_1251),
.Y(n_1385)
);

OR2x6_ASAP7_75t_L g1386 ( 
.A(n_1228),
.B(n_1348),
.Y(n_1386)
);

INVx4_ASAP7_75t_SL g1387 ( 
.A(n_1240),
.Y(n_1387)
);

INVx2_ASAP7_75t_L g1388 ( 
.A(n_1237),
.Y(n_1388)
);

O2A1O1Ixp33_ASAP7_75t_SL g1389 ( 
.A1(n_1231),
.A2(n_1364),
.B(n_1217),
.C(n_1244),
.Y(n_1389)
);

INVx3_ASAP7_75t_L g1390 ( 
.A(n_1233),
.Y(n_1390)
);

AND2x4_ASAP7_75t_L g1391 ( 
.A(n_1309),
.B(n_1305),
.Y(n_1391)
);

CKINVDCx11_ASAP7_75t_R g1392 ( 
.A(n_1280),
.Y(n_1392)
);

AOI22xp33_ASAP7_75t_L g1393 ( 
.A1(n_1349),
.A2(n_1328),
.B1(n_1343),
.B2(n_1245),
.Y(n_1393)
);

AOI22xp5_ASAP7_75t_L g1394 ( 
.A1(n_1240),
.A2(n_1352),
.B1(n_1299),
.B2(n_1328),
.Y(n_1394)
);

INVx1_ASAP7_75t_L g1395 ( 
.A(n_1288),
.Y(n_1395)
);

INVx1_ASAP7_75t_L g1396 ( 
.A(n_1248),
.Y(n_1396)
);

O2A1O1Ixp33_ASAP7_75t_SL g1397 ( 
.A1(n_1316),
.A2(n_1359),
.B(n_1267),
.C(n_1340),
.Y(n_1397)
);

OAI22xp5_ASAP7_75t_L g1398 ( 
.A1(n_1258),
.A2(n_1356),
.B1(n_1277),
.B2(n_1312),
.Y(n_1398)
);

INVx1_ASAP7_75t_L g1399 ( 
.A(n_1256),
.Y(n_1399)
);

OA21x2_ASAP7_75t_L g1400 ( 
.A1(n_1314),
.A2(n_1266),
.B(n_1262),
.Y(n_1400)
);

A2O1A1Ixp33_ASAP7_75t_L g1401 ( 
.A1(n_1340),
.A2(n_1310),
.B(n_1245),
.C(n_1315),
.Y(n_1401)
);

AO21x2_ASAP7_75t_L g1402 ( 
.A1(n_1272),
.A2(n_1238),
.B(n_1274),
.Y(n_1402)
);

BUFx2_ASAP7_75t_L g1403 ( 
.A(n_1276),
.Y(n_1403)
);

INVx1_ASAP7_75t_SL g1404 ( 
.A(n_1269),
.Y(n_1404)
);

NOR2xp33_ASAP7_75t_L g1405 ( 
.A(n_1293),
.B(n_1302),
.Y(n_1405)
);

INVx1_ASAP7_75t_L g1406 ( 
.A(n_1283),
.Y(n_1406)
);

OAI21x1_ASAP7_75t_L g1407 ( 
.A1(n_1230),
.A2(n_1289),
.B(n_1285),
.Y(n_1407)
);

OAI21xp5_ASAP7_75t_L g1408 ( 
.A1(n_1357),
.A2(n_1282),
.B(n_1310),
.Y(n_1408)
);

OAI22xp5_ASAP7_75t_L g1409 ( 
.A1(n_1253),
.A2(n_1354),
.B1(n_1302),
.B2(n_1321),
.Y(n_1409)
);

INVx2_ASAP7_75t_L g1410 ( 
.A(n_1287),
.Y(n_1410)
);

BUFx12f_ASAP7_75t_L g1411 ( 
.A(n_1227),
.Y(n_1411)
);

AO21x2_ASAP7_75t_L g1412 ( 
.A1(n_1272),
.A2(n_1238),
.B(n_1274),
.Y(n_1412)
);

AOI22xp33_ASAP7_75t_L g1413 ( 
.A1(n_1229),
.A2(n_1236),
.B1(n_1264),
.B2(n_1221),
.Y(n_1413)
);

OAI22xp5_ASAP7_75t_L g1414 ( 
.A1(n_1321),
.A2(n_1270),
.B1(n_1261),
.B2(n_1325),
.Y(n_1414)
);

A2O1A1Ixp33_ASAP7_75t_L g1415 ( 
.A1(n_1221),
.A2(n_1229),
.B(n_1236),
.C(n_1342),
.Y(n_1415)
);

HB1xp67_ASAP7_75t_L g1416 ( 
.A(n_1360),
.Y(n_1416)
);

OAI22xp5_ASAP7_75t_L g1417 ( 
.A1(n_1232),
.A2(n_1311),
.B1(n_1324),
.B2(n_1320),
.Y(n_1417)
);

O2A1O1Ixp33_ASAP7_75t_L g1418 ( 
.A1(n_1317),
.A2(n_1336),
.B(n_1318),
.C(n_1254),
.Y(n_1418)
);

AOI21xp33_ASAP7_75t_L g1419 ( 
.A1(n_1239),
.A2(n_1252),
.B(n_1235),
.Y(n_1419)
);

AOI22xp33_ASAP7_75t_SL g1420 ( 
.A1(n_1304),
.A2(n_1326),
.B1(n_1240),
.B2(n_1301),
.Y(n_1420)
);

O2A1O1Ixp33_ASAP7_75t_L g1421 ( 
.A1(n_1334),
.A2(n_1339),
.B(n_1338),
.C(n_1345),
.Y(n_1421)
);

OAI22xp33_ASAP7_75t_L g1422 ( 
.A1(n_1301),
.A2(n_1239),
.B1(n_1339),
.B2(n_1334),
.Y(n_1422)
);

AOI22xp33_ASAP7_75t_L g1423 ( 
.A1(n_1352),
.A2(n_1252),
.B1(n_1341),
.B2(n_1292),
.Y(n_1423)
);

BUFx3_ASAP7_75t_L g1424 ( 
.A(n_1352),
.Y(n_1424)
);

CKINVDCx8_ASAP7_75t_R g1425 ( 
.A(n_1352),
.Y(n_1425)
);

NAND2xp5_ASAP7_75t_SL g1426 ( 
.A(n_1281),
.B(n_1291),
.Y(n_1426)
);

HB1xp67_ASAP7_75t_L g1427 ( 
.A(n_1360),
.Y(n_1427)
);

INVx2_ASAP7_75t_L g1428 ( 
.A(n_1292),
.Y(n_1428)
);

AOI22x1_ASAP7_75t_L g1429 ( 
.A1(n_1361),
.A2(n_1323),
.B1(n_1297),
.B2(n_1332),
.Y(n_1429)
);

AO31x2_ASAP7_75t_L g1430 ( 
.A1(n_1300),
.A2(n_1281),
.A3(n_1291),
.B(n_1298),
.Y(n_1430)
);

NAND3xp33_ASAP7_75t_L g1431 ( 
.A(n_1338),
.B(n_1223),
.C(n_1306),
.Y(n_1431)
);

AND2x2_ASAP7_75t_L g1432 ( 
.A(n_1247),
.B(n_1271),
.Y(n_1432)
);

NAND3xp33_ASAP7_75t_L g1433 ( 
.A(n_1327),
.B(n_1333),
.C(n_1271),
.Y(n_1433)
);

OAI21x1_ASAP7_75t_L g1434 ( 
.A1(n_1284),
.A2(n_1303),
.B(n_1344),
.Y(n_1434)
);

BUFx6f_ASAP7_75t_L g1435 ( 
.A(n_1247),
.Y(n_1435)
);

OR2x6_ASAP7_75t_L g1436 ( 
.A(n_1296),
.B(n_1295),
.Y(n_1436)
);

NOR2xp67_ASAP7_75t_L g1437 ( 
.A(n_1361),
.B(n_1351),
.Y(n_1437)
);

INVx1_ASAP7_75t_L g1438 ( 
.A(n_1294),
.Y(n_1438)
);

NAND2x1_ASAP7_75t_L g1439 ( 
.A(n_1284),
.B(n_1350),
.Y(n_1439)
);

BUFx3_ASAP7_75t_L g1440 ( 
.A(n_1260),
.Y(n_1440)
);

INVx1_ASAP7_75t_SL g1441 ( 
.A(n_1319),
.Y(n_1441)
);

INVx5_ASAP7_75t_SL g1442 ( 
.A(n_1260),
.Y(n_1442)
);

AOI22xp33_ASAP7_75t_SL g1443 ( 
.A1(n_1301),
.A2(n_1335),
.B1(n_1286),
.B2(n_1337),
.Y(n_1443)
);

INVxp67_ASAP7_75t_L g1444 ( 
.A(n_1330),
.Y(n_1444)
);

AOI21xp5_ASAP7_75t_L g1445 ( 
.A1(n_1250),
.A2(n_1330),
.B(n_1286),
.Y(n_1445)
);

OAI21x1_ASAP7_75t_L g1446 ( 
.A1(n_1275),
.A2(n_1307),
.B(n_1322),
.Y(n_1446)
);

INVx1_ASAP7_75t_L g1447 ( 
.A(n_1335),
.Y(n_1447)
);

AOI221xp5_ASAP7_75t_SL g1448 ( 
.A1(n_1335),
.A2(n_1260),
.B1(n_1295),
.B2(n_1346),
.C(n_1307),
.Y(n_1448)
);

O2A1O1Ixp33_ASAP7_75t_SL g1449 ( 
.A1(n_1346),
.A2(n_1286),
.B(n_1307),
.C(n_1322),
.Y(n_1449)
);

OAI22xp5_ASAP7_75t_L g1450 ( 
.A1(n_1295),
.A2(n_1346),
.B1(n_1322),
.B2(n_1275),
.Y(n_1450)
);

NAND3xp33_ASAP7_75t_SL g1451 ( 
.A(n_1275),
.B(n_1358),
.C(n_747),
.Y(n_1451)
);

O2A1O1Ixp33_ASAP7_75t_L g1452 ( 
.A1(n_1358),
.A2(n_747),
.B(n_593),
.C(n_1279),
.Y(n_1452)
);

AND2x2_ASAP7_75t_L g1453 ( 
.A(n_1222),
.B(n_1072),
.Y(n_1453)
);

AOI21xp5_ASAP7_75t_L g1454 ( 
.A1(n_1358),
.A2(n_1148),
.B(n_1145),
.Y(n_1454)
);

OAI21x1_ASAP7_75t_L g1455 ( 
.A1(n_1363),
.A2(n_1265),
.B(n_1290),
.Y(n_1455)
);

OAI21x1_ASAP7_75t_SL g1456 ( 
.A1(n_1329),
.A2(n_1355),
.B(n_1279),
.Y(n_1456)
);

AND2x2_ASAP7_75t_L g1457 ( 
.A(n_1222),
.B(n_1072),
.Y(n_1457)
);

NOR2xp33_ASAP7_75t_L g1458 ( 
.A(n_1362),
.B(n_747),
.Y(n_1458)
);

BUFx3_ASAP7_75t_L g1459 ( 
.A(n_1347),
.Y(n_1459)
);

INVx1_ASAP7_75t_L g1460 ( 
.A(n_1220),
.Y(n_1460)
);

NAND2xp5_ASAP7_75t_L g1461 ( 
.A(n_1259),
.B(n_1021),
.Y(n_1461)
);

OAI21x1_ASAP7_75t_L g1462 ( 
.A1(n_1363),
.A2(n_1265),
.B(n_1290),
.Y(n_1462)
);

OA21x2_ASAP7_75t_L g1463 ( 
.A1(n_1265),
.A2(n_1363),
.B(n_1226),
.Y(n_1463)
);

OR2x2_ASAP7_75t_L g1464 ( 
.A(n_1257),
.B(n_1258),
.Y(n_1464)
);

AND2x4_ASAP7_75t_L g1465 ( 
.A(n_1309),
.B(n_1233),
.Y(n_1465)
);

NOR3xp33_ASAP7_75t_L g1466 ( 
.A(n_1358),
.B(n_747),
.C(n_1216),
.Y(n_1466)
);

AOI22xp5_ASAP7_75t_L g1467 ( 
.A1(n_1362),
.A2(n_747),
.B1(n_1023),
.B2(n_1021),
.Y(n_1467)
);

OAI21x1_ASAP7_75t_L g1468 ( 
.A1(n_1363),
.A2(n_1265),
.B(n_1290),
.Y(n_1468)
);

INVx5_ASAP7_75t_L g1469 ( 
.A(n_1352),
.Y(n_1469)
);

NAND2x1p5_ASAP7_75t_L g1470 ( 
.A(n_1313),
.B(n_1337),
.Y(n_1470)
);

OA21x2_ASAP7_75t_L g1471 ( 
.A1(n_1265),
.A2(n_1363),
.B(n_1226),
.Y(n_1471)
);

INVx1_ASAP7_75t_L g1472 ( 
.A(n_1220),
.Y(n_1472)
);

NAND2x1p5_ASAP7_75t_L g1473 ( 
.A(n_1313),
.B(n_1337),
.Y(n_1473)
);

HB1xp67_ASAP7_75t_L g1474 ( 
.A(n_1360),
.Y(n_1474)
);

AOI22xp33_ASAP7_75t_L g1475 ( 
.A1(n_1353),
.A2(n_974),
.B1(n_671),
.B2(n_785),
.Y(n_1475)
);

OAI21x1_ASAP7_75t_L g1476 ( 
.A1(n_1363),
.A2(n_1265),
.B(n_1290),
.Y(n_1476)
);

INVx1_ASAP7_75t_L g1477 ( 
.A(n_1220),
.Y(n_1477)
);

AOI22xp33_ASAP7_75t_SL g1478 ( 
.A1(n_1353),
.A2(n_785),
.B1(n_815),
.B2(n_671),
.Y(n_1478)
);

OAI21x1_ASAP7_75t_L g1479 ( 
.A1(n_1363),
.A2(n_1265),
.B(n_1290),
.Y(n_1479)
);

OAI21xp5_ASAP7_75t_L g1480 ( 
.A1(n_1358),
.A2(n_747),
.B(n_593),
.Y(n_1480)
);

OAI21x1_ASAP7_75t_L g1481 ( 
.A1(n_1363),
.A2(n_1265),
.B(n_1290),
.Y(n_1481)
);

OA21x2_ASAP7_75t_L g1482 ( 
.A1(n_1265),
.A2(n_1363),
.B(n_1226),
.Y(n_1482)
);

AND2x2_ASAP7_75t_L g1483 ( 
.A(n_1222),
.B(n_1072),
.Y(n_1483)
);

NOR2xp67_ASAP7_75t_L g1484 ( 
.A(n_1222),
.B(n_973),
.Y(n_1484)
);

OAI21x1_ASAP7_75t_L g1485 ( 
.A1(n_1363),
.A2(n_1265),
.B(n_1290),
.Y(n_1485)
);

NOR2xp67_ASAP7_75t_L g1486 ( 
.A(n_1222),
.B(n_973),
.Y(n_1486)
);

BUFx12f_ASAP7_75t_L g1487 ( 
.A(n_1227),
.Y(n_1487)
);

BUFx3_ASAP7_75t_L g1488 ( 
.A(n_1347),
.Y(n_1488)
);

INVx1_ASAP7_75t_L g1489 ( 
.A(n_1220),
.Y(n_1489)
);

CKINVDCx11_ASAP7_75t_R g1490 ( 
.A(n_1280),
.Y(n_1490)
);

INVx2_ASAP7_75t_L g1491 ( 
.A(n_1218),
.Y(n_1491)
);

NAND2xp5_ASAP7_75t_L g1492 ( 
.A(n_1259),
.B(n_1021),
.Y(n_1492)
);

BUFx3_ASAP7_75t_L g1493 ( 
.A(n_1347),
.Y(n_1493)
);

OAI211xp5_ASAP7_75t_SL g1494 ( 
.A1(n_1358),
.A2(n_593),
.B(n_747),
.C(n_571),
.Y(n_1494)
);

INVx2_ASAP7_75t_L g1495 ( 
.A(n_1218),
.Y(n_1495)
);

AOI22xp33_ASAP7_75t_L g1496 ( 
.A1(n_1353),
.A2(n_974),
.B1(n_671),
.B2(n_785),
.Y(n_1496)
);

AOI22xp33_ASAP7_75t_L g1497 ( 
.A1(n_1353),
.A2(n_974),
.B1(n_671),
.B2(n_785),
.Y(n_1497)
);

AOI222xp33_ASAP7_75t_SL g1498 ( 
.A1(n_1279),
.A2(n_562),
.B1(n_671),
.B2(n_534),
.C1(n_519),
.C2(n_385),
.Y(n_1498)
);

OAI21x1_ASAP7_75t_L g1499 ( 
.A1(n_1363),
.A2(n_1265),
.B(n_1290),
.Y(n_1499)
);

OAI21x1_ASAP7_75t_L g1500 ( 
.A1(n_1363),
.A2(n_1265),
.B(n_1290),
.Y(n_1500)
);

INVx1_ASAP7_75t_L g1501 ( 
.A(n_1220),
.Y(n_1501)
);

OAI21x1_ASAP7_75t_L g1502 ( 
.A1(n_1363),
.A2(n_1265),
.B(n_1290),
.Y(n_1502)
);

INVx3_ASAP7_75t_L g1503 ( 
.A(n_1347),
.Y(n_1503)
);

OAI21x1_ASAP7_75t_L g1504 ( 
.A1(n_1363),
.A2(n_1265),
.B(n_1290),
.Y(n_1504)
);

OAI21xp5_ASAP7_75t_L g1505 ( 
.A1(n_1358),
.A2(n_747),
.B(n_593),
.Y(n_1505)
);

NAND2xp5_ASAP7_75t_L g1506 ( 
.A(n_1259),
.B(n_1021),
.Y(n_1506)
);

BUFx6f_ASAP7_75t_L g1507 ( 
.A(n_1228),
.Y(n_1507)
);

OA21x2_ASAP7_75t_L g1508 ( 
.A1(n_1265),
.A2(n_1363),
.B(n_1226),
.Y(n_1508)
);

AOI22xp33_ASAP7_75t_SL g1509 ( 
.A1(n_1353),
.A2(n_785),
.B1(n_815),
.B2(n_671),
.Y(n_1509)
);

BUFx6f_ASAP7_75t_L g1510 ( 
.A(n_1228),
.Y(n_1510)
);

NOR2xp33_ASAP7_75t_L g1511 ( 
.A(n_1362),
.B(n_747),
.Y(n_1511)
);

OR2x2_ASAP7_75t_L g1512 ( 
.A(n_1257),
.B(n_1258),
.Y(n_1512)
);

OR2x2_ASAP7_75t_L g1513 ( 
.A(n_1257),
.B(n_1258),
.Y(n_1513)
);

AO31x2_ASAP7_75t_L g1514 ( 
.A1(n_1245),
.A2(n_1331),
.A3(n_1226),
.B(n_1231),
.Y(n_1514)
);

OAI22xp5_ASAP7_75t_L g1515 ( 
.A1(n_1355),
.A2(n_747),
.B1(n_1023),
.B2(n_1021),
.Y(n_1515)
);

NAND2x1p5_ASAP7_75t_L g1516 ( 
.A(n_1313),
.B(n_1337),
.Y(n_1516)
);

INVx2_ASAP7_75t_SL g1517 ( 
.A(n_1276),
.Y(n_1517)
);

NOR2xp33_ASAP7_75t_L g1518 ( 
.A(n_1362),
.B(n_747),
.Y(n_1518)
);

NOR2x1_ASAP7_75t_SL g1519 ( 
.A(n_1367),
.B(n_1469),
.Y(n_1519)
);

AND2x2_ASAP7_75t_L g1520 ( 
.A(n_1375),
.B(n_1370),
.Y(n_1520)
);

INVx2_ASAP7_75t_SL g1521 ( 
.A(n_1459),
.Y(n_1521)
);

OAI22xp5_ASAP7_75t_L g1522 ( 
.A1(n_1467),
.A2(n_1511),
.B1(n_1458),
.B2(n_1518),
.Y(n_1522)
);

BUFx6f_ASAP7_75t_L g1523 ( 
.A(n_1367),
.Y(n_1523)
);

O2A1O1Ixp33_ASAP7_75t_L g1524 ( 
.A1(n_1458),
.A2(n_1518),
.B(n_1511),
.C(n_1452),
.Y(n_1524)
);

OA21x2_ASAP7_75t_L g1525 ( 
.A1(n_1448),
.A2(n_1446),
.B(n_1454),
.Y(n_1525)
);

AOI21x1_ASAP7_75t_SL g1526 ( 
.A1(n_1461),
.A2(n_1506),
.B(n_1492),
.Y(n_1526)
);

HB1xp67_ASAP7_75t_L g1527 ( 
.A(n_1371),
.Y(n_1527)
);

AND2x2_ASAP7_75t_L g1528 ( 
.A(n_1405),
.B(n_1385),
.Y(n_1528)
);

OR2x2_ASAP7_75t_L g1529 ( 
.A(n_1464),
.B(n_1512),
.Y(n_1529)
);

O2A1O1Ixp33_ASAP7_75t_L g1530 ( 
.A1(n_1515),
.A2(n_1505),
.B(n_1480),
.C(n_1466),
.Y(n_1530)
);

O2A1O1Ixp33_ASAP7_75t_L g1531 ( 
.A1(n_1466),
.A2(n_1494),
.B(n_1384),
.C(n_1456),
.Y(n_1531)
);

O2A1O1Ixp33_ASAP7_75t_L g1532 ( 
.A1(n_1494),
.A2(n_1369),
.B(n_1365),
.C(n_1373),
.Y(n_1532)
);

AND2x2_ASAP7_75t_L g1533 ( 
.A(n_1405),
.B(n_1385),
.Y(n_1533)
);

OAI22xp5_ASAP7_75t_L g1534 ( 
.A1(n_1478),
.A2(n_1509),
.B1(n_1497),
.B2(n_1496),
.Y(n_1534)
);

HB1xp67_ASAP7_75t_L g1535 ( 
.A(n_1371),
.Y(n_1535)
);

AND2x2_ASAP7_75t_L g1536 ( 
.A(n_1453),
.B(n_1457),
.Y(n_1536)
);

AND2x4_ASAP7_75t_L g1537 ( 
.A(n_1469),
.B(n_1387),
.Y(n_1537)
);

INVx2_ASAP7_75t_L g1538 ( 
.A(n_1439),
.Y(n_1538)
);

AOI21xp5_ASAP7_75t_L g1539 ( 
.A1(n_1401),
.A2(n_1389),
.B(n_1397),
.Y(n_1539)
);

AND2x4_ASAP7_75t_L g1540 ( 
.A(n_1387),
.B(n_1424),
.Y(n_1540)
);

O2A1O1Ixp33_ASAP7_75t_L g1541 ( 
.A1(n_1373),
.A2(n_1389),
.B(n_1368),
.C(n_1401),
.Y(n_1541)
);

AND2x4_ASAP7_75t_L g1542 ( 
.A(n_1424),
.B(n_1372),
.Y(n_1542)
);

A2O1A1Ixp33_ASAP7_75t_L g1543 ( 
.A1(n_1368),
.A2(n_1420),
.B(n_1478),
.C(n_1509),
.Y(n_1543)
);

AND2x2_ASAP7_75t_SL g1544 ( 
.A(n_1393),
.B(n_1475),
.Y(n_1544)
);

NAND2xp5_ASAP7_75t_L g1545 ( 
.A(n_1513),
.B(n_1483),
.Y(n_1545)
);

O2A1O1Ixp33_ASAP7_75t_L g1546 ( 
.A1(n_1397),
.A2(n_1451),
.B(n_1418),
.C(n_1421),
.Y(n_1546)
);

O2A1O1Ixp33_ASAP7_75t_L g1547 ( 
.A1(n_1451),
.A2(n_1417),
.B(n_1398),
.C(n_1409),
.Y(n_1547)
);

OAI22xp5_ASAP7_75t_L g1548 ( 
.A1(n_1475),
.A2(n_1497),
.B1(n_1496),
.B2(n_1420),
.Y(n_1548)
);

NAND2xp5_ASAP7_75t_L g1549 ( 
.A(n_1404),
.B(n_1379),
.Y(n_1549)
);

OR2x2_ASAP7_75t_L g1550 ( 
.A(n_1381),
.B(n_1383),
.Y(n_1550)
);

AOI21x1_ASAP7_75t_SL g1551 ( 
.A1(n_1416),
.A2(n_1474),
.B(n_1427),
.Y(n_1551)
);

OAI22xp5_ASAP7_75t_L g1552 ( 
.A1(n_1393),
.A2(n_1394),
.B1(n_1486),
.B2(n_1484),
.Y(n_1552)
);

AOI21xp5_ASAP7_75t_SL g1553 ( 
.A1(n_1415),
.A2(n_1473),
.B(n_1470),
.Y(n_1553)
);

NAND2xp5_ASAP7_75t_L g1554 ( 
.A(n_1460),
.B(n_1472),
.Y(n_1554)
);

AOI21x1_ASAP7_75t_SL g1555 ( 
.A1(n_1416),
.A2(n_1427),
.B(n_1474),
.Y(n_1555)
);

INVx1_ASAP7_75t_L g1556 ( 
.A(n_1477),
.Y(n_1556)
);

A2O1A1Ixp33_ASAP7_75t_SL g1557 ( 
.A1(n_1408),
.A2(n_1376),
.B(n_1503),
.C(n_1423),
.Y(n_1557)
);

NAND2xp5_ASAP7_75t_L g1558 ( 
.A(n_1489),
.B(n_1501),
.Y(n_1558)
);

OAI22xp5_ASAP7_75t_L g1559 ( 
.A1(n_1425),
.A2(n_1414),
.B1(n_1413),
.B2(n_1443),
.Y(n_1559)
);

OR2x2_ASAP7_75t_L g1560 ( 
.A(n_1426),
.B(n_1438),
.Y(n_1560)
);

O2A1O1Ixp5_ASAP7_75t_L g1561 ( 
.A1(n_1422),
.A2(n_1415),
.B(n_1445),
.C(n_1426),
.Y(n_1561)
);

BUFx3_ASAP7_75t_L g1562 ( 
.A(n_1459),
.Y(n_1562)
);

O2A1O1Ixp33_ASAP7_75t_L g1563 ( 
.A1(n_1422),
.A2(n_1449),
.B(n_1423),
.C(n_1431),
.Y(n_1563)
);

CKINVDCx5p33_ASAP7_75t_R g1564 ( 
.A(n_1392),
.Y(n_1564)
);

INVx1_ASAP7_75t_L g1565 ( 
.A(n_1395),
.Y(n_1565)
);

OAI22xp5_ASAP7_75t_L g1566 ( 
.A1(n_1413),
.A2(n_1443),
.B1(n_1473),
.B2(n_1470),
.Y(n_1566)
);

HB1xp67_ASAP7_75t_L g1567 ( 
.A(n_1400),
.Y(n_1567)
);

AND2x2_ASAP7_75t_L g1568 ( 
.A(n_1432),
.B(n_1444),
.Y(n_1568)
);

NAND2xp5_ASAP7_75t_L g1569 ( 
.A(n_1444),
.B(n_1428),
.Y(n_1569)
);

NAND2xp5_ASAP7_75t_L g1570 ( 
.A(n_1465),
.B(n_1402),
.Y(n_1570)
);

OAI22xp5_ASAP7_75t_L g1571 ( 
.A1(n_1516),
.A2(n_1517),
.B1(n_1488),
.B2(n_1493),
.Y(n_1571)
);

O2A1O1Ixp5_ASAP7_75t_L g1572 ( 
.A1(n_1450),
.A2(n_1419),
.B(n_1447),
.C(n_1391),
.Y(n_1572)
);

HB1xp67_ASAP7_75t_L g1573 ( 
.A(n_1400),
.Y(n_1573)
);

INVx1_ASAP7_75t_L g1574 ( 
.A(n_1396),
.Y(n_1574)
);

AND2x2_ASAP7_75t_L g1575 ( 
.A(n_1390),
.B(n_1441),
.Y(n_1575)
);

AOI21xp5_ASAP7_75t_L g1576 ( 
.A1(n_1449),
.A2(n_1377),
.B(n_1508),
.Y(n_1576)
);

O2A1O1Ixp33_ASAP7_75t_L g1577 ( 
.A1(n_1498),
.A2(n_1503),
.B(n_1376),
.C(n_1516),
.Y(n_1577)
);

AND2x2_ASAP7_75t_L g1578 ( 
.A(n_1435),
.B(n_1372),
.Y(n_1578)
);

AND2x4_ASAP7_75t_L g1579 ( 
.A(n_1372),
.B(n_1386),
.Y(n_1579)
);

OAI22xp5_ASAP7_75t_L g1580 ( 
.A1(n_1488),
.A2(n_1493),
.B1(n_1429),
.B2(n_1433),
.Y(n_1580)
);

INVxp67_ASAP7_75t_L g1581 ( 
.A(n_1402),
.Y(n_1581)
);

NAND2xp5_ASAP7_75t_L g1582 ( 
.A(n_1412),
.B(n_1372),
.Y(n_1582)
);

OA21x2_ASAP7_75t_L g1583 ( 
.A1(n_1455),
.A2(n_1485),
.B(n_1481),
.Y(n_1583)
);

OR2x2_ASAP7_75t_L g1584 ( 
.A(n_1430),
.B(n_1412),
.Y(n_1584)
);

NAND2xp5_ASAP7_75t_L g1585 ( 
.A(n_1372),
.B(n_1437),
.Y(n_1585)
);

AND2x2_ASAP7_75t_L g1586 ( 
.A(n_1435),
.B(n_1440),
.Y(n_1586)
);

OAI31xp33_ASAP7_75t_L g1587 ( 
.A1(n_1440),
.A2(n_1399),
.A3(n_1406),
.B(n_1514),
.Y(n_1587)
);

INVx1_ASAP7_75t_SL g1588 ( 
.A(n_1392),
.Y(n_1588)
);

AND2x2_ASAP7_75t_L g1589 ( 
.A(n_1435),
.B(n_1442),
.Y(n_1589)
);

NAND2xp5_ASAP7_75t_L g1590 ( 
.A(n_1435),
.B(n_1495),
.Y(n_1590)
);

OA21x2_ASAP7_75t_L g1591 ( 
.A1(n_1462),
.A2(n_1468),
.B(n_1476),
.Y(n_1591)
);

AOI21xp5_ASAP7_75t_SL g1592 ( 
.A1(n_1436),
.A2(n_1386),
.B(n_1510),
.Y(n_1592)
);

AOI21x1_ASAP7_75t_SL g1593 ( 
.A1(n_1490),
.A2(n_1411),
.B(n_1487),
.Y(n_1593)
);

O2A1O1Ixp5_ASAP7_75t_L g1594 ( 
.A1(n_1380),
.A2(n_1410),
.B(n_1491),
.C(n_1388),
.Y(n_1594)
);

AOI21xp5_ASAP7_75t_L g1595 ( 
.A1(n_1377),
.A2(n_1463),
.B(n_1482),
.Y(n_1595)
);

OAI22xp5_ASAP7_75t_L g1596 ( 
.A1(n_1436),
.A2(n_1386),
.B1(n_1471),
.B2(n_1482),
.Y(n_1596)
);

HB1xp67_ASAP7_75t_L g1597 ( 
.A(n_1400),
.Y(n_1597)
);

INVx1_ASAP7_75t_L g1598 ( 
.A(n_1430),
.Y(n_1598)
);

OA21x2_ASAP7_75t_L g1599 ( 
.A1(n_1479),
.A2(n_1499),
.B(n_1504),
.Y(n_1599)
);

INVxp67_ASAP7_75t_L g1600 ( 
.A(n_1471),
.Y(n_1600)
);

OA21x2_ASAP7_75t_L g1601 ( 
.A1(n_1500),
.A2(n_1502),
.B(n_1378),
.Y(n_1601)
);

OA21x2_ASAP7_75t_L g1602 ( 
.A1(n_1382),
.A2(n_1434),
.B(n_1407),
.Y(n_1602)
);

AND2x2_ASAP7_75t_L g1603 ( 
.A(n_1507),
.B(n_1514),
.Y(n_1603)
);

NAND2xp5_ASAP7_75t_L g1604 ( 
.A(n_1507),
.B(n_1365),
.Y(n_1604)
);

AND2x2_ASAP7_75t_L g1605 ( 
.A(n_1375),
.B(n_1370),
.Y(n_1605)
);

CKINVDCx20_ASAP7_75t_R g1606 ( 
.A(n_1392),
.Y(n_1606)
);

O2A1O1Ixp5_ASAP7_75t_L g1607 ( 
.A1(n_1369),
.A2(n_1458),
.B(n_1518),
.C(n_1511),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_1374),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_1374),
.Y(n_1609)
);

OAI22xp5_ASAP7_75t_L g1610 ( 
.A1(n_1467),
.A2(n_1458),
.B1(n_1518),
.B2(n_1511),
.Y(n_1610)
);

CKINVDCx20_ASAP7_75t_R g1611 ( 
.A(n_1392),
.Y(n_1611)
);

NAND2xp5_ASAP7_75t_L g1612 ( 
.A(n_1365),
.B(n_1366),
.Y(n_1612)
);

OAI22xp5_ASAP7_75t_L g1613 ( 
.A1(n_1467),
.A2(n_1458),
.B1(n_1518),
.B2(n_1511),
.Y(n_1613)
);

AOI21xp5_ASAP7_75t_SL g1614 ( 
.A1(n_1367),
.A2(n_1452),
.B(n_1424),
.Y(n_1614)
);

AND2x2_ASAP7_75t_L g1615 ( 
.A(n_1375),
.B(n_1370),
.Y(n_1615)
);

NAND2xp5_ASAP7_75t_L g1616 ( 
.A(n_1365),
.B(n_1366),
.Y(n_1616)
);

AOI21x1_ASAP7_75t_SL g1617 ( 
.A1(n_1461),
.A2(n_1506),
.B(n_1492),
.Y(n_1617)
);

AOI221x1_ASAP7_75t_SL g1618 ( 
.A1(n_1515),
.A2(n_1518),
.B1(n_1511),
.B2(n_1458),
.C(n_1384),
.Y(n_1618)
);

AOI21xp5_ASAP7_75t_SL g1619 ( 
.A1(n_1367),
.A2(n_1452),
.B(n_1424),
.Y(n_1619)
);

O2A1O1Ixp5_ASAP7_75t_L g1620 ( 
.A1(n_1369),
.A2(n_1458),
.B(n_1518),
.C(n_1511),
.Y(n_1620)
);

AND2x4_ASAP7_75t_L g1621 ( 
.A(n_1469),
.B(n_1424),
.Y(n_1621)
);

OAI22xp5_ASAP7_75t_L g1622 ( 
.A1(n_1467),
.A2(n_1458),
.B1(n_1518),
.B2(n_1511),
.Y(n_1622)
);

BUFx8_ASAP7_75t_SL g1623 ( 
.A(n_1411),
.Y(n_1623)
);

OAI22xp5_ASAP7_75t_L g1624 ( 
.A1(n_1467),
.A2(n_1458),
.B1(n_1518),
.B2(n_1511),
.Y(n_1624)
);

AND2x2_ASAP7_75t_L g1625 ( 
.A(n_1375),
.B(n_1370),
.Y(n_1625)
);

O2A1O1Ixp33_ASAP7_75t_L g1626 ( 
.A1(n_1458),
.A2(n_747),
.B(n_1518),
.C(n_1511),
.Y(n_1626)
);

O2A1O1Ixp33_ASAP7_75t_L g1627 ( 
.A1(n_1458),
.A2(n_747),
.B(n_1518),
.C(n_1511),
.Y(n_1627)
);

AND2x2_ASAP7_75t_L g1628 ( 
.A(n_1375),
.B(n_1370),
.Y(n_1628)
);

OR2x2_ASAP7_75t_L g1629 ( 
.A(n_1464),
.B(n_1512),
.Y(n_1629)
);

INVx1_ASAP7_75t_L g1630 ( 
.A(n_1374),
.Y(n_1630)
);

BUFx3_ASAP7_75t_L g1631 ( 
.A(n_1403),
.Y(n_1631)
);

NAND2xp5_ASAP7_75t_L g1632 ( 
.A(n_1365),
.B(n_1366),
.Y(n_1632)
);

INVxp67_ASAP7_75t_L g1633 ( 
.A(n_1366),
.Y(n_1633)
);

INVx1_ASAP7_75t_SL g1634 ( 
.A(n_1392),
.Y(n_1634)
);

O2A1O1Ixp5_ASAP7_75t_L g1635 ( 
.A1(n_1369),
.A2(n_1458),
.B(n_1518),
.C(n_1511),
.Y(n_1635)
);

CKINVDCx5p33_ASAP7_75t_R g1636 ( 
.A(n_1392),
.Y(n_1636)
);

AOI21xp5_ASAP7_75t_SL g1637 ( 
.A1(n_1367),
.A2(n_1452),
.B(n_1424),
.Y(n_1637)
);

NAND2xp5_ASAP7_75t_L g1638 ( 
.A(n_1365),
.B(n_1366),
.Y(n_1638)
);

AND2x2_ASAP7_75t_L g1639 ( 
.A(n_1375),
.B(n_1370),
.Y(n_1639)
);

INVx1_ASAP7_75t_SL g1640 ( 
.A(n_1392),
.Y(n_1640)
);

OAI22xp5_ASAP7_75t_L g1641 ( 
.A1(n_1467),
.A2(n_1458),
.B1(n_1518),
.B2(n_1511),
.Y(n_1641)
);

O2A1O1Ixp33_ASAP7_75t_L g1642 ( 
.A1(n_1458),
.A2(n_747),
.B(n_1518),
.C(n_1511),
.Y(n_1642)
);

O2A1O1Ixp33_ASAP7_75t_L g1643 ( 
.A1(n_1458),
.A2(n_747),
.B(n_1518),
.C(n_1511),
.Y(n_1643)
);

AND2x2_ASAP7_75t_L g1644 ( 
.A(n_1375),
.B(n_1370),
.Y(n_1644)
);

NAND2xp5_ASAP7_75t_L g1645 ( 
.A(n_1365),
.B(n_1366),
.Y(n_1645)
);

BUFx2_ASAP7_75t_R g1646 ( 
.A(n_1564),
.Y(n_1646)
);

OA21x2_ASAP7_75t_L g1647 ( 
.A1(n_1595),
.A2(n_1576),
.B(n_1561),
.Y(n_1647)
);

OR2x2_ASAP7_75t_L g1648 ( 
.A(n_1529),
.B(n_1629),
.Y(n_1648)
);

OAI22xp5_ASAP7_75t_L g1649 ( 
.A1(n_1626),
.A2(n_1642),
.B1(n_1643),
.B2(n_1627),
.Y(n_1649)
);

OR2x6_ASAP7_75t_L g1650 ( 
.A(n_1579),
.B(n_1542),
.Y(n_1650)
);

AOI22xp33_ASAP7_75t_L g1651 ( 
.A1(n_1544),
.A2(n_1534),
.B1(n_1548),
.B2(n_1559),
.Y(n_1651)
);

INVx1_ASAP7_75t_L g1652 ( 
.A(n_1565),
.Y(n_1652)
);

AND2x2_ASAP7_75t_L g1653 ( 
.A(n_1603),
.B(n_1520),
.Y(n_1653)
);

INVx3_ASAP7_75t_L g1654 ( 
.A(n_1525),
.Y(n_1654)
);

AND2x2_ASAP7_75t_L g1655 ( 
.A(n_1605),
.B(n_1615),
.Y(n_1655)
);

CKINVDCx20_ASAP7_75t_R g1656 ( 
.A(n_1606),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1556),
.Y(n_1657)
);

AO21x2_ASAP7_75t_L g1658 ( 
.A1(n_1598),
.A2(n_1581),
.B(n_1543),
.Y(n_1658)
);

NAND2xp5_ASAP7_75t_L g1659 ( 
.A(n_1633),
.B(n_1645),
.Y(n_1659)
);

INVx1_ASAP7_75t_L g1660 ( 
.A(n_1608),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_1609),
.Y(n_1661)
);

OR2x6_ASAP7_75t_L g1662 ( 
.A(n_1579),
.B(n_1542),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_1630),
.Y(n_1663)
);

INVx1_ASAP7_75t_L g1664 ( 
.A(n_1560),
.Y(n_1664)
);

AO21x2_ASAP7_75t_L g1665 ( 
.A1(n_1581),
.A2(n_1543),
.B(n_1563),
.Y(n_1665)
);

AOI22xp33_ASAP7_75t_L g1666 ( 
.A1(n_1544),
.A2(n_1610),
.B1(n_1641),
.B2(n_1522),
.Y(n_1666)
);

INVx1_ASAP7_75t_L g1667 ( 
.A(n_1554),
.Y(n_1667)
);

INVx1_ASAP7_75t_L g1668 ( 
.A(n_1558),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_1574),
.Y(n_1669)
);

NAND2xp5_ASAP7_75t_L g1670 ( 
.A(n_1633),
.B(n_1612),
.Y(n_1670)
);

BUFx2_ASAP7_75t_L g1671 ( 
.A(n_1579),
.Y(n_1671)
);

INVx3_ASAP7_75t_L g1672 ( 
.A(n_1525),
.Y(n_1672)
);

AO21x2_ASAP7_75t_L g1673 ( 
.A1(n_1600),
.A2(n_1567),
.B(n_1597),
.Y(n_1673)
);

AOI22xp33_ASAP7_75t_L g1674 ( 
.A1(n_1613),
.A2(n_1622),
.B1(n_1624),
.B2(n_1566),
.Y(n_1674)
);

AND2x2_ASAP7_75t_L g1675 ( 
.A(n_1625),
.B(n_1628),
.Y(n_1675)
);

AND2x2_ASAP7_75t_L g1676 ( 
.A(n_1639),
.B(n_1644),
.Y(n_1676)
);

INVxp33_ASAP7_75t_L g1677 ( 
.A(n_1536),
.Y(n_1677)
);

INVx1_ASAP7_75t_L g1678 ( 
.A(n_1550),
.Y(n_1678)
);

INVx1_ASAP7_75t_L g1679 ( 
.A(n_1570),
.Y(n_1679)
);

INVx1_ASAP7_75t_L g1680 ( 
.A(n_1569),
.Y(n_1680)
);

AOI22xp33_ASAP7_75t_L g1681 ( 
.A1(n_1552),
.A2(n_1638),
.B1(n_1632),
.B2(n_1616),
.Y(n_1681)
);

AND2x2_ASAP7_75t_L g1682 ( 
.A(n_1582),
.B(n_1528),
.Y(n_1682)
);

BUFx2_ASAP7_75t_L g1683 ( 
.A(n_1578),
.Y(n_1683)
);

NAND2xp5_ASAP7_75t_L g1684 ( 
.A(n_1533),
.B(n_1524),
.Y(n_1684)
);

AO21x2_ASAP7_75t_L g1685 ( 
.A1(n_1567),
.A2(n_1573),
.B(n_1539),
.Y(n_1685)
);

NAND2xp5_ASAP7_75t_L g1686 ( 
.A(n_1532),
.B(n_1527),
.Y(n_1686)
);

OR2x2_ASAP7_75t_L g1687 ( 
.A(n_1545),
.B(n_1527),
.Y(n_1687)
);

OR2x2_ASAP7_75t_L g1688 ( 
.A(n_1535),
.B(n_1584),
.Y(n_1688)
);

BUFx2_ASAP7_75t_L g1689 ( 
.A(n_1535),
.Y(n_1689)
);

INVx1_ASAP7_75t_L g1690 ( 
.A(n_1573),
.Y(n_1690)
);

OAI22xp33_ASAP7_75t_L g1691 ( 
.A1(n_1604),
.A2(n_1585),
.B1(n_1580),
.B2(n_1523),
.Y(n_1691)
);

AND2x2_ASAP7_75t_L g1692 ( 
.A(n_1525),
.B(n_1607),
.Y(n_1692)
);

INVx1_ASAP7_75t_L g1693 ( 
.A(n_1538),
.Y(n_1693)
);

AND2x2_ASAP7_75t_L g1694 ( 
.A(n_1620),
.B(n_1635),
.Y(n_1694)
);

AND2x2_ASAP7_75t_L g1695 ( 
.A(n_1568),
.B(n_1596),
.Y(n_1695)
);

NAND2xp5_ASAP7_75t_L g1696 ( 
.A(n_1618),
.B(n_1549),
.Y(n_1696)
);

OAI21x1_ASAP7_75t_L g1697 ( 
.A1(n_1551),
.A2(n_1555),
.B(n_1602),
.Y(n_1697)
);

INVx1_ASAP7_75t_L g1698 ( 
.A(n_1590),
.Y(n_1698)
);

OAI21xp5_ASAP7_75t_L g1699 ( 
.A1(n_1541),
.A2(n_1530),
.B(n_1531),
.Y(n_1699)
);

AO21x2_ASAP7_75t_L g1700 ( 
.A1(n_1557),
.A2(n_1547),
.B(n_1546),
.Y(n_1700)
);

OAI21x1_ASAP7_75t_L g1701 ( 
.A1(n_1601),
.A2(n_1591),
.B(n_1583),
.Y(n_1701)
);

AND2x4_ASAP7_75t_L g1702 ( 
.A(n_1537),
.B(n_1519),
.Y(n_1702)
);

INVx1_ASAP7_75t_L g1703 ( 
.A(n_1572),
.Y(n_1703)
);

OR2x6_ASAP7_75t_L g1704 ( 
.A(n_1592),
.B(n_1553),
.Y(n_1704)
);

INVx1_ASAP7_75t_L g1705 ( 
.A(n_1594),
.Y(n_1705)
);

AND2x2_ASAP7_75t_L g1706 ( 
.A(n_1631),
.B(n_1575),
.Y(n_1706)
);

BUFx2_ASAP7_75t_L g1707 ( 
.A(n_1631),
.Y(n_1707)
);

CKINVDCx6p67_ASAP7_75t_R g1708 ( 
.A(n_1562),
.Y(n_1708)
);

AND2x2_ASAP7_75t_L g1709 ( 
.A(n_1586),
.B(n_1587),
.Y(n_1709)
);

INVx2_ASAP7_75t_L g1710 ( 
.A(n_1583),
.Y(n_1710)
);

AND2x2_ASAP7_75t_L g1711 ( 
.A(n_1583),
.B(n_1591),
.Y(n_1711)
);

OA21x2_ASAP7_75t_L g1712 ( 
.A1(n_1621),
.A2(n_1557),
.B(n_1537),
.Y(n_1712)
);

HB1xp67_ASAP7_75t_L g1713 ( 
.A(n_1562),
.Y(n_1713)
);

AND2x2_ASAP7_75t_L g1714 ( 
.A(n_1682),
.B(n_1599),
.Y(n_1714)
);

AND2x2_ASAP7_75t_L g1715 ( 
.A(n_1682),
.B(n_1599),
.Y(n_1715)
);

AND2x2_ASAP7_75t_L g1716 ( 
.A(n_1653),
.B(n_1599),
.Y(n_1716)
);

OR2x2_ASAP7_75t_L g1717 ( 
.A(n_1687),
.B(n_1688),
.Y(n_1717)
);

INVx2_ASAP7_75t_L g1718 ( 
.A(n_1710),
.Y(n_1718)
);

BUFx3_ASAP7_75t_L g1719 ( 
.A(n_1712),
.Y(n_1719)
);

AND2x2_ASAP7_75t_L g1720 ( 
.A(n_1653),
.B(n_1692),
.Y(n_1720)
);

AND2x2_ASAP7_75t_L g1721 ( 
.A(n_1692),
.B(n_1637),
.Y(n_1721)
);

AND2x4_ASAP7_75t_L g1722 ( 
.A(n_1650),
.B(n_1537),
.Y(n_1722)
);

INVxp67_ASAP7_75t_L g1723 ( 
.A(n_1686),
.Y(n_1723)
);

AND2x2_ASAP7_75t_L g1724 ( 
.A(n_1685),
.B(n_1619),
.Y(n_1724)
);

INVx1_ASAP7_75t_L g1725 ( 
.A(n_1690),
.Y(n_1725)
);

INVxp67_ASAP7_75t_SL g1726 ( 
.A(n_1686),
.Y(n_1726)
);

AND2x2_ASAP7_75t_L g1727 ( 
.A(n_1685),
.B(n_1614),
.Y(n_1727)
);

BUFx2_ASAP7_75t_SL g1728 ( 
.A(n_1712),
.Y(n_1728)
);

AND2x4_ASAP7_75t_L g1729 ( 
.A(n_1650),
.B(n_1540),
.Y(n_1729)
);

INVx1_ASAP7_75t_L g1730 ( 
.A(n_1652),
.Y(n_1730)
);

AND2x2_ASAP7_75t_L g1731 ( 
.A(n_1711),
.B(n_1521),
.Y(n_1731)
);

HB1xp67_ASAP7_75t_L g1732 ( 
.A(n_1689),
.Y(n_1732)
);

INVx1_ASAP7_75t_L g1733 ( 
.A(n_1652),
.Y(n_1733)
);

OR2x2_ASAP7_75t_L g1734 ( 
.A(n_1687),
.B(n_1688),
.Y(n_1734)
);

OAI21xp33_ASAP7_75t_L g1735 ( 
.A1(n_1666),
.A2(n_1636),
.B(n_1564),
.Y(n_1735)
);

BUFx3_ASAP7_75t_L g1736 ( 
.A(n_1712),
.Y(n_1736)
);

NOR2xp67_ASAP7_75t_L g1737 ( 
.A(n_1679),
.B(n_1571),
.Y(n_1737)
);

NAND3xp33_ASAP7_75t_SL g1738 ( 
.A(n_1699),
.B(n_1577),
.C(n_1606),
.Y(n_1738)
);

AND2x2_ASAP7_75t_L g1739 ( 
.A(n_1647),
.B(n_1654),
.Y(n_1739)
);

NAND2x1_ASAP7_75t_L g1740 ( 
.A(n_1650),
.B(n_1621),
.Y(n_1740)
);

BUFx3_ASAP7_75t_L g1741 ( 
.A(n_1712),
.Y(n_1741)
);

AOI22xp33_ASAP7_75t_L g1742 ( 
.A1(n_1651),
.A2(n_1523),
.B1(n_1640),
.B2(n_1588),
.Y(n_1742)
);

NAND4xp25_ASAP7_75t_L g1743 ( 
.A(n_1699),
.B(n_1634),
.C(n_1526),
.D(n_1617),
.Y(n_1743)
);

AND2x4_ASAP7_75t_L g1744 ( 
.A(n_1650),
.B(n_1589),
.Y(n_1744)
);

HB1xp67_ASAP7_75t_L g1745 ( 
.A(n_1673),
.Y(n_1745)
);

OR2x2_ASAP7_75t_L g1746 ( 
.A(n_1659),
.B(n_1636),
.Y(n_1746)
);

INVxp67_ASAP7_75t_L g1747 ( 
.A(n_1703),
.Y(n_1747)
);

AND2x2_ASAP7_75t_L g1748 ( 
.A(n_1654),
.B(n_1672),
.Y(n_1748)
);

OR2x2_ASAP7_75t_L g1749 ( 
.A(n_1659),
.B(n_1670),
.Y(n_1749)
);

INVx1_ASAP7_75t_L g1750 ( 
.A(n_1730),
.Y(n_1750)
);

OAI22xp33_ASAP7_75t_L g1751 ( 
.A1(n_1738),
.A2(n_1649),
.B1(n_1684),
.B2(n_1696),
.Y(n_1751)
);

NAND2xp5_ASAP7_75t_L g1752 ( 
.A(n_1726),
.B(n_1684),
.Y(n_1752)
);

HB1xp67_ASAP7_75t_L g1753 ( 
.A(n_1732),
.Y(n_1753)
);

INVx2_ASAP7_75t_L g1754 ( 
.A(n_1718),
.Y(n_1754)
);

AOI33xp33_ASAP7_75t_L g1755 ( 
.A1(n_1721),
.A2(n_1674),
.A3(n_1694),
.B1(n_1681),
.B2(n_1703),
.B3(n_1657),
.Y(n_1755)
);

AO21x2_ASAP7_75t_L g1756 ( 
.A1(n_1745),
.A2(n_1705),
.B(n_1665),
.Y(n_1756)
);

NAND2xp5_ASAP7_75t_L g1757 ( 
.A(n_1726),
.B(n_1694),
.Y(n_1757)
);

NOR2xp33_ASAP7_75t_R g1758 ( 
.A(n_1738),
.B(n_1611),
.Y(n_1758)
);

INVx4_ASAP7_75t_L g1759 ( 
.A(n_1719),
.Y(n_1759)
);

INVx1_ASAP7_75t_SL g1760 ( 
.A(n_1746),
.Y(n_1760)
);

INVx1_ASAP7_75t_L g1761 ( 
.A(n_1730),
.Y(n_1761)
);

OAI22xp5_ASAP7_75t_L g1762 ( 
.A1(n_1735),
.A2(n_1649),
.B1(n_1696),
.B2(n_1677),
.Y(n_1762)
);

NOR4xp25_ASAP7_75t_SL g1763 ( 
.A(n_1735),
.B(n_1707),
.C(n_1671),
.D(n_1683),
.Y(n_1763)
);

AOI221xp5_ASAP7_75t_L g1764 ( 
.A1(n_1723),
.A2(n_1665),
.B1(n_1670),
.B2(n_1679),
.C(n_1667),
.Y(n_1764)
);

NOR2xp33_ASAP7_75t_L g1765 ( 
.A(n_1743),
.B(n_1746),
.Y(n_1765)
);

INVx1_ASAP7_75t_L g1766 ( 
.A(n_1730),
.Y(n_1766)
);

AND2x4_ASAP7_75t_SL g1767 ( 
.A(n_1729),
.B(n_1708),
.Y(n_1767)
);

NAND2xp5_ASAP7_75t_L g1768 ( 
.A(n_1723),
.B(n_1664),
.Y(n_1768)
);

NAND2xp33_ASAP7_75t_SL g1769 ( 
.A(n_1740),
.B(n_1611),
.Y(n_1769)
);

AOI22xp5_ASAP7_75t_L g1770 ( 
.A1(n_1743),
.A2(n_1665),
.B1(n_1700),
.B2(n_1709),
.Y(n_1770)
);

AND2x4_ASAP7_75t_L g1771 ( 
.A(n_1729),
.B(n_1662),
.Y(n_1771)
);

OAI221xp5_ASAP7_75t_SL g1772 ( 
.A1(n_1719),
.A2(n_1691),
.B1(n_1695),
.B2(n_1655),
.C(n_1675),
.Y(n_1772)
);

BUFx2_ASAP7_75t_L g1773 ( 
.A(n_1744),
.Y(n_1773)
);

OAI211xp5_ASAP7_75t_L g1774 ( 
.A1(n_1747),
.A2(n_1707),
.B(n_1713),
.C(n_1672),
.Y(n_1774)
);

NAND3xp33_ASAP7_75t_L g1775 ( 
.A(n_1747),
.B(n_1664),
.C(n_1667),
.Y(n_1775)
);

INVx1_ASAP7_75t_L g1776 ( 
.A(n_1733),
.Y(n_1776)
);

BUFx2_ASAP7_75t_L g1777 ( 
.A(n_1744),
.Y(n_1777)
);

INVx3_ASAP7_75t_L g1778 ( 
.A(n_1719),
.Y(n_1778)
);

INVx1_ASAP7_75t_L g1779 ( 
.A(n_1733),
.Y(n_1779)
);

AOI22xp33_ASAP7_75t_L g1780 ( 
.A1(n_1742),
.A2(n_1700),
.B1(n_1658),
.B2(n_1704),
.Y(n_1780)
);

AND2x2_ASAP7_75t_L g1781 ( 
.A(n_1720),
.B(n_1683),
.Y(n_1781)
);

OAI221xp5_ASAP7_75t_L g1782 ( 
.A1(n_1736),
.A2(n_1680),
.B1(n_1668),
.B2(n_1698),
.C(n_1669),
.Y(n_1782)
);

NOR3xp33_ASAP7_75t_L g1783 ( 
.A(n_1736),
.B(n_1697),
.C(n_1672),
.Y(n_1783)
);

OR2x2_ASAP7_75t_L g1784 ( 
.A(n_1717),
.B(n_1648),
.Y(n_1784)
);

NAND3xp33_ASAP7_75t_L g1785 ( 
.A(n_1724),
.B(n_1668),
.C(n_1698),
.Y(n_1785)
);

INVxp67_ASAP7_75t_SL g1786 ( 
.A(n_1737),
.Y(n_1786)
);

INVx1_ASAP7_75t_SL g1787 ( 
.A(n_1746),
.Y(n_1787)
);

OAI221xp5_ASAP7_75t_L g1788 ( 
.A1(n_1736),
.A2(n_1669),
.B1(n_1678),
.B2(n_1693),
.C(n_1663),
.Y(n_1788)
);

AOI222xp33_ASAP7_75t_L g1789 ( 
.A1(n_1727),
.A2(n_1736),
.B1(n_1741),
.B2(n_1742),
.C1(n_1721),
.C2(n_1737),
.Y(n_1789)
);

CKINVDCx16_ASAP7_75t_R g1790 ( 
.A(n_1729),
.Y(n_1790)
);

AND2x2_ASAP7_75t_L g1791 ( 
.A(n_1720),
.B(n_1706),
.Y(n_1791)
);

AND2x2_ASAP7_75t_L g1792 ( 
.A(n_1720),
.B(n_1716),
.Y(n_1792)
);

OR2x2_ASAP7_75t_L g1793 ( 
.A(n_1717),
.B(n_1648),
.Y(n_1793)
);

AOI221xp5_ASAP7_75t_L g1794 ( 
.A1(n_1745),
.A2(n_1700),
.B1(n_1663),
.B2(n_1661),
.C(n_1660),
.Y(n_1794)
);

AOI31xp33_ASAP7_75t_L g1795 ( 
.A1(n_1721),
.A2(n_1706),
.A3(n_1676),
.B(n_1702),
.Y(n_1795)
);

OR2x6_ASAP7_75t_L g1796 ( 
.A(n_1728),
.B(n_1704),
.Y(n_1796)
);

AND2x2_ASAP7_75t_L g1797 ( 
.A(n_1716),
.B(n_1676),
.Y(n_1797)
);

INVx2_ASAP7_75t_SL g1798 ( 
.A(n_1778),
.Y(n_1798)
);

INVx1_ASAP7_75t_L g1799 ( 
.A(n_1750),
.Y(n_1799)
);

INVx1_ASAP7_75t_L g1800 ( 
.A(n_1761),
.Y(n_1800)
);

AND2x2_ASAP7_75t_L g1801 ( 
.A(n_1790),
.B(n_1716),
.Y(n_1801)
);

INVx2_ASAP7_75t_L g1802 ( 
.A(n_1754),
.Y(n_1802)
);

INVxp67_ASAP7_75t_SL g1803 ( 
.A(n_1786),
.Y(n_1803)
);

AOI21x1_ASAP7_75t_L g1804 ( 
.A1(n_1757),
.A2(n_1739),
.B(n_1748),
.Y(n_1804)
);

INVx1_ASAP7_75t_L g1805 ( 
.A(n_1766),
.Y(n_1805)
);

INVx1_ASAP7_75t_L g1806 ( 
.A(n_1776),
.Y(n_1806)
);

INVx1_ASAP7_75t_L g1807 ( 
.A(n_1779),
.Y(n_1807)
);

INVx2_ASAP7_75t_SL g1808 ( 
.A(n_1778),
.Y(n_1808)
);

INVx1_ASAP7_75t_L g1809 ( 
.A(n_1784),
.Y(n_1809)
);

INVx1_ASAP7_75t_L g1810 ( 
.A(n_1793),
.Y(n_1810)
);

OA21x2_ASAP7_75t_L g1811 ( 
.A1(n_1794),
.A2(n_1701),
.B(n_1739),
.Y(n_1811)
);

INVx1_ASAP7_75t_L g1812 ( 
.A(n_1768),
.Y(n_1812)
);

INVx1_ASAP7_75t_L g1813 ( 
.A(n_1753),
.Y(n_1813)
);

BUFx2_ASAP7_75t_L g1814 ( 
.A(n_1769),
.Y(n_1814)
);

NAND2xp5_ASAP7_75t_L g1815 ( 
.A(n_1752),
.B(n_1749),
.Y(n_1815)
);

INVx2_ASAP7_75t_SL g1816 ( 
.A(n_1778),
.Y(n_1816)
);

NAND2xp5_ASAP7_75t_SL g1817 ( 
.A(n_1795),
.B(n_1727),
.Y(n_1817)
);

INVx1_ASAP7_75t_L g1818 ( 
.A(n_1775),
.Y(n_1818)
);

INVx3_ASAP7_75t_L g1819 ( 
.A(n_1759),
.Y(n_1819)
);

NAND2xp5_ASAP7_75t_SL g1820 ( 
.A(n_1769),
.B(n_1727),
.Y(n_1820)
);

BUFx3_ASAP7_75t_L g1821 ( 
.A(n_1770),
.Y(n_1821)
);

OA21x2_ASAP7_75t_L g1822 ( 
.A1(n_1764),
.A2(n_1701),
.B(n_1739),
.Y(n_1822)
);

INVx2_ASAP7_75t_SL g1823 ( 
.A(n_1767),
.Y(n_1823)
);

INVx1_ASAP7_75t_L g1824 ( 
.A(n_1788),
.Y(n_1824)
);

HB1xp67_ASAP7_75t_L g1825 ( 
.A(n_1760),
.Y(n_1825)
);

BUFx2_ASAP7_75t_L g1826 ( 
.A(n_1759),
.Y(n_1826)
);

AND2x4_ASAP7_75t_L g1827 ( 
.A(n_1771),
.B(n_1722),
.Y(n_1827)
);

AND2x2_ASAP7_75t_L g1828 ( 
.A(n_1797),
.B(n_1763),
.Y(n_1828)
);

NAND2xp5_ASAP7_75t_L g1829 ( 
.A(n_1755),
.B(n_1725),
.Y(n_1829)
);

NAND2xp5_ASAP7_75t_L g1830 ( 
.A(n_1755),
.B(n_1725),
.Y(n_1830)
);

HB1xp67_ASAP7_75t_L g1831 ( 
.A(n_1787),
.Y(n_1831)
);

NAND2xp5_ASAP7_75t_SL g1832 ( 
.A(n_1789),
.B(n_1729),
.Y(n_1832)
);

NAND2xp5_ASAP7_75t_L g1833 ( 
.A(n_1765),
.B(n_1725),
.Y(n_1833)
);

BUFx2_ASAP7_75t_L g1834 ( 
.A(n_1759),
.Y(n_1834)
);

AND2x2_ASAP7_75t_L g1835 ( 
.A(n_1797),
.B(n_1731),
.Y(n_1835)
);

HB1xp67_ASAP7_75t_L g1836 ( 
.A(n_1782),
.Y(n_1836)
);

AND2x2_ASAP7_75t_L g1837 ( 
.A(n_1828),
.B(n_1792),
.Y(n_1837)
);

INVx2_ASAP7_75t_L g1838 ( 
.A(n_1811),
.Y(n_1838)
);

AND2x4_ASAP7_75t_L g1839 ( 
.A(n_1827),
.B(n_1771),
.Y(n_1839)
);

INVx1_ASAP7_75t_L g1840 ( 
.A(n_1799),
.Y(n_1840)
);

INVx1_ASAP7_75t_L g1841 ( 
.A(n_1799),
.Y(n_1841)
);

AND2x2_ASAP7_75t_L g1842 ( 
.A(n_1828),
.B(n_1792),
.Y(n_1842)
);

INVx2_ASAP7_75t_L g1843 ( 
.A(n_1811),
.Y(n_1843)
);

NAND4xp25_ASAP7_75t_L g1844 ( 
.A(n_1821),
.B(n_1765),
.C(n_1783),
.D(n_1762),
.Y(n_1844)
);

AND2x4_ASAP7_75t_L g1845 ( 
.A(n_1827),
.B(n_1796),
.Y(n_1845)
);

AND2x2_ASAP7_75t_L g1846 ( 
.A(n_1801),
.B(n_1773),
.Y(n_1846)
);

AND2x2_ASAP7_75t_L g1847 ( 
.A(n_1801),
.B(n_1777),
.Y(n_1847)
);

INVx1_ASAP7_75t_L g1848 ( 
.A(n_1800),
.Y(n_1848)
);

AND2x2_ASAP7_75t_L g1849 ( 
.A(n_1814),
.B(n_1781),
.Y(n_1849)
);

AND2x2_ASAP7_75t_L g1850 ( 
.A(n_1814),
.B(n_1714),
.Y(n_1850)
);

OR2x2_ASAP7_75t_L g1851 ( 
.A(n_1829),
.B(n_1717),
.Y(n_1851)
);

AND2x2_ASAP7_75t_L g1852 ( 
.A(n_1835),
.B(n_1817),
.Y(n_1852)
);

AND2x2_ASAP7_75t_L g1853 ( 
.A(n_1835),
.B(n_1803),
.Y(n_1853)
);

NOR2xp67_ASAP7_75t_L g1854 ( 
.A(n_1820),
.B(n_1774),
.Y(n_1854)
);

INVx2_ASAP7_75t_L g1855 ( 
.A(n_1811),
.Y(n_1855)
);

INVx1_ASAP7_75t_L g1856 ( 
.A(n_1800),
.Y(n_1856)
);

INVx1_ASAP7_75t_L g1857 ( 
.A(n_1805),
.Y(n_1857)
);

NAND2x1p5_ASAP7_75t_L g1858 ( 
.A(n_1819),
.B(n_1740),
.Y(n_1858)
);

AND2x2_ASAP7_75t_L g1859 ( 
.A(n_1804),
.B(n_1714),
.Y(n_1859)
);

INVx1_ASAP7_75t_L g1860 ( 
.A(n_1805),
.Y(n_1860)
);

INVx1_ASAP7_75t_L g1861 ( 
.A(n_1806),
.Y(n_1861)
);

BUFx3_ASAP7_75t_L g1862 ( 
.A(n_1826),
.Y(n_1862)
);

INVx1_ASAP7_75t_L g1863 ( 
.A(n_1806),
.Y(n_1863)
);

HB1xp67_ASAP7_75t_L g1864 ( 
.A(n_1825),
.Y(n_1864)
);

INVx1_ASAP7_75t_L g1865 ( 
.A(n_1807),
.Y(n_1865)
);

NAND2x1p5_ASAP7_75t_L g1866 ( 
.A(n_1819),
.B(n_1740),
.Y(n_1866)
);

INVx1_ASAP7_75t_L g1867 ( 
.A(n_1807),
.Y(n_1867)
);

AND2x2_ASAP7_75t_L g1868 ( 
.A(n_1823),
.B(n_1791),
.Y(n_1868)
);

INVx2_ASAP7_75t_L g1869 ( 
.A(n_1811),
.Y(n_1869)
);

HB1xp67_ASAP7_75t_L g1870 ( 
.A(n_1831),
.Y(n_1870)
);

OAI211xp5_ASAP7_75t_L g1871 ( 
.A1(n_1818),
.A2(n_1758),
.B(n_1780),
.C(n_1772),
.Y(n_1871)
);

AND2x2_ASAP7_75t_L g1872 ( 
.A(n_1804),
.B(n_1714),
.Y(n_1872)
);

INVx4_ASAP7_75t_L g1873 ( 
.A(n_1819),
.Y(n_1873)
);

INVx1_ASAP7_75t_L g1874 ( 
.A(n_1809),
.Y(n_1874)
);

NOR2xp67_ASAP7_75t_L g1875 ( 
.A(n_1819),
.B(n_1785),
.Y(n_1875)
);

NOR2xp33_ASAP7_75t_L g1876 ( 
.A(n_1818),
.B(n_1646),
.Y(n_1876)
);

OR2x2_ASAP7_75t_L g1877 ( 
.A(n_1829),
.B(n_1734),
.Y(n_1877)
);

INVx1_ASAP7_75t_L g1878 ( 
.A(n_1809),
.Y(n_1878)
);

AND2x2_ASAP7_75t_L g1879 ( 
.A(n_1811),
.B(n_1715),
.Y(n_1879)
);

AND2x2_ASAP7_75t_L g1880 ( 
.A(n_1826),
.B(n_1715),
.Y(n_1880)
);

INVx1_ASAP7_75t_SL g1881 ( 
.A(n_1834),
.Y(n_1881)
);

NAND3x1_ASAP7_75t_L g1882 ( 
.A(n_1830),
.B(n_1758),
.C(n_1751),
.Y(n_1882)
);

OR2x2_ASAP7_75t_L g1883 ( 
.A(n_1830),
.B(n_1734),
.Y(n_1883)
);

INVxp67_ASAP7_75t_L g1884 ( 
.A(n_1864),
.Y(n_1884)
);

AND2x2_ASAP7_75t_L g1885 ( 
.A(n_1854),
.B(n_1853),
.Y(n_1885)
);

OR2x2_ASAP7_75t_L g1886 ( 
.A(n_1851),
.B(n_1833),
.Y(n_1886)
);

AND2x4_ASAP7_75t_L g1887 ( 
.A(n_1839),
.B(n_1827),
.Y(n_1887)
);

INVx2_ASAP7_75t_L g1888 ( 
.A(n_1838),
.Y(n_1888)
);

HB1xp67_ASAP7_75t_L g1889 ( 
.A(n_1870),
.Y(n_1889)
);

OR2x2_ASAP7_75t_L g1890 ( 
.A(n_1851),
.B(n_1833),
.Y(n_1890)
);

AND2x2_ASAP7_75t_L g1891 ( 
.A(n_1853),
.B(n_1849),
.Y(n_1891)
);

INVx1_ASAP7_75t_L g1892 ( 
.A(n_1840),
.Y(n_1892)
);

NAND2x1p5_ASAP7_75t_L g1893 ( 
.A(n_1862),
.B(n_1823),
.Y(n_1893)
);

INVxp67_ASAP7_75t_SL g1894 ( 
.A(n_1882),
.Y(n_1894)
);

O2A1O1Ixp33_ASAP7_75t_L g1895 ( 
.A1(n_1844),
.A2(n_1836),
.B(n_1821),
.C(n_1824),
.Y(n_1895)
);

INVx1_ASAP7_75t_L g1896 ( 
.A(n_1840),
.Y(n_1896)
);

INVx1_ASAP7_75t_L g1897 ( 
.A(n_1841),
.Y(n_1897)
);

NAND2xp5_ASAP7_75t_L g1898 ( 
.A(n_1881),
.B(n_1824),
.Y(n_1898)
);

INVx1_ASAP7_75t_L g1899 ( 
.A(n_1841),
.Y(n_1899)
);

OR2x2_ASAP7_75t_L g1900 ( 
.A(n_1877),
.B(n_1810),
.Y(n_1900)
);

OR2x2_ASAP7_75t_L g1901 ( 
.A(n_1877),
.B(n_1883),
.Y(n_1901)
);

INVx2_ASAP7_75t_L g1902 ( 
.A(n_1838),
.Y(n_1902)
);

INVx1_ASAP7_75t_L g1903 ( 
.A(n_1848),
.Y(n_1903)
);

OR2x2_ASAP7_75t_L g1904 ( 
.A(n_1883),
.B(n_1810),
.Y(n_1904)
);

INVx1_ASAP7_75t_L g1905 ( 
.A(n_1848),
.Y(n_1905)
);

OR2x6_ASAP7_75t_L g1906 ( 
.A(n_1882),
.B(n_1728),
.Y(n_1906)
);

INVx1_ASAP7_75t_L g1907 ( 
.A(n_1856),
.Y(n_1907)
);

INVx1_ASAP7_75t_L g1908 ( 
.A(n_1856),
.Y(n_1908)
);

INVx1_ASAP7_75t_L g1909 ( 
.A(n_1857),
.Y(n_1909)
);

INVx1_ASAP7_75t_L g1910 ( 
.A(n_1857),
.Y(n_1910)
);

NAND2xp5_ASAP7_75t_L g1911 ( 
.A(n_1881),
.B(n_1853),
.Y(n_1911)
);

OR2x2_ASAP7_75t_L g1912 ( 
.A(n_1874),
.B(n_1815),
.Y(n_1912)
);

BUFx2_ASAP7_75t_SL g1913 ( 
.A(n_1854),
.Y(n_1913)
);

INVx1_ASAP7_75t_L g1914 ( 
.A(n_1860),
.Y(n_1914)
);

INVx1_ASAP7_75t_L g1915 ( 
.A(n_1860),
.Y(n_1915)
);

NAND2xp5_ASAP7_75t_L g1916 ( 
.A(n_1874),
.B(n_1812),
.Y(n_1916)
);

AND2x2_ASAP7_75t_L g1917 ( 
.A(n_1849),
.B(n_1823),
.Y(n_1917)
);

INVx1_ASAP7_75t_L g1918 ( 
.A(n_1861),
.Y(n_1918)
);

INVx2_ASAP7_75t_SL g1919 ( 
.A(n_1862),
.Y(n_1919)
);

NAND2xp5_ASAP7_75t_L g1920 ( 
.A(n_1878),
.B(n_1812),
.Y(n_1920)
);

NOR2x1_ASAP7_75t_L g1921 ( 
.A(n_1862),
.B(n_1656),
.Y(n_1921)
);

INVx2_ASAP7_75t_SL g1922 ( 
.A(n_1868),
.Y(n_1922)
);

OR2x2_ASAP7_75t_L g1923 ( 
.A(n_1889),
.B(n_1844),
.Y(n_1923)
);

NAND2xp5_ASAP7_75t_L g1924 ( 
.A(n_1891),
.B(n_1878),
.Y(n_1924)
);

INVx1_ASAP7_75t_L g1925 ( 
.A(n_1889),
.Y(n_1925)
);

OAI22xp33_ASAP7_75t_L g1926 ( 
.A1(n_1906),
.A2(n_1821),
.B1(n_1843),
.B2(n_1869),
.Y(n_1926)
);

INVx2_ASAP7_75t_L g1927 ( 
.A(n_1906),
.Y(n_1927)
);

AND2x2_ASAP7_75t_L g1928 ( 
.A(n_1913),
.B(n_1849),
.Y(n_1928)
);

INVx1_ASAP7_75t_L g1929 ( 
.A(n_1892),
.Y(n_1929)
);

INVx1_ASAP7_75t_L g1930 ( 
.A(n_1896),
.Y(n_1930)
);

OR2x2_ASAP7_75t_L g1931 ( 
.A(n_1884),
.B(n_1861),
.Y(n_1931)
);

HB1xp67_ASAP7_75t_L g1932 ( 
.A(n_1917),
.Y(n_1932)
);

NAND2xp5_ASAP7_75t_L g1933 ( 
.A(n_1884),
.B(n_1868),
.Y(n_1933)
);

INVxp67_ASAP7_75t_SL g1934 ( 
.A(n_1894),
.Y(n_1934)
);

INVx1_ASAP7_75t_L g1935 ( 
.A(n_1897),
.Y(n_1935)
);

INVx1_ASAP7_75t_SL g1936 ( 
.A(n_1885),
.Y(n_1936)
);

OR2x2_ASAP7_75t_L g1937 ( 
.A(n_1900),
.B(n_1904),
.Y(n_1937)
);

AOI22xp33_ASAP7_75t_L g1938 ( 
.A1(n_1906),
.A2(n_1843),
.B1(n_1855),
.B2(n_1838),
.Y(n_1938)
);

OR2x2_ASAP7_75t_L g1939 ( 
.A(n_1901),
.B(n_1863),
.Y(n_1939)
);

OR2x6_ASAP7_75t_L g1940 ( 
.A(n_1895),
.B(n_1882),
.Y(n_1940)
);

NOR2xp33_ASAP7_75t_L g1941 ( 
.A(n_1921),
.B(n_1876),
.Y(n_1941)
);

AND2x2_ASAP7_75t_L g1942 ( 
.A(n_1885),
.B(n_1852),
.Y(n_1942)
);

OAI22xp5_ASAP7_75t_L g1943 ( 
.A1(n_1894),
.A2(n_1871),
.B1(n_1875),
.B2(n_1879),
.Y(n_1943)
);

NAND2xp5_ASAP7_75t_L g1944 ( 
.A(n_1922),
.B(n_1852),
.Y(n_1944)
);

INVx1_ASAP7_75t_L g1945 ( 
.A(n_1899),
.Y(n_1945)
);

AND2x2_ASAP7_75t_L g1946 ( 
.A(n_1917),
.B(n_1852),
.Y(n_1946)
);

AOI22xp33_ASAP7_75t_L g1947 ( 
.A1(n_1888),
.A2(n_1855),
.B1(n_1869),
.B2(n_1843),
.Y(n_1947)
);

INVx4_ASAP7_75t_L g1948 ( 
.A(n_1919),
.Y(n_1948)
);

AND3x1_ASAP7_75t_L g1949 ( 
.A(n_1895),
.B(n_1842),
.C(n_1837),
.Y(n_1949)
);

INVx2_ASAP7_75t_L g1950 ( 
.A(n_1888),
.Y(n_1950)
);

INVx1_ASAP7_75t_SL g1951 ( 
.A(n_1911),
.Y(n_1951)
);

AND3x1_ASAP7_75t_L g1952 ( 
.A(n_1928),
.B(n_1941),
.C(n_1942),
.Y(n_1952)
);

OR2x2_ASAP7_75t_L g1953 ( 
.A(n_1923),
.B(n_1898),
.Y(n_1953)
);

INVx1_ASAP7_75t_L g1954 ( 
.A(n_1925),
.Y(n_1954)
);

INVx1_ASAP7_75t_L g1955 ( 
.A(n_1925),
.Y(n_1955)
);

AND2x2_ASAP7_75t_L g1956 ( 
.A(n_1928),
.B(n_1922),
.Y(n_1956)
);

INVx2_ASAP7_75t_L g1957 ( 
.A(n_1940),
.Y(n_1957)
);

OAI22xp33_ASAP7_75t_L g1958 ( 
.A1(n_1940),
.A2(n_1855),
.B1(n_1869),
.B2(n_1822),
.Y(n_1958)
);

INVx2_ASAP7_75t_SL g1959 ( 
.A(n_1942),
.Y(n_1959)
);

NAND4xp25_ASAP7_75t_L g1960 ( 
.A(n_1923),
.B(n_1873),
.C(n_1837),
.D(n_1842),
.Y(n_1960)
);

HB1xp67_ASAP7_75t_L g1961 ( 
.A(n_1932),
.Y(n_1961)
);

A2O1A1Ixp33_ASAP7_75t_L g1962 ( 
.A1(n_1943),
.A2(n_1871),
.B(n_1879),
.C(n_1875),
.Y(n_1962)
);

OAI211xp5_ASAP7_75t_SL g1963 ( 
.A1(n_1936),
.A2(n_1919),
.B(n_1908),
.C(n_1918),
.Y(n_1963)
);

AND2x2_ASAP7_75t_L g1964 ( 
.A(n_1946),
.B(n_1893),
.Y(n_1964)
);

INVx1_ASAP7_75t_L g1965 ( 
.A(n_1937),
.Y(n_1965)
);

INVx1_ASAP7_75t_L g1966 ( 
.A(n_1937),
.Y(n_1966)
);

AND2x2_ASAP7_75t_L g1967 ( 
.A(n_1946),
.B(n_1893),
.Y(n_1967)
);

AOI21xp33_ASAP7_75t_SL g1968 ( 
.A1(n_1940),
.A2(n_1866),
.B(n_1858),
.Y(n_1968)
);

AOI21xp5_ASAP7_75t_L g1969 ( 
.A1(n_1940),
.A2(n_1832),
.B(n_1916),
.Y(n_1969)
);

INVx2_ASAP7_75t_L g1970 ( 
.A(n_1949),
.Y(n_1970)
);

OAI21xp5_ASAP7_75t_L g1971 ( 
.A1(n_1926),
.A2(n_1934),
.B(n_1938),
.Y(n_1971)
);

OAI32xp33_ASAP7_75t_L g1972 ( 
.A1(n_1951),
.A2(n_1879),
.A3(n_1886),
.B1(n_1890),
.B2(n_1914),
.Y(n_1972)
);

AOI22xp5_ASAP7_75t_L g1973 ( 
.A1(n_1950),
.A2(n_1822),
.B1(n_1902),
.B2(n_1837),
.Y(n_1973)
);

NOR2xp33_ASAP7_75t_L g1974 ( 
.A(n_1948),
.B(n_1933),
.Y(n_1974)
);

NOR3xp33_ASAP7_75t_SL g1975 ( 
.A(n_1960),
.B(n_1962),
.C(n_1974),
.Y(n_1975)
);

INVx2_ASAP7_75t_L g1976 ( 
.A(n_1964),
.Y(n_1976)
);

INVx1_ASAP7_75t_L g1977 ( 
.A(n_1961),
.Y(n_1977)
);

NAND2xp5_ASAP7_75t_L g1978 ( 
.A(n_1959),
.B(n_1948),
.Y(n_1978)
);

NAND2xp5_ASAP7_75t_L g1979 ( 
.A(n_1959),
.B(n_1948),
.Y(n_1979)
);

NAND2x1p5_ASAP7_75t_L g1980 ( 
.A(n_1957),
.B(n_1623),
.Y(n_1980)
);

OR2x2_ASAP7_75t_L g1981 ( 
.A(n_1953),
.B(n_1944),
.Y(n_1981)
);

INVx1_ASAP7_75t_L g1982 ( 
.A(n_1965),
.Y(n_1982)
);

INVx1_ASAP7_75t_L g1983 ( 
.A(n_1966),
.Y(n_1983)
);

NAND2xp5_ASAP7_75t_L g1984 ( 
.A(n_1956),
.B(n_1939),
.Y(n_1984)
);

INVxp67_ASAP7_75t_L g1985 ( 
.A(n_1952),
.Y(n_1985)
);

INVx1_ASAP7_75t_SL g1986 ( 
.A(n_1953),
.Y(n_1986)
);

NOR2xp33_ASAP7_75t_L g1987 ( 
.A(n_1964),
.B(n_1646),
.Y(n_1987)
);

NAND2xp5_ASAP7_75t_L g1988 ( 
.A(n_1956),
.B(n_1939),
.Y(n_1988)
);

INVx1_ASAP7_75t_L g1989 ( 
.A(n_1954),
.Y(n_1989)
);

NAND2xp5_ASAP7_75t_L g1990 ( 
.A(n_1967),
.B(n_1924),
.Y(n_1990)
);

AND4x2_ASAP7_75t_L g1991 ( 
.A(n_1975),
.B(n_1969),
.C(n_1970),
.D(n_1963),
.Y(n_1991)
);

OAI22xp5_ASAP7_75t_L g1992 ( 
.A1(n_1985),
.A2(n_1962),
.B1(n_1970),
.B2(n_1973),
.Y(n_1992)
);

NOR2x1_ASAP7_75t_L g1993 ( 
.A(n_1986),
.B(n_1955),
.Y(n_1993)
);

O2A1O1Ixp33_ASAP7_75t_L g1994 ( 
.A1(n_1986),
.A2(n_1972),
.B(n_1971),
.C(n_1957),
.Y(n_1994)
);

OAI211xp5_ASAP7_75t_SL g1995 ( 
.A1(n_1981),
.A2(n_1958),
.B(n_1927),
.C(n_1931),
.Y(n_1995)
);

AOI221xp5_ASAP7_75t_L g1996 ( 
.A1(n_1982),
.A2(n_1972),
.B1(n_1947),
.B2(n_1968),
.C(n_1950),
.Y(n_1996)
);

OAI21xp33_ASAP7_75t_L g1997 ( 
.A1(n_1976),
.A2(n_1967),
.B(n_1927),
.Y(n_1997)
);

AOI211xp5_ASAP7_75t_L g1998 ( 
.A1(n_1987),
.A2(n_1931),
.B(n_1929),
.C(n_1945),
.Y(n_1998)
);

AOI22xp5_ASAP7_75t_L g1999 ( 
.A1(n_1980),
.A2(n_1902),
.B1(n_1822),
.B2(n_1842),
.Y(n_1999)
);

AOI211xp5_ASAP7_75t_L g2000 ( 
.A1(n_1984),
.A2(n_1988),
.B(n_1983),
.C(n_1990),
.Y(n_2000)
);

AOI221xp5_ASAP7_75t_L g2001 ( 
.A1(n_1989),
.A2(n_1945),
.B1(n_1930),
.B2(n_1929),
.C(n_1935),
.Y(n_2001)
);

AOI21xp5_ASAP7_75t_L g2002 ( 
.A1(n_1978),
.A2(n_1930),
.B(n_1920),
.Y(n_2002)
);

NAND2xp33_ASAP7_75t_SL g2003 ( 
.A(n_1979),
.B(n_1873),
.Y(n_2003)
);

AOI221xp5_ASAP7_75t_L g2004 ( 
.A1(n_1977),
.A2(n_1915),
.B1(n_1907),
.B2(n_1905),
.C(n_1910),
.Y(n_2004)
);

AOI221xp5_ASAP7_75t_L g2005 ( 
.A1(n_1980),
.A2(n_1909),
.B1(n_1903),
.B2(n_1859),
.C(n_1872),
.Y(n_2005)
);

INVx1_ASAP7_75t_L g2006 ( 
.A(n_1993),
.Y(n_2006)
);

AOI221xp5_ASAP7_75t_L g2007 ( 
.A1(n_1995),
.A2(n_1859),
.B1(n_1872),
.B2(n_1912),
.C(n_1850),
.Y(n_2007)
);

OA22x2_ASAP7_75t_L g2008 ( 
.A1(n_1997),
.A2(n_1992),
.B1(n_1999),
.B2(n_1991),
.Y(n_2008)
);

AOI321xp33_ASAP7_75t_L g2009 ( 
.A1(n_1994),
.A2(n_1780),
.A3(n_1872),
.B1(n_1859),
.B2(n_1887),
.C(n_1850),
.Y(n_2009)
);

AOI22xp5_ASAP7_75t_L g2010 ( 
.A1(n_1996),
.A2(n_1822),
.B1(n_1887),
.B2(n_1850),
.Y(n_2010)
);

NOR4xp25_ASAP7_75t_L g2011 ( 
.A(n_2001),
.B(n_2004),
.C(n_2005),
.D(n_2000),
.Y(n_2011)
);

AOI21xp33_ASAP7_75t_SL g2012 ( 
.A1(n_1998),
.A2(n_1866),
.B(n_1858),
.Y(n_2012)
);

OAI221xp5_ASAP7_75t_L g2013 ( 
.A1(n_2002),
.A2(n_1822),
.B1(n_1728),
.B2(n_1866),
.C(n_1858),
.Y(n_2013)
);

INVx2_ASAP7_75t_SL g2014 ( 
.A(n_2006),
.Y(n_2014)
);

AOI21xp33_ASAP7_75t_L g2015 ( 
.A1(n_2008),
.A2(n_2003),
.B(n_1865),
.Y(n_2015)
);

INVx1_ASAP7_75t_L g2016 ( 
.A(n_2009),
.Y(n_2016)
);

INVx1_ASAP7_75t_L g2017 ( 
.A(n_2010),
.Y(n_2017)
);

NAND2xp5_ASAP7_75t_L g2018 ( 
.A(n_2011),
.B(n_1887),
.Y(n_2018)
);

INVx2_ASAP7_75t_L g2019 ( 
.A(n_2013),
.Y(n_2019)
);

NAND2xp5_ASAP7_75t_L g2020 ( 
.A(n_2007),
.B(n_1880),
.Y(n_2020)
);

INVx1_ASAP7_75t_L g2021 ( 
.A(n_2012),
.Y(n_2021)
);

AOI21xp33_ASAP7_75t_SL g2022 ( 
.A1(n_2018),
.A2(n_1623),
.B(n_1858),
.Y(n_2022)
);

CKINVDCx5p33_ASAP7_75t_R g2023 ( 
.A(n_2014),
.Y(n_2023)
);

INVxp67_ASAP7_75t_SL g2024 ( 
.A(n_2016),
.Y(n_2024)
);

HB1xp67_ASAP7_75t_L g2025 ( 
.A(n_2021),
.Y(n_2025)
);

OR2x2_ASAP7_75t_L g2026 ( 
.A(n_2020),
.B(n_1873),
.Y(n_2026)
);

HB1xp67_ASAP7_75t_L g2027 ( 
.A(n_2017),
.Y(n_2027)
);

XOR2xp5_ASAP7_75t_L g2028 ( 
.A(n_2027),
.B(n_2019),
.Y(n_2028)
);

AOI221xp5_ASAP7_75t_L g2029 ( 
.A1(n_2024),
.A2(n_2015),
.B1(n_1865),
.B2(n_1863),
.C(n_1867),
.Y(n_2029)
);

AOI21xp5_ASAP7_75t_L g2030 ( 
.A1(n_2023),
.A2(n_2015),
.B(n_1873),
.Y(n_2030)
);

AOI22xp5_ASAP7_75t_L g2031 ( 
.A1(n_2025),
.A2(n_1845),
.B1(n_1880),
.B2(n_1839),
.Y(n_2031)
);

NOR2xp33_ASAP7_75t_L g2032 ( 
.A(n_2028),
.B(n_2022),
.Y(n_2032)
);

OAI322xp33_ASAP7_75t_L g2033 ( 
.A1(n_2032),
.A2(n_2030),
.A3(n_2026),
.B1(n_2031),
.B2(n_2029),
.C1(n_1867),
.C2(n_1866),
.Y(n_2033)
);

AOI22xp33_ASAP7_75t_L g2034 ( 
.A1(n_2033),
.A2(n_1756),
.B1(n_1845),
.B2(n_1834),
.Y(n_2034)
);

OA22x2_ASAP7_75t_L g2035 ( 
.A1(n_2033),
.A2(n_1798),
.B1(n_1808),
.B2(n_1816),
.Y(n_2035)
);

OAI22x1_ASAP7_75t_L g2036 ( 
.A1(n_2035),
.A2(n_1845),
.B1(n_1798),
.B2(n_1808),
.Y(n_2036)
);

AOI22xp33_ASAP7_75t_L g2037 ( 
.A1(n_2034),
.A2(n_1845),
.B1(n_1756),
.B2(n_1880),
.Y(n_2037)
);

INVx1_ASAP7_75t_SL g2038 ( 
.A(n_2036),
.Y(n_2038)
);

INVx2_ASAP7_75t_L g2039 ( 
.A(n_2037),
.Y(n_2039)
);

NAND2xp5_ASAP7_75t_L g2040 ( 
.A(n_2038),
.B(n_1802),
.Y(n_2040)
);

INVx1_ASAP7_75t_L g2041 ( 
.A(n_2040),
.Y(n_2041)
);

AO21x2_ASAP7_75t_L g2042 ( 
.A1(n_2041),
.A2(n_2039),
.B(n_1593),
.Y(n_2042)
);

AOI22x1_ASAP7_75t_L g2043 ( 
.A1(n_2042),
.A2(n_1808),
.B1(n_1798),
.B2(n_1816),
.Y(n_2043)
);

AOI22xp5_ASAP7_75t_L g2044 ( 
.A1(n_2043),
.A2(n_1847),
.B1(n_1846),
.B2(n_1839),
.Y(n_2044)
);

AOI211xp5_ASAP7_75t_L g2045 ( 
.A1(n_2044),
.A2(n_1847),
.B(n_1846),
.C(n_1813),
.Y(n_2045)
);


endmodule