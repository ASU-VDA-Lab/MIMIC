module real_jpeg_8595_n_6 (n_5, n_4, n_0, n_1, n_2, n_3, n_6);

input n_5;
input n_4;
input n_0;
input n_1;
input n_2;
input n_3;

output n_6;

wire n_17;
wire n_8;
wire n_43;
wire n_37;
wire n_21;
wire n_33;
wire n_35;
wire n_38;
wire n_50;
wire n_29;
wire n_49;
wire n_10;
wire n_31;
wire n_9;
wire n_12;
wire n_24;
wire n_34;
wire n_44;
wire n_28;
wire n_46;
wire n_23;
wire n_11;
wire n_14;
wire n_51;
wire n_47;
wire n_45;
wire n_25;
wire n_42;
wire n_7;
wire n_22;
wire n_18;
wire n_40;
wire n_39;
wire n_36;
wire n_41;
wire n_26;
wire n_27;
wire n_20;
wire n_19;
wire n_48;
wire n_32;
wire n_30;
wire n_16;
wire n_15;
wire n_13;

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_0),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_1),
.Y(n_16)
);

OR2x2_ASAP7_75t_SL g37 ( 
.A(n_1),
.B(n_17),
.Y(n_37)
);

OR2x2_ASAP7_75t_SL g42 ( 
.A(n_1),
.B(n_3),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g10 ( 
.A(n_2),
.B(n_11),
.Y(n_10)
);

NAND2xp5_ASAP7_75t_L g12 ( 
.A(n_2),
.B(n_11),
.Y(n_12)
);

AOI22xp5_ASAP7_75t_SL g28 ( 
.A1(n_2),
.A2(n_29),
.B1(n_30),
.B2(n_31),
.Y(n_28)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_3),
.Y(n_17)
);

OR2x2_ASAP7_75t_L g27 ( 
.A(n_3),
.B(n_16),
.Y(n_27)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_4),
.Y(n_11)
);

AND2x2_ASAP7_75t_L g24 ( 
.A(n_4),
.B(n_25),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_SL g30 ( 
.A1(n_4),
.A2(n_5),
.B1(n_9),
.B2(n_11),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_4),
.B(n_44),
.Y(n_43)
);

INVx1_ASAP7_75t_L g9 ( 
.A(n_5),
.Y(n_9)
);

AOI21xp5_ASAP7_75t_SL g20 ( 
.A1(n_5),
.A2(n_10),
.B(n_12),
.Y(n_20)
);

OAI211xp5_ASAP7_75t_L g6 ( 
.A1(n_7),
.A2(n_13),
.B(n_22),
.C(n_45),
.Y(n_6)
);

CKINVDCx20_ASAP7_75t_R g7 ( 
.A(n_8),
.Y(n_7)
);

OAI21xp33_ASAP7_75t_L g39 ( 
.A1(n_8),
.A2(n_40),
.B(n_43),
.Y(n_39)
);

OA21x2_ASAP7_75t_L g8 ( 
.A1(n_9),
.A2(n_10),
.B(n_12),
.Y(n_8)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_18),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_15),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_15),
.B(n_25),
.Y(n_48)
);

OR2x2_ASAP7_75t_SL g15 ( 
.A(n_16),
.B(n_17),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_19),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_21),
.Y(n_19)
);

AOI21xp5_ASAP7_75t_L g50 ( 
.A1(n_20),
.A2(n_25),
.B(n_51),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_20),
.B(n_25),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_21),
.Y(n_25)
);

AOI211xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_26),
.B(n_34),
.C(n_39),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_24),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_25),
.B(n_33),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_25),
.B(n_36),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_25),
.B(n_41),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_SL g44 ( 
.A(n_25),
.B(n_37),
.Y(n_44)
);

OAI21xp5_ASAP7_75t_SL g47 ( 
.A1(n_25),
.A2(n_41),
.B(n_48),
.Y(n_47)
);

OAI21xp5_ASAP7_75t_L g26 ( 
.A1(n_27),
.A2(n_28),
.B(n_32),
.Y(n_26)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_27),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_28),
.Y(n_38)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_35),
.B(n_38),
.Y(n_34)
);

INVx1_ASAP7_75t_SL g36 ( 
.A(n_37),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_42),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_46),
.B(n_49),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_47),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_50),
.Y(n_49)
);


endmodule