module fake_jpeg_14000_n_432 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_432);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_432;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_430;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_15),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_7),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_7),
.Y(n_22)
);

BUFx16f_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_2),
.B(n_11),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_12),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

INVx5_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_3),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_3),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_9),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_7),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_8),
.Y(n_36)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_10),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_15),
.Y(n_38)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_13),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_0),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_15),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_6),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_0),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_10),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_19),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_45),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_19),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_46),
.Y(n_102)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_23),
.Y(n_47)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_47),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_25),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_48),
.B(n_49),
.Y(n_95)
);

CKINVDCx16_ASAP7_75t_R g49 ( 
.A(n_23),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_33),
.Y(n_50)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_50),
.Y(n_97)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_19),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_51),
.Y(n_125)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_44),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_52),
.Y(n_127)
);

BUFx10_ASAP7_75t_L g53 ( 
.A(n_30),
.Y(n_53)
);

INVx3_ASAP7_75t_SL g110 ( 
.A(n_53),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_21),
.Y(n_54)
);

INVx6_ASAP7_75t_L g131 ( 
.A(n_54),
.Y(n_131)
);

INVx6_ASAP7_75t_SL g55 ( 
.A(n_23),
.Y(n_55)
);

INVx5_ASAP7_75t_L g91 ( 
.A(n_55),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_21),
.Y(n_56)
);

INVx8_ASAP7_75t_L g111 ( 
.A(n_56),
.Y(n_111)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_57),
.Y(n_118)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_58),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_21),
.Y(n_59)
);

INVx8_ASAP7_75t_L g112 ( 
.A(n_59),
.Y(n_112)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_33),
.Y(n_60)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_60),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_24),
.Y(n_61)
);

INVx5_ASAP7_75t_L g123 ( 
.A(n_61),
.Y(n_123)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_20),
.Y(n_62)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_62),
.Y(n_107)
);

INVx1_ASAP7_75t_SL g63 ( 
.A(n_40),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g119 ( 
.A(n_63),
.B(n_72),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_24),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g124 ( 
.A(n_64),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_28),
.B(n_20),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_65),
.B(n_82),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_28),
.B(n_18),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_66),
.B(n_42),
.Y(n_90)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_27),
.Y(n_67)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_67),
.Y(n_122)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_38),
.Y(n_68)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_68),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_24),
.Y(n_69)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_69),
.Y(n_100)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_29),
.Y(n_70)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_70),
.Y(n_104)
);

INVx5_ASAP7_75t_L g71 ( 
.A(n_38),
.Y(n_71)
);

INVx4_ASAP7_75t_L g117 ( 
.A(n_71),
.Y(n_117)
);

INVx1_ASAP7_75t_SL g72 ( 
.A(n_40),
.Y(n_72)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_26),
.Y(n_73)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_73),
.Y(n_103)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_27),
.Y(n_74)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_74),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_26),
.Y(n_75)
);

INVx4_ASAP7_75t_L g130 ( 
.A(n_75),
.Y(n_130)
);

CKINVDCx16_ASAP7_75t_R g76 ( 
.A(n_29),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_76),
.B(n_79),
.Y(n_98)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_40),
.Y(n_77)
);

HB1xp67_ASAP7_75t_L g138 ( 
.A(n_77),
.Y(n_138)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_40),
.Y(n_78)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_78),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_37),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_37),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_80),
.B(n_83),
.Y(n_116)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_26),
.Y(n_81)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_81),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_18),
.B(n_14),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_22),
.B(n_12),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_36),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_84),
.B(n_85),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_22),
.B(n_12),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_36),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_86),
.B(n_89),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_44),
.Y(n_87)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_87),
.Y(n_108)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_44),
.Y(n_88)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_88),
.Y(n_115)
);

BUFx16f_ASAP7_75t_L g89 ( 
.A(n_30),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g179 ( 
.A(n_90),
.B(n_94),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_51),
.A2(n_16),
.B1(n_41),
.B2(n_17),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_92),
.A2(n_114),
.B1(n_120),
.B2(n_126),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_55),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_50),
.B(n_42),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_101),
.B(n_109),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_60),
.B(n_32),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_L g114 ( 
.A1(n_81),
.A2(n_35),
.B1(n_41),
.B2(n_16),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_L g120 ( 
.A1(n_88),
.A2(n_35),
.B1(n_41),
.B2(n_16),
.Y(n_120)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_77),
.Y(n_121)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_121),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_L g126 ( 
.A1(n_52),
.A2(n_17),
.B1(n_32),
.B2(n_31),
.Y(n_126)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_78),
.Y(n_129)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_129),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_47),
.B(n_31),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_134),
.B(n_139),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_73),
.A2(n_17),
.B1(n_43),
.B2(n_34),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_136),
.A2(n_70),
.B1(n_34),
.B2(n_43),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_63),
.B(n_0),
.Y(n_139)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_57),
.Y(n_140)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_140),
.Y(n_162)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_58),
.Y(n_141)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_141),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_137),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_142),
.B(n_145),
.Y(n_193)
);

AO22x1_ASAP7_75t_SL g143 ( 
.A1(n_97),
.A2(n_72),
.B1(n_53),
.B2(n_75),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_143),
.B(n_188),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_SL g144 ( 
.A(n_122),
.B(n_53),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_144),
.B(n_149),
.C(n_170),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_133),
.B(n_89),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_106),
.Y(n_146)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_146),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_138),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_147),
.B(n_151),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_135),
.B(n_68),
.C(n_87),
.Y(n_149)
);

AND2x2_ASAP7_75t_L g150 ( 
.A(n_119),
.B(n_71),
.Y(n_150)
);

INVx1_ASAP7_75t_SL g233 ( 
.A(n_150),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_138),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_96),
.Y(n_152)
);

BUFx3_ASAP7_75t_L g208 ( 
.A(n_152),
.Y(n_208)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_115),
.Y(n_153)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_153),
.Y(n_214)
);

OR2x2_ASAP7_75t_SL g154 ( 
.A(n_128),
.B(n_89),
.Y(n_154)
);

AND2x2_ASAP7_75t_L g205 ( 
.A(n_154),
.B(n_191),
.Y(n_205)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_119),
.Y(n_156)
);

HB1xp67_ASAP7_75t_L g221 ( 
.A(n_156),
.Y(n_221)
);

INVx11_ASAP7_75t_L g157 ( 
.A(n_104),
.Y(n_157)
);

INVx11_ASAP7_75t_L g222 ( 
.A(n_157),
.Y(n_222)
);

CKINVDCx14_ASAP7_75t_R g158 ( 
.A(n_98),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_158),
.B(n_168),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_114),
.A2(n_56),
.B1(n_69),
.B2(n_64),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_L g234 ( 
.A1(n_160),
.A2(n_167),
.B1(n_11),
.B2(n_164),
.Y(n_234)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_96),
.Y(n_161)
);

BUFx3_ASAP7_75t_L g209 ( 
.A(n_161),
.Y(n_209)
);

INVx5_ASAP7_75t_L g163 ( 
.A(n_117),
.Y(n_163)
);

INVx3_ASAP7_75t_L g194 ( 
.A(n_163),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_102),
.Y(n_164)
);

INVx3_ASAP7_75t_L g218 ( 
.A(n_164),
.Y(n_218)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_99),
.Y(n_165)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_165),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_166),
.A2(n_175),
.B1(n_184),
.B2(n_123),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_120),
.A2(n_61),
.B1(n_59),
.B2(n_54),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_116),
.B(n_39),
.Y(n_168)
);

AND2x2_ASAP7_75t_L g170 ( 
.A(n_107),
.B(n_39),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g171 ( 
.A(n_95),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_171),
.B(n_185),
.Y(n_217)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_103),
.Y(n_173)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_173),
.Y(n_237)
);

AOI22xp33_ASAP7_75t_SL g174 ( 
.A1(n_110),
.A2(n_46),
.B1(n_45),
.B2(n_3),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_SL g211 ( 
.A1(n_174),
.A2(n_176),
.B1(n_112),
.B2(n_111),
.Y(n_211)
);

AOI22xp33_ASAP7_75t_L g175 ( 
.A1(n_126),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_SL g176 ( 
.A1(n_110),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_176)
);

HB1xp67_ASAP7_75t_L g177 ( 
.A(n_105),
.Y(n_177)
);

CKINVDCx16_ASAP7_75t_R g196 ( 
.A(n_177),
.Y(n_196)
);

INVx3_ASAP7_75t_L g178 ( 
.A(n_117),
.Y(n_178)
);

INVx3_ASAP7_75t_L g235 ( 
.A(n_178),
.Y(n_235)
);

INVx6_ASAP7_75t_SL g181 ( 
.A(n_91),
.Y(n_181)
);

CKINVDCx16_ASAP7_75t_R g210 ( 
.A(n_181),
.Y(n_210)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_93),
.Y(n_182)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_182),
.Y(n_230)
);

INVx4_ASAP7_75t_L g183 ( 
.A(n_93),
.Y(n_183)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_183),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_108),
.A2(n_1),
.B1(n_5),
.B2(n_6),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_113),
.B(n_5),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_100),
.Y(n_186)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_186),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_91),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_187),
.B(n_189),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_111),
.B(n_112),
.Y(n_188)
);

CKINVDCx16_ASAP7_75t_R g189 ( 
.A(n_118),
.Y(n_189)
);

INVx3_ASAP7_75t_L g190 ( 
.A(n_104),
.Y(n_190)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_190),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_132),
.B(n_5),
.Y(n_191)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_100),
.Y(n_192)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_192),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_181),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_197),
.B(n_212),
.Y(n_238)
);

A2O1A1Ixp33_ASAP7_75t_L g199 ( 
.A1(n_172),
.A2(n_5),
.B(n_6),
.C(n_8),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_199),
.B(n_216),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_201),
.A2(n_225),
.B1(n_232),
.B2(n_167),
.Y(n_246)
);

AND2x2_ASAP7_75t_SL g202 ( 
.A(n_144),
.B(n_130),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_202),
.B(n_207),
.C(n_229),
.Y(n_250)
);

FAx1_ASAP7_75t_SL g203 ( 
.A(n_172),
.B(n_6),
.CI(n_8),
.CON(n_203),
.SN(n_203)
);

NOR2xp33_ASAP7_75t_SL g249 ( 
.A(n_203),
.B(n_184),
.Y(n_249)
);

AND2x2_ASAP7_75t_SL g207 ( 
.A(n_149),
.B(n_130),
.Y(n_207)
);

AOI22xp33_ASAP7_75t_SL g269 ( 
.A1(n_211),
.A2(n_221),
.B1(n_218),
.B2(n_209),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_157),
.Y(n_212)
);

AOI21xp5_ASAP7_75t_L g215 ( 
.A1(n_156),
.A2(n_123),
.B(n_124),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_SL g265 ( 
.A1(n_215),
.A2(n_143),
.B(n_159),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_155),
.B(n_131),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_L g219 ( 
.A1(n_170),
.A2(n_124),
.B(n_127),
.Y(n_219)
);

INVxp67_ASAP7_75t_L g262 ( 
.A(n_219),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_188),
.B(n_131),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_220),
.B(n_228),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_166),
.A2(n_125),
.B1(n_127),
.B2(n_102),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_165),
.B(n_125),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_150),
.B(n_8),
.C(n_9),
.Y(n_229)
);

AOI22xp33_ASAP7_75t_SL g231 ( 
.A1(n_160),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_231)
);

INVxp67_ASAP7_75t_L g263 ( 
.A(n_231),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_169),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_234),
.A2(n_152),
.B1(n_161),
.B2(n_192),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_193),
.B(n_179),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_SL g278 ( 
.A(n_239),
.B(n_249),
.Y(n_278)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_228),
.Y(n_240)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_240),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_216),
.B(n_146),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_243),
.B(n_260),
.Y(n_298)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_204),
.Y(n_244)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_244),
.Y(n_297)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_204),
.Y(n_245)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_245),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_L g292 ( 
.A1(n_246),
.A2(n_247),
.B1(n_269),
.B2(n_208),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_206),
.A2(n_170),
.B1(n_143),
.B2(n_150),
.Y(n_247)
);

AOI22xp33_ASAP7_75t_SL g248 ( 
.A1(n_233),
.A2(n_190),
.B1(n_186),
.B2(n_182),
.Y(n_248)
);

INVxp67_ASAP7_75t_L g286 ( 
.A(n_248),
.Y(n_286)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_214),
.Y(n_251)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_251),
.Y(n_310)
);

INVx4_ASAP7_75t_L g252 ( 
.A(n_218),
.Y(n_252)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_252),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_217),
.B(n_171),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_253),
.B(n_254),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_200),
.B(n_148),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_198),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_255),
.B(n_259),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_197),
.B(n_153),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g281 ( 
.A(n_256),
.B(n_257),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_SL g257 ( 
.A(n_202),
.B(n_173),
.Y(n_257)
);

OR2x2_ASAP7_75t_L g258 ( 
.A(n_203),
.B(n_154),
.Y(n_258)
);

OAI21xp5_ASAP7_75t_L g300 ( 
.A1(n_258),
.A2(n_276),
.B(n_222),
.Y(n_300)
);

INVxp33_ASAP7_75t_L g259 ( 
.A(n_223),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_207),
.B(n_202),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_213),
.B(n_220),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_261),
.B(n_264),
.Y(n_305)
);

AOI21xp5_ASAP7_75t_L g294 ( 
.A1(n_265),
.A2(n_266),
.B(n_275),
.Y(n_294)
);

OAI21xp5_ASAP7_75t_SL g266 ( 
.A1(n_213),
.A2(n_159),
.B(n_162),
.Y(n_266)
);

OAI22xp33_ASAP7_75t_SL g267 ( 
.A1(n_206),
.A2(n_183),
.B1(n_178),
.B2(n_180),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_267),
.B(n_273),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_233),
.A2(n_162),
.B1(n_180),
.B2(n_163),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_268),
.B(n_272),
.Y(n_312)
);

CKINVDCx16_ASAP7_75t_R g270 ( 
.A(n_219),
.Y(n_270)
);

CKINVDCx16_ASAP7_75t_R g285 ( 
.A(n_270),
.Y(n_285)
);

INVx6_ASAP7_75t_L g271 ( 
.A(n_235),
.Y(n_271)
);

BUFx3_ASAP7_75t_L g303 ( 
.A(n_271),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_207),
.A2(n_201),
.B1(n_215),
.B2(n_232),
.Y(n_272)
);

CKINVDCx16_ASAP7_75t_R g273 ( 
.A(n_205),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_214),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_274),
.Y(n_290)
);

OAI21xp5_ASAP7_75t_SL g275 ( 
.A1(n_205),
.A2(n_210),
.B(n_203),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_205),
.B(n_230),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g277 ( 
.A(n_226),
.B(n_237),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_277),
.B(n_235),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_246),
.A2(n_225),
.B1(n_226),
.B2(n_237),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_279),
.A2(n_292),
.B1(n_295),
.B2(n_301),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_261),
.B(n_230),
.C(n_196),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_282),
.B(n_287),
.C(n_289),
.Y(n_330)
);

XOR2x2_ASAP7_75t_L g283 ( 
.A(n_260),
.B(n_229),
.Y(n_283)
);

XOR2xp5_ASAP7_75t_L g322 ( 
.A(n_283),
.B(n_253),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_266),
.B(n_212),
.C(n_224),
.Y(n_287)
);

OAI21xp5_ASAP7_75t_SL g288 ( 
.A1(n_270),
.A2(n_199),
.B(n_224),
.Y(n_288)
);

OAI21xp5_ASAP7_75t_SL g318 ( 
.A1(n_288),
.A2(n_293),
.B(n_256),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_250),
.B(n_227),
.C(n_195),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g320 ( 
.A(n_291),
.B(n_244),
.Y(n_320)
);

NOR2x1_ASAP7_75t_R g293 ( 
.A(n_275),
.B(n_227),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_L g295 ( 
.A1(n_240),
.A2(n_208),
.B1(n_209),
.B2(n_195),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_SL g337 ( 
.A(n_300),
.B(n_285),
.Y(n_337)
);

OAI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_247),
.A2(n_236),
.B1(n_194),
.B2(n_222),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_L g302 ( 
.A1(n_242),
.A2(n_194),
.B1(n_236),
.B2(n_262),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_302),
.A2(n_304),
.B1(n_309),
.B2(n_267),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_242),
.A2(n_243),
.B1(n_241),
.B2(n_272),
.Y(n_304)
);

OAI21xp5_ASAP7_75t_L g306 ( 
.A1(n_258),
.A2(n_241),
.B(n_238),
.Y(n_306)
);

AND2x2_ASAP7_75t_L g336 ( 
.A(n_306),
.B(n_311),
.Y(n_336)
);

OAI22xp5_ASAP7_75t_L g309 ( 
.A1(n_273),
.A2(n_249),
.B1(n_255),
.B2(n_258),
.Y(n_309)
);

OAI21xp5_ASAP7_75t_L g311 ( 
.A1(n_238),
.A2(n_257),
.B(n_276),
.Y(n_311)
);

BUFx6f_ASAP7_75t_L g314 ( 
.A(n_303),
.Y(n_314)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_314),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_280),
.B(n_239),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_SL g343 ( 
.A(n_315),
.B(n_324),
.Y(n_343)
);

AOI22xp5_ASAP7_75t_SL g316 ( 
.A1(n_292),
.A2(n_286),
.B1(n_263),
.B2(n_309),
.Y(n_316)
);

OAI21xp5_ASAP7_75t_SL g358 ( 
.A1(n_316),
.A2(n_288),
.B(n_290),
.Y(n_358)
);

OAI22xp5_ASAP7_75t_L g341 ( 
.A1(n_317),
.A2(n_319),
.B1(n_329),
.B2(n_332),
.Y(n_341)
);

OAI21xp5_ASAP7_75t_L g362 ( 
.A1(n_318),
.A2(n_290),
.B(n_291),
.Y(n_362)
);

AOI22xp5_ASAP7_75t_L g319 ( 
.A1(n_312),
.A2(n_264),
.B1(n_250),
.B2(n_265),
.Y(n_319)
);

INVxp67_ASAP7_75t_L g345 ( 
.A(n_320),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_296),
.B(n_277),
.Y(n_321)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_321),
.Y(n_342)
);

XNOR2xp5_ASAP7_75t_L g348 ( 
.A(n_322),
.B(n_283),
.Y(n_348)
);

OAI22xp5_ASAP7_75t_SL g323 ( 
.A1(n_312),
.A2(n_269),
.B1(n_254),
.B2(n_274),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_323),
.B(n_327),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_278),
.B(n_271),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_296),
.B(n_245),
.Y(n_325)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_325),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_SL g326 ( 
.A(n_284),
.B(n_251),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_SL g350 ( 
.A(n_326),
.B(n_338),
.Y(n_350)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_295),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_297),
.Y(n_328)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_328),
.Y(n_359)
);

OAI22xp5_ASAP7_75t_L g329 ( 
.A1(n_278),
.A2(n_252),
.B1(n_271),
.B2(n_268),
.Y(n_329)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_297),
.Y(n_331)
);

INVx2_ASAP7_75t_L g357 ( 
.A(n_331),
.Y(n_357)
);

OAI22xp5_ASAP7_75t_L g332 ( 
.A1(n_305),
.A2(n_252),
.B1(n_306),
.B2(n_307),
.Y(n_332)
);

AOI22xp5_ASAP7_75t_L g333 ( 
.A1(n_279),
.A2(n_304),
.B1(n_305),
.B2(n_302),
.Y(n_333)
);

OAI22xp5_ASAP7_75t_L g363 ( 
.A1(n_333),
.A2(n_303),
.B1(n_308),
.B2(n_313),
.Y(n_363)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_299),
.Y(n_334)
);

INVxp67_ASAP7_75t_L g347 ( 
.A(n_334),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_289),
.B(n_282),
.C(n_287),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g351 ( 
.A(n_335),
.B(n_294),
.C(n_298),
.Y(n_351)
);

INVxp67_ASAP7_75t_L g361 ( 
.A(n_337),
.Y(n_361)
);

NOR3xp33_ASAP7_75t_SL g338 ( 
.A(n_307),
.B(n_293),
.C(n_310),
.Y(n_338)
);

OAI21xp33_ASAP7_75t_SL g339 ( 
.A1(n_286),
.A2(n_294),
.B(n_300),
.Y(n_339)
);

AO21x1_ASAP7_75t_L g360 ( 
.A1(n_339),
.A2(n_301),
.B(n_310),
.Y(n_360)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_299),
.Y(n_340)
);

HB1xp67_ASAP7_75t_L g349 ( 
.A(n_340),
.Y(n_349)
);

OAI22xp5_ASAP7_75t_SL g346 ( 
.A1(n_333),
.A2(n_316),
.B1(n_317),
.B2(n_319),
.Y(n_346)
);

AOI22xp5_ASAP7_75t_L g365 ( 
.A1(n_346),
.A2(n_363),
.B1(n_323),
.B2(n_327),
.Y(n_365)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_348),
.B(n_351),
.C(n_355),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_336),
.B(n_281),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_SL g377 ( 
.A(n_353),
.B(n_328),
.Y(n_377)
);

MAJIxp5_ASAP7_75t_L g355 ( 
.A(n_330),
.B(n_298),
.C(n_311),
.Y(n_355)
);

CKINVDCx20_ASAP7_75t_R g356 ( 
.A(n_325),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_356),
.B(n_338),
.Y(n_378)
);

INVxp67_ASAP7_75t_L g381 ( 
.A(n_358),
.Y(n_381)
);

INVx1_ASAP7_75t_SL g367 ( 
.A(n_360),
.Y(n_367)
);

HB1xp67_ASAP7_75t_L g368 ( 
.A(n_362),
.Y(n_368)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_365),
.Y(n_398)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_349),
.Y(n_366)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_366),
.Y(n_390)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_357),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_369),
.B(n_370),
.Y(n_384)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_357),
.Y(n_370)
);

CKINVDCx20_ASAP7_75t_R g371 ( 
.A(n_343),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_SL g383 ( 
.A(n_371),
.B(n_379),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_350),
.B(n_336),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_SL g386 ( 
.A(n_372),
.B(n_377),
.Y(n_386)
);

AOI22xp5_ASAP7_75t_L g373 ( 
.A1(n_341),
.A2(n_336),
.B1(n_321),
.B2(n_337),
.Y(n_373)
);

HB1xp67_ASAP7_75t_L g388 ( 
.A(n_373),
.Y(n_388)
);

MAJIxp5_ASAP7_75t_L g374 ( 
.A(n_351),
.B(n_330),
.C(n_335),
.Y(n_374)
);

MAJIxp5_ASAP7_75t_L g391 ( 
.A(n_374),
.B(n_375),
.C(n_376),
.Y(n_391)
);

MAJIxp5_ASAP7_75t_L g375 ( 
.A(n_355),
.B(n_322),
.C(n_318),
.Y(n_375)
);

MAJIxp5_ASAP7_75t_L g376 ( 
.A(n_348),
.B(n_313),
.C(n_331),
.Y(n_376)
);

CKINVDCx20_ASAP7_75t_R g385 ( 
.A(n_378),
.Y(n_385)
);

CKINVDCx20_ASAP7_75t_R g379 ( 
.A(n_356),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_L g380 ( 
.A(n_345),
.B(n_314),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_L g393 ( 
.A(n_380),
.B(n_354),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_347),
.B(n_334),
.Y(n_382)
);

CKINVDCx20_ASAP7_75t_R g392 ( 
.A(n_382),
.Y(n_392)
);

OAI21xp5_ASAP7_75t_SL g387 ( 
.A1(n_381),
.A2(n_352),
.B(n_361),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_387),
.B(n_394),
.Y(n_401)
);

XOR2xp5_ASAP7_75t_L g389 ( 
.A(n_376),
.B(n_358),
.Y(n_389)
);

XOR2xp5_ASAP7_75t_L g399 ( 
.A(n_389),
.B(n_375),
.Y(n_399)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_393),
.Y(n_402)
);

INVxp33_ASAP7_75t_L g394 ( 
.A(n_382),
.Y(n_394)
);

AOI22xp5_ASAP7_75t_L g395 ( 
.A1(n_367),
.A2(n_346),
.B1(n_352),
.B2(n_361),
.Y(n_395)
);

OAI22xp5_ASAP7_75t_SL g409 ( 
.A1(n_395),
.A2(n_397),
.B1(n_360),
.B2(n_367),
.Y(n_409)
);

XNOR2xp5_ASAP7_75t_L g396 ( 
.A(n_364),
.B(n_362),
.Y(n_396)
);

XNOR2xp5_ASAP7_75t_L g400 ( 
.A(n_396),
.B(n_364),
.Y(n_400)
);

AOI22xp5_ASAP7_75t_SL g397 ( 
.A1(n_381),
.A2(n_344),
.B1(n_342),
.B2(n_345),
.Y(n_397)
);

MAJx2_ASAP7_75t_L g417 ( 
.A(n_399),
.B(n_400),
.C(n_407),
.Y(n_417)
);

MAJIxp5_ASAP7_75t_L g403 ( 
.A(n_391),
.B(n_374),
.C(n_396),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_403),
.B(n_404),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_SL g404 ( 
.A(n_383),
.B(n_378),
.Y(n_404)
);

MAJIxp5_ASAP7_75t_L g405 ( 
.A(n_391),
.B(n_368),
.C(n_373),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_405),
.B(n_406),
.Y(n_416)
);

INVxp67_ASAP7_75t_L g406 ( 
.A(n_387),
.Y(n_406)
);

MAJIxp5_ASAP7_75t_L g407 ( 
.A(n_389),
.B(n_365),
.C(n_369),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_SL g408 ( 
.A(n_386),
.B(n_366),
.Y(n_408)
);

OAI22xp5_ASAP7_75t_SL g411 ( 
.A1(n_408),
.A2(n_397),
.B1(n_390),
.B2(n_392),
.Y(n_411)
);

AOI22xp5_ASAP7_75t_L g415 ( 
.A1(n_409),
.A2(n_394),
.B1(n_384),
.B2(n_347),
.Y(n_415)
);

AOI22xp5_ASAP7_75t_L g410 ( 
.A1(n_406),
.A2(n_388),
.B1(n_398),
.B2(n_385),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_L g420 ( 
.A(n_410),
.B(n_415),
.Y(n_420)
);

NOR2xp67_ASAP7_75t_SL g422 ( 
.A(n_411),
.B(n_412),
.Y(n_422)
);

NOR2xp67_ASAP7_75t_L g412 ( 
.A(n_403),
.B(n_342),
.Y(n_412)
);

OAI22xp5_ASAP7_75t_SL g413 ( 
.A1(n_402),
.A2(n_398),
.B1(n_395),
.B2(n_344),
.Y(n_413)
);

MAJIxp5_ASAP7_75t_L g418 ( 
.A(n_413),
.B(n_407),
.C(n_401),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_418),
.B(n_419),
.Y(n_424)
);

MAJIxp5_ASAP7_75t_L g419 ( 
.A(n_414),
.B(n_400),
.C(n_405),
.Y(n_419)
);

MAJIxp5_ASAP7_75t_L g421 ( 
.A(n_417),
.B(n_399),
.C(n_384),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_SL g423 ( 
.A(n_421),
.B(n_416),
.Y(n_423)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_423),
.Y(n_427)
);

AOI21xp5_ASAP7_75t_L g425 ( 
.A1(n_422),
.A2(n_410),
.B(n_415),
.Y(n_425)
);

AO21x1_ASAP7_75t_L g426 ( 
.A1(n_425),
.A2(n_420),
.B(n_370),
.Y(n_426)
);

NOR2xp33_ASAP7_75t_L g428 ( 
.A(n_426),
.B(n_427),
.Y(n_428)
);

MAJIxp5_ASAP7_75t_L g429 ( 
.A(n_428),
.B(n_424),
.C(n_417),
.Y(n_429)
);

AOI21xp33_ASAP7_75t_L g430 ( 
.A1(n_429),
.A2(n_359),
.B(n_340),
.Y(n_430)
);

MAJIxp5_ASAP7_75t_L g431 ( 
.A(n_430),
.B(n_359),
.C(n_354),
.Y(n_431)
);

XNOR2xp5_ASAP7_75t_L g432 ( 
.A(n_431),
.B(n_308),
.Y(n_432)
);


endmodule