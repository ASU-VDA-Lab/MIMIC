module fake_jpeg_14866_n_111 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_111);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_111;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_30;
wire n_106;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_1),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_1),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_SL g15 ( 
.A(n_11),
.B(n_8),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_12),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_4),
.B(n_5),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_12),
.Y(n_21)
);

INVx11_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_SL g24 ( 
.A(n_2),
.B(n_4),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_17),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_SL g47 ( 
.A(n_26),
.B(n_32),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_17),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_27),
.Y(n_39)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_22),
.Y(n_28)
);

INVx5_ASAP7_75t_L g42 ( 
.A(n_28),
.Y(n_42)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_18),
.Y(n_29)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_29),
.Y(n_45)
);

OAI21xp33_ASAP7_75t_L g30 ( 
.A1(n_15),
.A2(n_0),
.B(n_2),
.Y(n_30)
);

AND2x2_ASAP7_75t_L g36 ( 
.A(n_30),
.B(n_34),
.Y(n_36)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_17),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_31),
.B(n_35),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_SL g32 ( 
.A1(n_18),
.A2(n_0),
.B1(n_3),
.B2(n_6),
.Y(n_32)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_19),
.Y(n_33)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_33),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_15),
.B(n_3),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_L g35 ( 
.A1(n_19),
.A2(n_6),
.B1(n_7),
.B2(n_9),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_37),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_34),
.B(n_24),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_40),
.B(n_21),
.Y(n_58)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_28),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_43),
.B(n_44),
.Y(n_52)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_27),
.Y(n_44)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_27),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_46),
.B(n_48),
.Y(n_54)
);

BUFx2_ASAP7_75t_L g48 ( 
.A(n_29),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_33),
.B(n_24),
.Y(n_49)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_49),
.Y(n_63)
);

XOR2xp5_ASAP7_75t_L g50 ( 
.A(n_36),
.B(n_35),
.Y(n_50)
);

XNOR2xp5_ASAP7_75t_L g68 ( 
.A(n_50),
.B(n_55),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_36),
.B(n_20),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_51),
.B(n_56),
.Y(n_74)
);

NOR2xp67_ASAP7_75t_L g53 ( 
.A(n_38),
.B(n_20),
.Y(n_53)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_53),
.B(n_57),
.Y(n_71)
);

XNOR2xp5_ASAP7_75t_L g55 ( 
.A(n_47),
.B(n_33),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_41),
.B(n_21),
.Y(n_56)
);

NOR2x1_ASAP7_75t_SL g57 ( 
.A(n_48),
.B(n_25),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_58),
.B(n_66),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_44),
.A2(n_31),
.B1(n_26),
.B2(n_46),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_59),
.A2(n_60),
.B1(n_62),
.B2(n_39),
.Y(n_73)
);

AND2x2_ASAP7_75t_L g60 ( 
.A(n_45),
.B(n_31),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g62 ( 
.A1(n_41),
.A2(n_43),
.B1(n_42),
.B2(n_39),
.Y(n_62)
);

INVxp67_ASAP7_75t_L g64 ( 
.A(n_37),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_64),
.B(n_22),
.Y(n_76)
);

OAI21xp5_ASAP7_75t_SL g65 ( 
.A1(n_42),
.A2(n_14),
.B(n_13),
.Y(n_65)
);

CKINVDCx16_ASAP7_75t_R g70 ( 
.A(n_65),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_37),
.B(n_14),
.Y(n_66)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_54),
.Y(n_69)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_69),
.Y(n_81)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_65),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_72),
.Y(n_83)
);

INVx1_ASAP7_75t_SL g79 ( 
.A(n_73),
.Y(n_79)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_52),
.Y(n_75)
);

OAI21xp5_ASAP7_75t_SL g82 ( 
.A1(n_75),
.A2(n_76),
.B(n_64),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_63),
.B(n_13),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_77),
.B(n_78),
.Y(n_86)
);

CKINVDCx16_ASAP7_75t_R g78 ( 
.A(n_61),
.Y(n_78)
);

XOR2xp5_ASAP7_75t_L g80 ( 
.A(n_68),
.B(n_50),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_80),
.B(n_84),
.C(n_85),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_82),
.B(n_88),
.Y(n_89)
);

XNOR2xp5_ASAP7_75t_SL g84 ( 
.A(n_68),
.B(n_55),
.Y(n_84)
);

XNOR2xp5_ASAP7_75t_L g85 ( 
.A(n_67),
.B(n_57),
.Y(n_85)
);

XOR2xp5_ASAP7_75t_L g87 ( 
.A(n_71),
.B(n_60),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_87),
.B(n_69),
.C(n_74),
.Y(n_93)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_75),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_79),
.A2(n_70),
.B1(n_71),
.B2(n_73),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_90),
.A2(n_92),
.B1(n_79),
.B2(n_83),
.Y(n_98)
);

CKINVDCx14_ASAP7_75t_R g92 ( 
.A(n_86),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_93),
.B(n_94),
.C(n_87),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_84),
.B(n_62),
.C(n_59),
.Y(n_94)
);

BUFx12_ASAP7_75t_L g95 ( 
.A(n_88),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_95),
.B(n_81),
.Y(n_99)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_89),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_96),
.B(n_97),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_98),
.A2(n_99),
.B1(n_7),
.B2(n_16),
.Y(n_104)
);

BUFx24_ASAP7_75t_SL g100 ( 
.A(n_92),
.Y(n_100)
);

MAJx2_ASAP7_75t_L g102 ( 
.A(n_100),
.B(n_91),
.C(n_95),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_102),
.B(n_25),
.Y(n_106)
);

MAJx2_ASAP7_75t_L g103 ( 
.A(n_97),
.B(n_60),
.C(n_10),
.Y(n_103)
);

AOI21xp5_ASAP7_75t_L g107 ( 
.A1(n_103),
.A2(n_16),
.B(n_23),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_104),
.B(n_16),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_105),
.A2(n_107),
.B1(n_101),
.B2(n_23),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_106),
.B(n_23),
.Y(n_109)
);

BUFx24_ASAP7_75t_SL g110 ( 
.A(n_108),
.Y(n_110)
);

XOR2xp5_ASAP7_75t_L g111 ( 
.A(n_110),
.B(n_109),
.Y(n_111)
);


endmodule