module fake_netlist_6_4663_n_742 (n_52, n_16, n_1, n_91, n_119, n_46, n_18, n_21, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_138, n_22, n_68, n_28, n_50, n_49, n_7, n_83, n_5, n_101, n_127, n_125, n_77, n_106, n_92, n_42, n_133, n_96, n_8, n_90, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_75, n_109, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_742);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_18;
input n_21;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_138;
input n_22;
input n_68;
input n_28;
input n_50;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_127;
input n_125;
input n_77;
input n_106;
input n_92;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_75;
input n_109;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_742;

wire n_591;
wire n_435;
wire n_326;
wire n_256;
wire n_440;
wire n_587;
wire n_695;
wire n_507;
wire n_580;
wire n_209;
wire n_367;
wire n_465;
wire n_680;
wire n_741;
wire n_590;
wire n_625;
wire n_661;
wire n_223;
wire n_278;
wire n_341;
wire n_362;
wire n_148;
wire n_226;
wire n_161;
wire n_208;
wire n_462;
wire n_671;
wire n_607;
wire n_726;
wire n_316;
wire n_419;
wire n_304;
wire n_212;
wire n_700;
wire n_694;
wire n_740;
wire n_578;
wire n_703;
wire n_144;
wire n_365;
wire n_168;
wire n_384;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_342;
wire n_725;
wire n_358;
wire n_160;
wire n_449;
wire n_188;
wire n_310;
wire n_509;
wire n_186;
wire n_245;
wire n_368;
wire n_575;
wire n_677;
wire n_396;
wire n_495;
wire n_350;
wire n_585;
wire n_732;
wire n_568;
wire n_392;
wire n_442;
wire n_480;
wire n_724;
wire n_382;
wire n_673;
wire n_180;
wire n_628;
wire n_557;
wire n_349;
wire n_643;
wire n_233;
wire n_698;
wire n_617;
wire n_255;
wire n_739;
wire n_284;
wire n_400;
wire n_337;
wire n_214;
wire n_485;
wire n_443;
wire n_246;
wire n_471;
wire n_289;
wire n_421;
wire n_424;
wire n_615;
wire n_181;
wire n_182;
wire n_238;
wire n_573;
wire n_202;
wire n_320;
wire n_639;
wire n_676;
wire n_327;
wire n_727;
wire n_369;
wire n_597;
wire n_685;
wire n_280;
wire n_287;
wire n_353;
wire n_610;
wire n_555;
wire n_389;
wire n_415;
wire n_230;
wire n_605;
wire n_461;
wire n_383;
wire n_669;
wire n_200;
wire n_447;
wire n_176;
wire n_198;
wire n_300;
wire n_222;
wire n_179;
wire n_248;
wire n_517;
wire n_718;
wire n_667;
wire n_229;
wire n_542;
wire n_644;
wire n_682;
wire n_621;
wire n_305;
wire n_721;
wire n_532;
wire n_173;
wire n_691;
wire n_535;
wire n_250;
wire n_372;
wire n_468;
wire n_544;
wire n_504;
wire n_314;
wire n_378;
wire n_413;
wire n_377;
wire n_183;
wire n_510;
wire n_375;
wire n_601;
wire n_338;
wire n_522;
wire n_466;
wire n_704;
wire n_506;
wire n_360;
wire n_603;
wire n_235;
wire n_536;
wire n_622;
wire n_147;
wire n_191;
wire n_340;
wire n_710;
wire n_387;
wire n_452;
wire n_616;
wire n_658;
wire n_344;
wire n_581;
wire n_428;
wire n_609;
wire n_432;
wire n_641;
wire n_693;
wire n_167;
wire n_631;
wire n_174;
wire n_516;
wire n_153;
wire n_720;
wire n_525;
wire n_611;
wire n_156;
wire n_491;
wire n_145;
wire n_656;
wire n_666;
wire n_371;
wire n_567;
wire n_189;
wire n_738;
wire n_405;
wire n_213;
wire n_538;
wire n_294;
wire n_302;
wire n_499;
wire n_380;
wire n_705;
wire n_647;
wire n_197;
wire n_343;
wire n_448;
wire n_494;
wire n_539;
wire n_493;
wire n_397;
wire n_155;
wire n_614;
wire n_529;
wire n_445;
wire n_425;
wire n_684;
wire n_454;
wire n_218;
wire n_638;
wire n_234;
wire n_486;
wire n_381;
wire n_236;
wire n_653;
wire n_172;
wire n_713;
wire n_648;
wire n_657;
wire n_576;
wire n_472;
wire n_270;
wire n_239;
wire n_414;
wire n_563;
wire n_490;
wire n_290;
wire n_220;
wire n_224;
wire n_734;
wire n_708;
wire n_196;
wire n_402;
wire n_352;
wire n_668;
wire n_478;
wire n_626;
wire n_574;
wire n_460;
wire n_417;
wire n_446;
wire n_498;
wire n_662;
wire n_374;
wire n_659;
wire n_709;
wire n_366;
wire n_407;
wire n_450;
wire n_272;
wire n_526;
wire n_185;
wire n_712;
wire n_348;
wire n_711;
wire n_579;
wire n_376;
wire n_390;
wire n_473;
wire n_293;
wire n_334;
wire n_559;
wire n_370;
wire n_458;
wire n_232;
wire n_650;
wire n_163;
wire n_717;
wire n_330;
wire n_470;
wire n_475;
wire n_298;
wire n_492;
wire n_281;
wire n_258;
wire n_551;
wire n_154;
wire n_699;
wire n_456;
wire n_564;
wire n_260;
wire n_265;
wire n_313;
wire n_451;
wire n_624;
wire n_279;
wire n_686;
wire n_252;
wire n_228;
wire n_594;
wire n_565;
wire n_719;
wire n_356;
wire n_577;
wire n_166;
wire n_184;
wire n_552;
wire n_619;
wire n_216;
wire n_455;
wire n_521;
wire n_363;
wire n_572;
wire n_395;
wire n_592;
wire n_654;
wire n_323;
wire n_606;
wire n_393;
wire n_411;
wire n_503;
wire n_716;
wire n_152;
wire n_623;
wire n_599;
wire n_513;
wire n_321;
wire n_645;
wire n_331;
wire n_227;
wire n_570;
wire n_731;
wire n_406;
wire n_483;
wire n_735;
wire n_204;
wire n_482;
wire n_474;
wire n_527;
wire n_261;
wire n_608;
wire n_620;
wire n_420;
wire n_683;
wire n_630;
wire n_312;
wire n_394;
wire n_519;
wire n_541;
wire n_512;
wire n_164;
wire n_292;
wire n_307;
wire n_469;
wire n_433;
wire n_500;
wire n_476;
wire n_714;
wire n_291;
wire n_219;
wire n_543;
wire n_357;
wire n_150;
wire n_264;
wire n_263;
wire n_589;
wire n_481;
wire n_325;
wire n_329;
wire n_464;
wire n_600;
wire n_561;
wire n_477;
wire n_549;
wire n_533;
wire n_408;
wire n_237;
wire n_584;
wire n_244;
wire n_399;
wire n_243;
wire n_548;
wire n_282;
wire n_436;
wire n_211;
wire n_523;
wire n_175;
wire n_322;
wire n_707;
wire n_345;
wire n_409;
wire n_231;
wire n_354;
wire n_689;
wire n_505;
wire n_240;
wire n_319;
wire n_547;
wire n_537;
wire n_273;
wire n_558;
wire n_635;
wire n_311;
wire n_403;
wire n_723;
wire n_253;
wire n_634;
wire n_583;
wire n_596;
wire n_546;
wire n_562;
wire n_249;
wire n_201;
wire n_386;
wire n_556;
wire n_159;
wire n_157;
wire n_162;
wire n_692;
wire n_733;
wire n_487;
wire n_550;
wire n_241;
wire n_275;
wire n_553;
wire n_652;
wire n_560;
wire n_642;
wire n_276;
wire n_569;
wire n_441;
wire n_221;
wire n_444;
wire n_586;
wire n_423;
wire n_146;
wire n_737;
wire n_318;
wire n_303;
wire n_511;
wire n_715;
wire n_467;
wire n_306;
wire n_193;
wire n_269;
wire n_359;
wire n_346;
wire n_416;
wire n_530;
wire n_277;
wire n_520;
wire n_418;
wire n_618;
wire n_582;
wire n_199;
wire n_266;
wire n_296;
wire n_674;
wire n_571;
wire n_268;
wire n_271;
wire n_404;
wire n_651;
wire n_439;
wire n_158;
wire n_217;
wire n_210;
wire n_299;
wire n_518;
wire n_206;
wire n_679;
wire n_453;
wire n_612;
wire n_633;
wire n_665;
wire n_333;
wire n_588;
wire n_215;
wire n_178;
wire n_247;
wire n_225;
wire n_308;
wire n_309;
wire n_355;
wire n_426;
wire n_317;
wire n_149;
wire n_632;
wire n_702;
wire n_431;
wire n_347;
wire n_459;
wire n_502;
wire n_328;
wire n_672;
wire n_534;
wire n_488;
wire n_429;
wire n_373;
wire n_195;
wire n_285;
wire n_497;
wire n_675;
wire n_257;
wire n_730;
wire n_655;
wire n_706;
wire n_670;
wire n_203;
wire n_286;
wire n_254;
wire n_207;
wire n_242;
wire n_690;
wire n_401;
wire n_324;
wire n_335;
wire n_430;
wire n_463;
wire n_545;
wire n_489;
wire n_205;
wire n_604;
wire n_251;
wire n_301;
wire n_274;
wire n_636;
wire n_728;
wire n_681;
wire n_729;
wire n_151;
wire n_412;
wire n_640;
wire n_660;
wire n_267;
wire n_438;
wire n_339;
wire n_315;
wire n_434;
wire n_515;
wire n_288;
wire n_427;
wire n_479;
wire n_496;
wire n_598;
wire n_422;
wire n_696;
wire n_688;
wire n_722;
wire n_165;
wire n_351;
wire n_437;
wire n_259;
wire n_177;
wire n_540;
wire n_593;
wire n_514;
wire n_646;
wire n_528;
wire n_391;
wire n_457;
wire n_687;
wire n_697;
wire n_364;
wire n_637;
wire n_295;
wire n_385;
wire n_701;
wire n_629;
wire n_388;
wire n_190;
wire n_262;
wire n_484;
wire n_613;
wire n_736;
wire n_187;
wire n_501;
wire n_531;
wire n_361;
wire n_508;
wire n_663;
wire n_379;
wire n_170;
wire n_332;
wire n_336;
wire n_398;
wire n_410;
wire n_566;
wire n_554;
wire n_602;
wire n_194;
wire n_664;
wire n_171;
wire n_678;
wire n_192;
wire n_169;
wire n_649;
wire n_283;

BUFx3_ASAP7_75t_L g144 ( 
.A(n_118),
.Y(n_144)
);

CKINVDCx5p33_ASAP7_75t_R g145 ( 
.A(n_76),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_130),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_17),
.Y(n_147)
);

CKINVDCx16_ASAP7_75t_R g148 ( 
.A(n_65),
.Y(n_148)
);

CKINVDCx5p33_ASAP7_75t_R g149 ( 
.A(n_20),
.Y(n_149)
);

CKINVDCx5p33_ASAP7_75t_R g150 ( 
.A(n_39),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_111),
.Y(n_151)
);

CKINVDCx5p33_ASAP7_75t_R g152 ( 
.A(n_53),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_85),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_81),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_95),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_90),
.Y(n_156)
);

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_115),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_100),
.Y(n_158)
);

NOR2xp67_ASAP7_75t_L g159 ( 
.A(n_78),
.B(n_73),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_9),
.Y(n_160)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_113),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_142),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_7),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_51),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_33),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_7),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_93),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_112),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_119),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_107),
.Y(n_170)
);

CKINVDCx16_ASAP7_75t_R g171 ( 
.A(n_101),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_59),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_0),
.Y(n_173)
);

INVxp67_ASAP7_75t_L g174 ( 
.A(n_94),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_79),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_63),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_124),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_42),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_132),
.Y(n_179)
);

OR2x2_ASAP7_75t_L g180 ( 
.A(n_136),
.B(n_88),
.Y(n_180)
);

NOR2xp67_ASAP7_75t_L g181 ( 
.A(n_122),
.B(n_2),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_98),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_89),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_24),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_80),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_75),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_43),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_99),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_11),
.Y(n_189)
);

BUFx3_ASAP7_75t_L g190 ( 
.A(n_97),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_11),
.Y(n_191)
);

NOR2xp67_ASAP7_75t_L g192 ( 
.A(n_127),
.B(n_52),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_120),
.Y(n_193)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_60),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_125),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_83),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_109),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_55),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_57),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_87),
.Y(n_200)
);

HB1xp67_ASAP7_75t_L g201 ( 
.A(n_163),
.Y(n_201)
);

OAI21x1_ASAP7_75t_L g202 ( 
.A1(n_161),
.A2(n_0),
.B(n_1),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g203 ( 
.A(n_151),
.Y(n_203)
);

OA21x2_ASAP7_75t_L g204 ( 
.A1(n_147),
.A2(n_1),
.B(n_2),
.Y(n_204)
);

BUFx6f_ASAP7_75t_L g205 ( 
.A(n_151),
.Y(n_205)
);

BUFx6f_ASAP7_75t_L g206 ( 
.A(n_151),
.Y(n_206)
);

CKINVDCx16_ASAP7_75t_R g207 ( 
.A(n_148),
.Y(n_207)
);

OA21x2_ASAP7_75t_L g208 ( 
.A1(n_160),
.A2(n_3),
.B(n_4),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_161),
.B(n_3),
.Y(n_209)
);

AND2x2_ASAP7_75t_L g210 ( 
.A(n_144),
.B(n_4),
.Y(n_210)
);

OAI22x1_ASAP7_75t_L g211 ( 
.A1(n_173),
.A2(n_5),
.B1(n_6),
.B2(n_8),
.Y(n_211)
);

BUFx2_ASAP7_75t_L g212 ( 
.A(n_189),
.Y(n_212)
);

INVx3_ASAP7_75t_L g213 ( 
.A(n_166),
.Y(n_213)
);

BUFx6f_ASAP7_75t_L g214 ( 
.A(n_151),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_166),
.Y(n_215)
);

INVx2_ASAP7_75t_SL g216 ( 
.A(n_166),
.Y(n_216)
);

AND2x2_ASAP7_75t_L g217 ( 
.A(n_144),
.B(n_190),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_166),
.Y(n_218)
);

BUFx12f_ASAP7_75t_L g219 ( 
.A(n_145),
.Y(n_219)
);

BUFx6f_ASAP7_75t_L g220 ( 
.A(n_190),
.Y(n_220)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_191),
.Y(n_221)
);

INVx5_ASAP7_75t_L g222 ( 
.A(n_194),
.Y(n_222)
);

BUFx6f_ASAP7_75t_L g223 ( 
.A(n_194),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_171),
.B(n_5),
.Y(n_224)
);

AND2x6_ASAP7_75t_L g225 ( 
.A(n_146),
.B(n_143),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_153),
.Y(n_226)
);

OA21x2_ASAP7_75t_L g227 ( 
.A1(n_154),
.A2(n_158),
.B(n_155),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_164),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_181),
.B(n_6),
.Y(n_229)
);

OAI22x1_ASAP7_75t_R g230 ( 
.A1(n_162),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_230)
);

INVx2_ASAP7_75t_SL g231 ( 
.A(n_165),
.Y(n_231)
);

CKINVDCx11_ASAP7_75t_R g232 ( 
.A(n_162),
.Y(n_232)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_167),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_168),
.Y(n_234)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_170),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_SL g236 ( 
.A(n_176),
.B(n_10),
.Y(n_236)
);

HB1xp67_ASAP7_75t_L g237 ( 
.A(n_175),
.Y(n_237)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_177),
.Y(n_238)
);

INVx2_ASAP7_75t_SL g239 ( 
.A(n_178),
.Y(n_239)
);

AND2x2_ASAP7_75t_L g240 ( 
.A(n_184),
.B(n_187),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_200),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_176),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_242)
);

BUFx12f_ASAP7_75t_L g243 ( 
.A(n_149),
.Y(n_243)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_223),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_224),
.B(n_186),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_232),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_215),
.Y(n_247)
);

AND2x2_ASAP7_75t_SL g248 ( 
.A(n_236),
.B(n_180),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_215),
.Y(n_249)
);

BUFx6f_ASAP7_75t_L g250 ( 
.A(n_203),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_217),
.B(n_150),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_218),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_218),
.Y(n_253)
);

NAND3xp33_ASAP7_75t_L g254 ( 
.A(n_237),
.B(n_174),
.C(n_198),
.Y(n_254)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_223),
.Y(n_255)
);

AND2x2_ASAP7_75t_L g256 ( 
.A(n_217),
.B(n_152),
.Y(n_256)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_223),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_213),
.Y(n_258)
);

AND2x6_ASAP7_75t_L g259 ( 
.A(n_210),
.B(n_240),
.Y(n_259)
);

INVx3_ASAP7_75t_L g260 ( 
.A(n_203),
.Y(n_260)
);

BUFx10_ASAP7_75t_L g261 ( 
.A(n_201),
.Y(n_261)
);

INVx3_ASAP7_75t_L g262 ( 
.A(n_203),
.Y(n_262)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_223),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_213),
.Y(n_264)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_223),
.Y(n_265)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_213),
.Y(n_266)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_203),
.Y(n_267)
);

OAI22xp33_ASAP7_75t_L g268 ( 
.A1(n_242),
.A2(n_199),
.B1(n_186),
.B2(n_156),
.Y(n_268)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_203),
.Y(n_269)
);

INVxp67_ASAP7_75t_SL g270 ( 
.A(n_220),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_216),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_243),
.Y(n_272)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_205),
.Y(n_273)
);

NAND3xp33_ASAP7_75t_L g274 ( 
.A(n_210),
.B(n_185),
.C(n_197),
.Y(n_274)
);

NOR3xp33_ASAP7_75t_L g275 ( 
.A(n_229),
.B(n_209),
.C(n_207),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_216),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_220),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_220),
.Y(n_278)
);

AND2x2_ASAP7_75t_L g279 ( 
.A(n_240),
.B(n_157),
.Y(n_279)
);

NAND3xp33_ASAP7_75t_L g280 ( 
.A(n_220),
.B(n_183),
.C(n_196),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_220),
.Y(n_281)
);

OAI22xp33_ASAP7_75t_SL g282 ( 
.A1(n_212),
.A2(n_182),
.B1(n_195),
.B2(n_193),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_233),
.Y(n_283)
);

INVxp67_ASAP7_75t_R g284 ( 
.A(n_230),
.Y(n_284)
);

NAND2xp33_ASAP7_75t_SL g285 ( 
.A(n_211),
.B(n_199),
.Y(n_285)
);

AND3x2_ASAP7_75t_L g286 ( 
.A(n_212),
.B(n_192),
.C(n_159),
.Y(n_286)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_205),
.Y(n_287)
);

AND3x2_ASAP7_75t_L g288 ( 
.A(n_226),
.B(n_12),
.C(n_13),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_227),
.B(n_169),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_248),
.B(n_219),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_SL g291 ( 
.A(n_248),
.B(n_172),
.Y(n_291)
);

INVx4_ASAP7_75t_L g292 ( 
.A(n_259),
.Y(n_292)
);

AND2x2_ASAP7_75t_L g293 ( 
.A(n_256),
.B(n_231),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_259),
.B(n_227),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_251),
.B(n_219),
.Y(n_295)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_244),
.Y(n_296)
);

AND2x2_ASAP7_75t_SL g297 ( 
.A(n_275),
.B(n_204),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_256),
.B(n_243),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_271),
.Y(n_299)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_244),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_279),
.B(n_226),
.Y(n_301)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_255),
.Y(n_302)
);

NOR2xp67_ASAP7_75t_L g303 ( 
.A(n_280),
.B(n_274),
.Y(n_303)
);

NOR2xp67_ASAP7_75t_SL g304 ( 
.A(n_250),
.B(n_204),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_245),
.A2(n_225),
.B1(n_188),
.B2(n_179),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_245),
.A2(n_225),
.B1(n_211),
.B2(n_239),
.Y(n_306)
);

INVxp67_ASAP7_75t_SL g307 ( 
.A(n_253),
.Y(n_307)
);

INVxp33_ASAP7_75t_L g308 ( 
.A(n_279),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_270),
.B(n_222),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_277),
.B(n_222),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_278),
.B(n_222),
.Y(n_311)
);

BUFx3_ASAP7_75t_L g312 ( 
.A(n_276),
.Y(n_312)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_255),
.Y(n_313)
);

INVx4_ASAP7_75t_L g314 ( 
.A(n_260),
.Y(n_314)
);

INVx2_ASAP7_75t_SL g315 ( 
.A(n_261),
.Y(n_315)
);

BUFx6f_ASAP7_75t_SL g316 ( 
.A(n_261),
.Y(n_316)
);

NAND2xp33_ASAP7_75t_SL g317 ( 
.A(n_289),
.B(n_231),
.Y(n_317)
);

NOR2x1p5_ASAP7_75t_L g318 ( 
.A(n_272),
.B(n_221),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_SL g319 ( 
.A(n_272),
.B(n_225),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_281),
.B(n_222),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_258),
.Y(n_321)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_257),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_257),
.B(n_228),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_263),
.B(n_228),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_SL g325 ( 
.A(n_282),
.B(n_235),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_263),
.B(n_234),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_265),
.B(n_234),
.Y(n_327)
);

INVxp67_ASAP7_75t_L g328 ( 
.A(n_285),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_265),
.B(n_241),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_254),
.B(n_247),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_264),
.Y(n_331)
);

INVx2_ASAP7_75t_SL g332 ( 
.A(n_261),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_SL g333 ( 
.A(n_268),
.B(n_235),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_249),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_SL g335 ( 
.A(n_266),
.B(n_238),
.Y(n_335)
);

INVx6_ASAP7_75t_L g336 ( 
.A(n_250),
.Y(n_336)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_260),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_252),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_260),
.B(n_241),
.Y(n_339)
);

AO221x1_ASAP7_75t_L g340 ( 
.A1(n_285),
.A2(n_208),
.B1(n_204),
.B2(n_202),
.C(n_206),
.Y(n_340)
);

AOI22xp33_ASAP7_75t_L g341 ( 
.A1(n_286),
.A2(n_204),
.B1(n_208),
.B2(n_225),
.Y(n_341)
);

BUFx6f_ASAP7_75t_L g342 ( 
.A(n_250),
.Y(n_342)
);

INVx2_ASAP7_75t_SL g343 ( 
.A(n_288),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_262),
.B(n_238),
.Y(n_344)
);

NAND2xp33_ASAP7_75t_L g345 ( 
.A(n_267),
.B(n_225),
.Y(n_345)
);

BUFx3_ASAP7_75t_L g346 ( 
.A(n_266),
.Y(n_346)
);

INVx2_ASAP7_75t_L g347 ( 
.A(n_262),
.Y(n_347)
);

AOI22xp5_ASAP7_75t_L g348 ( 
.A1(n_283),
.A2(n_225),
.B1(n_239),
.B2(n_208),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_262),
.B(n_267),
.Y(n_349)
);

INVx11_ASAP7_75t_L g350 ( 
.A(n_316),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_308),
.B(n_246),
.Y(n_351)
);

OAI21x1_ASAP7_75t_L g352 ( 
.A1(n_294),
.A2(n_269),
.B(n_287),
.Y(n_352)
);

AOI211xp5_ASAP7_75t_L g353 ( 
.A1(n_333),
.A2(n_284),
.B(n_221),
.C(n_230),
.Y(n_353)
);

INVx2_ASAP7_75t_SL g354 ( 
.A(n_312),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_301),
.B(n_269),
.Y(n_355)
);

INVx3_ASAP7_75t_L g356 ( 
.A(n_346),
.Y(n_356)
);

AOI21xp5_ASAP7_75t_L g357 ( 
.A1(n_317),
.A2(n_273),
.B(n_205),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_301),
.B(n_253),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_307),
.Y(n_359)
);

HB1xp67_ASAP7_75t_L g360 ( 
.A(n_328),
.Y(n_360)
);

AOI21xp5_ASAP7_75t_L g361 ( 
.A1(n_309),
.A2(n_206),
.B(n_214),
.Y(n_361)
);

CKINVDCx14_ASAP7_75t_R g362 ( 
.A(n_298),
.Y(n_362)
);

NOR2xp67_ASAP7_75t_L g363 ( 
.A(n_315),
.B(n_246),
.Y(n_363)
);

AOI21xp5_ASAP7_75t_L g364 ( 
.A1(n_345),
.A2(n_206),
.B(n_214),
.Y(n_364)
);

AND2x6_ASAP7_75t_L g365 ( 
.A(n_348),
.B(n_206),
.Y(n_365)
);

INVx2_ASAP7_75t_L g366 ( 
.A(n_296),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_307),
.B(n_208),
.Y(n_367)
);

AOI21xp5_ASAP7_75t_L g368 ( 
.A1(n_349),
.A2(n_206),
.B(n_214),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_L g369 ( 
.A(n_291),
.B(n_14),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_293),
.B(n_214),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_306),
.B(n_214),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_291),
.B(n_15),
.Y(n_372)
);

AND2x2_ASAP7_75t_L g373 ( 
.A(n_332),
.B(n_318),
.Y(n_373)
);

INVx2_ASAP7_75t_SL g374 ( 
.A(n_299),
.Y(n_374)
);

INVx2_ASAP7_75t_SL g375 ( 
.A(n_325),
.Y(n_375)
);

INVx2_ASAP7_75t_L g376 ( 
.A(n_300),
.Y(n_376)
);

INVx2_ASAP7_75t_L g377 ( 
.A(n_302),
.Y(n_377)
);

AOI22xp33_ASAP7_75t_SL g378 ( 
.A1(n_297),
.A2(n_284),
.B1(n_16),
.B2(n_17),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_297),
.B(n_21),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_L g380 ( 
.A(n_328),
.B(n_15),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_334),
.B(n_22),
.Y(n_381)
);

BUFx8_ASAP7_75t_L g382 ( 
.A(n_316),
.Y(n_382)
);

A2O1A1Ixp33_ASAP7_75t_L g383 ( 
.A1(n_330),
.A2(n_16),
.B(n_18),
.C(n_19),
.Y(n_383)
);

NAND3xp33_ASAP7_75t_L g384 ( 
.A(n_325),
.B(n_341),
.C(n_330),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_338),
.B(n_303),
.Y(n_385)
);

AOI21xp5_ASAP7_75t_L g386 ( 
.A1(n_292),
.A2(n_82),
.B(n_140),
.Y(n_386)
);

AOI21xp33_ASAP7_75t_L g387 ( 
.A1(n_333),
.A2(n_18),
.B(n_19),
.Y(n_387)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_313),
.Y(n_388)
);

AND2x2_ASAP7_75t_L g389 ( 
.A(n_295),
.B(n_23),
.Y(n_389)
);

AOI22xp5_ASAP7_75t_L g390 ( 
.A1(n_295),
.A2(n_25),
.B1(n_26),
.B2(n_27),
.Y(n_390)
);

OR2x2_ASAP7_75t_L g391 ( 
.A(n_290),
.B(n_28),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_341),
.B(n_29),
.Y(n_392)
);

AOI22xp5_ASAP7_75t_L g393 ( 
.A1(n_305),
.A2(n_30),
.B1(n_31),
.B2(n_32),
.Y(n_393)
);

AOI21xp5_ASAP7_75t_L g394 ( 
.A1(n_292),
.A2(n_34),
.B(n_35),
.Y(n_394)
);

NOR2xp33_ASAP7_75t_L g395 ( 
.A(n_298),
.B(n_36),
.Y(n_395)
);

INVx2_ASAP7_75t_SL g396 ( 
.A(n_343),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_L g397 ( 
.A(n_321),
.B(n_37),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_340),
.B(n_38),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_L g399 ( 
.A(n_331),
.B(n_40),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_304),
.B(n_41),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_323),
.Y(n_401)
);

AOI21xp5_ASAP7_75t_L g402 ( 
.A1(n_344),
.A2(n_44),
.B(n_45),
.Y(n_402)
);

AOI21xp5_ASAP7_75t_L g403 ( 
.A1(n_324),
.A2(n_46),
.B(n_47),
.Y(n_403)
);

AOI21xp5_ASAP7_75t_L g404 ( 
.A1(n_326),
.A2(n_48),
.B(n_49),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_327),
.B(n_50),
.Y(n_405)
);

OAI21x1_ASAP7_75t_L g406 ( 
.A1(n_337),
.A2(n_54),
.B(n_56),
.Y(n_406)
);

AOI21xp5_ASAP7_75t_L g407 ( 
.A1(n_329),
.A2(n_58),
.B(n_61),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_339),
.Y(n_408)
);

AOI21xp5_ASAP7_75t_L g409 ( 
.A1(n_310),
.A2(n_62),
.B(n_64),
.Y(n_409)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_322),
.Y(n_410)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_347),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_335),
.Y(n_412)
);

AO21x1_ASAP7_75t_L g413 ( 
.A1(n_319),
.A2(n_66),
.B(n_67),
.Y(n_413)
);

BUFx6f_ASAP7_75t_L g414 ( 
.A(n_354),
.Y(n_414)
);

OAI22x1_ASAP7_75t_L g415 ( 
.A1(n_369),
.A2(n_335),
.B1(n_314),
.B2(n_320),
.Y(n_415)
);

AOI21x1_ASAP7_75t_L g416 ( 
.A1(n_367),
.A2(n_311),
.B(n_314),
.Y(n_416)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_366),
.Y(n_417)
);

AND2x4_ASAP7_75t_L g418 ( 
.A(n_374),
.B(n_342),
.Y(n_418)
);

OAI21x1_ASAP7_75t_L g419 ( 
.A1(n_352),
.A2(n_336),
.B(n_342),
.Y(n_419)
);

A2O1A1Ixp33_ASAP7_75t_L g420 ( 
.A1(n_372),
.A2(n_342),
.B(n_69),
.C(n_70),
.Y(n_420)
);

OAI21xp5_ASAP7_75t_L g421 ( 
.A1(n_384),
.A2(n_336),
.B(n_71),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_359),
.B(n_68),
.Y(n_422)
);

OAI21xp5_ASAP7_75t_L g423 ( 
.A1(n_384),
.A2(n_398),
.B(n_392),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_412),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_SL g425 ( 
.A(n_385),
.B(n_375),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_401),
.B(n_72),
.Y(n_426)
);

OAI21x1_ASAP7_75t_SL g427 ( 
.A1(n_413),
.A2(n_74),
.B(n_77),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_SL g428 ( 
.A(n_395),
.B(n_84),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_408),
.B(n_86),
.Y(n_429)
);

AND2x2_ASAP7_75t_L g430 ( 
.A(n_360),
.B(n_91),
.Y(n_430)
);

OAI21xp33_ASAP7_75t_SL g431 ( 
.A1(n_392),
.A2(n_141),
.B(n_92),
.Y(n_431)
);

CKINVDCx6p67_ASAP7_75t_R g432 ( 
.A(n_373),
.Y(n_432)
);

BUFx12f_ASAP7_75t_L g433 ( 
.A(n_382),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_376),
.Y(n_434)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_377),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_358),
.B(n_96),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_388),
.Y(n_437)
);

OAI21x1_ASAP7_75t_L g438 ( 
.A1(n_406),
.A2(n_102),
.B(n_103),
.Y(n_438)
);

OAI21x1_ASAP7_75t_L g439 ( 
.A1(n_400),
.A2(n_104),
.B(n_105),
.Y(n_439)
);

BUFx3_ASAP7_75t_L g440 ( 
.A(n_396),
.Y(n_440)
);

AOI221xp5_ASAP7_75t_L g441 ( 
.A1(n_387),
.A2(n_106),
.B1(n_108),
.B2(n_110),
.C(n_114),
.Y(n_441)
);

AO21x2_ASAP7_75t_L g442 ( 
.A1(n_379),
.A2(n_398),
.B(n_371),
.Y(n_442)
);

BUFx6f_ASAP7_75t_L g443 ( 
.A(n_356),
.Y(n_443)
);

BUFx12f_ASAP7_75t_L g444 ( 
.A(n_382),
.Y(n_444)
);

BUFx4f_ASAP7_75t_SL g445 ( 
.A(n_391),
.Y(n_445)
);

BUFx6f_ASAP7_75t_L g446 ( 
.A(n_356),
.Y(n_446)
);

OAI21x1_ASAP7_75t_L g447 ( 
.A1(n_364),
.A2(n_116),
.B(n_117),
.Y(n_447)
);

INVx2_ASAP7_75t_SL g448 ( 
.A(n_370),
.Y(n_448)
);

OAI22xp5_ASAP7_75t_L g449 ( 
.A1(n_378),
.A2(n_121),
.B1(n_123),
.B2(n_126),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_355),
.B(n_128),
.Y(n_450)
);

BUFx6f_ASAP7_75t_L g451 ( 
.A(n_381),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_389),
.B(n_129),
.Y(n_452)
);

AOI21xp5_ASAP7_75t_L g453 ( 
.A1(n_405),
.A2(n_131),
.B(n_133),
.Y(n_453)
);

OR2x2_ASAP7_75t_L g454 ( 
.A(n_351),
.B(n_134),
.Y(n_454)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_410),
.Y(n_455)
);

INVx1_ASAP7_75t_SL g456 ( 
.A(n_380),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_365),
.B(n_135),
.Y(n_457)
);

AOI21xp5_ASAP7_75t_L g458 ( 
.A1(n_405),
.A2(n_137),
.B(n_138),
.Y(n_458)
);

AND2x2_ASAP7_75t_L g459 ( 
.A(n_362),
.B(n_139),
.Y(n_459)
);

NAND2x1p5_ASAP7_75t_L g460 ( 
.A(n_393),
.B(n_390),
.Y(n_460)
);

CKINVDCx20_ASAP7_75t_R g461 ( 
.A(n_350),
.Y(n_461)
);

AOI22xp33_ASAP7_75t_L g462 ( 
.A1(n_387),
.A2(n_365),
.B1(n_411),
.B2(n_399),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_365),
.B(n_397),
.Y(n_463)
);

AOI21xp5_ASAP7_75t_L g464 ( 
.A1(n_357),
.A2(n_361),
.B(n_368),
.Y(n_464)
);

OAI21xp5_ASAP7_75t_L g465 ( 
.A1(n_423),
.A2(n_365),
.B(n_386),
.Y(n_465)
);

OAI21x1_ASAP7_75t_L g466 ( 
.A1(n_419),
.A2(n_394),
.B(n_402),
.Y(n_466)
);

AO21x2_ASAP7_75t_L g467 ( 
.A1(n_423),
.A2(n_421),
.B(n_442),
.Y(n_467)
);

OAI21x1_ASAP7_75t_L g468 ( 
.A1(n_438),
.A2(n_403),
.B(n_404),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_424),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_434),
.Y(n_470)
);

AO21x2_ASAP7_75t_L g471 ( 
.A1(n_421),
.A2(n_383),
.B(n_407),
.Y(n_471)
);

OAI21x1_ASAP7_75t_L g472 ( 
.A1(n_416),
.A2(n_409),
.B(n_363),
.Y(n_472)
);

AND2x4_ASAP7_75t_L g473 ( 
.A(n_443),
.B(n_446),
.Y(n_473)
);

HB1xp67_ASAP7_75t_L g474 ( 
.A(n_414),
.Y(n_474)
);

OAI21xp5_ASAP7_75t_L g475 ( 
.A1(n_463),
.A2(n_353),
.B(n_436),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_437),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_417),
.Y(n_477)
);

BUFx6f_ASAP7_75t_L g478 ( 
.A(n_443),
.Y(n_478)
);

OAI21xp5_ASAP7_75t_L g479 ( 
.A1(n_463),
.A2(n_353),
.B(n_436),
.Y(n_479)
);

AOI22x1_ASAP7_75t_L g480 ( 
.A1(n_415),
.A2(n_460),
.B1(n_427),
.B2(n_464),
.Y(n_480)
);

OAI21x1_ASAP7_75t_SL g481 ( 
.A1(n_429),
.A2(n_426),
.B(n_457),
.Y(n_481)
);

OAI21x1_ASAP7_75t_L g482 ( 
.A1(n_447),
.A2(n_439),
.B(n_450),
.Y(n_482)
);

NOR2xp67_ASAP7_75t_L g483 ( 
.A(n_454),
.B(n_455),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_456),
.B(n_425),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_435),
.Y(n_485)
);

AOI21xp33_ASAP7_75t_L g486 ( 
.A1(n_456),
.A2(n_452),
.B(n_426),
.Y(n_486)
);

OAI21x1_ASAP7_75t_L g487 ( 
.A1(n_450),
.A2(n_452),
.B(n_457),
.Y(n_487)
);

OAI21x1_ASAP7_75t_L g488 ( 
.A1(n_422),
.A2(n_429),
.B(n_460),
.Y(n_488)
);

AOI21xp5_ASAP7_75t_L g489 ( 
.A1(n_422),
.A2(n_451),
.B(n_428),
.Y(n_489)
);

INVx3_ASAP7_75t_L g490 ( 
.A(n_443),
.Y(n_490)
);

BUFx3_ASAP7_75t_L g491 ( 
.A(n_414),
.Y(n_491)
);

OAI222xp33_ASAP7_75t_L g492 ( 
.A1(n_449),
.A2(n_445),
.B1(n_462),
.B2(n_430),
.C1(n_459),
.C2(n_448),
.Y(n_492)
);

CKINVDCx20_ASAP7_75t_R g493 ( 
.A(n_461),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_418),
.Y(n_494)
);

AO21x2_ASAP7_75t_L g495 ( 
.A1(n_442),
.A2(n_420),
.B(n_458),
.Y(n_495)
);

OA21x2_ASAP7_75t_L g496 ( 
.A1(n_441),
.A2(n_453),
.B(n_449),
.Y(n_496)
);

OAI21x1_ASAP7_75t_L g497 ( 
.A1(n_441),
.A2(n_451),
.B(n_431),
.Y(n_497)
);

OAI21x1_ASAP7_75t_L g498 ( 
.A1(n_451),
.A2(n_418),
.B(n_446),
.Y(n_498)
);

OR2x2_ASAP7_75t_L g499 ( 
.A(n_432),
.B(n_414),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_446),
.Y(n_500)
);

AOI21x1_ASAP7_75t_L g501 ( 
.A1(n_440),
.A2(n_433),
.B(n_444),
.Y(n_501)
);

OAI21x1_ASAP7_75t_L g502 ( 
.A1(n_419),
.A2(n_352),
.B(n_438),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_424),
.Y(n_503)
);

HB1xp67_ASAP7_75t_L g504 ( 
.A(n_414),
.Y(n_504)
);

BUFx2_ASAP7_75t_L g505 ( 
.A(n_431),
.Y(n_505)
);

INVx2_ASAP7_75t_L g506 ( 
.A(n_424),
.Y(n_506)
);

NAND2x1p5_ASAP7_75t_L g507 ( 
.A(n_443),
.B(n_446),
.Y(n_507)
);

OAI21xp5_ASAP7_75t_L g508 ( 
.A1(n_423),
.A2(n_384),
.B(n_392),
.Y(n_508)
);

AO31x2_ASAP7_75t_L g509 ( 
.A1(n_415),
.A2(n_398),
.A3(n_369),
.B(n_372),
.Y(n_509)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_506),
.Y(n_510)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_506),
.Y(n_511)
);

INVx2_ASAP7_75t_SL g512 ( 
.A(n_491),
.Y(n_512)
);

BUFx6f_ASAP7_75t_L g513 ( 
.A(n_478),
.Y(n_513)
);

INVx2_ASAP7_75t_L g514 ( 
.A(n_469),
.Y(n_514)
);

BUFx3_ASAP7_75t_L g515 ( 
.A(n_491),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_475),
.B(n_479),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_508),
.B(n_486),
.Y(n_517)
);

AND2x2_ASAP7_75t_L g518 ( 
.A(n_503),
.B(n_505),
.Y(n_518)
);

AND2x4_ASAP7_75t_L g519 ( 
.A(n_473),
.B(n_498),
.Y(n_519)
);

INVx2_ASAP7_75t_L g520 ( 
.A(n_502),
.Y(n_520)
);

OR2x2_ASAP7_75t_L g521 ( 
.A(n_484),
.B(n_505),
.Y(n_521)
);

AOI22xp33_ASAP7_75t_L g522 ( 
.A1(n_496),
.A2(n_471),
.B1(n_494),
.B2(n_483),
.Y(n_522)
);

BUFx2_ASAP7_75t_L g523 ( 
.A(n_474),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_470),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_SL g525 ( 
.A(n_499),
.B(n_473),
.Y(n_525)
);

INVx3_ASAP7_75t_L g526 ( 
.A(n_473),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_476),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_477),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_485),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_498),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_509),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_509),
.Y(n_532)
);

HB1xp67_ASAP7_75t_L g533 ( 
.A(n_504),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_509),
.Y(n_534)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_480),
.Y(n_535)
);

AOI22xp33_ASAP7_75t_L g536 ( 
.A1(n_496),
.A2(n_471),
.B1(n_467),
.B2(n_465),
.Y(n_536)
);

AND2x2_ASAP7_75t_L g537 ( 
.A(n_496),
.B(n_509),
.Y(n_537)
);

BUFx12f_ASAP7_75t_L g538 ( 
.A(n_499),
.Y(n_538)
);

HB1xp67_ASAP7_75t_L g539 ( 
.A(n_478),
.Y(n_539)
);

AOI22xp33_ASAP7_75t_L g540 ( 
.A1(n_471),
.A2(n_467),
.B1(n_497),
.B2(n_481),
.Y(n_540)
);

INVx2_ASAP7_75t_L g541 ( 
.A(n_467),
.Y(n_541)
);

INVx2_ASAP7_75t_L g542 ( 
.A(n_466),
.Y(n_542)
);

AND2x2_ASAP7_75t_L g543 ( 
.A(n_497),
.B(n_490),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_500),
.Y(n_544)
);

INVx3_ASAP7_75t_L g545 ( 
.A(n_478),
.Y(n_545)
);

INVx2_ASAP7_75t_L g546 ( 
.A(n_495),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_490),
.Y(n_547)
);

INVx4_ASAP7_75t_L g548 ( 
.A(n_478),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_L g549 ( 
.A(n_490),
.B(n_489),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_481),
.Y(n_550)
);

INVx2_ASAP7_75t_SL g551 ( 
.A(n_515),
.Y(n_551)
);

AND2x2_ASAP7_75t_L g552 ( 
.A(n_510),
.B(n_507),
.Y(n_552)
);

OR2x2_ASAP7_75t_L g553 ( 
.A(n_516),
.B(n_521),
.Y(n_553)
);

INVx2_ASAP7_75t_L g554 ( 
.A(n_546),
.Y(n_554)
);

OR2x2_ASAP7_75t_L g555 ( 
.A(n_516),
.B(n_495),
.Y(n_555)
);

HB1xp67_ASAP7_75t_L g556 ( 
.A(n_523),
.Y(n_556)
);

HB1xp67_ASAP7_75t_L g557 ( 
.A(n_523),
.Y(n_557)
);

INVx2_ASAP7_75t_L g558 ( 
.A(n_510),
.Y(n_558)
);

INVx2_ASAP7_75t_L g559 ( 
.A(n_510),
.Y(n_559)
);

INVx2_ASAP7_75t_L g560 ( 
.A(n_511),
.Y(n_560)
);

BUFx2_ASAP7_75t_L g561 ( 
.A(n_518),
.Y(n_561)
);

HB1xp67_ASAP7_75t_L g562 ( 
.A(n_533),
.Y(n_562)
);

INVx2_ASAP7_75t_SL g563 ( 
.A(n_515),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_L g564 ( 
.A(n_521),
.B(n_507),
.Y(n_564)
);

AND2x2_ASAP7_75t_L g565 ( 
.A(n_511),
.B(n_495),
.Y(n_565)
);

INVx6_ASAP7_75t_L g566 ( 
.A(n_538),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_L g567 ( 
.A(n_518),
.B(n_517),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_L g568 ( 
.A(n_517),
.B(n_493),
.Y(n_568)
);

AND2x2_ASAP7_75t_L g569 ( 
.A(n_511),
.B(n_488),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_530),
.Y(n_570)
);

INVx2_ASAP7_75t_L g571 ( 
.A(n_514),
.Y(n_571)
);

HB1xp67_ASAP7_75t_L g572 ( 
.A(n_515),
.Y(n_572)
);

AND2x2_ASAP7_75t_L g573 ( 
.A(n_514),
.B(n_488),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_530),
.Y(n_574)
);

NOR2xp33_ASAP7_75t_L g575 ( 
.A(n_525),
.B(n_493),
.Y(n_575)
);

AOI22xp33_ASAP7_75t_L g576 ( 
.A1(n_538),
.A2(n_492),
.B1(n_487),
.B2(n_472),
.Y(n_576)
);

HB1xp67_ASAP7_75t_L g577 ( 
.A(n_539),
.Y(n_577)
);

AND2x2_ASAP7_75t_L g578 ( 
.A(n_514),
.B(n_526),
.Y(n_578)
);

INVx2_ASAP7_75t_SL g579 ( 
.A(n_538),
.Y(n_579)
);

HB1xp67_ASAP7_75t_L g580 ( 
.A(n_512),
.Y(n_580)
);

INVx2_ASAP7_75t_L g581 ( 
.A(n_524),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_531),
.Y(n_582)
);

AND2x2_ASAP7_75t_L g583 ( 
.A(n_526),
.B(n_487),
.Y(n_583)
);

AND2x2_ASAP7_75t_L g584 ( 
.A(n_526),
.B(n_472),
.Y(n_584)
);

AND2x4_ASAP7_75t_SL g585 ( 
.A(n_519),
.B(n_526),
.Y(n_585)
);

INVx3_ASAP7_75t_L g586 ( 
.A(n_519),
.Y(n_586)
);

OR2x2_ASAP7_75t_L g587 ( 
.A(n_537),
.B(n_482),
.Y(n_587)
);

INVx3_ASAP7_75t_L g588 ( 
.A(n_519),
.Y(n_588)
);

OAI22xp5_ASAP7_75t_L g589 ( 
.A1(n_522),
.A2(n_501),
.B1(n_482),
.B2(n_468),
.Y(n_589)
);

AND2x2_ASAP7_75t_L g590 ( 
.A(n_519),
.B(n_468),
.Y(n_590)
);

AOI22xp5_ASAP7_75t_L g591 ( 
.A1(n_528),
.A2(n_529),
.B1(n_524),
.B2(n_527),
.Y(n_591)
);

AND2x2_ASAP7_75t_L g592 ( 
.A(n_537),
.B(n_527),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_531),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_532),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_532),
.Y(n_595)
);

OR2x2_ASAP7_75t_L g596 ( 
.A(n_534),
.B(n_541),
.Y(n_596)
);

AND2x2_ASAP7_75t_L g597 ( 
.A(n_528),
.B(n_529),
.Y(n_597)
);

AND2x2_ASAP7_75t_L g598 ( 
.A(n_592),
.B(n_534),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_570),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_570),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_581),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_574),
.Y(n_602)
);

AND2x2_ASAP7_75t_L g603 ( 
.A(n_592),
.B(n_543),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_SL g604 ( 
.A(n_568),
.B(n_575),
.Y(n_604)
);

AND2x2_ASAP7_75t_L g605 ( 
.A(n_586),
.B(n_543),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_574),
.Y(n_606)
);

INVx2_ASAP7_75t_L g607 ( 
.A(n_571),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_567),
.B(n_544),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_582),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_582),
.Y(n_610)
);

INVx2_ASAP7_75t_L g611 ( 
.A(n_571),
.Y(n_611)
);

BUFx2_ASAP7_75t_L g612 ( 
.A(n_586),
.Y(n_612)
);

BUFx2_ASAP7_75t_L g613 ( 
.A(n_586),
.Y(n_613)
);

OR2x2_ASAP7_75t_L g614 ( 
.A(n_555),
.B(n_541),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_593),
.Y(n_615)
);

INVx2_ASAP7_75t_SL g616 ( 
.A(n_566),
.Y(n_616)
);

INVx2_ASAP7_75t_L g617 ( 
.A(n_554),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_581),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_597),
.Y(n_619)
);

AND2x2_ASAP7_75t_L g620 ( 
.A(n_588),
.B(n_561),
.Y(n_620)
);

INVx2_ASAP7_75t_L g621 ( 
.A(n_554),
.Y(n_621)
);

NOR2xp67_ASAP7_75t_L g622 ( 
.A(n_579),
.B(n_512),
.Y(n_622)
);

AND2x2_ASAP7_75t_L g623 ( 
.A(n_588),
.B(n_536),
.Y(n_623)
);

NOR2xp33_ASAP7_75t_L g624 ( 
.A(n_562),
.B(n_544),
.Y(n_624)
);

AOI22xp33_ASAP7_75t_L g625 ( 
.A1(n_566),
.A2(n_550),
.B1(n_549),
.B2(n_540),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_593),
.Y(n_626)
);

OR2x2_ASAP7_75t_L g627 ( 
.A(n_555),
.B(n_550),
.Y(n_627)
);

HB1xp67_ASAP7_75t_L g628 ( 
.A(n_556),
.Y(n_628)
);

INVx2_ASAP7_75t_L g629 ( 
.A(n_554),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_L g630 ( 
.A(n_553),
.B(n_547),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_594),
.Y(n_631)
);

AND2x2_ASAP7_75t_L g632 ( 
.A(n_588),
.B(n_520),
.Y(n_632)
);

AND2x4_ASAP7_75t_L g633 ( 
.A(n_620),
.B(n_590),
.Y(n_633)
);

NAND2x1_ASAP7_75t_L g634 ( 
.A(n_616),
.B(n_566),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_599),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_599),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_600),
.Y(n_637)
);

AND2x2_ASAP7_75t_L g638 ( 
.A(n_603),
.B(n_587),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_L g639 ( 
.A(n_628),
.B(n_608),
.Y(n_639)
);

AND2x2_ASAP7_75t_L g640 ( 
.A(n_603),
.B(n_587),
.Y(n_640)
);

AND2x2_ASAP7_75t_SL g641 ( 
.A(n_612),
.B(n_561),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_L g642 ( 
.A(n_604),
.B(n_553),
.Y(n_642)
);

AND2x2_ASAP7_75t_L g643 ( 
.A(n_620),
.B(n_565),
.Y(n_643)
);

OR2x2_ASAP7_75t_L g644 ( 
.A(n_614),
.B(n_596),
.Y(n_644)
);

INVxp67_ASAP7_75t_L g645 ( 
.A(n_624),
.Y(n_645)
);

AND2x2_ASAP7_75t_L g646 ( 
.A(n_605),
.B(n_565),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_L g647 ( 
.A(n_630),
.B(n_557),
.Y(n_647)
);

INVx1_ASAP7_75t_SL g648 ( 
.A(n_612),
.Y(n_648)
);

AND2x4_ASAP7_75t_L g649 ( 
.A(n_613),
.B(n_590),
.Y(n_649)
);

NOR2xp33_ASAP7_75t_L g650 ( 
.A(n_623),
.B(n_564),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_600),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_602),
.Y(n_652)
);

AND2x2_ASAP7_75t_L g653 ( 
.A(n_605),
.B(n_573),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_L g654 ( 
.A(n_619),
.B(n_578),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_602),
.Y(n_655)
);

OR2x2_ASAP7_75t_L g656 ( 
.A(n_614),
.B(n_596),
.Y(n_656)
);

AND2x2_ASAP7_75t_L g657 ( 
.A(n_623),
.B(n_573),
.Y(n_657)
);

AND2x2_ASAP7_75t_L g658 ( 
.A(n_598),
.B(n_595),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_635),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_650),
.B(n_627),
.Y(n_660)
);

INVx2_ASAP7_75t_L g661 ( 
.A(n_636),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_637),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_L g663 ( 
.A(n_650),
.B(n_639),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_651),
.Y(n_664)
);

OAI32xp33_ASAP7_75t_L g665 ( 
.A1(n_642),
.A2(n_580),
.A3(n_627),
.B1(n_626),
.B2(n_615),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_652),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_655),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_SL g668 ( 
.A(n_641),
.B(n_616),
.Y(n_668)
);

AND2x2_ASAP7_75t_L g669 ( 
.A(n_657),
.B(n_613),
.Y(n_669)
);

AOI21xp5_ASAP7_75t_L g670 ( 
.A1(n_641),
.A2(n_589),
.B(n_576),
.Y(n_670)
);

OR2x2_ASAP7_75t_L g671 ( 
.A(n_657),
.B(n_610),
.Y(n_671)
);

AND2x2_ASAP7_75t_L g672 ( 
.A(n_653),
.B(n_598),
.Y(n_672)
);

AND2x2_ASAP7_75t_L g673 ( 
.A(n_672),
.B(n_638),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_661),
.Y(n_674)
);

A2O1A1Ixp33_ASAP7_75t_L g675 ( 
.A1(n_670),
.A2(n_645),
.B(n_579),
.C(n_634),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_663),
.B(n_647),
.Y(n_676)
);

NAND4xp75_ASAP7_75t_L g677 ( 
.A(n_668),
.B(n_622),
.C(n_563),
.D(n_551),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_661),
.Y(n_678)
);

AOI322xp5_ASAP7_75t_L g679 ( 
.A1(n_668),
.A2(n_638),
.A3(n_640),
.B1(n_658),
.B2(n_653),
.C1(n_646),
.C2(n_643),
.Y(n_679)
);

OAI21xp5_ASAP7_75t_L g680 ( 
.A1(n_665),
.A2(n_625),
.B(n_591),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_L g681 ( 
.A(n_660),
.B(n_640),
.Y(n_681)
);

AOI22xp5_ASAP7_75t_L g682 ( 
.A1(n_669),
.A2(n_566),
.B1(n_633),
.B2(n_649),
.Y(n_682)
);

OR2x2_ASAP7_75t_L g683 ( 
.A(n_669),
.B(n_656),
.Y(n_683)
);

AO21x1_ASAP7_75t_L g684 ( 
.A1(n_680),
.A2(n_676),
.B(n_674),
.Y(n_684)
);

AOI22xp5_ASAP7_75t_L g685 ( 
.A1(n_680),
.A2(n_633),
.B1(n_649),
.B2(n_585),
.Y(n_685)
);

AOI21xp5_ASAP7_75t_L g686 ( 
.A1(n_675),
.A2(n_549),
.B(n_654),
.Y(n_686)
);

INVxp67_ASAP7_75t_L g687 ( 
.A(n_681),
.Y(n_687)
);

AOI21xp5_ASAP7_75t_L g688 ( 
.A1(n_678),
.A2(n_659),
.B(n_667),
.Y(n_688)
);

AND2x2_ASAP7_75t_L g689 ( 
.A(n_687),
.B(n_673),
.Y(n_689)
);

OAI22x1_ASAP7_75t_L g690 ( 
.A1(n_685),
.A2(n_682),
.B1(n_683),
.B2(n_664),
.Y(n_690)
);

OAI221xp5_ASAP7_75t_L g691 ( 
.A1(n_688),
.A2(n_679),
.B1(n_662),
.B2(n_666),
.C(n_671),
.Y(n_691)
);

CKINVDCx5p33_ASAP7_75t_R g692 ( 
.A(n_686),
.Y(n_692)
);

NOR2xp33_ASAP7_75t_L g693 ( 
.A(n_684),
.B(n_677),
.Y(n_693)
);

O2A1O1Ixp33_ASAP7_75t_L g694 ( 
.A1(n_684),
.A2(n_577),
.B(n_572),
.C(n_648),
.Y(n_694)
);

NOR4xp25_ASAP7_75t_L g695 ( 
.A(n_694),
.B(n_597),
.C(n_563),
.D(n_551),
.Y(n_695)
);

AOI21xp5_ASAP7_75t_L g696 ( 
.A1(n_692),
.A2(n_672),
.B(n_649),
.Y(n_696)
);

NOR2xp33_ASAP7_75t_L g697 ( 
.A(n_691),
.B(n_633),
.Y(n_697)
);

HB1xp67_ASAP7_75t_L g698 ( 
.A(n_693),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_689),
.Y(n_699)
);

NOR3xp33_ASAP7_75t_L g700 ( 
.A(n_698),
.B(n_690),
.C(n_548),
.Y(n_700)
);

AOI22xp5_ASAP7_75t_L g701 ( 
.A1(n_697),
.A2(n_658),
.B1(n_646),
.B2(n_643),
.Y(n_701)
);

NAND4xp75_ASAP7_75t_L g702 ( 
.A(n_696),
.B(n_591),
.C(n_552),
.D(n_618),
.Y(n_702)
);

AOI21xp33_ASAP7_75t_SL g703 ( 
.A1(n_700),
.A2(n_695),
.B(n_699),
.Y(n_703)
);

AO22x1_ASAP7_75t_L g704 ( 
.A1(n_702),
.A2(n_535),
.B1(n_601),
.B2(n_606),
.Y(n_704)
);

NAND3xp33_ASAP7_75t_L g705 ( 
.A(n_701),
.B(n_535),
.C(n_552),
.Y(n_705)
);

OAI22xp5_ASAP7_75t_L g706 ( 
.A1(n_703),
.A2(n_644),
.B1(n_631),
.B2(n_626),
.Y(n_706)
);

NOR2x1_ASAP7_75t_L g707 ( 
.A(n_705),
.B(n_548),
.Y(n_707)
);

XOR2xp5_ASAP7_75t_L g708 ( 
.A(n_704),
.B(n_547),
.Y(n_708)
);

NAND4xp75_ASAP7_75t_L g709 ( 
.A(n_703),
.B(n_578),
.C(n_606),
.D(n_615),
.Y(n_709)
);

AND2x4_ASAP7_75t_L g710 ( 
.A(n_705),
.B(n_585),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_705),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_711),
.Y(n_712)
);

INVx4_ASAP7_75t_L g713 ( 
.A(n_710),
.Y(n_713)
);

OA22x2_ASAP7_75t_L g714 ( 
.A1(n_706),
.A2(n_631),
.B1(n_609),
.B2(n_610),
.Y(n_714)
);

AND3x4_ASAP7_75t_L g715 ( 
.A(n_707),
.B(n_535),
.C(n_611),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_708),
.Y(n_716)
);

XNOR2x1_ASAP7_75t_L g717 ( 
.A(n_709),
.B(n_545),
.Y(n_717)
);

BUFx2_ASAP7_75t_L g718 ( 
.A(n_707),
.Y(n_718)
);

OA22x2_ASAP7_75t_L g719 ( 
.A1(n_713),
.A2(n_609),
.B1(n_585),
.B2(n_548),
.Y(n_719)
);

AO21x2_ASAP7_75t_L g720 ( 
.A1(n_712),
.A2(n_595),
.B(n_594),
.Y(n_720)
);

OAI21xp5_ASAP7_75t_SL g721 ( 
.A1(n_716),
.A2(n_583),
.B(n_584),
.Y(n_721)
);

OAI22xp5_ASAP7_75t_L g722 ( 
.A1(n_715),
.A2(n_545),
.B1(n_548),
.B2(n_607),
.Y(n_722)
);

CKINVDCx14_ASAP7_75t_R g723 ( 
.A(n_718),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_L g724 ( 
.A(n_717),
.B(n_545),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_723),
.Y(n_725)
);

OA22x2_ASAP7_75t_L g726 ( 
.A1(n_721),
.A2(n_714),
.B1(n_545),
.B2(n_607),
.Y(n_726)
);

AO22x1_ASAP7_75t_L g727 ( 
.A1(n_724),
.A2(n_513),
.B1(n_611),
.B2(n_559),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_720),
.Y(n_728)
);

OAI21xp5_ASAP7_75t_L g729 ( 
.A1(n_722),
.A2(n_583),
.B(n_584),
.Y(n_729)
);

OAI22xp5_ASAP7_75t_SL g730 ( 
.A1(n_719),
.A2(n_513),
.B1(n_560),
.B2(n_559),
.Y(n_730)
);

OAI221xp5_ASAP7_75t_L g731 ( 
.A1(n_725),
.A2(n_513),
.B1(n_560),
.B2(n_558),
.C(n_542),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_728),
.Y(n_732)
);

OAI22xp5_ASAP7_75t_SL g733 ( 
.A1(n_730),
.A2(n_513),
.B1(n_558),
.B2(n_617),
.Y(n_733)
);

AOI221x1_ASAP7_75t_L g734 ( 
.A1(n_729),
.A2(n_513),
.B1(n_617),
.B2(n_621),
.C(n_629),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_726),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_732),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_735),
.Y(n_737)
);

OAI21xp33_ASAP7_75t_L g738 ( 
.A1(n_737),
.A2(n_731),
.B(n_733),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_736),
.B(n_727),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_L g740 ( 
.A(n_738),
.B(n_734),
.Y(n_740)
);

OR2x6_ASAP7_75t_L g741 ( 
.A(n_740),
.B(n_739),
.Y(n_741)
);

AOI211xp5_ASAP7_75t_L g742 ( 
.A1(n_741),
.A2(n_513),
.B(n_569),
.C(n_632),
.Y(n_742)
);


endmodule