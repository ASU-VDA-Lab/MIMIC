module fake_jpeg_18413_n_323 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_323);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_323;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_13;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_145;
wire n_18;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_12;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx12f_ASAP7_75t_L g12 ( 
.A(n_8),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_1),
.Y(n_13)
);

BUFx12_ASAP7_75t_L g14 ( 
.A(n_3),
.Y(n_14)
);

BUFx12f_ASAP7_75t_L g15 ( 
.A(n_9),
.Y(n_15)
);

BUFx5_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_9),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_0),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_9),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

INVx8_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_27),
.B(n_28),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g28 ( 
.A(n_20),
.B(n_11),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_23),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_SL g41 ( 
.A(n_29),
.B(n_30),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_23),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_17),
.B(n_11),
.Y(n_31)
);

CKINVDCx14_ASAP7_75t_R g45 ( 
.A(n_31),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_32),
.Y(n_38)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_33),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_34),
.Y(n_39)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_12),
.Y(n_35)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

INVx11_ASAP7_75t_L g42 ( 
.A(n_26),
.Y(n_42)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_SL g43 ( 
.A1(n_26),
.A2(n_24),
.B1(n_25),
.B2(n_20),
.Y(n_43)
);

INVx1_ASAP7_75t_SL g59 ( 
.A(n_43),
.Y(n_59)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_26),
.Y(n_46)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_46),
.Y(n_60)
);

OAI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_33),
.A2(n_24),
.B1(n_25),
.B2(n_13),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_47),
.A2(n_26),
.B1(n_35),
.B2(n_33),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_41),
.B(n_30),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_48),
.B(n_49),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_41),
.B(n_28),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_45),
.B(n_29),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_50),
.B(n_52),
.Y(n_73)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_51),
.Y(n_80)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_44),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_41),
.B(n_30),
.Y(n_53)
);

XNOR2xp5_ASAP7_75t_L g67 ( 
.A(n_53),
.B(n_61),
.Y(n_67)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_55),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_L g56 ( 
.A1(n_45),
.A2(n_37),
.B1(n_28),
.B2(n_30),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_56),
.A2(n_63),
.B1(n_64),
.B2(n_66),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_57),
.Y(n_72)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_58),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_37),
.B(n_29),
.Y(n_61)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_40),
.Y(n_62)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_62),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_45),
.B(n_31),
.Y(n_64)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_44),
.Y(n_65)
);

INVxp67_ASAP7_75t_L g69 ( 
.A(n_65),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_37),
.B(n_29),
.Y(n_66)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_55),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_68),
.Y(n_93)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_60),
.Y(n_74)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_74),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_55),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_76),
.B(n_79),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_59),
.A2(n_43),
.B1(n_47),
.B2(n_33),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_77),
.A2(n_47),
.B1(n_35),
.B2(n_27),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_55),
.Y(n_79)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_60),
.Y(n_81)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_81),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_50),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_83),
.B(n_87),
.Y(n_100)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_57),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_84),
.Y(n_94)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_57),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_85),
.B(n_62),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_L g86 ( 
.A1(n_61),
.A2(n_43),
.B(n_31),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_SL g101 ( 
.A1(n_86),
.A2(n_17),
.B(n_21),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_48),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_86),
.A2(n_59),
.B1(n_66),
.B2(n_63),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_88),
.A2(n_91),
.B1(n_109),
.B2(n_27),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_75),
.B(n_53),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_89),
.B(n_90),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_75),
.B(n_67),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_77),
.A2(n_59),
.B1(n_43),
.B2(n_49),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_95),
.A2(n_103),
.B1(n_36),
.B2(n_46),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_83),
.A2(n_64),
.B1(n_24),
.B2(n_35),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_96),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_73),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_99),
.B(n_102),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_L g139 ( 
.A(n_101),
.B(n_14),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_67),
.B(n_40),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_78),
.A2(n_44),
.B1(n_36),
.B2(n_46),
.Y(n_103)
);

INVx13_ASAP7_75t_L g104 ( 
.A(n_70),
.Y(n_104)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_104),
.Y(n_114)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_74),
.Y(n_105)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_105),
.Y(n_117)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_106),
.Y(n_131)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_71),
.Y(n_107)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_107),
.Y(n_123)
);

BUFx2_ASAP7_75t_L g108 ( 
.A(n_80),
.Y(n_108)
);

CKINVDCx14_ASAP7_75t_R g118 ( 
.A(n_108),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_87),
.A2(n_44),
.B1(n_51),
.B2(n_58),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_100),
.B(n_21),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_110),
.B(n_119),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_112),
.A2(n_121),
.B1(n_126),
.B2(n_128),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_107),
.A2(n_68),
.B1(n_54),
.B2(n_84),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_113),
.A2(n_116),
.B1(n_94),
.B2(n_39),
.Y(n_162)
);

AOI21xp33_ASAP7_75t_L g115 ( 
.A1(n_100),
.A2(n_81),
.B(n_76),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_SL g143 ( 
.A1(n_115),
.A2(n_14),
.B(n_19),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_97),
.A2(n_54),
.B1(n_85),
.B2(n_60),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_97),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_L g120 ( 
.A1(n_96),
.A2(n_69),
.B(n_79),
.Y(n_120)
);

AOI21xp5_ASAP7_75t_L g156 ( 
.A1(n_120),
.A2(n_129),
.B(n_80),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_95),
.A2(n_103),
.B1(n_91),
.B2(n_88),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_90),
.B(n_27),
.C(n_65),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_122),
.B(n_127),
.C(n_112),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_124),
.A2(n_130),
.B1(n_138),
.B2(n_38),
.Y(n_154)
);

MAJx2_ASAP7_75t_L g125 ( 
.A(n_101),
.B(n_69),
.C(n_14),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_125),
.B(n_19),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_89),
.A2(n_72),
.B1(n_65),
.B2(n_46),
.Y(n_126)
);

OA21x2_ASAP7_75t_L g127 ( 
.A1(n_92),
.A2(n_72),
.B(n_52),
.Y(n_127)
);

AO22x1_ASAP7_75t_L g158 ( 
.A1(n_127),
.A2(n_39),
.B1(n_94),
.B2(n_32),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_102),
.A2(n_36),
.B1(n_25),
.B2(n_42),
.Y(n_128)
);

OAI31xp33_ASAP7_75t_L g129 ( 
.A1(n_98),
.A2(n_42),
.A3(n_14),
.B(n_36),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_109),
.A2(n_42),
.B1(n_52),
.B2(n_71),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g132 ( 
.A(n_92),
.B(n_54),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_132),
.B(n_134),
.Y(n_152)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_98),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_105),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_135),
.B(n_137),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_93),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_108),
.A2(n_82),
.B1(n_34),
.B2(n_32),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_139),
.B(n_15),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_131),
.B(n_104),
.Y(n_140)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_140),
.Y(n_180)
);

OAI22x1_ASAP7_75t_L g141 ( 
.A1(n_120),
.A2(n_108),
.B1(n_104),
.B2(n_93),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_141),
.A2(n_163),
.B1(n_165),
.B2(n_118),
.Y(n_178)
);

INVx13_ASAP7_75t_L g142 ( 
.A(n_114),
.Y(n_142)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_142),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_143),
.B(n_146),
.Y(n_176)
);

AND2x2_ASAP7_75t_L g144 ( 
.A(n_124),
.B(n_93),
.Y(n_144)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_144),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g145 ( 
.A(n_133),
.B(n_82),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_SL g179 ( 
.A(n_145),
.B(n_172),
.Y(n_179)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_123),
.Y(n_146)
);

INVx13_ASAP7_75t_L g147 ( 
.A(n_114),
.Y(n_147)
);

CKINVDCx16_ASAP7_75t_R g183 ( 
.A(n_147),
.Y(n_183)
);

AND2x2_ASAP7_75t_L g150 ( 
.A(n_127),
.B(n_70),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_150),
.B(n_151),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_131),
.B(n_94),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_153),
.B(n_164),
.C(n_136),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_154),
.A2(n_162),
.B1(n_39),
.B2(n_38),
.Y(n_187)
);

INVx1_ASAP7_75t_SL g155 ( 
.A(n_117),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_155),
.B(n_157),
.Y(n_197)
);

CKINVDCx16_ASAP7_75t_R g184 ( 
.A(n_156),
.Y(n_184)
);

AND2x2_ASAP7_75t_SL g157 ( 
.A(n_117),
.B(n_16),
.Y(n_157)
);

OA21x2_ASAP7_75t_L g194 ( 
.A1(n_158),
.A2(n_167),
.B(n_16),
.Y(n_194)
);

INVx13_ASAP7_75t_L g159 ( 
.A(n_137),
.Y(n_159)
);

INVxp33_ASAP7_75t_SL g190 ( 
.A(n_159),
.Y(n_190)
);

AND2x2_ASAP7_75t_L g160 ( 
.A(n_111),
.B(n_12),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_160),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_111),
.A2(n_38),
.B1(n_34),
.B2(n_32),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_122),
.B(n_34),
.C(n_32),
.Y(n_164)
);

INVxp67_ASAP7_75t_L g165 ( 
.A(n_130),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_165),
.Y(n_198)
);

INVx1_ASAP7_75t_SL g166 ( 
.A(n_134),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_166),
.Y(n_200)
);

OAI21xp33_ASAP7_75t_L g167 ( 
.A1(n_125),
.A2(n_11),
.B(n_10),
.Y(n_167)
);

CKINVDCx16_ASAP7_75t_R g168 ( 
.A(n_135),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_168),
.Y(n_201)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_123),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_169),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_170),
.B(n_173),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_119),
.B(n_14),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_SL g188 ( 
.A(n_171),
.B(n_149),
.Y(n_188)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_136),
.B(n_139),
.Y(n_172)
);

AND2x2_ASAP7_75t_L g173 ( 
.A(n_129),
.B(n_15),
.Y(n_173)
);

MAJx2_ASAP7_75t_L g196 ( 
.A(n_174),
.B(n_19),
.C(n_15),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_175),
.B(n_196),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_178),
.A2(n_154),
.B1(n_150),
.B2(n_173),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_172),
.B(n_138),
.C(n_34),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_181),
.B(n_189),
.C(n_202),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_187),
.A2(n_193),
.B1(n_202),
.B2(n_181),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_188),
.B(n_157),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_145),
.B(n_153),
.C(n_174),
.Y(n_189)
);

AND2x6_ASAP7_75t_L g192 ( 
.A(n_141),
.B(n_16),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_192),
.B(n_194),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_144),
.A2(n_38),
.B1(n_39),
.B2(n_34),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_164),
.B(n_156),
.C(n_152),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_195),
.B(n_142),
.C(n_22),
.Y(n_227)
);

MAJx2_ASAP7_75t_L g199 ( 
.A(n_167),
.B(n_15),
.C(n_22),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_SL g213 ( 
.A(n_199),
.B(n_163),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_144),
.B(n_32),
.C(n_15),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_SL g204 ( 
.A(n_180),
.B(n_155),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_204),
.B(n_212),
.Y(n_235)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_190),
.Y(n_205)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_205),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_200),
.B(n_161),
.Y(n_206)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_206),
.Y(n_236)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_190),
.Y(n_207)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_207),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_182),
.B(n_166),
.Y(n_208)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_208),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_209),
.A2(n_198),
.B1(n_187),
.B2(n_175),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_210),
.A2(n_216),
.B1(n_178),
.B2(n_220),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_185),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_213),
.B(n_191),
.Y(n_237)
);

INVxp33_ASAP7_75t_L g214 ( 
.A(n_197),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_214),
.Y(n_228)
);

A2O1A1Ixp33_ASAP7_75t_L g215 ( 
.A1(n_192),
.A2(n_150),
.B(n_173),
.C(n_160),
.Y(n_215)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_215),
.Y(n_248)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_193),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_216),
.B(n_217),
.Y(n_233)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_176),
.Y(n_218)
);

AOI22xp33_ASAP7_75t_SL g240 ( 
.A1(n_218),
.A2(n_221),
.B1(n_224),
.B2(n_203),
.Y(n_240)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_186),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_L g222 ( 
.A1(n_184),
.A2(n_160),
.B(n_158),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_L g241 ( 
.A1(n_222),
.A2(n_223),
.B(n_199),
.Y(n_241)
);

AOI21xp5_ASAP7_75t_SL g223 ( 
.A1(n_194),
.A2(n_157),
.B(n_148),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_195),
.Y(n_224)
);

OAI21xp33_ASAP7_75t_L g225 ( 
.A1(n_177),
.A2(n_148),
.B(n_159),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_225),
.B(n_222),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_201),
.B(n_147),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_L g245 ( 
.A1(n_226),
.A2(n_5),
.B1(n_10),
.B2(n_2),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_227),
.B(n_179),
.C(n_189),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_229),
.B(n_232),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_230),
.A2(n_213),
.B1(n_219),
.B2(n_221),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g257 ( 
.A(n_234),
.B(n_239),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_237),
.B(n_243),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_211),
.B(n_179),
.C(n_191),
.Y(n_239)
);

CKINVDCx14_ASAP7_75t_R g263 ( 
.A(n_240),
.Y(n_263)
);

AOI21xp5_ASAP7_75t_L g265 ( 
.A1(n_241),
.A2(n_209),
.B(n_206),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_211),
.B(n_183),
.C(n_194),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_242),
.B(n_244),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_220),
.B(n_196),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_227),
.B(n_22),
.Y(n_244)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_245),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_210),
.B(n_18),
.C(n_1),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_SL g249 ( 
.A(n_246),
.B(n_244),
.Y(n_249)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_249),
.Y(n_268)
);

A2O1A1O1Ixp25_ASAP7_75t_L g250 ( 
.A1(n_241),
.A2(n_248),
.B(n_228),
.C(n_229),
.D(n_215),
.Y(n_250)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_250),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_235),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_252),
.B(n_258),
.Y(n_274)
);

BUFx2_ASAP7_75t_L g253 ( 
.A(n_228),
.Y(n_253)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_253),
.Y(n_271)
);

INVxp33_ASAP7_75t_SL g254 ( 
.A(n_231),
.Y(n_254)
);

OR2x2_ASAP7_75t_L g275 ( 
.A(n_254),
.B(n_262),
.Y(n_275)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_233),
.Y(n_256)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_256),
.Y(n_277)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_236),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_260),
.B(n_261),
.Y(n_278)
);

INVx13_ASAP7_75t_L g261 ( 
.A(n_238),
.Y(n_261)
);

BUFx2_ASAP7_75t_L g262 ( 
.A(n_247),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_265),
.B(n_234),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_266),
.B(n_250),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_251),
.A2(n_237),
.B1(n_208),
.B2(n_246),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_267),
.A2(n_271),
.B1(n_279),
.B2(n_269),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_257),
.B(n_232),
.C(n_239),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_270),
.B(n_272),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_255),
.B(n_242),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_SL g273 ( 
.A(n_255),
.B(n_243),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_273),
.B(n_259),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_264),
.B(n_214),
.C(n_223),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_276),
.B(n_279),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_263),
.B(n_259),
.C(n_254),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_SL g304 ( 
.A(n_281),
.B(n_4),
.Y(n_304)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_275),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_283),
.B(n_285),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_284),
.B(n_286),
.Y(n_293)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_275),
.Y(n_285)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_278),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_287),
.B(n_291),
.Y(n_295)
);

OAI21xp5_ASAP7_75t_L g288 ( 
.A1(n_274),
.A2(n_253),
.B(n_262),
.Y(n_288)
);

AOI21xp5_ASAP7_75t_L g296 ( 
.A1(n_288),
.A2(n_290),
.B(n_6),
.Y(n_296)
);

AOI22xp33_ASAP7_75t_SL g289 ( 
.A1(n_277),
.A2(n_261),
.B1(n_18),
.B2(n_2),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_L g298 ( 
.A1(n_289),
.A2(n_288),
.B1(n_7),
.B2(n_3),
.Y(n_298)
);

OAI21xp5_ASAP7_75t_L g290 ( 
.A1(n_268),
.A2(n_18),
.B(n_6),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_278),
.A2(n_273),
.B1(n_6),
.B2(n_3),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_277),
.B(n_5),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_292),
.B(n_0),
.Y(n_300)
);

AND2x2_ASAP7_75t_L g294 ( 
.A(n_284),
.B(n_280),
.Y(n_294)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_294),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_296),
.B(n_300),
.Y(n_310)
);

OAI21xp5_ASAP7_75t_SL g297 ( 
.A1(n_282),
.A2(n_6),
.B(n_8),
.Y(n_297)
);

AOI21xp5_ASAP7_75t_L g308 ( 
.A1(n_297),
.A2(n_304),
.B(n_4),
.Y(n_308)
);

INVxp67_ASAP7_75t_L g305 ( 
.A(n_298),
.Y(n_305)
);

INVxp67_ASAP7_75t_SL g299 ( 
.A(n_289),
.Y(n_299)
);

OR2x2_ASAP7_75t_L g306 ( 
.A(n_299),
.B(n_301),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_281),
.B(n_3),
.Y(n_301)
);

AOI21xp5_ASAP7_75t_L g302 ( 
.A1(n_280),
.A2(n_4),
.B(n_7),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_SL g307 ( 
.A(n_302),
.B(n_4),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_307),
.B(n_308),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_SL g309 ( 
.A(n_303),
.B(n_7),
.Y(n_309)
);

BUFx24_ASAP7_75t_SL g313 ( 
.A(n_309),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_295),
.B(n_7),
.Y(n_312)
);

AND2x2_ASAP7_75t_L g314 ( 
.A(n_312),
.B(n_298),
.Y(n_314)
);

AOI322xp5_ASAP7_75t_L g317 ( 
.A1(n_314),
.A2(n_315),
.A3(n_312),
.B1(n_311),
.B2(n_305),
.C1(n_310),
.C2(n_313),
.Y(n_317)
);

NAND2x1p5_ASAP7_75t_L g315 ( 
.A(n_306),
.B(n_293),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_L g319 ( 
.A(n_317),
.B(n_318),
.Y(n_319)
);

OAI21xp5_ASAP7_75t_SL g318 ( 
.A1(n_316),
.A2(n_8),
.B(n_10),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_319),
.Y(n_320)
);

AOI21xp5_ASAP7_75t_SL g321 ( 
.A1(n_320),
.A2(n_10),
.B(n_0),
.Y(n_321)
);

OAI21xp5_ASAP7_75t_L g322 ( 
.A1(n_321),
.A2(n_0),
.B(n_1),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_322),
.B(n_0),
.Y(n_323)
);


endmodule