module fake_netlist_1_2095_n_694 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_694);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_694;
wire n_117;
wire n_663;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_627;
wire n_532;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_563;
wire n_540;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_533;
wire n_506;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_446;
wire n_342;
wire n_423;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_90;
wire n_357;
wire n_653;
wire n_260;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_684;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_84;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_132;
wire n_99;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
CKINVDCx20_ASAP7_75t_R g79 ( .A(n_35), .Y(n_79) );
INVx1_ASAP7_75t_L g80 ( .A(n_55), .Y(n_80) );
INVx1_ASAP7_75t_L g81 ( .A(n_69), .Y(n_81) );
INVx2_ASAP7_75t_L g82 ( .A(n_57), .Y(n_82) );
NOR2xp33_ASAP7_75t_L g83 ( .A(n_38), .B(n_74), .Y(n_83) );
NOR2xp67_ASAP7_75t_L g84 ( .A(n_19), .B(n_59), .Y(n_84) );
INVxp67_ASAP7_75t_L g85 ( .A(n_50), .Y(n_85) );
HB1xp67_ASAP7_75t_L g86 ( .A(n_77), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_63), .Y(n_87) );
INVx1_ASAP7_75t_SL g88 ( .A(n_1), .Y(n_88) );
NOR2xp67_ASAP7_75t_L g89 ( .A(n_24), .B(n_42), .Y(n_89) );
CKINVDCx20_ASAP7_75t_R g90 ( .A(n_22), .Y(n_90) );
INVx2_ASAP7_75t_L g91 ( .A(n_32), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_41), .Y(n_92) );
CKINVDCx5p33_ASAP7_75t_R g93 ( .A(n_28), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_7), .Y(n_94) );
BUFx2_ASAP7_75t_L g95 ( .A(n_52), .Y(n_95) );
INVx2_ASAP7_75t_L g96 ( .A(n_47), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_49), .Y(n_97) );
CKINVDCx20_ASAP7_75t_R g98 ( .A(n_51), .Y(n_98) );
CKINVDCx5p33_ASAP7_75t_R g99 ( .A(n_56), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_3), .Y(n_100) );
CKINVDCx5p33_ASAP7_75t_R g101 ( .A(n_26), .Y(n_101) );
CKINVDCx20_ASAP7_75t_R g102 ( .A(n_11), .Y(n_102) );
INVxp67_ASAP7_75t_L g103 ( .A(n_16), .Y(n_103) );
CKINVDCx16_ASAP7_75t_R g104 ( .A(n_67), .Y(n_104) );
CKINVDCx5p33_ASAP7_75t_R g105 ( .A(n_29), .Y(n_105) );
HB1xp67_ASAP7_75t_L g106 ( .A(n_31), .Y(n_106) );
CKINVDCx5p33_ASAP7_75t_R g107 ( .A(n_46), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_53), .Y(n_108) );
CKINVDCx20_ASAP7_75t_R g109 ( .A(n_37), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_4), .Y(n_110) );
CKINVDCx20_ASAP7_75t_R g111 ( .A(n_54), .Y(n_111) );
INVx2_ASAP7_75t_L g112 ( .A(n_62), .Y(n_112) );
CKINVDCx5p33_ASAP7_75t_R g113 ( .A(n_19), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_34), .Y(n_114) );
INVx1_ASAP7_75t_SL g115 ( .A(n_3), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_1), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_48), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_72), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_12), .Y(n_119) );
INVxp67_ASAP7_75t_SL g120 ( .A(n_45), .Y(n_120) );
CKINVDCx5p33_ASAP7_75t_R g121 ( .A(n_40), .Y(n_121) );
CKINVDCx5p33_ASAP7_75t_R g122 ( .A(n_64), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_11), .Y(n_123) );
CKINVDCx5p33_ASAP7_75t_R g124 ( .A(n_60), .Y(n_124) );
CKINVDCx5p33_ASAP7_75t_R g125 ( .A(n_70), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_9), .Y(n_126) );
INVx1_ASAP7_75t_L g127 ( .A(n_80), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_80), .Y(n_128) );
INVx2_ASAP7_75t_L g129 ( .A(n_82), .Y(n_129) );
INVx2_ASAP7_75t_L g130 ( .A(n_82), .Y(n_130) );
NOR2x1_ASAP7_75t_L g131 ( .A(n_95), .B(n_23), .Y(n_131) );
INVx1_ASAP7_75t_L g132 ( .A(n_81), .Y(n_132) );
NAND2xp5_ASAP7_75t_L g133 ( .A(n_95), .B(n_0), .Y(n_133) );
AND2x4_ASAP7_75t_SL g134 ( .A(n_86), .B(n_25), .Y(n_134) );
INVx2_ASAP7_75t_L g135 ( .A(n_91), .Y(n_135) );
HB1xp67_ASAP7_75t_L g136 ( .A(n_103), .Y(n_136) );
BUFx8_ASAP7_75t_L g137 ( .A(n_81), .Y(n_137) );
BUFx6f_ASAP7_75t_L g138 ( .A(n_91), .Y(n_138) );
NAND2xp5_ASAP7_75t_L g139 ( .A(n_106), .B(n_0), .Y(n_139) );
NAND2xp33_ASAP7_75t_L g140 ( .A(n_93), .B(n_27), .Y(n_140) );
OAI22xp5_ASAP7_75t_SL g141 ( .A1(n_102), .A2(n_2), .B1(n_4), .B2(n_5), .Y(n_141) );
BUFx6f_ASAP7_75t_L g142 ( .A(n_96), .Y(n_142) );
BUFx6f_ASAP7_75t_L g143 ( .A(n_96), .Y(n_143) );
HB1xp67_ASAP7_75t_L g144 ( .A(n_113), .Y(n_144) );
INVx1_ASAP7_75t_L g145 ( .A(n_87), .Y(n_145) );
INVx2_ASAP7_75t_L g146 ( .A(n_112), .Y(n_146) );
INVx1_ASAP7_75t_L g147 ( .A(n_87), .Y(n_147) );
BUFx2_ASAP7_75t_L g148 ( .A(n_104), .Y(n_148) );
BUFx6f_ASAP7_75t_L g149 ( .A(n_112), .Y(n_149) );
BUFx6f_ASAP7_75t_L g150 ( .A(n_92), .Y(n_150) );
INVx1_ASAP7_75t_L g151 ( .A(n_92), .Y(n_151) );
INVx1_ASAP7_75t_L g152 ( .A(n_97), .Y(n_152) );
AND2x6_ASAP7_75t_L g153 ( .A(n_97), .B(n_30), .Y(n_153) );
INVx6_ASAP7_75t_L g154 ( .A(n_104), .Y(n_154) );
OAI22x1_ASAP7_75t_SL g155 ( .A1(n_94), .A2(n_2), .B1(n_5), .B2(n_6), .Y(n_155) );
AND2x2_ASAP7_75t_SL g156 ( .A(n_108), .B(n_78), .Y(n_156) );
INVx1_ASAP7_75t_L g157 ( .A(n_108), .Y(n_157) );
BUFx6f_ASAP7_75t_L g158 ( .A(n_114), .Y(n_158) );
AND2x2_ASAP7_75t_L g159 ( .A(n_94), .B(n_6), .Y(n_159) );
AND2x6_ASAP7_75t_L g160 ( .A(n_114), .B(n_33), .Y(n_160) );
INVx1_ASAP7_75t_L g161 ( .A(n_117), .Y(n_161) );
INVx2_ASAP7_75t_L g162 ( .A(n_117), .Y(n_162) );
INVx2_ASAP7_75t_L g163 ( .A(n_118), .Y(n_163) );
INVx1_ASAP7_75t_L g164 ( .A(n_118), .Y(n_164) );
NOR2x1_ASAP7_75t_L g165 ( .A(n_100), .B(n_36), .Y(n_165) );
INVx1_ASAP7_75t_L g166 ( .A(n_100), .Y(n_166) );
AND2x2_ASAP7_75t_SL g167 ( .A(n_83), .B(n_76), .Y(n_167) );
INVx1_ASAP7_75t_L g168 ( .A(n_110), .Y(n_168) );
AND2x2_ASAP7_75t_SL g169 ( .A(n_110), .B(n_75), .Y(n_169) );
INVx1_ASAP7_75t_L g170 ( .A(n_166), .Y(n_170) );
AOI22xp5_ASAP7_75t_L g171 ( .A1(n_154), .A2(n_126), .B1(n_123), .B2(n_119), .Y(n_171) );
BUFx10_ASAP7_75t_L g172 ( .A(n_154), .Y(n_172) );
CKINVDCx5p33_ASAP7_75t_R g173 ( .A(n_148), .Y(n_173) );
INVx1_ASAP7_75t_L g174 ( .A(n_166), .Y(n_174) );
NAND2xp5_ASAP7_75t_SL g175 ( .A(n_127), .B(n_85), .Y(n_175) );
INVx2_ASAP7_75t_L g176 ( .A(n_138), .Y(n_176) );
INVx1_ASAP7_75t_L g177 ( .A(n_168), .Y(n_177) );
NAND3xp33_ASAP7_75t_SL g178 ( .A(n_148), .B(n_88), .C(n_115), .Y(n_178) );
INVx4_ASAP7_75t_SL g179 ( .A(n_153), .Y(n_179) );
INVx1_ASAP7_75t_L g180 ( .A(n_168), .Y(n_180) );
AND2x6_ASAP7_75t_L g181 ( .A(n_131), .B(n_126), .Y(n_181) );
CKINVDCx5p33_ASAP7_75t_R g182 ( .A(n_154), .Y(n_182) );
NAND2xp5_ASAP7_75t_SL g183 ( .A(n_127), .B(n_89), .Y(n_183) );
HB1xp67_ASAP7_75t_L g184 ( .A(n_144), .Y(n_184) );
AOI22xp5_ASAP7_75t_L g185 ( .A1(n_154), .A2(n_156), .B1(n_169), .B2(n_136), .Y(n_185) );
AND2x2_ASAP7_75t_SL g186 ( .A(n_156), .B(n_116), .Y(n_186) );
BUFx3_ASAP7_75t_L g187 ( .A(n_153), .Y(n_187) );
INVx4_ASAP7_75t_L g188 ( .A(n_153), .Y(n_188) );
NOR2xp33_ASAP7_75t_L g189 ( .A(n_128), .B(n_120), .Y(n_189) );
XOR2x2_ASAP7_75t_L g190 ( .A(n_141), .B(n_84), .Y(n_190) );
BUFx3_ASAP7_75t_L g191 ( .A(n_153), .Y(n_191) );
NAND3xp33_ASAP7_75t_L g192 ( .A(n_133), .B(n_116), .C(n_119), .Y(n_192) );
BUFx3_ASAP7_75t_L g193 ( .A(n_153), .Y(n_193) );
INVx5_ASAP7_75t_L g194 ( .A(n_153), .Y(n_194) );
INVx2_ASAP7_75t_L g195 ( .A(n_138), .Y(n_195) );
BUFx10_ASAP7_75t_L g196 ( .A(n_134), .Y(n_196) );
INVx3_ASAP7_75t_L g197 ( .A(n_150), .Y(n_197) );
OR2x6_ASAP7_75t_L g198 ( .A(n_139), .B(n_123), .Y(n_198) );
OAI22xp33_ASAP7_75t_L g199 ( .A1(n_128), .A2(n_79), .B1(n_90), .B2(n_98), .Y(n_199) );
AND2x6_ASAP7_75t_L g200 ( .A(n_159), .B(n_84), .Y(n_200) );
NAND2xp5_ASAP7_75t_SL g201 ( .A(n_132), .B(n_125), .Y(n_201) );
INVx1_ASAP7_75t_SL g202 ( .A(n_134), .Y(n_202) );
NOR2xp33_ASAP7_75t_L g203 ( .A(n_132), .B(n_124), .Y(n_203) );
INVx1_ASAP7_75t_L g204 ( .A(n_159), .Y(n_204) );
AND2x2_ASAP7_75t_L g205 ( .A(n_145), .B(n_107), .Y(n_205) );
NOR2xp33_ASAP7_75t_L g206 ( .A(n_145), .B(n_122), .Y(n_206) );
INVx1_ASAP7_75t_L g207 ( .A(n_162), .Y(n_207) );
BUFx3_ASAP7_75t_L g208 ( .A(n_153), .Y(n_208) );
INVx2_ASAP7_75t_L g209 ( .A(n_138), .Y(n_209) );
NAND2xp5_ASAP7_75t_SL g210 ( .A(n_147), .B(n_121), .Y(n_210) );
AND2x2_ASAP7_75t_SL g211 ( .A(n_156), .B(n_111), .Y(n_211) );
NAND2xp5_ASAP7_75t_SL g212 ( .A(n_147), .B(n_105), .Y(n_212) );
NAND2xp5_ASAP7_75t_L g213 ( .A(n_151), .B(n_101), .Y(n_213) );
INVx4_ASAP7_75t_L g214 ( .A(n_160), .Y(n_214) );
INVx1_ASAP7_75t_L g215 ( .A(n_162), .Y(n_215) );
NAND2xp5_ASAP7_75t_SL g216 ( .A(n_151), .B(n_99), .Y(n_216) );
INVx2_ASAP7_75t_L g217 ( .A(n_138), .Y(n_217) );
INVxp67_ASAP7_75t_SL g218 ( .A(n_152), .Y(n_218) );
AND2x2_ASAP7_75t_L g219 ( .A(n_152), .B(n_109), .Y(n_219) );
INVx2_ASAP7_75t_L g220 ( .A(n_138), .Y(n_220) );
OR2x6_ASAP7_75t_L g221 ( .A(n_155), .B(n_7), .Y(n_221) );
INVx1_ASAP7_75t_L g222 ( .A(n_163), .Y(n_222) );
NAND2xp5_ASAP7_75t_L g223 ( .A(n_157), .B(n_8), .Y(n_223) );
INVx1_ASAP7_75t_L g224 ( .A(n_163), .Y(n_224) );
INVx4_ASAP7_75t_L g225 ( .A(n_160), .Y(n_225) );
INVx2_ASAP7_75t_L g226 ( .A(n_142), .Y(n_226) );
OR2x2_ASAP7_75t_L g227 ( .A(n_157), .B(n_8), .Y(n_227) );
NOR2xp33_ASAP7_75t_L g228 ( .A(n_161), .B(n_61), .Y(n_228) );
INVx1_ASAP7_75t_L g229 ( .A(n_161), .Y(n_229) );
INVxp33_ASAP7_75t_L g230 ( .A(n_164), .Y(n_230) );
NAND2xp5_ASAP7_75t_SL g231 ( .A(n_164), .B(n_73), .Y(n_231) );
CKINVDCx5p33_ASAP7_75t_R g232 ( .A(n_173), .Y(n_232) );
NAND2xp5_ASAP7_75t_SL g233 ( .A(n_188), .B(n_169), .Y(n_233) );
OAI22xp5_ASAP7_75t_SL g234 ( .A1(n_221), .A2(n_169), .B1(n_155), .B2(n_167), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g235 ( .A(n_230), .B(n_137), .Y(n_235) );
NAND2xp33_ASAP7_75t_L g236 ( .A(n_194), .B(n_160), .Y(n_236) );
AOI22xp33_ASAP7_75t_L g237 ( .A1(n_186), .A2(n_160), .B1(n_167), .B2(n_150), .Y(n_237) );
AOI21xp5_ASAP7_75t_L g238 ( .A1(n_188), .A2(n_140), .B(n_167), .Y(n_238) );
OR2x6_ASAP7_75t_L g239 ( .A(n_221), .B(n_165), .Y(n_239) );
NAND2xp5_ASAP7_75t_L g240 ( .A(n_230), .B(n_137), .Y(n_240) );
AND2x2_ASAP7_75t_L g241 ( .A(n_184), .B(n_129), .Y(n_241) );
OAI22xp5_ASAP7_75t_L g242 ( .A1(n_185), .A2(n_129), .B1(n_130), .B2(n_146), .Y(n_242) );
NAND2xp5_ASAP7_75t_L g243 ( .A(n_218), .B(n_137), .Y(n_243) );
NAND2xp5_ASAP7_75t_SL g244 ( .A(n_214), .B(n_158), .Y(n_244) );
INVx2_ASAP7_75t_SL g245 ( .A(n_172), .Y(n_245) );
INVx1_ASAP7_75t_L g246 ( .A(n_227), .Y(n_246) );
AOI22xp33_ASAP7_75t_L g247 ( .A1(n_186), .A2(n_160), .B1(n_158), .B2(n_150), .Y(n_247) );
INVx2_ASAP7_75t_L g248 ( .A(n_207), .Y(n_248) );
INVx2_ASAP7_75t_L g249 ( .A(n_215), .Y(n_249) );
NOR2xp33_ASAP7_75t_L g250 ( .A(n_205), .B(n_146), .Y(n_250) );
NAND2xp5_ASAP7_75t_SL g251 ( .A(n_214), .B(n_158), .Y(n_251) );
INVx1_ASAP7_75t_L g252 ( .A(n_222), .Y(n_252) );
INVx2_ASAP7_75t_L g253 ( .A(n_224), .Y(n_253) );
AOI22xp5_ASAP7_75t_L g254 ( .A1(n_211), .A2(n_160), .B1(n_130), .B2(n_135), .Y(n_254) );
NAND2xp5_ASAP7_75t_L g255 ( .A(n_203), .B(n_160), .Y(n_255) );
INVx2_ASAP7_75t_SL g256 ( .A(n_172), .Y(n_256) );
AOI22xp5_ASAP7_75t_L g257 ( .A1(n_211), .A2(n_135), .B1(n_150), .B2(n_158), .Y(n_257) );
NAND2x1p5_ASAP7_75t_L g258 ( .A(n_202), .B(n_158), .Y(n_258) );
INVx4_ASAP7_75t_L g259 ( .A(n_172), .Y(n_259) );
AND2x2_ASAP7_75t_L g260 ( .A(n_198), .B(n_150), .Y(n_260) );
INVx1_ASAP7_75t_L g261 ( .A(n_223), .Y(n_261) );
NAND2xp5_ASAP7_75t_L g262 ( .A(n_203), .B(n_149), .Y(n_262) );
AND2x6_ASAP7_75t_SL g263 ( .A(n_221), .B(n_9), .Y(n_263) );
NAND2xp5_ASAP7_75t_SL g264 ( .A(n_225), .B(n_149), .Y(n_264) );
OR2x6_ASAP7_75t_L g265 ( .A(n_219), .B(n_149), .Y(n_265) );
AND2x4_ASAP7_75t_L g266 ( .A(n_198), .B(n_149), .Y(n_266) );
INVx1_ASAP7_75t_L g267 ( .A(n_204), .Y(n_267) );
INVx1_ASAP7_75t_L g268 ( .A(n_170), .Y(n_268) );
AO22x1_ASAP7_75t_L g269 ( .A1(n_182), .A2(n_149), .B1(n_143), .B2(n_142), .Y(n_269) );
OAI22xp5_ASAP7_75t_L g270 ( .A1(n_198), .A2(n_143), .B1(n_142), .B2(n_13), .Y(n_270) );
OAI22xp5_ASAP7_75t_L g271 ( .A1(n_171), .A2(n_143), .B1(n_142), .B2(n_13), .Y(n_271) );
OR2x2_ASAP7_75t_SL g272 ( .A(n_178), .B(n_10), .Y(n_272) );
INVx2_ASAP7_75t_L g273 ( .A(n_197), .Y(n_273) );
AND2x4_ASAP7_75t_L g274 ( .A(n_192), .B(n_143), .Y(n_274) );
INVxp67_ASAP7_75t_L g275 ( .A(n_206), .Y(n_275) );
NAND2xp5_ASAP7_75t_SL g276 ( .A(n_225), .B(n_143), .Y(n_276) );
BUFx6f_ASAP7_75t_L g277 ( .A(n_187), .Y(n_277) );
NAND2x1_ASAP7_75t_L g278 ( .A(n_174), .B(n_142), .Y(n_278) );
NAND2xp5_ASAP7_75t_L g279 ( .A(n_206), .B(n_10), .Y(n_279) );
OAI22xp5_ASAP7_75t_L g280 ( .A1(n_229), .A2(n_12), .B1(n_14), .B2(n_15), .Y(n_280) );
O2A1O1Ixp33_ASAP7_75t_L g281 ( .A1(n_177), .A2(n_14), .B(n_15), .C(n_16), .Y(n_281) );
AOI22xp33_ASAP7_75t_SL g282 ( .A1(n_181), .A2(n_17), .B1(n_18), .B2(n_20), .Y(n_282) );
AND2x2_ASAP7_75t_L g283 ( .A(n_196), .B(n_17), .Y(n_283) );
OR2x2_ASAP7_75t_L g284 ( .A(n_199), .B(n_18), .Y(n_284) );
NAND2xp5_ASAP7_75t_L g285 ( .A(n_213), .B(n_20), .Y(n_285) );
AOI22xp33_ASAP7_75t_L g286 ( .A1(n_180), .A2(n_21), .B1(n_39), .B2(n_43), .Y(n_286) );
AND2x4_ASAP7_75t_L g287 ( .A(n_179), .B(n_21), .Y(n_287) );
AOI22xp33_ASAP7_75t_L g288 ( .A1(n_189), .A2(n_44), .B1(n_58), .B2(n_65), .Y(n_288) );
INVx1_ASAP7_75t_L g289 ( .A(n_183), .Y(n_289) );
AND2x2_ASAP7_75t_L g290 ( .A(n_196), .B(n_66), .Y(n_290) );
NOR2xp33_ASAP7_75t_L g291 ( .A(n_201), .B(n_68), .Y(n_291) );
AND2x2_ASAP7_75t_L g292 ( .A(n_196), .B(n_71), .Y(n_292) );
AND2x4_ASAP7_75t_L g293 ( .A(n_179), .B(n_175), .Y(n_293) );
NAND2xp5_ASAP7_75t_SL g294 ( .A(n_194), .B(n_208), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g295 ( .A(n_189), .B(n_216), .Y(n_295) );
AOI22xp5_ASAP7_75t_L g296 ( .A1(n_200), .A2(n_175), .B1(n_181), .B2(n_210), .Y(n_296) );
NAND2xp5_ASAP7_75t_SL g297 ( .A(n_194), .B(n_208), .Y(n_297) );
A2O1A1Ixp33_ASAP7_75t_SL g298 ( .A1(n_291), .A2(n_228), .B(n_197), .C(n_226), .Y(n_298) );
INVx1_ASAP7_75t_L g299 ( .A(n_268), .Y(n_299) );
NOR2xp33_ASAP7_75t_R g300 ( .A(n_232), .B(n_200), .Y(n_300) );
AOI21xp5_ASAP7_75t_L g301 ( .A1(n_236), .A2(n_191), .B(n_193), .Y(n_301) );
AOI21xp5_ASAP7_75t_L g302 ( .A1(n_255), .A2(n_191), .B(n_193), .Y(n_302) );
NAND2xp5_ASAP7_75t_L g303 ( .A(n_275), .B(n_200), .Y(n_303) );
BUFx2_ASAP7_75t_L g304 ( .A(n_265), .Y(n_304) );
INVx1_ASAP7_75t_L g305 ( .A(n_267), .Y(n_305) );
CKINVDCx5p33_ASAP7_75t_R g306 ( .A(n_263), .Y(n_306) );
INVx1_ASAP7_75t_L g307 ( .A(n_252), .Y(n_307) );
INVx1_ASAP7_75t_L g308 ( .A(n_260), .Y(n_308) );
BUFx6f_ASAP7_75t_L g309 ( .A(n_277), .Y(n_309) );
NAND2xp5_ASAP7_75t_L g310 ( .A(n_275), .B(n_200), .Y(n_310) );
AOI21xp5_ASAP7_75t_L g311 ( .A1(n_238), .A2(n_251), .B(n_244), .Y(n_311) );
OAI21xp5_ASAP7_75t_L g312 ( .A1(n_295), .A2(n_194), .B(n_187), .Y(n_312) );
INVx2_ASAP7_75t_SL g313 ( .A(n_283), .Y(n_313) );
OAI22xp5_ASAP7_75t_L g314 ( .A1(n_237), .A2(n_216), .B1(n_201), .B2(n_212), .Y(n_314) );
BUFx2_ASAP7_75t_L g315 ( .A(n_265), .Y(n_315) );
INVx1_ASAP7_75t_L g316 ( .A(n_246), .Y(n_316) );
OAI22xp5_ASAP7_75t_L g317 ( .A1(n_237), .A2(n_212), .B1(n_210), .B2(n_228), .Y(n_317) );
NAND2x1p5_ASAP7_75t_L g318 ( .A(n_259), .B(n_183), .Y(n_318) );
AOI21xp5_ASAP7_75t_L g319 ( .A1(n_244), .A2(n_231), .B(n_179), .Y(n_319) );
OAI22xp5_ASAP7_75t_L g320 ( .A1(n_233), .A2(n_231), .B1(n_200), .B2(n_176), .Y(n_320) );
O2A1O1Ixp33_ASAP7_75t_SL g321 ( .A1(n_276), .A2(n_176), .B(n_226), .C(n_220), .Y(n_321) );
NOR2xp33_ASAP7_75t_L g322 ( .A(n_235), .B(n_181), .Y(n_322) );
NOR2xp33_ASAP7_75t_L g323 ( .A(n_240), .B(n_181), .Y(n_323) );
OR2x2_ASAP7_75t_L g324 ( .A(n_241), .B(n_190), .Y(n_324) );
A2O1A1Ixp33_ASAP7_75t_L g325 ( .A1(n_261), .A2(n_195), .B(n_209), .C(n_217), .Y(n_325) );
INVx1_ASAP7_75t_SL g326 ( .A(n_259), .Y(n_326) );
INVx1_ASAP7_75t_L g327 ( .A(n_266), .Y(n_327) );
OAI21xp33_ASAP7_75t_L g328 ( .A1(n_243), .A2(n_190), .B(n_195), .Y(n_328) );
NOR2xp33_ASAP7_75t_L g329 ( .A(n_239), .B(n_181), .Y(n_329) );
AND2x4_ASAP7_75t_SL g330 ( .A(n_287), .B(n_220), .Y(n_330) );
NAND3xp33_ASAP7_75t_SL g331 ( .A(n_281), .B(n_209), .C(n_217), .Y(n_331) );
O2A1O1Ixp5_ASAP7_75t_L g332 ( .A1(n_279), .A2(n_285), .B(n_269), .C(n_233), .Y(n_332) );
INVx4_ASAP7_75t_L g333 ( .A(n_287), .Y(n_333) );
AOI21xp5_ASAP7_75t_L g334 ( .A1(n_251), .A2(n_276), .B(n_294), .Y(n_334) );
INVxp67_ASAP7_75t_L g335 ( .A(n_250), .Y(n_335) );
AOI22xp5_ASAP7_75t_L g336 ( .A1(n_234), .A2(n_254), .B1(n_257), .B2(n_265), .Y(n_336) );
OAI21xp33_ASAP7_75t_L g337 ( .A1(n_250), .A2(n_247), .B(n_284), .Y(n_337) );
NOR2xp33_ASAP7_75t_L g338 ( .A(n_239), .B(n_289), .Y(n_338) );
AOI21xp5_ASAP7_75t_L g339 ( .A1(n_294), .A2(n_264), .B(n_297), .Y(n_339) );
O2A1O1Ixp33_ASAP7_75t_L g340 ( .A1(n_242), .A2(n_271), .B(n_270), .C(n_280), .Y(n_340) );
AOI21xp5_ASAP7_75t_L g341 ( .A1(n_262), .A2(n_247), .B(n_293), .Y(n_341) );
CKINVDCx5p33_ASAP7_75t_R g342 ( .A(n_239), .Y(n_342) );
AOI222xp33_ASAP7_75t_L g343 ( .A1(n_266), .A2(n_274), .B1(n_248), .B2(n_249), .C1(n_253), .C2(n_286), .Y(n_343) );
A2O1A1Ixp33_ASAP7_75t_L g344 ( .A1(n_291), .A2(n_296), .B(n_274), .C(n_292), .Y(n_344) );
AOI22xp5_ASAP7_75t_L g345 ( .A1(n_245), .A2(n_256), .B1(n_293), .B2(n_290), .Y(n_345) );
NAND2xp5_ASAP7_75t_SL g346 ( .A(n_277), .B(n_258), .Y(n_346) );
INVx1_ASAP7_75t_L g347 ( .A(n_258), .Y(n_347) );
INVx1_ASAP7_75t_L g348 ( .A(n_272), .Y(n_348) );
AND2x4_ASAP7_75t_L g349 ( .A(n_277), .B(n_288), .Y(n_349) );
OAI22xp33_ASAP7_75t_SL g350 ( .A1(n_348), .A2(n_282), .B1(n_286), .B2(n_288), .Y(n_350) );
O2A1O1Ixp33_ASAP7_75t_SL g351 ( .A1(n_344), .A2(n_278), .B(n_273), .C(n_282), .Y(n_351) );
BUFx2_ASAP7_75t_L g352 ( .A(n_304), .Y(n_352) );
AOI21xp5_ASAP7_75t_L g353 ( .A1(n_311), .A2(n_277), .B(n_302), .Y(n_353) );
AO32x2_ASAP7_75t_L g354 ( .A1(n_317), .A2(n_314), .A3(n_320), .B1(n_313), .B2(n_333), .Y(n_354) );
BUFx6f_ASAP7_75t_L g355 ( .A(n_309), .Y(n_355) );
NAND2xp5_ASAP7_75t_L g356 ( .A(n_335), .B(n_316), .Y(n_356) );
INVx1_ASAP7_75t_SL g357 ( .A(n_326), .Y(n_357) );
NOR2xp33_ASAP7_75t_L g358 ( .A(n_324), .B(n_328), .Y(n_358) );
INVx1_ASAP7_75t_L g359 ( .A(n_305), .Y(n_359) );
AOI22xp33_ASAP7_75t_L g360 ( .A1(n_337), .A2(n_308), .B1(n_327), .B2(n_315), .Y(n_360) );
INVx1_ASAP7_75t_L g361 ( .A(n_299), .Y(n_361) );
NAND2xp5_ASAP7_75t_L g362 ( .A(n_307), .B(n_329), .Y(n_362) );
INVx1_ASAP7_75t_L g363 ( .A(n_318), .Y(n_363) );
AOI21xp5_ASAP7_75t_L g364 ( .A1(n_298), .A2(n_312), .B(n_334), .Y(n_364) );
INVx2_ASAP7_75t_L g365 ( .A(n_347), .Y(n_365) );
AOI21xp5_ASAP7_75t_L g366 ( .A1(n_303), .A2(n_310), .B(n_301), .Y(n_366) );
NAND3x1_ASAP7_75t_L g367 ( .A(n_338), .B(n_336), .C(n_306), .Y(n_367) );
AOI21xp5_ASAP7_75t_L g368 ( .A1(n_319), .A2(n_346), .B(n_321), .Y(n_368) );
NAND2xp5_ASAP7_75t_L g369 ( .A(n_326), .B(n_343), .Y(n_369) );
AOI22xp5_ASAP7_75t_L g370 ( .A1(n_342), .A2(n_333), .B1(n_322), .B2(n_323), .Y(n_370) );
NAND3xp33_ASAP7_75t_L g371 ( .A(n_343), .B(n_332), .C(n_340), .Y(n_371) );
AND2x2_ASAP7_75t_L g372 ( .A(n_300), .B(n_318), .Y(n_372) );
NOR2xp33_ASAP7_75t_L g373 ( .A(n_345), .B(n_349), .Y(n_373) );
AOI21xp5_ASAP7_75t_L g374 ( .A1(n_325), .A2(n_341), .B(n_339), .Y(n_374) );
AO31x2_ASAP7_75t_L g375 ( .A1(n_349), .A2(n_331), .A3(n_309), .B(n_330), .Y(n_375) );
AOI21xp5_ASAP7_75t_L g376 ( .A1(n_309), .A2(n_236), .B(n_255), .Y(n_376) );
AOI21xp5_ASAP7_75t_L g377 ( .A1(n_311), .A2(n_236), .B(n_255), .Y(n_377) );
O2A1O1Ixp33_ASAP7_75t_L g378 ( .A1(n_335), .A2(n_337), .B(n_275), .C(n_284), .Y(n_378) );
AOI21xp5_ASAP7_75t_L g379 ( .A1(n_311), .A2(n_236), .B(n_255), .Y(n_379) );
AOI22xp33_ASAP7_75t_L g380 ( .A1(n_324), .A2(n_234), .B1(n_211), .B2(n_186), .Y(n_380) );
BUFx12f_ASAP7_75t_L g381 ( .A(n_306), .Y(n_381) );
BUFx6f_ASAP7_75t_L g382 ( .A(n_309), .Y(n_382) );
AOI22xp33_ASAP7_75t_L g383 ( .A1(n_358), .A2(n_380), .B1(n_373), .B2(n_369), .Y(n_383) );
AO21x2_ASAP7_75t_L g384 ( .A1(n_364), .A2(n_371), .B(n_374), .Y(n_384) );
INVx1_ASAP7_75t_L g385 ( .A(n_359), .Y(n_385) );
AOI21xp5_ASAP7_75t_L g386 ( .A1(n_377), .A2(n_379), .B(n_368), .Y(n_386) );
INVx2_ASAP7_75t_L g387 ( .A(n_355), .Y(n_387) );
INVx2_ASAP7_75t_L g388 ( .A(n_355), .Y(n_388) );
INVx1_ASAP7_75t_L g389 ( .A(n_361), .Y(n_389) );
BUFx8_ASAP7_75t_L g390 ( .A(n_381), .Y(n_390) );
NAND2xp5_ASAP7_75t_L g391 ( .A(n_378), .B(n_356), .Y(n_391) );
AOI21xp5_ASAP7_75t_L g392 ( .A1(n_353), .A2(n_351), .B(n_376), .Y(n_392) );
INVx1_ASAP7_75t_L g393 ( .A(n_362), .Y(n_393) );
OAI21xp5_ASAP7_75t_L g394 ( .A1(n_371), .A2(n_366), .B(n_350), .Y(n_394) );
NAND2xp5_ASAP7_75t_L g395 ( .A(n_360), .B(n_350), .Y(n_395) );
OAI21x1_ASAP7_75t_L g396 ( .A1(n_363), .A2(n_354), .B(n_375), .Y(n_396) );
INVx1_ASAP7_75t_L g397 ( .A(n_365), .Y(n_397) );
OAI22xp5_ASAP7_75t_SL g398 ( .A1(n_357), .A2(n_352), .B1(n_370), .B2(n_367), .Y(n_398) );
INVx1_ASAP7_75t_L g399 ( .A(n_375), .Y(n_399) );
INVx1_ASAP7_75t_L g400 ( .A(n_375), .Y(n_400) );
INVx2_ASAP7_75t_SL g401 ( .A(n_357), .Y(n_401) );
INVx1_ASAP7_75t_L g402 ( .A(n_354), .Y(n_402) );
AOI21xp5_ASAP7_75t_L g403 ( .A1(n_355), .A2(n_382), .B(n_354), .Y(n_403) );
OR2x2_ASAP7_75t_L g404 ( .A(n_372), .B(n_382), .Y(n_404) );
BUFx3_ASAP7_75t_L g405 ( .A(n_382), .Y(n_405) );
OA21x2_ASAP7_75t_L g406 ( .A1(n_364), .A2(n_374), .B(n_371), .Y(n_406) );
OAI21xp5_ASAP7_75t_L g407 ( .A1(n_371), .A2(n_344), .B(n_364), .Y(n_407) );
OAI21x1_ASAP7_75t_L g408 ( .A1(n_364), .A2(n_374), .B(n_368), .Y(n_408) );
OA21x2_ASAP7_75t_L g409 ( .A1(n_364), .A2(n_374), .B(n_371), .Y(n_409) );
A2O1A1Ixp33_ASAP7_75t_L g410 ( .A1(n_378), .A2(n_373), .B(n_371), .C(n_185), .Y(n_410) );
INVx2_ASAP7_75t_L g411 ( .A(n_384), .Y(n_411) );
INVx1_ASAP7_75t_L g412 ( .A(n_399), .Y(n_412) );
AND2x2_ASAP7_75t_SL g413 ( .A(n_395), .B(n_399), .Y(n_413) );
AND2x2_ASAP7_75t_L g414 ( .A(n_394), .B(n_395), .Y(n_414) );
HB1xp67_ASAP7_75t_L g415 ( .A(n_401), .Y(n_415) );
AO21x2_ASAP7_75t_L g416 ( .A1(n_386), .A2(n_407), .B(n_394), .Y(n_416) );
OR2x2_ASAP7_75t_L g417 ( .A(n_391), .B(n_383), .Y(n_417) );
INVx1_ASAP7_75t_L g418 ( .A(n_400), .Y(n_418) );
INVx3_ASAP7_75t_L g419 ( .A(n_405), .Y(n_419) );
INVx4_ASAP7_75t_L g420 ( .A(n_405), .Y(n_420) );
INVx2_ASAP7_75t_L g421 ( .A(n_384), .Y(n_421) );
INVx1_ASAP7_75t_L g422 ( .A(n_400), .Y(n_422) );
AO21x2_ASAP7_75t_L g423 ( .A1(n_407), .A2(n_392), .B(n_408), .Y(n_423) );
AOI22xp33_ASAP7_75t_L g424 ( .A1(n_398), .A2(n_391), .B1(n_393), .B2(n_385), .Y(n_424) );
INVx3_ASAP7_75t_L g425 ( .A(n_405), .Y(n_425) );
BUFx2_ASAP7_75t_L g426 ( .A(n_401), .Y(n_426) );
INVx2_ASAP7_75t_SL g427 ( .A(n_404), .Y(n_427) );
HB1xp67_ASAP7_75t_L g428 ( .A(n_387), .Y(n_428) );
HB1xp67_ASAP7_75t_L g429 ( .A(n_387), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_384), .Y(n_430) );
OAI22xp5_ASAP7_75t_L g431 ( .A1(n_410), .A2(n_398), .B1(n_393), .B2(n_389), .Y(n_431) );
NAND2xp5_ASAP7_75t_L g432 ( .A(n_385), .B(n_389), .Y(n_432) );
AND2x2_ASAP7_75t_L g433 ( .A(n_384), .B(n_409), .Y(n_433) );
INVx2_ASAP7_75t_SL g434 ( .A(n_404), .Y(n_434) );
INVx1_ASAP7_75t_L g435 ( .A(n_406), .Y(n_435) );
OAI21xp5_ASAP7_75t_L g436 ( .A1(n_408), .A2(n_396), .B(n_406), .Y(n_436) );
AO21x2_ASAP7_75t_L g437 ( .A1(n_403), .A2(n_402), .B(n_396), .Y(n_437) );
BUFx2_ASAP7_75t_L g438 ( .A(n_387), .Y(n_438) );
AOI22xp5_ASAP7_75t_L g439 ( .A1(n_397), .A2(n_406), .B1(n_409), .B2(n_402), .Y(n_439) );
INVx2_ASAP7_75t_L g440 ( .A(n_406), .Y(n_440) );
INVxp67_ASAP7_75t_L g441 ( .A(n_397), .Y(n_441) );
AO21x2_ASAP7_75t_L g442 ( .A1(n_388), .A2(n_409), .B(n_390), .Y(n_442) );
INVx4_ASAP7_75t_L g443 ( .A(n_388), .Y(n_443) );
OR2x2_ASAP7_75t_L g444 ( .A(n_409), .B(n_388), .Y(n_444) );
INVx1_ASAP7_75t_L g445 ( .A(n_390), .Y(n_445) );
INVx1_ASAP7_75t_L g446 ( .A(n_412), .Y(n_446) );
BUFx3_ASAP7_75t_L g447 ( .A(n_420), .Y(n_447) );
INVx1_ASAP7_75t_SL g448 ( .A(n_426), .Y(n_448) );
AND2x2_ASAP7_75t_L g449 ( .A(n_433), .B(n_390), .Y(n_449) );
AND2x2_ASAP7_75t_L g450 ( .A(n_433), .B(n_390), .Y(n_450) );
NAND2xp5_ASAP7_75t_L g451 ( .A(n_414), .B(n_417), .Y(n_451) );
AND2x4_ASAP7_75t_L g452 ( .A(n_442), .B(n_433), .Y(n_452) );
INVx1_ASAP7_75t_L g453 ( .A(n_412), .Y(n_453) );
AND2x2_ASAP7_75t_L g454 ( .A(n_414), .B(n_416), .Y(n_454) );
INVx2_ASAP7_75t_L g455 ( .A(n_440), .Y(n_455) );
AND2x2_ASAP7_75t_L g456 ( .A(n_414), .B(n_416), .Y(n_456) );
BUFx2_ASAP7_75t_L g457 ( .A(n_442), .Y(n_457) );
INVx1_ASAP7_75t_L g458 ( .A(n_412), .Y(n_458) );
AND2x2_ASAP7_75t_L g459 ( .A(n_416), .B(n_430), .Y(n_459) );
AOI22xp5_ASAP7_75t_L g460 ( .A1(n_431), .A2(n_417), .B1(n_424), .B2(n_441), .Y(n_460) );
AND2x2_ASAP7_75t_L g461 ( .A(n_416), .B(n_430), .Y(n_461) );
AND2x2_ASAP7_75t_L g462 ( .A(n_416), .B(n_430), .Y(n_462) );
AOI22xp33_ASAP7_75t_L g463 ( .A1(n_417), .A2(n_431), .B1(n_424), .B2(n_445), .Y(n_463) );
BUFx2_ASAP7_75t_L g464 ( .A(n_442), .Y(n_464) );
NOR2xp33_ASAP7_75t_L g465 ( .A(n_445), .B(n_427), .Y(n_465) );
AND2x2_ASAP7_75t_L g466 ( .A(n_439), .B(n_435), .Y(n_466) );
NAND2xp5_ASAP7_75t_L g467 ( .A(n_432), .B(n_441), .Y(n_467) );
NAND2xp5_ASAP7_75t_L g468 ( .A(n_432), .B(n_418), .Y(n_468) );
AND2x2_ASAP7_75t_L g469 ( .A(n_439), .B(n_435), .Y(n_469) );
NOR2x1_ASAP7_75t_SL g470 ( .A(n_442), .B(n_420), .Y(n_470) );
AND2x4_ASAP7_75t_L g471 ( .A(n_442), .B(n_440), .Y(n_471) );
CKINVDCx5p33_ASAP7_75t_R g472 ( .A(n_445), .Y(n_472) );
INVx1_ASAP7_75t_L g473 ( .A(n_418), .Y(n_473) );
INVx1_ASAP7_75t_L g474 ( .A(n_418), .Y(n_474) );
HB1xp67_ASAP7_75t_L g475 ( .A(n_428), .Y(n_475) );
INVx1_ASAP7_75t_L g476 ( .A(n_422), .Y(n_476) );
BUFx2_ASAP7_75t_L g477 ( .A(n_420), .Y(n_477) );
INVx2_ASAP7_75t_L g478 ( .A(n_444), .Y(n_478) );
INVx1_ASAP7_75t_L g479 ( .A(n_422), .Y(n_479) );
AND2x2_ASAP7_75t_L g480 ( .A(n_435), .B(n_422), .Y(n_480) );
AND2x4_ASAP7_75t_L g481 ( .A(n_436), .B(n_444), .Y(n_481) );
BUFx2_ASAP7_75t_L g482 ( .A(n_444), .Y(n_482) );
INVx1_ASAP7_75t_L g483 ( .A(n_411), .Y(n_483) );
INVx1_ASAP7_75t_L g484 ( .A(n_411), .Y(n_484) );
NAND2xp5_ASAP7_75t_L g485 ( .A(n_413), .B(n_429), .Y(n_485) );
INVx1_ASAP7_75t_L g486 ( .A(n_411), .Y(n_486) );
INVx1_ASAP7_75t_L g487 ( .A(n_421), .Y(n_487) );
INVx3_ASAP7_75t_SL g488 ( .A(n_420), .Y(n_488) );
BUFx3_ASAP7_75t_L g489 ( .A(n_420), .Y(n_489) );
OR2x2_ASAP7_75t_L g490 ( .A(n_421), .B(n_415), .Y(n_490) );
INVx2_ASAP7_75t_L g491 ( .A(n_455), .Y(n_491) );
AND2x2_ASAP7_75t_L g492 ( .A(n_454), .B(n_413), .Y(n_492) );
INVx1_ASAP7_75t_L g493 ( .A(n_446), .Y(n_493) );
NOR2xp33_ASAP7_75t_L g494 ( .A(n_472), .B(n_434), .Y(n_494) );
OR2x2_ASAP7_75t_L g495 ( .A(n_482), .B(n_423), .Y(n_495) );
AND2x2_ASAP7_75t_L g496 ( .A(n_454), .B(n_413), .Y(n_496) );
OR2x2_ASAP7_75t_L g497 ( .A(n_482), .B(n_423), .Y(n_497) );
INVx1_ASAP7_75t_L g498 ( .A(n_446), .Y(n_498) );
INVx1_ASAP7_75t_L g499 ( .A(n_453), .Y(n_499) );
AND2x2_ASAP7_75t_L g500 ( .A(n_454), .B(n_413), .Y(n_500) );
AND2x2_ASAP7_75t_L g501 ( .A(n_456), .B(n_480), .Y(n_501) );
OR2x2_ASAP7_75t_L g502 ( .A(n_482), .B(n_423), .Y(n_502) );
AND2x2_ASAP7_75t_L g503 ( .A(n_456), .B(n_436), .Y(n_503) );
AND2x4_ASAP7_75t_L g504 ( .A(n_452), .B(n_423), .Y(n_504) );
AND2x2_ASAP7_75t_L g505 ( .A(n_456), .B(n_437), .Y(n_505) );
INVx1_ASAP7_75t_L g506 ( .A(n_453), .Y(n_506) );
AND2x2_ASAP7_75t_L g507 ( .A(n_480), .B(n_437), .Y(n_507) );
NAND2xp5_ASAP7_75t_L g508 ( .A(n_465), .B(n_434), .Y(n_508) );
HB1xp67_ASAP7_75t_L g509 ( .A(n_475), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_465), .B(n_434), .Y(n_510) );
OR2x2_ASAP7_75t_L g511 ( .A(n_451), .B(n_423), .Y(n_511) );
AND2x4_ASAP7_75t_L g512 ( .A(n_452), .B(n_437), .Y(n_512) );
BUFx6f_ASAP7_75t_L g513 ( .A(n_471), .Y(n_513) );
INVx2_ASAP7_75t_SL g514 ( .A(n_488), .Y(n_514) );
AND2x4_ASAP7_75t_L g515 ( .A(n_452), .B(n_437), .Y(n_515) );
INVx2_ASAP7_75t_L g516 ( .A(n_455), .Y(n_516) );
AND2x2_ASAP7_75t_L g517 ( .A(n_480), .B(n_437), .Y(n_517) );
AND2x4_ASAP7_75t_L g518 ( .A(n_452), .B(n_443), .Y(n_518) );
INVx2_ASAP7_75t_SL g519 ( .A(n_488), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_449), .B(n_427), .Y(n_520) );
INVx1_ASAP7_75t_L g521 ( .A(n_458), .Y(n_521) );
INVx1_ASAP7_75t_L g522 ( .A(n_458), .Y(n_522) );
INVx1_ASAP7_75t_L g523 ( .A(n_473), .Y(n_523) );
HB1xp67_ASAP7_75t_SL g524 ( .A(n_449), .Y(n_524) );
NAND2xp5_ASAP7_75t_L g525 ( .A(n_449), .B(n_427), .Y(n_525) );
INVx1_ASAP7_75t_L g526 ( .A(n_473), .Y(n_526) );
NOR2x1_ASAP7_75t_L g527 ( .A(n_450), .B(n_426), .Y(n_527) );
AND2x2_ASAP7_75t_L g528 ( .A(n_466), .B(n_428), .Y(n_528) );
AND2x4_ASAP7_75t_L g529 ( .A(n_452), .B(n_443), .Y(n_529) );
OR2x2_ASAP7_75t_L g530 ( .A(n_451), .B(n_415), .Y(n_530) );
AND2x2_ASAP7_75t_L g531 ( .A(n_466), .B(n_429), .Y(n_531) );
INVx1_ASAP7_75t_L g532 ( .A(n_474), .Y(n_532) );
BUFx3_ASAP7_75t_L g533 ( .A(n_488), .Y(n_533) );
INVx1_ASAP7_75t_L g534 ( .A(n_474), .Y(n_534) );
INVx1_ASAP7_75t_L g535 ( .A(n_476), .Y(n_535) );
INVx1_ASAP7_75t_L g536 ( .A(n_476), .Y(n_536) );
OR2x2_ASAP7_75t_L g537 ( .A(n_475), .B(n_426), .Y(n_537) );
AND2x2_ASAP7_75t_L g538 ( .A(n_466), .B(n_438), .Y(n_538) );
AND2x2_ASAP7_75t_L g539 ( .A(n_469), .B(n_438), .Y(n_539) );
NAND2x1p5_ASAP7_75t_L g540 ( .A(n_477), .B(n_419), .Y(n_540) );
NAND2xp5_ASAP7_75t_L g541 ( .A(n_450), .B(n_438), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_450), .B(n_443), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_463), .B(n_443), .Y(n_543) );
NOR2xp33_ASAP7_75t_L g544 ( .A(n_488), .B(n_419), .Y(n_544) );
AND2x2_ASAP7_75t_L g545 ( .A(n_501), .B(n_461), .Y(n_545) );
OR2x2_ASAP7_75t_L g546 ( .A(n_501), .B(n_530), .Y(n_546) );
AND2x2_ASAP7_75t_L g547 ( .A(n_503), .B(n_461), .Y(n_547) );
INVx1_ASAP7_75t_L g548 ( .A(n_493), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g549 ( .A(n_530), .B(n_460), .Y(n_549) );
OR2x2_ASAP7_75t_L g550 ( .A(n_511), .B(n_490), .Y(n_550) );
OR2x2_ASAP7_75t_L g551 ( .A(n_511), .B(n_490), .Y(n_551) );
OR2x2_ASAP7_75t_L g552 ( .A(n_503), .B(n_490), .Y(n_552) );
AOI222xp33_ASAP7_75t_L g553 ( .A1(n_492), .A2(n_463), .B1(n_462), .B2(n_461), .C1(n_459), .C2(n_469), .Y(n_553) );
OR2x2_ASAP7_75t_L g554 ( .A(n_507), .B(n_478), .Y(n_554) );
AND2x4_ASAP7_75t_L g555 ( .A(n_512), .B(n_470), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g556 ( .A(n_505), .B(n_460), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g557 ( .A(n_505), .B(n_528), .Y(n_557) );
NOR2xp33_ASAP7_75t_L g558 ( .A(n_524), .B(n_467), .Y(n_558) );
OA21x2_ASAP7_75t_L g559 ( .A1(n_543), .A2(n_464), .B(n_457), .Y(n_559) );
OR2x2_ASAP7_75t_L g560 ( .A(n_507), .B(n_478), .Y(n_560) );
INVx4_ASAP7_75t_L g561 ( .A(n_533), .Y(n_561) );
AND2x4_ASAP7_75t_L g562 ( .A(n_512), .B(n_470), .Y(n_562) );
NAND2x1p5_ASAP7_75t_L g563 ( .A(n_533), .B(n_477), .Y(n_563) );
AND2x2_ASAP7_75t_L g564 ( .A(n_517), .B(n_462), .Y(n_564) );
AND2x2_ASAP7_75t_L g565 ( .A(n_517), .B(n_462), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g566 ( .A(n_528), .B(n_479), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_531), .B(n_479), .Y(n_567) );
AND3x2_ASAP7_75t_L g568 ( .A(n_544), .B(n_464), .C(n_457), .Y(n_568) );
NAND2xp5_ASAP7_75t_L g569 ( .A(n_531), .B(n_459), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g570 ( .A(n_509), .B(n_459), .Y(n_570) );
INVx1_ASAP7_75t_L g571 ( .A(n_493), .Y(n_571) );
INVx1_ASAP7_75t_L g572 ( .A(n_498), .Y(n_572) );
INVx2_ASAP7_75t_L g573 ( .A(n_491), .Y(n_573) );
AND2x2_ASAP7_75t_L g574 ( .A(n_492), .B(n_469), .Y(n_574) );
AND2x2_ASAP7_75t_L g575 ( .A(n_496), .B(n_481), .Y(n_575) );
HB1xp67_ASAP7_75t_L g576 ( .A(n_537), .Y(n_576) );
INVx2_ASAP7_75t_L g577 ( .A(n_516), .Y(n_577) );
INVxp33_ASAP7_75t_L g578 ( .A(n_527), .Y(n_578) );
AND2x2_ASAP7_75t_L g579 ( .A(n_496), .B(n_481), .Y(n_579) );
OAI21xp5_ASAP7_75t_SL g580 ( .A1(n_514), .A2(n_467), .B(n_448), .Y(n_580) );
AND2x2_ASAP7_75t_SL g581 ( .A(n_518), .B(n_485), .Y(n_581) );
NOR2xp33_ASAP7_75t_L g582 ( .A(n_494), .B(n_447), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g583 ( .A(n_521), .B(n_468), .Y(n_583) );
HB1xp67_ASAP7_75t_L g584 ( .A(n_537), .Y(n_584) );
AND2x2_ASAP7_75t_L g585 ( .A(n_500), .B(n_481), .Y(n_585) );
INVx1_ASAP7_75t_L g586 ( .A(n_498), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g587 ( .A(n_536), .B(n_468), .Y(n_587) );
INVx1_ASAP7_75t_L g588 ( .A(n_499), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g589 ( .A(n_538), .B(n_478), .Y(n_589) );
AND2x4_ASAP7_75t_L g590 ( .A(n_512), .B(n_481), .Y(n_590) );
NAND4xp25_ASAP7_75t_L g591 ( .A(n_508), .B(n_485), .C(n_481), .D(n_471), .Y(n_591) );
AND2x2_ASAP7_75t_L g592 ( .A(n_500), .B(n_471), .Y(n_592) );
INVx1_ASAP7_75t_L g593 ( .A(n_499), .Y(n_593) );
INVxp67_ASAP7_75t_L g594 ( .A(n_514), .Y(n_594) );
NAND2x1p5_ASAP7_75t_L g595 ( .A(n_561), .B(n_519), .Y(n_595) );
NAND4xp25_ASAP7_75t_L g596 ( .A(n_553), .B(n_510), .C(n_504), .D(n_515), .Y(n_596) );
NAND2xp5_ASAP7_75t_L g597 ( .A(n_564), .B(n_526), .Y(n_597) );
AOI22xp5_ASAP7_75t_L g598 ( .A1(n_558), .A2(n_519), .B1(n_515), .B2(n_504), .Y(n_598) );
AND2x2_ASAP7_75t_L g599 ( .A(n_545), .B(n_529), .Y(n_599) );
INVx1_ASAP7_75t_L g600 ( .A(n_576), .Y(n_600) );
NAND2x1_ASAP7_75t_L g601 ( .A(n_561), .B(n_529), .Y(n_601) );
INVx1_ASAP7_75t_L g602 ( .A(n_584), .Y(n_602) );
OAI21xp33_ASAP7_75t_L g603 ( .A1(n_591), .A2(n_515), .B(n_504), .Y(n_603) );
INVxp67_ASAP7_75t_SL g604 ( .A(n_563), .Y(n_604) );
INVx1_ASAP7_75t_L g605 ( .A(n_546), .Y(n_605) );
NAND2x2_ASAP7_75t_L g606 ( .A(n_556), .B(n_489), .Y(n_606) );
INVx1_ASAP7_75t_L g607 ( .A(n_546), .Y(n_607) );
INVx1_ASAP7_75t_L g608 ( .A(n_548), .Y(n_608) );
OR2x2_ASAP7_75t_L g609 ( .A(n_552), .B(n_539), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g610 ( .A(n_564), .B(n_538), .Y(n_610) );
AOI21xp33_ASAP7_75t_SL g611 ( .A1(n_563), .A2(n_540), .B(n_542), .Y(n_611) );
AND2x2_ASAP7_75t_L g612 ( .A(n_545), .B(n_529), .Y(n_612) );
INVx2_ASAP7_75t_L g613 ( .A(n_561), .Y(n_613) );
INVx2_ASAP7_75t_L g614 ( .A(n_563), .Y(n_614) );
NAND2x1p5_ASAP7_75t_L g615 ( .A(n_581), .B(n_447), .Y(n_615) );
NAND2xp5_ASAP7_75t_L g616 ( .A(n_565), .B(n_506), .Y(n_616) );
NAND3xp33_ASAP7_75t_L g617 ( .A(n_580), .B(n_513), .C(n_502), .Y(n_617) );
OR2x2_ASAP7_75t_L g618 ( .A(n_552), .B(n_539), .Y(n_618) );
NAND2xp5_ASAP7_75t_L g619 ( .A(n_565), .B(n_506), .Y(n_619) );
NAND2x1p5_ASAP7_75t_L g620 ( .A(n_581), .B(n_447), .Y(n_620) );
INVx1_ASAP7_75t_L g621 ( .A(n_571), .Y(n_621) );
INVx1_ASAP7_75t_L g622 ( .A(n_572), .Y(n_622) );
NAND2xp5_ASAP7_75t_L g623 ( .A(n_547), .B(n_523), .Y(n_623) );
OAI21xp5_ASAP7_75t_L g624 ( .A1(n_578), .A2(n_540), .B(n_448), .Y(n_624) );
AND2x2_ASAP7_75t_L g625 ( .A(n_547), .B(n_518), .Y(n_625) );
NOR2xp67_ASAP7_75t_L g626 ( .A(n_555), .B(n_518), .Y(n_626) );
NAND2xp5_ASAP7_75t_L g627 ( .A(n_569), .B(n_526), .Y(n_627) );
AND2x2_ASAP7_75t_SL g628 ( .A(n_555), .B(n_513), .Y(n_628) );
INVx1_ASAP7_75t_L g629 ( .A(n_586), .Y(n_629) );
OAI222xp33_ASAP7_75t_L g630 ( .A1(n_594), .A2(n_541), .B1(n_540), .B2(n_525), .C1(n_520), .C2(n_502), .Y(n_630) );
INVx1_ASAP7_75t_L g631 ( .A(n_588), .Y(n_631) );
NAND2xp5_ASAP7_75t_L g632 ( .A(n_549), .B(n_535), .Y(n_632) );
OR2x2_ASAP7_75t_L g633 ( .A(n_609), .B(n_570), .Y(n_633) );
INVx1_ASAP7_75t_L g634 ( .A(n_600), .Y(n_634) );
INVx1_ASAP7_75t_L g635 ( .A(n_602), .Y(n_635) );
AND2x2_ASAP7_75t_L g636 ( .A(n_605), .B(n_592), .Y(n_636) );
NAND2xp5_ASAP7_75t_L g637 ( .A(n_607), .B(n_574), .Y(n_637) );
OAI32xp33_ASAP7_75t_L g638 ( .A1(n_596), .A2(n_578), .A3(n_582), .B1(n_550), .B2(n_551), .Y(n_638) );
INVx1_ASAP7_75t_L g639 ( .A(n_597), .Y(n_639) );
INVx1_ASAP7_75t_L g640 ( .A(n_608), .Y(n_640) );
NOR2xp33_ASAP7_75t_L g641 ( .A(n_596), .B(n_557), .Y(n_641) );
INVx1_ASAP7_75t_L g642 ( .A(n_597), .Y(n_642) );
AND2x2_ASAP7_75t_L g643 ( .A(n_599), .B(n_592), .Y(n_643) );
AND2x2_ASAP7_75t_L g644 ( .A(n_612), .B(n_575), .Y(n_644) );
A2O1A1Ixp33_ASAP7_75t_SL g645 ( .A1(n_624), .A2(n_614), .B(n_613), .C(n_604), .Y(n_645) );
NAND2xp5_ASAP7_75t_L g646 ( .A(n_632), .B(n_574), .Y(n_646) );
NOR2xp33_ASAP7_75t_L g647 ( .A(n_616), .B(n_567), .Y(n_647) );
OAI31xp33_ASAP7_75t_L g648 ( .A1(n_615), .A2(n_562), .A3(n_555), .B(n_590), .Y(n_648) );
NAND2xp5_ASAP7_75t_L g649 ( .A(n_616), .B(n_585), .Y(n_649) );
INVx1_ASAP7_75t_L g650 ( .A(n_619), .Y(n_650) );
AOI221xp5_ASAP7_75t_L g651 ( .A1(n_603), .A2(n_575), .B1(n_585), .B2(n_579), .C(n_566), .Y(n_651) );
AOI221x1_ASAP7_75t_L g652 ( .A1(n_611), .A2(n_562), .B1(n_593), .B2(n_535), .C(n_534), .Y(n_652) );
OAI22xp5_ASAP7_75t_L g653 ( .A1(n_606), .A2(n_562), .B1(n_590), .B2(n_551), .Y(n_653) );
AND2x2_ASAP7_75t_L g654 ( .A(n_625), .B(n_579), .Y(n_654) );
AND2x2_ASAP7_75t_L g655 ( .A(n_619), .B(n_590), .Y(n_655) );
OAI22xp5_ASAP7_75t_L g656 ( .A1(n_641), .A2(n_626), .B1(n_615), .B2(n_620), .Y(n_656) );
INVx2_ASAP7_75t_L g657 ( .A(n_640), .Y(n_657) );
OAI211xp5_ASAP7_75t_SL g658 ( .A1(n_651), .A2(n_598), .B(n_624), .C(n_617), .Y(n_658) );
OAI211xp5_ASAP7_75t_SL g659 ( .A1(n_648), .A2(n_627), .B(n_623), .C(n_629), .Y(n_659) );
AOI22xp5_ASAP7_75t_L g660 ( .A1(n_653), .A2(n_628), .B1(n_627), .B2(n_620), .Y(n_660) );
AOI221xp5_ASAP7_75t_SL g661 ( .A1(n_638), .A2(n_630), .B1(n_610), .B2(n_618), .C(n_621), .Y(n_661) );
INVx1_ASAP7_75t_SL g662 ( .A(n_634), .Y(n_662) );
AOI21xp5_ASAP7_75t_L g663 ( .A1(n_638), .A2(n_601), .B(n_595), .Y(n_663) );
INVx1_ASAP7_75t_SL g664 ( .A(n_635), .Y(n_664) );
OAI221xp5_ASAP7_75t_L g665 ( .A1(n_645), .A2(n_595), .B1(n_622), .B2(n_631), .C(n_550), .Y(n_665) );
A2O1A1Ixp33_ASAP7_75t_L g666 ( .A1(n_647), .A2(n_489), .B(n_554), .C(n_560), .Y(n_666) );
NAND3xp33_ASAP7_75t_SL g667 ( .A(n_652), .B(n_495), .C(n_497), .Y(n_667) );
AOI322xp5_ASAP7_75t_L g668 ( .A1(n_637), .A2(n_589), .A3(n_587), .B1(n_583), .B2(n_522), .C1(n_523), .C2(n_532), .Y(n_668) );
AOI22xp5_ASAP7_75t_L g669 ( .A1(n_639), .A2(n_568), .B1(n_513), .B2(n_559), .Y(n_669) );
AOI221xp5_ASAP7_75t_L g670 ( .A1(n_661), .A2(n_650), .B1(n_642), .B2(n_640), .C(n_655), .Y(n_670) );
INVx1_ASAP7_75t_L g671 ( .A(n_657), .Y(n_671) );
OAI22x1_ASAP7_75t_L g672 ( .A1(n_660), .A2(n_652), .B1(n_655), .B2(n_643), .Y(n_672) );
OA22x2_ASAP7_75t_L g673 ( .A1(n_669), .A2(n_654), .B1(n_644), .B2(n_643), .Y(n_673) );
NAND2xp5_ASAP7_75t_SL g674 ( .A(n_663), .B(n_513), .Y(n_674) );
OAI32xp33_ASAP7_75t_L g675 ( .A1(n_659), .A2(n_633), .A3(n_646), .B1(n_649), .B2(n_644), .Y(n_675) );
OAI22xp33_ASAP7_75t_L g676 ( .A1(n_656), .A2(n_633), .B1(n_654), .B2(n_513), .Y(n_676) );
NAND2xp33_ASAP7_75t_SL g677 ( .A(n_667), .B(n_636), .Y(n_677) );
NAND2xp5_ASAP7_75t_L g678 ( .A(n_670), .B(n_668), .Y(n_678) );
OAI211xp5_ASAP7_75t_SL g679 ( .A1(n_674), .A2(n_665), .B(n_664), .C(n_662), .Y(n_679) );
NAND2xp5_ASAP7_75t_SL g680 ( .A(n_677), .B(n_666), .Y(n_680) );
AOI22xp33_ASAP7_75t_L g681 ( .A1(n_673), .A2(n_658), .B1(n_667), .B2(n_559), .Y(n_681) );
NAND2xp5_ASAP7_75t_SL g682 ( .A(n_676), .B(n_636), .Y(n_682) );
NOR5xp2_ASAP7_75t_L g683 ( .A(n_679), .B(n_675), .C(n_672), .D(n_671), .E(n_522), .Y(n_683) );
AND2x4_ASAP7_75t_L g684 ( .A(n_682), .B(n_554), .Y(n_684) );
NAND2xp5_ASAP7_75t_SL g685 ( .A(n_681), .B(n_489), .Y(n_685) );
AOI22xp33_ASAP7_75t_L g686 ( .A1(n_685), .A2(n_680), .B1(n_678), .B2(n_559), .Y(n_686) );
NAND3xp33_ASAP7_75t_L g687 ( .A(n_683), .B(n_534), .C(n_532), .Y(n_687) );
AOI22x1_ASAP7_75t_L g688 ( .A1(n_686), .A2(n_684), .B1(n_425), .B2(n_419), .Y(n_688) );
INVx2_ASAP7_75t_L g689 ( .A(n_687), .Y(n_689) );
AOI22xp5_ASAP7_75t_L g690 ( .A1(n_689), .A2(n_471), .B1(n_419), .B2(n_425), .Y(n_690) );
AOI222xp33_ASAP7_75t_SL g691 ( .A1(n_690), .A2(n_688), .B1(n_425), .B2(n_419), .C1(n_573), .C2(n_577), .Y(n_691) );
AOI222xp33_ASAP7_75t_L g692 ( .A1(n_691), .A2(n_425), .B1(n_487), .B2(n_486), .C1(n_484), .C2(n_483), .Y(n_692) );
OR2x2_ASAP7_75t_L g693 ( .A(n_692), .B(n_560), .Y(n_693) );
AOI22xp5_ASAP7_75t_L g694 ( .A1(n_693), .A2(n_425), .B1(n_471), .B2(n_495), .Y(n_694) );
endmodule