module fake_jpeg_20234_n_237 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_237);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_237;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_233;
wire n_102;
wire n_121;
wire n_130;
wire n_99;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx3_ASAP7_75t_L g15 ( 
.A(n_1),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_13),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

INVx6_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

BUFx12_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

INVx5_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_2),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_0),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_9),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_22),
.Y(n_33)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_33),
.Y(n_56)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_22),
.Y(n_34)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_34),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_19),
.B(n_0),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_SL g54 ( 
.A(n_35),
.B(n_37),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_22),
.Y(n_36)
);

BUFx2_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g37 ( 
.A(n_24),
.B(n_0),
.Y(n_37)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_19),
.Y(n_38)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g39 ( 
.A(n_16),
.B(n_1),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_39),
.B(n_42),
.Y(n_60)
);

INVx11_ASAP7_75t_L g40 ( 
.A(n_19),
.Y(n_40)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_40),
.Y(n_61)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_23),
.Y(n_41)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_41),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_16),
.B(n_1),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_43),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_32),
.Y(n_44)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_44),
.Y(n_52)
);

INVx5_ASAP7_75t_L g45 ( 
.A(n_15),
.Y(n_45)
);

INVx11_ASAP7_75t_L g65 ( 
.A(n_45),
.Y(n_65)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_32),
.Y(n_46)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_46),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g47 ( 
.A1(n_34),
.A2(n_18),
.B1(n_15),
.B2(n_20),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_47),
.A2(n_53),
.B1(n_67),
.B2(n_71),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_34),
.A2(n_18),
.B1(n_20),
.B2(n_15),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_48),
.A2(n_59),
.B1(n_29),
.B2(n_23),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_45),
.A2(n_18),
.B1(n_20),
.B2(n_31),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_39),
.B(n_31),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_55),
.B(n_68),
.Y(n_87)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_58),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_41),
.A2(n_30),
.B1(n_28),
.B2(n_25),
.Y(n_59)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_46),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_63),
.B(n_64),
.Y(n_81)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_33),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_35),
.B(n_30),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_66),
.B(n_69),
.Y(n_92)
);

OAI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_45),
.A2(n_28),
.B1(n_17),
.B2(n_27),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_37),
.B(n_27),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_37),
.B(n_25),
.Y(n_69)
);

A2O1A1Ixp33_ASAP7_75t_L g70 ( 
.A1(n_38),
.A2(n_21),
.B(n_17),
.C(n_19),
.Y(n_70)
);

A2O1A1Ixp33_ASAP7_75t_L g95 ( 
.A1(n_70),
.A2(n_3),
.B(n_6),
.C(n_7),
.Y(n_95)
);

OAI22xp33_ASAP7_75t_L g71 ( 
.A1(n_33),
.A2(n_19),
.B1(n_26),
.B2(n_24),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_40),
.B(n_21),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_72),
.B(n_73),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_40),
.B(n_14),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_41),
.B(n_26),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_74),
.B(n_76),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_36),
.B(n_26),
.Y(n_76)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_36),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_77),
.B(n_78),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_36),
.B(n_24),
.Y(n_78)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_36),
.Y(n_79)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_79),
.Y(n_91)
);

AO22x1_ASAP7_75t_SL g80 ( 
.A1(n_43),
.A2(n_23),
.B1(n_29),
.B2(n_4),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_80),
.A2(n_13),
.B1(n_7),
.B2(n_8),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_L g82 ( 
.A1(n_56),
.A2(n_44),
.B1(n_43),
.B2(n_46),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_82),
.A2(n_88),
.B1(n_96),
.B2(n_52),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_60),
.B(n_44),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_83),
.B(n_85),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_60),
.B(n_46),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_86),
.Y(n_129)
);

OAI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_70),
.A2(n_46),
.B1(n_29),
.B2(n_4),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_65),
.A2(n_2),
.B1(n_3),
.B2(n_5),
.Y(n_89)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_89),
.Y(n_131)
);

AOI21xp33_ASAP7_75t_L g90 ( 
.A1(n_54),
.A2(n_3),
.B(n_5),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g115 ( 
.A(n_90),
.B(n_107),
.Y(n_115)
);

BUFx2_ASAP7_75t_L g93 ( 
.A(n_49),
.Y(n_93)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_93),
.Y(n_132)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_71),
.Y(n_94)
);

INVx1_ASAP7_75t_SL g119 ( 
.A(n_94),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_95),
.B(n_97),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_58),
.B(n_6),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_54),
.B(n_6),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_100),
.B(n_102),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g101 ( 
.A(n_47),
.B(n_9),
.Y(n_101)
);

AO21x1_ASAP7_75t_L g125 ( 
.A1(n_101),
.A2(n_104),
.B(n_50),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_80),
.B(n_11),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_53),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_103),
.B(n_52),
.Y(n_113)
);

OA22x2_ASAP7_75t_L g104 ( 
.A1(n_56),
.A2(n_11),
.B1(n_12),
.B2(n_75),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_51),
.B(n_12),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_105),
.B(n_64),
.Y(n_126)
);

CKINVDCx16_ASAP7_75t_R g106 ( 
.A(n_51),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_106),
.B(n_62),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_80),
.B(n_12),
.Y(n_107)
);

AND2x2_ASAP7_75t_L g143 ( 
.A(n_110),
.B(n_113),
.Y(n_143)
);

NAND2x1_ASAP7_75t_L g111 ( 
.A(n_95),
.B(n_75),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_SL g149 ( 
.A1(n_111),
.A2(n_114),
.B(n_130),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_112),
.A2(n_127),
.B1(n_119),
.B2(n_96),
.Y(n_157)
);

NAND2x1_ASAP7_75t_SL g114 ( 
.A(n_104),
.B(n_49),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_98),
.B(n_57),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g156 ( 
.A(n_116),
.B(n_118),
.Y(n_156)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_91),
.Y(n_117)
);

INVxp67_ASAP7_75t_SL g158 ( 
.A(n_117),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_98),
.B(n_57),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_84),
.B(n_62),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_121),
.B(n_106),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_93),
.Y(n_123)
);

INVx2_ASAP7_75t_SL g159 ( 
.A(n_123),
.Y(n_159)
);

XOR2xp5_ASAP7_75t_L g124 ( 
.A(n_85),
.B(n_65),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_124),
.B(n_134),
.C(n_105),
.Y(n_150)
);

AO22x1_ASAP7_75t_L g140 ( 
.A1(n_125),
.A2(n_102),
.B1(n_104),
.B2(n_101),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_126),
.B(n_128),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_109),
.A2(n_63),
.B1(n_77),
.B2(n_79),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_87),
.B(n_50),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_84),
.A2(n_61),
.B1(n_104),
.B2(n_91),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_87),
.B(n_61),
.Y(n_133)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_133),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_83),
.B(n_99),
.C(n_108),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_99),
.B(n_92),
.Y(n_135)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_135),
.Y(n_144)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_81),
.Y(n_137)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_137),
.Y(n_145)
);

INVx5_ASAP7_75t_L g138 ( 
.A(n_93),
.Y(n_138)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_138),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_140),
.B(n_148),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_141),
.B(n_151),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g142 ( 
.A(n_124),
.B(n_100),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_142),
.B(n_150),
.C(n_152),
.Y(n_168)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_110),
.Y(n_147)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_147),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_134),
.A2(n_109),
.B1(n_107),
.B2(n_101),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_132),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g152 ( 
.A(n_120),
.B(n_97),
.Y(n_152)
);

NOR3xp33_ASAP7_75t_L g153 ( 
.A(n_111),
.B(n_92),
.C(n_108),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_153),
.B(n_115),
.Y(n_174)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_132),
.Y(n_154)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_154),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_157),
.B(n_160),
.Y(n_166)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_123),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_123),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_161),
.B(n_162),
.Y(n_170)
);

NOR2x1_ASAP7_75t_L g162 ( 
.A(n_111),
.B(n_104),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_121),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_163),
.B(n_126),
.Y(n_169)
);

AOI322xp5_ASAP7_75t_SL g164 ( 
.A1(n_144),
.A2(n_115),
.A3(n_136),
.B1(n_112),
.B2(n_122),
.C1(n_131),
.C2(n_137),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_SL g182 ( 
.A(n_164),
.B(n_148),
.Y(n_182)
);

O2A1O1Ixp33_ASAP7_75t_R g165 ( 
.A1(n_162),
.A2(n_114),
.B(n_125),
.C(n_122),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_165),
.B(n_174),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_169),
.B(n_173),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_150),
.B(n_120),
.C(n_127),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_156),
.B(n_117),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_176),
.B(n_177),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_145),
.B(n_139),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_L g178 ( 
.A1(n_149),
.A2(n_136),
.B(n_129),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_L g194 ( 
.A1(n_178),
.A2(n_143),
.B(n_155),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_152),
.B(n_125),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_179),
.B(n_180),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_142),
.B(n_81),
.C(n_114),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_149),
.B(n_138),
.C(n_129),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_181),
.B(n_143),
.Y(n_193)
);

AOI321xp33_ASAP7_75t_L g202 ( 
.A1(n_182),
.A2(n_194),
.A3(n_184),
.B1(n_188),
.B2(n_186),
.C(n_187),
.Y(n_202)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_175),
.Y(n_183)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_183),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_166),
.A2(n_157),
.B1(n_163),
.B2(n_131),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_185),
.B(n_189),
.Y(n_205)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_171),
.Y(n_187)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_187),
.Y(n_208)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_172),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_165),
.A2(n_167),
.B1(n_179),
.B2(n_170),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_190),
.A2(n_195),
.B1(n_140),
.B2(n_178),
.Y(n_201)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_169),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_191),
.Y(n_199)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_193),
.B(n_194),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_167),
.A2(n_147),
.B1(n_143),
.B2(n_140),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_173),
.B(n_141),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_196),
.B(n_168),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_197),
.B(n_201),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_186),
.B(n_168),
.C(n_180),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_200),
.B(n_204),
.C(n_183),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_SL g211 ( 
.A(n_202),
.B(n_206),
.Y(n_211)
);

CKINVDCx16_ASAP7_75t_R g203 ( 
.A(n_192),
.Y(n_203)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_203),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_188),
.B(n_181),
.Y(n_204)
);

OA21x2_ASAP7_75t_SL g206 ( 
.A1(n_195),
.A2(n_158),
.B(n_119),
.Y(n_206)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_207),
.Y(n_209)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_209),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_205),
.A2(n_185),
.B1(n_190),
.B2(n_189),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_213),
.B(n_215),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_214),
.B(n_204),
.Y(n_223)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_207),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_200),
.B(n_146),
.C(n_159),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_216),
.B(n_201),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_SL g217 ( 
.A1(n_205),
.A2(n_146),
.B(n_159),
.Y(n_217)
);

AOI21xp5_ASAP7_75t_L g222 ( 
.A1(n_217),
.A2(n_208),
.B(n_199),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_219),
.B(n_222),
.C(n_217),
.Y(n_227)
);

INVx11_ASAP7_75t_L g221 ( 
.A(n_210),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_221),
.A2(n_224),
.B1(n_208),
.B2(n_209),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_223),
.B(n_198),
.C(n_212),
.Y(n_228)
);

NOR2x1_ASAP7_75t_L g224 ( 
.A(n_211),
.B(n_199),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_225),
.B(n_226),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_218),
.A2(n_216),
.B1(n_214),
.B2(n_202),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_227),
.B(n_228),
.Y(n_231)
);

AOI21xp33_ASAP7_75t_L g229 ( 
.A1(n_224),
.A2(n_198),
.B(n_159),
.Y(n_229)
);

A2O1A1Ixp33_ASAP7_75t_SL g232 ( 
.A1(n_229),
.A2(n_222),
.B(n_221),
.C(n_218),
.Y(n_232)
);

BUFx24_ASAP7_75t_SL g234 ( 
.A(n_232),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_231),
.B(n_220),
.Y(n_233)
);

AOI21xp5_ASAP7_75t_L g236 ( 
.A1(n_233),
.A2(n_230),
.B(n_219),
.Y(n_236)
);

FAx1_ASAP7_75t_SL g235 ( 
.A(n_234),
.B(n_223),
.CI(n_227),
.CON(n_235),
.SN(n_235)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_235),
.B(n_236),
.Y(n_237)
);


endmodule