module real_jpeg_7908_n_16 (n_333, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_334, n_7, n_3, n_10, n_9, n_16);

input n_333;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_334;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_216;
wire n_128;
wire n_202;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_288;
wire n_83;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_330;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_299;
wire n_243;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx24_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

BUFx12_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

BUFx10_ASAP7_75t_L g111 ( 
.A(n_2),
.Y(n_111)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_3),
.Y(n_62)
);

BUFx10_ASAP7_75t_L g57 ( 
.A(n_4),
.Y(n_57)
);

BUFx6f_ASAP7_75t_SL g43 ( 
.A(n_5),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_6),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g35 ( 
.A1(n_7),
.A2(n_24),
.B1(n_33),
.B2(n_36),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_7),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_7),
.A2(n_29),
.B1(n_30),
.B2(n_36),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_7),
.A2(n_36),
.B1(n_60),
.B2(n_61),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_7),
.A2(n_36),
.B1(n_44),
.B2(n_46),
.Y(n_259)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_8),
.A2(n_60),
.B1(n_61),
.B2(n_109),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_8),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_8),
.A2(n_44),
.B1(n_46),
.B2(n_109),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_SL g179 ( 
.A1(n_8),
.A2(n_29),
.B1(n_30),
.B2(n_109),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_SL g234 ( 
.A1(n_8),
.A2(n_24),
.B1(n_33),
.B2(n_109),
.Y(n_234)
);

AOI21xp5_ASAP7_75t_L g118 ( 
.A1(n_9),
.A2(n_46),
.B(n_119),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_9),
.B(n_46),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_9),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_9),
.A2(n_132),
.B1(n_133),
.B2(n_134),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_9),
.B(n_91),
.Y(n_185)
);

AOI21xp33_ASAP7_75t_L g205 ( 
.A1(n_9),
.A2(n_26),
.B(n_30),
.Y(n_205)
);

OAI22xp33_ASAP7_75t_SL g223 ( 
.A1(n_9),
.A2(n_24),
.B1(n_33),
.B2(n_130),
.Y(n_223)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_10),
.A2(n_60),
.B1(n_61),
.B2(n_114),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_10),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g157 ( 
.A1(n_10),
.A2(n_44),
.B1(n_46),
.B2(n_114),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_SL g221 ( 
.A1(n_10),
.A2(n_29),
.B1(n_30),
.B2(n_114),
.Y(n_221)
);

AOI22xp33_ASAP7_75t_SL g253 ( 
.A1(n_10),
.A2(n_24),
.B1(n_33),
.B2(n_114),
.Y(n_253)
);

BUFx10_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_L g47 ( 
.A1(n_12),
.A2(n_29),
.B1(n_30),
.B2(n_48),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_12),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_12),
.A2(n_44),
.B1(n_46),
.B2(n_48),
.Y(n_65)
);

OAI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_12),
.A2(n_48),
.B1(n_60),
.B2(n_61),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_12),
.A2(n_24),
.B1(n_33),
.B2(n_48),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_13),
.A2(n_44),
.B1(n_46),
.B2(n_121),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_13),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_13),
.A2(n_60),
.B1(n_61),
.B2(n_121),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_13),
.A2(n_29),
.B1(n_30),
.B2(n_121),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_L g225 ( 
.A1(n_13),
.A2(n_24),
.B1(n_33),
.B2(n_121),
.Y(n_225)
);

AOI22xp33_ASAP7_75t_SL g32 ( 
.A1(n_14),
.A2(n_24),
.B1(n_33),
.B2(n_34),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_14),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_SL g183 ( 
.A1(n_14),
.A2(n_34),
.B1(n_60),
.B2(n_61),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_14),
.A2(n_34),
.B1(n_44),
.B2(n_46),
.Y(n_240)
);

AOI22xp33_ASAP7_75t_SL g281 ( 
.A1(n_14),
.A2(n_29),
.B1(n_30),
.B2(n_34),
.Y(n_281)
);

AOI22xp33_ASAP7_75t_L g53 ( 
.A1(n_15),
.A2(n_29),
.B1(n_30),
.B2(n_54),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_15),
.Y(n_54)
);

OAI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_15),
.A2(n_24),
.B1(n_33),
.B2(n_54),
.Y(n_71)
);

OAI22xp33_ASAP7_75t_SL g169 ( 
.A1(n_15),
.A2(n_54),
.B1(n_60),
.B2(n_61),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_L g218 ( 
.A1(n_15),
.A2(n_44),
.B1(n_46),
.B2(n_54),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_97),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_SL g17 ( 
.A(n_18),
.B(n_95),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_82),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_19),
.B(n_82),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_69),
.C(n_73),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_SL g324 ( 
.A1(n_20),
.A2(n_21),
.B1(n_69),
.B2(n_318),
.Y(n_324)
);

CKINVDCx14_ASAP7_75t_R g20 ( 
.A(n_21),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_37),
.B1(n_38),
.B2(n_68),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_22),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g22 ( 
.A1(n_23),
.A2(n_28),
.B1(n_32),
.B2(n_35),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_23),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_23),
.A2(n_28),
.B1(n_225),
.B2(n_234),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_23),
.A2(n_28),
.B1(n_234),
.B2(n_253),
.Y(n_252)
);

OAI21xp5_ASAP7_75t_SL g277 ( 
.A1(n_23),
.A2(n_253),
.B(n_278),
.Y(n_277)
);

OAI21xp5_ASAP7_75t_SL g298 ( 
.A1(n_23),
.A2(n_90),
.B(n_299),
.Y(n_298)
);

A2O1A1Ixp33_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_25),
.B(n_27),
.C(n_28),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_24),
.B(n_25),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_24),
.Y(n_33)
);

A2O1A1Ixp33_ASAP7_75t_L g204 ( 
.A1(n_24),
.A2(n_25),
.B(n_130),
.C(n_205),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g28 ( 
.A1(n_25),
.A2(n_26),
.B1(n_29),
.B2(n_30),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_26),
.Y(n_25)
);

OAI21xp5_ASAP7_75t_L g69 ( 
.A1(n_28),
.A2(n_32),
.B(n_70),
.Y(n_69)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_28),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_30),
.Y(n_29)
);

O2A1O1Ixp33_ASAP7_75t_L g50 ( 
.A1(n_30),
.A2(n_41),
.B(n_42),
.C(n_51),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_30),
.B(n_42),
.Y(n_51)
);

HAxp5_ASAP7_75t_SL g159 ( 
.A(n_30),
.B(n_130),
.CON(n_159),
.SN(n_159)
);

BUFx10_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_35),
.Y(n_88)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_SL g38 ( 
.A1(n_39),
.A2(n_55),
.B1(n_66),
.B2(n_67),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_39),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_40),
.B(n_49),
.Y(n_39)
);

OAI21xp5_ASAP7_75t_SL g235 ( 
.A1(n_40),
.A2(n_76),
.B(n_221),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_41),
.B(n_47),
.Y(n_40)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_41),
.Y(n_81)
);

OAI21xp5_ASAP7_75t_L g85 ( 
.A1(n_41),
.A2(n_47),
.B(n_50),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_41),
.A2(n_50),
.B1(n_159),
.B2(n_160),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_41),
.A2(n_50),
.B1(n_78),
.B2(n_304),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_SL g41 ( 
.A1(n_42),
.A2(n_43),
.B1(n_44),
.B2(n_46),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_SL g165 ( 
.A(n_42),
.B(n_46),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_43),
.Y(n_42)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_44),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_44),
.A2(n_51),
.B1(n_159),
.B2(n_165),
.Y(n_164)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

A2O1A1Ixp33_ASAP7_75t_SL g56 ( 
.A1(n_46),
.A2(n_57),
.B(n_58),
.C(n_59),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_46),
.B(n_57),
.Y(n_58)
);

AOI21xp5_ASAP7_75t_L g255 ( 
.A1(n_47),
.A2(n_50),
.B(n_80),
.Y(n_255)
);

OAI21xp5_ASAP7_75t_L g280 ( 
.A1(n_49),
.A2(n_81),
.B(n_281),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_50),
.B(n_52),
.Y(n_49)
);

CKINVDCx16_ASAP7_75t_R g76 ( 
.A(n_50),
.Y(n_76)
);

INVxp67_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_53),
.B(n_81),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_55),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_55),
.B(n_66),
.C(n_68),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g320 ( 
.A1(n_55),
.A2(n_67),
.B1(n_74),
.B2(n_75),
.Y(n_320)
);

AOI21xp5_ASAP7_75t_SL g55 ( 
.A1(n_56),
.A2(n_59),
.B(n_64),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_56),
.A2(n_59),
.B1(n_118),
.B2(n_120),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_56),
.A2(n_59),
.B1(n_120),
.B2(n_147),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_56),
.A2(n_59),
.B1(n_147),
.B2(n_157),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_SL g192 ( 
.A1(n_56),
.A2(n_157),
.B(n_193),
.Y(n_192)
);

CKINVDCx16_ASAP7_75t_R g216 ( 
.A(n_56),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g258 ( 
.A1(n_56),
.A2(n_59),
.B1(n_240),
.B2(n_259),
.Y(n_258)
);

OAI21xp5_ASAP7_75t_SL g287 ( 
.A1(n_56),
.A2(n_259),
.B(n_288),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_57),
.A2(n_60),
.B1(n_61),
.B2(n_63),
.Y(n_59)
);

CKINVDCx16_ASAP7_75t_R g63 ( 
.A(n_57),
.Y(n_63)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_58),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g129 ( 
.A(n_59),
.B(n_130),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g194 ( 
.A(n_59),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_59),
.B(n_218),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_L g239 ( 
.A1(n_59),
.A2(n_240),
.B(n_241),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_60),
.B(n_111),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_60),
.B(n_63),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_60),
.B(n_138),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_61),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_61),
.A2(n_123),
.B1(n_124),
.B2(n_125),
.Y(n_122)
);

BUFx24_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVxp67_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_65),
.B(n_194),
.Y(n_193)
);

AOI21xp5_ASAP7_75t_L g215 ( 
.A1(n_65),
.A2(n_216),
.B(n_217),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_67),
.B(n_69),
.C(n_74),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_69),
.A2(n_318),
.B1(n_319),
.B2(n_320),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_69),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_71),
.B(n_72),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_71),
.B(n_91),
.Y(n_90)
);

AOI21xp5_ASAP7_75t_L g87 ( 
.A1(n_72),
.A2(n_88),
.B(n_89),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_72),
.A2(n_91),
.B1(n_223),
.B2(n_224),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g323 ( 
.A(n_73),
.B(n_324),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_75),
.Y(n_74)
);

OAI21xp5_ASAP7_75t_SL g75 ( 
.A1(n_76),
.A2(n_77),
.B(n_79),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_76),
.A2(n_81),
.B1(n_178),
.B2(n_179),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_76),
.A2(n_81),
.B1(n_179),
.B2(n_221),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_78),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_80),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_81),
.B(n_130),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_83),
.A2(n_92),
.B1(n_93),
.B2(n_94),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_83),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_84),
.A2(n_85),
.B1(n_86),
.B2(n_87),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_85),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_87),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_90),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_91),
.B(n_279),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_93),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

OAI321xp33_ASAP7_75t_L g97 ( 
.A1(n_98),
.A2(n_315),
.A3(n_325),
.B1(n_330),
.B2(n_331),
.C(n_333),
.Y(n_97)
);

AOI321xp33_ASAP7_75t_L g98 ( 
.A1(n_99),
.A2(n_267),
.A3(n_291),
.B1(n_308),
.B2(n_314),
.C(n_334),
.Y(n_98)
);

NOR3xp33_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_227),
.C(n_263),
.Y(n_99)
);

AOI21xp5_ASAP7_75t_L g100 ( 
.A1(n_101),
.A2(n_198),
.B(n_226),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_SL g101 ( 
.A1(n_102),
.A2(n_172),
.B(n_197),
.Y(n_101)
);

AOI21xp5_ASAP7_75t_L g102 ( 
.A1(n_103),
.A2(n_152),
.B(n_171),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_SL g103 ( 
.A1(n_104),
.A2(n_141),
.B(n_151),
.Y(n_103)
);

AOI21xp5_ASAP7_75t_L g104 ( 
.A1(n_105),
.A2(n_127),
.B(n_140),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_106),
.B(n_115),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_106),
.B(n_115),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_107),
.A2(n_110),
.B1(n_111),
.B2(n_112),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_108),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_108),
.A2(n_132),
.B1(n_133),
.B2(n_134),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_110),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_110),
.B(n_169),
.Y(n_184)
);

CKINVDCx16_ASAP7_75t_R g134 ( 
.A(n_111),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_111),
.B(n_150),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_111),
.B(n_169),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_113),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_L g148 ( 
.A1(n_113),
.A2(n_133),
.B(n_149),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_116),
.A2(n_117),
.B1(n_122),
.B2(n_126),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g142 ( 
.A(n_116),
.B(n_126),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_117),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_119),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_122),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_SL g127 ( 
.A1(n_128),
.A2(n_135),
.B(n_139),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_131),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_129),
.B(n_131),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_130),
.B(n_134),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_SL g166 ( 
.A1(n_133),
.A2(n_167),
.B(n_168),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_133),
.A2(n_134),
.B1(n_183),
.B2(n_208),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_SL g243 ( 
.A1(n_133),
.A2(n_168),
.B(n_208),
.Y(n_243)
);

AOI21xp5_ASAP7_75t_L g286 ( 
.A1(n_133),
.A2(n_134),
.B(n_167),
.Y(n_286)
);

OAI21xp5_ASAP7_75t_L g182 ( 
.A1(n_134),
.A2(n_183),
.B(n_184),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_136),
.B(n_137),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_143),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_142),
.B(n_143),
.Y(n_151)
);

CKINVDCx5p33_ASAP7_75t_R g143 ( 
.A(n_144),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_144),
.B(n_153),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g171 ( 
.A(n_144),
.B(n_153),
.Y(n_171)
);

FAx1_ASAP7_75t_SL g144 ( 
.A(n_145),
.B(n_146),
.CI(n_148),
.CON(n_144),
.SN(n_144)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_149),
.B(n_184),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_150),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_154),
.A2(n_155),
.B1(n_163),
.B2(n_170),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_156),
.A2(n_158),
.B1(n_161),
.B2(n_162),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_156),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_158),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_158),
.B(n_162),
.C(n_170),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_160),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_163),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_166),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_164),
.B(n_166),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_173),
.B(n_174),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_173),
.B(n_174),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_175),
.A2(n_176),
.B1(n_189),
.B2(n_190),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_175),
.B(n_192),
.C(n_195),
.Y(n_199)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_177),
.A2(n_180),
.B1(n_181),
.B2(n_188),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_177),
.Y(n_188)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_182),
.A2(n_185),
.B1(n_186),
.B2(n_187),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_182),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_185),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_185),
.B(n_186),
.C(n_188),
.Y(n_209)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_191),
.A2(n_192),
.B1(n_195),
.B2(n_196),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_191),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_192),
.Y(n_196)
);

AND2x2_ASAP7_75t_L g305 ( 
.A(n_193),
.B(n_241),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_200),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_SL g226 ( 
.A(n_199),
.B(n_200),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_212),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_202),
.A2(n_209),
.B1(n_210),
.B2(n_211),
.Y(n_201)
);

CKINVDCx16_ASAP7_75t_R g210 ( 
.A(n_202),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_202),
.B(n_211),
.C(n_212),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_203),
.A2(n_204),
.B1(n_206),
.B2(n_207),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_203),
.B(n_207),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_204),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_207),
.Y(n_206)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_209),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_222),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_214),
.A2(n_215),
.B1(n_219),
.B2(n_220),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_215),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_215),
.B(n_219),
.C(n_222),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_216),
.B(n_242),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_217),
.Y(n_288)
);

INVxp67_ASAP7_75t_L g242 ( 
.A(n_218),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_220),
.Y(n_219)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_227),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_246),
.Y(n_227)
);

AND2x2_ASAP7_75t_L g312 ( 
.A(n_228),
.B(n_246),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_237),
.C(n_244),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_229),
.B(n_266),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_231),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_230),
.B(n_232),
.C(n_236),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_232),
.A2(n_233),
.B1(n_235),
.B2(n_236),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_233),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_235),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_237),
.A2(n_238),
.B1(n_244),
.B2(n_245),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_238),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_243),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_239),
.B(n_243),
.Y(n_249)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_247),
.A2(n_260),
.B1(n_261),
.B2(n_262),
.Y(n_246)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_247),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_256),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_248),
.B(n_256),
.C(n_260),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_250),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_249),
.B(n_251),
.C(n_255),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_251),
.A2(n_252),
.B1(n_254),
.B2(n_255),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_252),
.Y(n_251)
);

CKINVDCx14_ASAP7_75t_R g254 ( 
.A(n_255),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_257),
.B(n_258),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_257),
.B(n_258),
.Y(n_274)
);

CKINVDCx14_ASAP7_75t_R g260 ( 
.A(n_261),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_264),
.B(n_265),
.Y(n_263)
);

AND2x2_ASAP7_75t_L g311 ( 
.A(n_264),
.B(n_265),
.Y(n_311)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

OAI21xp5_ASAP7_75t_SL g308 ( 
.A1(n_268),
.A2(n_309),
.B(n_313),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_270),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_SL g313 ( 
.A(n_269),
.B(n_270),
.Y(n_313)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_271),
.B(n_290),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_272),
.A2(n_273),
.B1(n_283),
.B2(n_284),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_272),
.B(n_284),
.C(n_290),
.Y(n_292)
);

CKINVDCx14_ASAP7_75t_R g272 ( 
.A(n_273),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_274),
.B(n_275),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_274),
.B(n_276),
.C(n_282),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_L g275 ( 
.A1(n_276),
.A2(n_277),
.B1(n_280),
.B2(n_282),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_277),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_279),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_280),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_281),
.Y(n_304)
);

CKINVDCx16_ASAP7_75t_R g283 ( 
.A(n_284),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_L g284 ( 
.A1(n_285),
.A2(n_286),
.B1(n_287),
.B2(n_289),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_285),
.A2(n_286),
.B1(n_297),
.B2(n_298),
.Y(n_296)
);

OAI21xp5_ASAP7_75t_L g322 ( 
.A1(n_285),
.A2(n_298),
.B(n_301),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_286),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_286),
.B(n_287),
.Y(n_300)
);

CKINVDCx14_ASAP7_75t_R g289 ( 
.A(n_287),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_292),
.B(n_293),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_SL g314 ( 
.A(n_292),
.B(n_293),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_293),
.Y(n_326)
);

FAx1_ASAP7_75t_SL g293 ( 
.A(n_294),
.B(n_302),
.CI(n_307),
.CON(n_293),
.SN(n_293)
);

OAI22xp5_ASAP7_75t_L g294 ( 
.A1(n_295),
.A2(n_296),
.B1(n_300),
.B2(n_301),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_298),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_300),
.Y(n_301)
);

OAI21xp5_ASAP7_75t_L g302 ( 
.A1(n_303),
.A2(n_305),
.B(n_306),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_303),
.B(n_305),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_306),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_SL g328 ( 
.A1(n_306),
.A2(n_317),
.B1(n_321),
.B2(n_329),
.Y(n_328)
);

AOI21xp5_ASAP7_75t_L g309 ( 
.A1(n_310),
.A2(n_311),
.B(n_312),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_316),
.B(n_323),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_316),
.B(n_323),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_317),
.B(n_321),
.C(n_322),
.Y(n_316)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_317),
.Y(n_329)
);

CKINVDCx14_ASAP7_75t_R g319 ( 
.A(n_320),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_L g327 ( 
.A(n_322),
.B(n_328),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_326),
.B(n_327),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_SL g330 ( 
.A(n_326),
.B(n_327),
.Y(n_330)
);


endmodule