module fake_jpeg_16628_n_373 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_373);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_373;

wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_327;
wire n_122;
wire n_75;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx3_ASAP7_75t_L g14 ( 
.A(n_10),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_8),
.Y(n_15)
);

BUFx4f_ASAP7_75t_SL g16 ( 
.A(n_12),
.Y(n_16)
);

BUFx24_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

INVx4_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_3),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_2),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_2),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_4),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

BUFx12_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

CKINVDCx14_ASAP7_75t_R g29 ( 
.A(n_2),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_13),
.Y(n_32)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_11),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_5),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_18),
.Y(n_37)
);

INVx5_ASAP7_75t_L g83 ( 
.A(n_37),
.Y(n_83)
);

BUFx12f_ASAP7_75t_SL g38 ( 
.A(n_17),
.Y(n_38)
);

OR2x2_ASAP7_75t_L g98 ( 
.A(n_38),
.B(n_26),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_39),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_31),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_40),
.B(n_43),
.Y(n_76)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_19),
.Y(n_41)
);

BUFx2_ASAP7_75t_SL g70 ( 
.A(n_41),
.Y(n_70)
);

BUFx10_ASAP7_75t_L g42 ( 
.A(n_16),
.Y(n_42)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_42),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_32),
.B(n_13),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_31),
.B(n_0),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_44),
.B(n_45),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_16),
.Y(n_45)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_46),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_32),
.B(n_12),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_47),
.B(n_51),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_18),
.Y(n_48)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_48),
.Y(n_79)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_23),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_49),
.Y(n_69)
);

INVx4_ASAP7_75t_SL g50 ( 
.A(n_16),
.Y(n_50)
);

INVx13_ASAP7_75t_L g84 ( 
.A(n_50),
.Y(n_84)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_14),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_14),
.Y(n_52)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_52),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_23),
.Y(n_53)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_53),
.Y(n_80)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_23),
.Y(n_54)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_54),
.Y(n_102)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_19),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_55),
.B(n_58),
.Y(n_74)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_28),
.Y(n_56)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_56),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_25),
.Y(n_57)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_57),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_16),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_34),
.Y(n_59)
);

HB1xp67_ASAP7_75t_L g72 ( 
.A(n_59),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_25),
.Y(n_60)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_60),
.Y(n_110)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_25),
.Y(n_61)
);

INVx8_ASAP7_75t_L g86 ( 
.A(n_61),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_26),
.B(n_0),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_62),
.B(n_64),
.Y(n_75)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_33),
.Y(n_63)
);

INVx11_ASAP7_75t_L g89 ( 
.A(n_63),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_28),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_28),
.Y(n_65)
);

HB1xp67_ASAP7_75t_L g113 ( 
.A(n_65),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_15),
.B(n_0),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_66),
.B(n_36),
.Y(n_77)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_59),
.Y(n_67)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_67),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_66),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_68),
.B(n_96),
.Y(n_127)
);

AOI21xp5_ASAP7_75t_L g71 ( 
.A1(n_38),
.A2(n_17),
.B(n_28),
.Y(n_71)
);

OAI21xp33_ASAP7_75t_L g125 ( 
.A1(n_71),
.A2(n_100),
.B(n_4),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_61),
.A2(n_46),
.B1(n_19),
.B2(n_33),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_73),
.A2(n_88),
.B1(n_92),
.B2(n_108),
.Y(n_118)
);

AND2x2_ASAP7_75t_L g141 ( 
.A(n_77),
.B(n_105),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_40),
.B(n_36),
.Y(n_81)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_81),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_50),
.A2(n_33),
.B1(n_29),
.B2(n_24),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_85),
.A2(n_87),
.B1(n_90),
.B2(n_91),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_51),
.A2(n_29),
.B1(n_2),
.B2(n_3),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_52),
.A2(n_30),
.B1(n_27),
.B2(n_15),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_L g90 ( 
.A1(n_63),
.A2(n_24),
.B1(n_20),
.B2(n_21),
.Y(n_90)
);

OAI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_56),
.A2(n_22),
.B1(n_20),
.B2(n_21),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_44),
.A2(n_57),
.B1(n_53),
.B2(n_60),
.Y(n_92)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_37),
.Y(n_94)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_94),
.Y(n_133)
);

INVx8_ASAP7_75t_L g95 ( 
.A(n_37),
.Y(n_95)
);

INVx4_ASAP7_75t_L g117 ( 
.A(n_95),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_65),
.Y(n_96)
);

INVx1_ASAP7_75t_SL g135 ( 
.A(n_98),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_45),
.B(n_22),
.Y(n_99)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_99),
.Y(n_136)
);

AND2x4_ASAP7_75t_SL g100 ( 
.A(n_42),
.B(n_35),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_58),
.B(n_26),
.Y(n_101)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_101),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_64),
.B(n_35),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_39),
.A2(n_17),
.B1(n_30),
.B2(n_27),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_106),
.A2(n_17),
.B1(n_41),
.B2(n_6),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_48),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_49),
.B(n_35),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_109),
.B(n_112),
.Y(n_140)
);

OR2x2_ASAP7_75t_L g112 ( 
.A(n_42),
.B(n_26),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_49),
.A2(n_30),
.B1(n_27),
.B2(n_35),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_114),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_147)
);

INVx11_ASAP7_75t_L g115 ( 
.A(n_54),
.Y(n_115)
);

INVx6_ASAP7_75t_L g120 ( 
.A(n_115),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_42),
.B(n_4),
.Y(n_116)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_116),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_82),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g203 ( 
.A(n_119),
.Y(n_203)
);

CKINVDCx14_ASAP7_75t_R g121 ( 
.A(n_71),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_121),
.B(n_124),
.Y(n_173)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_67),
.Y(n_122)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_122),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_123),
.A2(n_131),
.B1(n_147),
.B2(n_151),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_72),
.Y(n_124)
);

AND2x2_ASAP7_75t_L g179 ( 
.A(n_125),
.B(n_139),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_76),
.B(n_55),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_SL g201 ( 
.A(n_126),
.B(n_145),
.Y(n_201)
);

INVx6_ASAP7_75t_L g128 ( 
.A(n_82),
.Y(n_128)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_128),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_100),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_104),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_132),
.B(n_142),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_SL g134 ( 
.A(n_77),
.B(n_5),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_134),
.B(n_150),
.C(n_143),
.Y(n_176)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_94),
.Y(n_138)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_138),
.Y(n_193)
);

OA22x2_ASAP7_75t_SL g139 ( 
.A1(n_100),
.A2(n_54),
.B1(n_6),
.B2(n_7),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_70),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_107),
.B(n_5),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_143),
.B(n_152),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_111),
.B(n_7),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_111),
.B(n_7),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_SL g202 ( 
.A(n_146),
.B(n_162),
.Y(n_202)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_78),
.Y(n_148)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_148),
.Y(n_198)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_78),
.Y(n_149)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_149),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_105),
.B(n_8),
.C(n_10),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_100),
.A2(n_8),
.B1(n_11),
.B2(n_68),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_107),
.B(n_11),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_89),
.A2(n_11),
.B1(n_86),
.B2(n_110),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_153),
.A2(n_110),
.B1(n_80),
.B2(n_103),
.Y(n_187)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_104),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_155),
.B(n_157),
.Y(n_183)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_82),
.Y(n_156)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_156),
.Y(n_205)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_79),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_98),
.A2(n_108),
.B1(n_87),
.B2(n_88),
.Y(n_158)
);

OR2x2_ASAP7_75t_L g191 ( 
.A(n_158),
.B(n_89),
.Y(n_191)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_79),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_159),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g160 ( 
.A(n_80),
.Y(n_160)
);

BUFx3_ASAP7_75t_L g177 ( 
.A(n_160),
.Y(n_177)
);

BUFx2_ASAP7_75t_L g161 ( 
.A(n_113),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_161),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_74),
.Y(n_162)
);

INVx3_ASAP7_75t_L g163 ( 
.A(n_97),
.Y(n_163)
);

INVx13_ASAP7_75t_L g195 ( 
.A(n_163),
.Y(n_195)
);

CKINVDCx16_ASAP7_75t_R g164 ( 
.A(n_109),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_164),
.B(n_75),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_96),
.B(n_92),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_165),
.B(n_166),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_112),
.B(n_76),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_165),
.A2(n_73),
.B1(n_114),
.B2(n_86),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_169),
.A2(n_182),
.B1(n_190),
.B2(n_150),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_129),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_170),
.B(n_186),
.Y(n_219)
);

INVx2_ASAP7_75t_SL g171 ( 
.A(n_160),
.Y(n_171)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_171),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_176),
.B(n_134),
.Y(n_213)
);

INVxp67_ASAP7_75t_L g180 ( 
.A(n_138),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_180),
.B(n_69),
.Y(n_230)
);

AND2x6_ASAP7_75t_L g181 ( 
.A(n_125),
.B(n_98),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_181),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_158),
.A2(n_137),
.B1(n_118),
.B2(n_141),
.Y(n_182)
);

O2A1O1Ixp33_ASAP7_75t_L g184 ( 
.A1(n_139),
.A2(n_93),
.B(n_102),
.C(n_95),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_L g233 ( 
.A1(n_184),
.A2(n_187),
.B(n_191),
.Y(n_233)
);

AND2x2_ASAP7_75t_L g185 ( 
.A(n_140),
.B(n_112),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_SL g212 ( 
.A1(n_185),
.A2(n_197),
.B(n_210),
.Y(n_212)
);

BUFx5_ASAP7_75t_L g186 ( 
.A(n_117),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_118),
.A2(n_103),
.B1(n_97),
.B2(n_83),
.Y(n_190)
);

AND2x6_ASAP7_75t_L g192 ( 
.A(n_135),
.B(n_141),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_192),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_133),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_194),
.B(n_196),
.Y(n_220)
);

INVx6_ASAP7_75t_L g196 ( 
.A(n_119),
.Y(n_196)
);

AND2x2_ASAP7_75t_L g197 ( 
.A(n_140),
.B(n_84),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_SL g216 ( 
.A(n_199),
.B(n_206),
.Y(n_216)
);

INVx13_ASAP7_75t_L g200 ( 
.A(n_142),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_200),
.B(n_208),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_127),
.B(n_141),
.Y(n_206)
);

BUFx8_ASAP7_75t_L g207 ( 
.A(n_163),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_207),
.Y(n_235)
);

INVx13_ASAP7_75t_L g208 ( 
.A(n_161),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_152),
.B(n_115),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_SL g218 ( 
.A(n_209),
.B(n_154),
.Y(n_218)
);

AND2x6_ASAP7_75t_L g210 ( 
.A(n_135),
.B(n_84),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_213),
.B(n_228),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_182),
.A2(n_166),
.B1(n_139),
.B2(n_128),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_L g256 ( 
.A1(n_214),
.A2(n_217),
.B1(n_226),
.B2(n_242),
.Y(n_256)
);

INVxp67_ASAP7_75t_L g215 ( 
.A(n_175),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_215),
.B(n_218),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_172),
.A2(n_147),
.B1(n_122),
.B2(n_148),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_221),
.A2(n_234),
.B1(n_244),
.B2(n_241),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_189),
.B(n_149),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_222),
.B(n_227),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_191),
.A2(n_156),
.B1(n_144),
.B2(n_83),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_223),
.A2(n_245),
.B1(n_246),
.B2(n_247),
.Y(n_250)
);

AOI21xp5_ASAP7_75t_L g224 ( 
.A1(n_179),
.A2(n_117),
.B(n_120),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_SL g266 ( 
.A1(n_224),
.A2(n_238),
.B(n_240),
.Y(n_266)
);

CKINVDCx16_ASAP7_75t_R g225 ( 
.A(n_183),
.Y(n_225)
);

CKINVDCx14_ASAP7_75t_R g261 ( 
.A(n_225),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_189),
.A2(n_120),
.B1(n_102),
.B2(n_93),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_SL g227 ( 
.A(n_178),
.B(n_130),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_185),
.B(n_136),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_228),
.B(n_239),
.Y(n_263)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_198),
.Y(n_229)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_229),
.Y(n_268)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_230),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_202),
.B(n_84),
.Y(n_231)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_231),
.Y(n_251)
);

CKINVDCx16_ASAP7_75t_R g237 ( 
.A(n_198),
.Y(n_237)
);

INVx1_ASAP7_75t_SL g258 ( 
.A(n_237),
.Y(n_258)
);

OAI21xp5_ASAP7_75t_SL g238 ( 
.A1(n_179),
.A2(n_185),
.B(n_197),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_178),
.B(n_69),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_197),
.B(n_179),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_240),
.B(n_244),
.Y(n_279)
);

AOI21xp5_ASAP7_75t_SL g241 ( 
.A1(n_181),
.A2(n_173),
.B(n_184),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_L g252 ( 
.A1(n_241),
.A2(n_193),
.B(n_207),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_190),
.A2(n_169),
.B1(n_192),
.B2(n_210),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_201),
.B(n_167),
.Y(n_243)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_243),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_176),
.B(n_167),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_187),
.A2(n_180),
.B1(n_174),
.B2(n_204),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_204),
.A2(n_188),
.B1(n_168),
.B2(n_174),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_168),
.A2(n_171),
.B1(n_188),
.B2(n_205),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_200),
.B(n_207),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_248),
.B(n_213),
.C(n_212),
.Y(n_275)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_205),
.Y(n_249)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_249),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_252),
.A2(n_211),
.B1(n_216),
.B2(n_279),
.Y(n_306)
);

OAI21xp5_ASAP7_75t_SL g294 ( 
.A1(n_253),
.A2(n_266),
.B(n_281),
.Y(n_294)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_212),
.B(n_195),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_255),
.B(n_260),
.C(n_275),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_234),
.A2(n_171),
.B1(n_193),
.B2(n_196),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_L g300 ( 
.A1(n_257),
.A2(n_262),
.B1(n_265),
.B2(n_247),
.Y(n_300)
);

OAI22xp33_ASAP7_75t_SL g259 ( 
.A1(n_245),
.A2(n_195),
.B1(n_208),
.B2(n_177),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g291 ( 
.A(n_259),
.B(n_264),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_241),
.A2(n_232),
.B1(n_221),
.B2(n_217),
.Y(n_262)
);

OAI22xp33_ASAP7_75t_SL g264 ( 
.A1(n_223),
.A2(n_177),
.B1(n_186),
.B2(n_203),
.Y(n_264)
);

OA22x2_ASAP7_75t_L g265 ( 
.A1(n_233),
.A2(n_203),
.B1(n_224),
.B2(n_226),
.Y(n_265)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_249),
.Y(n_269)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_269),
.Y(n_289)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_220),
.Y(n_273)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_273),
.Y(n_290)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_229),
.Y(n_274)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_274),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_232),
.B(n_238),
.C(n_222),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_276),
.B(n_243),
.Y(n_283)
);

INVxp67_ASAP7_75t_L g277 ( 
.A(n_236),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_277),
.B(n_280),
.Y(n_284)
);

FAx1_ASAP7_75t_SL g278 ( 
.A(n_214),
.B(n_233),
.CI(n_242),
.CON(n_278),
.SN(n_278)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_278),
.B(n_262),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_219),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_L g281 ( 
.A1(n_239),
.A2(n_231),
.B(n_218),
.Y(n_281)
);

AOI21xp5_ASAP7_75t_L g282 ( 
.A1(n_266),
.A2(n_248),
.B(n_235),
.Y(n_282)
);

OAI21xp5_ASAP7_75t_SL g311 ( 
.A1(n_282),
.A2(n_285),
.B(n_295),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_283),
.B(n_288),
.C(n_260),
.Y(n_316)
);

XNOR2x2_ASAP7_75t_L g285 ( 
.A(n_252),
.B(n_278),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_261),
.B(n_225),
.Y(n_286)
);

CKINVDCx14_ASAP7_75t_R g317 ( 
.A(n_286),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_268),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_287),
.B(n_296),
.Y(n_324)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_275),
.B(n_216),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_268),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_269),
.Y(n_297)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_297),
.Y(n_308)
);

INVxp67_ASAP7_75t_L g298 ( 
.A(n_257),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_298),
.B(n_299),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_254),
.B(n_227),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_300),
.A2(n_265),
.B1(n_263),
.B2(n_279),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_271),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_L g312 ( 
.A1(n_301),
.A2(n_303),
.B1(n_304),
.B2(n_258),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_270),
.B(n_246),
.Y(n_302)
);

INVxp67_ASAP7_75t_L g326 ( 
.A(n_302),
.Y(n_326)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_272),
.Y(n_303)
);

AOI21xp5_ASAP7_75t_L g304 ( 
.A1(n_255),
.A2(n_235),
.B(n_230),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_251),
.B(n_237),
.Y(n_305)
);

NAND3xp33_ASAP7_75t_L g310 ( 
.A(n_305),
.B(n_307),
.C(n_254),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_306),
.B(n_263),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_272),
.B(n_211),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_L g331 ( 
.A1(n_309),
.A2(n_313),
.B1(n_318),
.B2(n_322),
.Y(n_331)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_310),
.Y(n_328)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_312),
.Y(n_338)
);

OAI22xp5_ASAP7_75t_L g313 ( 
.A1(n_302),
.A2(n_253),
.B1(n_276),
.B2(n_256),
.Y(n_313)
);

AOI22x1_ASAP7_75t_L g314 ( 
.A1(n_285),
.A2(n_265),
.B1(n_250),
.B2(n_278),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_SL g342 ( 
.A1(n_314),
.A2(n_320),
.B1(n_318),
.B2(n_325),
.Y(n_342)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_316),
.B(n_321),
.C(n_323),
.Y(n_341)
);

AOI322xp5_ASAP7_75t_L g319 ( 
.A1(n_300),
.A2(n_281),
.A3(n_265),
.B1(n_267),
.B2(n_250),
.C1(n_277),
.C2(n_258),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_319),
.B(n_314),
.Y(n_343)
);

OAI22xp5_ASAP7_75t_SL g320 ( 
.A1(n_295),
.A2(n_304),
.B1(n_285),
.B2(n_294),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_292),
.B(n_288),
.C(n_283),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_L g322 ( 
.A1(n_291),
.A2(n_284),
.B1(n_305),
.B2(n_303),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_292),
.B(n_282),
.C(n_294),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_306),
.B(n_299),
.C(n_307),
.Y(n_325)
);

XNOR2xp5_ASAP7_75t_L g332 ( 
.A(n_325),
.B(n_327),
.Y(n_332)
);

XNOR2xp5_ASAP7_75t_L g327 ( 
.A(n_284),
.B(n_286),
.Y(n_327)
);

AOI21xp5_ASAP7_75t_SL g329 ( 
.A1(n_311),
.A2(n_291),
.B(n_287),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_L g352 ( 
.A1(n_329),
.A2(n_328),
.B1(n_331),
.B2(n_335),
.Y(n_352)
);

CKINVDCx20_ASAP7_75t_R g330 ( 
.A(n_324),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_330),
.B(n_339),
.Y(n_348)
);

AOI21xp5_ASAP7_75t_L g333 ( 
.A1(n_311),
.A2(n_296),
.B(n_301),
.Y(n_333)
);

OAI22xp5_ASAP7_75t_SL g350 ( 
.A1(n_333),
.A2(n_321),
.B1(n_338),
.B2(n_334),
.Y(n_350)
);

AOI22xp5_ASAP7_75t_L g334 ( 
.A1(n_326),
.A2(n_289),
.B1(n_297),
.B2(n_293),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_L g344 ( 
.A1(n_334),
.A2(n_317),
.B1(n_309),
.B2(n_323),
.Y(n_344)
);

OAI21xp33_ASAP7_75t_L g335 ( 
.A1(n_315),
.A2(n_293),
.B(n_289),
.Y(n_335)
);

AOI21xp5_ASAP7_75t_L g347 ( 
.A1(n_335),
.A2(n_340),
.B(n_316),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_SL g336 ( 
.A(n_327),
.B(n_290),
.Y(n_336)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_336),
.Y(n_351)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_308),
.Y(n_337)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_337),
.Y(n_353)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_315),
.Y(n_339)
);

OAI21xp5_ASAP7_75t_L g340 ( 
.A1(n_326),
.A2(n_290),
.B(n_314),
.Y(n_340)
);

XNOR2xp5_ASAP7_75t_L g345 ( 
.A(n_342),
.B(n_343),
.Y(n_345)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_344),
.Y(n_357)
);

XNOR2xp5_ASAP7_75t_L g346 ( 
.A(n_332),
.B(n_320),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g355 ( 
.A(n_346),
.B(n_354),
.C(n_341),
.Y(n_355)
);

XNOR2xp5_ASAP7_75t_L g358 ( 
.A(n_347),
.B(n_350),
.Y(n_358)
);

OA21x2_ASAP7_75t_L g349 ( 
.A1(n_329),
.A2(n_333),
.B(n_340),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_L g360 ( 
.A(n_349),
.B(n_352),
.Y(n_360)
);

AOI21xp5_ASAP7_75t_L g359 ( 
.A1(n_352),
.A2(n_337),
.B(n_349),
.Y(n_359)
);

XNOR2xp5_ASAP7_75t_L g354 ( 
.A(n_332),
.B(n_341),
.Y(n_354)
);

XOR2xp5_ASAP7_75t_L g362 ( 
.A(n_355),
.B(n_359),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_SL g356 ( 
.A(n_351),
.B(n_342),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_356),
.B(n_350),
.Y(n_364)
);

AOI21xp5_ASAP7_75t_L g363 ( 
.A1(n_360),
.A2(n_345),
.B(n_346),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_SL g361 ( 
.A(n_357),
.B(n_348),
.Y(n_361)
);

OAI21xp5_ASAP7_75t_L g367 ( 
.A1(n_361),
.A2(n_363),
.B(n_355),
.Y(n_367)
);

OAI22xp5_ASAP7_75t_SL g366 ( 
.A1(n_364),
.A2(n_349),
.B1(n_358),
.B2(n_345),
.Y(n_366)
);

OAI21xp5_ASAP7_75t_SL g365 ( 
.A1(n_362),
.A2(n_353),
.B(n_358),
.Y(n_365)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_365),
.Y(n_368)
);

INVxp33_ASAP7_75t_L g369 ( 
.A(n_366),
.Y(n_369)
);

AOI21xp5_ASAP7_75t_L g370 ( 
.A1(n_368),
.A2(n_367),
.B(n_362),
.Y(n_370)
);

BUFx24_ASAP7_75t_SL g371 ( 
.A(n_370),
.Y(n_371)
);

XOR2xp5_ASAP7_75t_L g372 ( 
.A(n_371),
.B(n_354),
.Y(n_372)
);

XOR2xp5_ASAP7_75t_L g373 ( 
.A(n_372),
.B(n_369),
.Y(n_373)
);


endmodule