module real_aes_3966_n_422 (n_76, n_113, n_187, n_90, n_257, n_390, n_65, n_74, n_185, n_285, n_30, n_222, n_61, n_20, n_287, n_357, n_386, n_64, n_254, n_207, n_10, n_83, n_181, n_362, n_124, n_191, n_209, n_299, n_322, n_328, n_19, n_40, n_318, n_355, n_239, n_100, n_54, n_112, n_319, n_364, n_35, n_42, n_421, n_329, n_132, n_131, n_144, n_169, n_242, n_376, n_308, n_172, n_341, n_232, n_6, n_401, n_69, n_317, n_353, n_321, n_73, n_320, n_77, n_260, n_37, n_97, n_186, n_138, n_379, n_374, n_26, n_235, n_399, n_378, n_245, n_161, n_189, n_271, n_2, n_145, n_415, n_227, n_92, n_330, n_388, n_395, n_332, n_292, n_400, n_116, n_94, n_289, n_280, n_333, n_213, n_356, n_408, n_184, n_28, n_372, n_202, n_56, n_370, n_34, n_98, n_384, n_121, n_352, n_125, n_216, n_82, n_327, n_47, n_106, n_32, n_263, n_230, n_51, n_248, n_301, n_27, n_343, n_369, n_174, n_18, n_104, n_211, n_281, n_173, n_234, n_284, n_153, n_316, n_75, n_178, n_409, n_298, n_49, n_43, n_297, n_383, n_9, n_119, n_310, n_164, n_231, n_44, n_102, n_122, n_141, n_128, n_111, n_167, n_80, n_179, n_12, n_68, n_129, n_345, n_304, n_381, n_311, n_324, n_25, n_278, n_236, n_367, n_267, n_218, n_48, n_204, n_339, n_398, n_89, n_277, n_331, n_93, n_182, n_363, n_417, n_323, n_199, n_350, n_142, n_223, n_67, n_405, n_368, n_250, n_85, n_406, n_45, n_5, n_244, n_118, n_139, n_402, n_87, n_171, n_78, n_146, n_17, n_226, n_255, n_286, n_416, n_410, n_120, n_261, n_238, n_391, n_360, n_58, n_165, n_361, n_246, n_176, n_412, n_163, n_29, n_52, n_251, n_220, n_387, n_197, n_296, n_3, n_41, n_1405, n_256, n_71, n_302, n_351, n_126, n_200, n_115, n_96, n_110, n_392, n_150, n_147, n_288, n_404, n_23, n_334, n_274, n_160, n_303, n_95, n_188, n_269, n_201, n_413, n_306, n_158, n_4, n_366, n_346, n_193, n_397, n_293, n_162, n_358, n_385, n_275, n_214, n_46, n_109, n_59, n_203, n_81, n_133, n_377, n_273, n_114, n_276, n_295, n_382, n_265, n_354, n_154, n_127, n_326, n_24, n_407, n_217, n_419, n_55, n_62, n_411, n_291, n_148, n_88, n_159, n_11, n_108, n_373, n_60, n_233, n_290, n_365, n_155, n_243, n_268, n_136, n_157, n_282, n_389, n_101, n_309, n_344, n_229, n_107, n_33, n_53, n_36, n_149, n_190, n_262, n_134, n_349, n_336, n_420, n_195, n_300, n_252, n_283, n_314, n_249, n_221, n_156, n_359, n_57, n_66, n_21, n_31, n_8, n_312, n_183, n_266, n_205, n_335, n_177, n_313, n_22, n_140, n_418, n_219, n_180, n_212, n_210, n_325, n_338, n_371, n_103, n_166, n_224, n_151, n_130, n_253, n_99, n_15, n_72, n_152, n_198, n_7, n_228, n_272, n_196, n_347, n_315, n_414, n_123, n_279, n_79, n_270, n_305, n_117, n_208, n_215, n_135, n_70, n_50, n_170, n_86, n_375, n_340, n_13, n_380, n_394, n_168, n_175, n_241, n_105, n_84, n_294, n_393, n_258, n_206, n_307, n_396, n_342, n_348, n_14, n_403, n_194, n_137, n_225, n_16, n_39, n_337, n_247, n_240, n_38, n_259, n_143, n_192, n_0, n_264, n_63, n_1, n_237, n_91, n_422);
input n_76;
input n_113;
input n_187;
input n_90;
input n_257;
input n_390;
input n_65;
input n_74;
input n_185;
input n_285;
input n_30;
input n_222;
input n_61;
input n_20;
input n_287;
input n_357;
input n_386;
input n_64;
input n_254;
input n_207;
input n_10;
input n_83;
input n_181;
input n_362;
input n_124;
input n_191;
input n_209;
input n_299;
input n_322;
input n_328;
input n_19;
input n_40;
input n_318;
input n_355;
input n_239;
input n_100;
input n_54;
input n_112;
input n_319;
input n_364;
input n_35;
input n_42;
input n_421;
input n_329;
input n_132;
input n_131;
input n_144;
input n_169;
input n_242;
input n_376;
input n_308;
input n_172;
input n_341;
input n_232;
input n_6;
input n_401;
input n_69;
input n_317;
input n_353;
input n_321;
input n_73;
input n_320;
input n_77;
input n_260;
input n_37;
input n_97;
input n_186;
input n_138;
input n_379;
input n_374;
input n_26;
input n_235;
input n_399;
input n_378;
input n_245;
input n_161;
input n_189;
input n_271;
input n_2;
input n_145;
input n_415;
input n_227;
input n_92;
input n_330;
input n_388;
input n_395;
input n_332;
input n_292;
input n_400;
input n_116;
input n_94;
input n_289;
input n_280;
input n_333;
input n_213;
input n_356;
input n_408;
input n_184;
input n_28;
input n_372;
input n_202;
input n_56;
input n_370;
input n_34;
input n_98;
input n_384;
input n_121;
input n_352;
input n_125;
input n_216;
input n_82;
input n_327;
input n_47;
input n_106;
input n_32;
input n_263;
input n_230;
input n_51;
input n_248;
input n_301;
input n_27;
input n_343;
input n_369;
input n_174;
input n_18;
input n_104;
input n_211;
input n_281;
input n_173;
input n_234;
input n_284;
input n_153;
input n_316;
input n_75;
input n_178;
input n_409;
input n_298;
input n_49;
input n_43;
input n_297;
input n_383;
input n_9;
input n_119;
input n_310;
input n_164;
input n_231;
input n_44;
input n_102;
input n_122;
input n_141;
input n_128;
input n_111;
input n_167;
input n_80;
input n_179;
input n_12;
input n_68;
input n_129;
input n_345;
input n_304;
input n_381;
input n_311;
input n_324;
input n_25;
input n_278;
input n_236;
input n_367;
input n_267;
input n_218;
input n_48;
input n_204;
input n_339;
input n_398;
input n_89;
input n_277;
input n_331;
input n_93;
input n_182;
input n_363;
input n_417;
input n_323;
input n_199;
input n_350;
input n_142;
input n_223;
input n_67;
input n_405;
input n_368;
input n_250;
input n_85;
input n_406;
input n_45;
input n_5;
input n_244;
input n_118;
input n_139;
input n_402;
input n_87;
input n_171;
input n_78;
input n_146;
input n_17;
input n_226;
input n_255;
input n_286;
input n_416;
input n_410;
input n_120;
input n_261;
input n_238;
input n_391;
input n_360;
input n_58;
input n_165;
input n_361;
input n_246;
input n_176;
input n_412;
input n_163;
input n_29;
input n_52;
input n_251;
input n_220;
input n_387;
input n_197;
input n_296;
input n_3;
input n_41;
input n_1405;
input n_256;
input n_71;
input n_302;
input n_351;
input n_126;
input n_200;
input n_115;
input n_96;
input n_110;
input n_392;
input n_150;
input n_147;
input n_288;
input n_404;
input n_23;
input n_334;
input n_274;
input n_160;
input n_303;
input n_95;
input n_188;
input n_269;
input n_201;
input n_413;
input n_306;
input n_158;
input n_4;
input n_366;
input n_346;
input n_193;
input n_397;
input n_293;
input n_162;
input n_358;
input n_385;
input n_275;
input n_214;
input n_46;
input n_109;
input n_59;
input n_203;
input n_81;
input n_133;
input n_377;
input n_273;
input n_114;
input n_276;
input n_295;
input n_382;
input n_265;
input n_354;
input n_154;
input n_127;
input n_326;
input n_24;
input n_407;
input n_217;
input n_419;
input n_55;
input n_62;
input n_411;
input n_291;
input n_148;
input n_88;
input n_159;
input n_11;
input n_108;
input n_373;
input n_60;
input n_233;
input n_290;
input n_365;
input n_155;
input n_243;
input n_268;
input n_136;
input n_157;
input n_282;
input n_389;
input n_101;
input n_309;
input n_344;
input n_229;
input n_107;
input n_33;
input n_53;
input n_36;
input n_149;
input n_190;
input n_262;
input n_134;
input n_349;
input n_336;
input n_420;
input n_195;
input n_300;
input n_252;
input n_283;
input n_314;
input n_249;
input n_221;
input n_156;
input n_359;
input n_57;
input n_66;
input n_21;
input n_31;
input n_8;
input n_312;
input n_183;
input n_266;
input n_205;
input n_335;
input n_177;
input n_313;
input n_22;
input n_140;
input n_418;
input n_219;
input n_180;
input n_212;
input n_210;
input n_325;
input n_338;
input n_371;
input n_103;
input n_166;
input n_224;
input n_151;
input n_130;
input n_253;
input n_99;
input n_15;
input n_72;
input n_152;
input n_198;
input n_7;
input n_228;
input n_272;
input n_196;
input n_347;
input n_315;
input n_414;
input n_123;
input n_279;
input n_79;
input n_270;
input n_305;
input n_117;
input n_208;
input n_215;
input n_135;
input n_70;
input n_50;
input n_170;
input n_86;
input n_375;
input n_340;
input n_13;
input n_380;
input n_394;
input n_168;
input n_175;
input n_241;
input n_105;
input n_84;
input n_294;
input n_393;
input n_258;
input n_206;
input n_307;
input n_396;
input n_342;
input n_348;
input n_14;
input n_403;
input n_194;
input n_137;
input n_225;
input n_16;
input n_39;
input n_337;
input n_247;
input n_240;
input n_38;
input n_259;
input n_143;
input n_192;
input n_0;
input n_264;
input n_63;
input n_1;
input n_237;
input n_91;
output n_422;
wire n_476;
wire n_599;
wire n_887;
wire n_1279;
wire n_1314;
wire n_830;
wire n_1371;
wire n_624;
wire n_618;
wire n_933;
wire n_485;
wire n_822;
wire n_750;
wire n_503;
wire n_469;
wire n_1310;
wire n_1376;
wire n_592;
wire n_761;
wire n_919;
wire n_1217;
wire n_571;
wire n_549;
wire n_1034;
wire n_1328;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_593;
wire n_989;
wire n_431;
wire n_1044;
wire n_963;
wire n_551;
wire n_884;
wire n_814;
wire n_944;
wire n_1283;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_1313;
wire n_870;
wire n_1248;
wire n_548;
wire n_572;
wire n_815;
wire n_1140;
wire n_786;
wire n_512;
wire n_795;
wire n_1379;
wire n_1160;
wire n_1287;
wire n_883;
wire n_478;
wire n_553;
wire n_744;
wire n_1367;
wire n_1325;
wire n_1382;
wire n_1225;
wire n_875;
wire n_951;
wire n_1199;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_595;
wire n_1282;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_962;
wire n_755;
wire n_781;
wire n_576;
wire n_956;
wire n_1242;
wire n_796;
wire n_874;
wire n_1126;
wire n_455;
wire n_682;
wire n_812;
wire n_817;
wire n_782;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_1020;
wire n_885;
wire n_950;
wire n_1196;
wire n_1013;
wire n_808;
wire n_1224;
wire n_688;
wire n_1042;
wire n_1317;
wire n_690;
wire n_499;
wire n_1142;
wire n_947;
wire n_970;
wire n_1149;
wire n_527;
wire n_1342;
wire n_552;
wire n_1383;
wire n_1346;
wire n_590;
wire n_1293;
wire n_432;
wire n_1131;
wire n_1008;
wire n_805;
wire n_619;
wire n_1095;
wire n_1250;
wire n_1284;
wire n_859;
wire n_1304;
wire n_685;
wire n_1080;
wire n_917;
wire n_1247;
wire n_501;
wire n_488;
wire n_1380;
wire n_954;
wire n_702;
wire n_1007;
wire n_898;
wire n_562;
wire n_1022;
wire n_1073;
wire n_728;
wire n_1301;
wire n_1201;
wire n_997;
wire n_1105;
wire n_1243;
wire n_1003;
wire n_749;
wire n_914;
wire n_1286;
wire n_494;
wire n_927;
wire n_723;
wire n_972;
wire n_1351;
wire n_1209;
wire n_498;
wire n_1397;
wire n_765;
wire n_648;
wire n_939;
wire n_928;
wire n_1384;
wire n_789;
wire n_738;
wire n_1387;
wire n_922;
wire n_1048;
wire n_787;
wire n_1214;
wire n_806;
wire n_715;
wire n_1258;
wire n_873;
wire n_438;
wire n_446;
wire n_1281;
wire n_712;
wire n_861;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_724;
wire n_440;
wire n_1231;
wire n_1305;
wire n_1161;
wire n_686;
wire n_1299;
wire n_949;
wire n_586;
wire n_788;
wire n_441;
wire n_1045;
wire n_1339;
wire n_837;
wire n_1349;
wire n_829;
wire n_1030;
wire n_1348;
wire n_1391;
wire n_597;
wire n_1036;
wire n_687;
wire n_652;
wire n_500;
wire n_804;
wire n_1173;
wire n_854;
wire n_424;
wire n_877;
wire n_802;
wire n_480;
wire n_684;
wire n_1178;
wire n_821;
wire n_1018;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_635;
wire n_792;
wire n_1392;
wire n_665;
wire n_667;
wire n_991;
wire n_580;
wire n_1004;
wire n_1370;
wire n_979;
wire n_445;
wire n_596;
wire n_1197;
wire n_657;
wire n_1260;
wire n_1129;
wire n_1285;
wire n_742;
wire n_1014;
wire n_1385;
wire n_461;
wire n_1047;
wire n_1016;
wire n_694;
wire n_1350;
wire n_894;
wire n_545;
wire n_538;
wire n_537;
wire n_560;
wire n_1094;
wire n_1220;
wire n_696;
wire n_1147;
wire n_704;
wire n_453;
wire n_647;
wire n_948;
wire n_700;
wire n_677;
wire n_1269;
wire n_591;
wire n_1366;
wire n_678;
wire n_1400;
wire n_564;
wire n_638;
wire n_510;
wire n_1361;
wire n_1358;
wire n_550;
wire n_966;
wire n_1368;
wire n_994;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_992;
wire n_813;
wire n_981;
wire n_1338;
wire n_1182;
wire n_872;
wire n_1401;
wire n_1086;
wire n_1070;
wire n_1189;
wire n_535;
wire n_882;
wire n_1210;
wire n_746;
wire n_656;
wire n_1148;
wire n_860;
wire n_748;
wire n_1261;
wire n_1062;
wire n_651;
wire n_801;
wire n_1271;
wire n_529;
wire n_504;
wire n_973;
wire n_1364;
wire n_659;
wire n_634;
wire n_903;
wire n_565;
wire n_925;
wire n_1389;
wire n_1393;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_1362;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_754;
wire n_508;
wire n_1141;
wire n_1112;
wire n_428;
wire n_783;
wire n_1107;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1386;
wire n_617;
wire n_733;
wire n_602;
wire n_658;
wire n_676;
wire n_531;
wire n_1031;
wire n_1394;
wire n_807;
wire n_1011;
wire n_895;
wire n_799;
wire n_490;
wire n_695;
wire n_1181;
wire n_881;
wire n_645;
wire n_1145;
wire n_557;
wire n_777;
wire n_985;
wire n_910;
wire n_642;
wire n_613;
wire n_1125;
wire n_1347;
wire n_1163;
wire n_1278;
wire n_734;
wire n_735;
wire n_1179;
wire n_569;
wire n_1171;
wire n_785;
wire n_1203;
wire n_1232;
wire n_471;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1187;
wire n_1000;
wire n_649;
wire n_1234;
wire n_622;
wire n_1353;
wire n_1002;
wire n_1165;
wire n_1058;
wire n_1216;
wire n_662;
wire n_850;
wire n_720;
wire n_1026;
wire n_492;
wire n_1023;
wire n_730;
wire n_643;
wire n_1403;
wire n_486;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_526;
wire n_1194;
wire n_701;
wire n_809;
wire n_520;
wire n_679;
wire n_926;
wire n_942;
wire n_1374;
wire n_1120;
wire n_689;
wire n_946;
wire n_753;
wire n_1188;
wire n_623;
wire n_1032;
wire n_721;
wire n_1133;
wire n_739;
wire n_1322;
wire n_1162;
wire n_762;
wire n_1298;
wire n_442;
wire n_740;
wire n_1357;
wire n_639;
wire n_1186;
wire n_1365;
wire n_459;
wire n_1172;
wire n_998;
wire n_1395;
wire n_1276;
wire n_836;
wire n_1184;
wire n_583;
wire n_1336;
wire n_776;
wire n_1138;
wire n_890;
wire n_1306;
wire n_1266;
wire n_497;
wire n_911;
wire n_450;
wire n_473;
wire n_967;
wire n_474;
wire n_1159;
wire n_1315;
wire n_1055;
wire n_611;
wire n_844;
wire n_968;
wire n_710;
wire n_1040;
wire n_1102;
wire n_661;
wire n_1185;
wire n_447;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1069;
wire n_842;
wire n_798;
wire n_668;
wire n_862;
wire n_869;
wire n_1066;
wire n_1377;
wire n_800;
wire n_1175;
wire n_778;
wire n_1170;
wire n_522;
wire n_943;
wire n_977;
wire n_905;
wire n_878;
wire n_1333;
wire n_577;
wire n_759;
wire n_1235;
wire n_900;
wire n_841;
wire n_1218;
wire n_736;
wire n_766;
wire n_852;
wire n_1113;
wire n_1268;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_1302;
wire n_1289;
wire n_937;
wire n_773;
wire n_865;
wire n_594;
wire n_856;
wire n_1146;
wire n_932;
wire n_958;
wire n_775;
wire n_763;
wire n_1093;
wire n_427;
wire n_519;
wire n_1116;
wire n_709;
wire n_816;
wire n_625;
wire n_953;
wire n_1373;
wire n_716;
wire n_584;
wire n_896;
wire n_528;
wire n_1078;
wire n_495;
wire n_1072;
wire n_935;
wire n_467;
wire n_1213;
wire n_1053;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_1168;
wire n_1309;
wire n_909;
wire n_523;
wire n_996;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1332;
wire n_1263;
wire n_1115;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_454;
wire n_1303;
wire n_443;
wire n_1029;
wire n_1207;
wire n_664;
wire n_1017;
wire n_581;
wire n_936;
wire n_1215;
wire n_582;
wire n_641;
wire n_940;
wire n_745;
wire n_1167;
wire n_1327;
wire n_609;
wire n_1006;
wire n_1259;
wire n_561;
wire n_437;
wire n_1223;
wire n_621;
wire n_1012;
wire n_1241;
wire n_502;
wire n_434;
wire n_769;
wire n_1212;
wire n_1054;
wire n_1308;
wire n_1050;
wire n_426;
wire n_1134;
wire n_1319;
wire n_1363;
wire n_616;
wire n_880;
wire n_1103;
wire n_1274;
wire n_832;
wire n_1321;
wire n_1060;
wire n_1154;
wire n_632;
wire n_1344;
wire n_714;
wire n_1331;
wire n_1222;
wire n_1041;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_1335;
wire n_912;
wire n_464;
wire n_1227;
wire n_945;
wire n_563;
wire n_891;
wire n_568;
wire n_1157;
wire n_902;
wire n_1158;
wire n_1079;
wire n_1330;
wire n_1033;
wire n_1028;
wire n_727;
wire n_1083;
wire n_1056;
wire n_663;
wire n_588;
wire n_707;
wire n_915;
wire n_1001;
wire n_711;
wire n_864;
wire n_1169;
wire n_1139;
wire n_1038;
wire n_1085;
wire n_845;
wire n_1127;
wire n_484;
wire n_893;
wire n_1068;
wire n_747;
wire n_1244;
wire n_697;
wire n_978;
wire n_847;
wire n_826;
wire n_628;
wire n_487;
wire n_831;
wire n_653;
wire n_692;
wire n_1051;
wire n_1355;
wire n_827;
wire n_472;
wire n_866;
wire n_452;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_858;
wire n_764;
wire n_741;
wire n_1090;
wire n_456;
wire n_1164;
wire n_433;
wire n_627;
wire n_771;
wire n_524;
wire n_1378;
wire n_705;
wire n_1191;
wire n_1206;
wire n_1270;
wire n_1399;
wire n_546;
wire n_1010;
wire n_1375;
wire n_1015;
wire n_863;
wire n_525;
wire n_1226;
wire n_644;
wire n_1150;
wire n_1341;
wire n_833;
wire n_1229;
wire n_929;
wire n_1143;
wire n_1190;
wire n_543;
wire n_585;
wire n_465;
wire n_719;
wire n_1343;
wire n_1156;
wire n_988;
wire n_1396;
wire n_921;
wire n_640;
wire n_1176;
wire n_1151;
wire n_1254;
wire n_646;
wire n_650;
wire n_1211;
wire n_743;
wire n_823;
wire n_1101;
wire n_1076;
wire n_1251;
wire n_1104;
wire n_849;
wire n_1061;
wire n_554;
wire n_1153;
wire n_1337;
wire n_797;
wire n_1177;
wire n_758;
wire n_436;
wire n_1096;
wire n_1316;
wire n_1092;
wire n_846;
wire n_631;
wire n_673;
wire n_1067;
wire n_518;
wire n_1192;
wire n_1292;
wire n_1240;
wire n_987;
wire n_1065;
wire n_540;
wire n_1064;
wire n_1075;
wire n_718;
wire n_669;
wire n_1091;
wire n_423;
wire n_1221;
wire n_458;
wire n_1200;
wire n_444;
wire n_555;
wire n_1295;
wire n_974;
wire n_1329;
wire n_857;
wire n_491;
wire n_1294;
wire n_1110;
wire n_1137;
wire n_460;
wire n_666;
wire n_660;
wire n_1359;
wire n_886;
wire n_767;
wire n_889;
wire n_1398;
wire n_1021;
wire n_1297;
wire n_1046;
wire n_1109;
wire n_961;
wire n_489;
wire n_1381;
wire n_573;
wire n_1099;
wire n_626;
wire n_539;
wire n_462;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_1272;
wire n_578;
wire n_892;
wire n_938;
wire n_774;
wire n_466;
wire n_559;
wire n_1049;
wire n_1277;
wire n_984;
wire n_726;
wire n_517;
wire n_931;
wire n_780;
wire n_530;
wire n_834;
wire n_693;
wire n_496;
wire n_1360;
wire n_1082;
wire n_1257;
wire n_468;
wire n_532;
wire n_1025;
wire n_924;
wire n_1264;
wire n_1245;
wire n_1152;
wire n_1081;
wire n_547;
wire n_1324;
wire n_1198;
wire n_1307;
wire n_993;
wire n_819;
wire n_737;
wire n_1318;
wire n_1290;
wire n_1135;
wire n_1063;
wire n_828;
wire n_770;
wire n_867;
wire n_1100;
wire n_425;
wire n_879;
wire n_449;
wire n_1340;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_655;
wire n_654;
wire n_672;
wire n_567;
wire n_916;
wire n_1354;
wire n_1334;
wire n_1291;
wire n_986;
wire n_451;
wire n_1037;
wire n_1267;
wire n_790;
wire n_1262;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_1356;
wire n_768;
wire n_542;
wire n_1256;
wire n_1077;
wire n_1111;
wire n_1249;
wire n_1239;
wire n_969;
wire n_1009;
wire n_1202;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_430;
wire n_1252;
wire n_1132;
wire n_1275;
wire n_843;
wire n_579;
wire n_533;
wire n_536;
wire n_470;
wire n_851;
wire n_1155;
wire n_934;
wire n_1027;
wire n_965;
wire n_1296;
wire n_1043;
wire n_435;
wire n_511;
wire n_509;
wire n_1204;
wire n_930;
wire n_1265;
wire n_1057;
wire n_907;
wire n_1005;
wire n_1312;
wire n_899;
wire n_637;
wire n_544;
wire n_1087;
wire n_482;
wire n_633;
wire n_971;
wire n_1052;
wire n_1071;
wire n_1311;
wire n_1273;
wire n_959;
wire n_1130;
wire n_794;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1253;
wire n_1183;
wire n_516;
wire n_521;
wire n_1195;
wire n_575;
wire n_1300;
wire n_1372;
wire n_698;
wire n_1345;
wire n_587;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_793;
wire n_1390;
wire n_757;
wire n_803;
wire n_514;
wire n_507;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1088;
wire n_1230;
wire n_1326;
wire n_1402;
wire n_1388;
wire n_483;
wire n_729;
wire n_1280;
wire n_1323;
wire n_1352;
wire n_1369;
wire n_703;
wire n_1097;
wire n_601;
wire n_463;
wire n_1236;
wire n_603;
wire n_1288;
wire n_868;
wire n_1024;
wire n_1144;
wire n_475;
wire n_897;
wire n_1320;
wire n_855;
wire n_429;
INVx1_ASAP7_75t_L g1359 ( .A(n_0), .Y(n_1359) );
AOI22xp5_ASAP7_75t_L g1365 ( .A1(n_1), .A2(n_342), .B1(n_477), .B2(n_802), .Y(n_1365) );
AOI22xp33_ASAP7_75t_L g488 ( .A1(n_2), .A2(n_121), .B1(n_489), .B2(n_491), .Y(n_488) );
AOI22x1_ASAP7_75t_L g1003 ( .A1(n_3), .A2(n_269), .B1(n_635), .B2(n_828), .Y(n_1003) );
AOI22xp33_ASAP7_75t_L g597 ( .A1(n_4), .A2(n_171), .B1(n_598), .B2(n_599), .Y(n_597) );
AOI22xp33_ASAP7_75t_L g928 ( .A1(n_5), .A2(n_385), .B1(n_501), .B2(n_929), .Y(n_928) );
AOI22xp33_ASAP7_75t_L g740 ( .A1(n_6), .A2(n_326), .B1(n_741), .B2(n_742), .Y(n_740) );
AOI22xp33_ASAP7_75t_L g899 ( .A1(n_7), .A2(n_218), .B1(n_477), .B2(n_542), .Y(n_899) );
AOI22xp33_ASAP7_75t_L g973 ( .A1(n_8), .A2(n_386), .B1(n_555), .B2(n_974), .Y(n_973) );
CKINVDCx20_ASAP7_75t_R g1221 ( .A(n_9), .Y(n_1221) );
AO22x1_ASAP7_75t_L g1050 ( .A1(n_10), .A2(n_222), .B1(n_1051), .B2(n_1052), .Y(n_1050) );
AOI221xp5_ASAP7_75t_L g675 ( .A1(n_11), .A2(n_341), .B1(n_554), .B2(n_676), .C(n_678), .Y(n_675) );
AOI22xp33_ASAP7_75t_L g714 ( .A1(n_12), .A2(n_363), .B1(n_576), .B2(n_578), .Y(n_714) );
AOI22xp5_ASAP7_75t_L g1015 ( .A1(n_13), .A2(n_354), .B1(n_780), .B2(n_934), .Y(n_1015) );
AOI22xp5_ASAP7_75t_L g969 ( .A1(n_14), .A2(n_98), .B1(n_970), .B2(n_971), .Y(n_969) );
AOI22xp33_ASAP7_75t_L g591 ( .A1(n_15), .A2(n_241), .B1(n_592), .B2(n_593), .Y(n_591) );
NAND2xp5_ASAP7_75t_SL g451 ( .A(n_16), .B(n_439), .Y(n_451) );
AOI22xp33_ASAP7_75t_L g830 ( .A1(n_17), .A2(n_356), .B1(n_458), .B2(n_544), .Y(n_830) );
AOI22xp33_ASAP7_75t_L g925 ( .A1(n_18), .A2(n_232), .B1(n_489), .B2(n_635), .Y(n_925) );
AOI22xp33_ASAP7_75t_L g682 ( .A1(n_19), .A2(n_323), .B1(n_516), .B2(n_551), .Y(n_682) );
AOI22xp33_ASAP7_75t_SL g1394 ( .A1(n_20), .A2(n_204), .B1(n_489), .B2(n_635), .Y(n_1394) );
AOI22xp33_ASAP7_75t_L g692 ( .A1(n_21), .A2(n_108), .B1(n_477), .B2(n_658), .Y(n_692) );
INVx1_ASAP7_75t_SL g619 ( .A(n_22), .Y(n_619) );
INVx1_ASAP7_75t_L g1070 ( .A(n_23), .Y(n_1070) );
INVx1_ASAP7_75t_L g781 ( .A(n_24), .Y(n_781) );
BUFx6f_ASAP7_75t_L g439 ( .A(n_25), .Y(n_439) );
AOI22xp5_ASAP7_75t_L g978 ( .A1(n_26), .A2(n_398), .B1(n_473), .B2(n_667), .Y(n_978) );
AOI22xp33_ASAP7_75t_L g810 ( .A1(n_27), .A2(n_39), .B1(n_595), .B2(n_598), .Y(n_810) );
AOI22xp33_ASAP7_75t_L g836 ( .A1(n_28), .A2(n_147), .B1(n_555), .B2(n_837), .Y(n_836) );
INVx1_ASAP7_75t_L g957 ( .A(n_29), .Y(n_957) );
AOI22xp33_ASAP7_75t_L g722 ( .A1(n_30), .A2(n_85), .B1(n_596), .B2(n_599), .Y(n_722) );
AOI22xp33_ASAP7_75t_L g833 ( .A1(n_31), .A2(n_169), .B1(n_477), .B2(n_542), .Y(n_833) );
AOI22xp33_ASAP7_75t_L g882 ( .A1(n_32), .A2(n_270), .B1(n_579), .B2(n_589), .Y(n_882) );
AOI22xp33_ASAP7_75t_L g856 ( .A1(n_33), .A2(n_76), .B1(n_655), .B2(n_658), .Y(n_856) );
NAND2xp5_ASAP7_75t_L g813 ( .A(n_34), .B(n_560), .Y(n_813) );
AOI22xp33_ASAP7_75t_L g930 ( .A1(n_35), .A2(n_340), .B1(n_931), .B2(n_933), .Y(n_930) );
AOI22xp5_ASAP7_75t_L g691 ( .A1(n_36), .A2(n_193), .B1(n_548), .B2(n_635), .Y(n_691) );
AOI22xp33_ASAP7_75t_L g671 ( .A1(n_37), .A2(n_214), .B1(n_658), .B2(n_672), .Y(n_671) );
AOI22xp33_ASAP7_75t_L g1352 ( .A1(n_38), .A2(n_133), .B1(n_701), .B2(n_1353), .Y(n_1352) );
AOI21xp33_ASAP7_75t_L g1080 ( .A1(n_40), .A2(n_560), .B(n_1081), .Y(n_1080) );
AO22x1_ASAP7_75t_L g773 ( .A1(n_41), .A2(n_61), .B1(n_774), .B2(n_775), .Y(n_773) );
AOI22xp33_ASAP7_75t_L g862 ( .A1(n_42), .A2(n_63), .B1(n_787), .B2(n_863), .Y(n_862) );
INVx1_ASAP7_75t_L g1358 ( .A(n_43), .Y(n_1358) );
AOI21xp5_ASAP7_75t_L g557 ( .A1(n_44), .A2(n_558), .B(n_561), .Y(n_557) );
AOI22xp33_ASAP7_75t_L g1020 ( .A1(n_45), .A2(n_229), .B1(n_516), .B2(n_776), .Y(n_1020) );
INVx1_ASAP7_75t_L g585 ( .A(n_46), .Y(n_585) );
AOI22xp33_ASAP7_75t_L g950 ( .A1(n_47), .A2(n_125), .B1(n_544), .B2(n_795), .Y(n_950) );
AOI22xp33_ASAP7_75t_L g1122 ( .A1(n_48), .A2(n_184), .B1(n_1114), .B2(n_1116), .Y(n_1122) );
AOI22xp33_ASAP7_75t_L g962 ( .A1(n_49), .A2(n_57), .B1(n_516), .B2(n_758), .Y(n_962) );
AOI22xp33_ASAP7_75t_L g515 ( .A1(n_50), .A2(n_256), .B1(n_516), .B2(n_526), .Y(n_515) );
AOI22xp33_ASAP7_75t_L g818 ( .A1(n_51), .A2(n_115), .B1(n_579), .B2(n_819), .Y(n_818) );
AOI22xp5_ASAP7_75t_L g1085 ( .A1(n_52), .A2(n_399), .B1(n_743), .B2(n_878), .Y(n_1085) );
AOI22xp33_ASAP7_75t_SL g1395 ( .A1(n_53), .A2(n_303), .B1(n_458), .B2(n_544), .Y(n_1395) );
AOI22xp33_ASAP7_75t_L g1042 ( .A1(n_54), .A2(n_404), .B1(n_590), .B2(n_596), .Y(n_1042) );
AOI22xp33_ASAP7_75t_L g689 ( .A1(n_55), .A2(n_158), .B1(n_458), .B2(n_473), .Y(n_689) );
CKINVDCx20_ASAP7_75t_R g873 ( .A(n_56), .Y(n_873) );
AOI22xp33_ASAP7_75t_L g1035 ( .A1(n_58), .A2(n_346), .B1(n_578), .B2(n_579), .Y(n_1035) );
NAND2xp5_ASAP7_75t_L g752 ( .A(n_59), .B(n_566), .Y(n_752) );
NAND2xp5_ASAP7_75t_L g942 ( .A(n_60), .B(n_943), .Y(n_942) );
OA22x2_ASAP7_75t_L g445 ( .A1(n_62), .A2(n_181), .B1(n_439), .B2(n_443), .Y(n_445) );
INVx1_ASAP7_75t_L g464 ( .A(n_62), .Y(n_464) );
AOI22xp33_ASAP7_75t_L g897 ( .A1(n_64), .A2(n_142), .B1(n_489), .B2(n_635), .Y(n_897) );
AOI221xp5_ASAP7_75t_L g694 ( .A1(n_65), .A2(n_78), .B1(n_695), .B2(n_697), .C(n_698), .Y(n_694) );
AOI22xp33_ASAP7_75t_L g980 ( .A1(n_66), .A2(n_357), .B1(n_658), .B2(n_672), .Y(n_980) );
AOI221x1_ASAP7_75t_L g1012 ( .A1(n_67), .A2(n_308), .B1(n_655), .B2(n_885), .C(n_1013), .Y(n_1012) );
AOI22xp33_ASAP7_75t_L g922 ( .A1(n_68), .A2(n_368), .B1(n_458), .B2(n_544), .Y(n_922) );
INVx1_ASAP7_75t_L g1136 ( .A(n_69), .Y(n_1136) );
AOI22xp33_ASAP7_75t_L g1178 ( .A1(n_70), .A2(n_167), .B1(n_1127), .B2(n_1135), .Y(n_1178) );
AOI221xp5_ASAP7_75t_L g1001 ( .A1(n_71), .A2(n_288), .B1(n_800), .B2(n_802), .C(n_1002), .Y(n_1001) );
AOI22xp33_ASAP7_75t_L g906 ( .A1(n_72), .A2(n_333), .B1(n_552), .B2(n_703), .Y(n_906) );
AOI22xp5_ASAP7_75t_L g854 ( .A1(n_73), .A2(n_166), .B1(n_473), .B2(n_855), .Y(n_854) );
AOI22xp33_ASAP7_75t_L g577 ( .A1(n_74), .A2(n_388), .B1(n_578), .B2(n_579), .Y(n_577) );
INVx1_ASAP7_75t_SL g1138 ( .A(n_75), .Y(n_1138) );
INVx1_ASAP7_75t_L g442 ( .A(n_77), .Y(n_442) );
OAI21xp33_ASAP7_75t_L g465 ( .A1(n_77), .A2(n_181), .B(n_466), .Y(n_465) );
NOR2xp33_ASAP7_75t_L g532 ( .A(n_77), .B(n_206), .Y(n_532) );
AOI22xp33_ASAP7_75t_L g799 ( .A1(n_79), .A2(n_365), .B1(n_800), .B2(n_802), .Y(n_799) );
INVx1_ASAP7_75t_L g1031 ( .A(n_80), .Y(n_1031) );
AOI22xp33_ASAP7_75t_L g979 ( .A1(n_81), .A2(n_118), .B1(n_433), .B2(n_634), .Y(n_979) );
INVx1_ASAP7_75t_L g538 ( .A(n_82), .Y(n_538) );
AOI22xp5_ASAP7_75t_L g1106 ( .A1(n_82), .A2(n_122), .B1(n_1107), .B2(n_1111), .Y(n_1106) );
AOI22xp33_ASAP7_75t_L g753 ( .A1(n_83), .A2(n_197), .B1(n_754), .B2(n_755), .Y(n_753) );
AOI22xp33_ASAP7_75t_L g808 ( .A1(n_84), .A2(n_275), .B1(n_575), .B2(n_599), .Y(n_808) );
NOR3xp33_ASAP7_75t_L g1009 ( .A(n_86), .B(n_1010), .C(n_1014), .Y(n_1009) );
AOI22xp5_ASAP7_75t_L g1027 ( .A1(n_86), .A2(n_1014), .B1(n_1019), .B2(n_1405), .Y(n_1027) );
OAI21xp5_ASAP7_75t_L g1028 ( .A1(n_86), .A2(n_1010), .B(n_1022), .Y(n_1028) );
INVx1_ASAP7_75t_SL g647 ( .A(n_87), .Y(n_647) );
INVx1_ASAP7_75t_L g1382 ( .A(n_88), .Y(n_1382) );
AOI22xp33_ASAP7_75t_L g811 ( .A1(n_89), .A2(n_189), .B1(n_592), .B2(n_593), .Y(n_811) );
AOI21xp33_ASAP7_75t_L g815 ( .A1(n_90), .A2(n_589), .B(n_816), .Y(n_815) );
AOI22xp33_ASAP7_75t_L g949 ( .A1(n_91), .A2(n_94), .B1(n_548), .B2(n_736), .Y(n_949) );
AOI22xp33_ASAP7_75t_L g797 ( .A1(n_92), .A2(n_238), .B1(n_741), .B2(n_798), .Y(n_797) );
INVx1_ASAP7_75t_L g1109 ( .A(n_93), .Y(n_1109) );
AND2x4_ASAP7_75t_L g1112 ( .A(n_93), .B(n_321), .Y(n_1112) );
HB1xp67_ASAP7_75t_L g1402 ( .A(n_93), .Y(n_1402) );
AOI22xp33_ASAP7_75t_L g496 ( .A1(n_95), .A2(n_107), .B1(n_497), .B2(n_501), .Y(n_496) );
AOI22xp33_ASAP7_75t_L g809 ( .A1(n_96), .A2(n_102), .B1(n_590), .B2(n_596), .Y(n_809) );
AOI22xp33_ASAP7_75t_L g1129 ( .A1(n_97), .A2(n_377), .B1(n_1107), .B2(n_1124), .Y(n_1129) );
AOI22xp33_ASAP7_75t_L g553 ( .A1(n_99), .A2(n_276), .B1(n_554), .B2(n_555), .Y(n_553) );
AOI21xp33_ASAP7_75t_L g582 ( .A1(n_100), .A2(n_583), .B(n_584), .Y(n_582) );
AOI21xp5_ASAP7_75t_L g903 ( .A1(n_101), .A2(n_776), .B(n_904), .Y(n_903) );
XOR2xp5_ASAP7_75t_L g946 ( .A(n_103), .B(n_947), .Y(n_946) );
AOI211xp5_ASAP7_75t_L g992 ( .A1(n_104), .A2(n_993), .B(n_995), .C(n_999), .Y(n_992) );
XNOR2x1_ASAP7_75t_L g711 ( .A(n_105), .B(n_712), .Y(n_711) );
AO22x2_ASAP7_75t_L g1152 ( .A1(n_105), .A2(n_349), .B1(n_1107), .B2(n_1124), .Y(n_1152) );
AOI22xp33_ASAP7_75t_L g1043 ( .A1(n_106), .A2(n_129), .B1(n_595), .B2(n_598), .Y(n_1043) );
AOI22xp33_ASAP7_75t_L g476 ( .A1(n_109), .A2(n_177), .B1(n_477), .B2(n_481), .Y(n_476) );
AOI22xp5_ASAP7_75t_L g996 ( .A1(n_110), .A2(n_224), .B1(n_501), .B2(n_695), .Y(n_996) );
AOI22xp33_ASAP7_75t_L g1146 ( .A1(n_111), .A2(n_150), .B1(n_1135), .B2(n_1147), .Y(n_1146) );
AOI22xp33_ASAP7_75t_L g1366 ( .A1(n_112), .A2(n_355), .B1(n_468), .B2(n_829), .Y(n_1366) );
AOI22xp5_ASAP7_75t_L g881 ( .A1(n_113), .A2(n_182), .B1(n_578), .B2(n_787), .Y(n_881) );
AOI22xp5_ASAP7_75t_L g1113 ( .A1(n_114), .A2(n_152), .B1(n_1114), .B2(n_1116), .Y(n_1113) );
INVx1_ASAP7_75t_L g1039 ( .A(n_116), .Y(n_1039) );
INVx1_ASAP7_75t_SL g614 ( .A(n_117), .Y(n_614) );
AOI22xp5_ASAP7_75t_L g541 ( .A1(n_119), .A2(n_296), .B1(n_477), .B2(n_542), .Y(n_541) );
INVx1_ASAP7_75t_L g871 ( .A(n_120), .Y(n_871) );
INVx1_ASAP7_75t_SL g621 ( .A(n_123), .Y(n_621) );
AOI22xp33_ASAP7_75t_L g858 ( .A1(n_124), .A2(n_148), .B1(n_548), .B2(n_792), .Y(n_858) );
AND2x4_ASAP7_75t_L g1110 ( .A(n_126), .B(n_1095), .Y(n_1110) );
INVx1_ASAP7_75t_SL g1115 ( .A(n_126), .Y(n_1115) );
INVx1_ASAP7_75t_L g1118 ( .A(n_126), .Y(n_1118) );
AOI22xp33_ASAP7_75t_L g892 ( .A1(n_127), .A2(n_414), .B1(n_655), .B2(n_658), .Y(n_892) );
AOI22xp33_ASAP7_75t_L g690 ( .A1(n_128), .A2(n_131), .B1(n_433), .B2(n_634), .Y(n_690) );
AOI22xp33_ASAP7_75t_L g724 ( .A1(n_130), .A2(n_319), .B1(n_590), .B2(n_598), .Y(n_724) );
INVx1_ASAP7_75t_L g1377 ( .A(n_132), .Y(n_1377) );
AOI22xp33_ASAP7_75t_L g835 ( .A1(n_134), .A2(n_394), .B1(n_507), .B2(n_551), .Y(n_835) );
XNOR2x1_ASAP7_75t_L g571 ( .A(n_135), .B(n_572), .Y(n_571) );
AOI22xp33_ASAP7_75t_L g1123 ( .A1(n_135), .A2(n_159), .B1(n_1107), .B2(n_1124), .Y(n_1123) );
AOI22xp33_ASAP7_75t_L g814 ( .A1(n_136), .A2(n_352), .B1(n_576), .B2(n_578), .Y(n_814) );
AOI22xp33_ASAP7_75t_L g827 ( .A1(n_137), .A2(n_178), .B1(n_828), .B2(n_829), .Y(n_827) );
NAND2xp5_ASAP7_75t_L g1077 ( .A(n_138), .B(n_554), .Y(n_1077) );
AOI22xp5_ASAP7_75t_L g1148 ( .A1(n_139), .A2(n_421), .B1(n_1107), .B2(n_1127), .Y(n_1148) );
AOI22xp33_ASAP7_75t_L g877 ( .A1(n_140), .A2(n_272), .B1(n_878), .B2(n_879), .Y(n_877) );
AOI22xp5_ASAP7_75t_L g908 ( .A1(n_141), .A2(n_325), .B1(n_497), .B2(n_501), .Y(n_908) );
AOI22xp33_ASAP7_75t_L g550 ( .A1(n_143), .A2(n_364), .B1(n_551), .B2(n_552), .Y(n_550) );
AOI22xp33_ASAP7_75t_L g547 ( .A1(n_144), .A2(n_188), .B1(n_473), .B2(n_548), .Y(n_547) );
AOI22xp33_ASAP7_75t_L g594 ( .A1(n_145), .A2(n_194), .B1(n_595), .B2(n_596), .Y(n_594) );
AOI22xp33_ASAP7_75t_L g737 ( .A1(n_146), .A2(n_400), .B1(n_738), .B2(n_739), .Y(n_737) );
INVx1_ASAP7_75t_L g749 ( .A(n_149), .Y(n_749) );
NAND2xp5_ASAP7_75t_L g580 ( .A(n_151), .B(n_581), .Y(n_580) );
NAND2xp33_ASAP7_75t_L g1011 ( .A(n_153), .B(n_795), .Y(n_1011) );
AOI22xp33_ASAP7_75t_L g1388 ( .A1(n_154), .A2(n_401), .B1(n_566), .B2(n_751), .Y(n_1388) );
AOI22xp5_ASAP7_75t_L g898 ( .A1(n_155), .A2(n_411), .B1(n_468), .B2(n_473), .Y(n_898) );
AOI22xp33_ASAP7_75t_L g1054 ( .A1(n_156), .A2(n_316), .B1(n_800), .B2(n_1024), .Y(n_1054) );
INVx1_ASAP7_75t_L g1062 ( .A(n_157), .Y(n_1062) );
INVx1_ASAP7_75t_L g612 ( .A(n_160), .Y(n_612) );
AOI22xp5_ASAP7_75t_L g880 ( .A1(n_161), .A2(n_199), .B1(n_634), .B2(n_670), .Y(n_880) );
AOI22xp33_ASAP7_75t_L g859 ( .A1(n_162), .A2(n_207), .B1(n_433), .B2(n_860), .Y(n_859) );
AOI22xp33_ASAP7_75t_L g1363 ( .A1(n_163), .A2(n_165), .B1(n_458), .B2(n_473), .Y(n_1363) );
INVxp67_ASAP7_75t_SL g918 ( .A(n_164), .Y(n_918) );
AOI22xp5_ASAP7_75t_L g730 ( .A1(n_168), .A2(n_268), .B1(n_637), .B2(n_731), .Y(n_730) );
AOI22xp33_ASAP7_75t_L g923 ( .A1(n_170), .A2(n_417), .B1(n_468), .B2(n_473), .Y(n_923) );
INVx1_ASAP7_75t_L g817 ( .A(n_172), .Y(n_817) );
XNOR2x1_ASAP7_75t_L g824 ( .A(n_173), .B(n_825), .Y(n_824) );
INVx1_ASAP7_75t_L g562 ( .A(n_174), .Y(n_562) );
AOI22xp33_ASAP7_75t_L g668 ( .A1(n_175), .A2(n_309), .B1(n_473), .B2(n_548), .Y(n_668) );
AO22x1_ASAP7_75t_L g1005 ( .A1(n_176), .A2(n_266), .B1(n_468), .B2(n_650), .Y(n_1005) );
AOI22xp33_ASAP7_75t_L g924 ( .A1(n_179), .A2(n_198), .B1(n_477), .B2(n_802), .Y(n_924) );
INVx1_ASAP7_75t_L g457 ( .A(n_180), .Y(n_457) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_180), .B(n_254), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_180), .B(n_462), .Y(n_534) );
NOR2xp33_ASAP7_75t_L g531 ( .A(n_181), .B(n_337), .Y(n_531) );
AND2x2_ASAP7_75t_L g1013 ( .A(n_183), .B(n_734), .Y(n_1013) );
AOI22xp33_ASAP7_75t_SL g1391 ( .A1(n_185), .A2(n_225), .B1(n_468), .B2(n_650), .Y(n_1391) );
AOI22xp33_ASAP7_75t_SL g1036 ( .A1(n_186), .A2(n_344), .B1(n_576), .B2(n_589), .Y(n_1036) );
AOI22xp33_ASAP7_75t_L g702 ( .A1(n_187), .A2(n_192), .B1(n_507), .B2(n_703), .Y(n_702) );
AOI21xp33_ASAP7_75t_L g955 ( .A1(n_190), .A2(n_581), .B(n_956), .Y(n_955) );
XNOR2x1_ASAP7_75t_L g874 ( .A(n_191), .B(n_875), .Y(n_874) );
CKINVDCx5p33_ASAP7_75t_R g1141 ( .A(n_195), .Y(n_1141) );
AOI22xp33_ASAP7_75t_L g1371 ( .A1(n_195), .A2(n_1372), .B1(n_1398), .B2(n_1400), .Y(n_1371) );
AOI22xp33_ASAP7_75t_L g503 ( .A1(n_196), .A2(n_324), .B1(n_504), .B2(n_507), .Y(n_503) );
AO22x1_ASAP7_75t_L g999 ( .A1(n_200), .A2(n_362), .B1(n_544), .B2(n_1000), .Y(n_999) );
AOI22xp33_ASAP7_75t_L g704 ( .A1(n_201), .A2(n_420), .B1(n_501), .B2(n_551), .Y(n_704) );
NAND2xp5_ASAP7_75t_L g565 ( .A(n_202), .B(n_566), .Y(n_565) );
AOI22xp5_ASAP7_75t_L g959 ( .A1(n_203), .A2(n_244), .B1(n_655), .B2(n_658), .Y(n_959) );
INVx1_ASAP7_75t_L g1355 ( .A(n_205), .Y(n_1355) );
NAND2xp5_ASAP7_75t_L g449 ( .A(n_206), .B(n_450), .Y(n_449) );
AOI22xp33_ASAP7_75t_SL g1087 ( .A1(n_208), .A2(n_391), .B1(n_655), .B2(n_1024), .Y(n_1087) );
AOI22xp5_ASAP7_75t_L g1086 ( .A1(n_209), .A2(n_396), .B1(n_860), .B2(n_885), .Y(n_1086) );
NAND2xp5_ASAP7_75t_L g907 ( .A(n_210), .B(n_626), .Y(n_907) );
AOI22xp5_ASAP7_75t_L g1084 ( .A1(n_211), .A2(n_359), .B1(n_736), .B2(n_795), .Y(n_1084) );
INVx1_ASAP7_75t_L g1356 ( .A(n_212), .Y(n_1356) );
AOI22xp5_ASAP7_75t_L g1392 ( .A1(n_213), .A2(n_300), .B1(n_800), .B2(n_802), .Y(n_1392) );
INVx1_ASAP7_75t_L g952 ( .A(n_215), .Y(n_952) );
INVx1_ASAP7_75t_L g842 ( .A(n_216), .Y(n_842) );
AOI22xp33_ASAP7_75t_L g884 ( .A1(n_217), .A2(n_317), .B1(n_795), .B2(n_885), .Y(n_884) );
AOI21xp33_ASAP7_75t_SL g869 ( .A1(n_219), .A2(n_551), .B(n_870), .Y(n_869) );
AOI22xp33_ASAP7_75t_L g669 ( .A1(n_220), .A2(n_372), .B1(n_634), .B2(n_670), .Y(n_669) );
AOI22xp33_ASAP7_75t_L g975 ( .A1(n_221), .A2(n_304), .B1(n_863), .B2(n_976), .Y(n_975) );
INVxp33_ASAP7_75t_SL g1143 ( .A(n_223), .Y(n_1143) );
INVx1_ASAP7_75t_L g1381 ( .A(n_226), .Y(n_1381) );
INVx1_ASAP7_75t_SL g624 ( .A(n_227), .Y(n_624) );
INVx1_ASAP7_75t_L g820 ( .A(n_228), .Y(n_820) );
AOI22xp33_ASAP7_75t_L g786 ( .A1(n_230), .A2(n_237), .B1(n_566), .B2(n_787), .Y(n_786) );
AOI221xp5_ASAP7_75t_L g1004 ( .A1(n_231), .A2(n_245), .B1(n_775), .B2(n_933), .C(n_1005), .Y(n_1004) );
INVx1_ASAP7_75t_L g610 ( .A(n_233), .Y(n_610) );
AOI22xp33_ASAP7_75t_L g1174 ( .A1(n_233), .A2(n_408), .B1(n_1124), .B2(n_1175), .Y(n_1174) );
AOI21xp5_ASAP7_75t_L g718 ( .A1(n_234), .A2(n_583), .B(n_719), .Y(n_718) );
INVx1_ASAP7_75t_L g1386 ( .A(n_235), .Y(n_1386) );
AOI22xp33_ASAP7_75t_L g832 ( .A1(n_236), .A2(n_397), .B1(n_468), .B2(n_473), .Y(n_832) );
AOI22xp33_ASAP7_75t_L g1078 ( .A1(n_239), .A2(n_419), .B1(n_863), .B2(n_976), .Y(n_1078) );
INVx1_ASAP7_75t_L g1066 ( .A(n_240), .Y(n_1066) );
AOI22xp33_ASAP7_75t_L g732 ( .A1(n_242), .A2(n_294), .B1(n_733), .B2(n_735), .Y(n_732) );
AOI21xp33_ASAP7_75t_L g1037 ( .A1(n_243), .A2(n_819), .B(n_1038), .Y(n_1037) );
INVx1_ASAP7_75t_L g966 ( .A(n_246), .Y(n_966) );
AOI22xp5_ASAP7_75t_L g636 ( .A1(n_247), .A2(n_350), .B1(n_637), .B2(n_640), .Y(n_636) );
AOI22xp33_ASAP7_75t_L g725 ( .A1(n_248), .A2(n_406), .B1(n_592), .B2(n_593), .Y(n_725) );
AOI22xp33_ASAP7_75t_SL g1373 ( .A1(n_249), .A2(n_1374), .B1(n_1396), .B2(n_1397), .Y(n_1373) );
INVx1_ASAP7_75t_L g1396 ( .A(n_249), .Y(n_1396) );
INVx1_ASAP7_75t_L g1063 ( .A(n_250), .Y(n_1063) );
AOI21x1_ASAP7_75t_SL g838 ( .A1(n_251), .A2(n_839), .B(n_841), .Y(n_838) );
INVx1_ASAP7_75t_L g720 ( .A(n_252), .Y(n_720) );
AOI22xp33_ASAP7_75t_L g866 ( .A1(n_253), .A2(n_302), .B1(n_867), .B2(n_868), .Y(n_866) );
INVx1_ASAP7_75t_L g440 ( .A(n_254), .Y(n_440) );
OAI22x1_ASAP7_75t_L g894 ( .A1(n_255), .A2(n_895), .B1(n_900), .B2(n_909), .Y(n_894) );
NAND5xp2_ASAP7_75t_SL g895 ( .A(n_255), .B(n_896), .C(n_897), .D(n_898), .E(n_899), .Y(n_895) );
AOI21xp5_ASAP7_75t_L g935 ( .A1(n_257), .A2(n_936), .B(n_938), .Y(n_935) );
AOI22xp5_ASAP7_75t_L g631 ( .A1(n_258), .A2(n_301), .B1(n_632), .B2(n_635), .Y(n_631) );
AOI22xp33_ASAP7_75t_L g1079 ( .A1(n_259), .A2(n_378), .B1(n_758), .B2(n_780), .Y(n_1079) );
AOI22xp33_ASAP7_75t_L g997 ( .A1(n_260), .A2(n_407), .B1(n_701), .B2(n_998), .Y(n_997) );
AOI22xp33_ASAP7_75t_L g467 ( .A1(n_261), .A2(n_412), .B1(n_468), .B2(n_473), .Y(n_467) );
AOI22xp33_ASAP7_75t_L g628 ( .A1(n_262), .A2(n_271), .B1(n_516), .B2(n_526), .Y(n_628) );
AOI22xp33_ASAP7_75t_L g1044 ( .A1(n_263), .A2(n_287), .B1(n_592), .B2(n_593), .Y(n_1044) );
AOI22xp33_ASAP7_75t_L g896 ( .A1(n_264), .A2(n_307), .B1(n_458), .B2(n_544), .Y(n_896) );
AOI22xp33_ASAP7_75t_L g960 ( .A1(n_265), .A2(n_389), .B1(n_491), .B2(n_860), .Y(n_960) );
INVx1_ASAP7_75t_L g844 ( .A(n_267), .Y(n_844) );
AOI22xp33_ASAP7_75t_L g1041 ( .A1(n_273), .A2(n_413), .B1(n_575), .B2(n_599), .Y(n_1041) );
AOI22xp33_ASAP7_75t_L g1071 ( .A1(n_274), .A2(n_280), .B1(n_701), .B2(n_976), .Y(n_1071) );
XNOR2x1_ASAP7_75t_L g1074 ( .A(n_277), .B(n_1075), .Y(n_1074) );
INVx1_ASAP7_75t_L g778 ( .A(n_278), .Y(n_778) );
XOR2x2_ASAP7_75t_L g1047 ( .A(n_279), .B(n_1048), .Y(n_1047) );
AOI22xp33_ASAP7_75t_L g574 ( .A1(n_281), .A2(n_293), .B1(n_575), .B2(n_576), .Y(n_574) );
INVx1_ASAP7_75t_L g699 ( .A(n_282), .Y(n_699) );
AOI22xp5_ASAP7_75t_L g1021 ( .A1(n_283), .A2(n_375), .B1(n_512), .B2(n_943), .Y(n_1021) );
AOI22xp5_ASAP7_75t_L g1023 ( .A1(n_284), .A2(n_402), .B1(n_546), .B2(n_1024), .Y(n_1023) );
AOI22xp33_ASAP7_75t_L g963 ( .A1(n_285), .A2(n_409), .B1(n_863), .B2(n_868), .Y(n_963) );
AOI22xp33_ASAP7_75t_L g723 ( .A1(n_286), .A2(n_390), .B1(n_575), .B2(n_595), .Y(n_723) );
AOI22xp5_ASAP7_75t_L g683 ( .A1(n_289), .A2(n_381), .B1(n_555), .B2(n_684), .Y(n_683) );
AOI22xp5_ASAP7_75t_L g793 ( .A1(n_290), .A2(n_383), .B1(n_473), .B2(n_794), .Y(n_793) );
AOI22xp33_ASAP7_75t_L g1126 ( .A1(n_291), .A2(n_403), .B1(n_1127), .B2(n_1128), .Y(n_1126) );
INVx1_ASAP7_75t_SL g656 ( .A(n_292), .Y(n_656) );
AOI22xp33_ASAP7_75t_L g666 ( .A1(n_295), .A2(n_322), .B1(n_433), .B2(n_667), .Y(n_666) );
INVx1_ASAP7_75t_L g890 ( .A(n_297), .Y(n_890) );
NAND2xp5_ASAP7_75t_L g864 ( .A(n_298), .B(n_697), .Y(n_864) );
NAND2xp5_ASAP7_75t_L g1016 ( .A(n_299), .B(n_1017), .Y(n_1016) );
AOI22xp33_ASAP7_75t_L g1364 ( .A1(n_305), .A2(n_374), .B1(n_489), .B2(n_544), .Y(n_1364) );
AOI22xp33_ASAP7_75t_L g790 ( .A1(n_306), .A2(n_345), .B1(n_646), .B2(n_791), .Y(n_790) );
INVx1_ASAP7_75t_L g428 ( .A(n_310), .Y(n_428) );
AOI22xp33_ASAP7_75t_L g715 ( .A1(n_311), .A2(n_361), .B1(n_579), .B2(n_589), .Y(n_715) );
INVx1_ASAP7_75t_L g1059 ( .A(n_312), .Y(n_1059) );
INVx1_ASAP7_75t_L g1350 ( .A(n_313), .Y(n_1350) );
AOI22xp5_ASAP7_75t_L g981 ( .A1(n_314), .A2(n_415), .B1(n_548), .B2(n_982), .Y(n_981) );
AOI22xp33_ASAP7_75t_L g543 ( .A1(n_315), .A2(n_332), .B1(n_458), .B2(n_544), .Y(n_543) );
AOI22xp33_ASAP7_75t_SL g756 ( .A1(n_318), .A2(n_351), .B1(n_757), .B2(n_759), .Y(n_756) );
AO22x1_ASAP7_75t_L g1153 ( .A1(n_320), .A2(n_328), .B1(n_1114), .B2(n_1128), .Y(n_1153) );
HB1xp67_ASAP7_75t_L g1097 ( .A(n_321), .Y(n_1097) );
AND2x4_ASAP7_75t_L g1108 ( .A(n_321), .B(n_1109), .Y(n_1108) );
AOI22xp33_ASAP7_75t_L g432 ( .A1(n_327), .A2(n_343), .B1(n_433), .B2(n_458), .Y(n_432) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_329), .B(n_511), .Y(n_510) );
AOI22xp5_ASAP7_75t_L g1025 ( .A1(n_330), .A2(n_382), .B1(n_634), .B2(n_879), .Y(n_1025) );
INVx1_ASAP7_75t_L g1057 ( .A(n_331), .Y(n_1057) );
INVx1_ASAP7_75t_L g1068 ( .A(n_334), .Y(n_1068) );
INVx1_ASAP7_75t_L g679 ( .A(n_335), .Y(n_679) );
AOI22xp33_ASAP7_75t_L g1055 ( .A1(n_336), .A2(n_338), .B1(n_828), .B2(n_829), .Y(n_1055) );
INVx1_ASAP7_75t_L g455 ( .A(n_337), .Y(n_455) );
INVxp67_ASAP7_75t_L g525 ( .A(n_337), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g972 ( .A(n_339), .B(n_695), .Y(n_972) );
INVx2_ASAP7_75t_L g1095 ( .A(n_347), .Y(n_1095) );
INVxp33_ASAP7_75t_SL g1222 ( .A(n_348), .Y(n_1222) );
INVx1_ASAP7_75t_L g1082 ( .A(n_353), .Y(n_1082) );
AOI22xp33_ASAP7_75t_L g545 ( .A1(n_358), .A2(n_376), .B1(n_489), .B2(n_546), .Y(n_545) );
OAI22x1_ASAP7_75t_L g803 ( .A1(n_360), .A2(n_804), .B1(n_805), .B2(n_821), .Y(n_803) );
INVx1_ASAP7_75t_L g821 ( .A(n_360), .Y(n_821) );
AOI221xp5_ASAP7_75t_L g886 ( .A1(n_366), .A2(n_392), .B1(n_867), .B2(n_887), .C(n_889), .Y(n_886) );
INVx1_ASAP7_75t_SL g648 ( .A(n_367), .Y(n_648) );
AO221x2_ASAP7_75t_L g1218 ( .A1(n_369), .A2(n_370), .B1(n_1175), .B2(n_1219), .C(n_1220), .Y(n_1218) );
CKINVDCx14_ASAP7_75t_R g990 ( .A(n_371), .Y(n_990) );
NAND2xp5_ASAP7_75t_L g1034 ( .A(n_373), .B(n_512), .Y(n_1034) );
INVx1_ASAP7_75t_L g686 ( .A(n_377), .Y(n_686) );
INVx1_ASAP7_75t_L g941 ( .A(n_379), .Y(n_941) );
AOI21xp33_ASAP7_75t_SL g745 ( .A1(n_380), .A2(n_746), .B(n_748), .Y(n_745) );
AOI22xp33_ASAP7_75t_L g588 ( .A1(n_384), .A2(n_416), .B1(n_589), .B2(n_590), .Y(n_588) );
INVx1_ASAP7_75t_L g905 ( .A(n_387), .Y(n_905) );
OAI22x1_ASAP7_75t_L g726 ( .A1(n_393), .A2(n_727), .B1(n_728), .B2(n_761), .Y(n_726) );
INVx1_ASAP7_75t_L g761 ( .A(n_393), .Y(n_761) );
AOI22x1_ASAP7_75t_L g763 ( .A1(n_393), .A2(n_727), .B1(n_728), .B2(n_761), .Y(n_763) );
INVx1_ASAP7_75t_L g1378 ( .A(n_395), .Y(n_1378) );
INVx1_ASAP7_75t_L g784 ( .A(n_405), .Y(n_784) );
CKINVDCx5p33_ASAP7_75t_R g652 ( .A(n_410), .Y(n_652) );
NAND2xp5_ASAP7_75t_L g716 ( .A(n_418), .B(n_717), .Y(n_716) );
XNOR2x1_ASAP7_75t_L g663 ( .A(n_421), .B(n_664), .Y(n_663) );
AOI21xp5_ASAP7_75t_L g422 ( .A1(n_423), .A2(n_1091), .B(n_1098), .Y(n_422) );
XNOR2xp5_ASAP7_75t_L g423 ( .A(n_424), .B(n_764), .Y(n_423) );
XNOR2x2_ASAP7_75t_SL g424 ( .A(n_425), .B(n_603), .Y(n_424) );
AOI22xp5_ASAP7_75t_L g425 ( .A1(n_426), .A2(n_536), .B1(n_601), .B2(n_602), .Y(n_425) );
INVx2_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
BUFx2_ASAP7_75t_L g601 ( .A(n_427), .Y(n_601) );
AO21x2_ASAP7_75t_L g427 ( .A1(n_428), .A2(n_429), .B(n_535), .Y(n_427) );
NOR3xp33_ASAP7_75t_SL g535 ( .A(n_428), .B(n_431), .C(n_495), .Y(n_535) );
NAND2xp5_ASAP7_75t_L g429 ( .A(n_430), .B(n_494), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
NAND4xp25_ASAP7_75t_SL g431 ( .A(n_432), .B(n_467), .C(n_476), .D(n_488), .Y(n_431) );
BUFx6f_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
BUFx6f_ASAP7_75t_L g544 ( .A(n_434), .Y(n_544) );
BUFx6f_ASAP7_75t_L g639 ( .A(n_434), .Y(n_639) );
BUFx6f_ASAP7_75t_L g885 ( .A(n_434), .Y(n_885) );
AND2x4_ASAP7_75t_L g434 ( .A(n_435), .B(n_446), .Y(n_434) );
AND2x4_ASAP7_75t_L g478 ( .A(n_435), .B(n_479), .Y(n_478) );
AND2x2_ASAP7_75t_L g485 ( .A(n_435), .B(n_486), .Y(n_485) );
AND2x4_ASAP7_75t_L g490 ( .A(n_435), .B(n_471), .Y(n_490) );
AND2x4_ASAP7_75t_L g575 ( .A(n_435), .B(n_475), .Y(n_575) );
AND2x4_ASAP7_75t_L g592 ( .A(n_435), .B(n_479), .Y(n_592) );
AND2x4_ASAP7_75t_L g593 ( .A(n_435), .B(n_486), .Y(n_593) );
AND2x4_ASAP7_75t_L g595 ( .A(n_435), .B(n_471), .Y(n_595) );
AND2x4_ASAP7_75t_L g435 ( .A(n_436), .B(n_444), .Y(n_435) );
AND2x2_ASAP7_75t_L g500 ( .A(n_436), .B(n_445), .Y(n_500) );
INVx1_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
AND2x2_ASAP7_75t_L g470 ( .A(n_437), .B(n_445), .Y(n_470) );
NAND2xp5_ASAP7_75t_L g437 ( .A(n_438), .B(n_441), .Y(n_437) );
NAND2xp33_ASAP7_75t_L g438 ( .A(n_439), .B(n_440), .Y(n_438) );
INVx2_ASAP7_75t_L g443 ( .A(n_439), .Y(n_443) );
INVx3_ASAP7_75t_L g450 ( .A(n_439), .Y(n_450) );
NAND2xp33_ASAP7_75t_L g456 ( .A(n_439), .B(n_457), .Y(n_456) );
INVx1_ASAP7_75t_L g466 ( .A(n_439), .Y(n_466) );
HB1xp67_ASAP7_75t_L g521 ( .A(n_439), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g463 ( .A(n_440), .B(n_464), .Y(n_463) );
NAND2xp5_ASAP7_75t_L g441 ( .A(n_442), .B(n_443), .Y(n_441) );
OAI21xp5_ASAP7_75t_L g524 ( .A1(n_442), .A2(n_466), .B(n_525), .Y(n_524) );
INVx1_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
AND2x2_ASAP7_75t_L g523 ( .A(n_445), .B(n_524), .Y(n_523) );
AND2x4_ASAP7_75t_L g459 ( .A(n_446), .B(n_460), .Y(n_459) );
AND2x4_ASAP7_75t_L g596 ( .A(n_446), .B(n_470), .Y(n_596) );
AND2x4_ASAP7_75t_L g599 ( .A(n_446), .B(n_460), .Y(n_599) );
INVx2_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
INVx2_ASAP7_75t_L g475 ( .A(n_447), .Y(n_475) );
OR2x2_ASAP7_75t_L g447 ( .A(n_448), .B(n_452), .Y(n_447) );
AND2x4_ASAP7_75t_L g471 ( .A(n_448), .B(n_472), .Y(n_471) );
AND2x4_ASAP7_75t_L g479 ( .A(n_448), .B(n_480), .Y(n_479) );
INVx2_ASAP7_75t_L g487 ( .A(n_448), .Y(n_487) );
AND2x2_ASAP7_75t_L g519 ( .A(n_448), .B(n_520), .Y(n_519) );
AND2x4_ASAP7_75t_L g448 ( .A(n_449), .B(n_451), .Y(n_448) );
NAND2xp5_ASAP7_75t_L g454 ( .A(n_450), .B(n_455), .Y(n_454) );
INVxp67_ASAP7_75t_L g462 ( .A(n_450), .Y(n_462) );
NAND3xp33_ASAP7_75t_L g533 ( .A(n_451), .B(n_461), .C(n_534), .Y(n_533) );
INVx1_ASAP7_75t_L g472 ( .A(n_452), .Y(n_472) );
INVx1_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
INVx1_ASAP7_75t_L g480 ( .A(n_453), .Y(n_480) );
AND2x2_ASAP7_75t_L g453 ( .A(n_454), .B(n_456), .Y(n_453) );
BUFx3_ASAP7_75t_L g731 ( .A(n_458), .Y(n_731) );
BUFx12f_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
INVx6_ASAP7_75t_L g643 ( .A(n_459), .Y(n_643) );
AND2x4_ASAP7_75t_L g493 ( .A(n_460), .B(n_471), .Y(n_493) );
AND2x4_ASAP7_75t_L g502 ( .A(n_460), .B(n_486), .Y(n_502) );
AND2x4_ASAP7_75t_L g579 ( .A(n_460), .B(n_486), .Y(n_579) );
AND2x4_ASAP7_75t_L g598 ( .A(n_460), .B(n_471), .Y(n_598) );
AND2x2_ASAP7_75t_L g460 ( .A(n_461), .B(n_465), .Y(n_460) );
NAND2xp5_ASAP7_75t_L g461 ( .A(n_462), .B(n_463), .Y(n_461) );
BUFx8_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
BUFx6f_ASAP7_75t_L g548 ( .A(n_469), .Y(n_548) );
AND2x2_ASAP7_75t_L g469 ( .A(n_470), .B(n_471), .Y(n_469) );
AND2x4_ASAP7_75t_L g474 ( .A(n_470), .B(n_475), .Y(n_474) );
AND2x2_ASAP7_75t_L g509 ( .A(n_470), .B(n_479), .Y(n_509) );
AND2x2_ASAP7_75t_L g514 ( .A(n_470), .B(n_486), .Y(n_514) );
AND2x4_ASAP7_75t_L g578 ( .A(n_470), .B(n_479), .Y(n_578) );
AND2x2_ASAP7_75t_L g583 ( .A(n_470), .B(n_486), .Y(n_583) );
AND2x4_ASAP7_75t_L g590 ( .A(n_470), .B(n_471), .Y(n_590) );
AND2x2_ASAP7_75t_L g734 ( .A(n_470), .B(n_471), .Y(n_734) );
BUFx6f_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
BUFx3_ASAP7_75t_L g650 ( .A(n_474), .Y(n_650) );
BUFx12f_ASAP7_75t_L g736 ( .A(n_474), .Y(n_736) );
BUFx6f_ASAP7_75t_L g879 ( .A(n_474), .Y(n_879) );
BUFx6f_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
BUFx12f_ASAP7_75t_L g655 ( .A(n_478), .Y(n_655) );
INVx3_ASAP7_75t_L g673 ( .A(n_478), .Y(n_673) );
AND2x4_ASAP7_75t_L g506 ( .A(n_479), .B(n_500), .Y(n_506) );
AND2x4_ASAP7_75t_L g589 ( .A(n_479), .B(n_500), .Y(n_589) );
AND2x4_ASAP7_75t_L g486 ( .A(n_480), .B(n_487), .Y(n_486) );
INVx1_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
INVx1_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
BUFx6f_ASAP7_75t_L g802 ( .A(n_483), .Y(n_802) );
INVx2_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
INVx1_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
BUFx5_ASAP7_75t_L g542 ( .A(n_485), .Y(n_542) );
BUFx6f_ASAP7_75t_L g658 ( .A(n_485), .Y(n_658) );
BUFx3_ASAP7_75t_L g1024 ( .A(n_485), .Y(n_1024) );
AND2x4_ASAP7_75t_L g499 ( .A(n_486), .B(n_500), .Y(n_499) );
AND2x2_ASAP7_75t_L g819 ( .A(n_486), .B(n_500), .Y(n_819) );
BUFx6f_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
BUFx12f_ASAP7_75t_L g634 ( .A(n_490), .Y(n_634) );
BUFx6f_ASAP7_75t_L g860 ( .A(n_490), .Y(n_860) );
INVx4_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
INVx4_ASAP7_75t_L g546 ( .A(n_492), .Y(n_546) );
INVx4_ASAP7_75t_L g635 ( .A(n_492), .Y(n_635) );
INVx2_ASAP7_75t_SL g670 ( .A(n_492), .Y(n_670) );
INVx2_ASAP7_75t_L g743 ( .A(n_492), .Y(n_743) );
INVx1_ASAP7_75t_L g792 ( .A(n_492), .Y(n_792) );
INVx1_ASAP7_75t_L g829 ( .A(n_492), .Y(n_829) );
INVx2_ASAP7_75t_L g982 ( .A(n_492), .Y(n_982) );
INVx8_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
INVx1_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
NAND4xp25_ASAP7_75t_L g495 ( .A(n_496), .B(n_503), .C(n_510), .D(n_515), .Y(n_495) );
INVx2_ASAP7_75t_L g620 ( .A(n_497), .Y(n_620) );
INVx2_ASAP7_75t_SL g497 ( .A(n_498), .Y(n_497) );
INVx2_ASAP7_75t_SL g867 ( .A(n_498), .Y(n_867) );
INVx2_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
BUFx8_ASAP7_75t_SL g554 ( .A(n_499), .Y(n_554) );
BUFx6f_ASAP7_75t_L g581 ( .A(n_499), .Y(n_581) );
INVx2_ASAP7_75t_L g696 ( .A(n_499), .Y(n_696) );
BUFx6f_ASAP7_75t_L g717 ( .A(n_499), .Y(n_717) );
BUFx3_ASAP7_75t_L g1017 ( .A(n_499), .Y(n_1017) );
INVx4_ASAP7_75t_L g622 ( .A(n_501), .Y(n_622) );
BUFx3_ASAP7_75t_L g755 ( .A(n_501), .Y(n_755) );
BUFx6f_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
INVx3_ASAP7_75t_L g556 ( .A(n_502), .Y(n_556) );
BUFx6f_ASAP7_75t_L g780 ( .A(n_502), .Y(n_780) );
INVx2_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
INVx2_ASAP7_75t_L g974 ( .A(n_505), .Y(n_974) );
INVx1_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
BUFx6f_ASAP7_75t_L g551 ( .A(n_506), .Y(n_551) );
BUFx3_ASAP7_75t_L g758 ( .A(n_506), .Y(n_758) );
BUFx3_ASAP7_75t_L g776 ( .A(n_506), .Y(n_776) );
INVx2_ASAP7_75t_L g1379 ( .A(n_507), .Y(n_1379) );
INVx1_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
BUFx6f_ASAP7_75t_L g617 ( .A(n_508), .Y(n_617) );
INVx2_ASAP7_75t_L g934 ( .A(n_508), .Y(n_934) );
INVx2_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
BUFx3_ASAP7_75t_L g552 ( .A(n_509), .Y(n_552) );
BUFx6f_ASAP7_75t_L g863 ( .A(n_509), .Y(n_863) );
BUFx3_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
INVx2_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
BUFx6f_ASAP7_75t_L g627 ( .A(n_513), .Y(n_627) );
INVx2_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
BUFx3_ASAP7_75t_L g560 ( .A(n_514), .Y(n_560) );
INVx3_ASAP7_75t_L g677 ( .A(n_514), .Y(n_677) );
INVx4_ASAP7_75t_L g516 ( .A(n_517), .Y(n_516) );
INVx2_ASAP7_75t_L g703 ( .A(n_517), .Y(n_703) );
INVx2_ASAP7_75t_L g787 ( .A(n_517), .Y(n_787) );
INVx3_ASAP7_75t_L g998 ( .A(n_517), .Y(n_998) );
INVx2_ASAP7_75t_L g1353 ( .A(n_517), .Y(n_1353) );
INVx5_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
BUFx4f_ASAP7_75t_L g751 ( .A(n_518), .Y(n_751) );
BUFx2_ASAP7_75t_L g940 ( .A(n_518), .Y(n_940) );
BUFx2_ASAP7_75t_L g976 ( .A(n_518), .Y(n_976) );
AND2x4_ASAP7_75t_L g518 ( .A(n_519), .B(n_523), .Y(n_518) );
AND2x4_ASAP7_75t_L g564 ( .A(n_519), .B(n_523), .Y(n_564) );
AND2x2_ASAP7_75t_L g576 ( .A(n_519), .B(n_523), .Y(n_576) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_521), .B(n_522), .Y(n_520) );
INVx1_ASAP7_75t_L g529 ( .A(n_521), .Y(n_529) );
INVx2_ASAP7_75t_SL g845 ( .A(n_526), .Y(n_845) );
INVx2_ASAP7_75t_SL g526 ( .A(n_527), .Y(n_526) );
INVx2_ASAP7_75t_L g681 ( .A(n_527), .Y(n_681) );
NOR2xp33_ASAP7_75t_L g719 ( .A(n_527), .B(n_720), .Y(n_719) );
BUFx6f_ASAP7_75t_L g872 ( .A(n_527), .Y(n_872) );
BUFx6f_ASAP7_75t_L g891 ( .A(n_527), .Y(n_891) );
INVx1_ASAP7_75t_L g971 ( .A(n_527), .Y(n_971) );
BUFx6f_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
INVx3_ASAP7_75t_L g568 ( .A(n_528), .Y(n_568) );
AO21x2_ASAP7_75t_L g528 ( .A1(n_529), .A2(n_530), .B(n_533), .Y(n_528) );
HB1xp67_ASAP7_75t_L g1096 ( .A(n_530), .Y(n_1096) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_531), .B(n_532), .Y(n_530) );
INVx2_ASAP7_75t_L g602 ( .A(n_536), .Y(n_602) );
OA22x2_ASAP7_75t_L g536 ( .A1(n_537), .A2(n_569), .B1(n_570), .B2(n_600), .Y(n_536) );
INVx1_ASAP7_75t_L g600 ( .A(n_537), .Y(n_600) );
XNOR2x1_ASAP7_75t_L g537 ( .A(n_538), .B(n_539), .Y(n_537) );
NOR2x1_ASAP7_75t_L g539 ( .A(n_540), .B(n_549), .Y(n_539) );
NAND4xp25_ASAP7_75t_L g540 ( .A(n_541), .B(n_543), .C(n_545), .D(n_547), .Y(n_540) );
BUFx3_ASAP7_75t_L g646 ( .A(n_548), .Y(n_646) );
NAND3xp33_ASAP7_75t_L g549 ( .A(n_550), .B(n_553), .C(n_557), .Y(n_549) );
INVx4_ASAP7_75t_L g613 ( .A(n_551), .Y(n_613) );
INVx2_ASAP7_75t_L g760 ( .A(n_552), .Y(n_760) );
INVx3_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
INVx2_ASAP7_75t_L g868 ( .A(n_556), .Y(n_868) );
INVx2_ASAP7_75t_L g1384 ( .A(n_556), .Y(n_1384) );
INVx1_ASAP7_75t_L g1351 ( .A(n_558), .Y(n_1351) );
INVx2_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
INVx2_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
BUFx3_ASAP7_75t_L g747 ( .A(n_560), .Y(n_747) );
INVx1_ASAP7_75t_L g937 ( .A(n_560), .Y(n_937) );
OAI21xp5_ASAP7_75t_L g561 ( .A1(n_562), .A2(n_563), .B(n_565), .Y(n_561) );
INVx4_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
INVx4_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
NOR2xp33_ASAP7_75t_L g816 ( .A(n_567), .B(n_817), .Y(n_816) );
INVx3_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
INVx4_ASAP7_75t_L g586 ( .A(n_568), .Y(n_586) );
INVx1_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
INVx1_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
OAI22xp5_ASAP7_75t_L g708 ( .A1(n_571), .A2(n_709), .B1(n_710), .B2(n_711), .Y(n_708) );
INVx1_ASAP7_75t_SL g709 ( .A(n_571), .Y(n_709) );
NOR2x1_ASAP7_75t_L g572 ( .A(n_573), .B(n_587), .Y(n_572) );
NAND4xp25_ASAP7_75t_L g573 ( .A(n_574), .B(n_577), .C(n_580), .D(n_582), .Y(n_573) );
BUFx3_ASAP7_75t_L g929 ( .A(n_581), .Y(n_929) );
INVx2_ASAP7_75t_L g888 ( .A(n_583), .Y(n_888) );
NOR2xp33_ASAP7_75t_L g584 ( .A(n_585), .B(n_586), .Y(n_584) );
INVx4_ASAP7_75t_L g701 ( .A(n_586), .Y(n_701) );
NOR2xp33_ASAP7_75t_L g904 ( .A(n_586), .B(n_905), .Y(n_904) );
NOR2xp33_ASAP7_75t_L g1038 ( .A(n_586), .B(n_1039), .Y(n_1038) );
NAND4xp25_ASAP7_75t_L g587 ( .A(n_588), .B(n_591), .C(n_594), .D(n_597), .Y(n_587) );
XNOR2xp5_ASAP7_75t_L g603 ( .A(n_604), .B(n_705), .Y(n_603) );
INVx1_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
OA22x2_ASAP7_75t_L g605 ( .A1(n_606), .A2(n_607), .B1(n_661), .B2(n_662), .Y(n_605) );
INVx4_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
AO22x2_ASAP7_75t_L g607 ( .A1(n_608), .A2(n_609), .B1(n_629), .B2(n_659), .Y(n_607) );
NOR4xp25_ASAP7_75t_L g608 ( .A(n_609), .B(n_611), .C(n_618), .D(n_623), .Y(n_608) );
CKINVDCx5p33_ASAP7_75t_R g609 ( .A(n_610), .Y(n_609) );
NOR3xp33_ASAP7_75t_SL g660 ( .A(n_611), .B(n_618), .C(n_623), .Y(n_660) );
OAI22xp33_ASAP7_75t_L g611 ( .A1(n_612), .A2(n_613), .B1(n_614), .B2(n_615), .Y(n_611) );
OAI22xp5_ASAP7_75t_L g1061 ( .A1(n_613), .A2(n_1062), .B1(n_1063), .B2(n_1064), .Y(n_1061) );
OAI22xp5_ASAP7_75t_L g1357 ( .A1(n_613), .A2(n_1358), .B1(n_1359), .B2(n_1360), .Y(n_1357) );
INVx1_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
INVx2_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
INVx2_ASAP7_75t_L g684 ( .A(n_617), .Y(n_684) );
INVx2_ASAP7_75t_L g774 ( .A(n_617), .Y(n_774) );
INVx1_ASAP7_75t_L g1361 ( .A(n_617), .Y(n_1361) );
OAI22xp33_ASAP7_75t_L g618 ( .A1(n_619), .A2(n_620), .B1(n_621), .B2(n_622), .Y(n_618) );
OAI22xp5_ASAP7_75t_L g1065 ( .A1(n_622), .A2(n_1066), .B1(n_1067), .B2(n_1068), .Y(n_1065) );
OAI22xp33_ASAP7_75t_L g1354 ( .A1(n_622), .A2(n_1067), .B1(n_1355), .B2(n_1356), .Y(n_1354) );
OAI21xp33_ASAP7_75t_L g623 ( .A1(n_624), .A2(n_625), .B(n_628), .Y(n_623) );
INVx1_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
INVx2_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
INVx1_ASAP7_75t_L g840 ( .A(n_627), .Y(n_840) );
INVx2_ASAP7_75t_L g954 ( .A(n_627), .Y(n_954) );
NAND2xp5_ASAP7_75t_SL g659 ( .A(n_629), .B(n_660), .Y(n_659) );
NOR3xp33_ASAP7_75t_L g629 ( .A(n_630), .B(n_644), .C(n_651), .Y(n_629) );
NAND2xp5_ASAP7_75t_L g630 ( .A(n_631), .B(n_636), .Y(n_630) );
INVx1_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
INVx1_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
BUFx6f_ASAP7_75t_L g741 ( .A(n_634), .Y(n_741) );
BUFx12f_ASAP7_75t_L g828 ( .A(n_634), .Y(n_828) );
INVx1_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
INVx1_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
BUFx3_ASAP7_75t_L g798 ( .A(n_639), .Y(n_798) );
INVx1_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
INVx1_ASAP7_75t_L g641 ( .A(n_642), .Y(n_641) );
HB1xp67_ASAP7_75t_L g1052 ( .A(n_642), .Y(n_1052) );
INVx2_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
INVx3_ASAP7_75t_L g667 ( .A(n_643), .Y(n_667) );
INVx5_ASAP7_75t_L g795 ( .A(n_643), .Y(n_795) );
INVx1_ASAP7_75t_L g855 ( .A(n_643), .Y(n_855) );
INVx1_ASAP7_75t_L g1000 ( .A(n_643), .Y(n_1000) );
OAI22xp5_ASAP7_75t_L g644 ( .A1(n_645), .A2(n_647), .B1(n_648), .B2(n_649), .Y(n_644) );
INVx1_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
OAI22xp5_ASAP7_75t_L g1056 ( .A1(n_649), .A2(n_1057), .B1(n_1058), .B2(n_1059), .Y(n_1056) );
INVx1_ASAP7_75t_L g649 ( .A(n_650), .Y(n_649) );
OAI22x1_ASAP7_75t_SL g651 ( .A1(n_652), .A2(n_653), .B1(n_656), .B2(n_657), .Y(n_651) );
INVx1_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
HB1xp67_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
INVx1_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
BUFx2_ASAP7_75t_SL g739 ( .A(n_658), .Y(n_739) );
INVx1_ASAP7_75t_SL g661 ( .A(n_662), .Y(n_661) );
XNOR2xp5_ASAP7_75t_L g662 ( .A(n_663), .B(n_685), .Y(n_662) );
NOR2x1_ASAP7_75t_L g664 ( .A(n_665), .B(n_674), .Y(n_664) );
NAND4xp25_ASAP7_75t_L g665 ( .A(n_666), .B(n_668), .C(n_669), .D(n_671), .Y(n_665) );
INVx1_ASAP7_75t_L g672 ( .A(n_673), .Y(n_672) );
INVx1_ASAP7_75t_L g738 ( .A(n_673), .Y(n_738) );
INVx2_ASAP7_75t_L g801 ( .A(n_673), .Y(n_801) );
NAND3xp33_ASAP7_75t_L g674 ( .A(n_675), .B(n_682), .C(n_683), .Y(n_674) );
INVx2_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
INVx3_ASAP7_75t_SL g697 ( .A(n_677), .Y(n_697) );
INVx2_ASAP7_75t_L g970 ( .A(n_677), .Y(n_970) );
INVx2_ASAP7_75t_L g994 ( .A(n_677), .Y(n_994) );
NOR2xp33_ASAP7_75t_L g678 ( .A(n_679), .B(n_680), .Y(n_678) );
NOR2xp33_ASAP7_75t_L g956 ( .A(n_680), .B(n_957), .Y(n_956) );
INVx3_ASAP7_75t_L g680 ( .A(n_681), .Y(n_680) );
INVx2_ASAP7_75t_L g707 ( .A(n_685), .Y(n_707) );
XNOR2x1_ASAP7_75t_L g685 ( .A(n_686), .B(n_687), .Y(n_685) );
NOR2x1_ASAP7_75t_L g687 ( .A(n_688), .B(n_693), .Y(n_687) );
NAND4xp25_ASAP7_75t_L g688 ( .A(n_689), .B(n_690), .C(n_691), .D(n_692), .Y(n_688) );
NAND3xp33_ASAP7_75t_L g693 ( .A(n_694), .B(n_702), .C(n_704), .Y(n_693) );
INVx2_ASAP7_75t_L g782 ( .A(n_695), .Y(n_782) );
INVx3_ASAP7_75t_L g695 ( .A(n_696), .Y(n_695) );
INVx2_ASAP7_75t_L g837 ( .A(n_696), .Y(n_837) );
INVx1_ASAP7_75t_L g785 ( .A(n_697), .Y(n_785) );
NOR2xp33_ASAP7_75t_L g698 ( .A(n_699), .B(n_700), .Y(n_698) );
INVx2_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
INVx1_ASAP7_75t_L g843 ( .A(n_703), .Y(n_843) );
AO22x2_ASAP7_75t_L g705 ( .A1(n_706), .A2(n_726), .B1(n_762), .B2(n_763), .Y(n_705) );
INVx1_ASAP7_75t_L g762 ( .A(n_706), .Y(n_762) );
XNOR2xp5_ASAP7_75t_L g706 ( .A(n_707), .B(n_708), .Y(n_706) );
INVx2_ASAP7_75t_L g710 ( .A(n_711), .Y(n_710) );
OR2x2_ASAP7_75t_L g712 ( .A(n_713), .B(n_721), .Y(n_712) );
NAND4xp25_ASAP7_75t_L g713 ( .A(n_714), .B(n_715), .C(n_716), .D(n_718), .Y(n_713) );
BUFx3_ASAP7_75t_L g754 ( .A(n_717), .Y(n_754) );
NAND4xp25_ASAP7_75t_L g721 ( .A(n_722), .B(n_723), .C(n_724), .D(n_725), .Y(n_721) );
INVx2_ASAP7_75t_L g727 ( .A(n_728), .Y(n_727) );
OR2x2_ASAP7_75t_L g728 ( .A(n_729), .B(n_744), .Y(n_728) );
NAND4xp25_ASAP7_75t_SL g729 ( .A(n_730), .B(n_732), .C(n_737), .D(n_740), .Y(n_729) );
INVxp67_ASAP7_75t_L g1058 ( .A(n_733), .Y(n_1058) );
BUFx6f_ASAP7_75t_L g733 ( .A(n_734), .Y(n_733) );
BUFx4f_ASAP7_75t_L g878 ( .A(n_734), .Y(n_878) );
BUFx3_ASAP7_75t_L g735 ( .A(n_736), .Y(n_735) );
BUFx2_ASAP7_75t_SL g742 ( .A(n_743), .Y(n_742) );
NAND3xp33_ASAP7_75t_L g744 ( .A(n_745), .B(n_753), .C(n_756), .Y(n_744) );
HB1xp67_ASAP7_75t_L g746 ( .A(n_747), .Y(n_746) );
OAI21xp33_ASAP7_75t_L g748 ( .A1(n_749), .A2(n_750), .B(n_752), .Y(n_748) );
INVx2_ASAP7_75t_SL g750 ( .A(n_751), .Y(n_750) );
BUFx2_ASAP7_75t_L g757 ( .A(n_758), .Y(n_757) );
INVx2_ASAP7_75t_L g759 ( .A(n_760), .Y(n_759) );
XNOR2xp5_ASAP7_75t_L g764 ( .A(n_765), .B(n_914), .Y(n_764) );
AOI22xp5_ASAP7_75t_L g765 ( .A1(n_766), .A2(n_767), .B1(n_848), .B2(n_913), .Y(n_765) );
INVx2_ASAP7_75t_L g766 ( .A(n_767), .Y(n_766) );
OAI21xp5_ASAP7_75t_L g767 ( .A1(n_768), .A2(n_822), .B(n_846), .Y(n_767) );
NAND2xp5_ASAP7_75t_L g846 ( .A(n_768), .B(n_847), .Y(n_846) );
INVx1_ASAP7_75t_L g768 ( .A(n_769), .Y(n_768) );
XNOR2xp5_ASAP7_75t_L g769 ( .A(n_770), .B(n_803), .Y(n_769) );
INVx2_ASAP7_75t_L g770 ( .A(n_771), .Y(n_770) );
AND2x4_ASAP7_75t_L g771 ( .A(n_772), .B(n_788), .Y(n_771) );
NOR3xp33_ASAP7_75t_L g772 ( .A(n_773), .B(n_777), .C(n_783), .Y(n_772) );
INVxp67_ASAP7_75t_L g1064 ( .A(n_774), .Y(n_1064) );
HB1xp67_ASAP7_75t_L g775 ( .A(n_776), .Y(n_775) );
INVx2_ASAP7_75t_L g932 ( .A(n_776), .Y(n_932) );
OAI22xp5_ASAP7_75t_L g777 ( .A1(n_778), .A2(n_779), .B1(n_781), .B2(n_782), .Y(n_777) );
INVx3_ASAP7_75t_L g779 ( .A(n_780), .Y(n_779) );
OAI22xp5_ASAP7_75t_L g1380 ( .A1(n_782), .A2(n_1381), .B1(n_1382), .B2(n_1383), .Y(n_1380) );
OAI21xp33_ASAP7_75t_L g783 ( .A1(n_784), .A2(n_785), .B(n_786), .Y(n_783) );
OAI21xp33_ASAP7_75t_L g1069 ( .A1(n_785), .A2(n_1070), .B(n_1071), .Y(n_1069) );
NOR2x1_ASAP7_75t_L g788 ( .A(n_789), .B(n_796), .Y(n_788) );
NAND2xp5_ASAP7_75t_L g789 ( .A(n_790), .B(n_793), .Y(n_789) );
BUFx2_ASAP7_75t_L g791 ( .A(n_792), .Y(n_791) );
HB1xp67_ASAP7_75t_L g794 ( .A(n_795), .Y(n_794) );
NAND2xp5_ASAP7_75t_L g796 ( .A(n_797), .B(n_799), .Y(n_796) );
BUFx4f_ASAP7_75t_L g800 ( .A(n_801), .Y(n_800) );
INVx2_ASAP7_75t_L g804 ( .A(n_805), .Y(n_804) );
XOR2x2_ASAP7_75t_L g805 ( .A(n_806), .B(n_820), .Y(n_805) );
NOR2xp67_ASAP7_75t_L g806 ( .A(n_807), .B(n_812), .Y(n_806) );
NAND4xp25_ASAP7_75t_L g807 ( .A(n_808), .B(n_809), .C(n_810), .D(n_811), .Y(n_807) );
NAND4xp25_ASAP7_75t_L g812 ( .A(n_813), .B(n_814), .C(n_815), .D(n_818), .Y(n_812) );
INVx1_ASAP7_75t_L g822 ( .A(n_823), .Y(n_822) );
BUFx3_ASAP7_75t_L g823 ( .A(n_824), .Y(n_823) );
INVx1_ASAP7_75t_L g847 ( .A(n_824), .Y(n_847) );
NAND4xp75_ASAP7_75t_SL g825 ( .A(n_826), .B(n_831), .C(n_834), .D(n_838), .Y(n_825) );
AND2x2_ASAP7_75t_L g826 ( .A(n_827), .B(n_830), .Y(n_826) );
AND2x2_ASAP7_75t_L g831 ( .A(n_832), .B(n_833), .Y(n_831) );
AND2x2_ASAP7_75t_L g834 ( .A(n_835), .B(n_836), .Y(n_834) );
HB1xp67_ASAP7_75t_L g839 ( .A(n_840), .Y(n_839) );
OAI22xp5_ASAP7_75t_L g841 ( .A1(n_842), .A2(n_843), .B1(n_844), .B2(n_845), .Y(n_841) );
HB1xp67_ASAP7_75t_L g848 ( .A(n_849), .Y(n_848) );
INVx2_ASAP7_75t_L g913 ( .A(n_849), .Y(n_913) );
XNOR2x1_ASAP7_75t_L g849 ( .A(n_850), .B(n_893), .Y(n_849) );
XNOR2xp5_ASAP7_75t_L g850 ( .A(n_851), .B(n_874), .Y(n_850) );
XNOR2x1_ASAP7_75t_L g851 ( .A(n_852), .B(n_873), .Y(n_851) );
NOR4xp75_ASAP7_75t_L g852 ( .A(n_853), .B(n_857), .C(n_861), .D(n_865), .Y(n_852) );
NAND2xp5_ASAP7_75t_L g853 ( .A(n_854), .B(n_856), .Y(n_853) );
NAND2xp5_ASAP7_75t_L g857 ( .A(n_858), .B(n_859), .Y(n_857) );
NAND2xp5_ASAP7_75t_L g861 ( .A(n_862), .B(n_864), .Y(n_861) );
NAND2xp5_ASAP7_75t_SL g865 ( .A(n_866), .B(n_869), .Y(n_865) );
NOR2xp33_ASAP7_75t_L g870 ( .A(n_871), .B(n_872), .Y(n_870) );
INVx2_ASAP7_75t_L g943 ( .A(n_872), .Y(n_943) );
NOR2x1_ASAP7_75t_L g875 ( .A(n_876), .B(n_883), .Y(n_875) );
NAND4xp25_ASAP7_75t_L g876 ( .A(n_877), .B(n_880), .C(n_881), .D(n_882), .Y(n_876) );
NAND3xp33_ASAP7_75t_L g883 ( .A(n_884), .B(n_886), .C(n_892), .Y(n_883) );
BUFx3_ASAP7_75t_L g1051 ( .A(n_885), .Y(n_1051) );
INVx2_ASAP7_75t_L g887 ( .A(n_888), .Y(n_887) );
NOR2xp33_ASAP7_75t_L g889 ( .A(n_890), .B(n_891), .Y(n_889) );
NOR2xp33_ASAP7_75t_L g1081 ( .A(n_891), .B(n_1082), .Y(n_1081) );
BUFx3_ASAP7_75t_L g893 ( .A(n_894), .Y(n_893) );
NAND4xp25_ASAP7_75t_L g910 ( .A(n_896), .B(n_897), .C(n_899), .D(n_907), .Y(n_910) );
NAND2xp5_ASAP7_75t_L g912 ( .A(n_898), .B(n_908), .Y(n_912) );
NAND3xp33_ASAP7_75t_L g900 ( .A(n_901), .B(n_907), .C(n_908), .Y(n_900) );
INVxp67_ASAP7_75t_L g901 ( .A(n_902), .Y(n_901) );
OR2x2_ASAP7_75t_L g911 ( .A(n_902), .B(n_912), .Y(n_911) );
NAND2xp5_ASAP7_75t_L g902 ( .A(n_903), .B(n_906), .Y(n_902) );
NOR2x1_ASAP7_75t_L g909 ( .A(n_910), .B(n_911), .Y(n_909) );
OAI22xp5_ASAP7_75t_L g914 ( .A1(n_915), .A2(n_985), .B1(n_1089), .B2(n_1090), .Y(n_914) );
INVx1_ASAP7_75t_L g1090 ( .A(n_915), .Y(n_1090) );
HB1xp67_ASAP7_75t_L g915 ( .A(n_916), .Y(n_915) );
OA22x2_ASAP7_75t_L g916 ( .A1(n_917), .A2(n_945), .B1(n_983), .B2(n_984), .Y(n_916) );
INVx2_ASAP7_75t_L g984 ( .A(n_917), .Y(n_984) );
AO21x2_ASAP7_75t_L g917 ( .A1(n_918), .A2(n_919), .B(n_944), .Y(n_917) );
NOR3xp33_ASAP7_75t_L g944 ( .A(n_918), .B(n_921), .C(n_927), .Y(n_944) );
NAND2xp5_ASAP7_75t_L g919 ( .A(n_920), .B(n_926), .Y(n_919) );
INVx1_ASAP7_75t_L g920 ( .A(n_921), .Y(n_920) );
NAND4xp25_ASAP7_75t_SL g921 ( .A(n_922), .B(n_923), .C(n_924), .D(n_925), .Y(n_921) );
INVx1_ASAP7_75t_L g926 ( .A(n_927), .Y(n_926) );
NAND3xp33_ASAP7_75t_L g927 ( .A(n_928), .B(n_930), .C(n_935), .Y(n_927) );
INVx1_ASAP7_75t_L g1067 ( .A(n_929), .Y(n_1067) );
INVx2_ASAP7_75t_L g931 ( .A(n_932), .Y(n_931) );
OAI22xp5_ASAP7_75t_L g1376 ( .A1(n_932), .A2(n_1377), .B1(n_1378), .B2(n_1379), .Y(n_1376) );
BUFx3_ASAP7_75t_L g933 ( .A(n_934), .Y(n_933) );
INVx2_ASAP7_75t_L g936 ( .A(n_937), .Y(n_936) );
OAI21xp5_ASAP7_75t_SL g938 ( .A1(n_939), .A2(n_941), .B(n_942), .Y(n_938) );
INVxp67_ASAP7_75t_L g939 ( .A(n_940), .Y(n_939) );
INVx1_ASAP7_75t_L g983 ( .A(n_945), .Y(n_983) );
XNOR2xp5_ASAP7_75t_L g945 ( .A(n_946), .B(n_964), .Y(n_945) );
NAND4xp75_ASAP7_75t_L g947 ( .A(n_948), .B(n_951), .C(n_958), .D(n_961), .Y(n_947) );
AND2x2_ASAP7_75t_L g948 ( .A(n_949), .B(n_950), .Y(n_948) );
OA21x2_ASAP7_75t_L g951 ( .A1(n_952), .A2(n_953), .B(n_955), .Y(n_951) );
INVx1_ASAP7_75t_L g953 ( .A(n_954), .Y(n_953) );
AND2x2_ASAP7_75t_L g958 ( .A(n_959), .B(n_960), .Y(n_958) );
AND2x2_ASAP7_75t_L g961 ( .A(n_962), .B(n_963), .Y(n_961) );
XNOR2xp5_ASAP7_75t_L g964 ( .A(n_965), .B(n_967), .Y(n_964) );
CKINVDCx5p33_ASAP7_75t_R g965 ( .A(n_966), .Y(n_965) );
NOR2x1_ASAP7_75t_L g967 ( .A(n_968), .B(n_977), .Y(n_967) );
NAND4xp25_ASAP7_75t_L g968 ( .A(n_969), .B(n_972), .C(n_973), .D(n_975), .Y(n_968) );
INVx2_ASAP7_75t_L g1387 ( .A(n_970), .Y(n_1387) );
NAND4xp25_ASAP7_75t_L g977 ( .A(n_978), .B(n_979), .C(n_980), .D(n_981), .Y(n_977) );
INVx2_ASAP7_75t_L g1089 ( .A(n_985), .Y(n_1089) );
AO22x2_ASAP7_75t_L g985 ( .A1(n_986), .A2(n_987), .B1(n_1046), .B2(n_1088), .Y(n_985) );
INVx1_ASAP7_75t_L g986 ( .A(n_987), .Y(n_986) );
XNOR2x1_ASAP7_75t_L g987 ( .A(n_988), .B(n_1006), .Y(n_987) );
INVx2_ASAP7_75t_L g988 ( .A(n_989), .Y(n_988) );
XNOR2x2_ASAP7_75t_L g989 ( .A(n_990), .B(n_991), .Y(n_989) );
NAND3xp33_ASAP7_75t_L g991 ( .A(n_992), .B(n_1001), .C(n_1004), .Y(n_991) );
HB1xp67_ASAP7_75t_L g993 ( .A(n_994), .Y(n_993) );
NAND2xp5_ASAP7_75t_L g995 ( .A(n_996), .B(n_997), .Y(n_995) );
INVx1_ASAP7_75t_L g1002 ( .A(n_1003), .Y(n_1002) );
AO22x2_ASAP7_75t_L g1006 ( .A1(n_1007), .A2(n_1008), .B1(n_1029), .B2(n_1030), .Y(n_1006) );
INVx2_ASAP7_75t_SL g1007 ( .A(n_1008), .Y(n_1007) );
AO21x2_ASAP7_75t_L g1008 ( .A1(n_1009), .A2(n_1018), .B(n_1026), .Y(n_1008) );
NAND2xp5_ASAP7_75t_L g1010 ( .A(n_1011), .B(n_1012), .Y(n_1010) );
NAND2xp5_ASAP7_75t_SL g1014 ( .A(n_1015), .B(n_1016), .Y(n_1014) );
NOR2xp33_ASAP7_75t_L g1018 ( .A(n_1019), .B(n_1022), .Y(n_1018) );
NAND2xp5_ASAP7_75t_L g1019 ( .A(n_1020), .B(n_1021), .Y(n_1019) );
NAND2x1_ASAP7_75t_SL g1022 ( .A(n_1023), .B(n_1025), .Y(n_1022) );
NAND2xp5_ASAP7_75t_L g1026 ( .A(n_1027), .B(n_1028), .Y(n_1026) );
OA22x2_ASAP7_75t_L g1072 ( .A1(n_1029), .A2(n_1030), .B1(n_1073), .B2(n_1074), .Y(n_1072) );
INVx2_ASAP7_75t_L g1029 ( .A(n_1030), .Y(n_1029) );
AO21x2_ASAP7_75t_L g1030 ( .A1(n_1031), .A2(n_1032), .B(n_1045), .Y(n_1030) );
NOR3xp33_ASAP7_75t_SL g1045 ( .A(n_1031), .B(n_1033), .C(n_1040), .Y(n_1045) );
OR2x2_ASAP7_75t_L g1032 ( .A(n_1033), .B(n_1040), .Y(n_1032) );
NAND4xp75_ASAP7_75t_L g1033 ( .A(n_1034), .B(n_1035), .C(n_1036), .D(n_1037), .Y(n_1033) );
NAND4xp25_ASAP7_75t_L g1040 ( .A(n_1041), .B(n_1042), .C(n_1043), .D(n_1044), .Y(n_1040) );
INVx2_ASAP7_75t_L g1088 ( .A(n_1046), .Y(n_1088) );
XNOR2x1_ASAP7_75t_L g1046 ( .A(n_1047), .B(n_1072), .Y(n_1046) );
NAND2xp5_ASAP7_75t_L g1048 ( .A(n_1049), .B(n_1060), .Y(n_1048) );
NOR3xp33_ASAP7_75t_L g1049 ( .A(n_1050), .B(n_1053), .C(n_1056), .Y(n_1049) );
NAND2xp5_ASAP7_75t_L g1053 ( .A(n_1054), .B(n_1055), .Y(n_1053) );
NOR3xp33_ASAP7_75t_L g1060 ( .A(n_1061), .B(n_1065), .C(n_1069), .Y(n_1060) );
INVx2_ASAP7_75t_L g1073 ( .A(n_1074), .Y(n_1073) );
NOR2x1_ASAP7_75t_L g1075 ( .A(n_1076), .B(n_1083), .Y(n_1075) );
NAND4xp25_ASAP7_75t_L g1076 ( .A(n_1077), .B(n_1078), .C(n_1079), .D(n_1080), .Y(n_1076) );
NAND4xp25_ASAP7_75t_L g1083 ( .A(n_1084), .B(n_1085), .C(n_1086), .D(n_1087), .Y(n_1083) );
INVx2_ASAP7_75t_SL g1091 ( .A(n_1092), .Y(n_1091) );
NAND3xp33_ASAP7_75t_L g1092 ( .A(n_1093), .B(n_1096), .C(n_1097), .Y(n_1092) );
AND2x2_ASAP7_75t_L g1368 ( .A(n_1093), .B(n_1369), .Y(n_1368) );
AND2x2_ASAP7_75t_L g1399 ( .A(n_1093), .B(n_1370), .Y(n_1399) );
AOI21xp5_ASAP7_75t_L g1403 ( .A1(n_1093), .A2(n_1097), .B(n_1115), .Y(n_1403) );
INVx1_ASAP7_75t_L g1093 ( .A(n_1094), .Y(n_1093) );
AO21x1_ASAP7_75t_L g1401 ( .A1(n_1094), .A2(n_1402), .B(n_1403), .Y(n_1401) );
HB1xp67_ASAP7_75t_L g1094 ( .A(n_1095), .Y(n_1094) );
AND3x4_ASAP7_75t_L g1114 ( .A(n_1095), .B(n_1108), .C(n_1115), .Y(n_1114) );
AND2x2_ASAP7_75t_L g1117 ( .A(n_1095), .B(n_1118), .Y(n_1117) );
NOR2xp33_ASAP7_75t_L g1369 ( .A(n_1096), .B(n_1370), .Y(n_1369) );
INVx1_ASAP7_75t_L g1370 ( .A(n_1097), .Y(n_1370) );
OAI221xp5_ASAP7_75t_L g1098 ( .A1(n_1099), .A2(n_1342), .B1(n_1344), .B2(n_1367), .C(n_1371), .Y(n_1098) );
O2A1O1Ixp33_ASAP7_75t_SL g1099 ( .A1(n_1100), .A2(n_1223), .B(n_1247), .C(n_1313), .Y(n_1099) );
NAND5xp2_ASAP7_75t_L g1100 ( .A(n_1101), .B(n_1189), .C(n_1204), .D(n_1213), .E(n_1218), .Y(n_1100) );
AOI221xp5_ASAP7_75t_L g1101 ( .A1(n_1102), .A2(n_1149), .B1(n_1154), .B2(n_1162), .C(n_1165), .Y(n_1101) );
INVxp67_ASAP7_75t_SL g1102 ( .A(n_1103), .Y(n_1102) );
NAND2xp5_ASAP7_75t_L g1103 ( .A(n_1104), .B(n_1119), .Y(n_1103) );
NAND2xp5_ASAP7_75t_L g1251 ( .A(n_1104), .B(n_1252), .Y(n_1251) );
NAND2xp5_ASAP7_75t_L g1305 ( .A(n_1104), .B(n_1267), .Y(n_1305) );
HB1xp67_ASAP7_75t_L g1104 ( .A(n_1105), .Y(n_1104) );
NOR2xp33_ASAP7_75t_L g1184 ( .A(n_1105), .B(n_1132), .Y(n_1184) );
OR2x2_ASAP7_75t_L g1187 ( .A(n_1105), .B(n_1151), .Y(n_1187) );
CKINVDCx5p33_ASAP7_75t_R g1199 ( .A(n_1105), .Y(n_1199) );
HB1xp67_ASAP7_75t_L g1207 ( .A(n_1105), .Y(n_1207) );
NAND2xp5_ASAP7_75t_L g1217 ( .A(n_1105), .B(n_1193), .Y(n_1217) );
BUFx2_ASAP7_75t_L g1231 ( .A(n_1105), .Y(n_1231) );
NAND2xp5_ASAP7_75t_L g1234 ( .A(n_1105), .B(n_1132), .Y(n_1234) );
NOR2xp33_ASAP7_75t_L g1266 ( .A(n_1105), .B(n_1239), .Y(n_1266) );
AND2x2_ASAP7_75t_L g1285 ( .A(n_1105), .B(n_1151), .Y(n_1285) );
AND2x4_ASAP7_75t_L g1105 ( .A(n_1106), .B(n_1113), .Y(n_1105) );
AND2x4_ASAP7_75t_L g1107 ( .A(n_1108), .B(n_1110), .Y(n_1107) );
AND2x4_ASAP7_75t_L g1127 ( .A(n_1108), .B(n_1117), .Y(n_1127) );
NAND2xp5_ASAP7_75t_L g1142 ( .A(n_1108), .B(n_1110), .Y(n_1142) );
AND2x4_ASAP7_75t_L g1177 ( .A(n_1108), .B(n_1110), .Y(n_1177) );
AND2x2_ASAP7_75t_L g1111 ( .A(n_1110), .B(n_1112), .Y(n_1111) );
AND2x4_ASAP7_75t_L g1124 ( .A(n_1110), .B(n_1112), .Y(n_1124) );
AND2x2_ASAP7_75t_L g1147 ( .A(n_1110), .B(n_1112), .Y(n_1147) );
AND2x2_ASAP7_75t_L g1116 ( .A(n_1112), .B(n_1117), .Y(n_1116) );
AND2x2_ASAP7_75t_L g1128 ( .A(n_1112), .B(n_1117), .Y(n_1128) );
AND2x4_ASAP7_75t_L g1135 ( .A(n_1112), .B(n_1117), .Y(n_1135) );
AND2x2_ASAP7_75t_L g1119 ( .A(n_1120), .B(n_1130), .Y(n_1119) );
INVx1_ASAP7_75t_L g1168 ( .A(n_1120), .Y(n_1168) );
AND2x2_ASAP7_75t_L g1208 ( .A(n_1120), .B(n_1159), .Y(n_1208) );
AND2x2_ASAP7_75t_L g1273 ( .A(n_1120), .B(n_1156), .Y(n_1273) );
AND2x2_ASAP7_75t_L g1291 ( .A(n_1120), .B(n_1144), .Y(n_1291) );
AND2x2_ASAP7_75t_L g1120 ( .A(n_1121), .B(n_1125), .Y(n_1120) );
CKINVDCx5p33_ASAP7_75t_R g1161 ( .A(n_1121), .Y(n_1161) );
OR2x2_ASAP7_75t_L g1169 ( .A(n_1121), .B(n_1125), .Y(n_1169) );
AND2x2_ASAP7_75t_L g1121 ( .A(n_1122), .B(n_1123), .Y(n_1121) );
INVx2_ASAP7_75t_L g1137 ( .A(n_1124), .Y(n_1137) );
OR2x2_ASAP7_75t_L g1160 ( .A(n_1125), .B(n_1161), .Y(n_1160) );
AND2x2_ASAP7_75t_L g1181 ( .A(n_1125), .B(n_1161), .Y(n_1181) );
NAND2xp5_ASAP7_75t_L g1201 ( .A(n_1125), .B(n_1156), .Y(n_1201) );
AND2x2_ASAP7_75t_L g1214 ( .A(n_1125), .B(n_1215), .Y(n_1214) );
OR2x2_ASAP7_75t_L g1320 ( .A(n_1125), .B(n_1145), .Y(n_1320) );
AND2x2_ASAP7_75t_L g1125 ( .A(n_1126), .B(n_1129), .Y(n_1125) );
INVx3_ASAP7_75t_L g1140 ( .A(n_1127), .Y(n_1140) );
AND2x2_ASAP7_75t_L g1188 ( .A(n_1130), .B(n_1181), .Y(n_1188) );
INVx1_ASAP7_75t_L g1130 ( .A(n_1131), .Y(n_1130) );
NOR2xp33_ASAP7_75t_L g1295 ( .A(n_1131), .B(n_1160), .Y(n_1295) );
NAND2xp5_ASAP7_75t_L g1131 ( .A(n_1132), .B(n_1144), .Y(n_1131) );
INVx2_ASAP7_75t_L g1159 ( .A(n_1132), .Y(n_1159) );
INVx3_ASAP7_75t_L g1193 ( .A(n_1132), .Y(n_1193) );
NAND2xp5_ASAP7_75t_L g1264 ( .A(n_1132), .B(n_1198), .Y(n_1264) );
NOR2xp33_ASAP7_75t_L g1269 ( .A(n_1132), .B(n_1160), .Y(n_1269) );
NAND2xp5_ASAP7_75t_L g1284 ( .A(n_1132), .B(n_1285), .Y(n_1284) );
HB1xp67_ASAP7_75t_L g1289 ( .A(n_1132), .Y(n_1289) );
NOR2xp33_ASAP7_75t_L g1334 ( .A(n_1132), .B(n_1151), .Y(n_1334) );
OR2x2_ASAP7_75t_L g1132 ( .A(n_1133), .B(n_1139), .Y(n_1132) );
OAI22xp5_ASAP7_75t_L g1133 ( .A1(n_1134), .A2(n_1136), .B1(n_1137), .B2(n_1138), .Y(n_1133) );
OAI22xp5_ASAP7_75t_L g1220 ( .A1(n_1134), .A2(n_1137), .B1(n_1221), .B2(n_1222), .Y(n_1220) );
INVx3_ASAP7_75t_L g1134 ( .A(n_1135), .Y(n_1134) );
OAI22xp5_ASAP7_75t_L g1139 ( .A1(n_1140), .A2(n_1141), .B1(n_1142), .B2(n_1143), .Y(n_1139) );
INVx1_ASAP7_75t_L g1219 ( .A(n_1140), .Y(n_1219) );
XNOR2x1_ASAP7_75t_L g1346 ( .A(n_1141), .B(n_1347), .Y(n_1346) );
OAI311xp33_ASAP7_75t_L g1165 ( .A1(n_1144), .A2(n_1166), .A3(n_1170), .B1(n_1179), .C1(n_1185), .Y(n_1165) );
A2O1A1Ixp33_ASAP7_75t_L g1179 ( .A1(n_1144), .A2(n_1180), .B(n_1181), .C(n_1182), .Y(n_1179) );
NAND2xp5_ASAP7_75t_L g1195 ( .A(n_1144), .B(n_1161), .Y(n_1195) );
HB1xp67_ASAP7_75t_L g1215 ( .A(n_1144), .Y(n_1215) );
OR2x2_ASAP7_75t_L g1228 ( .A(n_1144), .B(n_1169), .Y(n_1228) );
AND2x2_ASAP7_75t_L g1236 ( .A(n_1144), .B(n_1237), .Y(n_1236) );
NAND2xp5_ASAP7_75t_L g1242 ( .A(n_1144), .B(n_1243), .Y(n_1242) );
OR2x2_ASAP7_75t_L g1282 ( .A(n_1144), .B(n_1161), .Y(n_1282) );
NAND2xp5_ASAP7_75t_L g1298 ( .A(n_1144), .B(n_1212), .Y(n_1298) );
NOR2xp33_ASAP7_75t_L g1307 ( .A(n_1144), .B(n_1160), .Y(n_1307) );
NAND2xp5_ASAP7_75t_L g1322 ( .A(n_1144), .B(n_1269), .Y(n_1322) );
INVx3_ASAP7_75t_L g1144 ( .A(n_1145), .Y(n_1144) );
INVx1_ASAP7_75t_L g1157 ( .A(n_1145), .Y(n_1157) );
NAND2xp5_ASAP7_75t_L g1255 ( .A(n_1145), .B(n_1193), .Y(n_1255) );
AND2x2_ASAP7_75t_L g1145 ( .A(n_1146), .B(n_1148), .Y(n_1145) );
NAND2xp5_ASAP7_75t_L g1183 ( .A(n_1149), .B(n_1184), .Y(n_1183) );
AND2x2_ASAP7_75t_L g1240 ( .A(n_1149), .B(n_1172), .Y(n_1240) );
INVx2_ASAP7_75t_L g1149 ( .A(n_1150), .Y(n_1149) );
INVx1_ASAP7_75t_L g1150 ( .A(n_1151), .Y(n_1150) );
CKINVDCx6p67_ASAP7_75t_R g1164 ( .A(n_1151), .Y(n_1164) );
AND2x2_ASAP7_75t_L g1198 ( .A(n_1151), .B(n_1199), .Y(n_1198) );
OR2x2_ASAP7_75t_L g1239 ( .A(n_1151), .B(n_1172), .Y(n_1239) );
OR2x6_ASAP7_75t_L g1151 ( .A(n_1152), .B(n_1153), .Y(n_1151) );
INVx1_ASAP7_75t_L g1154 ( .A(n_1155), .Y(n_1154) );
NAND2xp5_ASAP7_75t_L g1155 ( .A(n_1156), .B(n_1158), .Y(n_1155) );
AND2x2_ASAP7_75t_L g1246 ( .A(n_1156), .B(n_1181), .Y(n_1246) );
AND2x2_ASAP7_75t_L g1262 ( .A(n_1156), .B(n_1161), .Y(n_1262) );
AOI211xp5_ASAP7_75t_L g1318 ( .A1(n_1156), .A2(n_1159), .B(n_1160), .C(n_1319), .Y(n_1318) );
AND3x1_ASAP7_75t_L g1335 ( .A(n_1156), .B(n_1210), .C(n_1212), .Y(n_1335) );
INVx3_ASAP7_75t_L g1156 ( .A(n_1157), .Y(n_1156) );
NOR2xp33_ASAP7_75t_L g1158 ( .A(n_1159), .B(n_1160), .Y(n_1158) );
NAND2xp5_ASAP7_75t_L g1170 ( .A(n_1159), .B(n_1171), .Y(n_1170) );
INVx1_ASAP7_75t_L g1226 ( .A(n_1159), .Y(n_1226) );
NAND2xp5_ASAP7_75t_L g1290 ( .A(n_1159), .B(n_1291), .Y(n_1290) );
NAND2xp5_ASAP7_75t_L g1331 ( .A(n_1159), .B(n_1273), .Y(n_1331) );
INVx1_ASAP7_75t_L g1243 ( .A(n_1160), .Y(n_1243) );
AOI21xp33_ASAP7_75t_L g1304 ( .A1(n_1162), .A2(n_1305), .B(n_1306), .Y(n_1304) );
CKINVDCx14_ASAP7_75t_R g1162 ( .A(n_1163), .Y(n_1162) );
INVx1_ASAP7_75t_L g1163 ( .A(n_1164), .Y(n_1163) );
NAND3xp33_ASAP7_75t_L g1213 ( .A(n_1164), .B(n_1214), .C(n_1216), .Y(n_1213) );
NAND2xp5_ASAP7_75t_L g1276 ( .A(n_1164), .B(n_1172), .Y(n_1276) );
AND2x2_ASAP7_75t_L g1296 ( .A(n_1164), .B(n_1231), .Y(n_1296) );
INVx1_ASAP7_75t_L g1166 ( .A(n_1167), .Y(n_1166) );
NAND2xp5_ASAP7_75t_L g1167 ( .A(n_1168), .B(n_1169), .Y(n_1167) );
INVx1_ASAP7_75t_L g1237 ( .A(n_1169), .Y(n_1237) );
NOR2xp33_ASAP7_75t_L g1278 ( .A(n_1169), .B(n_1193), .Y(n_1278) );
NOR2xp33_ASAP7_75t_L g1337 ( .A(n_1169), .B(n_1289), .Y(n_1337) );
INVx3_ASAP7_75t_L g1180 ( .A(n_1171), .Y(n_1180) );
NAND2xp5_ASAP7_75t_L g1197 ( .A(n_1171), .B(n_1198), .Y(n_1197) );
NAND2xp5_ASAP7_75t_L g1206 ( .A(n_1171), .B(n_1207), .Y(n_1206) );
INVx5_ASAP7_75t_L g1260 ( .A(n_1171), .Y(n_1260) );
AOI22xp5_ASAP7_75t_L g1323 ( .A1(n_1171), .A2(n_1312), .B1(n_1324), .B2(n_1327), .Y(n_1323) );
NAND2xp5_ASAP7_75t_L g1328 ( .A(n_1171), .B(n_1285), .Y(n_1328) );
INVx3_ASAP7_75t_L g1171 ( .A(n_1172), .Y(n_1171) );
AND2x2_ASAP7_75t_L g1209 ( .A(n_1172), .B(n_1210), .Y(n_1209) );
AND2x2_ASAP7_75t_L g1230 ( .A(n_1172), .B(n_1231), .Y(n_1230) );
INVx3_ASAP7_75t_L g1172 ( .A(n_1173), .Y(n_1172) );
OR2x2_ASAP7_75t_L g1300 ( .A(n_1173), .B(n_1301), .Y(n_1300) );
OR2x2_ASAP7_75t_L g1317 ( .A(n_1173), .B(n_1187), .Y(n_1317) );
NAND2xp5_ASAP7_75t_L g1173 ( .A(n_1174), .B(n_1178), .Y(n_1173) );
INVx2_ASAP7_75t_L g1175 ( .A(n_1176), .Y(n_1175) );
INVx2_ASAP7_75t_SL g1176 ( .A(n_1177), .Y(n_1176) );
NAND2xp5_ASAP7_75t_L g1203 ( .A(n_1180), .B(n_1198), .Y(n_1203) );
AND2x2_ASAP7_75t_L g1212 ( .A(n_1181), .B(n_1193), .Y(n_1212) );
AND2x2_ASAP7_75t_L g1270 ( .A(n_1181), .B(n_1192), .Y(n_1270) );
INVx1_ASAP7_75t_L g1293 ( .A(n_1181), .Y(n_1293) );
AND2x2_ASAP7_75t_L g1341 ( .A(n_1181), .B(n_1215), .Y(n_1341) );
INVx1_ASAP7_75t_L g1182 ( .A(n_1183), .Y(n_1182) );
OAI21xp33_ASAP7_75t_L g1324 ( .A1(n_1183), .A2(n_1282), .B(n_1325), .Y(n_1324) );
NAND2xp5_ASAP7_75t_L g1185 ( .A(n_1186), .B(n_1188), .Y(n_1185) );
AOI222xp33_ASAP7_75t_L g1265 ( .A1(n_1186), .A2(n_1205), .B1(n_1237), .B2(n_1266), .C1(n_1267), .C2(n_1270), .Y(n_1265) );
INVx2_ASAP7_75t_L g1186 ( .A(n_1187), .Y(n_1186) );
INVx1_ASAP7_75t_L g1224 ( .A(n_1188), .Y(n_1224) );
AOI22xp33_ASAP7_75t_L g1189 ( .A1(n_1190), .A2(n_1196), .B1(n_1200), .B2(n_1202), .Y(n_1189) );
INVxp33_ASAP7_75t_SL g1190 ( .A(n_1191), .Y(n_1190) );
NAND2xp5_ASAP7_75t_L g1191 ( .A(n_1192), .B(n_1194), .Y(n_1191) );
INVx1_ASAP7_75t_SL g1192 ( .A(n_1193), .Y(n_1192) );
AND2x2_ASAP7_75t_L g1312 ( .A(n_1193), .B(n_1236), .Y(n_1312) );
INVx1_ASAP7_75t_L g1194 ( .A(n_1195), .Y(n_1194) );
INVx1_ASAP7_75t_L g1196 ( .A(n_1197), .Y(n_1196) );
OAI32xp33_ASAP7_75t_L g1338 ( .A1(n_1197), .A2(n_1217), .A3(n_1239), .B1(n_1339), .B2(n_1340), .Y(n_1338) );
INVx1_ASAP7_75t_L g1211 ( .A(n_1199), .Y(n_1211) );
INVx1_ASAP7_75t_L g1200 ( .A(n_1201), .Y(n_1200) );
AOI222xp33_ASAP7_75t_L g1314 ( .A1(n_1202), .A2(n_1296), .B1(n_1315), .B2(n_1316), .C1(n_1318), .C2(n_1321), .Y(n_1314) );
INVx1_ASAP7_75t_L g1202 ( .A(n_1203), .Y(n_1202) );
AOI22xp5_ASAP7_75t_L g1204 ( .A1(n_1205), .A2(n_1208), .B1(n_1209), .B2(n_1212), .Y(n_1204) );
INVx1_ASAP7_75t_L g1205 ( .A(n_1206), .Y(n_1205) );
NOR2xp33_ASAP7_75t_L g1302 ( .A(n_1207), .B(n_1253), .Y(n_1302) );
NAND2xp5_ASAP7_75t_L g1245 ( .A(n_1209), .B(n_1246), .Y(n_1245) );
INVx1_ASAP7_75t_L g1210 ( .A(n_1211), .Y(n_1210) );
A2O1A1Ixp33_ASAP7_75t_L g1303 ( .A1(n_1214), .A2(n_1263), .B(n_1304), .C(n_1308), .Y(n_1303) );
INVx1_ASAP7_75t_L g1339 ( .A(n_1214), .Y(n_1339) );
INVx1_ASAP7_75t_L g1216 ( .A(n_1217), .Y(n_1216) );
INVx2_ASAP7_75t_L g1279 ( .A(n_1218), .Y(n_1279) );
HB1xp67_ASAP7_75t_L g1343 ( .A(n_1219), .Y(n_1343) );
A2O1A1Ixp33_ASAP7_75t_L g1223 ( .A1(n_1224), .A2(n_1225), .B(n_1229), .C(n_1232), .Y(n_1223) );
AOI21xp33_ASAP7_75t_L g1332 ( .A1(n_1224), .A2(n_1276), .B(n_1305), .Y(n_1332) );
NAND2xp5_ASAP7_75t_L g1225 ( .A(n_1226), .B(n_1227), .Y(n_1225) );
O2A1O1Ixp33_ASAP7_75t_L g1336 ( .A1(n_1227), .A2(n_1266), .B(n_1337), .C(n_1338), .Y(n_1336) );
INVx1_ASAP7_75t_L g1227 ( .A(n_1228), .Y(n_1227) );
INVx1_ASAP7_75t_L g1229 ( .A(n_1230), .Y(n_1229) );
AOI221xp5_ASAP7_75t_SL g1232 ( .A1(n_1233), .A2(n_1238), .B1(n_1240), .B2(n_1241), .C(n_1244), .Y(n_1232) );
NOR2xp33_ASAP7_75t_L g1233 ( .A(n_1234), .B(n_1235), .Y(n_1233) );
INVx1_ASAP7_75t_L g1259 ( .A(n_1234), .Y(n_1259) );
NAND2xp5_ASAP7_75t_L g1281 ( .A(n_1235), .B(n_1282), .Y(n_1281) );
INVx1_ASAP7_75t_L g1235 ( .A(n_1236), .Y(n_1235) );
NAND3xp33_ASAP7_75t_L g1258 ( .A(n_1236), .B(n_1259), .C(n_1260), .Y(n_1258) );
AOI221xp5_ASAP7_75t_L g1280 ( .A1(n_1238), .A2(n_1281), .B1(n_1283), .B2(n_1286), .C(n_1292), .Y(n_1280) );
INVx1_ASAP7_75t_L g1238 ( .A(n_1239), .Y(n_1238) );
INVx1_ASAP7_75t_L g1249 ( .A(n_1240), .Y(n_1249) );
NOR2xp33_ASAP7_75t_L g1287 ( .A(n_1241), .B(n_1262), .Y(n_1287) );
INVx1_ASAP7_75t_L g1241 ( .A(n_1242), .Y(n_1241) );
NAND2xp5_ASAP7_75t_L g1253 ( .A(n_1243), .B(n_1254), .Y(n_1253) );
INVxp67_ASAP7_75t_SL g1244 ( .A(n_1245), .Y(n_1244) );
INVx1_ASAP7_75t_L g1256 ( .A(n_1246), .Y(n_1256) );
NAND5xp2_ASAP7_75t_L g1247 ( .A(n_1248), .B(n_1280), .C(n_1294), .D(n_1303), .E(n_1309), .Y(n_1247) );
AOI211xp5_ASAP7_75t_L g1248 ( .A1(n_1249), .A2(n_1250), .B(n_1257), .C(n_1271), .Y(n_1248) );
OAI221xp5_ASAP7_75t_L g1271 ( .A1(n_1249), .A2(n_1272), .B1(n_1274), .B2(n_1277), .C(n_1279), .Y(n_1271) );
INVxp67_ASAP7_75t_L g1250 ( .A(n_1251), .Y(n_1250) );
NAND2xp5_ASAP7_75t_L g1252 ( .A(n_1253), .B(n_1256), .Y(n_1252) );
INVx1_ASAP7_75t_L g1254 ( .A(n_1255), .Y(n_1254) );
NAND3xp33_ASAP7_75t_L g1257 ( .A(n_1258), .B(n_1261), .C(n_1265), .Y(n_1257) );
NOR2xp33_ASAP7_75t_L g1274 ( .A(n_1259), .B(n_1275), .Y(n_1274) );
CKINVDCx14_ASAP7_75t_R g1308 ( .A(n_1260), .Y(n_1308) );
NOR2xp33_ASAP7_75t_L g1310 ( .A(n_1260), .B(n_1311), .Y(n_1310) );
A2O1A1Ixp33_ASAP7_75t_L g1333 ( .A1(n_1260), .A2(n_1262), .B(n_1334), .C(n_1335), .Y(n_1333) );
NAND2xp5_ASAP7_75t_L g1261 ( .A(n_1262), .B(n_1263), .Y(n_1261) );
INVx1_ASAP7_75t_L g1263 ( .A(n_1264), .Y(n_1263) );
NOR2xp33_ASAP7_75t_L g1292 ( .A(n_1264), .B(n_1293), .Y(n_1292) );
INVx2_ASAP7_75t_L g1267 ( .A(n_1268), .Y(n_1267) );
INVx1_ASAP7_75t_L g1268 ( .A(n_1269), .Y(n_1268) );
INVx1_ASAP7_75t_L g1272 ( .A(n_1273), .Y(n_1272) );
INVx1_ASAP7_75t_L g1275 ( .A(n_1276), .Y(n_1275) );
INVxp67_ASAP7_75t_L g1277 ( .A(n_1278), .Y(n_1277) );
O2A1O1Ixp33_ASAP7_75t_L g1329 ( .A1(n_1278), .A2(n_1299), .B(n_1330), .C(n_1332), .Y(n_1329) );
INVx1_ASAP7_75t_L g1283 ( .A(n_1284), .Y(n_1283) );
INVx2_ASAP7_75t_L g1301 ( .A(n_1285), .Y(n_1301) );
OAI21xp33_ASAP7_75t_L g1286 ( .A1(n_1287), .A2(n_1288), .B(n_1290), .Y(n_1286) );
INVx1_ASAP7_75t_L g1288 ( .A(n_1289), .Y(n_1288) );
INVx1_ASAP7_75t_L g1315 ( .A(n_1290), .Y(n_1315) );
AOI221xp5_ASAP7_75t_L g1294 ( .A1(n_1295), .A2(n_1296), .B1(n_1297), .B2(n_1299), .C(n_1302), .Y(n_1294) );
INVx1_ASAP7_75t_L g1297 ( .A(n_1298), .Y(n_1297) );
INVx1_ASAP7_75t_L g1299 ( .A(n_1300), .Y(n_1299) );
INVx1_ASAP7_75t_L g1326 ( .A(n_1301), .Y(n_1326) );
INVx1_ASAP7_75t_L g1306 ( .A(n_1307), .Y(n_1306) );
NAND2xp5_ASAP7_75t_L g1325 ( .A(n_1307), .B(n_1326), .Y(n_1325) );
INVxp67_ASAP7_75t_L g1309 ( .A(n_1310), .Y(n_1309) );
INVx1_ASAP7_75t_L g1311 ( .A(n_1312), .Y(n_1311) );
NAND5xp2_ASAP7_75t_SL g1313 ( .A(n_1314), .B(n_1323), .C(n_1329), .D(n_1333), .E(n_1336), .Y(n_1313) );
INVx1_ASAP7_75t_L g1316 ( .A(n_1317), .Y(n_1316) );
INVx1_ASAP7_75t_L g1319 ( .A(n_1320), .Y(n_1319) );
INVx1_ASAP7_75t_L g1321 ( .A(n_1322), .Y(n_1321) );
INVx1_ASAP7_75t_L g1327 ( .A(n_1328), .Y(n_1327) );
INVxp67_ASAP7_75t_SL g1330 ( .A(n_1331), .Y(n_1330) );
INVx1_ASAP7_75t_L g1340 ( .A(n_1341), .Y(n_1340) );
CKINVDCx5p33_ASAP7_75t_R g1342 ( .A(n_1343), .Y(n_1342) );
INVx1_ASAP7_75t_L g1344 ( .A(n_1345), .Y(n_1344) );
INVx4_ASAP7_75t_R g1345 ( .A(n_1346), .Y(n_1345) );
AND2x4_ASAP7_75t_L g1347 ( .A(n_1348), .B(n_1362), .Y(n_1347) );
NOR3xp33_ASAP7_75t_L g1348 ( .A(n_1349), .B(n_1354), .C(n_1357), .Y(n_1348) );
OAI21xp5_ASAP7_75t_L g1349 ( .A1(n_1350), .A2(n_1351), .B(n_1352), .Y(n_1349) );
INVxp67_ASAP7_75t_L g1360 ( .A(n_1361), .Y(n_1360) );
AND4x1_ASAP7_75t_L g1362 ( .A(n_1363), .B(n_1364), .C(n_1365), .D(n_1366), .Y(n_1362) );
CKINVDCx16_ASAP7_75t_R g1367 ( .A(n_1368), .Y(n_1367) );
INVxp33_ASAP7_75t_SL g1372 ( .A(n_1373), .Y(n_1372) );
INVxp67_ASAP7_75t_SL g1397 ( .A(n_1374), .Y(n_1397) );
AND2x2_ASAP7_75t_L g1374 ( .A(n_1375), .B(n_1389), .Y(n_1374) );
NOR3xp33_ASAP7_75t_L g1375 ( .A(n_1376), .B(n_1380), .C(n_1385), .Y(n_1375) );
INVx1_ASAP7_75t_L g1383 ( .A(n_1384), .Y(n_1383) );
OAI21xp33_ASAP7_75t_L g1385 ( .A1(n_1386), .A2(n_1387), .B(n_1388), .Y(n_1385) );
NOR2xp33_ASAP7_75t_L g1389 ( .A(n_1390), .B(n_1393), .Y(n_1389) );
NAND2xp5_ASAP7_75t_L g1390 ( .A(n_1391), .B(n_1392), .Y(n_1390) );
NAND2xp5_ASAP7_75t_L g1393 ( .A(n_1394), .B(n_1395), .Y(n_1393) );
BUFx2_ASAP7_75t_SL g1398 ( .A(n_1399), .Y(n_1398) );
HB1xp67_ASAP7_75t_L g1400 ( .A(n_1401), .Y(n_1400) );
endmodule