module fake_netlist_5_1268_n_1236 (n_137, n_168, n_164, n_91, n_82, n_122, n_142, n_176, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_165, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_177, n_60, n_155, n_152, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_125, n_35, n_167, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_157, n_29, n_79, n_131, n_151, n_47, n_173, n_25, n_53, n_160, n_8, n_158, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_159, n_163, n_95, n_119, n_175, n_169, n_59, n_26, n_133, n_55, n_99, n_2, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_178, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_162, n_27, n_170, n_64, n_77, n_102, n_106, n_161, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_174, n_134, n_32, n_41, n_104, n_172, n_103, n_56, n_51, n_63, n_97, n_141, n_166, n_11, n_171, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_1236);

input n_137;
input n_168;
input n_164;
input n_91;
input n_82;
input n_122;
input n_142;
input n_176;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_165;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_177;
input n_60;
input n_155;
input n_152;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_125;
input n_35;
input n_167;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_157;
input n_29;
input n_79;
input n_131;
input n_151;
input n_47;
input n_173;
input n_25;
input n_53;
input n_160;
input n_8;
input n_158;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_159;
input n_163;
input n_95;
input n_119;
input n_175;
input n_169;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_178;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_162;
input n_27;
input n_170;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_174;
input n_134;
input n_32;
input n_41;
input n_104;
input n_172;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_166;
input n_11;
input n_171;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_1236;

wire n_924;
wire n_977;
wire n_611;
wire n_1126;
wire n_1166;
wire n_469;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1150;
wire n_226;
wire n_667;
wire n_790;
wire n_1055;
wire n_880;
wire n_544;
wire n_1007;
wire n_552;
wire n_1198;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1021;
wire n_551;
wire n_688;
wire n_800;
wire n_671;
wire n_819;
wire n_1022;
wire n_915;
wire n_864;
wire n_859;
wire n_951;
wire n_447;
wire n_247;
wire n_292;
wire n_625;
wire n_854;
wire n_674;
wire n_417;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_606;
wire n_275;
wire n_877;
wire n_755;
wire n_1118;
wire n_947;
wire n_373;
wire n_307;
wire n_530;
wire n_1107;
wire n_556;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_929;
wire n_1124;
wire n_902;
wire n_191;
wire n_1104;
wire n_659;
wire n_1182;
wire n_579;
wire n_938;
wire n_1098;
wire n_320;
wire n_1154;
wire n_1135;
wire n_406;
wire n_519;
wire n_1016;
wire n_546;
wire n_281;
wire n_240;
wire n_291;
wire n_231;
wire n_257;
wire n_731;
wire n_371;
wire n_709;
wire n_317;
wire n_569;
wire n_227;
wire n_920;
wire n_335;
wire n_370;
wire n_976;
wire n_343;
wire n_308;
wire n_297;
wire n_1078;
wire n_775;
wire n_219;
wire n_600;
wire n_223;
wire n_264;
wire n_955;
wire n_339;
wire n_1146;
wire n_882;
wire n_183;
wire n_243;
wire n_1036;
wire n_1097;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_215;
wire n_350;
wire n_196;
wire n_798;
wire n_646;
wire n_436;
wire n_1216;
wire n_290;
wire n_580;
wire n_1040;
wire n_578;
wire n_926;
wire n_344;
wire n_1218;
wire n_422;
wire n_475;
wire n_777;
wire n_1070;
wire n_1030;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_496;
wire n_958;
wire n_1034;
wire n_670;
wire n_521;
wire n_663;
wire n_845;
wire n_673;
wire n_837;
wire n_528;
wire n_680;
wire n_395;
wire n_553;
wire n_901;
wire n_813;
wire n_214;
wire n_675;
wire n_888;
wire n_1167;
wire n_637;
wire n_184;
wire n_446;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_468;
wire n_213;
wire n_342;
wire n_464;
wire n_363;
wire n_197;
wire n_1069;
wire n_1075;
wire n_460;
wire n_889;
wire n_973;
wire n_477;
wire n_571;
wire n_461;
wire n_1211;
wire n_1197;
wire n_907;
wire n_190;
wire n_989;
wire n_1039;
wire n_228;
wire n_283;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1002;
wire n_310;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_230;
wire n_953;
wire n_279;
wire n_1014;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_440;
wire n_793;
wire n_478;
wire n_476;
wire n_534;
wire n_884;
wire n_345;
wire n_944;
wire n_182;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_832;
wire n_857;
wire n_207;
wire n_561;
wire n_1027;
wire n_971;
wire n_1156;
wire n_794;
wire n_326;
wire n_404;
wire n_686;
wire n_847;
wire n_596;
wire n_558;
wire n_702;
wire n_822;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1199;
wire n_352;
wire n_1038;
wire n_520;
wire n_409;
wire n_887;
wire n_300;
wire n_809;
wire n_870;
wire n_931;
wire n_599;
wire n_434;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_965;
wire n_935;
wire n_1175;
wire n_817;
wire n_360;
wire n_759;
wire n_806;
wire n_324;
wire n_187;
wire n_1189;
wire n_706;
wire n_746;
wire n_747;
wire n_784;
wire n_431;
wire n_1194;
wire n_615;
wire n_851;
wire n_843;
wire n_523;
wire n_913;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_776;
wire n_367;
wire n_452;
wire n_525;
wire n_649;
wire n_547;
wire n_1191;
wire n_284;
wire n_1128;
wire n_744;
wire n_590;
wire n_629;
wire n_254;
wire n_1233;
wire n_526;
wire n_372;
wire n_293;
wire n_677;
wire n_244;
wire n_1121;
wire n_314;
wire n_368;
wire n_433;
wire n_604;
wire n_949;
wire n_1008;
wire n_946;
wire n_1001;
wire n_498;
wire n_689;
wire n_738;
wire n_640;
wire n_252;
wire n_624;
wire n_295;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1195;
wire n_610;
wire n_936;
wire n_568;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_259;
wire n_448;
wire n_758;
wire n_999;
wire n_1158;
wire n_563;
wire n_1145;
wire n_878;
wire n_524;
wire n_204;
wire n_394;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1068;
wire n_331;
wire n_906;
wire n_1163;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_658;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_592;
wire n_1169;
wire n_1017;
wire n_978;
wire n_1054;
wire n_1095;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_484;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1009;
wire n_1148;
wire n_742;
wire n_750;
wire n_995;
wire n_454;
wire n_374;
wire n_185;
wire n_396;
wire n_1073;
wire n_255;
wire n_662;
wire n_459;
wire n_218;
wire n_962;
wire n_1215;
wire n_1171;
wire n_723;
wire n_1065;
wire n_473;
wire n_1043;
wire n_355;
wire n_486;
wire n_614;
wire n_337;
wire n_1177;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_208;
wire n_743;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_829;
wire n_361;
wire n_700;
wire n_573;
wire n_1132;
wire n_388;
wire n_1127;
wire n_761;
wire n_1006;
wire n_329;
wire n_274;
wire n_582;
wire n_309;
wire n_512;
wire n_322;
wire n_652;
wire n_1111;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_224;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_239;
wire n_630;
wire n_504;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_987;
wire n_261;
wire n_767;
wire n_993;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_729;
wire n_1131;
wire n_1084;
wire n_970;
wire n_911;
wire n_513;
wire n_1094;
wire n_560;
wire n_340;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_495;
wire n_602;
wire n_574;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_490;
wire n_996;
wire n_921;
wire n_233;
wire n_572;
wire n_366;
wire n_815;
wire n_327;
wire n_1037;
wire n_1080;
wire n_426;
wire n_1082;
wire n_589;
wire n_716;
wire n_562;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_531;
wire n_890;
wire n_764;
wire n_1056;
wire n_960;
wire n_222;
wire n_1123;
wire n_1047;
wire n_634;
wire n_199;
wire n_348;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_256;
wire n_950;
wire n_380;
wire n_419;
wire n_444;
wire n_1060;
wire n_1141;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_912;
wire n_968;
wire n_315;
wire n_451;
wire n_619;
wire n_408;
wire n_376;
wire n_967;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_483;
wire n_683;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_983;
wire n_280;
wire n_873;
wire n_378;
wire n_1112;
wire n_762;
wire n_690;
wire n_583;
wire n_302;
wire n_1203;
wire n_821;
wire n_321;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_212;
wire n_385;
wire n_507;
wire n_330;
wire n_1228;
wire n_972;
wire n_692;
wire n_820;
wire n_1200;
wire n_1185;
wire n_991;
wire n_828;
wire n_779;
wire n_576;
wire n_1143;
wire n_804;
wire n_537;
wire n_945;
wire n_492;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_286;
wire n_883;
wire n_470;
wire n_449;
wire n_325;
wire n_1214;
wire n_900;
wire n_856;
wire n_918;
wire n_942;
wire n_189;
wire n_1147;
wire n_1077;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_195;
wire n_356;
wire n_894;
wire n_831;
wire n_964;
wire n_1096;
wire n_234;
wire n_833;
wire n_225;
wire n_988;
wire n_814;
wire n_192;
wire n_1201;
wire n_1114;
wire n_655;
wire n_669;
wire n_472;
wire n_1176;
wire n_387;
wire n_1149;
wire n_398;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_211;
wire n_1219;
wire n_1204;
wire n_1035;
wire n_287;
wire n_555;
wire n_783;
wire n_1188;
wire n_661;
wire n_849;
wire n_336;
wire n_584;
wire n_681;
wire n_430;
wire n_510;
wire n_216;
wire n_311;
wire n_830;
wire n_801;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_445;
wire n_749;
wire n_1134;
wire n_717;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1019;
wire n_1105;
wire n_249;
wire n_304;
wire n_577;
wire n_338;
wire n_693;
wire n_836;
wire n_990;
wire n_975;
wire n_567;
wire n_778;
wire n_1122;
wire n_306;
wire n_458;
wire n_770;
wire n_1102;
wire n_711;
wire n_1187;
wire n_1164;
wire n_489;
wire n_1174;
wire n_617;
wire n_876;
wire n_1190;
wire n_601;
wire n_917;
wire n_966;
wire n_253;
wire n_1116;
wire n_1212;
wire n_206;
wire n_217;
wire n_726;
wire n_982;
wire n_818;
wire n_861;
wire n_1183;
wire n_899;
wire n_210;
wire n_774;
wire n_1059;
wire n_1133;
wire n_557;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_1168;
wire n_707;
wire n_937;
wire n_393;
wire n_487;
wire n_665;
wire n_421;
wire n_910;
wire n_768;
wire n_205;
wire n_1136;
wire n_754;
wire n_179;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_735;
wire n_232;
wire n_1109;
wire n_895;
wire n_202;
wire n_427;
wire n_791;
wire n_732;
wire n_193;
wire n_808;
wire n_797;
wire n_1025;
wire n_500;
wire n_1067;
wire n_435;
wire n_766;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1213;
wire n_536;
wire n_872;
wire n_594;
wire n_200;
wire n_1155;
wire n_1011;
wire n_1184;
wire n_985;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_626;
wire n_1144;
wire n_1137;
wire n_1170;
wire n_305;
wire n_676;
wire n_294;
wire n_318;
wire n_653;
wire n_642;
wire n_194;
wire n_855;
wire n_1178;
wire n_850;
wire n_684;
wire n_268;
wire n_664;
wire n_503;
wire n_235;
wire n_605;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_1115;
wire n_980;
wire n_780;
wire n_998;
wire n_467;
wire n_1227;
wire n_840;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_672;
wire n_581;
wire n_382;
wire n_554;
wire n_898;
wire n_1013;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_198;
wire n_714;
wire n_909;
wire n_997;
wire n_932;
wire n_612;
wire n_788;
wire n_559;
wire n_825;
wire n_508;
wire n_506;
wire n_737;
wire n_986;
wire n_509;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_209;
wire n_733;
wire n_941;
wire n_981;
wire n_867;
wire n_186;
wire n_587;
wire n_792;
wire n_756;
wire n_399;
wire n_548;
wire n_812;
wire n_298;
wire n_518;
wire n_505;
wire n_282;
wire n_752;
wire n_905;
wire n_1108;
wire n_782;
wire n_1100;
wire n_862;
wire n_760;
wire n_381;
wire n_220;
wire n_390;
wire n_481;
wire n_769;
wire n_1046;
wire n_271;
wire n_934;
wire n_826;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_379;
wire n_428;
wire n_570;
wire n_853;
wire n_377;
wire n_751;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_704;
wire n_787;
wire n_961;
wire n_771;
wire n_276;
wire n_1225;
wire n_522;
wire n_400;
wire n_930;
wire n_181;
wire n_221;
wire n_622;
wire n_1087;
wire n_386;
wire n_994;
wire n_848;
wire n_1223;
wire n_682;
wire n_922;
wire n_816;
wire n_591;
wire n_313;
wire n_631;
wire n_479;
wire n_432;
wire n_839;
wire n_1210;
wire n_328;
wire n_369;
wire n_871;
wire n_598;
wire n_685;
wire n_608;
wire n_928;
wire n_772;
wire n_499;
wire n_517;
wire n_402;
wire n_413;
wire n_1086;
wire n_796;
wire n_236;
wire n_1012;
wire n_903;
wire n_740;
wire n_203;
wire n_384;
wire n_277;
wire n_1061;
wire n_333;
wire n_462;
wire n_1193;
wire n_258;
wire n_1113;
wire n_1226;
wire n_722;
wire n_188;
wire n_844;
wire n_201;
wire n_471;
wire n_852;
wire n_1028;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_632;
wire n_699;
wire n_979;
wire n_846;
wire n_465;
wire n_362;
wire n_273;
wire n_585;
wire n_270;
wire n_616;
wire n_745;
wire n_1103;
wire n_648;
wire n_312;
wire n_1076;
wire n_1091;
wire n_494;
wire n_641;
wire n_730;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_180;
wire n_656;
wire n_1220;
wire n_229;
wire n_437;
wire n_453;
wire n_403;
wire n_1130;
wire n_720;
wire n_863;
wire n_805;
wire n_712;
wire n_246;
wire n_1042;
wire n_269;
wire n_285;
wire n_412;
wire n_657;
wire n_644;
wire n_1160;
wire n_491;
wire n_1074;
wire n_251;
wire n_566;
wire n_565;
wire n_597;
wire n_1181;
wire n_1196;
wire n_651;
wire n_334;
wire n_811;
wire n_807;
wire n_835;
wire n_666;
wire n_262;
wire n_1026;
wire n_1234;
wire n_319;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_1004;
wire n_1186;
wire n_242;
wire n_1032;
wire n_1018;
wire n_438;
wire n_713;
wire n_904;
wire n_1180;
wire n_533;
wire n_278;

INVx1_ASAP7_75t_L g179 ( 
.A(n_88),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g180 ( 
.A(n_177),
.Y(n_180)
);

INVx2_ASAP7_75t_SL g181 ( 
.A(n_1),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_54),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_127),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_116),
.Y(n_184)
);

BUFx3_ASAP7_75t_L g185 ( 
.A(n_132),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_157),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_67),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_47),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_57),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_53),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_32),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_38),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_129),
.Y(n_193)
);

BUFx10_ASAP7_75t_L g194 ( 
.A(n_118),
.Y(n_194)
);

BUFx3_ASAP7_75t_L g195 ( 
.A(n_151),
.Y(n_195)
);

INVxp67_ASAP7_75t_L g196 ( 
.A(n_92),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_42),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_11),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_28),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_9),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_69),
.Y(n_201)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_142),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_9),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_65),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_115),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_123),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_159),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_101),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_58),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_23),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_61),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_56),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_106),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_62),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_24),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_17),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_6),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_149),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_11),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_96),
.Y(n_220)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_16),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_27),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_134),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_110),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_10),
.Y(n_225)
);

INVx1_ASAP7_75t_SL g226 ( 
.A(n_141),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_136),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_73),
.Y(n_228)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_166),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_87),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_19),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_144),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_85),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_160),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_147),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_16),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_186),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_188),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_189),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_190),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_197),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_201),
.Y(n_242)
);

HB1xp67_ASAP7_75t_L g243 ( 
.A(n_236),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_221),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_206),
.Y(n_245)
);

INVx1_ASAP7_75t_SL g246 ( 
.A(n_198),
.Y(n_246)
);

CKINVDCx16_ASAP7_75t_R g247 ( 
.A(n_194),
.Y(n_247)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_221),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_191),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_216),
.Y(n_250)
);

BUFx3_ASAP7_75t_L g251 ( 
.A(n_185),
.Y(n_251)
);

BUFx2_ASAP7_75t_SL g252 ( 
.A(n_184),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_209),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_231),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_211),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_212),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_181),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_214),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_218),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_220),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_223),
.Y(n_261)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_180),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_181),
.Y(n_263)
);

BUFx10_ASAP7_75t_L g264 ( 
.A(n_180),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_224),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_228),
.Y(n_266)
);

BUFx3_ASAP7_75t_L g267 ( 
.A(n_251),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_237),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_248),
.Y(n_269)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_262),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_238),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_239),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_248),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_240),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_262),
.Y(n_275)
);

INVx1_ASAP7_75t_SL g276 ( 
.A(n_246),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_241),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_242),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_245),
.Y(n_279)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_262),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_253),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_249),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_255),
.Y(n_283)
);

INVxp67_ASAP7_75t_SL g284 ( 
.A(n_251),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_256),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_258),
.Y(n_286)
);

INVx2_ASAP7_75t_SL g287 ( 
.A(n_251),
.Y(n_287)
);

INVx1_ASAP7_75t_SL g288 ( 
.A(n_252),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_249),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_250),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_257),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_250),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_259),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_254),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_260),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_254),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_244),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_261),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_265),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_266),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_252),
.Y(n_301)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_244),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_247),
.Y(n_303)
);

BUFx2_ASAP7_75t_L g304 ( 
.A(n_243),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_257),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_263),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_247),
.Y(n_307)
);

BUFx2_ASAP7_75t_L g308 ( 
.A(n_263),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_264),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_264),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_264),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_264),
.Y(n_312)
);

CKINVDCx16_ASAP7_75t_R g313 ( 
.A(n_247),
.Y(n_313)
);

INVxp67_ASAP7_75t_SL g314 ( 
.A(n_251),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_248),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_248),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_248),
.Y(n_317)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_262),
.Y(n_318)
);

INVxp67_ASAP7_75t_SL g319 ( 
.A(n_267),
.Y(n_319)
);

INVx2_ASAP7_75t_L g320 ( 
.A(n_270),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_313),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_270),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_280),
.Y(n_323)
);

INVx2_ASAP7_75t_L g324 ( 
.A(n_280),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_318),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_318),
.Y(n_326)
);

INVx2_ASAP7_75t_L g327 ( 
.A(n_275),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_268),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_282),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_282),
.Y(n_330)
);

INVx2_ASAP7_75t_L g331 ( 
.A(n_302),
.Y(n_331)
);

INVxp67_ASAP7_75t_L g332 ( 
.A(n_276),
.Y(n_332)
);

BUFx2_ASAP7_75t_L g333 ( 
.A(n_267),
.Y(n_333)
);

CKINVDCx14_ASAP7_75t_R g334 ( 
.A(n_303),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_284),
.B(n_226),
.Y(n_335)
);

INVxp33_ASAP7_75t_SL g336 ( 
.A(n_301),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_289),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_289),
.Y(n_338)
);

INVx3_ASAP7_75t_L g339 ( 
.A(n_302),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_290),
.Y(n_340)
);

INVx2_ASAP7_75t_L g341 ( 
.A(n_269),
.Y(n_341)
);

INVxp33_ASAP7_75t_L g342 ( 
.A(n_304),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_271),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_290),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_292),
.Y(n_345)
);

INVx1_ASAP7_75t_SL g346 ( 
.A(n_288),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_292),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_294),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_294),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_296),
.Y(n_350)
);

HB1xp67_ASAP7_75t_L g351 ( 
.A(n_287),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_296),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_297),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_297),
.Y(n_354)
);

INVx2_ASAP7_75t_L g355 ( 
.A(n_269),
.Y(n_355)
);

CKINVDCx16_ASAP7_75t_R g356 ( 
.A(n_310),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_273),
.Y(n_357)
);

BUFx2_ASAP7_75t_L g358 ( 
.A(n_314),
.Y(n_358)
);

CKINVDCx16_ASAP7_75t_R g359 ( 
.A(n_304),
.Y(n_359)
);

INVxp67_ASAP7_75t_L g360 ( 
.A(n_308),
.Y(n_360)
);

CKINVDCx20_ASAP7_75t_R g361 ( 
.A(n_272),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_274),
.Y(n_362)
);

BUFx3_ASAP7_75t_L g363 ( 
.A(n_287),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_273),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_315),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_315),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_316),
.Y(n_367)
);

CKINVDCx20_ASAP7_75t_R g368 ( 
.A(n_361),
.Y(n_368)
);

INVxp67_ASAP7_75t_L g369 ( 
.A(n_332),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_L g370 ( 
.A(n_346),
.B(n_277),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_R g371 ( 
.A(n_328),
.B(n_278),
.Y(n_371)
);

INVx2_ASAP7_75t_L g372 ( 
.A(n_341),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_329),
.Y(n_373)
);

NOR2xp67_ASAP7_75t_L g374 ( 
.A(n_343),
.B(n_279),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_329),
.Y(n_375)
);

CKINVDCx16_ASAP7_75t_R g376 ( 
.A(n_356),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_330),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_330),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_362),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_334),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_321),
.Y(n_381)
);

CKINVDCx20_ASAP7_75t_R g382 ( 
.A(n_356),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_337),
.Y(n_383)
);

HB1xp67_ASAP7_75t_L g384 ( 
.A(n_360),
.Y(n_384)
);

INVxp67_ASAP7_75t_L g385 ( 
.A(n_351),
.Y(n_385)
);

NAND2xp33_ASAP7_75t_R g386 ( 
.A(n_358),
.B(n_307),
.Y(n_386)
);

CKINVDCx20_ASAP7_75t_R g387 ( 
.A(n_359),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_336),
.Y(n_388)
);

CKINVDCx20_ASAP7_75t_R g389 ( 
.A(n_359),
.Y(n_389)
);

INVxp67_ASAP7_75t_L g390 ( 
.A(n_333),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_337),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_338),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_338),
.Y(n_393)
);

INVxp67_ASAP7_75t_SL g394 ( 
.A(n_363),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_340),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_333),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_358),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_340),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_344),
.Y(n_399)
);

CKINVDCx20_ASAP7_75t_R g400 ( 
.A(n_335),
.Y(n_400)
);

HB1xp67_ASAP7_75t_L g401 ( 
.A(n_342),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_363),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_344),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_L g404 ( 
.A(n_319),
.B(n_281),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_363),
.Y(n_405)
);

CKINVDCx20_ASAP7_75t_R g406 ( 
.A(n_345),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_345),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_347),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_347),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_L g410 ( 
.A(n_348),
.B(n_283),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_348),
.Y(n_411)
);

CKINVDCx20_ASAP7_75t_R g412 ( 
.A(n_349),
.Y(n_412)
);

CKINVDCx20_ASAP7_75t_R g413 ( 
.A(n_349),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_350),
.Y(n_414)
);

INVx3_ASAP7_75t_L g415 ( 
.A(n_372),
.Y(n_415)
);

BUFx2_ASAP7_75t_L g416 ( 
.A(n_396),
.Y(n_416)
);

CKINVDCx6p67_ASAP7_75t_R g417 ( 
.A(n_368),
.Y(n_417)
);

OAI21x1_ASAP7_75t_L g418 ( 
.A1(n_372),
.A2(n_352),
.B(n_350),
.Y(n_418)
);

BUFx6f_ASAP7_75t_L g419 ( 
.A(n_373),
.Y(n_419)
);

AND2x6_ASAP7_75t_L g420 ( 
.A(n_375),
.B(n_352),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_377),
.Y(n_421)
);

AND2x2_ASAP7_75t_L g422 ( 
.A(n_370),
.B(n_285),
.Y(n_422)
);

INVx2_ASAP7_75t_L g423 ( 
.A(n_378),
.Y(n_423)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_383),
.Y(n_424)
);

OAI22x1_ASAP7_75t_R g425 ( 
.A1(n_382),
.A2(n_225),
.B1(n_215),
.B2(n_286),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_391),
.Y(n_426)
);

AOI22xp5_ASAP7_75t_L g427 ( 
.A1(n_400),
.A2(n_295),
.B1(n_298),
.B2(n_293),
.Y(n_427)
);

INVx2_ASAP7_75t_SL g428 ( 
.A(n_401),
.Y(n_428)
);

BUFx6f_ASAP7_75t_L g429 ( 
.A(n_392),
.Y(n_429)
);

OAI21x1_ASAP7_75t_L g430 ( 
.A1(n_393),
.A2(n_354),
.B(n_353),
.Y(n_430)
);

OAI22xp5_ASAP7_75t_L g431 ( 
.A1(n_402),
.A2(n_207),
.B1(n_204),
.B2(n_299),
.Y(n_431)
);

INVx2_ASAP7_75t_L g432 ( 
.A(n_395),
.Y(n_432)
);

INVx2_ASAP7_75t_L g433 ( 
.A(n_398),
.Y(n_433)
);

AOI22x1_ASAP7_75t_SL g434 ( 
.A1(n_379),
.A2(n_380),
.B1(n_389),
.B2(n_387),
.Y(n_434)
);

INVx3_ASAP7_75t_L g435 ( 
.A(n_399),
.Y(n_435)
);

AOI22xp5_ASAP7_75t_L g436 ( 
.A1(n_410),
.A2(n_300),
.B1(n_354),
.B2(n_353),
.Y(n_436)
);

BUFx2_ASAP7_75t_L g437 ( 
.A(n_396),
.Y(n_437)
);

CKINVDCx11_ASAP7_75t_R g438 ( 
.A(n_376),
.Y(n_438)
);

AOI22xp5_ASAP7_75t_L g439 ( 
.A1(n_407),
.A2(n_312),
.B1(n_366),
.B2(n_365),
.Y(n_439)
);

INVx2_ASAP7_75t_L g440 ( 
.A(n_403),
.Y(n_440)
);

CKINVDCx8_ASAP7_75t_R g441 ( 
.A(n_379),
.Y(n_441)
);

INVx2_ASAP7_75t_L g442 ( 
.A(n_408),
.Y(n_442)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_409),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_414),
.Y(n_444)
);

INVx2_ASAP7_75t_L g445 ( 
.A(n_407),
.Y(n_445)
);

BUFx6f_ASAP7_75t_L g446 ( 
.A(n_402),
.Y(n_446)
);

BUFx8_ASAP7_75t_L g447 ( 
.A(n_371),
.Y(n_447)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_411),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_394),
.B(n_357),
.Y(n_449)
);

AND2x4_ASAP7_75t_L g450 ( 
.A(n_390),
.B(n_357),
.Y(n_450)
);

AOI22xp5_ASAP7_75t_L g451 ( 
.A1(n_411),
.A2(n_312),
.B1(n_366),
.B2(n_365),
.Y(n_451)
);

OAI22x1_ASAP7_75t_L g452 ( 
.A1(n_397),
.A2(n_308),
.B1(n_236),
.B2(n_217),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_405),
.Y(n_453)
);

BUFx2_ASAP7_75t_L g454 ( 
.A(n_397),
.Y(n_454)
);

HB1xp67_ASAP7_75t_L g455 ( 
.A(n_406),
.Y(n_455)
);

OAI22xp5_ASAP7_75t_L g456 ( 
.A1(n_405),
.A2(n_202),
.B1(n_229),
.B2(n_367),
.Y(n_456)
);

BUFx6f_ASAP7_75t_L g457 ( 
.A(n_404),
.Y(n_457)
);

CKINVDCx5p33_ASAP7_75t_R g458 ( 
.A(n_380),
.Y(n_458)
);

INVx2_ASAP7_75t_L g459 ( 
.A(n_412),
.Y(n_459)
);

AND2x2_ASAP7_75t_SL g460 ( 
.A(n_384),
.B(n_202),
.Y(n_460)
);

AOI22xp5_ASAP7_75t_L g461 ( 
.A1(n_413),
.A2(n_367),
.B1(n_364),
.B2(n_311),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_385),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_369),
.Y(n_463)
);

BUFx6f_ASAP7_75t_L g464 ( 
.A(n_388),
.Y(n_464)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_388),
.Y(n_465)
);

INVx2_ASAP7_75t_L g466 ( 
.A(n_381),
.Y(n_466)
);

CKINVDCx20_ASAP7_75t_R g467 ( 
.A(n_381),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_374),
.Y(n_468)
);

INVx2_ASAP7_75t_L g469 ( 
.A(n_386),
.Y(n_469)
);

INVx5_ASAP7_75t_L g470 ( 
.A(n_372),
.Y(n_470)
);

CKINVDCx5p33_ASAP7_75t_R g471 ( 
.A(n_371),
.Y(n_471)
);

INVx2_ASAP7_75t_L g472 ( 
.A(n_372),
.Y(n_472)
);

INVx4_ASAP7_75t_L g473 ( 
.A(n_402),
.Y(n_473)
);

AND2x4_ASAP7_75t_L g474 ( 
.A(n_373),
.B(n_364),
.Y(n_474)
);

BUFx3_ASAP7_75t_L g475 ( 
.A(n_368),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_373),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_373),
.Y(n_477)
);

AND2x2_ASAP7_75t_L g478 ( 
.A(n_370),
.B(n_291),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_373),
.Y(n_479)
);

INVx2_ASAP7_75t_L g480 ( 
.A(n_372),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_373),
.Y(n_481)
);

AND2x2_ASAP7_75t_L g482 ( 
.A(n_370),
.B(n_305),
.Y(n_482)
);

INVxp67_ASAP7_75t_L g483 ( 
.A(n_401),
.Y(n_483)
);

BUFx12f_ASAP7_75t_L g484 ( 
.A(n_380),
.Y(n_484)
);

INVx2_ASAP7_75t_L g485 ( 
.A(n_372),
.Y(n_485)
);

BUFx6f_ASAP7_75t_L g486 ( 
.A(n_372),
.Y(n_486)
);

CKINVDCx5p33_ASAP7_75t_R g487 ( 
.A(n_371),
.Y(n_487)
);

INVx2_ASAP7_75t_L g488 ( 
.A(n_372),
.Y(n_488)
);

INVx2_ASAP7_75t_SL g489 ( 
.A(n_401),
.Y(n_489)
);

CKINVDCx11_ASAP7_75t_R g490 ( 
.A(n_387),
.Y(n_490)
);

BUFx6f_ASAP7_75t_L g491 ( 
.A(n_372),
.Y(n_491)
);

AND2x4_ASAP7_75t_L g492 ( 
.A(n_373),
.B(n_355),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_373),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_373),
.Y(n_494)
);

OAI22xp5_ASAP7_75t_L g495 ( 
.A1(n_402),
.A2(n_229),
.B1(n_196),
.B2(n_309),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_373),
.Y(n_496)
);

INVx5_ASAP7_75t_L g497 ( 
.A(n_372),
.Y(n_497)
);

HB1xp67_ASAP7_75t_L g498 ( 
.A(n_428),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_472),
.Y(n_499)
);

HB1xp67_ASAP7_75t_L g500 ( 
.A(n_489),
.Y(n_500)
);

AND2x2_ASAP7_75t_L g501 ( 
.A(n_482),
.B(n_355),
.Y(n_501)
);

AND2x4_ASAP7_75t_L g502 ( 
.A(n_423),
.B(n_331),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_472),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_480),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_457),
.B(n_331),
.Y(n_505)
);

HB1xp67_ASAP7_75t_L g506 ( 
.A(n_459),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_480),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_485),
.Y(n_508)
);

OA21x2_ASAP7_75t_L g509 ( 
.A1(n_418),
.A2(n_327),
.B(n_323),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_457),
.B(n_339),
.Y(n_510)
);

AND2x2_ASAP7_75t_L g511 ( 
.A(n_423),
.B(n_305),
.Y(n_511)
);

AND2x4_ASAP7_75t_L g512 ( 
.A(n_424),
.B(n_339),
.Y(n_512)
);

HB1xp67_ASAP7_75t_L g513 ( 
.A(n_459),
.Y(n_513)
);

AND2x4_ASAP7_75t_L g514 ( 
.A(n_424),
.B(n_306),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_485),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_457),
.B(n_327),
.Y(n_516)
);

AND2x4_ASAP7_75t_L g517 ( 
.A(n_432),
.B(n_306),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_457),
.B(n_322),
.Y(n_518)
);

BUFx2_ASAP7_75t_L g519 ( 
.A(n_455),
.Y(n_519)
);

INVx3_ASAP7_75t_L g520 ( 
.A(n_486),
.Y(n_520)
);

HB1xp67_ASAP7_75t_L g521 ( 
.A(n_483),
.Y(n_521)
);

AND2x2_ASAP7_75t_L g522 ( 
.A(n_432),
.B(n_320),
.Y(n_522)
);

INVx2_ASAP7_75t_L g523 ( 
.A(n_488),
.Y(n_523)
);

BUFx6f_ASAP7_75t_L g524 ( 
.A(n_486),
.Y(n_524)
);

BUFx6f_ASAP7_75t_L g525 ( 
.A(n_486),
.Y(n_525)
);

BUFx2_ASAP7_75t_L g526 ( 
.A(n_455),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_SL g527 ( 
.A(n_460),
.B(n_182),
.Y(n_527)
);

XNOR2xp5_ASAP7_75t_L g528 ( 
.A(n_431),
.B(n_199),
.Y(n_528)
);

AND2x4_ASAP7_75t_L g529 ( 
.A(n_433),
.B(n_179),
.Y(n_529)
);

BUFx6f_ASAP7_75t_L g530 ( 
.A(n_486),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_L g531 ( 
.A(n_478),
.B(n_322),
.Y(n_531)
);

AND2x2_ASAP7_75t_L g532 ( 
.A(n_433),
.B(n_320),
.Y(n_532)
);

AND2x6_ASAP7_75t_L g533 ( 
.A(n_419),
.B(n_180),
.Y(n_533)
);

INVx2_ASAP7_75t_L g534 ( 
.A(n_418),
.Y(n_534)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_415),
.Y(n_535)
);

INVx2_ASAP7_75t_L g536 ( 
.A(n_430),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_440),
.B(n_323),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_430),
.Y(n_538)
);

BUFx6f_ASAP7_75t_L g539 ( 
.A(n_491),
.Y(n_539)
);

INVx2_ASAP7_75t_L g540 ( 
.A(n_491),
.Y(n_540)
);

CKINVDCx5p33_ASAP7_75t_R g541 ( 
.A(n_471),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_440),
.Y(n_542)
);

BUFx6f_ASAP7_75t_L g543 ( 
.A(n_470),
.Y(n_543)
);

INVx2_ASAP7_75t_L g544 ( 
.A(n_442),
.Y(n_544)
);

AND2x4_ASAP7_75t_L g545 ( 
.A(n_442),
.B(n_187),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_443),
.Y(n_546)
);

AND2x2_ASAP7_75t_L g547 ( 
.A(n_506),
.B(n_445),
.Y(n_547)
);

AND2x2_ASAP7_75t_L g548 ( 
.A(n_513),
.B(n_445),
.Y(n_548)
);

AO22x2_ASAP7_75t_L g549 ( 
.A1(n_527),
.A2(n_448),
.B1(n_469),
.B2(n_466),
.Y(n_549)
);

AO22x2_ASAP7_75t_L g550 ( 
.A1(n_538),
.A2(n_448),
.B1(n_469),
.B2(n_466),
.Y(n_550)
);

NOR2xp33_ASAP7_75t_L g551 ( 
.A(n_528),
.B(n_422),
.Y(n_551)
);

INVx2_ASAP7_75t_L g552 ( 
.A(n_544),
.Y(n_552)
);

OAI22xp33_ASAP7_75t_L g553 ( 
.A1(n_519),
.A2(n_427),
.B1(n_436),
.B2(n_461),
.Y(n_553)
);

NAND2xp33_ASAP7_75t_SL g554 ( 
.A(n_541),
.B(n_446),
.Y(n_554)
);

OAI22xp33_ASAP7_75t_SL g555 ( 
.A1(n_519),
.A2(n_453),
.B1(n_495),
.B2(n_451),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_L g556 ( 
.A(n_501),
.B(n_460),
.Y(n_556)
);

INVx3_ASAP7_75t_L g557 ( 
.A(n_543),
.Y(n_557)
);

BUFx3_ASAP7_75t_L g558 ( 
.A(n_526),
.Y(n_558)
);

OAI22xp33_ASAP7_75t_SL g559 ( 
.A1(n_526),
.A2(n_439),
.B1(n_473),
.B2(n_421),
.Y(n_559)
);

AOI22xp5_ASAP7_75t_L g560 ( 
.A1(n_501),
.A2(n_450),
.B1(n_474),
.B2(n_435),
.Y(n_560)
);

AND2x2_ASAP7_75t_L g561 ( 
.A(n_521),
.B(n_454),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_SL g562 ( 
.A(n_498),
.B(n_446),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_544),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_SL g564 ( 
.A(n_500),
.B(n_446),
.Y(n_564)
);

AO22x2_ASAP7_75t_L g565 ( 
.A1(n_538),
.A2(n_456),
.B1(n_473),
.B2(n_443),
.Y(n_565)
);

OAI22xp5_ASAP7_75t_L g566 ( 
.A1(n_531),
.A2(n_473),
.B1(n_446),
.B2(n_419),
.Y(n_566)
);

AO22x2_ASAP7_75t_L g567 ( 
.A1(n_536),
.A2(n_426),
.B1(n_476),
.B2(n_444),
.Y(n_567)
);

OAI22xp5_ASAP7_75t_SL g568 ( 
.A1(n_528),
.A2(n_452),
.B1(n_467),
.B2(n_425),
.Y(n_568)
);

AND2x2_ASAP7_75t_L g569 ( 
.A(n_511),
.B(n_416),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_523),
.Y(n_570)
);

OA22x2_ASAP7_75t_L g571 ( 
.A1(n_542),
.A2(n_465),
.B1(n_463),
.B2(n_462),
.Y(n_571)
);

OR2x6_ASAP7_75t_L g572 ( 
.A(n_543),
.B(n_464),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_523),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_523),
.Y(n_574)
);

OAI22xp33_ASAP7_75t_SL g575 ( 
.A1(n_516),
.A2(n_479),
.B1(n_481),
.B2(n_477),
.Y(n_575)
);

AOI22xp5_ASAP7_75t_L g576 ( 
.A1(n_529),
.A2(n_450),
.B1(n_474),
.B2(n_435),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_499),
.Y(n_577)
);

AND2x2_ASAP7_75t_L g578 ( 
.A(n_511),
.B(n_437),
.Y(n_578)
);

AOI22xp5_ASAP7_75t_L g579 ( 
.A1(n_529),
.A2(n_450),
.B1(n_474),
.B2(n_493),
.Y(n_579)
);

AO22x2_ASAP7_75t_L g580 ( 
.A1(n_536),
.A2(n_534),
.B1(n_546),
.B2(n_542),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_499),
.Y(n_581)
);

NOR2xp33_ASAP7_75t_L g582 ( 
.A(n_518),
.B(n_471),
.Y(n_582)
);

NOR2xp33_ASAP7_75t_L g583 ( 
.A(n_505),
.B(n_487),
.Y(n_583)
);

AO22x2_ASAP7_75t_L g584 ( 
.A1(n_536),
.A2(n_496),
.B1(n_494),
.B2(n_465),
.Y(n_584)
);

OA22x2_ASAP7_75t_L g585 ( 
.A1(n_546),
.A2(n_458),
.B1(n_468),
.B2(n_487),
.Y(n_585)
);

AO22x2_ASAP7_75t_L g586 ( 
.A1(n_534),
.A2(n_434),
.B1(n_449),
.B2(n_475),
.Y(n_586)
);

OAI22xp33_ASAP7_75t_L g587 ( 
.A1(n_510),
.A2(n_441),
.B1(n_464),
.B2(n_458),
.Y(n_587)
);

OAI22xp5_ASAP7_75t_L g588 ( 
.A1(n_543),
.A2(n_419),
.B1(n_429),
.B2(n_497),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_580),
.Y(n_589)
);

BUFx6f_ASAP7_75t_L g590 ( 
.A(n_572),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_L g591 ( 
.A(n_582),
.B(n_514),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_L g592 ( 
.A(n_569),
.B(n_578),
.Y(n_592)
);

BUFx3_ASAP7_75t_L g593 ( 
.A(n_558),
.Y(n_593)
);

INVx2_ASAP7_75t_L g594 ( 
.A(n_570),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_570),
.Y(n_595)
);

INVx2_ASAP7_75t_L g596 ( 
.A(n_573),
.Y(n_596)
);

INVx4_ASAP7_75t_L g597 ( 
.A(n_572),
.Y(n_597)
);

INVx2_ASAP7_75t_L g598 ( 
.A(n_574),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_580),
.Y(n_599)
);

NAND2xp33_ASAP7_75t_L g600 ( 
.A(n_566),
.B(n_543),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_SL g601 ( 
.A(n_553),
.B(n_441),
.Y(n_601)
);

CKINVDCx6p67_ASAP7_75t_R g602 ( 
.A(n_561),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_567),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_567),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_L g605 ( 
.A(n_583),
.B(n_514),
.Y(n_605)
);

INVx2_ASAP7_75t_L g606 ( 
.A(n_552),
.Y(n_606)
);

INVx2_ASAP7_75t_SL g607 ( 
.A(n_547),
.Y(n_607)
);

INVx2_ASAP7_75t_L g608 ( 
.A(n_563),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_SL g609 ( 
.A(n_556),
.B(n_464),
.Y(n_609)
);

INVx8_ASAP7_75t_L g610 ( 
.A(n_557),
.Y(n_610)
);

INVx2_ASAP7_75t_L g611 ( 
.A(n_577),
.Y(n_611)
);

INVxp67_ASAP7_75t_SL g612 ( 
.A(n_548),
.Y(n_612)
);

INVx2_ASAP7_75t_L g613 ( 
.A(n_577),
.Y(n_613)
);

OR2x2_ASAP7_75t_L g614 ( 
.A(n_581),
.B(n_529),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_581),
.Y(n_615)
);

NAND2xp33_ASAP7_75t_L g616 ( 
.A(n_576),
.B(n_543),
.Y(n_616)
);

BUFx10_ASAP7_75t_L g617 ( 
.A(n_551),
.Y(n_617)
);

INVx2_ASAP7_75t_SL g618 ( 
.A(n_571),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_SL g619 ( 
.A(n_587),
.B(n_464),
.Y(n_619)
);

OAI21xp33_ASAP7_75t_SL g620 ( 
.A1(n_579),
.A2(n_504),
.B(n_503),
.Y(n_620)
);

INVx2_ASAP7_75t_L g621 ( 
.A(n_584),
.Y(n_621)
);

NOR2xp33_ASAP7_75t_L g622 ( 
.A(n_568),
.B(n_475),
.Y(n_622)
);

BUFx3_ASAP7_75t_L g623 ( 
.A(n_557),
.Y(n_623)
);

NAND3xp33_ASAP7_75t_L g624 ( 
.A(n_579),
.B(n_447),
.C(n_438),
.Y(n_624)
);

INVx2_ASAP7_75t_L g625 ( 
.A(n_584),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_550),
.Y(n_626)
);

AND2x2_ASAP7_75t_L g627 ( 
.A(n_560),
.B(n_529),
.Y(n_627)
);

INVx2_ASAP7_75t_L g628 ( 
.A(n_550),
.Y(n_628)
);

INVx2_ASAP7_75t_L g629 ( 
.A(n_565),
.Y(n_629)
);

BUFx3_ASAP7_75t_L g630 ( 
.A(n_585),
.Y(n_630)
);

INVx2_ASAP7_75t_L g631 ( 
.A(n_565),
.Y(n_631)
);

NOR2xp33_ASAP7_75t_L g632 ( 
.A(n_568),
.B(n_467),
.Y(n_632)
);

HB1xp67_ASAP7_75t_L g633 ( 
.A(n_562),
.Y(n_633)
);

INVx2_ASAP7_75t_L g634 ( 
.A(n_560),
.Y(n_634)
);

INVx2_ASAP7_75t_L g635 ( 
.A(n_576),
.Y(n_635)
);

BUFx2_ASAP7_75t_L g636 ( 
.A(n_549),
.Y(n_636)
);

BUFx6f_ASAP7_75t_L g637 ( 
.A(n_564),
.Y(n_637)
);

INVx2_ASAP7_75t_L g638 ( 
.A(n_549),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_575),
.Y(n_639)
);

BUFx2_ASAP7_75t_L g640 ( 
.A(n_554),
.Y(n_640)
);

INVxp67_ASAP7_75t_SL g641 ( 
.A(n_588),
.Y(n_641)
);

CKINVDCx20_ASAP7_75t_R g642 ( 
.A(n_586),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_559),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_L g644 ( 
.A(n_555),
.B(n_514),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_586),
.Y(n_645)
);

INVx2_ASAP7_75t_L g646 ( 
.A(n_570),
.Y(n_646)
);

BUFx6f_ASAP7_75t_L g647 ( 
.A(n_572),
.Y(n_647)
);

INVx2_ASAP7_75t_L g648 ( 
.A(n_570),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_580),
.Y(n_649)
);

BUFx3_ASAP7_75t_L g650 ( 
.A(n_558),
.Y(n_650)
);

AOI22xp5_ASAP7_75t_L g651 ( 
.A1(n_551),
.A2(n_438),
.B1(n_447),
.B2(n_417),
.Y(n_651)
);

INVx2_ASAP7_75t_L g652 ( 
.A(n_570),
.Y(n_652)
);

INVx2_ASAP7_75t_L g653 ( 
.A(n_570),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_580),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_SL g655 ( 
.A(n_582),
.B(n_419),
.Y(n_655)
);

NAND3xp33_ASAP7_75t_L g656 ( 
.A(n_551),
.B(n_447),
.C(n_490),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_577),
.Y(n_657)
);

AND3x2_ASAP7_75t_L g658 ( 
.A(n_551),
.B(n_545),
.C(n_517),
.Y(n_658)
);

OR2x6_ASAP7_75t_L g659 ( 
.A(n_567),
.B(n_534),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_SL g660 ( 
.A(n_582),
.B(n_429),
.Y(n_660)
);

NAND2xp33_ASAP7_75t_L g661 ( 
.A(n_566),
.B(n_543),
.Y(n_661)
);

CKINVDCx5p33_ASAP7_75t_R g662 ( 
.A(n_558),
.Y(n_662)
);

BUFx4f_ASAP7_75t_L g663 ( 
.A(n_572),
.Y(n_663)
);

INVx4_ASAP7_75t_L g664 ( 
.A(n_572),
.Y(n_664)
);

AND3x2_ASAP7_75t_L g665 ( 
.A(n_551),
.B(n_545),
.C(n_517),
.Y(n_665)
);

INVx2_ASAP7_75t_L g666 ( 
.A(n_570),
.Y(n_666)
);

INVx2_ASAP7_75t_L g667 ( 
.A(n_570),
.Y(n_667)
);

INVx1_ASAP7_75t_SL g668 ( 
.A(n_561),
.Y(n_668)
);

AND2x2_ASAP7_75t_L g669 ( 
.A(n_552),
.B(n_545),
.Y(n_669)
);

BUFx3_ASAP7_75t_L g670 ( 
.A(n_558),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_577),
.Y(n_671)
);

BUFx3_ASAP7_75t_L g672 ( 
.A(n_558),
.Y(n_672)
);

INVx2_ASAP7_75t_L g673 ( 
.A(n_570),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_582),
.B(n_514),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_615),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_639),
.B(n_503),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_SL g677 ( 
.A(n_591),
.B(n_429),
.Y(n_677)
);

BUFx4f_ASAP7_75t_L g678 ( 
.A(n_602),
.Y(n_678)
);

OR2x2_ASAP7_75t_SL g679 ( 
.A(n_656),
.B(n_192),
.Y(n_679)
);

INVxp33_ASAP7_75t_L g680 ( 
.A(n_592),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_657),
.Y(n_681)
);

INVx4_ASAP7_75t_L g682 ( 
.A(n_662),
.Y(n_682)
);

BUFx3_ASAP7_75t_L g683 ( 
.A(n_593),
.Y(n_683)
);

AND2x2_ASAP7_75t_L g684 ( 
.A(n_607),
.B(n_545),
.Y(n_684)
);

INVx2_ASAP7_75t_L g685 ( 
.A(n_611),
.Y(n_685)
);

AND2x4_ASAP7_75t_L g686 ( 
.A(n_597),
.B(n_540),
.Y(n_686)
);

INVx2_ASAP7_75t_SL g687 ( 
.A(n_662),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_671),
.Y(n_688)
);

NOR2xp33_ASAP7_75t_L g689 ( 
.A(n_674),
.B(n_429),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_611),
.Y(n_690)
);

CKINVDCx5p33_ASAP7_75t_R g691 ( 
.A(n_602),
.Y(n_691)
);

INVx3_ASAP7_75t_L g692 ( 
.A(n_623),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_L g693 ( 
.A(n_639),
.B(n_504),
.Y(n_693)
);

HB1xp67_ASAP7_75t_L g694 ( 
.A(n_659),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_613),
.Y(n_695)
);

INVx1_ASAP7_75t_SL g696 ( 
.A(n_607),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_613),
.Y(n_697)
);

AND2x2_ASAP7_75t_L g698 ( 
.A(n_668),
.B(n_517),
.Y(n_698)
);

BUFx4f_ASAP7_75t_L g699 ( 
.A(n_590),
.Y(n_699)
);

INVx2_ASAP7_75t_L g700 ( 
.A(n_606),
.Y(n_700)
);

BUFx6f_ASAP7_75t_L g701 ( 
.A(n_593),
.Y(n_701)
);

INVx2_ASAP7_75t_SL g702 ( 
.A(n_650),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_589),
.Y(n_703)
);

INVx4_ASAP7_75t_L g704 ( 
.A(n_610),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_L g705 ( 
.A(n_634),
.B(n_507),
.Y(n_705)
);

NOR2xp33_ASAP7_75t_L g706 ( 
.A(n_601),
.B(n_517),
.Y(n_706)
);

INVx2_ASAP7_75t_L g707 ( 
.A(n_606),
.Y(n_707)
);

AND2x2_ASAP7_75t_L g708 ( 
.A(n_612),
.B(n_512),
.Y(n_708)
);

INVx2_ASAP7_75t_L g709 ( 
.A(n_608),
.Y(n_709)
);

AND2x2_ASAP7_75t_L g710 ( 
.A(n_605),
.B(n_512),
.Y(n_710)
);

OAI22xp33_ASAP7_75t_SL g711 ( 
.A1(n_619),
.A2(n_203),
.B1(n_210),
.B2(n_200),
.Y(n_711)
);

NOR2xp33_ASAP7_75t_L g712 ( 
.A(n_609),
.B(n_417),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_589),
.Y(n_713)
);

INVxp67_ASAP7_75t_SL g714 ( 
.A(n_603),
.Y(n_714)
);

CKINVDCx11_ASAP7_75t_R g715 ( 
.A(n_617),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_599),
.Y(n_716)
);

INVx4_ASAP7_75t_L g717 ( 
.A(n_610),
.Y(n_717)
);

OR2x6_ASAP7_75t_L g718 ( 
.A(n_659),
.B(n_634),
.Y(n_718)
);

NOR2xp33_ASAP7_75t_L g719 ( 
.A(n_655),
.B(n_540),
.Y(n_719)
);

AND2x4_ASAP7_75t_L g720 ( 
.A(n_597),
.B(n_540),
.Y(n_720)
);

AND2x2_ASAP7_75t_L g721 ( 
.A(n_643),
.B(n_512),
.Y(n_721)
);

BUFx10_ASAP7_75t_L g722 ( 
.A(n_622),
.Y(n_722)
);

BUFx10_ASAP7_75t_L g723 ( 
.A(n_632),
.Y(n_723)
);

NOR2xp33_ASAP7_75t_L g724 ( 
.A(n_660),
.B(n_520),
.Y(n_724)
);

INVx2_ASAP7_75t_SL g725 ( 
.A(n_650),
.Y(n_725)
);

INVx2_ASAP7_75t_SL g726 ( 
.A(n_670),
.Y(n_726)
);

BUFx6f_ASAP7_75t_L g727 ( 
.A(n_670),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_SL g728 ( 
.A(n_640),
.B(n_502),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_L g729 ( 
.A(n_635),
.B(n_643),
.Y(n_729)
);

OR2x6_ASAP7_75t_L g730 ( 
.A(n_659),
.B(n_524),
.Y(n_730)
);

AND2x4_ASAP7_75t_L g731 ( 
.A(n_597),
.B(n_520),
.Y(n_731)
);

OAI21xp33_ASAP7_75t_L g732 ( 
.A1(n_644),
.A2(n_195),
.B(n_185),
.Y(n_732)
);

INVx4_ASAP7_75t_L g733 ( 
.A(n_610),
.Y(n_733)
);

INVx4_ASAP7_75t_L g734 ( 
.A(n_610),
.Y(n_734)
);

INVx2_ASAP7_75t_L g735 ( 
.A(n_596),
.Y(n_735)
);

INVx2_ASAP7_75t_L g736 ( 
.A(n_596),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_599),
.Y(n_737)
);

INVx3_ASAP7_75t_L g738 ( 
.A(n_623),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_649),
.Y(n_739)
);

OR2x2_ASAP7_75t_L g740 ( 
.A(n_614),
.B(n_508),
.Y(n_740)
);

AND2x2_ASAP7_75t_L g741 ( 
.A(n_618),
.B(n_512),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_649),
.Y(n_742)
);

BUFx2_ASAP7_75t_L g743 ( 
.A(n_672),
.Y(n_743)
);

NOR2xp33_ASAP7_75t_L g744 ( 
.A(n_618),
.B(n_520),
.Y(n_744)
);

NOR2xp33_ASAP7_75t_L g745 ( 
.A(n_633),
.B(n_520),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_654),
.Y(n_746)
);

INVx2_ASAP7_75t_L g747 ( 
.A(n_598),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_594),
.B(n_508),
.Y(n_748)
);

OR2x2_ASAP7_75t_L g749 ( 
.A(n_614),
.B(n_515),
.Y(n_749)
);

NOR2xp33_ASAP7_75t_L g750 ( 
.A(n_630),
.B(n_535),
.Y(n_750)
);

BUFx3_ASAP7_75t_L g751 ( 
.A(n_672),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_654),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_603),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_604),
.Y(n_754)
);

AND2x2_ASAP7_75t_L g755 ( 
.A(n_669),
.B(n_502),
.Y(n_755)
);

AOI22xp33_ASAP7_75t_L g756 ( 
.A1(n_642),
.A2(n_194),
.B1(n_195),
.B2(n_219),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_604),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_L g758 ( 
.A(n_594),
.B(n_515),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_729),
.B(n_636),
.Y(n_759)
);

NAND2xp33_ASAP7_75t_L g760 ( 
.A(n_756),
.B(n_637),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_729),
.B(n_636),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_703),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_675),
.B(n_638),
.Y(n_763)
);

AND2x4_ASAP7_75t_L g764 ( 
.A(n_730),
.B(n_621),
.Y(n_764)
);

NAND3xp33_ASAP7_75t_L g765 ( 
.A(n_756),
.B(n_624),
.C(n_645),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_713),
.Y(n_766)
);

AOI22xp33_ASAP7_75t_L g767 ( 
.A1(n_732),
.A2(n_642),
.B1(n_645),
.B2(n_630),
.Y(n_767)
);

INVx2_ASAP7_75t_SL g768 ( 
.A(n_701),
.Y(n_768)
);

INVx2_ASAP7_75t_SL g769 ( 
.A(n_701),
.Y(n_769)
);

NOR2xp33_ASAP7_75t_L g770 ( 
.A(n_680),
.B(n_617),
.Y(n_770)
);

NAND3xp33_ASAP7_75t_L g771 ( 
.A(n_706),
.B(n_665),
.C(n_658),
.Y(n_771)
);

INVx2_ASAP7_75t_L g772 ( 
.A(n_685),
.Y(n_772)
);

NOR2xp33_ASAP7_75t_L g773 ( 
.A(n_680),
.B(n_617),
.Y(n_773)
);

NOR3xp33_ASAP7_75t_L g774 ( 
.A(n_711),
.B(n_640),
.C(n_664),
.Y(n_774)
);

NAND3xp33_ASAP7_75t_L g775 ( 
.A(n_706),
.B(n_637),
.C(n_638),
.Y(n_775)
);

INVx2_ASAP7_75t_L g776 ( 
.A(n_681),
.Y(n_776)
);

AND2x2_ASAP7_75t_L g777 ( 
.A(n_696),
.B(n_627),
.Y(n_777)
);

NOR2xp33_ASAP7_75t_L g778 ( 
.A(n_687),
.B(n_490),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_L g779 ( 
.A(n_696),
.B(n_627),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_688),
.B(n_716),
.Y(n_780)
);

INVx2_ASAP7_75t_L g781 ( 
.A(n_700),
.Y(n_781)
);

BUFx3_ASAP7_75t_L g782 ( 
.A(n_701),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_737),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_739),
.B(n_621),
.Y(n_784)
);

AND2x2_ASAP7_75t_L g785 ( 
.A(n_698),
.B(n_637),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_SL g786 ( 
.A(n_678),
.B(n_637),
.Y(n_786)
);

BUFx6f_ASAP7_75t_L g787 ( 
.A(n_727),
.Y(n_787)
);

INVxp33_ASAP7_75t_L g788 ( 
.A(n_715),
.Y(n_788)
);

BUFx12f_ASAP7_75t_L g789 ( 
.A(n_691),
.Y(n_789)
);

INVxp33_ASAP7_75t_L g790 ( 
.A(n_727),
.Y(n_790)
);

NOR2xp33_ASAP7_75t_L g791 ( 
.A(n_682),
.B(n_722),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_SL g792 ( 
.A(n_678),
.B(n_637),
.Y(n_792)
);

NOR2xp33_ASAP7_75t_L g793 ( 
.A(n_682),
.B(n_651),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_742),
.Y(n_794)
);

NOR2xp33_ASAP7_75t_L g795 ( 
.A(n_722),
.B(n_484),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_L g796 ( 
.A(n_746),
.B(n_625),
.Y(n_796)
);

NOR3xp33_ASAP7_75t_L g797 ( 
.A(n_712),
.B(n_664),
.C(n_661),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_752),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_714),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_L g800 ( 
.A(n_690),
.B(n_625),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_L g801 ( 
.A(n_695),
.B(n_697),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_714),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_753),
.Y(n_803)
);

INVx2_ASAP7_75t_L g804 ( 
.A(n_707),
.Y(n_804)
);

BUFx3_ASAP7_75t_L g805 ( 
.A(n_727),
.Y(n_805)
);

NOR3xp33_ASAP7_75t_L g806 ( 
.A(n_712),
.B(n_689),
.C(n_677),
.Y(n_806)
);

INVx2_ASAP7_75t_L g807 ( 
.A(n_709),
.Y(n_807)
);

NOR2xp33_ASAP7_75t_L g808 ( 
.A(n_723),
.B(n_679),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_L g809 ( 
.A(n_754),
.B(n_626),
.Y(n_809)
);

INVxp67_ASAP7_75t_L g810 ( 
.A(n_743),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_L g811 ( 
.A(n_757),
.B(n_626),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_676),
.Y(n_812)
);

BUFx6f_ASAP7_75t_L g813 ( 
.A(n_683),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_L g814 ( 
.A(n_676),
.B(n_629),
.Y(n_814)
);

BUFx6f_ASAP7_75t_L g815 ( 
.A(n_751),
.Y(n_815)
);

NAND2xp33_ASAP7_75t_L g816 ( 
.A(n_702),
.B(n_590),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_L g817 ( 
.A(n_693),
.B(n_629),
.Y(n_817)
);

AOI221xp5_ASAP7_75t_L g818 ( 
.A1(n_689),
.A2(n_222),
.B1(n_227),
.B2(n_213),
.C(n_208),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_SL g819 ( 
.A(n_723),
.B(n_663),
.Y(n_819)
);

NOR2xp33_ASAP7_75t_SL g820 ( 
.A(n_704),
.B(n_484),
.Y(n_820)
);

INVx2_ASAP7_75t_L g821 ( 
.A(n_735),
.Y(n_821)
);

BUFx6f_ASAP7_75t_L g822 ( 
.A(n_725),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_693),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_L g824 ( 
.A(n_677),
.B(n_736),
.Y(n_824)
);

NOR2xp67_ASAP7_75t_SL g825 ( 
.A(n_704),
.B(n_590),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_694),
.Y(n_826)
);

INVx2_ASAP7_75t_L g827 ( 
.A(n_747),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_SL g828 ( 
.A(n_726),
.B(n_663),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_SL g829 ( 
.A(n_699),
.B(n_663),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_694),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_718),
.Y(n_831)
);

AOI22xp33_ASAP7_75t_L g832 ( 
.A1(n_760),
.A2(n_710),
.B1(n_194),
.B2(n_721),
.Y(n_832)
);

INVx2_ASAP7_75t_SL g833 ( 
.A(n_813),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_812),
.B(n_719),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_SL g835 ( 
.A(n_774),
.B(n_699),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_L g836 ( 
.A(n_823),
.B(n_719),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_780),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_777),
.B(n_708),
.Y(n_838)
);

AND2x4_ASAP7_75t_L g839 ( 
.A(n_831),
.B(n_730),
.Y(n_839)
);

NOR2xp33_ASAP7_75t_L g840 ( 
.A(n_770),
.B(n_692),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_L g841 ( 
.A(n_779),
.B(n_806),
.Y(n_841)
);

BUFx3_ASAP7_75t_L g842 ( 
.A(n_813),
.Y(n_842)
);

AND2x2_ASAP7_75t_L g843 ( 
.A(n_810),
.B(n_718),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_L g844 ( 
.A(n_773),
.B(n_684),
.Y(n_844)
);

INVxp67_ASAP7_75t_L g845 ( 
.A(n_780),
.Y(n_845)
);

CKINVDCx5p33_ASAP7_75t_R g846 ( 
.A(n_789),
.Y(n_846)
);

NOR2xp33_ASAP7_75t_L g847 ( 
.A(n_808),
.B(n_692),
.Y(n_847)
);

INVx2_ASAP7_75t_L g848 ( 
.A(n_776),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_762),
.Y(n_849)
);

INVx2_ASAP7_75t_L g850 ( 
.A(n_772),
.Y(n_850)
);

NOR2xp67_ASAP7_75t_L g851 ( 
.A(n_791),
.B(n_717),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_SL g852 ( 
.A(n_771),
.B(n_717),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_L g853 ( 
.A(n_759),
.B(n_761),
.Y(n_853)
);

INVxp67_ASAP7_75t_L g854 ( 
.A(n_826),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_L g855 ( 
.A(n_759),
.B(n_631),
.Y(n_855)
);

NOR2xp33_ASAP7_75t_L g856 ( 
.A(n_790),
.B(n_765),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_761),
.B(n_631),
.Y(n_857)
);

HB1xp67_ASAP7_75t_L g858 ( 
.A(n_799),
.Y(n_858)
);

INVx2_ASAP7_75t_L g859 ( 
.A(n_766),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_L g860 ( 
.A(n_824),
.B(n_718),
.Y(n_860)
);

INVx2_ASAP7_75t_SL g861 ( 
.A(n_813),
.Y(n_861)
);

AOI22xp33_ASAP7_75t_L g862 ( 
.A1(n_818),
.A2(n_755),
.B1(n_193),
.B2(n_205),
.Y(n_862)
);

OR2x6_ASAP7_75t_L g863 ( 
.A(n_775),
.B(n_730),
.Y(n_863)
);

BUFx3_ASAP7_75t_L g864 ( 
.A(n_815),
.Y(n_864)
);

OAI22xp33_ASAP7_75t_L g865 ( 
.A1(n_788),
.A2(n_728),
.B1(n_641),
.B2(n_659),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_L g866 ( 
.A(n_824),
.B(n_724),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_814),
.B(n_724),
.Y(n_867)
);

NOR2xp33_ASAP7_75t_L g868 ( 
.A(n_793),
.B(n_738),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_L g869 ( 
.A(n_814),
.B(n_745),
.Y(n_869)
);

NOR2xp33_ASAP7_75t_L g870 ( 
.A(n_795),
.B(n_738),
.Y(n_870)
);

NOR2xp33_ASAP7_75t_L g871 ( 
.A(n_819),
.B(n_728),
.Y(n_871)
);

NOR3xp33_ASAP7_75t_L g872 ( 
.A(n_797),
.B(n_750),
.C(n_744),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_783),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_794),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_L g875 ( 
.A(n_817),
.B(n_745),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_817),
.B(n_628),
.Y(n_876)
);

INVx2_ASAP7_75t_SL g877 ( 
.A(n_815),
.Y(n_877)
);

INVxp67_ASAP7_75t_L g878 ( 
.A(n_830),
.Y(n_878)
);

INVx2_ASAP7_75t_L g879 ( 
.A(n_798),
.Y(n_879)
);

INVxp67_ASAP7_75t_SL g880 ( 
.A(n_802),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_803),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_L g882 ( 
.A(n_801),
.B(n_628),
.Y(n_882)
);

INVx2_ASAP7_75t_L g883 ( 
.A(n_781),
.Y(n_883)
);

NOR2xp33_ASAP7_75t_L g884 ( 
.A(n_815),
.B(n_750),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_809),
.Y(n_885)
);

AOI22xp5_ASAP7_75t_L g886 ( 
.A1(n_767),
.A2(n_828),
.B1(n_820),
.B2(n_786),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_809),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_801),
.B(n_740),
.Y(n_888)
);

NOR2xp67_ASAP7_75t_L g889 ( 
.A(n_768),
.B(n_769),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_L g890 ( 
.A(n_804),
.B(n_749),
.Y(n_890)
);

INVx2_ASAP7_75t_L g891 ( 
.A(n_807),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_811),
.Y(n_892)
);

NOR2xp33_ASAP7_75t_L g893 ( 
.A(n_778),
.B(n_733),
.Y(n_893)
);

NAND2x1_ASAP7_75t_L g894 ( 
.A(n_825),
.B(n_733),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_L g895 ( 
.A(n_821),
.B(n_705),
.Y(n_895)
);

NOR2xp33_ASAP7_75t_L g896 ( 
.A(n_822),
.B(n_734),
.Y(n_896)
);

INVxp67_ASAP7_75t_L g897 ( 
.A(n_811),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_L g898 ( 
.A(n_827),
.B(n_705),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_SL g899 ( 
.A(n_822),
.B(n_734),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_L g900 ( 
.A(n_785),
.B(n_620),
.Y(n_900)
);

INVx2_ASAP7_75t_L g901 ( 
.A(n_800),
.Y(n_901)
);

AND2x2_ASAP7_75t_L g902 ( 
.A(n_782),
.B(n_686),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_L g903 ( 
.A(n_763),
.B(n_748),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_SL g904 ( 
.A(n_822),
.B(n_686),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_L g905 ( 
.A(n_763),
.B(n_748),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_784),
.Y(n_906)
);

INVx2_ASAP7_75t_SL g907 ( 
.A(n_787),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_L g908 ( 
.A(n_800),
.B(n_758),
.Y(n_908)
);

AND2x4_ASAP7_75t_L g909 ( 
.A(n_839),
.B(n_843),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_858),
.Y(n_910)
);

AO22x2_ASAP7_75t_L g911 ( 
.A1(n_849),
.A2(n_784),
.B1(n_796),
.B2(n_764),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_858),
.Y(n_912)
);

INVx2_ASAP7_75t_L g913 ( 
.A(n_837),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_873),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_L g915 ( 
.A(n_897),
.B(n_845),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_874),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_881),
.Y(n_917)
);

OAI221xp5_ASAP7_75t_L g918 ( 
.A1(n_852),
.A2(n_792),
.B1(n_816),
.B2(n_796),
.C(n_805),
.Y(n_918)
);

OR2x2_ASAP7_75t_SL g919 ( 
.A(n_841),
.B(n_787),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_859),
.Y(n_920)
);

OAI221xp5_ASAP7_75t_L g921 ( 
.A1(n_832),
.A2(n_829),
.B1(n_787),
.B2(n_744),
.C(n_616),
.Y(n_921)
);

BUFx8_ASAP7_75t_L g922 ( 
.A(n_833),
.Y(n_922)
);

CKINVDCx16_ASAP7_75t_R g923 ( 
.A(n_842),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_879),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_L g925 ( 
.A(n_853),
.B(n_764),
.Y(n_925)
);

OAI221xp5_ASAP7_75t_L g926 ( 
.A1(n_832),
.A2(n_616),
.B1(n_234),
.B2(n_182),
.C(n_183),
.Y(n_926)
);

CKINVDCx5p33_ASAP7_75t_R g927 ( 
.A(n_846),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_880),
.Y(n_928)
);

AO22x2_ASAP7_75t_L g929 ( 
.A1(n_880),
.A2(n_885),
.B1(n_892),
.B2(n_887),
.Y(n_929)
);

AOI22xp5_ASAP7_75t_L g930 ( 
.A1(n_862),
.A2(n_872),
.B1(n_856),
.B2(n_865),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_854),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_854),
.Y(n_932)
);

NAND3xp33_ASAP7_75t_L g933 ( 
.A(n_856),
.B(n_180),
.C(n_741),
.Y(n_933)
);

AO22x2_ASAP7_75t_L g934 ( 
.A1(n_906),
.A2(n_720),
.B1(n_664),
.B2(n_731),
.Y(n_934)
);

OAI22xp33_ASAP7_75t_L g935 ( 
.A1(n_886),
.A2(n_590),
.B1(n_647),
.B2(n_758),
.Y(n_935)
);

AO22x2_ASAP7_75t_L g936 ( 
.A1(n_845),
.A2(n_720),
.B1(n_731),
.B2(n_646),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_878),
.Y(n_937)
);

OAI221xp5_ASAP7_75t_L g938 ( 
.A1(n_835),
.A2(n_234),
.B1(n_183),
.B2(n_235),
.C(n_233),
.Y(n_938)
);

AOI22xp33_ASAP7_75t_L g939 ( 
.A1(n_872),
.A2(n_600),
.B1(n_661),
.B2(n_180),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_878),
.Y(n_940)
);

AND2x4_ASAP7_75t_L g941 ( 
.A(n_839),
.B(n_590),
.Y(n_941)
);

INVx2_ASAP7_75t_L g942 ( 
.A(n_848),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_901),
.Y(n_943)
);

INVx5_ASAP7_75t_L g944 ( 
.A(n_863),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_L g945 ( 
.A(n_897),
.B(n_595),
.Y(n_945)
);

INVx2_ASAP7_75t_L g946 ( 
.A(n_850),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_883),
.Y(n_947)
);

INVx2_ASAP7_75t_L g948 ( 
.A(n_891),
.Y(n_948)
);

INVx3_ASAP7_75t_L g949 ( 
.A(n_864),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_890),
.Y(n_950)
);

INVx2_ASAP7_75t_L g951 ( 
.A(n_860),
.Y(n_951)
);

INVx2_ASAP7_75t_L g952 ( 
.A(n_866),
.Y(n_952)
);

INVx2_ASAP7_75t_L g953 ( 
.A(n_861),
.Y(n_953)
);

INVx2_ASAP7_75t_L g954 ( 
.A(n_877),
.Y(n_954)
);

NOR2xp67_ASAP7_75t_L g955 ( 
.A(n_851),
.B(n_595),
.Y(n_955)
);

AND2x4_ASAP7_75t_L g956 ( 
.A(n_889),
.B(n_647),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_895),
.Y(n_957)
);

INVx1_ASAP7_75t_L g958 ( 
.A(n_898),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_L g959 ( 
.A(n_869),
.B(n_646),
.Y(n_959)
);

INVx2_ASAP7_75t_L g960 ( 
.A(n_907),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_888),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_834),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_836),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_L g964 ( 
.A(n_962),
.B(n_875),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_SL g965 ( 
.A(n_944),
.B(n_865),
.Y(n_965)
);

OAI21xp33_ASAP7_75t_L g966 ( 
.A1(n_930),
.A2(n_871),
.B(n_867),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_SL g967 ( 
.A(n_944),
.B(n_868),
.Y(n_967)
);

INVx5_ASAP7_75t_L g968 ( 
.A(n_944),
.Y(n_968)
);

CKINVDCx8_ASAP7_75t_R g969 ( 
.A(n_927),
.Y(n_969)
);

A2O1A1Ixp33_ASAP7_75t_L g970 ( 
.A1(n_930),
.A2(n_871),
.B(n_862),
.C(n_847),
.Y(n_970)
);

OAI21xp33_ASAP7_75t_L g971 ( 
.A1(n_933),
.A2(n_900),
.B(n_857),
.Y(n_971)
);

OAI22xp5_ASAP7_75t_L g972 ( 
.A1(n_939),
.A2(n_863),
.B1(n_884),
.B2(n_844),
.Y(n_972)
);

BUFx6f_ASAP7_75t_L g973 ( 
.A(n_956),
.Y(n_973)
);

AOI21xp5_ASAP7_75t_L g974 ( 
.A1(n_933),
.A2(n_894),
.B(n_863),
.Y(n_974)
);

AND2x4_ASAP7_75t_L g975 ( 
.A(n_909),
.B(n_904),
.Y(n_975)
);

AOI22xp33_ASAP7_75t_L g976 ( 
.A1(n_926),
.A2(n_840),
.B1(n_870),
.B2(n_893),
.Y(n_976)
);

INVx4_ASAP7_75t_L g977 ( 
.A(n_923),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_914),
.Y(n_978)
);

NAND2xp5_ASAP7_75t_L g979 ( 
.A(n_963),
.B(n_855),
.Y(n_979)
);

BUFx6f_ASAP7_75t_L g980 ( 
.A(n_956),
.Y(n_980)
);

AO21x1_ASAP7_75t_L g981 ( 
.A1(n_915),
.A2(n_899),
.B(n_896),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_L g982 ( 
.A(n_952),
.B(n_903),
.Y(n_982)
);

BUFx4f_ASAP7_75t_L g983 ( 
.A(n_949),
.Y(n_983)
);

OAI22xp5_ASAP7_75t_L g984 ( 
.A1(n_921),
.A2(n_919),
.B1(n_918),
.B2(n_923),
.Y(n_984)
);

OAI21xp5_ASAP7_75t_L g985 ( 
.A1(n_938),
.A2(n_915),
.B(n_935),
.Y(n_985)
);

A2O1A1Ixp33_ASAP7_75t_L g986 ( 
.A1(n_955),
.A2(n_905),
.B(n_876),
.C(n_838),
.Y(n_986)
);

BUFx4f_ASAP7_75t_L g987 ( 
.A(n_949),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_L g988 ( 
.A(n_961),
.B(n_908),
.Y(n_988)
);

A2O1A1Ixp33_ASAP7_75t_L g989 ( 
.A1(n_955),
.A2(n_882),
.B(n_902),
.C(n_600),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_SL g990 ( 
.A(n_950),
.B(n_647),
.Y(n_990)
);

AOI21xp5_ASAP7_75t_L g991 ( 
.A1(n_934),
.A2(n_669),
.B(n_647),
.Y(n_991)
);

NOR2xp33_ASAP7_75t_L g992 ( 
.A(n_909),
.B(n_0),
.Y(n_992)
);

O2A1O1Ixp33_ASAP7_75t_L g993 ( 
.A1(n_959),
.A2(n_0),
.B(n_1),
.C(n_2),
.Y(n_993)
);

AOI21xp5_ASAP7_75t_L g994 ( 
.A1(n_934),
.A2(n_647),
.B(n_648),
.Y(n_994)
);

AND2x2_ASAP7_75t_L g995 ( 
.A(n_951),
.B(n_673),
.Y(n_995)
);

AOI21xp33_ASAP7_75t_L g996 ( 
.A1(n_911),
.A2(n_2),
.B(n_3),
.Y(n_996)
);

INVx2_ASAP7_75t_L g997 ( 
.A(n_913),
.Y(n_997)
);

AOI21xp5_ASAP7_75t_L g998 ( 
.A1(n_911),
.A2(n_653),
.B(n_652),
.Y(n_998)
);

NOR2x1p5_ASAP7_75t_L g999 ( 
.A(n_925),
.B(n_957),
.Y(n_999)
);

OAI22xp5_ASAP7_75t_L g1000 ( 
.A1(n_958),
.A2(n_673),
.B1(n_667),
.B2(n_666),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_L g1001 ( 
.A(n_931),
.B(n_666),
.Y(n_1001)
);

AOI22xp33_ASAP7_75t_L g1002 ( 
.A1(n_941),
.A2(n_533),
.B1(n_420),
.B2(n_235),
.Y(n_1002)
);

O2A1O1Ixp33_ASAP7_75t_L g1003 ( 
.A1(n_932),
.A2(n_3),
.B(n_4),
.C(n_5),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_L g1004 ( 
.A(n_937),
.B(n_667),
.Y(n_1004)
);

INVx3_ASAP7_75t_L g1005 ( 
.A(n_922),
.Y(n_1005)
);

BUFx6f_ASAP7_75t_L g1006 ( 
.A(n_960),
.Y(n_1006)
);

AOI21xp5_ASAP7_75t_L g1007 ( 
.A1(n_936),
.A2(n_537),
.B(n_233),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_L g1008 ( 
.A(n_940),
.B(n_916),
.Y(n_1008)
);

INVx3_ASAP7_75t_L g1009 ( 
.A(n_922),
.Y(n_1009)
);

AOI21xp5_ASAP7_75t_L g1010 ( 
.A1(n_936),
.A2(n_232),
.B(n_230),
.Y(n_1010)
);

OAI321xp33_ASAP7_75t_L g1011 ( 
.A1(n_945),
.A2(n_316),
.A3(n_317),
.B1(n_6),
.B2(n_7),
.C(n_8),
.Y(n_1011)
);

AND2x4_ASAP7_75t_L g1012 ( 
.A(n_941),
.B(n_4),
.Y(n_1012)
);

O2A1O1Ixp33_ASAP7_75t_L g1013 ( 
.A1(n_945),
.A2(n_5),
.B(n_7),
.C(n_8),
.Y(n_1013)
);

INVx1_ASAP7_75t_L g1014 ( 
.A(n_917),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_910),
.Y(n_1015)
);

INVx3_ASAP7_75t_L g1016 ( 
.A(n_953),
.Y(n_1016)
);

BUFx3_ASAP7_75t_L g1017 ( 
.A(n_954),
.Y(n_1017)
);

AOI21xp5_ASAP7_75t_L g1018 ( 
.A1(n_929),
.A2(n_928),
.B(n_947),
.Y(n_1018)
);

NOR2x1_ASAP7_75t_L g1019 ( 
.A(n_912),
.B(n_509),
.Y(n_1019)
);

INVx1_ASAP7_75t_L g1020 ( 
.A(n_920),
.Y(n_1020)
);

AOI21xp5_ASAP7_75t_L g1021 ( 
.A1(n_929),
.A2(n_502),
.B(n_492),
.Y(n_1021)
);

NAND2xp5_ASAP7_75t_SL g1022 ( 
.A(n_946),
.B(n_502),
.Y(n_1022)
);

AOI21xp5_ASAP7_75t_L g1023 ( 
.A1(n_924),
.A2(n_492),
.B(n_317),
.Y(n_1023)
);

HB1xp67_ASAP7_75t_L g1024 ( 
.A(n_942),
.Y(n_1024)
);

NAND2xp5_ASAP7_75t_L g1025 ( 
.A(n_943),
.B(n_10),
.Y(n_1025)
);

OAI21xp5_ASAP7_75t_L g1026 ( 
.A1(n_948),
.A2(n_533),
.B(n_492),
.Y(n_1026)
);

INVx2_ASAP7_75t_L g1027 ( 
.A(n_997),
.Y(n_1027)
);

INVx2_ASAP7_75t_L g1028 ( 
.A(n_978),
.Y(n_1028)
);

AND3x1_ASAP7_75t_SL g1029 ( 
.A(n_999),
.B(n_12),
.C(n_13),
.Y(n_1029)
);

INVx6_ASAP7_75t_L g1030 ( 
.A(n_968),
.Y(n_1030)
);

INVx2_ASAP7_75t_L g1031 ( 
.A(n_1014),
.Y(n_1031)
);

INVx5_ASAP7_75t_L g1032 ( 
.A(n_968),
.Y(n_1032)
);

BUFx10_ASAP7_75t_L g1033 ( 
.A(n_1012),
.Y(n_1033)
);

INVx3_ASAP7_75t_L g1034 ( 
.A(n_968),
.Y(n_1034)
);

BUFx3_ASAP7_75t_L g1035 ( 
.A(n_1005),
.Y(n_1035)
);

HB1xp67_ASAP7_75t_L g1036 ( 
.A(n_1024),
.Y(n_1036)
);

AND2x6_ASAP7_75t_SL g1037 ( 
.A(n_992),
.B(n_12),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_SL g1038 ( 
.A(n_977),
.B(n_981),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_1020),
.Y(n_1039)
);

INVx1_ASAP7_75t_L g1040 ( 
.A(n_1015),
.Y(n_1040)
);

NAND2xp5_ASAP7_75t_L g1041 ( 
.A(n_966),
.B(n_13),
.Y(n_1041)
);

OAI22xp33_ASAP7_75t_L g1042 ( 
.A1(n_984),
.A2(n_539),
.B1(n_524),
.B2(n_525),
.Y(n_1042)
);

NAND2xp5_ASAP7_75t_L g1043 ( 
.A(n_971),
.B(n_14),
.Y(n_1043)
);

BUFx6f_ASAP7_75t_L g1044 ( 
.A(n_1009),
.Y(n_1044)
);

INVx5_ASAP7_75t_L g1045 ( 
.A(n_1032),
.Y(n_1045)
);

BUFx6f_ASAP7_75t_L g1046 ( 
.A(n_1044),
.Y(n_1046)
);

NAND2xp33_ASAP7_75t_L g1047 ( 
.A(n_1038),
.B(n_970),
.Y(n_1047)
);

NAND2x1_ASAP7_75t_L g1048 ( 
.A(n_1030),
.B(n_973),
.Y(n_1048)
);

A2O1A1Ixp33_ASAP7_75t_L g1049 ( 
.A1(n_1041),
.A2(n_1013),
.B(n_993),
.C(n_1003),
.Y(n_1049)
);

NAND2xp5_ASAP7_75t_SL g1050 ( 
.A(n_1032),
.B(n_983),
.Y(n_1050)
);

AND2x2_ASAP7_75t_L g1051 ( 
.A(n_1035),
.B(n_973),
.Y(n_1051)
);

NAND2xp5_ASAP7_75t_SL g1052 ( 
.A(n_1032),
.B(n_987),
.Y(n_1052)
);

NOR2xp33_ASAP7_75t_L g1053 ( 
.A(n_1035),
.B(n_969),
.Y(n_1053)
);

AND2x2_ASAP7_75t_L g1054 ( 
.A(n_1044),
.B(n_973),
.Y(n_1054)
);

OAI21xp5_ASAP7_75t_L g1055 ( 
.A1(n_1043),
.A2(n_996),
.B(n_985),
.Y(n_1055)
);

INVx1_ASAP7_75t_SL g1056 ( 
.A(n_1030),
.Y(n_1056)
);

INVx2_ASAP7_75t_L g1057 ( 
.A(n_1030),
.Y(n_1057)
);

NAND2xp5_ASAP7_75t_L g1058 ( 
.A(n_1036),
.B(n_986),
.Y(n_1058)
);

AOI22xp5_ASAP7_75t_L g1059 ( 
.A1(n_1044),
.A2(n_965),
.B1(n_967),
.B2(n_972),
.Y(n_1059)
);

NOR3xp33_ASAP7_75t_L g1060 ( 
.A(n_1034),
.B(n_1011),
.C(n_1025),
.Y(n_1060)
);

BUFx2_ASAP7_75t_SL g1061 ( 
.A(n_1032),
.Y(n_1061)
);

AOI21xp5_ASAP7_75t_L g1062 ( 
.A1(n_1042),
.A2(n_974),
.B(n_989),
.Y(n_1062)
);

INVx3_ASAP7_75t_L g1063 ( 
.A(n_1032),
.Y(n_1063)
);

AOI21xp5_ASAP7_75t_L g1064 ( 
.A1(n_1044),
.A2(n_1010),
.B(n_1018),
.Y(n_1064)
);

OAI22xp5_ASAP7_75t_L g1065 ( 
.A1(n_1044),
.A2(n_1030),
.B1(n_976),
.B2(n_1034),
.Y(n_1065)
);

INVx1_ASAP7_75t_SL g1066 ( 
.A(n_1034),
.Y(n_1066)
);

AOI21xp5_ASAP7_75t_L g1067 ( 
.A1(n_1040),
.A2(n_1007),
.B(n_990),
.Y(n_1067)
);

INVx2_ASAP7_75t_L g1068 ( 
.A(n_1033),
.Y(n_1068)
);

INVx2_ASAP7_75t_L g1069 ( 
.A(n_1033),
.Y(n_1069)
);

BUFx2_ASAP7_75t_R g1070 ( 
.A(n_1050),
.Y(n_1070)
);

INVx2_ASAP7_75t_SL g1071 ( 
.A(n_1045),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_L g1072 ( 
.A(n_1060),
.B(n_1037),
.Y(n_1072)
);

INVxp67_ASAP7_75t_SL g1073 ( 
.A(n_1047),
.Y(n_1073)
);

INVx1_ASAP7_75t_L g1074 ( 
.A(n_1066),
.Y(n_1074)
);

BUFx3_ASAP7_75t_L g1075 ( 
.A(n_1046),
.Y(n_1075)
);

OAI21x1_ASAP7_75t_L g1076 ( 
.A1(n_1048),
.A2(n_1027),
.B(n_1028),
.Y(n_1076)
);

BUFx6f_ASAP7_75t_L g1077 ( 
.A(n_1075),
.Y(n_1077)
);

AOI21xp5_ASAP7_75t_L g1078 ( 
.A1(n_1072),
.A2(n_1055),
.B(n_1073),
.Y(n_1078)
);

INVx2_ASAP7_75t_L g1079 ( 
.A(n_1071),
.Y(n_1079)
);

INVx1_ASAP7_75t_SL g1080 ( 
.A(n_1077),
.Y(n_1080)
);

BUFx2_ASAP7_75t_L g1081 ( 
.A(n_1077),
.Y(n_1081)
);

INVx1_ASAP7_75t_L g1082 ( 
.A(n_1079),
.Y(n_1082)
);

OAI21x1_ASAP7_75t_SL g1083 ( 
.A1(n_1082),
.A2(n_1078),
.B(n_1055),
.Y(n_1083)
);

BUFx6f_ASAP7_75t_L g1084 ( 
.A(n_1081),
.Y(n_1084)
);

INVx6_ASAP7_75t_L g1085 ( 
.A(n_1084),
.Y(n_1085)
);

INVx6_ASAP7_75t_L g1086 ( 
.A(n_1084),
.Y(n_1086)
);

OAI22xp5_ASAP7_75t_L g1087 ( 
.A1(n_1085),
.A2(n_1070),
.B1(n_1059),
.B2(n_1058),
.Y(n_1087)
);

BUFx6f_ASAP7_75t_L g1088 ( 
.A(n_1086),
.Y(n_1088)
);

INVx1_ASAP7_75t_L g1089 ( 
.A(n_1088),
.Y(n_1089)
);

AND2x2_ASAP7_75t_L g1090 ( 
.A(n_1087),
.B(n_1081),
.Y(n_1090)
);

AOI22xp33_ASAP7_75t_L g1091 ( 
.A1(n_1090),
.A2(n_1083),
.B1(n_1080),
.B2(n_1074),
.Y(n_1091)
);

OAI22xp5_ASAP7_75t_L g1092 ( 
.A1(n_1089),
.A2(n_1068),
.B1(n_1069),
.B2(n_1056),
.Y(n_1092)
);

INVx2_ASAP7_75t_L g1093 ( 
.A(n_1092),
.Y(n_1093)
);

INVx4_ASAP7_75t_L g1094 ( 
.A(n_1091),
.Y(n_1094)
);

AND2x2_ASAP7_75t_L g1095 ( 
.A(n_1093),
.B(n_1090),
.Y(n_1095)
);

BUFx6f_ASAP7_75t_L g1096 ( 
.A(n_1094),
.Y(n_1096)
);

OAI21x1_ASAP7_75t_L g1097 ( 
.A1(n_1093),
.A2(n_1074),
.B(n_1076),
.Y(n_1097)
);

AOI22xp33_ASAP7_75t_L g1098 ( 
.A1(n_1096),
.A2(n_1071),
.B1(n_1075),
.B2(n_1056),
.Y(n_1098)
);

AO31x2_ASAP7_75t_L g1099 ( 
.A1(n_1095),
.A2(n_1057),
.A3(n_1053),
.B(n_1065),
.Y(n_1099)
);

AND2x2_ASAP7_75t_L g1100 ( 
.A(n_1096),
.B(n_1066),
.Y(n_1100)
);

OR2x2_ASAP7_75t_L g1101 ( 
.A(n_1099),
.B(n_1097),
.Y(n_1101)
);

HB1xp67_ASAP7_75t_L g1102 ( 
.A(n_1100),
.Y(n_1102)
);

AND2x2_ASAP7_75t_L g1103 ( 
.A(n_1102),
.B(n_1098),
.Y(n_1103)
);

BUFx6f_ASAP7_75t_L g1104 ( 
.A(n_1101),
.Y(n_1104)
);

OA21x2_ASAP7_75t_L g1105 ( 
.A1(n_1103),
.A2(n_1096),
.B(n_1104),
.Y(n_1105)
);

OAI21xp5_ASAP7_75t_L g1106 ( 
.A1(n_1104),
.A2(n_1076),
.B(n_1063),
.Y(n_1106)
);

INVx2_ASAP7_75t_L g1107 ( 
.A(n_1105),
.Y(n_1107)
);

OAI21xp33_ASAP7_75t_L g1108 ( 
.A1(n_1106),
.A2(n_1063),
.B(n_1052),
.Y(n_1108)
);

INVx2_ASAP7_75t_L g1109 ( 
.A(n_1107),
.Y(n_1109)
);

NOR3xp33_ASAP7_75t_L g1110 ( 
.A(n_1108),
.B(n_1049),
.C(n_1064),
.Y(n_1110)
);

NAND2xp5_ASAP7_75t_L g1111 ( 
.A(n_1110),
.B(n_1045),
.Y(n_1111)
);

INVx2_ASAP7_75t_L g1112 ( 
.A(n_1109),
.Y(n_1112)
);

INVx1_ASAP7_75t_L g1113 ( 
.A(n_1111),
.Y(n_1113)
);

INVx1_ASAP7_75t_L g1114 ( 
.A(n_1112),
.Y(n_1114)
);

INVx1_ASAP7_75t_SL g1115 ( 
.A(n_1111),
.Y(n_1115)
);

AOI31xp33_ASAP7_75t_L g1116 ( 
.A1(n_1114),
.A2(n_1051),
.A3(n_1054),
.B(n_1067),
.Y(n_1116)
);

AND2x2_ASAP7_75t_L g1117 ( 
.A(n_1115),
.B(n_1061),
.Y(n_1117)
);

OA21x2_ASAP7_75t_L g1118 ( 
.A1(n_1113),
.A2(n_1045),
.B(n_1062),
.Y(n_1118)
);

NAND2xp5_ASAP7_75t_L g1119 ( 
.A(n_1117),
.B(n_1116),
.Y(n_1119)
);

OR2x2_ASAP7_75t_L g1120 ( 
.A(n_1118),
.B(n_1045),
.Y(n_1120)
);

INVx1_ASAP7_75t_L g1121 ( 
.A(n_1120),
.Y(n_1121)
);

AND2x2_ASAP7_75t_L g1122 ( 
.A(n_1119),
.B(n_1046),
.Y(n_1122)
);

NAND2xp5_ASAP7_75t_L g1123 ( 
.A(n_1122),
.B(n_1046),
.Y(n_1123)
);

AND2x2_ASAP7_75t_L g1124 ( 
.A(n_1121),
.B(n_1027),
.Y(n_1124)
);

INVx1_ASAP7_75t_L g1125 ( 
.A(n_1123),
.Y(n_1125)
);

INVx1_ASAP7_75t_L g1126 ( 
.A(n_1124),
.Y(n_1126)
);

INVx2_ASAP7_75t_L g1127 ( 
.A(n_1126),
.Y(n_1127)
);

NAND2xp5_ASAP7_75t_L g1128 ( 
.A(n_1125),
.B(n_14),
.Y(n_1128)
);

AOI22xp5_ASAP7_75t_L g1129 ( 
.A1(n_1127),
.A2(n_1040),
.B1(n_1039),
.B2(n_1028),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_1128),
.Y(n_1130)
);

INVx1_ASAP7_75t_L g1131 ( 
.A(n_1130),
.Y(n_1131)
);

AND2x2_ASAP7_75t_L g1132 ( 
.A(n_1129),
.B(n_1031),
.Y(n_1132)
);

OAI322xp33_ASAP7_75t_L g1133 ( 
.A1(n_1130),
.A2(n_15),
.A3(n_17),
.B1(n_18),
.B2(n_19),
.C1(n_20),
.C2(n_21),
.Y(n_1133)
);

OAI22xp5_ASAP7_75t_L g1134 ( 
.A1(n_1131),
.A2(n_1039),
.B1(n_1031),
.B2(n_20),
.Y(n_1134)
);

INVx1_ASAP7_75t_L g1135 ( 
.A(n_1132),
.Y(n_1135)
);

AOI22xp5_ASAP7_75t_L g1136 ( 
.A1(n_1133),
.A2(n_1029),
.B1(n_1033),
.B2(n_1012),
.Y(n_1136)
);

INVx1_ASAP7_75t_L g1137 ( 
.A(n_1135),
.Y(n_1137)
);

INVx1_ASAP7_75t_L g1138 ( 
.A(n_1134),
.Y(n_1138)
);

INVx1_ASAP7_75t_L g1139 ( 
.A(n_1137),
.Y(n_1139)
);

NAND2xp5_ASAP7_75t_L g1140 ( 
.A(n_1138),
.B(n_1136),
.Y(n_1140)
);

NAND3xp33_ASAP7_75t_L g1141 ( 
.A(n_1139),
.B(n_326),
.C(n_325),
.Y(n_1141)
);

OAI221xp5_ASAP7_75t_L g1142 ( 
.A1(n_1140),
.A2(n_15),
.B1(n_18),
.B2(n_21),
.C(n_22),
.Y(n_1142)
);

NOR2xp33_ASAP7_75t_L g1143 ( 
.A(n_1141),
.B(n_22),
.Y(n_1143)
);

AOI21xp5_ASAP7_75t_L g1144 ( 
.A1(n_1142),
.A2(n_326),
.B(n_325),
.Y(n_1144)
);

NAND3xp33_ASAP7_75t_L g1145 ( 
.A(n_1144),
.B(n_324),
.C(n_23),
.Y(n_1145)
);

NAND2xp5_ASAP7_75t_L g1146 ( 
.A(n_1143),
.B(n_24),
.Y(n_1146)
);

AOI211xp5_ASAP7_75t_L g1147 ( 
.A1(n_1145),
.A2(n_25),
.B(n_26),
.C(n_27),
.Y(n_1147)
);

INVxp67_ASAP7_75t_SL g1148 ( 
.A(n_1146),
.Y(n_1148)
);

AOI31xp33_ASAP7_75t_L g1149 ( 
.A1(n_1148),
.A2(n_25),
.A3(n_26),
.B(n_28),
.Y(n_1149)
);

OAI321xp33_ASAP7_75t_L g1150 ( 
.A1(n_1147),
.A2(n_29),
.A3(n_30),
.B1(n_31),
.B2(n_32),
.C(n_33),
.Y(n_1150)
);

AOI221xp5_ASAP7_75t_L g1151 ( 
.A1(n_1148),
.A2(n_324),
.B1(n_30),
.B2(n_31),
.C(n_33),
.Y(n_1151)
);

NOR2x1_ASAP7_75t_L g1152 ( 
.A(n_1150),
.B(n_29),
.Y(n_1152)
);

OAI22xp33_ASAP7_75t_L g1153 ( 
.A1(n_1149),
.A2(n_34),
.B1(n_35),
.B2(n_36),
.Y(n_1153)
);

AOI221xp5_ASAP7_75t_L g1154 ( 
.A1(n_1151),
.A2(n_34),
.B1(n_35),
.B2(n_36),
.C(n_1037),
.Y(n_1154)
);

NOR4xp25_ASAP7_75t_L g1155 ( 
.A(n_1152),
.B(n_37),
.C(n_39),
.D(n_40),
.Y(n_1155)
);

OAI221xp5_ASAP7_75t_L g1156 ( 
.A1(n_1153),
.A2(n_41),
.B1(n_43),
.B2(n_44),
.C(n_45),
.Y(n_1156)
);

INVx1_ASAP7_75t_L g1157 ( 
.A(n_1155),
.Y(n_1157)
);

AND2x2_ASAP7_75t_SL g1158 ( 
.A(n_1156),
.B(n_1154),
.Y(n_1158)
);

A2O1A1Ixp33_ASAP7_75t_SL g1159 ( 
.A1(n_1157),
.A2(n_46),
.B(n_48),
.C(n_49),
.Y(n_1159)
);

OAI211xp5_ASAP7_75t_SL g1160 ( 
.A1(n_1158),
.A2(n_50),
.B(n_51),
.C(n_52),
.Y(n_1160)
);

INVx1_ASAP7_75t_L g1161 ( 
.A(n_1160),
.Y(n_1161)
);

INVxp33_ASAP7_75t_L g1162 ( 
.A(n_1159),
.Y(n_1162)
);

NOR2x1_ASAP7_75t_L g1163 ( 
.A(n_1161),
.B(n_55),
.Y(n_1163)
);

NAND2xp5_ASAP7_75t_L g1164 ( 
.A(n_1162),
.B(n_59),
.Y(n_1164)
);

AND2x2_ASAP7_75t_L g1165 ( 
.A(n_1163),
.B(n_60),
.Y(n_1165)
);

INVx1_ASAP7_75t_L g1166 ( 
.A(n_1164),
.Y(n_1166)
);

NAND4xp25_ASAP7_75t_SL g1167 ( 
.A(n_1166),
.B(n_63),
.C(n_64),
.D(n_66),
.Y(n_1167)
);

OR5x1_ASAP7_75t_L g1168 ( 
.A(n_1165),
.B(n_68),
.C(n_70),
.D(n_71),
.E(n_72),
.Y(n_1168)
);

NOR2x1_ASAP7_75t_L g1169 ( 
.A(n_1166),
.B(n_74),
.Y(n_1169)
);

OAI22xp5_ASAP7_75t_L g1170 ( 
.A1(n_1168),
.A2(n_75),
.B1(n_76),
.B2(n_77),
.Y(n_1170)
);

HB1xp67_ASAP7_75t_L g1171 ( 
.A(n_1169),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_1167),
.Y(n_1172)
);

AOI32xp33_ASAP7_75t_L g1173 ( 
.A1(n_1172),
.A2(n_78),
.A3(n_79),
.B1(n_80),
.B2(n_81),
.Y(n_1173)
);

AOI322xp5_ASAP7_75t_L g1174 ( 
.A1(n_1171),
.A2(n_82),
.A3(n_83),
.B1(n_84),
.B2(n_86),
.C1(n_89),
.C2(n_90),
.Y(n_1174)
);

OAI22xp5_ASAP7_75t_L g1175 ( 
.A1(n_1173),
.A2(n_1170),
.B1(n_93),
.B2(n_94),
.Y(n_1175)
);

HB1xp67_ASAP7_75t_L g1176 ( 
.A(n_1174),
.Y(n_1176)
);

OAI22xp5_ASAP7_75t_L g1177 ( 
.A1(n_1176),
.A2(n_91),
.B1(n_95),
.B2(n_97),
.Y(n_1177)
);

OAI22x1_ASAP7_75t_L g1178 ( 
.A1(n_1175),
.A2(n_98),
.B1(n_99),
.B2(n_100),
.Y(n_1178)
);

INVx1_ASAP7_75t_L g1179 ( 
.A(n_1178),
.Y(n_1179)
);

INVx2_ASAP7_75t_L g1180 ( 
.A(n_1177),
.Y(n_1180)
);

NAND2xp5_ASAP7_75t_L g1181 ( 
.A(n_1180),
.B(n_1179),
.Y(n_1181)
);

OAI22xp5_ASAP7_75t_SL g1182 ( 
.A1(n_1180),
.A2(n_102),
.B1(n_103),
.B2(n_104),
.Y(n_1182)
);

AND3x4_ASAP7_75t_L g1183 ( 
.A(n_1181),
.B(n_105),
.C(n_107),
.Y(n_1183)
);

INVx1_ASAP7_75t_SL g1184 ( 
.A(n_1182),
.Y(n_1184)
);

NAND2xp5_ASAP7_75t_L g1185 ( 
.A(n_1184),
.B(n_108),
.Y(n_1185)
);

AOI22xp5_ASAP7_75t_L g1186 ( 
.A1(n_1183),
.A2(n_533),
.B1(n_1006),
.B2(n_980),
.Y(n_1186)
);

AND2x2_ASAP7_75t_L g1187 ( 
.A(n_1184),
.B(n_109),
.Y(n_1187)
);

OAI22xp5_ASAP7_75t_L g1188 ( 
.A1(n_1184),
.A2(n_1006),
.B1(n_980),
.B2(n_1017),
.Y(n_1188)
);

AOI22xp5_ASAP7_75t_L g1189 ( 
.A1(n_1186),
.A2(n_533),
.B1(n_1006),
.B2(n_980),
.Y(n_1189)
);

OAI21xp5_ASAP7_75t_L g1190 ( 
.A1(n_1185),
.A2(n_1187),
.B(n_1188),
.Y(n_1190)
);

OAI22xp5_ASAP7_75t_L g1191 ( 
.A1(n_1186),
.A2(n_111),
.B1(n_112),
.B2(n_113),
.Y(n_1191)
);

NAND2xp5_ASAP7_75t_L g1192 ( 
.A(n_1186),
.B(n_114),
.Y(n_1192)
);

CKINVDCx20_ASAP7_75t_R g1193 ( 
.A(n_1190),
.Y(n_1193)
);

HB1xp67_ASAP7_75t_L g1194 ( 
.A(n_1192),
.Y(n_1194)
);

AND2x4_ASAP7_75t_L g1195 ( 
.A(n_1189),
.B(n_117),
.Y(n_1195)
);

HB1xp67_ASAP7_75t_L g1196 ( 
.A(n_1193),
.Y(n_1196)
);

OAI22xp5_ASAP7_75t_L g1197 ( 
.A1(n_1194),
.A2(n_1191),
.B1(n_120),
.B2(n_121),
.Y(n_1197)
);

AOI22xp33_ASAP7_75t_L g1198 ( 
.A1(n_1195),
.A2(n_533),
.B1(n_122),
.B2(n_124),
.Y(n_1198)
);

AOI22xp5_ASAP7_75t_L g1199 ( 
.A1(n_1193),
.A2(n_533),
.B1(n_125),
.B2(n_126),
.Y(n_1199)
);

AOI21xp5_ASAP7_75t_L g1200 ( 
.A1(n_1193),
.A2(n_119),
.B(n_128),
.Y(n_1200)
);

OAI21x1_ASAP7_75t_L g1201 ( 
.A1(n_1193),
.A2(n_130),
.B(n_131),
.Y(n_1201)
);

OAI22xp33_ASAP7_75t_L g1202 ( 
.A1(n_1193),
.A2(n_133),
.B1(n_135),
.B2(n_137),
.Y(n_1202)
);

AOI21xp33_ASAP7_75t_L g1203 ( 
.A1(n_1193),
.A2(n_138),
.B(n_139),
.Y(n_1203)
);

OAI22xp5_ASAP7_75t_L g1204 ( 
.A1(n_1193),
.A2(n_140),
.B1(n_143),
.B2(n_145),
.Y(n_1204)
);

AO21x1_ASAP7_75t_SL g1205 ( 
.A1(n_1193),
.A2(n_146),
.B(n_148),
.Y(n_1205)
);

XNOR2xp5_ASAP7_75t_L g1206 ( 
.A(n_1193),
.B(n_150),
.Y(n_1206)
);

AOI221x1_ASAP7_75t_L g1207 ( 
.A1(n_1193),
.A2(n_152),
.B1(n_153),
.B2(n_154),
.C(n_155),
.Y(n_1207)
);

BUFx2_ASAP7_75t_SL g1208 ( 
.A(n_1196),
.Y(n_1208)
);

AOI21xp5_ASAP7_75t_L g1209 ( 
.A1(n_1197),
.A2(n_156),
.B(n_158),
.Y(n_1209)
);

OR3x1_ASAP7_75t_L g1210 ( 
.A(n_1201),
.B(n_161),
.C(n_162),
.Y(n_1210)
);

O2A1O1Ixp33_ASAP7_75t_L g1211 ( 
.A1(n_1198),
.A2(n_163),
.B(n_164),
.C(n_165),
.Y(n_1211)
);

AOI211xp5_ASAP7_75t_L g1212 ( 
.A1(n_1200),
.A2(n_167),
.B(n_168),
.C(n_169),
.Y(n_1212)
);

INVx1_ASAP7_75t_SL g1213 ( 
.A(n_1206),
.Y(n_1213)
);

OAI322xp33_ASAP7_75t_L g1214 ( 
.A1(n_1202),
.A2(n_170),
.A3(n_171),
.B1(n_172),
.B2(n_173),
.C1(n_174),
.C2(n_175),
.Y(n_1214)
);

AOI211xp5_ASAP7_75t_L g1215 ( 
.A1(n_1205),
.A2(n_176),
.B(n_178),
.C(n_1023),
.Y(n_1215)
);

AOI22xp5_ASAP7_75t_L g1216 ( 
.A1(n_1204),
.A2(n_533),
.B1(n_420),
.B2(n_1016),
.Y(n_1216)
);

AOI22xp5_ASAP7_75t_L g1217 ( 
.A1(n_1208),
.A2(n_1213),
.B1(n_1210),
.B2(n_1209),
.Y(n_1217)
);

OR2x6_ASAP7_75t_L g1218 ( 
.A(n_1211),
.B(n_1207),
.Y(n_1218)
);

AOI21xp33_ASAP7_75t_L g1219 ( 
.A1(n_1216),
.A2(n_1203),
.B(n_1199),
.Y(n_1219)
);

OAI22xp5_ASAP7_75t_L g1220 ( 
.A1(n_1212),
.A2(n_1002),
.B1(n_539),
.B2(n_530),
.Y(n_1220)
);

AOI22xp5_ASAP7_75t_L g1221 ( 
.A1(n_1215),
.A2(n_420),
.B1(n_524),
.B2(n_525),
.Y(n_1221)
);

AOI21xp5_ASAP7_75t_L g1222 ( 
.A1(n_1214),
.A2(n_532),
.B(n_522),
.Y(n_1222)
);

AOI21xp5_ASAP7_75t_L g1223 ( 
.A1(n_1208),
.A2(n_532),
.B(n_522),
.Y(n_1223)
);

XOR2xp5_ASAP7_75t_L g1224 ( 
.A(n_1217),
.B(n_975),
.Y(n_1224)
);

NAND2xp5_ASAP7_75t_L g1225 ( 
.A(n_1218),
.B(n_420),
.Y(n_1225)
);

NAND2xp5_ASAP7_75t_L g1226 ( 
.A(n_1219),
.B(n_420),
.Y(n_1226)
);

OAI21xp5_ASAP7_75t_L g1227 ( 
.A1(n_1225),
.A2(n_1222),
.B(n_1221),
.Y(n_1227)
);

OAI21xp5_ASAP7_75t_L g1228 ( 
.A1(n_1227),
.A2(n_1220),
.B(n_1223),
.Y(n_1228)
);

INVx1_ASAP7_75t_L g1229 ( 
.A(n_1228),
.Y(n_1229)
);

INVx1_ASAP7_75t_L g1230 ( 
.A(n_1229),
.Y(n_1230)
);

OA21x2_ASAP7_75t_L g1231 ( 
.A1(n_1230),
.A2(n_1226),
.B(n_1224),
.Y(n_1231)
);

OAI221xp5_ASAP7_75t_R g1232 ( 
.A1(n_1231),
.A2(n_991),
.B1(n_994),
.B2(n_1008),
.C(n_1019),
.Y(n_1232)
);

AOI22xp5_ASAP7_75t_L g1233 ( 
.A1(n_1232),
.A2(n_964),
.B1(n_979),
.B2(n_982),
.Y(n_1233)
);

AOI22xp5_ASAP7_75t_L g1234 ( 
.A1(n_1233),
.A2(n_988),
.B1(n_995),
.B2(n_1001),
.Y(n_1234)
);

AOI211xp5_ASAP7_75t_L g1235 ( 
.A1(n_1234),
.A2(n_998),
.B(n_1004),
.C(n_1021),
.Y(n_1235)
);

AOI211xp5_ASAP7_75t_L g1236 ( 
.A1(n_1235),
.A2(n_1022),
.B(n_1026),
.C(n_1000),
.Y(n_1236)
);


endmodule