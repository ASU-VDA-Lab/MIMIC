module real_jpeg_6004_n_20 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_19, n_16, n_15, n_13, n_20);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_19;
input n_16;
input n_15;
input n_13;

output n_20;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_456;
wire n_259;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_233;
wire n_73;
wire n_532;
wire n_516;
wire n_348;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_525;
wire n_288;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_469;
wire n_378;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_533;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_215;
wire n_176;
wire n_166;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_531;
wire n_112;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_537;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_534;
wire n_256;
wire n_520;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_343;
wire n_292;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_444;
wire n_178;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

CKINVDCx16_ASAP7_75t_R g171 ( 
.A(n_0),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_0),
.B(n_176),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_0),
.B(n_206),
.Y(n_205)
);

AND2x2_ASAP7_75t_SL g233 ( 
.A(n_0),
.B(n_234),
.Y(n_233)
);

AND2x2_ASAP7_75t_L g248 ( 
.A(n_0),
.B(n_249),
.Y(n_248)
);

AND2x2_ASAP7_75t_L g307 ( 
.A(n_0),
.B(n_308),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_0),
.B(n_267),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_SL g443 ( 
.A(n_0),
.B(n_444),
.Y(n_443)
);

INVx8_ASAP7_75t_L g169 ( 
.A(n_1),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g276 ( 
.A(n_1),
.Y(n_276)
);

INVx2_ASAP7_75t_L g326 ( 
.A(n_1),
.Y(n_326)
);

BUFx6f_ASAP7_75t_L g343 ( 
.A(n_1),
.Y(n_343)
);

BUFx6f_ASAP7_75t_L g403 ( 
.A(n_1),
.Y(n_403)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_2),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_2),
.Y(n_65)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_2),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g176 ( 
.A(n_2),
.Y(n_176)
);

INVx6_ASAP7_75t_L g472 ( 
.A(n_2),
.Y(n_472)
);

BUFx6f_ASAP7_75t_L g495 ( 
.A(n_2),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_3),
.B(n_217),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_3),
.B(n_229),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_3),
.B(n_258),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_3),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_3),
.B(n_147),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_3),
.B(n_350),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_3),
.B(n_140),
.Y(n_365)
);

CKINVDCx14_ASAP7_75t_R g92 ( 
.A(n_4),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g178 ( 
.A(n_4),
.B(n_179),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_4),
.B(n_211),
.Y(n_210)
);

AND2x2_ASAP7_75t_SL g236 ( 
.A(n_4),
.B(n_237),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_4),
.B(n_415),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_4),
.B(n_458),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_5),
.B(n_223),
.Y(n_222)
);

AND2x2_ASAP7_75t_L g245 ( 
.A(n_5),
.B(n_246),
.Y(n_245)
);

AND2x2_ASAP7_75t_L g260 ( 
.A(n_5),
.B(n_261),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_5),
.B(n_325),
.Y(n_324)
);

AND2x2_ASAP7_75t_L g338 ( 
.A(n_5),
.B(n_339),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_5),
.B(n_304),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_5),
.B(n_421),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_5),
.B(n_471),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_6),
.B(n_63),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_6),
.B(n_82),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_6),
.B(n_36),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_6),
.B(n_88),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_6),
.B(n_142),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_6),
.B(n_211),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_6),
.B(n_406),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_SL g442 ( 
.A(n_6),
.B(n_331),
.Y(n_442)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_7),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_7),
.Y(n_55)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_7),
.Y(n_106)
);

BUFx5_ASAP7_75t_L g173 ( 
.A(n_7),
.Y(n_173)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_9),
.B(n_34),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_9),
.B(n_49),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_9),
.B(n_86),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_9),
.B(n_98),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_9),
.B(n_132),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_9),
.B(n_145),
.Y(n_144)
);

AND2x2_ASAP7_75t_SL g402 ( 
.A(n_9),
.B(n_403),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_9),
.B(n_467),
.Y(n_466)
);

BUFx3_ASAP7_75t_L g110 ( 
.A(n_10),
.Y(n_110)
);

INVx3_ASAP7_75t_L g148 ( 
.A(n_10),
.Y(n_148)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_10),
.Y(n_239)
);

BUFx5_ASAP7_75t_L g331 ( 
.A(n_10),
.Y(n_331)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_11),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g20 ( 
.A1(n_12),
.A2(n_21),
.B1(n_24),
.B2(n_25),
.Y(n_20)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_13),
.Y(n_159)
);

BUFx3_ASAP7_75t_L g272 ( 
.A(n_13),
.Y(n_272)
);

BUFx6f_ASAP7_75t_L g323 ( 
.A(n_13),
.Y(n_323)
);

AND2x2_ASAP7_75t_SL g38 ( 
.A(n_14),
.B(n_39),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_14),
.B(n_43),
.Y(n_42)
);

INVx1_ASAP7_75t_SL g53 ( 
.A(n_14),
.Y(n_53)
);

AND2x2_ASAP7_75t_SL g72 ( 
.A(n_14),
.B(n_73),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_14),
.B(n_109),
.Y(n_108)
);

AND2x2_ASAP7_75t_SL g167 ( 
.A(n_14),
.B(n_168),
.Y(n_167)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_15),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_16),
.B(n_69),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_16),
.B(n_105),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_16),
.B(n_138),
.Y(n_137)
);

AND2x2_ASAP7_75t_L g150 ( 
.A(n_16),
.B(n_151),
.Y(n_150)
);

AND2x2_ASAP7_75t_L g273 ( 
.A(n_16),
.B(n_274),
.Y(n_273)
);

AND2x2_ASAP7_75t_L g286 ( 
.A(n_16),
.B(n_287),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_16),
.B(n_331),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_16),
.B(n_453),
.Y(n_452)
);

AND2x2_ASAP7_75t_L g251 ( 
.A(n_17),
.B(n_252),
.Y(n_251)
);

AND2x2_ASAP7_75t_L g279 ( 
.A(n_17),
.B(n_280),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_SL g301 ( 
.A(n_17),
.B(n_302),
.Y(n_301)
);

AND2x2_ASAP7_75t_L g311 ( 
.A(n_17),
.B(n_312),
.Y(n_311)
);

AND2x2_ASAP7_75t_L g342 ( 
.A(n_17),
.B(n_343),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_17),
.B(n_258),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_17),
.B(n_456),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_17),
.B(n_495),
.Y(n_494)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_18),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_19),
.B(n_215),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_19),
.B(n_267),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_19),
.B(n_283),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_19),
.B(n_322),
.Y(n_321)
);

AND2x2_ASAP7_75t_L g330 ( 
.A(n_19),
.B(n_331),
.Y(n_330)
);

CKINVDCx14_ASAP7_75t_R g361 ( 
.A(n_19),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_19),
.B(n_231),
.Y(n_399)
);

INVx3_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_22),
.Y(n_24)
);

INVx13_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

XNOR2xp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_121),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_120),
.Y(n_26)
);

INVxp67_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_77),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_29),
.B(n_77),
.Y(n_120)
);

XNOR2xp5_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_57),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_L g30 ( 
.A1(n_31),
.A2(n_32),
.B1(n_46),
.B2(n_47),
.Y(n_30)
);

CKINVDCx14_ASAP7_75t_R g31 ( 
.A(n_32),
.Y(n_31)
);

MAJIxp5_ASAP7_75t_L g32 ( 
.A(n_33),
.B(n_38),
.C(n_42),
.Y(n_32)
);

XOR2xp5_ASAP7_75t_L g59 ( 
.A(n_33),
.B(n_60),
.Y(n_59)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx5_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx3_ASAP7_75t_L g456 ( 
.A(n_37),
.Y(n_456)
);

OAI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_38),
.A2(n_42),
.B1(n_56),
.B2(n_61),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_38),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_38),
.A2(n_61),
.B1(n_72),
.B2(n_111),
.Y(n_115)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_41),
.Y(n_90)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_41),
.Y(n_140)
);

INVx3_ASAP7_75t_L g247 ( 
.A(n_41),
.Y(n_247)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_41),
.Y(n_460)
);

OAI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_42),
.A2(n_51),
.B1(n_52),
.B2(n_56),
.Y(n_50)
);

CKINVDCx16_ASAP7_75t_R g56 ( 
.A(n_42),
.Y(n_56)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_44),
.Y(n_84)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_44),
.Y(n_101)
);

BUFx5_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_45),
.Y(n_153)
);

INVx3_ASAP7_75t_L g181 ( 
.A(n_45),
.Y(n_181)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_45),
.Y(n_225)
);

INVx6_ASAP7_75t_L g447 ( 
.A(n_45),
.Y(n_447)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

XNOR2xp5_ASAP7_75t_L g47 ( 
.A(n_48),
.B(n_50),
.Y(n_47)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_49),
.Y(n_93)
);

CKINVDCx16_ASAP7_75t_R g51 ( 
.A(n_52),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_53),
.B(n_54),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_53),
.B(n_156),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_54),
.B(n_92),
.Y(n_127)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g285 ( 
.A(n_55),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g57 ( 
.A(n_58),
.B(n_62),
.C(n_66),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_58),
.A2(n_59),
.B1(n_118),
.B2(n_119),
.Y(n_117)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

MAJIxp5_ASAP7_75t_L g66 ( 
.A(n_61),
.B(n_67),
.C(n_72),
.Y(n_66)
);

XOR2xp5_ASAP7_75t_L g119 ( 
.A(n_62),
.B(n_66),
.Y(n_119)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_67),
.A2(n_68),
.B1(n_114),
.B2(n_115),
.Y(n_113)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_71),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_72),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_72),
.A2(n_107),
.B1(n_108),
.B2(n_111),
.Y(n_184)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx5_ASAP7_75t_L g335 ( 
.A(n_74),
.Y(n_335)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx5_ASAP7_75t_L g134 ( 
.A(n_75),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_75),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g363 ( 
.A(n_75),
.Y(n_363)
);

INVx6_ASAP7_75t_L g417 ( 
.A(n_75),
.Y(n_417)
);

INVx11_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

BUFx5_ASAP7_75t_L g235 ( 
.A(n_76),
.Y(n_235)
);

INVx3_ASAP7_75t_L g253 ( 
.A(n_76),
.Y(n_253)
);

BUFx3_ASAP7_75t_L g264 ( 
.A(n_76),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_116),
.C(n_117),
.Y(n_77)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_78),
.B(n_191),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_103),
.C(n_112),
.Y(n_78)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_79),
.B(n_188),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_SL g79 ( 
.A(n_80),
.B(n_94),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_80),
.B(n_96),
.C(n_102),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_85),
.C(n_91),
.Y(n_80)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_81),
.B(n_85),
.Y(n_162)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx6_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx8_ASAP7_75t_L g267 ( 
.A(n_89),
.Y(n_267)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_91),
.B(n_162),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_93),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_92),
.B(n_270),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_95),
.A2(n_96),
.B1(n_97),
.B2(n_102),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_95),
.Y(n_102)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

HB1xp67_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_103),
.A2(n_112),
.B1(n_113),
.B2(n_189),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_103),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_107),
.C(n_111),
.Y(n_103)
);

XOR2xp5_ASAP7_75t_L g183 ( 
.A(n_104),
.B(n_184),
.Y(n_183)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_107),
.A2(n_108),
.B1(n_155),
.B2(n_160),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_107),
.B(n_150),
.C(n_160),
.Y(n_185)
);

CKINVDCx14_ASAP7_75t_R g107 ( 
.A(n_108),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_116),
.B(n_117),
.Y(n_191)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

AO21x1_ASAP7_75t_L g121 ( 
.A1(n_122),
.A2(n_192),
.B(n_536),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_190),
.Y(n_122)
);

OR2x2_ASAP7_75t_L g537 ( 
.A(n_123),
.B(n_190),
.Y(n_537)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_182),
.C(n_187),
.Y(n_123)
);

XOR2xp5_ASAP7_75t_L g521 ( 
.A(n_124),
.B(n_522),
.Y(n_521)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_161),
.C(n_163),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_SL g524 ( 
.A(n_125),
.B(n_525),
.Y(n_524)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_136),
.C(n_149),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_L g514 ( 
.A(n_126),
.B(n_136),
.Y(n_514)
);

XNOR2xp5_ASAP7_75t_SL g126 ( 
.A(n_127),
.B(n_128),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_127),
.B(n_130),
.C(n_135),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_129),
.A2(n_130),
.B1(n_131),
.B2(n_135),
.Y(n_128)
);

CKINVDCx14_ASAP7_75t_R g135 ( 
.A(n_129),
.Y(n_135)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

BUFx3_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx5_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_SL g484 ( 
.A(n_136),
.B(n_485),
.Y(n_484)
);

MAJIxp5_ASAP7_75t_L g506 ( 
.A(n_136),
.B(n_481),
.C(n_485),
.Y(n_506)
);

FAx1_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_141),
.CI(n_144),
.CON(n_136),
.SN(n_136)
);

INVx4_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVx6_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

BUFx3_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVx4_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVx4_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g250 ( 
.A(n_148),
.Y(n_250)
);

INVx5_ASAP7_75t_L g305 ( 
.A(n_148),
.Y(n_305)
);

XOR2xp5_ASAP7_75t_L g513 ( 
.A(n_149),
.B(n_514),
.Y(n_513)
);

XNOR2xp5_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_154),
.Y(n_149)
);

INVx5_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_152),
.Y(n_215)
);

INVx6_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_155),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_155),
.B(n_166),
.C(n_170),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g483 ( 
.A1(n_155),
.A2(n_160),
.B1(n_166),
.B2(n_167),
.Y(n_483)
);

INVx3_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

INVx4_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g208 ( 
.A(n_159),
.Y(n_208)
);

BUFx3_ASAP7_75t_L g341 ( 
.A(n_159),
.Y(n_341)
);

AOI22xp5_ASAP7_75t_L g525 ( 
.A1(n_161),
.A2(n_163),
.B1(n_164),
.B2(n_526),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_161),
.Y(n_526)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_174),
.C(n_177),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g511 ( 
.A(n_165),
.B(n_512),
.Y(n_511)
);

AOI22xp5_ASAP7_75t_L g465 ( 
.A1(n_166),
.A2(n_167),
.B1(n_466),
.B2(n_468),
.Y(n_465)
);

MAJIxp5_ASAP7_75t_L g485 ( 
.A(n_166),
.B(n_466),
.C(n_469),
.Y(n_485)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_167),
.Y(n_166)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

INVx3_ASAP7_75t_L g213 ( 
.A(n_169),
.Y(n_213)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_169),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_SL g482 ( 
.A(n_170),
.B(n_483),
.Y(n_482)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_172),
.Y(n_170)
);

INVx4_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_173),
.Y(n_218)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_173),
.Y(n_422)
);

OAI22xp5_ASAP7_75t_L g512 ( 
.A1(n_174),
.A2(n_175),
.B1(n_177),
.B2(n_178),
.Y(n_512)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g493 ( 
.A1(n_177),
.A2(n_178),
.B1(n_494),
.B2(n_496),
.Y(n_493)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_178),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g509 ( 
.A(n_178),
.B(n_496),
.C(n_510),
.Y(n_509)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

INVx4_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

INVx4_ASAP7_75t_L g259 ( 
.A(n_181),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g522 ( 
.A(n_182),
.B(n_187),
.Y(n_522)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_185),
.C(n_186),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g527 ( 
.A(n_183),
.B(n_528),
.Y(n_527)
);

XNOR2xp5_ASAP7_75t_L g528 ( 
.A(n_185),
.B(n_186),
.Y(n_528)
);

AO21x1_ASAP7_75t_L g192 ( 
.A1(n_193),
.A2(n_517),
.B(n_533),
.Y(n_192)
);

OAI21x1_ASAP7_75t_L g193 ( 
.A1(n_194),
.A2(n_501),
.B(n_516),
.Y(n_193)
);

AOI21x1_ASAP7_75t_L g194 ( 
.A1(n_195),
.A2(n_476),
.B(n_500),
.Y(n_194)
);

OAI21x1_ASAP7_75t_L g195 ( 
.A1(n_196),
.A2(n_430),
.B(n_475),
.Y(n_195)
);

AOI21x1_ASAP7_75t_L g196 ( 
.A1(n_197),
.A2(n_392),
.B(n_429),
.Y(n_196)
);

AO21x1_ASAP7_75t_L g197 ( 
.A1(n_198),
.A2(n_315),
.B(n_391),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_199),
.B(n_295),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g391 ( 
.A(n_199),
.B(n_295),
.Y(n_391)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_200),
.A2(n_201),
.B1(n_242),
.B2(n_294),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g428 ( 
.A(n_200),
.B(n_243),
.C(n_277),
.Y(n_428)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_219),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g395 ( 
.A(n_202),
.B(n_220),
.C(n_241),
.Y(n_395)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_214),
.C(n_216),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g313 ( 
.A(n_203),
.B(n_314),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_209),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_204),
.A2(n_205),
.B1(n_209),
.B2(n_210),
.Y(n_300)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

INVx6_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

BUFx6f_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

INVx3_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_214),
.B(n_216),
.Y(n_314)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_220),
.A2(n_227),
.B1(n_240),
.B2(n_241),
.Y(n_219)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_220),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_L g220 ( 
.A1(n_221),
.A2(n_222),
.B(n_226),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_221),
.B(n_222),
.Y(n_226)
);

INVx4_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

INVx3_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_SL g407 ( 
.A(n_226),
.B(n_408),
.Y(n_407)
);

MAJIxp5_ASAP7_75t_L g437 ( 
.A(n_226),
.B(n_397),
.C(n_408),
.Y(n_437)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_227),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_232),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g427 ( 
.A(n_228),
.B(n_233),
.C(n_236),
.Y(n_427)
);

INVx3_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

INVx4_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_236),
.Y(n_232)
);

INVx5_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

INVx8_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

BUFx5_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_242),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_SL g242 ( 
.A(n_243),
.B(n_277),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_254),
.C(n_268),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g296 ( 
.A(n_244),
.B(n_297),
.Y(n_296)
);

BUFx24_ASAP7_75t_SL g539 ( 
.A(n_244),
.Y(n_539)
);

FAx1_ASAP7_75t_SL g244 ( 
.A(n_245),
.B(n_248),
.CI(n_251),
.CON(n_244),
.SN(n_244)
);

MAJx2_ASAP7_75t_L g293 ( 
.A(n_245),
.B(n_248),
.C(n_251),
.Y(n_293)
);

BUFx6f_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

BUFx6f_ASAP7_75t_L g280 ( 
.A(n_247),
.Y(n_280)
);

INVx4_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

BUFx6f_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

INVx3_ASAP7_75t_L g454 ( 
.A(n_253),
.Y(n_454)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_254),
.A2(n_255),
.B1(n_268),
.B2(n_298),
.Y(n_297)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

MAJx2_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_260),
.C(n_265),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g384 ( 
.A1(n_256),
.A2(n_257),
.B1(n_265),
.B2(n_266),
.Y(n_384)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

INVx8_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g383 ( 
.A(n_260),
.B(n_384),
.Y(n_383)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_268),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_273),
.Y(n_268)
);

AND2x2_ASAP7_75t_L g292 ( 
.A(n_269),
.B(n_273),
.Y(n_292)
);

INVx8_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

BUFx8_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

INVx2_ASAP7_75t_L g288 ( 
.A(n_272),
.Y(n_288)
);

BUFx5_ASAP7_75t_L g312 ( 
.A(n_272),
.Y(n_312)
);

BUFx3_ASAP7_75t_L g406 ( 
.A(n_272),
.Y(n_406)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

INVx3_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

INVx2_ASAP7_75t_L g351 ( 
.A(n_276),
.Y(n_351)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_278),
.B(n_291),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g411 ( 
.A(n_278),
.B(n_292),
.C(n_293),
.Y(n_411)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_279),
.B(n_281),
.Y(n_278)
);

MAJx2_ASAP7_75t_L g408 ( 
.A(n_279),
.B(n_286),
.C(n_289),
.Y(n_408)
);

AOI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_282),
.A2(n_286),
.B1(n_289),
.B2(n_290),
.Y(n_281)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_282),
.Y(n_289)
);

INVx3_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

INVx8_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

CKINVDCx16_ASAP7_75t_R g290 ( 
.A(n_286),
.Y(n_290)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

XOR2xp5_ASAP7_75t_L g291 ( 
.A(n_292),
.B(n_293),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_296),
.B(n_299),
.C(n_313),
.Y(n_295)
);

XOR2xp5_ASAP7_75t_L g388 ( 
.A(n_296),
.B(n_389),
.Y(n_388)
);

XOR2xp5_ASAP7_75t_L g389 ( 
.A(n_299),
.B(n_313),
.Y(n_389)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_300),
.B(n_301),
.C(n_306),
.Y(n_299)
);

XOR2xp5_ASAP7_75t_L g377 ( 
.A(n_300),
.B(n_301),
.Y(n_377)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

BUFx6f_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g376 ( 
.A(n_306),
.B(n_377),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_SL g306 ( 
.A(n_307),
.B(n_311),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g357 ( 
.A(n_307),
.B(n_311),
.Y(n_357)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

OAI21x1_ASAP7_75t_L g315 ( 
.A1(n_316),
.A2(n_386),
.B(n_390),
.Y(n_315)
);

OA21x2_ASAP7_75t_L g316 ( 
.A1(n_317),
.A2(n_371),
.B(n_385),
.Y(n_316)
);

AOI21xp5_ASAP7_75t_L g317 ( 
.A1(n_318),
.A2(n_354),
.B(n_370),
.Y(n_317)
);

OAI21xp5_ASAP7_75t_SL g318 ( 
.A1(n_319),
.A2(n_344),
.B(n_353),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_320),
.B(n_327),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_320),
.B(n_327),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_321),
.B(n_324),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_L g346 ( 
.A(n_321),
.B(n_324),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_L g348 ( 
.A(n_321),
.B(n_349),
.Y(n_348)
);

BUFx6f_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

BUFx5_ASAP7_75t_L g467 ( 
.A(n_323),
.Y(n_467)
);

INVx3_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_L g327 ( 
.A1(n_328),
.A2(n_329),
.B1(n_336),
.B2(n_337),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

XOR2xp5_ASAP7_75t_L g329 ( 
.A(n_330),
.B(n_332),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g369 ( 
.A(n_330),
.B(n_332),
.C(n_336),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_333),
.B(n_334),
.Y(n_332)
);

INVx3_ASAP7_75t_L g334 ( 
.A(n_335),
.Y(n_334)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_337),
.Y(n_336)
);

XNOR2xp5_ASAP7_75t_SL g337 ( 
.A(n_338),
.B(n_342),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_338),
.B(n_342),
.Y(n_358)
);

BUFx3_ASAP7_75t_L g339 ( 
.A(n_340),
.Y(n_339)
);

INVx2_ASAP7_75t_L g340 ( 
.A(n_341),
.Y(n_340)
);

AOI21xp5_ASAP7_75t_L g344 ( 
.A1(n_345),
.A2(n_348),
.B(n_352),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_SL g345 ( 
.A(n_346),
.B(n_347),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_L g352 ( 
.A(n_346),
.B(n_347),
.Y(n_352)
);

INVx2_ASAP7_75t_L g350 ( 
.A(n_351),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_SL g354 ( 
.A(n_355),
.B(n_369),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_L g370 ( 
.A(n_355),
.B(n_369),
.Y(n_370)
);

XNOR2xp5_ASAP7_75t_L g355 ( 
.A(n_356),
.B(n_359),
.Y(n_355)
);

XOR2xp5_ASAP7_75t_L g356 ( 
.A(n_357),
.B(n_358),
.Y(n_356)
);

MAJIxp5_ASAP7_75t_L g372 ( 
.A(n_357),
.B(n_358),
.C(n_373),
.Y(n_372)
);

INVxp67_ASAP7_75t_L g373 ( 
.A(n_359),
.Y(n_373)
);

XNOR2xp5_ASAP7_75t_SL g359 ( 
.A(n_360),
.B(n_364),
.Y(n_359)
);

MAJIxp5_ASAP7_75t_L g381 ( 
.A(n_360),
.B(n_366),
.C(n_368),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_L g360 ( 
.A(n_361),
.B(n_362),
.Y(n_360)
);

INVx11_ASAP7_75t_L g362 ( 
.A(n_363),
.Y(n_362)
);

AOI22xp5_ASAP7_75t_L g364 ( 
.A1(n_365),
.A2(n_366),
.B1(n_367),
.B2(n_368),
.Y(n_364)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_365),
.Y(n_368)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_367),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_L g371 ( 
.A(n_372),
.B(n_374),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_372),
.B(n_374),
.Y(n_385)
);

OAI22xp5_ASAP7_75t_SL g374 ( 
.A1(n_375),
.A2(n_376),
.B1(n_378),
.B2(n_379),
.Y(n_374)
);

MAJIxp5_ASAP7_75t_L g387 ( 
.A(n_375),
.B(n_381),
.C(n_382),
.Y(n_387)
);

INVx1_ASAP7_75t_SL g375 ( 
.A(n_376),
.Y(n_375)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_379),
.Y(n_378)
);

AOI22xp5_ASAP7_75t_L g379 ( 
.A1(n_380),
.A2(n_381),
.B1(n_382),
.B2(n_383),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_381),
.Y(n_380)
);

INVx1_ASAP7_75t_SL g382 ( 
.A(n_383),
.Y(n_382)
);

NOR2xp33_ASAP7_75t_L g386 ( 
.A(n_387),
.B(n_388),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_387),
.B(n_388),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_SL g392 ( 
.A(n_393),
.B(n_428),
.Y(n_392)
);

NOR2xp33_ASAP7_75t_L g429 ( 
.A(n_393),
.B(n_428),
.Y(n_429)
);

XNOR2xp5_ASAP7_75t_L g393 ( 
.A(n_394),
.B(n_410),
.Y(n_393)
);

XNOR2xp5_ASAP7_75t_L g394 ( 
.A(n_395),
.B(n_396),
.Y(n_394)
);

MAJIxp5_ASAP7_75t_L g431 ( 
.A(n_395),
.B(n_396),
.C(n_410),
.Y(n_431)
);

AOI22xp5_ASAP7_75t_L g396 ( 
.A1(n_397),
.A2(n_398),
.B1(n_407),
.B2(n_409),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_398),
.Y(n_397)
);

XNOR2xp5_ASAP7_75t_SL g398 ( 
.A(n_399),
.B(n_400),
.Y(n_398)
);

MAJIxp5_ASAP7_75t_L g448 ( 
.A(n_399),
.B(n_402),
.C(n_404),
.Y(n_448)
);

OAI22xp5_ASAP7_75t_SL g400 ( 
.A1(n_401),
.A2(n_402),
.B1(n_404),
.B2(n_405),
.Y(n_400)
);

CKINVDCx20_ASAP7_75t_R g401 ( 
.A(n_402),
.Y(n_401)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_405),
.Y(n_404)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_407),
.Y(n_409)
);

XNOR2xp5_ASAP7_75t_SL g410 ( 
.A(n_411),
.B(n_412),
.Y(n_410)
);

MAJIxp5_ASAP7_75t_L g433 ( 
.A(n_411),
.B(n_413),
.C(n_423),
.Y(n_433)
);

XNOR2xp5_ASAP7_75t_L g412 ( 
.A(n_413),
.B(n_423),
.Y(n_412)
);

XNOR2xp5_ASAP7_75t_L g413 ( 
.A(n_414),
.B(n_418),
.Y(n_413)
);

MAJIxp5_ASAP7_75t_L g462 ( 
.A(n_414),
.B(n_419),
.C(n_420),
.Y(n_462)
);

BUFx2_ASAP7_75t_L g415 ( 
.A(n_416),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_417),
.Y(n_416)
);

XNOR2xp5_ASAP7_75t_L g418 ( 
.A(n_419),
.B(n_420),
.Y(n_418)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_422),
.Y(n_421)
);

XNOR2xp5_ASAP7_75t_L g423 ( 
.A(n_424),
.B(n_427),
.Y(n_423)
);

XNOR2xp5_ASAP7_75t_L g424 ( 
.A(n_425),
.B(n_426),
.Y(n_424)
);

MAJIxp5_ASAP7_75t_L g439 ( 
.A(n_425),
.B(n_426),
.C(n_427),
.Y(n_439)
);

NOR2xp33_ASAP7_75t_L g430 ( 
.A(n_431),
.B(n_432),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_431),
.B(n_432),
.Y(n_475)
);

XNOR2xp5_ASAP7_75t_L g432 ( 
.A(n_433),
.B(n_434),
.Y(n_432)
);

MAJIxp5_ASAP7_75t_L g499 ( 
.A(n_433),
.B(n_450),
.C(n_473),
.Y(n_499)
);

AOI22xp5_ASAP7_75t_SL g434 ( 
.A1(n_435),
.A2(n_450),
.B1(n_473),
.B2(n_474),
.Y(n_434)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_435),
.Y(n_473)
);

AOI22xp5_ASAP7_75t_L g435 ( 
.A1(n_436),
.A2(n_437),
.B1(n_438),
.B2(n_449),
.Y(n_435)
);

MAJIxp5_ASAP7_75t_L g478 ( 
.A(n_436),
.B(n_439),
.C(n_440),
.Y(n_478)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_437),
.Y(n_436)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_438),
.Y(n_449)
);

XNOR2xp5_ASAP7_75t_SL g438 ( 
.A(n_439),
.B(n_440),
.Y(n_438)
);

XNOR2xp5_ASAP7_75t_L g440 ( 
.A(n_441),
.B(n_448),
.Y(n_440)
);

XOR2xp5_ASAP7_75t_L g441 ( 
.A(n_442),
.B(n_443),
.Y(n_441)
);

MAJIxp5_ASAP7_75t_L g491 ( 
.A(n_442),
.B(n_443),
.C(n_448),
.Y(n_491)
);

INVx6_ASAP7_75t_L g444 ( 
.A(n_445),
.Y(n_444)
);

INVx5_ASAP7_75t_L g445 ( 
.A(n_446),
.Y(n_445)
);

BUFx6f_ASAP7_75t_L g446 ( 
.A(n_447),
.Y(n_446)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_450),
.Y(n_474)
);

XNOR2xp5_ASAP7_75t_L g450 ( 
.A(n_451),
.B(n_461),
.Y(n_450)
);

MAJIxp5_ASAP7_75t_L g489 ( 
.A(n_451),
.B(n_462),
.C(n_463),
.Y(n_489)
);

BUFx24_ASAP7_75t_SL g542 ( 
.A(n_451),
.Y(n_542)
);

FAx1_ASAP7_75t_SL g451 ( 
.A(n_452),
.B(n_455),
.CI(n_457),
.CON(n_451),
.SN(n_451)
);

MAJIxp5_ASAP7_75t_L g497 ( 
.A(n_452),
.B(n_455),
.C(n_457),
.Y(n_497)
);

INVx5_ASAP7_75t_L g453 ( 
.A(n_454),
.Y(n_453)
);

INVx2_ASAP7_75t_L g458 ( 
.A(n_459),
.Y(n_458)
);

INVx2_ASAP7_75t_L g459 ( 
.A(n_460),
.Y(n_459)
);

XNOR2xp5_ASAP7_75t_L g461 ( 
.A(n_462),
.B(n_463),
.Y(n_461)
);

OAI22xp5_ASAP7_75t_SL g463 ( 
.A1(n_464),
.A2(n_465),
.B1(n_469),
.B2(n_470),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_465),
.Y(n_464)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_466),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_470),
.Y(n_469)
);

INVx2_ASAP7_75t_L g471 ( 
.A(n_472),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_SL g476 ( 
.A(n_477),
.B(n_499),
.Y(n_476)
);

NOR2xp33_ASAP7_75t_L g500 ( 
.A(n_477),
.B(n_499),
.Y(n_500)
);

XNOR2xp5_ASAP7_75t_L g477 ( 
.A(n_478),
.B(n_479),
.Y(n_477)
);

MAJIxp5_ASAP7_75t_L g515 ( 
.A(n_478),
.B(n_480),
.C(n_487),
.Y(n_515)
);

XNOR2xp5_ASAP7_75t_L g479 ( 
.A(n_480),
.B(n_487),
.Y(n_479)
);

AOI22xp5_ASAP7_75t_L g480 ( 
.A1(n_481),
.A2(n_482),
.B1(n_484),
.B2(n_486),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_482),
.Y(n_481)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_484),
.Y(n_486)
);

AOI22xp5_ASAP7_75t_L g487 ( 
.A1(n_488),
.A2(n_489),
.B1(n_490),
.B2(n_498),
.Y(n_487)
);

MAJIxp5_ASAP7_75t_L g503 ( 
.A(n_488),
.B(n_491),
.C(n_492),
.Y(n_503)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_489),
.Y(n_488)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_490),
.Y(n_498)
);

XNOR2xp5_ASAP7_75t_SL g490 ( 
.A(n_491),
.B(n_492),
.Y(n_490)
);

XNOR2xp5_ASAP7_75t_L g492 ( 
.A(n_493),
.B(n_497),
.Y(n_492)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_494),
.Y(n_496)
);

INVxp67_ASAP7_75t_L g510 ( 
.A(n_497),
.Y(n_510)
);

NOR2xp33_ASAP7_75t_SL g501 ( 
.A(n_502),
.B(n_515),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_502),
.B(n_515),
.Y(n_516)
);

BUFx24_ASAP7_75t_SL g540 ( 
.A(n_502),
.Y(n_540)
);

FAx1_ASAP7_75t_L g502 ( 
.A(n_503),
.B(n_504),
.CI(n_513),
.CON(n_502),
.SN(n_502)
);

MAJIxp5_ASAP7_75t_L g532 ( 
.A(n_503),
.B(n_504),
.C(n_513),
.Y(n_532)
);

AOI22xp5_ASAP7_75t_L g504 ( 
.A1(n_505),
.A2(n_506),
.B1(n_507),
.B2(n_508),
.Y(n_504)
);

MAJIxp5_ASAP7_75t_L g529 ( 
.A(n_505),
.B(n_509),
.C(n_511),
.Y(n_529)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_506),
.Y(n_505)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_508),
.Y(n_507)
);

XOR2xp5_ASAP7_75t_L g508 ( 
.A(n_509),
.B(n_511),
.Y(n_508)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_518),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_519),
.B(n_530),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_520),
.Y(n_519)
);

OAI21xp5_ASAP7_75t_L g533 ( 
.A1(n_520),
.A2(n_534),
.B(n_535),
.Y(n_533)
);

NOR2xp33_ASAP7_75t_SL g520 ( 
.A(n_521),
.B(n_523),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_521),
.B(n_523),
.Y(n_535)
);

MAJIxp5_ASAP7_75t_L g523 ( 
.A(n_524),
.B(n_527),
.C(n_529),
.Y(n_523)
);

FAx1_ASAP7_75t_SL g531 ( 
.A(n_524),
.B(n_527),
.CI(n_529),
.CON(n_531),
.SN(n_531)
);

OR2x2_ASAP7_75t_L g530 ( 
.A(n_531),
.B(n_532),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_L g534 ( 
.A(n_531),
.B(n_532),
.Y(n_534)
);

BUFx24_ASAP7_75t_SL g538 ( 
.A(n_531),
.Y(n_538)
);

CKINVDCx20_ASAP7_75t_R g536 ( 
.A(n_537),
.Y(n_536)
);


endmodule