module real_jpeg_24432_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_288;
wire n_83;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_312;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

AOI22xp33_ASAP7_75t_SL g33 ( 
.A1(n_0),
.A2(n_26),
.B1(n_27),
.B2(n_34),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

AOI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_0),
.A2(n_34),
.B1(n_39),
.B2(n_41),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_1),
.A2(n_55),
.B1(n_56),
.B2(n_57),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_1),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_1),
.A2(n_57),
.B1(n_60),
.B2(n_65),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_1),
.A2(n_39),
.B1(n_41),
.B2(n_57),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_L g211 ( 
.A1(n_1),
.A2(n_26),
.B1(n_27),
.B2(n_57),
.Y(n_211)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_2),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_3),
.A2(n_60),
.B1(n_65),
.B2(n_86),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_3),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_3),
.A2(n_39),
.B1(n_41),
.B2(n_86),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_3),
.A2(n_55),
.B1(n_86),
.B2(n_132),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_L g178 ( 
.A1(n_3),
.A2(n_26),
.B1(n_27),
.B2(n_86),
.Y(n_178)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_4),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_L g37 ( 
.A1(n_6),
.A2(n_38),
.B1(n_39),
.B2(n_41),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_6),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_6),
.A2(n_38),
.B1(n_60),
.B2(n_65),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_6),
.A2(n_26),
.B1(n_27),
.B2(n_38),
.Y(n_156)
);

INVx8_ASAP7_75t_SL g64 ( 
.A(n_7),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g47 ( 
.A1(n_8),
.A2(n_39),
.B1(n_41),
.B2(n_48),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_8),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_8),
.A2(n_26),
.B1(n_27),
.B2(n_48),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_8),
.A2(n_48),
.B1(n_60),
.B2(n_65),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_9),
.A2(n_56),
.B1(n_75),
.B2(n_108),
.Y(n_107)
);

CKINVDCx16_ASAP7_75t_R g108 ( 
.A(n_9),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_9),
.A2(n_60),
.B1(n_65),
.B2(n_108),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g236 ( 
.A1(n_9),
.A2(n_39),
.B1(n_41),
.B2(n_108),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_9),
.A2(n_26),
.B1(n_27),
.B2(n_108),
.Y(n_261)
);

BUFx5_ASAP7_75t_L g82 ( 
.A(n_10),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_11),
.B(n_173),
.Y(n_172)
);

INVx1_ASAP7_75t_SL g202 ( 
.A(n_11),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_11),
.B(n_59),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_11),
.B(n_39),
.C(n_82),
.Y(n_227)
);

AOI22xp33_ASAP7_75t_SL g239 ( 
.A1(n_11),
.A2(n_60),
.B1(n_65),
.B2(n_202),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_11),
.B(n_123),
.Y(n_257)
);

AOI22xp33_ASAP7_75t_SL g267 ( 
.A1(n_11),
.A2(n_39),
.B1(n_41),
.B2(n_202),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_11),
.B(n_26),
.C(n_44),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_L g290 ( 
.A1(n_11),
.A2(n_25),
.B(n_262),
.Y(n_290)
);

INVx13_ASAP7_75t_L g55 ( 
.A(n_12),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_L g69 ( 
.A1(n_13),
.A2(n_70),
.B1(n_71),
.B2(n_72),
.Y(n_69)
);

CKINVDCx16_ASAP7_75t_R g71 ( 
.A(n_13),
.Y(n_71)
);

OAI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_13),
.A2(n_60),
.B1(n_65),
.B2(n_71),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_13),
.A2(n_39),
.B1(n_41),
.B2(n_71),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_13),
.A2(n_26),
.B1(n_27),
.B2(n_71),
.Y(n_232)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_14),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_15),
.A2(n_70),
.B1(n_76),
.B2(n_148),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_15),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_15),
.A2(n_60),
.B1(n_65),
.B2(n_148),
.Y(n_195)
);

AOI22xp33_ASAP7_75t_L g235 ( 
.A1(n_15),
.A2(n_39),
.B1(n_41),
.B2(n_148),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_15),
.A2(n_26),
.B1(n_27),
.B2(n_148),
.Y(n_274)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_16),
.Y(n_29)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_16),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_16),
.B(n_263),
.Y(n_262)
);

INVx3_ASAP7_75t_L g284 ( 
.A(n_16),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_138),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_136),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_112),
.Y(n_20)
);

AND2x2_ASAP7_75t_L g137 ( 
.A(n_21),
.B(n_112),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_77),
.C(n_93),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_22),
.A2(n_77),
.B1(n_78),
.B2(n_317),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_22),
.Y(n_317)
);

XOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_50),
.Y(n_22)
);

AOI21xp33_ASAP7_75t_L g113 ( 
.A1(n_23),
.A2(n_24),
.B(n_52),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_35),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_24),
.A2(n_51),
.B1(n_52),
.B2(n_53),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_24),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_24),
.A2(n_35),
.B1(n_36),
.B2(n_51),
.Y(n_182)
);

AOI21xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_30),
.B(n_33),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_25),
.A2(n_30),
.B1(n_33),
.B2(n_98),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_25),
.A2(n_98),
.B1(n_155),
.B2(n_157),
.Y(n_154)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_25),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_25),
.A2(n_178),
.B1(n_211),
.B2(n_212),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_25),
.B(n_232),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_L g260 ( 
.A1(n_25),
.A2(n_261),
.B(n_262),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_29),
.Y(n_25)
);

OA22x2_ASAP7_75t_L g46 ( 
.A1(n_26),
.A2(n_27),
.B1(n_44),
.B2(n_45),
.Y(n_46)
);

INVx2_ASAP7_75t_SL g26 ( 
.A(n_27),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_27),
.B(n_288),
.Y(n_287)
);

INVx6_ASAP7_75t_SL g27 ( 
.A(n_28),
.Y(n_27)
);

INVx8_ASAP7_75t_L g158 ( 
.A(n_29),
.Y(n_158)
);

INVx5_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx5_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_32),
.Y(n_230)
);

CKINVDCx16_ASAP7_75t_R g35 ( 
.A(n_36),
.Y(n_35)
);

AOI22xp5_ASAP7_75t_L g36 ( 
.A1(n_37),
.A2(n_42),
.B1(n_47),
.B2(n_49),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_37),
.A2(n_42),
.B1(n_49),
.B2(n_101),
.Y(n_100)
);

INVx4_ASAP7_75t_SL g41 ( 
.A(n_39),
.Y(n_41)
);

OAI22xp33_ASAP7_75t_L g43 ( 
.A1(n_39),
.A2(n_41),
.B1(n_44),
.B2(n_45),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_39),
.A2(n_41),
.B1(n_82),
.B2(n_83),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_39),
.B(n_269),
.Y(n_268)
);

BUFx4f_ASAP7_75t_SL g39 ( 
.A(n_40),
.Y(n_39)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_42),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_L g127 ( 
.A1(n_42),
.A2(n_49),
.B(n_128),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_42),
.B(n_199),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_42),
.A2(n_49),
.B1(n_234),
.B2(n_236),
.Y(n_233)
);

AND2x2_ASAP7_75t_L g42 ( 
.A(n_43),
.B(n_46),
.Y(n_42)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_44),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_46),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_46),
.A2(n_89),
.B1(n_90),
.B2(n_91),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_46),
.A2(n_89),
.B1(n_102),
.B2(n_160),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_L g197 ( 
.A1(n_46),
.A2(n_160),
.B(n_198),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_L g259 ( 
.A1(n_46),
.A2(n_198),
.B(n_235),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_46),
.B(n_202),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_47),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_49),
.B(n_199),
.Y(n_250)
);

CKINVDCx14_ASAP7_75t_R g52 ( 
.A(n_53),
.Y(n_52)
);

OAI21xp5_ASAP7_75t_L g53 ( 
.A1(n_54),
.A2(n_58),
.B(n_67),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_54),
.A2(n_58),
.B1(n_109),
.B2(n_131),
.Y(n_130)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_55),
.Y(n_56)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_55),
.Y(n_72)
);

INVx11_ASAP7_75t_L g76 ( 
.A(n_55),
.Y(n_76)
);

INVx6_ASAP7_75t_L g134 ( 
.A(n_55),
.Y(n_134)
);

INVx11_ASAP7_75t_L g70 ( 
.A(n_56),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_58),
.B(n_74),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_58),
.B(n_69),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_L g164 ( 
.A1(n_58),
.A2(n_67),
.B(n_165),
.Y(n_164)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_59),
.A2(n_73),
.B1(n_107),
.B2(n_147),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_60),
.A2(n_63),
.B1(n_65),
.B2(n_66),
.Y(n_59)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_60),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_60),
.A2(n_65),
.B1(n_82),
.B2(n_83),
.Y(n_84)
);

NAND2xp33_ASAP7_75t_SL g174 ( 
.A(n_60),
.B(n_66),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_60),
.B(n_227),
.Y(n_226)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_63),
.Y(n_66)
);

OAI22xp33_ASAP7_75t_L g74 ( 
.A1(n_63),
.A2(n_66),
.B1(n_75),
.B2(n_76),
.Y(n_74)
);

AOI32xp33_ASAP7_75t_L g171 ( 
.A1(n_63),
.A2(n_65),
.A3(n_76),
.B1(n_172),
.B2(n_174),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_68),
.B(n_73),
.Y(n_67)
);

INVxp67_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx4_ASAP7_75t_L g173 ( 
.A(n_72),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_73),
.Y(n_109)
);

AOI21xp5_ASAP7_75t_L g200 ( 
.A1(n_73),
.A2(n_111),
.B(n_201),
.Y(n_200)
);

INVx8_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

OAI21xp33_ASAP7_75t_L g201 ( 
.A1(n_76),
.A2(n_202),
.B(n_203),
.Y(n_201)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

AOI21xp5_ASAP7_75t_L g78 ( 
.A1(n_79),
.A2(n_88),
.B(n_92),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_79),
.B(n_88),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_80),
.A2(n_81),
.B1(n_85),
.B2(n_87),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_80),
.A2(n_81),
.B1(n_85),
.B2(n_104),
.Y(n_103)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_80),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_SL g166 ( 
.A1(n_80),
.A2(n_167),
.B(n_169),
.Y(n_166)
);

OAI21xp33_ASAP7_75t_L g238 ( 
.A1(n_80),
.A2(n_169),
.B(n_239),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_84),
.Y(n_80)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_81),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_L g150 ( 
.A1(n_81),
.A2(n_104),
.B(n_151),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_SL g206 ( 
.A1(n_81),
.A2(n_151),
.B(n_207),
.Y(n_206)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_82),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_87),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_SL g248 ( 
.A1(n_89),
.A2(n_249),
.B(n_250),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_SL g266 ( 
.A1(n_89),
.A2(n_250),
.B(n_267),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_91),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_92),
.A2(n_115),
.B1(n_116),
.B2(n_117),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_92),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_93),
.A2(n_94),
.B1(n_316),
.B2(n_318),
.Y(n_315)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_103),
.C(n_105),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_95),
.A2(n_96),
.B1(n_184),
.B2(n_185),
.Y(n_183)
);

CKINVDCx16_ASAP7_75t_R g95 ( 
.A(n_96),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_99),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_97),
.A2(n_99),
.B1(n_100),
.B2(n_162),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_97),
.Y(n_162)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_102),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_SL g185 ( 
.A(n_103),
.B(n_105),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_L g105 ( 
.A1(n_106),
.A2(n_109),
.B(n_110),
.Y(n_105)
);

CKINVDCx16_ASAP7_75t_R g106 ( 
.A(n_107),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

XOR2xp5_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_114),
.Y(n_112)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_118),
.A2(n_119),
.B1(n_130),
.B2(n_135),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_120),
.A2(n_126),
.B1(n_127),
.B2(n_129),
.Y(n_119)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_120),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_121),
.A2(n_122),
.B1(n_123),
.B2(n_124),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_122),
.B(n_152),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_122),
.A2(n_123),
.B1(n_168),
.B2(n_195),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_123),
.B(n_152),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_125),
.Y(n_124)
);

CKINVDCx16_ASAP7_75t_R g126 ( 
.A(n_127),
.Y(n_126)
);

CKINVDCx14_ASAP7_75t_R g135 ( 
.A(n_130),
.Y(n_135)
);

INVx8_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx8_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

CKINVDCx16_ASAP7_75t_R g136 ( 
.A(n_137),
.Y(n_136)
);

AOI21xp5_ASAP7_75t_L g138 ( 
.A1(n_139),
.A2(n_314),
.B(n_320),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_L g139 ( 
.A1(n_140),
.A2(n_187),
.B(n_313),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_180),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_141),
.B(n_180),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_161),
.C(n_163),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_142),
.A2(n_143),
.B1(n_161),
.B2(n_311),
.Y(n_310)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

XOR2xp5_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_153),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_145),
.A2(n_146),
.B1(n_149),
.B2(n_150),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_146),
.B(n_149),
.C(n_153),
.Y(n_186)
);

CKINVDCx16_ASAP7_75t_R g165 ( 
.A(n_147),
.Y(n_165)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_159),
.Y(n_153)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_154),
.B(n_159),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_156),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_156),
.A2(n_176),
.B1(n_177),
.B2(n_179),
.Y(n_175)
);

INVx3_ASAP7_75t_L g179 ( 
.A(n_157),
.Y(n_179)
);

INVx5_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_161),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_163),
.B(n_310),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_166),
.C(n_170),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_164),
.B(n_166),
.Y(n_215)
);

CKINVDCx16_ASAP7_75t_R g167 ( 
.A(n_168),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_SL g214 ( 
.A(n_170),
.B(n_215),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_175),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_171),
.B(n_175),
.Y(n_204)
);

INVxp33_ASAP7_75t_L g203 ( 
.A(n_172),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_176),
.A2(n_273),
.B1(n_275),
.B2(n_277),
.Y(n_272)
);

CKINVDCx14_ASAP7_75t_R g177 ( 
.A(n_178),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_186),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_183),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_182),
.B(n_183),
.C(n_186),
.Y(n_319)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

O2A1O1Ixp33_ASAP7_75t_SL g187 ( 
.A1(n_188),
.A2(n_219),
.B(n_307),
.C(n_312),
.Y(n_187)
);

AND2x2_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_213),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_189),
.B(n_213),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_204),
.C(n_205),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_190),
.A2(n_191),
.B1(n_303),
.B2(n_304),
.Y(n_302)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_200),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_193),
.A2(n_194),
.B1(n_196),
.B2(n_197),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_194),
.B(n_196),
.C(n_200),
.Y(n_218)
);

CKINVDCx16_ASAP7_75t_R g207 ( 
.A(n_195),
.Y(n_207)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_202),
.B(n_289),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_SL g304 ( 
.A(n_204),
.B(n_205),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_208),
.C(n_210),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_206),
.B(n_243),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_208),
.A2(n_209),
.B1(n_210),
.B2(n_244),
.Y(n_243)
);

CKINVDCx16_ASAP7_75t_R g208 ( 
.A(n_209),
.Y(n_208)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_210),
.Y(n_244)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_211),
.Y(n_229)
);

BUFx2_ASAP7_75t_L g276 ( 
.A(n_212),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_216),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_214),
.B(n_217),
.C(n_218),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_218),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_221),
.Y(n_219)
);

AOI21xp5_ASAP7_75t_SL g221 ( 
.A1(n_222),
.A2(n_301),
.B(n_306),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_L g222 ( 
.A1(n_223),
.A2(n_251),
.B(n_300),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_240),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_224),
.B(n_240),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_233),
.C(n_237),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_225),
.B(n_296),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_SL g225 ( 
.A(n_226),
.B(n_228),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_226),
.B(n_228),
.Y(n_247)
);

AOI21xp5_ASAP7_75t_L g228 ( 
.A1(n_229),
.A2(n_230),
.B(n_231),
.Y(n_228)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_230),
.Y(n_289)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_231),
.Y(n_285)
);

INVxp67_ASAP7_75t_L g263 ( 
.A(n_232),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_233),
.A2(n_237),
.B1(n_238),
.B2(n_297),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_233),
.Y(n_297)
);

INVxp67_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_236),
.Y(n_249)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_241),
.A2(n_242),
.B1(n_245),
.B2(n_246),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_241),
.B(n_247),
.C(n_248),
.Y(n_305)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_248),
.Y(n_246)
);

AOI21xp5_ASAP7_75t_L g251 ( 
.A1(n_252),
.A2(n_294),
.B(n_299),
.Y(n_251)
);

OAI21xp5_ASAP7_75t_SL g252 ( 
.A1(n_253),
.A2(n_270),
.B(n_293),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_SL g253 ( 
.A(n_254),
.B(n_264),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_254),
.B(n_264),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_260),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_256),
.A2(n_257),
.B1(n_258),
.B2(n_259),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_256),
.B(n_259),
.C(n_260),
.Y(n_298)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

INVxp67_ASAP7_75t_L g277 ( 
.A(n_261),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_SL g264 ( 
.A(n_265),
.B(n_268),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_265),
.A2(n_266),
.B1(n_268),
.B2(n_279),
.Y(n_278)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_268),
.Y(n_279)
);

AOI21xp5_ASAP7_75t_L g270 ( 
.A1(n_271),
.A2(n_280),
.B(n_292),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_278),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_272),
.B(n_278),
.Y(n_292)
);

INVxp67_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

OAI21xp5_ASAP7_75t_L g283 ( 
.A1(n_274),
.A2(n_284),
.B(n_285),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_276),
.Y(n_275)
);

OAI21xp5_ASAP7_75t_SL g280 ( 
.A1(n_281),
.A2(n_286),
.B(n_291),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_282),
.B(n_283),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_282),
.B(n_283),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_287),
.B(n_290),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_295),
.B(n_298),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_295),
.B(n_298),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_SL g301 ( 
.A(n_302),
.B(n_305),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_302),
.B(n_305),
.Y(n_306)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_308),
.B(n_309),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_308),
.B(n_309),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_SL g314 ( 
.A(n_315),
.B(n_319),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_315),
.B(n_319),
.Y(n_320)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_316),
.Y(n_318)
);


endmodule