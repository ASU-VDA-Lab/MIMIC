module fake_jpeg_1685_n_152 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_152);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_152;

wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_73;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_15;
wire n_124;
wire n_141;
wire n_57;
wire n_21;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_6),
.Y(n_15)
);

INVx2_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_12),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_0),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_3),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_3),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_10),
.Y(n_26)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_10),
.Y(n_30)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_31),
.Y(n_52)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_28),
.Y(n_32)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_32),
.Y(n_51)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_33),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_18),
.B(n_0),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_SL g41 ( 
.A(n_34),
.B(n_39),
.Y(n_41)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_18),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

INVxp33_ASAP7_75t_L g42 ( 
.A(n_37),
.Y(n_42)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_27),
.Y(n_38)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_15),
.Y(n_39)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_27),
.Y(n_40)
);

BUFx10_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

OR2x2_ASAP7_75t_L g43 ( 
.A(n_32),
.B(n_37),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_43),
.B(n_45),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_39),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_40),
.B(n_29),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_46),
.B(n_47),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_34),
.B(n_29),
.Y(n_47)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_48),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_33),
.B(n_24),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_49),
.B(n_20),
.Y(n_57)
);

NAND3xp33_ASAP7_75t_L g50 ( 
.A(n_38),
.B(n_15),
.C(n_26),
.Y(n_50)
);

INVxp67_ASAP7_75t_L g59 ( 
.A(n_50),
.Y(n_59)
);

OAI21xp33_ASAP7_75t_L g91 ( 
.A1(n_57),
.A2(n_58),
.B(n_70),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_43),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_52),
.Y(n_60)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_60),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_49),
.B(n_31),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_62),
.B(n_74),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_L g65 ( 
.A1(n_41),
.A2(n_20),
.B(n_25),
.Y(n_65)
);

AOI21xp5_ASAP7_75t_L g92 ( 
.A1(n_65),
.A2(n_19),
.B(n_22),
.Y(n_92)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_52),
.Y(n_66)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_66),
.Y(n_86)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_51),
.Y(n_67)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_67),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_51),
.A2(n_21),
.B1(n_25),
.B2(n_30),
.Y(n_68)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_68),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_56),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_69),
.B(n_72),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_56),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_55),
.A2(n_35),
.B1(n_36),
.B2(n_21),
.Y(n_71)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_71),
.B(n_73),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_44),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_55),
.A2(n_24),
.B1(n_23),
.B2(n_22),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_42),
.B(n_23),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_42),
.Y(n_75)
);

INVxp33_ASAP7_75t_L g77 ( 
.A(n_75),
.Y(n_77)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_44),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_76),
.B(n_75),
.Y(n_83)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_83),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_62),
.B(n_48),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_84),
.B(n_85),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_57),
.B(n_53),
.Y(n_85)
);

CKINVDCx16_ASAP7_75t_R g88 ( 
.A(n_61),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_88),
.B(n_89),
.Y(n_95)
);

A2O1A1Ixp33_ASAP7_75t_L g89 ( 
.A1(n_58),
.A2(n_30),
.B(n_26),
.C(n_19),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_74),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_90),
.B(n_59),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_92),
.B(n_0),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_67),
.B(n_17),
.C(n_54),
.Y(n_93)
);

XNOR2xp5_ASAP7_75t_L g101 ( 
.A(n_93),
.B(n_76),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_84),
.A2(n_65),
.B1(n_63),
.B2(n_59),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_94),
.A2(n_105),
.B1(n_87),
.B2(n_79),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_97),
.B(n_98),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_83),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_91),
.B(n_17),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_99),
.B(n_106),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_80),
.Y(n_100)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_100),
.Y(n_109)
);

XOR2xp5_ASAP7_75t_L g120 ( 
.A(n_101),
.B(n_79),
.Y(n_120)
);

OAI21xp33_ASAP7_75t_L g103 ( 
.A1(n_82),
.A2(n_70),
.B(n_1),
.Y(n_103)
);

INVx1_ASAP7_75t_SL g116 ( 
.A(n_103),
.Y(n_116)
);

OAI32xp33_ASAP7_75t_L g104 ( 
.A1(n_82),
.A2(n_64),
.A3(n_54),
.B1(n_60),
.B2(n_66),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_104),
.B(n_93),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_85),
.A2(n_64),
.B1(n_53),
.B2(n_54),
.Y(n_105)
);

NOR4xp25_ASAP7_75t_L g106 ( 
.A(n_89),
.B(n_8),
.C(n_14),
.D(n_13),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_107),
.B(n_92),
.Y(n_118)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_81),
.Y(n_108)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_108),
.Y(n_113)
);

CKINVDCx16_ASAP7_75t_R g110 ( 
.A(n_95),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_110),
.B(n_94),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_111),
.A2(n_87),
.B1(n_105),
.B2(n_81),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_101),
.B(n_96),
.C(n_102),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_112),
.B(n_77),
.C(n_78),
.Y(n_126)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_114),
.Y(n_125)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_100),
.Y(n_115)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_115),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_118),
.B(n_86),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_SL g129 ( 
.A(n_120),
.B(n_54),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_121),
.B(n_122),
.Y(n_130)
);

AOI31xp33_ASAP7_75t_L g122 ( 
.A1(n_119),
.A2(n_103),
.A3(n_104),
.B(n_79),
.Y(n_122)
);

XNOR2xp5_ASAP7_75t_L g135 ( 
.A(n_124),
.B(n_126),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_127),
.B(n_116),
.Y(n_133)
);

AOI21xp5_ASAP7_75t_L g128 ( 
.A1(n_111),
.A2(n_86),
.B(n_78),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_L g136 ( 
.A1(n_128),
.A2(n_1),
.B1(n_4),
.B2(n_6),
.Y(n_136)
);

AOI321xp33_ASAP7_75t_L g132 ( 
.A1(n_129),
.A2(n_109),
.A3(n_113),
.B1(n_112),
.B2(n_116),
.C(n_117),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_125),
.A2(n_114),
.B1(n_120),
.B2(n_109),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_131),
.B(n_132),
.Y(n_140)
);

OR2x2_ASAP7_75t_L g137 ( 
.A(n_133),
.B(n_136),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_125),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_134)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_134),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_135),
.B(n_126),
.C(n_123),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_139),
.B(n_141),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_135),
.B(n_128),
.C(n_129),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_137),
.B(n_134),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_143),
.A2(n_144),
.B1(n_13),
.B2(n_14),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_138),
.B(n_131),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_140),
.A2(n_124),
.B1(n_130),
.B2(n_11),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_145),
.A2(n_7),
.B1(n_9),
.B2(n_11),
.Y(n_147)
);

BUFx24_ASAP7_75t_SL g146 ( 
.A(n_145),
.Y(n_146)
);

INVxp67_ASAP7_75t_L g150 ( 
.A(n_146),
.Y(n_150)
);

HB1xp67_ASAP7_75t_L g149 ( 
.A(n_147),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_150),
.B(n_142),
.C(n_148),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_151),
.B(n_149),
.Y(n_152)
);


endmodule