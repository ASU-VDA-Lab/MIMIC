module real_aes_4300_n_267 (n_17, n_28, n_226, n_76, n_202, n_255, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_257, n_261, n_262, n_238, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_263, n_230, n_165, n_51, n_195, n_246, n_248, n_252, n_176, n_27, n_163, n_222, n_249, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_254, n_18, n_207, n_104, n_21, n_31, n_8, n_251, n_183, n_266, n_205, n_220, n_211, n_10, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_234, n_153, n_75, n_178, n_219, n_256, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_239, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_253, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_95, n_131, n_144, n_164, n_231, n_169, n_242, n_44, n_102, n_188, n_152, n_198, n_201, n_122, n_7, n_228, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_69, n_46, n_109, n_59, n_25, n_203, n_236, n_73, n_77, n_218, n_81, n_133, n_48, n_260, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_138, n_50, n_114, n_89, n_170, n_26, n_235, n_265, n_86, n_93, n_182, n_154, n_127, n_199, n_245, n_161, n_189, n_13, n_24, n_217, n_2, n_142, n_55, n_168, n_175, n_241, n_145, n_62, n_105, n_223, n_84, n_227, n_67, n_92, n_33, n_206, n_258, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_250, n_116, n_94, n_229, n_39, n_5, n_45, n_60, n_233, n_240, n_247, n_38, n_259, n_155, n_243, n_118, n_143, n_139, n_244, n_192, n_213, n_136, n_87, n_171, n_0, n_157, n_78, n_264, n_101, n_63, n_1, n_146, n_237, n_107, n_184, n_53, n_36, n_267);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_255;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_257;
input n_261;
input n_262;
input n_238;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_263;
input n_230;
input n_165;
input n_51;
input n_195;
input n_246;
input n_248;
input n_252;
input n_176;
input n_27;
input n_163;
input n_222;
input n_249;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_254;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_251;
input n_183;
input n_266;
input n_205;
input n_220;
input n_211;
input n_10;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_234;
input n_153;
input n_75;
input n_178;
input n_219;
input n_256;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_239;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_253;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_242;
input n_44;
input n_102;
input n_188;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_69;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_236;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_260;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_138;
input n_50;
input n_114;
input n_89;
input n_170;
input n_26;
input n_235;
input n_265;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_245;
input n_161;
input n_189;
input n_13;
input n_24;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_241;
input n_145;
input n_62;
input n_105;
input n_223;
input n_84;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_258;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_250;
input n_116;
input n_94;
input n_229;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_240;
input n_247;
input n_38;
input n_259;
input n_155;
input n_243;
input n_118;
input n_143;
input n_139;
input n_244;
input n_192;
input n_213;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_264;
input n_101;
input n_63;
input n_1;
input n_146;
input n_237;
input n_107;
input n_184;
input n_53;
input n_36;
output n_267;
wire n_480;
wire n_476;
wire n_758;
wire n_599;
wire n_436;
wire n_887;
wire n_684;
wire n_390;
wire n_821;
wire n_830;
wire n_285;
wire n_624;
wire n_980;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_838;
wire n_933;
wire n_485;
wire n_822;
wire n_846;
wire n_750;
wire n_631;
wire n_943;
wire n_977;
wire n_357;
wire n_287;
wire n_503;
wire n_635;
wire n_673;
wire n_386;
wire n_792;
wire n_518;
wire n_905;
wire n_878;
wire n_665;
wire n_667;
wire n_991;
wire n_1004;
wire n_577;
wire n_580;
wire n_469;
wire n_987;
wire n_362;
wire n_759;
wire n_979;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_900;
wire n_328;
wire n_718;
wire n_318;
wire n_841;
wire n_355;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_364;
wire n_421;
wire n_319;
wire n_555;
wire n_329;
wire n_766;
wire n_852;
wire n_974;
wire n_919;
wire n_857;
wire n_461;
wire n_908;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_923;
wire n_894;
wire n_952;
wire n_429;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_460;
wire n_937;
wire n_773;
wire n_989;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_963;
wire n_865;
wire n_537;
wire n_551;
wire n_666;
wire n_320;
wire n_884;
wire n_560;
wire n_660;
wire n_814;
wire n_944;
wire n_886;
wire n_594;
wire n_856;
wire n_983;
wire n_767;
wire n_696;
wire n_889;
wire n_955;
wire n_975;
wire n_704;
wire n_941;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_932;
wire n_399;
wire n_948;
wire n_700;
wire n_677;
wire n_958;
wire n_378;
wire n_591;
wire n_775;
wire n_763;
wire n_961;
wire n_870;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_415;
wire n_572;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_625;
wire n_953;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_990;
wire n_550;
wire n_966;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_918;
wire n_356;
wire n_478;
wire n_883;
wire n_584;
wire n_896;
wire n_408;
wire n_553;
wire n_372;
wire n_994;
wire n_528;
wire n_578;
wire n_495;
wire n_892;
wire n_370;
wire n_744;
wire n_384;
wire n_938;
wire n_352;
wire n_935;
wire n_824;
wire n_467;
wire n_951;
wire n_875;
wire n_327;
wire n_774;
wire n_992;
wire n_813;
wire n_981;
wire n_791;
wire n_466;
wire n_559;
wire n_976;
wire n_636;
wire n_872;
wire n_906;
wire n_477;
wire n_515;
wire n_984;
wire n_680;
wire n_595;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_931;
wire n_780;
wire n_904;
wire n_570;
wire n_675;
wire n_840;
wire n_920;
wire n_530;
wire n_835;
wire n_535;
wire n_732;
wire n_834;
wire n_882;
wire n_784;
wire n_281;
wire n_496;
wire n_962;
wire n_693;
wire n_468;
wire n_746;
wire n_284;
wire n_532;
wire n_316;
wire n_656;
wire n_755;
wire n_409;
wire n_748;
wire n_781;
wire n_860;
wire n_996;
wire n_298;
wire n_523;
wire n_909;
wire n_439;
wire n_576;
wire n_924;
wire n_956;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_874;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_310;
wire n_455;
wire n_973;
wire n_725;
wire n_504;
wire n_671;
wire n_960;
wire n_659;
wire n_547;
wire n_634;
wire n_682;
wire n_903;
wire n_454;
wire n_812;
wire n_782;
wire n_443;
wire n_565;
wire n_817;
wire n_760;
wire n_608;
wire n_925;
wire n_534;
wire n_708;
wire n_457;
wire n_345;
wire n_304;
wire n_885;
wire n_950;
wire n_381;
wire n_993;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_664;
wire n_367;
wire n_819;
wire n_737;
wire n_581;
wire n_610;
wire n_936;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_940;
wire n_722;
wire n_745;
wire n_867;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_879;
wire n_331;
wire n_417;
wire n_363;
wire n_754;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_901;
wire n_561;
wire n_947;
wire n_970;
wire n_876;
wire n_437;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_672;
wire n_567;
wire n_916;
wire n_406;
wire n_426;
wire n_617;
wire n_402;
wire n_552;
wire n_602;
wire n_733;
wire n_658;
wire n_676;
wire n_986;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_880;
wire n_807;
wire n_286;
wire n_416;
wire n_790;
wire n_895;
wire n_832;
wire n_410;
wire n_799;
wire n_805;
wire n_751;
wire n_999;
wire n_490;
wire n_913;
wire n_619;
wire n_391;
wire n_360;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_361;
wire n_917;
wire n_632;
wire n_768;
wire n_412;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_985;
wire n_488;
wire n_501;
wire n_910;
wire n_642;
wire n_613;
wire n_869;
wire n_387;
wire n_957;
wire n_995;
wire n_296;
wire n_702;
wire n_954;
wire n_969;
wire n_912;
wire n_302;
wire n_464;
wire n_351;
wire n_945;
wire n_604;
wire n_734;
wire n_898;
wire n_848;
wire n_392;
wire n_562;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_997;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_891;
wire n_269;
wire n_430;
wire n_568;
wire n_413;
wire n_471;
wire n_902;
wire n_853;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_699;
wire n_533;
wire n_1000;
wire n_1003;
wire n_366;
wire n_346;
wire n_727;
wire n_397;
wire n_293;
wire n_749;
wire n_358;
wire n_275;
wire n_385;
wire n_649;
wire n_663;
wire n_588;
wire n_536;
wire n_914;
wire n_707;
wire n_622;
wire n_470;
wire n_915;
wire n_851;
wire n_1002;
wire n_934;
wire n_494;
wire n_1001;
wire n_711;
wire n_864;
wire n_377;
wire n_273;
wire n_927;
wire n_965;
wire n_723;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_845;
wire n_850;
wire n_720;
wire n_354;
wire n_972;
wire n_435;
wire n_511;
wire n_484;
wire n_326;
wire n_893;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_930;
wire n_411;
wire n_697;
wire n_291;
wire n_978;
wire n_847;
wire n_907;
wire n_779;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_826;
wire n_648;
wire n_373;
wire n_589;
wire n_628;
wire n_939;
wire n_487;
wire n_831;
wire n_290;
wire n_365;
wire n_653;
wire n_637;
wire n_526;
wire n_928;
wire n_899;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_922;
wire n_926;
wire n_942;
wire n_472;
wire n_971;
wire n_866;
wire n_452;
wire n_787;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_959;
wire n_946;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_858;
wire n_873;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_623;
wire n_446;
wire n_721;
wire n_681;
wire n_982;
wire n_456;
wire n_717;
wire n_359;
wire n_312;
wire n_712;
wire n_433;
wire n_335;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_524;
wire n_861;
wire n_705;
wire n_762;
wire n_325;
wire n_575;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_541;
wire n_839;
wire n_639;
wire n_546;
wire n_587;
wire n_811;
wire n_459;
wire n_558;
wire n_863;
wire n_998;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_888;
wire n_836;
wire n_793;
wire n_272;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_929;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_890;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_949;
wire n_614;
wire n_305;
wire n_586;
wire n_911;
wire n_772;
wire n_450;
wire n_788;
wire n_441;
wire n_585;
wire n_719;
wire n_473;
wire n_465;
wire n_566;
wire n_967;
wire n_837;
wire n_871;
wire n_474;
wire n_829;
wire n_988;
wire n_921;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_687;
wire n_729;
wire n_844;
wire n_968;
wire n_710;
wire n_646;
wire n_650;
wire n_743;
wire n_393;
wire n_294;
wire n_652;
wire n_703;
wire n_823;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_854;
wire n_424;
wire n_877;
wire n_802;
wire n_868;
wire n_574;
wire n_337;
wire n_842;
wire n_849;
wire n_475;
wire n_554;
wire n_897;
wire n_855;
wire n_798;
wire n_668;
wire n_797;
wire n_862;
AOI22xp33_ASAP7_75t_L g503 ( .A1(n_0), .A2(n_111), .B1(n_418), .B2(n_456), .Y(n_503) );
HB1xp67_ASAP7_75t_L g278 ( .A(n_1), .Y(n_278) );
AND2x4_ASAP7_75t_L g747 ( .A(n_1), .B(n_748), .Y(n_747) );
AND2x4_ASAP7_75t_L g753 ( .A(n_1), .B(n_258), .Y(n_753) );
AOI22xp33_ASAP7_75t_L g499 ( .A1(n_2), .A2(n_217), .B1(n_451), .B2(n_454), .Y(n_499) );
AO22x1_ASAP7_75t_L g751 ( .A1(n_3), .A2(n_5), .B1(n_752), .B2(n_754), .Y(n_751) );
INVx1_ASAP7_75t_L g405 ( .A(n_4), .Y(n_405) );
AOI22xp33_ASAP7_75t_L g776 ( .A1(n_6), .A2(n_199), .B1(n_744), .B2(n_759), .Y(n_776) );
AOI22xp33_ASAP7_75t_L g510 ( .A1(n_7), .A2(n_58), .B1(n_425), .B2(n_511), .Y(n_510) );
AOI22xp5_ASAP7_75t_L g436 ( .A1(n_8), .A2(n_34), .B1(n_437), .B2(n_439), .Y(n_436) );
AOI22xp33_ASAP7_75t_L g705 ( .A1(n_9), .A2(n_266), .B1(n_402), .B2(n_561), .Y(n_705) );
AOI22xp33_ASAP7_75t_L g719 ( .A1(n_10), .A2(n_22), .B1(n_334), .B2(n_537), .Y(n_719) );
AOI21xp33_ASAP7_75t_SL g638 ( .A1(n_11), .A2(n_511), .B(n_639), .Y(n_638) );
AOI21xp33_ASAP7_75t_L g475 ( .A1(n_12), .A2(n_476), .B(n_477), .Y(n_475) );
AOI22xp5_ASAP7_75t_L g730 ( .A1(n_13), .A2(n_109), .B1(n_357), .B2(n_581), .Y(n_730) );
AOI22xp33_ASAP7_75t_L g491 ( .A1(n_14), .A2(n_183), .B1(n_492), .B2(n_493), .Y(n_491) );
AOI22xp33_ASAP7_75t_L g501 ( .A1(n_15), .A2(n_121), .B1(n_453), .B2(n_502), .Y(n_501) );
AOI21xp5_ASAP7_75t_L g723 ( .A1(n_16), .A2(n_362), .B(n_724), .Y(n_723) );
AOI22xp33_ASAP7_75t_L g447 ( .A1(n_17), .A2(n_234), .B1(n_428), .B2(n_448), .Y(n_447) );
XOR2xp5_ASAP7_75t_L g395 ( .A(n_18), .B(n_396), .Y(n_395) );
AOI22xp33_ASAP7_75t_L g651 ( .A1(n_19), .A2(n_158), .B1(n_486), .B2(n_487), .Y(n_651) );
AOI22xp33_ASAP7_75t_L g352 ( .A1(n_20), .A2(n_137), .B1(n_353), .B2(n_357), .Y(n_352) );
AOI22xp33_ASAP7_75t_L g443 ( .A1(n_21), .A2(n_141), .B1(n_444), .B2(n_446), .Y(n_443) );
AO22x1_ASAP7_75t_L g967 ( .A1(n_23), .A2(n_25), .B1(n_968), .B2(n_969), .Y(n_967) );
AOI22xp5_ASAP7_75t_L g760 ( .A1(n_24), .A2(n_122), .B1(n_761), .B2(n_762), .Y(n_760) );
INVx1_ASAP7_75t_L g975 ( .A(n_26), .Y(n_975) );
AOI22xp33_ASAP7_75t_L g726 ( .A1(n_27), .A2(n_205), .B1(n_727), .B2(n_728), .Y(n_726) );
AOI221xp5_ASAP7_75t_L g505 ( .A1(n_28), .A2(n_48), .B1(n_506), .B2(n_507), .C(n_508), .Y(n_505) );
INVx1_ASAP7_75t_SL g586 ( .A(n_29), .Y(n_586) );
INVx1_ASAP7_75t_L g988 ( .A(n_30), .Y(n_988) );
INVx1_ASAP7_75t_L g509 ( .A(n_31), .Y(n_509) );
AOI22xp33_ASAP7_75t_L g534 ( .A1(n_32), .A2(n_178), .B1(n_535), .B2(n_537), .Y(n_534) );
AOI22xp33_ASAP7_75t_L g972 ( .A1(n_33), .A2(n_40), .B1(n_539), .B2(n_973), .Y(n_972) );
NOR2xp33_ASAP7_75t_L g276 ( .A(n_35), .B(n_202), .Y(n_276) );
INVx1_ASAP7_75t_L g312 ( .A(n_35), .Y(n_312) );
INVxp67_ASAP7_75t_L g383 ( .A(n_35), .Y(n_383) );
OA22x2_ASAP7_75t_L g647 ( .A1(n_36), .A2(n_648), .B1(n_659), .B2(n_660), .Y(n_647) );
INVx1_ASAP7_75t_L g660 ( .A(n_36), .Y(n_660) );
AOI22xp5_ASAP7_75t_L g702 ( .A1(n_37), .A2(n_204), .B1(n_472), .B2(n_632), .Y(n_702) );
AOI22xp33_ASAP7_75t_L g344 ( .A1(n_38), .A2(n_52), .B1(n_345), .B2(n_347), .Y(n_344) );
INVx1_ASAP7_75t_L g571 ( .A(n_39), .Y(n_571) );
AOI22xp33_ASAP7_75t_L g485 ( .A1(n_41), .A2(n_55), .B1(n_486), .B2(n_487), .Y(n_485) );
NAND2xp5_ASAP7_75t_L g440 ( .A(n_42), .B(n_441), .Y(n_440) );
XOR2xp5_ASAP7_75t_L g998 ( .A(n_43), .B(n_999), .Y(n_998) );
AOI22xp5_ASAP7_75t_L g682 ( .A1(n_44), .A2(n_97), .B1(n_290), .B2(n_683), .Y(n_682) );
NAND2xp5_ASAP7_75t_SL g308 ( .A(n_45), .B(n_296), .Y(n_308) );
AOI22xp33_ASAP7_75t_L g359 ( .A1(n_46), .A2(n_105), .B1(n_360), .B2(n_364), .Y(n_359) );
AOI22xp33_ASAP7_75t_L g681 ( .A1(n_47), .A2(n_230), .B1(n_334), .B2(n_537), .Y(n_681) );
INVx1_ASAP7_75t_SL g575 ( .A(n_49), .Y(n_575) );
AOI22xp33_ASAP7_75t_L g547 ( .A1(n_50), .A2(n_257), .B1(n_428), .B2(n_448), .Y(n_547) );
AOI22xp33_ASAP7_75t_L g452 ( .A1(n_51), .A2(n_227), .B1(n_453), .B2(n_454), .Y(n_452) );
INVx1_ASAP7_75t_L g640 ( .A(n_53), .Y(n_640) );
AOI22xp5_ASAP7_75t_L g668 ( .A1(n_54), .A2(n_93), .B1(n_511), .B2(n_669), .Y(n_668) );
INVx1_ASAP7_75t_L g986 ( .A(n_56), .Y(n_986) );
AOI22xp5_ASAP7_75t_L g785 ( .A1(n_57), .A2(n_171), .B1(n_754), .B2(n_770), .Y(n_785) );
AOI22xp5_ASAP7_75t_L g416 ( .A1(n_59), .A2(n_246), .B1(n_417), .B2(n_418), .Y(n_416) );
INVx1_ASAP7_75t_SL g583 ( .A(n_60), .Y(n_583) );
INVx2_ASAP7_75t_L g273 ( .A(n_61), .Y(n_273) );
AOI22xp33_ASAP7_75t_L g627 ( .A1(n_62), .A2(n_119), .B1(n_399), .B2(n_628), .Y(n_627) );
AOI22xp33_ASAP7_75t_L g401 ( .A1(n_63), .A2(n_131), .B1(n_290), .B2(n_402), .Y(n_401) );
INVx1_ASAP7_75t_L g746 ( .A(n_64), .Y(n_746) );
AND2x4_ASAP7_75t_L g750 ( .A(n_64), .B(n_273), .Y(n_750) );
INVx1_ASAP7_75t_SL g758 ( .A(n_64), .Y(n_758) );
INVx1_ASAP7_75t_SL g579 ( .A(n_65), .Y(n_579) );
AOI22xp5_ASAP7_75t_L g596 ( .A1(n_66), .A2(n_75), .B1(n_597), .B2(n_600), .Y(n_596) );
AOI22xp33_ASAP7_75t_L g849 ( .A1(n_67), .A2(n_187), .B1(n_752), .B2(n_771), .Y(n_849) );
AOI22xp33_ASAP7_75t_L g538 ( .A1(n_68), .A2(n_194), .B1(n_347), .B2(n_539), .Y(n_538) );
INVx1_ASAP7_75t_L g990 ( .A(n_69), .Y(n_990) );
INVx1_ASAP7_75t_L g552 ( .A(n_70), .Y(n_552) );
AOI22xp5_ASAP7_75t_L g670 ( .A1(n_71), .A2(n_181), .B1(n_671), .B2(n_673), .Y(n_670) );
INVx1_ASAP7_75t_L g433 ( .A(n_72), .Y(n_433) );
AOI22xp33_ASAP7_75t_L g711 ( .A1(n_73), .A2(n_238), .B1(n_417), .B2(n_418), .Y(n_711) );
BUFx6f_ASAP7_75t_L g296 ( .A(n_74), .Y(n_296) );
AOI22xp33_ASAP7_75t_L g455 ( .A1(n_76), .A2(n_190), .B1(n_418), .B2(n_456), .Y(n_455) );
AOI22xp5_ASAP7_75t_L g555 ( .A1(n_77), .A2(n_262), .B1(n_400), .B2(n_402), .Y(n_555) );
INVx1_ASAP7_75t_L g982 ( .A(n_78), .Y(n_982) );
INVx1_ASAP7_75t_L g667 ( .A(n_79), .Y(n_667) );
AOI22xp5_ASAP7_75t_L g790 ( .A1(n_80), .A2(n_162), .B1(n_744), .B2(n_749), .Y(n_790) );
AOI22xp5_ASAP7_75t_L g450 ( .A1(n_81), .A2(n_165), .B1(n_330), .B2(n_451), .Y(n_450) );
AOI22xp33_ASAP7_75t_L g541 ( .A1(n_82), .A2(n_136), .B1(n_325), .B2(n_330), .Y(n_541) );
AOI22xp33_ASAP7_75t_L g775 ( .A1(n_83), .A2(n_197), .B1(n_754), .B2(n_770), .Y(n_775) );
AOI22xp33_ASAP7_75t_L g540 ( .A1(n_84), .A2(n_256), .B1(n_290), .B2(n_315), .Y(n_540) );
AOI22xp33_ASAP7_75t_L g636 ( .A1(n_85), .A2(n_231), .B1(n_429), .B2(n_637), .Y(n_636) );
INVx1_ASAP7_75t_L g297 ( .A(n_86), .Y(n_297) );
NAND2xp5_ASAP7_75t_L g380 ( .A(n_86), .B(n_201), .Y(n_380) );
AOI22xp33_ASAP7_75t_L g652 ( .A1(n_87), .A2(n_229), .B1(n_469), .B2(n_489), .Y(n_652) );
AOI22xp33_ASAP7_75t_L g779 ( .A1(n_88), .A2(n_176), .B1(n_752), .B2(n_754), .Y(n_779) );
INVx1_ASAP7_75t_L g412 ( .A(n_89), .Y(n_412) );
OAI22x1_ASAP7_75t_L g714 ( .A1(n_90), .A2(n_715), .B1(n_720), .B2(n_731), .Y(n_714) );
NAND5xp2_ASAP7_75t_SL g715 ( .A(n_90), .B(n_716), .C(n_717), .D(n_718), .E(n_719), .Y(n_715) );
AO22x1_ASAP7_75t_L g528 ( .A1(n_91), .A2(n_113), .B1(n_439), .B2(n_448), .Y(n_528) );
XNOR2x1_ASAP7_75t_L g465 ( .A(n_92), .B(n_466), .Y(n_465) );
AOI21xp5_ASAP7_75t_L g368 ( .A1(n_94), .A2(n_369), .B(n_373), .Y(n_368) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_95), .B(n_506), .Y(n_546) );
INVx1_ASAP7_75t_SL g607 ( .A(n_96), .Y(n_607) );
AOI22xp33_ASAP7_75t_L g625 ( .A1(n_98), .A2(n_214), .B1(n_417), .B2(n_418), .Y(n_625) );
AOI22xp33_ASAP7_75t_L g289 ( .A1(n_99), .A2(n_195), .B1(n_290), .B2(n_315), .Y(n_289) );
AOI22xp5_ASAP7_75t_L g593 ( .A1(n_100), .A2(n_228), .B1(n_347), .B2(n_594), .Y(n_593) );
AOI22xp5_ASAP7_75t_L g650 ( .A1(n_101), .A2(n_260), .B1(n_484), .B2(n_490), .Y(n_650) );
AOI22xp33_ASAP7_75t_L g703 ( .A1(n_102), .A2(n_147), .B1(n_473), .B2(n_483), .Y(n_703) );
AOI221xp5_ASAP7_75t_L g706 ( .A1(n_103), .A2(n_152), .B1(n_637), .B2(n_707), .C(n_709), .Y(n_706) );
AOI22xp33_ASAP7_75t_L g548 ( .A1(n_104), .A2(n_129), .B1(n_424), .B2(n_549), .Y(n_548) );
AOI221xp5_ASAP7_75t_SL g654 ( .A1(n_106), .A2(n_235), .B1(n_354), .B2(n_483), .C(n_655), .Y(n_654) );
AOI22xp33_ASAP7_75t_L g699 ( .A1(n_107), .A2(n_153), .B1(n_558), .B2(n_700), .Y(n_699) );
AOI22xp33_ASAP7_75t_L g780 ( .A1(n_108), .A2(n_117), .B1(n_744), .B2(n_759), .Y(n_780) );
AOI22xp33_ASAP7_75t_L g717 ( .A1(n_110), .A2(n_185), .B1(n_345), .B2(n_347), .Y(n_717) );
CKINVDCx5p33_ASAP7_75t_R g656 ( .A(n_112), .Y(n_656) );
AOI22xp33_ASAP7_75t_L g488 ( .A1(n_114), .A2(n_232), .B1(n_489), .B2(n_490), .Y(n_488) );
AOI221xp5_ASAP7_75t_L g657 ( .A1(n_115), .A2(n_180), .B1(n_470), .B2(n_472), .C(n_658), .Y(n_657) );
AOI21xp33_ASAP7_75t_L g550 ( .A1(n_116), .A2(n_371), .B(n_551), .Y(n_550) );
AOI22xp33_ASAP7_75t_L g846 ( .A1(n_118), .A2(n_203), .B1(n_767), .B2(n_847), .Y(n_846) );
AOI22xp33_ASAP7_75t_L g589 ( .A1(n_120), .A2(n_148), .B1(n_425), .B2(n_590), .Y(n_589) );
NAND2xp5_ASAP7_75t_L g474 ( .A(n_123), .B(n_354), .Y(n_474) );
AOI22xp33_ASAP7_75t_L g631 ( .A1(n_124), .A2(n_184), .B1(n_428), .B2(n_632), .Y(n_631) );
AOI22xp5_ASAP7_75t_L g786 ( .A1(n_125), .A2(n_247), .B1(n_744), .B2(n_759), .Y(n_786) );
AOI22xp5_ASAP7_75t_L g653 ( .A1(n_126), .A2(n_157), .B1(n_492), .B2(n_493), .Y(n_653) );
AOI22xp33_ASAP7_75t_L g677 ( .A1(n_127), .A2(n_160), .B1(n_330), .B2(n_399), .Y(n_677) );
INVx1_ASAP7_75t_L g478 ( .A(n_128), .Y(n_478) );
AOI22xp33_ASAP7_75t_L g716 ( .A1(n_130), .A2(n_237), .B1(n_290), .B2(n_315), .Y(n_716) );
INVx1_ASAP7_75t_L g384 ( .A(n_132), .Y(n_384) );
AOI22xp5_ASAP7_75t_L g718 ( .A1(n_133), .A2(n_218), .B1(n_325), .B2(n_330), .Y(n_718) );
AOI22xp33_ASAP7_75t_L g419 ( .A1(n_134), .A2(n_146), .B1(n_420), .B2(n_421), .Y(n_419) );
AOI22xp5_ASAP7_75t_L g512 ( .A1(n_135), .A2(n_193), .B1(n_446), .B2(n_513), .Y(n_512) );
AOI22xp33_ASAP7_75t_L g423 ( .A1(n_138), .A2(n_166), .B1(n_424), .B2(n_425), .Y(n_423) );
AOI22xp33_ASAP7_75t_L g482 ( .A1(n_139), .A2(n_245), .B1(n_483), .B2(n_484), .Y(n_482) );
AOI22xp5_ASAP7_75t_L g556 ( .A1(n_140), .A2(n_172), .B1(n_557), .B2(n_558), .Y(n_556) );
INVx1_ASAP7_75t_L g725 ( .A(n_142), .Y(n_725) );
AOI22xp33_ASAP7_75t_L g971 ( .A1(n_143), .A2(n_263), .B1(n_535), .B2(n_563), .Y(n_971) );
AOI22xp33_ASAP7_75t_L g471 ( .A1(n_144), .A2(n_210), .B1(n_472), .B2(n_473), .Y(n_471) );
INVx1_ASAP7_75t_L g981 ( .A(n_145), .Y(n_981) );
AOI22xp33_ASAP7_75t_SL g562 ( .A1(n_149), .A2(n_254), .B1(n_417), .B2(n_563), .Y(n_562) );
INVx1_ASAP7_75t_L g573 ( .A(n_150), .Y(n_573) );
AOI22xp5_ASAP7_75t_L g701 ( .A1(n_151), .A2(n_239), .B1(n_453), .B2(n_502), .Y(n_701) );
AOI22xp5_ASAP7_75t_L g756 ( .A1(n_154), .A2(n_243), .B1(n_757), .B2(n_759), .Y(n_756) );
AOI22xp33_ASAP7_75t_L g629 ( .A1(n_155), .A2(n_253), .B1(n_420), .B2(n_454), .Y(n_629) );
AO22x1_ASAP7_75t_L g658 ( .A1(n_156), .A2(n_226), .B1(n_473), .B2(n_476), .Y(n_658) );
AOI22xp33_ASAP7_75t_L g992 ( .A1(n_159), .A2(n_173), .B1(n_448), .B2(n_993), .Y(n_992) );
AOI22xp5_ASAP7_75t_L g560 ( .A1(n_161), .A2(n_255), .B1(n_420), .B2(n_561), .Y(n_560) );
XNOR2x1_ASAP7_75t_L g543 ( .A(n_162), .B(n_544), .Y(n_543) );
CKINVDCx20_ASAP7_75t_R g641 ( .A(n_163), .Y(n_641) );
INVxp67_ASAP7_75t_SL g285 ( .A(n_164), .Y(n_285) );
AOI22xp5_ASAP7_75t_L g791 ( .A1(n_167), .A2(n_207), .B1(n_762), .B2(n_770), .Y(n_791) );
AOI22xp5_ASAP7_75t_L g623 ( .A1(n_168), .A2(n_209), .B1(n_330), .B2(n_624), .Y(n_623) );
AOI22xp33_ASAP7_75t_L g766 ( .A1(n_169), .A2(n_200), .B1(n_744), .B2(n_767), .Y(n_766) );
AOI222xp33_ASAP7_75t_L g961 ( .A1(n_169), .A2(n_962), .B1(n_994), .B2(n_998), .C1(n_1000), .C2(n_1002), .Y(n_961) );
XOR2x2_ASAP7_75t_L g964 ( .A(n_169), .B(n_965), .Y(n_964) );
NAND2xp5_ASAP7_75t_L g385 ( .A(n_170), .B(n_386), .Y(n_385) );
AOI22xp33_ASAP7_75t_L g324 ( .A1(n_174), .A2(n_244), .B1(n_325), .B2(n_330), .Y(n_324) );
AO221x2_ASAP7_75t_L g743 ( .A1(n_175), .A2(n_223), .B1(n_744), .B2(n_749), .C(n_751), .Y(n_743) );
AOI22xp33_ASAP7_75t_L g468 ( .A1(n_177), .A2(n_211), .B1(n_469), .B2(n_470), .Y(n_468) );
AOI22xp33_ASAP7_75t_L g529 ( .A1(n_179), .A2(n_233), .B1(n_511), .B2(n_530), .Y(n_529) );
OA22x2_ASAP7_75t_L g302 ( .A1(n_182), .A2(n_202), .B1(n_296), .B2(n_300), .Y(n_302) );
INVx1_ASAP7_75t_L g321 ( .A(n_182), .Y(n_321) );
AOI22xp33_ASAP7_75t_L g427 ( .A1(n_186), .A2(n_212), .B1(n_428), .B2(n_429), .Y(n_427) );
AOI221x1_ASAP7_75t_L g664 ( .A1(n_188), .A2(n_222), .B1(n_581), .B2(n_665), .C(n_666), .Y(n_664) );
AOI22xp33_ASAP7_75t_L g500 ( .A1(n_189), .A2(n_240), .B1(n_330), .B2(n_399), .Y(n_500) );
AOI22xp33_ASAP7_75t_L g678 ( .A1(n_191), .A2(n_196), .B1(n_345), .B2(n_347), .Y(n_678) );
AOI22xp33_ASAP7_75t_L g769 ( .A1(n_192), .A2(n_251), .B1(n_770), .B2(n_771), .Y(n_769) );
AOI22xp33_ASAP7_75t_L g333 ( .A1(n_198), .A2(n_236), .B1(n_334), .B2(n_338), .Y(n_333) );
INVx1_ASAP7_75t_L g314 ( .A(n_201), .Y(n_314) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_201), .B(n_319), .Y(n_392) );
OAI21xp33_ASAP7_75t_L g322 ( .A1(n_202), .A2(n_213), .B(n_323), .Y(n_322) );
CKINVDCx20_ASAP7_75t_R g524 ( .A(n_203), .Y(n_524) );
AOI22xp33_ASAP7_75t_L g531 ( .A1(n_206), .A2(n_219), .B1(n_357), .B2(n_532), .Y(n_531) );
INVx1_ASAP7_75t_SL g614 ( .A(n_208), .Y(n_614) );
NOR2xp33_ASAP7_75t_L g277 ( .A(n_213), .B(n_249), .Y(n_277) );
INVx1_ASAP7_75t_L g299 ( .A(n_213), .Y(n_299) );
AOI21xp33_ASAP7_75t_L g410 ( .A1(n_215), .A2(n_354), .B(n_411), .Y(n_410) );
CKINVDCx5p33_ASAP7_75t_R g611 ( .A(n_216), .Y(n_611) );
INVx1_ASAP7_75t_L g710 ( .A(n_220), .Y(n_710) );
NAND2xp5_ASAP7_75t_L g633 ( .A(n_221), .B(n_634), .Y(n_633) );
OAI21x1_ASAP7_75t_L g661 ( .A1(n_224), .A2(n_662), .B(n_684), .Y(n_661) );
INVx1_ASAP7_75t_L g687 ( .A(n_224), .Y(n_687) );
XNOR2x1_ASAP7_75t_L g696 ( .A(n_225), .B(n_697), .Y(n_696) );
AOI22xp5_ASAP7_75t_L g458 ( .A1(n_241), .A2(n_252), .B1(n_399), .B2(n_459), .Y(n_458) );
INVx1_ASAP7_75t_SL g606 ( .A(n_242), .Y(n_606) );
INVx1_ASAP7_75t_L g978 ( .A(n_248), .Y(n_978) );
NAND2xp5_ASAP7_75t_L g306 ( .A(n_249), .B(n_307), .Y(n_306) );
AOI22xp33_ASAP7_75t_L g398 ( .A1(n_250), .A2(n_259), .B1(n_399), .B2(n_400), .Y(n_398) );
INVx1_ASAP7_75t_L g748 ( .A(n_258), .Y(n_748) );
NAND2xp5_ASAP7_75t_L g729 ( .A(n_261), .B(n_588), .Y(n_729) );
XNOR2x1_ASAP7_75t_L g496 ( .A(n_264), .B(n_497), .Y(n_496) );
AOI21xp5_ASAP7_75t_L g527 ( .A1(n_265), .A2(n_369), .B(n_528), .Y(n_527) );
AOI21xp5_ASAP7_75t_L g267 ( .A1(n_268), .A2(n_279), .B(n_737), .Y(n_267) );
INVx1_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
BUFx4_ASAP7_75t_SL g269 ( .A(n_270), .Y(n_269) );
NAND3xp33_ASAP7_75t_L g270 ( .A(n_271), .B(n_274), .C(n_278), .Y(n_270) );
AND2x2_ASAP7_75t_L g995 ( .A(n_271), .B(n_996), .Y(n_995) );
AND2x2_ASAP7_75t_L g1001 ( .A(n_271), .B(n_997), .Y(n_1001) );
INVx1_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
OA21x2_ASAP7_75t_L g1003 ( .A1(n_272), .A2(n_758), .B(n_1004), .Y(n_1003) );
HB1xp67_ASAP7_75t_L g272 ( .A(n_273), .Y(n_272) );
AND2x2_ASAP7_75t_L g745 ( .A(n_273), .B(n_746), .Y(n_745) );
AND3x4_ASAP7_75t_L g757 ( .A(n_273), .B(n_747), .C(n_758), .Y(n_757) );
NOR2xp33_ASAP7_75t_L g996 ( .A(n_274), .B(n_997), .Y(n_996) );
HB1xp67_ASAP7_75t_L g274 ( .A(n_275), .Y(n_274) );
AO21x2_ASAP7_75t_L g389 ( .A1(n_275), .A2(n_390), .B(n_391), .Y(n_389) );
NAND2xp5_ASAP7_75t_L g275 ( .A(n_276), .B(n_277), .Y(n_275) );
INVx1_ASAP7_75t_L g997 ( .A(n_278), .Y(n_997) );
XNOR2xp5_ASAP7_75t_L g279 ( .A(n_280), .B(n_518), .Y(n_279) );
HB1xp67_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
OAI22xp5_ASAP7_75t_L g281 ( .A1(n_282), .A2(n_283), .B1(n_462), .B2(n_463), .Y(n_281) );
INVx2_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
OA22x2_ASAP7_75t_L g283 ( .A1(n_284), .A2(n_394), .B1(n_460), .B2(n_461), .Y(n_283) );
INVx2_ASAP7_75t_L g461 ( .A(n_284), .Y(n_461) );
AO21x2_ASAP7_75t_L g284 ( .A1(n_285), .A2(n_286), .B(n_393), .Y(n_284) );
NOR3xp33_ASAP7_75t_L g393 ( .A(n_285), .B(n_288), .C(n_351), .Y(n_393) );
NAND2xp5_ASAP7_75t_L g286 ( .A(n_287), .B(n_350), .Y(n_286) );
INVx1_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
NAND4xp25_ASAP7_75t_SL g288 ( .A(n_289), .B(n_324), .C(n_333), .D(n_344), .Y(n_288) );
BUFx6f_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
BUFx6f_ASAP7_75t_L g454 ( .A(n_291), .Y(n_454) );
BUFx6f_ASAP7_75t_L g561 ( .A(n_291), .Y(n_561) );
BUFx6f_ASAP7_75t_L g599 ( .A(n_291), .Y(n_599) );
AND2x4_ASAP7_75t_L g291 ( .A(n_292), .B(n_303), .Y(n_291) );
AND2x4_ASAP7_75t_L g335 ( .A(n_292), .B(n_336), .Y(n_335) );
AND2x2_ASAP7_75t_L g341 ( .A(n_292), .B(n_342), .Y(n_341) );
AND2x4_ASAP7_75t_L g346 ( .A(n_292), .B(n_328), .Y(n_346) );
AND2x4_ASAP7_75t_L g469 ( .A(n_292), .B(n_332), .Y(n_469) );
AND2x4_ASAP7_75t_L g486 ( .A(n_292), .B(n_336), .Y(n_486) );
AND2x4_ASAP7_75t_L g487 ( .A(n_292), .B(n_342), .Y(n_487) );
AND2x4_ASAP7_75t_L g489 ( .A(n_292), .B(n_328), .Y(n_489) );
AND2x4_ASAP7_75t_L g292 ( .A(n_293), .B(n_301), .Y(n_292) );
AND2x2_ASAP7_75t_L g356 ( .A(n_293), .B(n_302), .Y(n_356) );
INVx1_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
AND2x2_ASAP7_75t_L g327 ( .A(n_294), .B(n_302), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g294 ( .A(n_295), .B(n_298), .Y(n_294) );
NAND2xp33_ASAP7_75t_L g295 ( .A(n_296), .B(n_297), .Y(n_295) );
INVx2_ASAP7_75t_L g300 ( .A(n_296), .Y(n_300) );
INVx3_ASAP7_75t_L g307 ( .A(n_296), .Y(n_307) );
NAND2xp33_ASAP7_75t_L g313 ( .A(n_296), .B(n_314), .Y(n_313) );
INVx1_ASAP7_75t_L g323 ( .A(n_296), .Y(n_323) );
HB1xp67_ASAP7_75t_L g379 ( .A(n_296), .Y(n_379) );
NAND2xp5_ASAP7_75t_L g320 ( .A(n_297), .B(n_321), .Y(n_320) );
NAND2xp5_ASAP7_75t_L g298 ( .A(n_299), .B(n_300), .Y(n_298) );
OAI21xp5_ASAP7_75t_L g382 ( .A1(n_299), .A2(n_323), .B(n_383), .Y(n_382) );
INVx1_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
AND2x2_ASAP7_75t_L g381 ( .A(n_302), .B(n_382), .Y(n_381) );
AND2x4_ASAP7_75t_L g316 ( .A(n_303), .B(n_317), .Y(n_316) );
AND2x4_ASAP7_75t_L g490 ( .A(n_303), .B(n_327), .Y(n_490) );
AND2x4_ASAP7_75t_L g493 ( .A(n_303), .B(n_317), .Y(n_493) );
INVx2_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
INVx2_ASAP7_75t_L g332 ( .A(n_304), .Y(n_332) );
OR2x2_ASAP7_75t_L g304 ( .A(n_305), .B(n_309), .Y(n_304) );
AND2x4_ASAP7_75t_L g328 ( .A(n_305), .B(n_329), .Y(n_328) );
AND2x4_ASAP7_75t_L g336 ( .A(n_305), .B(n_337), .Y(n_336) );
INVx2_ASAP7_75t_L g343 ( .A(n_305), .Y(n_343) );
AND2x2_ASAP7_75t_L g377 ( .A(n_305), .B(n_378), .Y(n_377) );
AND2x4_ASAP7_75t_L g305 ( .A(n_306), .B(n_308), .Y(n_305) );
NAND2xp5_ASAP7_75t_L g311 ( .A(n_307), .B(n_312), .Y(n_311) );
INVxp67_ASAP7_75t_L g319 ( .A(n_307), .Y(n_319) );
NAND3xp33_ASAP7_75t_L g391 ( .A(n_308), .B(n_318), .C(n_392), .Y(n_391) );
INVx1_ASAP7_75t_L g329 ( .A(n_309), .Y(n_329) );
INVx1_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
INVx1_ASAP7_75t_L g337 ( .A(n_310), .Y(n_337) );
AND2x2_ASAP7_75t_L g310 ( .A(n_311), .B(n_313), .Y(n_310) );
BUFx12f_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
INVx6_ASAP7_75t_L g403 ( .A(n_316), .Y(n_403) );
AND2x4_ASAP7_75t_L g349 ( .A(n_317), .B(n_328), .Y(n_349) );
AND2x4_ASAP7_75t_L g358 ( .A(n_317), .B(n_342), .Y(n_358) );
AND2x4_ASAP7_75t_L g473 ( .A(n_317), .B(n_342), .Y(n_473) );
AND2x4_ASAP7_75t_L g492 ( .A(n_317), .B(n_328), .Y(n_492) );
AND2x2_ASAP7_75t_L g317 ( .A(n_318), .B(n_322), .Y(n_317) );
NAND2xp5_ASAP7_75t_L g318 ( .A(n_319), .B(n_320), .Y(n_318) );
BUFx8_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
BUFx6f_ASAP7_75t_L g399 ( .A(n_326), .Y(n_399) );
AND2x2_ASAP7_75t_L g326 ( .A(n_327), .B(n_328), .Y(n_326) );
AND2x4_ASAP7_75t_L g331 ( .A(n_327), .B(n_332), .Y(n_331) );
AND2x2_ASAP7_75t_L g367 ( .A(n_327), .B(n_336), .Y(n_367) );
AND2x2_ASAP7_75t_L g372 ( .A(n_327), .B(n_342), .Y(n_372) );
AND2x4_ASAP7_75t_L g472 ( .A(n_327), .B(n_336), .Y(n_472) );
AND2x2_ASAP7_75t_L g476 ( .A(n_327), .B(n_342), .Y(n_476) );
AND2x4_ASAP7_75t_L g484 ( .A(n_327), .B(n_328), .Y(n_484) );
AND2x2_ASAP7_75t_L g559 ( .A(n_327), .B(n_328), .Y(n_559) );
BUFx6f_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
BUFx12f_ASAP7_75t_L g400 ( .A(n_331), .Y(n_400) );
BUFx3_ASAP7_75t_L g609 ( .A(n_331), .Y(n_609) );
BUFx6f_ASAP7_75t_L g700 ( .A(n_331), .Y(n_700) );
BUFx6f_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
BUFx12f_ASAP7_75t_L g417 ( .A(n_335), .Y(n_417) );
INVx3_ASAP7_75t_L g457 ( .A(n_335), .Y(n_457) );
AND2x4_ASAP7_75t_L g363 ( .A(n_336), .B(n_356), .Y(n_363) );
AND2x4_ASAP7_75t_L g483 ( .A(n_336), .B(n_356), .Y(n_483) );
AND2x4_ASAP7_75t_L g342 ( .A(n_337), .B(n_343), .Y(n_342) );
BUFx6f_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
INVx2_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
INVx1_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
BUFx6f_ASAP7_75t_L g418 ( .A(n_341), .Y(n_418) );
BUFx5_ASAP7_75t_L g537 ( .A(n_341), .Y(n_537) );
BUFx3_ASAP7_75t_L g563 ( .A(n_341), .Y(n_563) );
AND2x4_ASAP7_75t_L g355 ( .A(n_342), .B(n_356), .Y(n_355) );
BUFx6f_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
BUFx6f_ASAP7_75t_L g420 ( .A(n_346), .Y(n_420) );
BUFx12f_ASAP7_75t_L g453 ( .A(n_346), .Y(n_453) );
INVx4_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
INVx4_ASAP7_75t_L g421 ( .A(n_348), .Y(n_421) );
INVx2_ASAP7_75t_L g459 ( .A(n_348), .Y(n_459) );
INVx2_ASAP7_75t_SL g502 ( .A(n_348), .Y(n_502) );
INVx2_ASAP7_75t_L g557 ( .A(n_348), .Y(n_557) );
INVx1_ASAP7_75t_L g628 ( .A(n_348), .Y(n_628) );
INVx1_ASAP7_75t_L g973 ( .A(n_348), .Y(n_973) );
INVx8_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
INVx1_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
NAND3xp33_ASAP7_75t_L g351 ( .A(n_352), .B(n_359), .C(n_368), .Y(n_351) );
INVx1_ASAP7_75t_L g987 ( .A(n_353), .Y(n_987) );
BUFx3_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
BUFx6f_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
INVx2_ASAP7_75t_L g442 ( .A(n_355), .Y(n_442) );
BUFx8_ASAP7_75t_SL g506 ( .A(n_355), .Y(n_506) );
INVx2_ASAP7_75t_L g582 ( .A(n_355), .Y(n_582) );
INVx4_ASAP7_75t_L g584 ( .A(n_357), .Y(n_584) );
BUFx6f_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
INVx3_ASAP7_75t_L g430 ( .A(n_358), .Y(n_430) );
BUFx6f_ASAP7_75t_L g549 ( .A(n_358), .Y(n_549) );
INVx2_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
INVx2_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
BUFx3_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
BUFx3_ASAP7_75t_L g424 ( .A(n_363), .Y(n_424) );
INVx1_ASAP7_75t_L g445 ( .A(n_363), .Y(n_445) );
BUFx6f_ASAP7_75t_L g511 ( .A(n_363), .Y(n_511) );
BUFx3_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
INVx1_ASAP7_75t_L g672 ( .A(n_365), .Y(n_672) );
INVx2_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
BUFx6f_ASAP7_75t_L g514 ( .A(n_366), .Y(n_514) );
INVx2_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
BUFx6f_ASAP7_75t_L g428 ( .A(n_367), .Y(n_428) );
BUFx3_ASAP7_75t_L g727 ( .A(n_367), .Y(n_727) );
INVx2_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
INVx1_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
BUFx3_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
INVx2_ASAP7_75t_L g409 ( .A(n_372), .Y(n_409) );
INVx3_ASAP7_75t_L g438 ( .A(n_372), .Y(n_438) );
OAI21xp5_ASAP7_75t_SL g373 ( .A1(n_374), .A2(n_384), .B(n_385), .Y(n_373) );
INVxp67_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
BUFx2_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
INVx5_ASAP7_75t_L g426 ( .A(n_376), .Y(n_426) );
BUFx2_ASAP7_75t_L g448 ( .A(n_376), .Y(n_448) );
AND2x4_ASAP7_75t_L g376 ( .A(n_377), .B(n_381), .Y(n_376) );
AND2x2_ASAP7_75t_L g470 ( .A(n_377), .B(n_381), .Y(n_470) );
NAND2xp5_ASAP7_75t_L g378 ( .A(n_379), .B(n_380), .Y(n_378) );
INVx1_ASAP7_75t_L g390 ( .A(n_379), .Y(n_390) );
INVx2_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
NOR2xp33_ASAP7_75t_L g639 ( .A(n_387), .B(n_640), .Y(n_639) );
BUFx6f_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
INVx2_ASAP7_75t_L g414 ( .A(n_388), .Y(n_414) );
INVx1_ASAP7_75t_L g439 ( .A(n_388), .Y(n_439) );
BUFx6f_ASAP7_75t_L g553 ( .A(n_388), .Y(n_553) );
INVx2_ASAP7_75t_SL g590 ( .A(n_388), .Y(n_590) );
NOR2xp33_ASAP7_75t_L g655 ( .A(n_388), .B(n_656), .Y(n_655) );
BUFx6f_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
INVx3_ASAP7_75t_L g480 ( .A(n_389), .Y(n_480) );
INVx1_ASAP7_75t_L g460 ( .A(n_394), .Y(n_460) );
XNOR2xp5_ASAP7_75t_L g394 ( .A(n_395), .B(n_431), .Y(n_394) );
NAND4xp75_ASAP7_75t_L g396 ( .A(n_397), .B(n_404), .C(n_415), .D(n_422), .Y(n_396) );
AND2x2_ASAP7_75t_L g397 ( .A(n_398), .B(n_401), .Y(n_397) );
BUFx3_ASAP7_75t_L g605 ( .A(n_399), .Y(n_605) );
INVx5_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
INVx3_ASAP7_75t_L g451 ( .A(n_403), .Y(n_451) );
INVx2_ASAP7_75t_L g602 ( .A(n_403), .Y(n_602) );
INVx1_ASAP7_75t_L g624 ( .A(n_403), .Y(n_624) );
INVx1_ASAP7_75t_L g683 ( .A(n_403), .Y(n_683) );
OA21x2_ASAP7_75t_L g404 ( .A1(n_405), .A2(n_406), .B(n_410), .Y(n_404) );
INVx1_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
INVx2_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
INVx2_ASAP7_75t_L g588 ( .A(n_408), .Y(n_588) );
INVx2_ASAP7_75t_L g665 ( .A(n_408), .Y(n_665) );
BUFx6f_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
NOR2xp33_ASAP7_75t_L g411 ( .A(n_412), .B(n_413), .Y(n_411) );
NOR2xp33_ASAP7_75t_L g508 ( .A(n_413), .B(n_509), .Y(n_508) );
INVx3_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
AND2x2_ASAP7_75t_L g415 ( .A(n_416), .B(n_419), .Y(n_415) );
HB1xp67_ASAP7_75t_L g613 ( .A(n_417), .Y(n_613) );
INVx1_ASAP7_75t_L g615 ( .A(n_418), .Y(n_615) );
AND2x2_ASAP7_75t_L g422 ( .A(n_423), .B(n_427), .Y(n_422) );
INVx4_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
INVx2_ASAP7_75t_L g632 ( .A(n_426), .Y(n_632) );
INVx3_ASAP7_75t_L g673 ( .A(n_426), .Y(n_673) );
INVx2_ASAP7_75t_L g728 ( .A(n_426), .Y(n_728) );
INVx2_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
INVx3_ASAP7_75t_L g446 ( .A(n_430), .Y(n_446) );
XNOR2xp5_ASAP7_75t_L g431 ( .A(n_432), .B(n_434), .Y(n_431) );
CKINVDCx5p33_ASAP7_75t_R g432 ( .A(n_433), .Y(n_432) );
NOR2x1_ASAP7_75t_L g434 ( .A(n_435), .B(n_449), .Y(n_434) );
NAND4xp25_ASAP7_75t_L g435 ( .A(n_436), .B(n_440), .C(n_443), .D(n_447), .Y(n_435) );
INVx2_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
INVx2_ASAP7_75t_L g507 ( .A(n_438), .Y(n_507) );
INVx3_ASAP7_75t_SL g634 ( .A(n_438), .Y(n_634) );
INVx3_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
INVx2_ASAP7_75t_L g532 ( .A(n_442), .Y(n_532) );
INVx2_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
NAND4xp25_ASAP7_75t_L g449 ( .A(n_450), .B(n_452), .C(n_455), .D(n_458), .Y(n_449) );
BUFx12f_ASAP7_75t_L g539 ( .A(n_453), .Y(n_539) );
INVx1_ASAP7_75t_L g595 ( .A(n_453), .Y(n_595) );
INVx1_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
INVx2_ASAP7_75t_L g536 ( .A(n_457), .Y(n_536) );
INVx1_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
AO22x1_ASAP7_75t_L g463 ( .A1(n_464), .A2(n_494), .B1(n_515), .B2(n_516), .Y(n_463) );
INVx1_ASAP7_75t_L g515 ( .A(n_464), .Y(n_515) );
INVx1_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
NOR2x1_ASAP7_75t_L g466 ( .A(n_467), .B(n_481), .Y(n_466) );
NAND4xp25_ASAP7_75t_L g467 ( .A(n_468), .B(n_471), .C(n_474), .D(n_475), .Y(n_467) );
INVx2_ASAP7_75t_L g708 ( .A(n_476), .Y(n_708) );
NOR2xp33_ASAP7_75t_L g477 ( .A(n_478), .B(n_479), .Y(n_477) );
NOR2xp33_ASAP7_75t_L g666 ( .A(n_479), .B(n_667), .Y(n_666) );
NOR2xp33_ASAP7_75t_L g724 ( .A(n_479), .B(n_725), .Y(n_724) );
INVx4_ASAP7_75t_L g993 ( .A(n_479), .Y(n_993) );
INVx4_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
NAND4xp25_ASAP7_75t_L g481 ( .A(n_482), .B(n_485), .C(n_488), .D(n_491), .Y(n_481) );
INVx1_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
INVx2_ASAP7_75t_L g517 ( .A(n_495), .Y(n_517) );
INVx2_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
NOR2x1_ASAP7_75t_L g497 ( .A(n_498), .B(n_504), .Y(n_497) );
NAND4xp25_ASAP7_75t_L g498 ( .A(n_499), .B(n_500), .C(n_501), .D(n_503), .Y(n_498) );
NAND3xp33_ASAP7_75t_L g504 ( .A(n_505), .B(n_510), .C(n_512), .Y(n_504) );
INVx4_ASAP7_75t_L g574 ( .A(n_511), .Y(n_574) );
INVx2_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
INVx1_ASAP7_75t_L g530 ( .A(n_514), .Y(n_530) );
INVx2_ASAP7_75t_L g577 ( .A(n_514), .Y(n_577) );
INVx2_ASAP7_75t_L g984 ( .A(n_514), .Y(n_984) );
INVx1_ASAP7_75t_L g516 ( .A(n_517), .Y(n_516) );
XNOR2xp5_ASAP7_75t_L g518 ( .A(n_519), .B(n_644), .Y(n_518) );
OAI22xp5_ASAP7_75t_L g519 ( .A1(n_520), .A2(n_566), .B1(n_642), .B2(n_643), .Y(n_519) );
INVx1_ASAP7_75t_L g642 ( .A(n_520), .Y(n_642) );
AOI22xp5_ASAP7_75t_L g520 ( .A1(n_521), .A2(n_542), .B1(n_564), .B2(n_565), .Y(n_520) );
INVx1_ASAP7_75t_L g564 ( .A(n_521), .Y(n_564) );
INVx1_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
INVx2_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
XNOR2xp5_ASAP7_75t_L g523 ( .A(n_524), .B(n_525), .Y(n_523) );
NOR2xp67_ASAP7_75t_L g525 ( .A(n_526), .B(n_533), .Y(n_525) );
NAND3xp33_ASAP7_75t_L g526 ( .A(n_527), .B(n_529), .C(n_531), .Y(n_526) );
NAND4xp25_ASAP7_75t_L g533 ( .A(n_534), .B(n_538), .C(n_540), .D(n_541), .Y(n_533) );
BUFx4f_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
INVx2_ASAP7_75t_L g565 ( .A(n_542), .Y(n_565) );
INVx1_ASAP7_75t_SL g542 ( .A(n_543), .Y(n_542) );
NOR2x1_ASAP7_75t_L g544 ( .A(n_545), .B(n_554), .Y(n_544) );
NAND4xp25_ASAP7_75t_L g545 ( .A(n_546), .B(n_547), .C(n_548), .D(n_550), .Y(n_545) );
BUFx3_ASAP7_75t_L g669 ( .A(n_549), .Y(n_669) );
NOR2xp33_ASAP7_75t_L g551 ( .A(n_552), .B(n_553), .Y(n_551) );
NOR2xp33_ASAP7_75t_L g709 ( .A(n_553), .B(n_710), .Y(n_709) );
NAND4xp25_ASAP7_75t_L g554 ( .A(n_555), .B(n_556), .C(n_560), .D(n_562), .Y(n_554) );
BUFx4f_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
BUFx6f_ASAP7_75t_L g977 ( .A(n_559), .Y(n_977) );
BUFx3_ASAP7_75t_L g968 ( .A(n_561), .Y(n_968) );
INVx1_ASAP7_75t_L g643 ( .A(n_566), .Y(n_643) );
OAI22xp5_ASAP7_75t_L g566 ( .A1(n_567), .A2(n_568), .B1(n_618), .B2(n_619), .Y(n_566) );
INVx4_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
AO22x2_ASAP7_75t_L g568 ( .A1(n_569), .A2(n_570), .B1(n_591), .B2(n_616), .Y(n_568) );
NOR4xp25_ASAP7_75t_L g569 ( .A(n_570), .B(n_572), .C(n_578), .D(n_585), .Y(n_569) );
CKINVDCx5p33_ASAP7_75t_R g570 ( .A(n_571), .Y(n_570) );
NOR3xp33_ASAP7_75t_SL g617 ( .A(n_572), .B(n_578), .C(n_585), .Y(n_617) );
OAI22xp33_ASAP7_75t_L g572 ( .A1(n_573), .A2(n_574), .B1(n_575), .B2(n_576), .Y(n_572) );
OAI22xp5_ASAP7_75t_L g980 ( .A1(n_574), .A2(n_981), .B1(n_982), .B2(n_983), .Y(n_980) );
INVx1_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
OAI22xp33_ASAP7_75t_L g578 ( .A1(n_579), .A2(n_580), .B1(n_583), .B2(n_584), .Y(n_578) );
INVx2_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
INVx2_ASAP7_75t_SL g581 ( .A(n_582), .Y(n_581) );
INVx2_ASAP7_75t_SL g637 ( .A(n_582), .Y(n_637) );
OAI22xp5_ASAP7_75t_L g985 ( .A1(n_584), .A2(n_986), .B1(n_987), .B2(n_988), .Y(n_985) );
OAI21xp33_ASAP7_75t_L g585 ( .A1(n_586), .A2(n_587), .B(n_589), .Y(n_585) );
INVx1_ASAP7_75t_L g587 ( .A(n_588), .Y(n_587) );
NAND2xp5_ASAP7_75t_SL g616 ( .A(n_591), .B(n_617), .Y(n_616) );
NOR3xp33_ASAP7_75t_L g591 ( .A(n_592), .B(n_603), .C(n_610), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g592 ( .A(n_593), .B(n_596), .Y(n_592) );
INVx1_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
INVx1_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
INVx1_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
INVx1_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
INVx1_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
HB1xp67_ASAP7_75t_L g969 ( .A(n_602), .Y(n_969) );
OAI22xp5_ASAP7_75t_L g603 ( .A1(n_604), .A2(n_606), .B1(n_607), .B2(n_608), .Y(n_603) );
INVx1_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
OAI22xp5_ASAP7_75t_L g974 ( .A1(n_608), .A2(n_975), .B1(n_976), .B2(n_978), .Y(n_974) );
INVx1_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
OAI22x1_ASAP7_75t_SL g610 ( .A1(n_611), .A2(n_612), .B1(n_614), .B2(n_615), .Y(n_610) );
INVx1_ASAP7_75t_L g612 ( .A(n_613), .Y(n_612) );
INVx1_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
BUFx2_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
XNOR2x1_ASAP7_75t_L g620 ( .A(n_621), .B(n_641), .Y(n_620) );
NOR4xp75_ASAP7_75t_L g621 ( .A(n_622), .B(n_626), .C(n_630), .D(n_635), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g622 ( .A(n_623), .B(n_625), .Y(n_622) );
NAND2xp5_ASAP7_75t_L g626 ( .A(n_627), .B(n_629), .Y(n_626) );
NAND2xp5_ASAP7_75t_L g630 ( .A(n_631), .B(n_633), .Y(n_630) );
INVx1_ASAP7_75t_L g991 ( .A(n_634), .Y(n_991) );
NAND2xp5_ASAP7_75t_SL g635 ( .A(n_636), .B(n_638), .Y(n_635) );
XOR2xp5_ASAP7_75t_L g644 ( .A(n_645), .B(n_691), .Y(n_644) );
HB1xp67_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
XNOR2xp5_ASAP7_75t_L g646 ( .A(n_647), .B(n_661), .Y(n_646) );
INVx1_ASAP7_75t_L g659 ( .A(n_648), .Y(n_659) );
NAND3xp33_ASAP7_75t_L g648 ( .A(n_649), .B(n_654), .C(n_657), .Y(n_648) );
AND4x1_ASAP7_75t_L g649 ( .A(n_650), .B(n_651), .C(n_652), .D(n_653), .Y(n_649) );
NOR2x1_ASAP7_75t_L g662 ( .A(n_663), .B(n_674), .Y(n_662) );
NAND3xp33_ASAP7_75t_L g663 ( .A(n_664), .B(n_668), .C(n_670), .Y(n_663) );
INVx1_ASAP7_75t_L g689 ( .A(n_664), .Y(n_689) );
INVxp67_ASAP7_75t_SL g690 ( .A(n_668), .Y(n_690) );
INVx1_ASAP7_75t_L g686 ( .A(n_670), .Y(n_686) );
INVx1_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
NAND2xp5_ASAP7_75t_L g674 ( .A(n_675), .B(n_679), .Y(n_674) );
INVx1_ASAP7_75t_L g675 ( .A(n_676), .Y(n_675) );
NOR3xp33_ASAP7_75t_L g685 ( .A(n_676), .B(n_686), .C(n_687), .Y(n_685) );
NAND2xp5_ASAP7_75t_L g676 ( .A(n_677), .B(n_678), .Y(n_676) );
INVx1_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
NOR3xp33_ASAP7_75t_L g688 ( .A(n_680), .B(n_689), .C(n_690), .Y(n_688) );
NAND2xp5_ASAP7_75t_L g680 ( .A(n_681), .B(n_682), .Y(n_680) );
NAND2xp5_ASAP7_75t_L g684 ( .A(n_685), .B(n_688), .Y(n_684) );
AOI22x1_ASAP7_75t_L g691 ( .A1(n_692), .A2(n_712), .B1(n_735), .B2(n_736), .Y(n_691) );
INVx1_ASAP7_75t_L g692 ( .A(n_693), .Y(n_692) );
INVx1_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
INVx1_ASAP7_75t_L g736 ( .A(n_694), .Y(n_736) );
INVx1_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
INVx1_ASAP7_75t_L g695 ( .A(n_696), .Y(n_695) );
NOR2x1_ASAP7_75t_L g697 ( .A(n_698), .B(n_704), .Y(n_697) );
NAND4xp25_ASAP7_75t_L g698 ( .A(n_699), .B(n_701), .C(n_702), .D(n_703), .Y(n_698) );
NAND3xp33_ASAP7_75t_L g704 ( .A(n_705), .B(n_706), .C(n_711), .Y(n_704) );
INVx2_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
INVx2_ASAP7_75t_L g735 ( .A(n_712), .Y(n_735) );
INVx2_ASAP7_75t_L g712 ( .A(n_713), .Y(n_712) );
BUFx3_ASAP7_75t_L g713 ( .A(n_714), .Y(n_713) );
NAND4xp25_ASAP7_75t_L g732 ( .A(n_716), .B(n_717), .C(n_719), .D(n_729), .Y(n_732) );
NAND2xp5_ASAP7_75t_L g734 ( .A(n_718), .B(n_730), .Y(n_734) );
NAND3xp33_ASAP7_75t_L g720 ( .A(n_721), .B(n_729), .C(n_730), .Y(n_720) );
INVxp67_ASAP7_75t_L g721 ( .A(n_722), .Y(n_721) );
OR2x2_ASAP7_75t_L g733 ( .A(n_722), .B(n_734), .Y(n_733) );
NAND2xp5_ASAP7_75t_L g722 ( .A(n_723), .B(n_726), .Y(n_722) );
NOR2x1_ASAP7_75t_L g731 ( .A(n_732), .B(n_733), .Y(n_731) );
OAI21xp5_ASAP7_75t_L g737 ( .A1(n_738), .A2(n_959), .B(n_961), .Y(n_737) );
NOR3xp33_ASAP7_75t_L g738 ( .A(n_739), .B(n_886), .C(n_924), .Y(n_738) );
OAI221xp5_ASAP7_75t_SL g739 ( .A1(n_740), .A2(n_844), .B1(n_845), .B2(n_850), .C(n_870), .Y(n_739) );
NOR4xp25_ASAP7_75t_L g740 ( .A(n_741), .B(n_815), .C(n_829), .D(n_837), .Y(n_740) );
OAI211xp5_ASAP7_75t_SL g741 ( .A1(n_742), .A2(n_763), .B(n_781), .C(n_808), .Y(n_741) );
INVx1_ASAP7_75t_L g813 ( .A(n_742), .Y(n_813) );
NOR2x1_ASAP7_75t_L g912 ( .A(n_742), .B(n_818), .Y(n_912) );
OR2x2_ASAP7_75t_L g742 ( .A(n_743), .B(n_755), .Y(n_742) );
INVx1_ASAP7_75t_L g799 ( .A(n_743), .Y(n_799) );
AND2x2_ASAP7_75t_L g828 ( .A(n_743), .B(n_792), .Y(n_828) );
AND2x2_ASAP7_75t_L g834 ( .A(n_743), .B(n_755), .Y(n_834) );
NAND2xp5_ASAP7_75t_L g922 ( .A(n_743), .B(n_789), .Y(n_922) );
OAI321xp33_ASAP7_75t_L g943 ( .A1(n_743), .A2(n_826), .A3(n_918), .B1(n_944), .B2(n_945), .C(n_947), .Y(n_943) );
AND2x2_ASAP7_75t_L g957 ( .A(n_743), .B(n_788), .Y(n_957) );
INVx3_ASAP7_75t_L g848 ( .A(n_744), .Y(n_848) );
AND2x4_ASAP7_75t_L g744 ( .A(n_745), .B(n_747), .Y(n_744) );
AND2x4_ASAP7_75t_L g752 ( .A(n_745), .B(n_753), .Y(n_752) );
AND2x2_ASAP7_75t_L g761 ( .A(n_745), .B(n_753), .Y(n_761) );
AND2x2_ASAP7_75t_L g770 ( .A(n_745), .B(n_753), .Y(n_770) );
AND2x4_ASAP7_75t_L g749 ( .A(n_747), .B(n_750), .Y(n_749) );
AND2x4_ASAP7_75t_L g759 ( .A(n_747), .B(n_750), .Y(n_759) );
NAND2xp5_ASAP7_75t_L g960 ( .A(n_747), .B(n_750), .Y(n_960) );
CKINVDCx5p33_ASAP7_75t_R g1004 ( .A(n_747), .Y(n_1004) );
AND2x2_ASAP7_75t_L g754 ( .A(n_750), .B(n_753), .Y(n_754) );
AND2x2_ASAP7_75t_L g762 ( .A(n_750), .B(n_753), .Y(n_762) );
AND2x4_ASAP7_75t_L g771 ( .A(n_750), .B(n_753), .Y(n_771) );
INVx1_ASAP7_75t_L g792 ( .A(n_755), .Y(n_792) );
AND2x2_ASAP7_75t_L g804 ( .A(n_755), .B(n_789), .Y(n_804) );
AND2x2_ASAP7_75t_L g823 ( .A(n_755), .B(n_799), .Y(n_823) );
AND2x2_ASAP7_75t_L g755 ( .A(n_756), .B(n_760), .Y(n_755) );
INVx2_ASAP7_75t_SL g768 ( .A(n_759), .Y(n_768) );
INVx1_ASAP7_75t_L g940 ( .A(n_763), .Y(n_940) );
NAND2xp5_ASAP7_75t_L g763 ( .A(n_764), .B(n_772), .Y(n_763) );
AND2x2_ASAP7_75t_L g800 ( .A(n_764), .B(n_777), .Y(n_800) );
NAND2xp5_ASAP7_75t_L g824 ( .A(n_764), .B(n_802), .Y(n_824) );
AND2x2_ASAP7_75t_L g836 ( .A(n_764), .B(n_826), .Y(n_836) );
OR2x2_ASAP7_75t_L g862 ( .A(n_764), .B(n_863), .Y(n_862) );
NAND2xp5_ASAP7_75t_L g918 ( .A(n_764), .B(n_784), .Y(n_918) );
NOR2xp33_ASAP7_75t_L g938 ( .A(n_764), .B(n_844), .Y(n_938) );
NOR2xp33_ASAP7_75t_L g954 ( .A(n_764), .B(n_843), .Y(n_954) );
INVx4_ASAP7_75t_L g764 ( .A(n_765), .Y(n_764) );
AND2x2_ASAP7_75t_L g853 ( .A(n_765), .B(n_854), .Y(n_853) );
AND2x2_ASAP7_75t_L g859 ( .A(n_765), .B(n_778), .Y(n_859) );
NAND3xp33_ASAP7_75t_L g864 ( .A(n_765), .B(n_823), .C(n_865), .Y(n_864) );
INVx1_ASAP7_75t_L g876 ( .A(n_765), .Y(n_876) );
NOR2xp33_ASAP7_75t_L g898 ( .A(n_765), .B(n_845), .Y(n_898) );
AND2x2_ASAP7_75t_L g901 ( .A(n_765), .B(n_826), .Y(n_901) );
NOR2xp33_ASAP7_75t_L g946 ( .A(n_765), .B(n_855), .Y(n_946) );
NOR3xp33_ASAP7_75t_SL g948 ( .A(n_765), .B(n_879), .C(n_915), .Y(n_948) );
AND2x2_ASAP7_75t_L g765 ( .A(n_766), .B(n_769), .Y(n_765) );
INVx2_ASAP7_75t_L g767 ( .A(n_768), .Y(n_767) );
INVx1_ASAP7_75t_L g772 ( .A(n_773), .Y(n_772) );
OAI332xp33_ASAP7_75t_L g913 ( .A1(n_773), .A2(n_858), .A3(n_914), .B1(n_917), .B2(n_918), .B3(n_919), .C1(n_920), .C2(n_923), .Y(n_913) );
OAI222xp33_ASAP7_75t_SL g930 ( .A1(n_773), .A2(n_788), .B1(n_843), .B2(n_931), .C1(n_935), .C2(n_936), .Y(n_930) );
OR2x2_ASAP7_75t_L g773 ( .A(n_774), .B(n_777), .Y(n_773) );
INVx4_ASAP7_75t_L g797 ( .A(n_774), .Y(n_797) );
OR2x2_ASAP7_75t_L g843 ( .A(n_774), .B(n_778), .Y(n_843) );
NOR2xp33_ASAP7_75t_L g861 ( .A(n_774), .B(n_807), .Y(n_861) );
NOR2xp33_ASAP7_75t_L g865 ( .A(n_774), .B(n_784), .Y(n_865) );
AND2x2_ASAP7_75t_L g868 ( .A(n_774), .B(n_777), .Y(n_868) );
NAND2xp5_ASAP7_75t_L g879 ( .A(n_774), .B(n_807), .Y(n_879) );
AND2x2_ASAP7_75t_L g774 ( .A(n_775), .B(n_776), .Y(n_774) );
INVx2_ASAP7_75t_L g802 ( .A(n_777), .Y(n_802) );
OR2x2_ASAP7_75t_L g855 ( .A(n_777), .B(n_797), .Y(n_855) );
INVxp67_ASAP7_75t_L g863 ( .A(n_777), .Y(n_863) );
INVx2_ASAP7_75t_L g777 ( .A(n_778), .Y(n_777) );
NAND2xp5_ASAP7_75t_L g778 ( .A(n_779), .B(n_780), .Y(n_778) );
O2A1O1Ixp33_ASAP7_75t_L g781 ( .A1(n_782), .A2(n_793), .B(n_800), .C(n_801), .Y(n_781) );
NOR2xp33_ASAP7_75t_L g782 ( .A(n_783), .B(n_787), .Y(n_782) );
AND2x2_ASAP7_75t_L g831 ( .A(n_783), .B(n_827), .Y(n_831) );
NAND2xp5_ASAP7_75t_L g891 ( .A(n_783), .B(n_892), .Y(n_891) );
NAND2xp5_ASAP7_75t_L g905 ( .A(n_783), .B(n_822), .Y(n_905) );
AND2x2_ASAP7_75t_L g958 ( .A(n_783), .B(n_854), .Y(n_958) );
INVx2_ASAP7_75t_L g783 ( .A(n_784), .Y(n_783) );
INVx2_ASAP7_75t_L g807 ( .A(n_784), .Y(n_807) );
AND2x2_ASAP7_75t_L g814 ( .A(n_784), .B(n_788), .Y(n_814) );
INVx3_ASAP7_75t_L g819 ( .A(n_784), .Y(n_819) );
AOI211xp5_ASAP7_75t_L g850 ( .A1(n_784), .A2(n_851), .B(n_856), .C(n_866), .Y(n_850) );
NOR2xp33_ASAP7_75t_L g921 ( .A(n_784), .B(n_922), .Y(n_921) );
NAND2xp5_ASAP7_75t_L g935 ( .A(n_784), .B(n_868), .Y(n_935) );
AND2x2_ASAP7_75t_L g784 ( .A(n_785), .B(n_786), .Y(n_784) );
INVx1_ASAP7_75t_L g892 ( .A(n_787), .Y(n_892) );
NAND2xp5_ASAP7_75t_L g787 ( .A(n_788), .B(n_792), .Y(n_787) );
AND2x2_ASAP7_75t_L g821 ( .A(n_788), .B(n_813), .Y(n_821) );
AND2x2_ASAP7_75t_L g833 ( .A(n_788), .B(n_834), .Y(n_833) );
NAND2xp5_ASAP7_75t_L g840 ( .A(n_788), .B(n_823), .Y(n_840) );
NAND2xp5_ASAP7_75t_L g873 ( .A(n_788), .B(n_874), .Y(n_873) );
AND2x2_ASAP7_75t_L g880 ( .A(n_788), .B(n_828), .Y(n_880) );
NAND2xp5_ASAP7_75t_L g911 ( .A(n_788), .B(n_912), .Y(n_911) );
CKINVDCx6p67_ASAP7_75t_R g788 ( .A(n_789), .Y(n_788) );
NAND2xp5_ASAP7_75t_L g798 ( .A(n_789), .B(n_799), .Y(n_798) );
AND2x2_ASAP7_75t_L g822 ( .A(n_789), .B(n_823), .Y(n_822) );
AND2x2_ASAP7_75t_L g827 ( .A(n_789), .B(n_828), .Y(n_827) );
AND2x2_ASAP7_75t_L g842 ( .A(n_789), .B(n_813), .Y(n_842) );
AND2x2_ASAP7_75t_L g884 ( .A(n_789), .B(n_818), .Y(n_884) );
AND2x2_ASAP7_75t_L g928 ( .A(n_789), .B(n_874), .Y(n_928) );
NOR2xp33_ASAP7_75t_L g934 ( .A(n_789), .B(n_792), .Y(n_934) );
AND2x2_ASAP7_75t_L g941 ( .A(n_789), .B(n_792), .Y(n_941) );
AND2x2_ASAP7_75t_L g789 ( .A(n_790), .B(n_791), .Y(n_789) );
NAND2xp5_ASAP7_75t_L g860 ( .A(n_792), .B(n_861), .Y(n_860) );
NOR2xp33_ASAP7_75t_L g793 ( .A(n_794), .B(n_798), .Y(n_793) );
NAND2xp5_ASAP7_75t_L g882 ( .A(n_794), .B(n_883), .Y(n_882) );
AOI221xp5_ASAP7_75t_L g925 ( .A1(n_794), .A2(n_926), .B1(n_928), .B2(n_929), .C(n_930), .Y(n_925) );
INVx2_ASAP7_75t_L g794 ( .A(n_795), .Y(n_794) );
HB1xp67_ASAP7_75t_L g929 ( .A(n_795), .Y(n_929) );
INVx1_ASAP7_75t_L g795 ( .A(n_796), .Y(n_795) );
INVx1_ASAP7_75t_L g806 ( .A(n_796), .Y(n_806) );
INVx1_ASAP7_75t_L g796 ( .A(n_797), .Y(n_796) );
INVx2_ASAP7_75t_L g826 ( .A(n_797), .Y(n_826) );
AOI221xp5_ASAP7_75t_L g887 ( .A1(n_799), .A2(n_817), .B1(n_888), .B2(n_890), .C(n_893), .Y(n_887) );
AOI221xp5_ASAP7_75t_L g906 ( .A1(n_800), .A2(n_907), .B1(n_908), .B2(n_910), .C(n_913), .Y(n_906) );
NAND2xp5_ASAP7_75t_L g923 ( .A(n_800), .B(n_904), .Y(n_923) );
NOR2xp33_ASAP7_75t_L g801 ( .A(n_802), .B(n_803), .Y(n_801) );
INVx3_ASAP7_75t_SL g817 ( .A(n_802), .Y(n_817) );
NAND2xp5_ASAP7_75t_L g885 ( .A(n_802), .B(n_844), .Y(n_885) );
NAND2xp5_ASAP7_75t_L g909 ( .A(n_802), .B(n_845), .Y(n_909) );
NAND2xp5_ASAP7_75t_L g803 ( .A(n_804), .B(n_805), .Y(n_803) );
INVx1_ASAP7_75t_L g919 ( .A(n_804), .Y(n_919) );
NOR2xp33_ASAP7_75t_L g805 ( .A(n_806), .B(n_807), .Y(n_805) );
INVx1_ASAP7_75t_L g811 ( .A(n_806), .Y(n_811) );
NOR2xp33_ASAP7_75t_L g932 ( .A(n_807), .B(n_933), .Y(n_932) );
NAND2xp5_ASAP7_75t_L g808 ( .A(n_809), .B(n_812), .Y(n_808) );
NOR2xp33_ASAP7_75t_L g910 ( .A(n_809), .B(n_911), .Y(n_910) );
HB1xp67_ASAP7_75t_L g809 ( .A(n_810), .Y(n_809) );
INVx1_ASAP7_75t_L g810 ( .A(n_811), .Y(n_810) );
INVx1_ASAP7_75t_L g904 ( .A(n_811), .Y(n_904) );
AND2x2_ASAP7_75t_L g812 ( .A(n_813), .B(n_814), .Y(n_812) );
AND2x2_ASAP7_75t_L g883 ( .A(n_813), .B(n_884), .Y(n_883) );
INVxp67_ASAP7_75t_L g917 ( .A(n_814), .Y(n_917) );
OAI22xp33_ASAP7_75t_SL g815 ( .A1(n_816), .A2(n_820), .B1(n_824), .B2(n_825), .Y(n_815) );
NAND2xp5_ASAP7_75t_L g816 ( .A(n_817), .B(n_818), .Y(n_816) );
AOI221xp5_ASAP7_75t_L g939 ( .A1(n_817), .A2(n_940), .B1(n_941), .B2(n_942), .C(n_943), .Y(n_939) );
NOR2x1_ASAP7_75t_L g839 ( .A(n_818), .B(n_840), .Y(n_839) );
NOR2xp33_ASAP7_75t_L g888 ( .A(n_818), .B(n_889), .Y(n_888) );
AND2x2_ASAP7_75t_L g907 ( .A(n_818), .B(n_869), .Y(n_907) );
INVx3_ASAP7_75t_L g818 ( .A(n_819), .Y(n_818) );
AND2x2_ASAP7_75t_L g874 ( .A(n_819), .B(n_834), .Y(n_874) );
NOR2xp33_ASAP7_75t_L g820 ( .A(n_821), .B(n_822), .Y(n_820) );
INVx1_ASAP7_75t_L g955 ( .A(n_821), .Y(n_955) );
INVx1_ASAP7_75t_L g857 ( .A(n_822), .Y(n_857) );
OAI21xp5_ASAP7_75t_L g956 ( .A1(n_822), .A2(n_957), .B(n_958), .Y(n_956) );
INVx1_ASAP7_75t_L g915 ( .A(n_823), .Y(n_915) );
INVx1_ASAP7_75t_L g871 ( .A(n_824), .Y(n_871) );
NAND2xp5_ASAP7_75t_L g825 ( .A(n_826), .B(n_827), .Y(n_825) );
O2A1O1Ixp33_ASAP7_75t_L g881 ( .A1(n_826), .A2(n_832), .B(n_882), .C(n_885), .Y(n_881) );
INVx1_ASAP7_75t_L g936 ( .A(n_827), .Y(n_936) );
NAND2xp5_ASAP7_75t_L g852 ( .A(n_828), .B(n_853), .Y(n_852) );
NAND2xp5_ASAP7_75t_L g896 ( .A(n_828), .B(n_884), .Y(n_896) );
INVx1_ASAP7_75t_L g916 ( .A(n_828), .Y(n_916) );
AOI21xp5_ASAP7_75t_L g829 ( .A1(n_830), .A2(n_832), .B(n_835), .Y(n_829) );
INVx1_ASAP7_75t_L g830 ( .A(n_831), .Y(n_830) );
INVx1_ASAP7_75t_L g832 ( .A(n_833), .Y(n_832) );
NAND2xp5_ASAP7_75t_L g927 ( .A(n_834), .B(n_884), .Y(n_927) );
INVx1_ASAP7_75t_L g944 ( .A(n_834), .Y(n_944) );
INVx1_ASAP7_75t_L g835 ( .A(n_836), .Y(n_835) );
AOI21xp33_ASAP7_75t_L g837 ( .A1(n_838), .A2(n_841), .B(n_843), .Y(n_837) );
INVx1_ASAP7_75t_L g838 ( .A(n_839), .Y(n_838) );
INVx1_ASAP7_75t_L g869 ( .A(n_840), .Y(n_869) );
NAND2xp5_ASAP7_75t_L g926 ( .A(n_841), .B(n_927), .Y(n_926) );
INVx1_ASAP7_75t_L g841 ( .A(n_842), .Y(n_841) );
CKINVDCx5p33_ASAP7_75t_R g844 ( .A(n_845), .Y(n_844) );
OAI221xp5_ASAP7_75t_SL g886 ( .A1(n_845), .A2(n_887), .B1(n_897), .B2(n_899), .C(n_906), .Y(n_886) );
OAI221xp5_ASAP7_75t_SL g924 ( .A1(n_845), .A2(n_925), .B1(n_937), .B2(n_939), .C(n_949), .Y(n_924) );
AND2x2_ASAP7_75t_L g845 ( .A(n_846), .B(n_849), .Y(n_845) );
INVx1_ASAP7_75t_L g847 ( .A(n_848), .Y(n_847) );
INVxp67_ASAP7_75t_SL g851 ( .A(n_852), .Y(n_851) );
AOI221xp5_ASAP7_75t_L g949 ( .A1(n_853), .A2(n_890), .B1(n_950), .B2(n_951), .C(n_952), .Y(n_949) );
INVx1_ASAP7_75t_L g854 ( .A(n_855), .Y(n_854) );
OAI221xp5_ASAP7_75t_L g856 ( .A1(n_857), .A2(n_858), .B1(n_860), .B2(n_862), .C(n_864), .Y(n_856) );
INVx1_ASAP7_75t_L g858 ( .A(n_859), .Y(n_858) );
INVxp67_ASAP7_75t_SL g866 ( .A(n_867), .Y(n_866) );
NAND2xp5_ASAP7_75t_L g867 ( .A(n_868), .B(n_869), .Y(n_867) );
INVx1_ASAP7_75t_L g889 ( .A(n_868), .Y(n_889) );
NAND2xp5_ASAP7_75t_L g894 ( .A(n_868), .B(n_895), .Y(n_894) );
AOI211xp5_ASAP7_75t_L g870 ( .A1(n_871), .A2(n_872), .B(n_875), .C(n_881), .Y(n_870) );
AOI21xp5_ASAP7_75t_L g899 ( .A1(n_872), .A2(n_900), .B(n_902), .Y(n_899) );
INVx1_ASAP7_75t_L g872 ( .A(n_873), .Y(n_872) );
NOR2xp33_ASAP7_75t_L g875 ( .A(n_876), .B(n_877), .Y(n_875) );
NAND2xp5_ASAP7_75t_L g877 ( .A(n_878), .B(n_880), .Y(n_877) );
INVx1_ASAP7_75t_L g878 ( .A(n_879), .Y(n_878) );
INVxp67_ASAP7_75t_SL g951 ( .A(n_885), .Y(n_951) );
INVx1_ASAP7_75t_L g890 ( .A(n_891), .Y(n_890) );
INVxp67_ASAP7_75t_SL g893 ( .A(n_894), .Y(n_893) );
INVx1_ASAP7_75t_L g895 ( .A(n_896), .Y(n_895) );
INVx1_ASAP7_75t_L g897 ( .A(n_898), .Y(n_897) );
INVx1_ASAP7_75t_L g900 ( .A(n_901), .Y(n_900) );
NOR2xp33_ASAP7_75t_L g902 ( .A(n_903), .B(n_905), .Y(n_902) );
HB1xp67_ASAP7_75t_L g903 ( .A(n_904), .Y(n_903) );
INVx1_ASAP7_75t_L g950 ( .A(n_905), .Y(n_950) );
INVxp67_ASAP7_75t_SL g908 ( .A(n_909), .Y(n_908) );
INVx1_ASAP7_75t_L g942 ( .A(n_911), .Y(n_942) );
AND2x2_ASAP7_75t_L g914 ( .A(n_915), .B(n_916), .Y(n_914) );
INVx1_ASAP7_75t_L g920 ( .A(n_921), .Y(n_920) );
INVxp67_ASAP7_75t_L g931 ( .A(n_932), .Y(n_931) );
INVx1_ASAP7_75t_L g933 ( .A(n_934), .Y(n_933) );
INVx1_ASAP7_75t_L g937 ( .A(n_938), .Y(n_937) );
INVx1_ASAP7_75t_L g945 ( .A(n_946), .Y(n_945) );
INVxp67_ASAP7_75t_L g947 ( .A(n_948), .Y(n_947) );
OAI21xp5_ASAP7_75t_L g952 ( .A1(n_953), .A2(n_955), .B(n_956), .Y(n_952) );
INVx1_ASAP7_75t_L g953 ( .A(n_954), .Y(n_953) );
BUFx2_ASAP7_75t_L g959 ( .A(n_960), .Y(n_959) );
INVx1_ASAP7_75t_L g962 ( .A(n_963), .Y(n_962) );
INVx2_ASAP7_75t_L g963 ( .A(n_964), .Y(n_963) );
HB1xp67_ASAP7_75t_L g999 ( .A(n_965), .Y(n_999) );
NAND2xp5_ASAP7_75t_L g965 ( .A(n_966), .B(n_979), .Y(n_965) );
NOR3xp33_ASAP7_75t_L g966 ( .A(n_967), .B(n_970), .C(n_974), .Y(n_966) );
NAND2xp5_ASAP7_75t_L g970 ( .A(n_971), .B(n_972), .Y(n_970) );
INVxp67_ASAP7_75t_L g976 ( .A(n_977), .Y(n_976) );
NOR3xp33_ASAP7_75t_L g979 ( .A(n_980), .B(n_985), .C(n_989), .Y(n_979) );
INVxp67_ASAP7_75t_L g983 ( .A(n_984), .Y(n_983) );
OAI21xp33_ASAP7_75t_L g989 ( .A1(n_990), .A2(n_991), .B(n_992), .Y(n_989) );
HB1xp67_ASAP7_75t_L g994 ( .A(n_995), .Y(n_994) );
HB1xp67_ASAP7_75t_L g1000 ( .A(n_1001), .Y(n_1000) );
BUFx2_ASAP7_75t_L g1002 ( .A(n_1003), .Y(n_1002) );
endmodule