module fake_ariane_2010_n_157 (n_8, n_24, n_7, n_22, n_1, n_6, n_13, n_20, n_27, n_29, n_17, n_4, n_41, n_38, n_2, n_18, n_32, n_28, n_37, n_9, n_11, n_34, n_26, n_3, n_14, n_0, n_36, n_33, n_19, n_30, n_39, n_40, n_31, n_16, n_5, n_12, n_15, n_21, n_23, n_35, n_10, n_25, n_157);

input n_8;
input n_24;
input n_7;
input n_22;
input n_1;
input n_6;
input n_13;
input n_20;
input n_27;
input n_29;
input n_17;
input n_4;
input n_41;
input n_38;
input n_2;
input n_18;
input n_32;
input n_28;
input n_37;
input n_9;
input n_11;
input n_34;
input n_26;
input n_3;
input n_14;
input n_0;
input n_36;
input n_33;
input n_19;
input n_30;
input n_39;
input n_40;
input n_31;
input n_16;
input n_5;
input n_12;
input n_15;
input n_21;
input n_23;
input n_35;
input n_10;
input n_25;

output n_157;

wire n_83;
wire n_56;
wire n_60;
wire n_64;
wire n_124;
wire n_119;
wire n_90;
wire n_47;
wire n_110;
wire n_153;
wire n_86;
wire n_75;
wire n_89;
wire n_67;
wire n_149;
wire n_69;
wire n_95;
wire n_92;
wire n_143;
wire n_150;
wire n_98;
wire n_74;
wire n_113;
wire n_114;
wire n_152;
wire n_120;
wire n_106;
wire n_53;
wire n_111;
wire n_115;
wire n_133;
wire n_66;
wire n_71;
wire n_109;
wire n_96;
wire n_156;
wire n_49;
wire n_100;
wire n_50;
wire n_132;
wire n_62;
wire n_147;
wire n_51;
wire n_76;
wire n_103;
wire n_79;
wire n_46;
wire n_84;
wire n_91;
wire n_107;
wire n_72;
wire n_105;
wire n_128;
wire n_44;
wire n_82;
wire n_42;
wire n_57;
wire n_131;
wire n_70;
wire n_117;
wire n_139;
wire n_85;
wire n_130;
wire n_144;
wire n_48;
wire n_94;
wire n_101;
wire n_134;
wire n_58;
wire n_65;
wire n_123;
wire n_138;
wire n_112;
wire n_45;
wire n_129;
wire n_126;
wire n_137;
wire n_122;
wire n_148;
wire n_52;
wire n_135;
wire n_73;
wire n_77;
wire n_121;
wire n_93;
wire n_118;
wire n_61;
wire n_108;
wire n_102;
wire n_125;
wire n_43;
wire n_87;
wire n_81;
wire n_140;
wire n_55;
wire n_151;
wire n_136;
wire n_80;
wire n_146;
wire n_97;
wire n_154;
wire n_142;
wire n_88;
wire n_141;
wire n_68;
wire n_116;
wire n_104;
wire n_145;
wire n_78;
wire n_63;
wire n_59;
wire n_99;
wire n_155;
wire n_127;
wire n_54;

INVx1_ASAP7_75t_L g42 ( 
.A(n_21),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_16),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_39),
.Y(n_44)
);

CKINVDCx5p33_ASAP7_75t_R g45 ( 
.A(n_9),
.Y(n_45)
);

INVxp33_ASAP7_75t_L g46 ( 
.A(n_19),
.Y(n_46)
);

INVxp33_ASAP7_75t_SL g47 ( 
.A(n_17),
.Y(n_47)
);

CKINVDCx16_ASAP7_75t_R g48 ( 
.A(n_7),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_14),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_8),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_32),
.Y(n_51)
);

HB1xp67_ASAP7_75t_L g52 ( 
.A(n_30),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_41),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_4),
.Y(n_55)
);

CKINVDCx16_ASAP7_75t_R g56 ( 
.A(n_2),
.Y(n_56)
);

CKINVDCx5p33_ASAP7_75t_R g57 ( 
.A(n_38),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_34),
.Y(n_58)
);

INVxp67_ASAP7_75t_L g59 ( 
.A(n_29),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_3),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_31),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_15),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_22),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_5),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_40),
.Y(n_65)
);

CKINVDCx5p33_ASAP7_75t_R g66 ( 
.A(n_4),
.Y(n_66)
);

CKINVDCx14_ASAP7_75t_R g67 ( 
.A(n_13),
.Y(n_67)
);

INVxp67_ASAP7_75t_SL g68 ( 
.A(n_27),
.Y(n_68)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_55),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_60),
.Y(n_70)
);

OAI21xp33_ASAP7_75t_SL g71 ( 
.A1(n_46),
.A2(n_64),
.B(n_47),
.Y(n_71)
);

AND2x2_ASAP7_75t_SL g72 ( 
.A(n_48),
.B(n_0),
.Y(n_72)
);

NAND3xp33_ASAP7_75t_L g73 ( 
.A(n_66),
.B(n_0),
.C(n_1),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_46),
.B(n_1),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_45),
.Y(n_75)
);

BUFx10_ASAP7_75t_L g76 ( 
.A(n_52),
.Y(n_76)
);

NAND2xp33_ASAP7_75t_SL g77 ( 
.A(n_50),
.B(n_2),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_42),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_43),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_44),
.Y(n_80)
);

INVx2_ASAP7_75t_SL g81 ( 
.A(n_56),
.Y(n_81)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_49),
.Y(n_82)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_51),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_53),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_47),
.B(n_3),
.Y(n_85)
);

INVx8_ASAP7_75t_L g86 ( 
.A(n_57),
.Y(n_86)
);

NAND3xp33_ASAP7_75t_L g87 ( 
.A(n_67),
.B(n_5),
.C(n_6),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_54),
.Y(n_88)
);

AND2x6_ASAP7_75t_L g89 ( 
.A(n_74),
.B(n_62),
.Y(n_89)
);

NOR2x1p5_ASAP7_75t_L g90 ( 
.A(n_87),
.B(n_45),
.Y(n_90)
);

OR2x2_ASAP7_75t_L g91 ( 
.A(n_81),
.B(n_65),
.Y(n_91)
);

BUFx2_ASAP7_75t_L g92 ( 
.A(n_75),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_78),
.B(n_67),
.Y(n_93)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_76),
.B(n_63),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_79),
.B(n_61),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_71),
.B(n_59),
.Y(n_96)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_69),
.Y(n_97)
);

AND2x4_ASAP7_75t_L g98 ( 
.A(n_80),
.B(n_58),
.Y(n_98)
);

AO22x1_ASAP7_75t_L g99 ( 
.A1(n_74),
.A2(n_68),
.B1(n_63),
.B2(n_50),
.Y(n_99)
);

NOR2x1_ASAP7_75t_R g100 ( 
.A(n_85),
.B(n_72),
.Y(n_100)
);

NAND2x2_ASAP7_75t_L g101 ( 
.A(n_85),
.B(n_6),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_73),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_102)
);

INVx1_ASAP7_75t_SL g103 ( 
.A(n_94),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_89),
.B(n_86),
.Y(n_104)
);

AO21x1_ASAP7_75t_L g105 ( 
.A1(n_96),
.A2(n_77),
.B(n_84),
.Y(n_105)
);

OA21x2_ASAP7_75t_L g106 ( 
.A1(n_95),
.A2(n_93),
.B(n_82),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_L g107 ( 
.A1(n_93),
.A2(n_83),
.B(n_87),
.Y(n_107)
);

AND2x4_ASAP7_75t_L g108 ( 
.A(n_90),
.B(n_73),
.Y(n_108)
);

CKINVDCx16_ASAP7_75t_R g109 ( 
.A(n_92),
.Y(n_109)
);

OAI21x1_ASAP7_75t_L g110 ( 
.A1(n_95),
.A2(n_70),
.B(n_88),
.Y(n_110)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_97),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_91),
.A2(n_86),
.B1(n_88),
.B2(n_76),
.Y(n_112)
);

AND2x4_ASAP7_75t_L g113 ( 
.A(n_98),
.B(n_88),
.Y(n_113)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_98),
.Y(n_114)
);

NAND2x1_ASAP7_75t_L g115 ( 
.A(n_106),
.B(n_89),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_111),
.Y(n_116)
);

CKINVDCx5p33_ASAP7_75t_R g117 ( 
.A(n_109),
.Y(n_117)
);

AOI21x1_ASAP7_75t_SL g118 ( 
.A1(n_104),
.A2(n_101),
.B(n_89),
.Y(n_118)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_110),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_111),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_106),
.B(n_89),
.Y(n_121)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_110),
.Y(n_122)
);

AOI221x1_ASAP7_75t_SL g123 ( 
.A1(n_108),
.A2(n_100),
.B1(n_99),
.B2(n_102),
.C(n_86),
.Y(n_123)
);

INVx2_ASAP7_75t_SL g124 ( 
.A(n_113),
.Y(n_124)
);

AND2x2_ASAP7_75t_L g125 ( 
.A(n_117),
.B(n_109),
.Y(n_125)
);

HB1xp67_ASAP7_75t_L g126 ( 
.A(n_117),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_124),
.A2(n_108),
.B1(n_106),
.B2(n_114),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_121),
.B(n_106),
.Y(n_128)
);

AND2x2_ASAP7_75t_L g129 ( 
.A(n_124),
.B(n_103),
.Y(n_129)
);

HB1xp67_ASAP7_75t_L g130 ( 
.A(n_116),
.Y(n_130)
);

AND2x2_ASAP7_75t_L g131 ( 
.A(n_120),
.B(n_114),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_115),
.Y(n_132)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_119),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_119),
.Y(n_134)
);

BUFx2_ASAP7_75t_L g135 ( 
.A(n_125),
.Y(n_135)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_131),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_127),
.B(n_108),
.Y(n_137)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_130),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_129),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_127),
.Y(n_140)
);

NOR2x1_ASAP7_75t_L g141 ( 
.A(n_138),
.B(n_113),
.Y(n_141)
);

BUFx2_ASAP7_75t_L g142 ( 
.A(n_135),
.Y(n_142)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_136),
.Y(n_143)
);

OR2x2_ASAP7_75t_L g144 ( 
.A(n_139),
.B(n_126),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_141),
.A2(n_108),
.B1(n_112),
.B2(n_137),
.Y(n_145)
);

AOI221xp5_ASAP7_75t_SL g146 ( 
.A1(n_142),
.A2(n_102),
.B1(n_107),
.B2(n_137),
.C(n_123),
.Y(n_146)
);

NAND2x1p5_ASAP7_75t_L g147 ( 
.A(n_144),
.B(n_113),
.Y(n_147)
);

AOI21xp33_ASAP7_75t_L g148 ( 
.A1(n_146),
.A2(n_140),
.B(n_143),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_145),
.A2(n_105),
.B1(n_113),
.B2(n_132),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_147),
.A2(n_105),
.B1(n_132),
.B2(n_128),
.Y(n_150)
);

OAI221xp5_ASAP7_75t_L g151 ( 
.A1(n_149),
.A2(n_118),
.B1(n_132),
.B2(n_134),
.C(n_133),
.Y(n_151)
);

NOR4xp75_ASAP7_75t_L g152 ( 
.A(n_151),
.B(n_148),
.C(n_150),
.D(n_128),
.Y(n_152)
);

AOI322xp5_ASAP7_75t_L g153 ( 
.A1(n_152),
.A2(n_122),
.A3(n_20),
.B1(n_23),
.B2(n_24),
.C1(n_25),
.C2(n_18),
.Y(n_153)
);

NOR3xp33_ASAP7_75t_L g154 ( 
.A(n_153),
.B(n_122),
.C(n_28),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_154),
.Y(n_155)
);

OR2x2_ASAP7_75t_L g156 ( 
.A(n_155),
.B(n_26),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_156),
.A2(n_33),
.B1(n_35),
.B2(n_36),
.Y(n_157)
);


endmodule