module fake_jpeg_4586_n_284 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_284);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_284;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_14;
wire n_182;
wire n_19;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_272;
wire n_280;
wire n_171;
wire n_263;
wire n_119;
wire n_23;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_8),
.Y(n_13)
);

BUFx10_ASAP7_75t_L g14 ( 
.A(n_0),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

INVx3_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_0),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

INVx8_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_5),
.Y(n_26)
);

INVx5_ASAP7_75t_L g27 ( 
.A(n_22),
.Y(n_27)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_27),
.Y(n_41)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_20),
.Y(n_28)
);

INVx5_ASAP7_75t_L g42 ( 
.A(n_28),
.Y(n_42)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_20),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_19),
.Y(n_30)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_30),
.Y(n_43)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_22),
.Y(n_31)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_31),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_22),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_32),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_16),
.B(n_6),
.Y(n_33)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_33),
.Y(n_39)
);

INVx3_ASAP7_75t_SL g34 ( 
.A(n_22),
.Y(n_34)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_15),
.Y(n_35)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_35),
.Y(n_40)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_19),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_L g37 ( 
.A1(n_36),
.A2(n_28),
.B1(n_25),
.B2(n_31),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_37),
.B(n_35),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_L g44 ( 
.A1(n_28),
.A2(n_25),
.B1(n_17),
.B2(n_26),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_44),
.A2(n_25),
.B1(n_17),
.B2(n_26),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_30),
.A2(n_25),
.B1(n_17),
.B2(n_18),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_48),
.A2(n_16),
.B1(n_24),
.B2(n_13),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_42),
.Y(n_49)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_49),
.Y(n_76)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_42),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_50),
.B(n_52),
.Y(n_83)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_45),
.Y(n_51)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_51),
.Y(n_68)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_42),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_53),
.B(n_54),
.Y(n_73)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_48),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_41),
.B(n_33),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_55),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_39),
.A2(n_31),
.B1(n_17),
.B2(n_34),
.Y(n_56)
);

INVxp67_ASAP7_75t_L g80 ( 
.A(n_56),
.Y(n_80)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

INVx3_ASAP7_75t_SL g78 ( 
.A(n_57),
.Y(n_78)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

INVx1_ASAP7_75t_SL g72 ( 
.A(n_58),
.Y(n_72)
);

INVx2_ASAP7_75t_SL g59 ( 
.A(n_40),
.Y(n_59)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_59),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_L g60 ( 
.A1(n_39),
.A2(n_36),
.B1(n_30),
.B2(n_27),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_60),
.A2(n_65),
.B1(n_37),
.B2(n_64),
.Y(n_82)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_40),
.Y(n_61)
);

INVx4_ASAP7_75t_SL g81 ( 
.A(n_61),
.Y(n_81)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_62),
.Y(n_69)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_40),
.Y(n_63)
);

BUFx2_ASAP7_75t_L g74 ( 
.A(n_63),
.Y(n_74)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_44),
.Y(n_64)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_64),
.Y(n_75)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_49),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_67),
.B(n_45),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_SL g70 ( 
.A1(n_54),
.A2(n_34),
.B(n_39),
.Y(n_70)
);

XOR2xp5_ASAP7_75t_L g99 ( 
.A(n_70),
.B(n_47),
.Y(n_99)
);

OR2x2_ASAP7_75t_L g77 ( 
.A(n_65),
.B(n_34),
.Y(n_77)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_77),
.B(n_27),
.Y(n_96)
);

BUFx2_ASAP7_75t_L g79 ( 
.A(n_51),
.Y(n_79)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_79),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_82),
.A2(n_73),
.B1(n_69),
.B2(n_71),
.Y(n_90)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_74),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_85),
.B(n_91),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_73),
.A2(n_53),
.B1(n_58),
.B2(n_57),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_86),
.A2(n_93),
.B1(n_94),
.B2(n_69),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_76),
.A2(n_52),
.B1(n_47),
.B2(n_46),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_87),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_76),
.A2(n_47),
.B1(n_46),
.B2(n_50),
.Y(n_88)
);

AOI21xp5_ASAP7_75t_L g117 ( 
.A1(n_88),
.A2(n_78),
.B(n_35),
.Y(n_117)
);

INVxp33_ASAP7_75t_L g116 ( 
.A(n_89),
.Y(n_116)
);

CKINVDCx16_ASAP7_75t_R g111 ( 
.A(n_90),
.Y(n_111)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_83),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_74),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_92),
.B(n_95),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_82),
.A2(n_43),
.B1(n_36),
.B2(n_46),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_70),
.A2(n_75),
.B1(n_80),
.B2(n_77),
.Y(n_94)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_83),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_96),
.B(n_97),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_71),
.B(n_61),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_81),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_98),
.B(n_101),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_99),
.B(n_96),
.Y(n_115)
);

OAI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_77),
.A2(n_43),
.B1(n_63),
.B2(n_29),
.Y(n_100)
);

OAI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_100),
.A2(n_78),
.B1(n_67),
.B2(n_66),
.Y(n_110)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_81),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_81),
.Y(n_102)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_102),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_103),
.A2(n_123),
.B1(n_59),
.B2(n_101),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_SL g104 ( 
.A1(n_99),
.A2(n_75),
.B(n_66),
.Y(n_104)
);

AOI21xp5_ASAP7_75t_L g145 ( 
.A1(n_104),
.A2(n_117),
.B(n_118),
.Y(n_145)
);

INVx6_ASAP7_75t_L g105 ( 
.A(n_84),
.Y(n_105)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_105),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_94),
.A2(n_43),
.B1(n_59),
.B2(n_76),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_106),
.A2(n_84),
.B1(n_68),
.B2(n_72),
.Y(n_142)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_97),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_109),
.B(n_102),
.Y(n_129)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_110),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_L g143 ( 
.A(n_115),
.B(n_121),
.Y(n_143)
);

AOI21xp5_ASAP7_75t_L g118 ( 
.A1(n_96),
.A2(n_100),
.B(n_91),
.Y(n_118)
);

CKINVDCx16_ASAP7_75t_R g120 ( 
.A(n_89),
.Y(n_120)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_120),
.Y(n_131)
);

MAJx2_ASAP7_75t_L g121 ( 
.A(n_90),
.B(n_78),
.C(n_32),
.Y(n_121)
);

OR2x2_ASAP7_75t_L g122 ( 
.A(n_86),
.B(n_18),
.Y(n_122)
);

AO22x1_ASAP7_75t_SL g144 ( 
.A1(n_122),
.A2(n_32),
.B1(n_15),
.B2(n_45),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_L g123 ( 
.A1(n_93),
.A2(n_29),
.B1(n_49),
.B2(n_68),
.Y(n_123)
);

NOR2xp67_ASAP7_75t_R g125 ( 
.A(n_122),
.B(n_95),
.Y(n_125)
);

FAx1_ASAP7_75t_L g159 ( 
.A(n_125),
.B(n_144),
.CI(n_110),
.CON(n_159),
.SN(n_159)
);

CKINVDCx16_ASAP7_75t_R g157 ( 
.A(n_127),
.Y(n_157)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_119),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_128),
.B(n_136),
.Y(n_161)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_129),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_109),
.B(n_98),
.Y(n_130)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_130),
.Y(n_156)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_119),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_132),
.B(n_134),
.Y(n_151)
);

OAI32xp33_ASAP7_75t_L g133 ( 
.A1(n_111),
.A2(n_24),
.A3(n_16),
.B1(n_32),
.B2(n_15),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_133),
.Y(n_154)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_113),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_111),
.A2(n_92),
.B1(n_72),
.B2(n_85),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_135),
.A2(n_117),
.B1(n_120),
.B2(n_107),
.Y(n_147)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_113),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_106),
.A2(n_118),
.B1(n_103),
.B2(n_122),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_137),
.A2(n_142),
.B1(n_108),
.B2(n_106),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_112),
.B(n_74),
.Y(n_138)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_138),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_108),
.A2(n_121),
.B1(n_122),
.B2(n_118),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g158 ( 
.A(n_139),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_L g140 ( 
.A1(n_115),
.A2(n_112),
.B(n_104),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g152 ( 
.A(n_140),
.B(n_141),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_L g141 ( 
.A1(n_115),
.A2(n_13),
.B(n_26),
.Y(n_141)
);

XOR2x2_ASAP7_75t_L g146 ( 
.A(n_104),
.B(n_121),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_SL g168 ( 
.A(n_146),
.B(n_20),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_147),
.A2(n_163),
.B1(n_144),
.B2(n_125),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_148),
.A2(n_133),
.B1(n_23),
.B2(n_15),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_146),
.A2(n_103),
.B1(n_117),
.B2(n_107),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_149),
.A2(n_169),
.B1(n_14),
.B2(n_23),
.Y(n_192)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_126),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_153),
.B(n_155),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_128),
.B(n_114),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_159),
.B(n_162),
.Y(n_172)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_129),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_124),
.A2(n_123),
.B1(n_114),
.B2(n_116),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_142),
.B(n_105),
.Y(n_164)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_164),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_130),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_165),
.B(n_170),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_136),
.B(n_105),
.Y(n_166)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_166),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_140),
.B(n_45),
.C(n_38),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_167),
.B(n_135),
.C(n_145),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_168),
.B(n_14),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_124),
.A2(n_18),
.B1(n_13),
.B2(n_24),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_138),
.Y(n_170)
);

INVxp33_ASAP7_75t_L g174 ( 
.A(n_161),
.Y(n_174)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_174),
.Y(n_195)
);

CKINVDCx16_ASAP7_75t_R g175 ( 
.A(n_151),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_175),
.B(n_171),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g176 ( 
.A(n_149),
.B(n_143),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_176),
.B(n_187),
.Y(n_194)
);

BUFx2_ASAP7_75t_L g177 ( 
.A(n_153),
.Y(n_177)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_177),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_L g193 ( 
.A1(n_178),
.A2(n_181),
.B(n_189),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_179),
.B(n_180),
.C(n_182),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_168),
.B(n_145),
.C(n_143),
.Y(n_180)
);

AOI21xp5_ASAP7_75t_L g181 ( 
.A1(n_158),
.A2(n_139),
.B(n_144),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_160),
.B(n_141),
.C(n_131),
.Y(n_182)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_183),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_157),
.A2(n_68),
.B1(n_79),
.B2(n_23),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_186),
.A2(n_148),
.B1(n_150),
.B2(n_156),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_152),
.B(n_79),
.Y(n_187)
);

XOR2x2_ASAP7_75t_L g188 ( 
.A(n_158),
.B(n_20),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_SL g206 ( 
.A(n_188),
.B(n_169),
.Y(n_206)
);

AOI21xp5_ASAP7_75t_L g189 ( 
.A1(n_165),
.A2(n_19),
.B(n_1),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_190),
.B(n_191),
.Y(n_210)
);

AOI21xp5_ASAP7_75t_L g191 ( 
.A1(n_160),
.A2(n_19),
.B(n_1),
.Y(n_191)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_192),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_176),
.B(n_152),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_197),
.B(n_206),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_187),
.B(n_167),
.C(n_170),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_199),
.B(n_200),
.C(n_207),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_180),
.B(n_150),
.C(n_162),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_185),
.B(n_156),
.Y(n_201)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_201),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_204),
.B(n_209),
.Y(n_215)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_173),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_205),
.B(n_208),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_179),
.B(n_154),
.C(n_159),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_173),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_SL g209 ( 
.A(n_174),
.B(n_154),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_182),
.B(n_159),
.C(n_21),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_211),
.B(n_184),
.C(n_172),
.Y(n_214)
);

AOI21xp5_ASAP7_75t_L g223 ( 
.A1(n_212),
.A2(n_177),
.B(n_190),
.Y(n_223)
);

AOI21xp5_ASAP7_75t_L g239 ( 
.A1(n_214),
.A2(n_220),
.B(n_223),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_200),
.B(n_171),
.C(n_172),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_216),
.B(n_219),
.C(n_221),
.Y(n_236)
);

BUFx24_ASAP7_75t_SL g217 ( 
.A(n_197),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_217),
.B(n_21),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_203),
.A2(n_178),
.B1(n_188),
.B2(n_181),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_218),
.A2(n_227),
.B1(n_229),
.B2(n_193),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_196),
.B(n_199),
.C(n_194),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_L g220 ( 
.A1(n_196),
.A2(n_189),
.B(n_191),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_194),
.B(n_192),
.C(n_186),
.Y(n_221)
);

HB1xp67_ASAP7_75t_L g224 ( 
.A(n_198),
.Y(n_224)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_224),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_207),
.B(n_21),
.C(n_14),
.Y(n_226)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_226),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_202),
.A2(n_23),
.B1(n_8),
.B2(n_12),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_211),
.A2(n_193),
.B1(n_204),
.B2(n_195),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_230),
.B(n_7),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_215),
.A2(n_198),
.B1(n_206),
.B2(n_210),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_233),
.B(n_234),
.C(n_237),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_222),
.B(n_210),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_228),
.Y(n_235)
);

AOI21xp5_ASAP7_75t_L g246 ( 
.A1(n_235),
.A2(n_38),
.B(n_7),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_214),
.A2(n_225),
.B1(n_221),
.B2(n_216),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_238),
.B(n_240),
.C(n_241),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_226),
.A2(n_8),
.B1(n_9),
.B2(n_12),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_222),
.B(n_38),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_219),
.B(n_14),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_SL g247 ( 
.A(n_242),
.B(n_14),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_213),
.B(n_38),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g255 ( 
.A(n_243),
.B(n_5),
.Y(n_255)
);

OAI21xp5_ASAP7_75t_SL g244 ( 
.A1(n_236),
.A2(n_213),
.B(n_8),
.Y(n_244)
);

AOI21xp5_ASAP7_75t_L g262 ( 
.A1(n_244),
.A2(n_246),
.B(n_247),
.Y(n_262)
);

HB1xp67_ASAP7_75t_L g249 ( 
.A(n_231),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_249),
.B(n_252),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_L g259 ( 
.A1(n_250),
.A2(n_251),
.B1(n_254),
.B2(n_240),
.Y(n_259)
);

AOI21xp5_ASAP7_75t_SL g251 ( 
.A1(n_232),
.A2(n_14),
.B(n_7),
.Y(n_251)
);

OAI221xp5_ASAP7_75t_L g252 ( 
.A1(n_241),
.A2(n_21),
.B1(n_14),
.B2(n_6),
.C(n_10),
.Y(n_252)
);

INVx1_ASAP7_75t_SL g253 ( 
.A(n_243),
.Y(n_253)
);

OR2x2_ASAP7_75t_L g263 ( 
.A(n_253),
.B(n_9),
.Y(n_263)
);

AOI21xp5_ASAP7_75t_L g254 ( 
.A1(n_239),
.A2(n_21),
.B(n_6),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_255),
.B(n_4),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_SL g256 ( 
.A(n_245),
.B(n_236),
.Y(n_256)
);

AOI21xp5_ASAP7_75t_L g269 ( 
.A1(n_256),
.A2(n_264),
.B(n_4),
.Y(n_269)
);

INVxp67_ASAP7_75t_L g258 ( 
.A(n_255),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_258),
.B(n_259),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_L g260 ( 
.A1(n_248),
.A2(n_242),
.B1(n_9),
.B2(n_10),
.Y(n_260)
);

INVxp67_ASAP7_75t_L g267 ( 
.A(n_260),
.Y(n_267)
);

OA21x2_ASAP7_75t_SL g261 ( 
.A1(n_249),
.A2(n_21),
.B(n_5),
.Y(n_261)
);

NOR2xp67_ASAP7_75t_SL g272 ( 
.A(n_261),
.B(n_10),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_L g273 ( 
.A1(n_263),
.A2(n_11),
.B1(n_1),
.B2(n_2),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_249),
.B(n_9),
.Y(n_264)
);

OAI321xp33_ASAP7_75t_L g271 ( 
.A1(n_265),
.A2(n_10),
.A3(n_11),
.B1(n_12),
.B2(n_3),
.C(n_0),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_SL g268 ( 
.A(n_262),
.B(n_21),
.Y(n_268)
);

AOI21xp5_ASAP7_75t_L g278 ( 
.A1(n_268),
.A2(n_270),
.B(n_271),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_269),
.Y(n_277)
);

AOI21xp5_ASAP7_75t_L g270 ( 
.A1(n_257),
.A2(n_4),
.B(n_11),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_272),
.B(n_273),
.Y(n_276)
);

NOR3xp33_ASAP7_75t_SL g274 ( 
.A(n_266),
.B(n_257),
.C(n_2),
.Y(n_274)
);

AOI21x1_ASAP7_75t_L g279 ( 
.A1(n_274),
.A2(n_275),
.B(n_2),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_267),
.B(n_0),
.Y(n_275)
);

AO21x1_ASAP7_75t_L g281 ( 
.A1(n_279),
.A2(n_280),
.B(n_277),
.Y(n_281)
);

AOI21xp5_ASAP7_75t_L g280 ( 
.A1(n_276),
.A2(n_2),
.B(n_3),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_281),
.B(n_278),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_282),
.B(n_3),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_283),
.B(n_3),
.Y(n_284)
);


endmodule