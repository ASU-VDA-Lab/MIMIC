module fake_jpeg_19640_n_323 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_323);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_323;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_13;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_11;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_12;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx12f_ASAP7_75t_L g11 ( 
.A(n_4),
.Y(n_11)
);

INVx2_ASAP7_75t_L g12 ( 
.A(n_3),
.Y(n_12)
);

INVx11_ASAP7_75t_SL g13 ( 
.A(n_1),
.Y(n_13)
);

BUFx12f_ASAP7_75t_L g14 ( 
.A(n_4),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_6),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_0),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_6),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_4),
.Y(n_21)
);

INVxp67_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_1),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_24),
.Y(n_35)
);

CKINVDCx14_ASAP7_75t_R g25 ( 
.A(n_13),
.Y(n_25)
);

CKINVDCx14_ASAP7_75t_R g42 ( 
.A(n_25),
.Y(n_42)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_26),
.Y(n_39)
);

INVx5_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_27),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_15),
.B(n_10),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_SL g36 ( 
.A(n_28),
.B(n_32),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

BUFx2_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_30),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_18),
.Y(n_31)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_31),
.Y(n_43)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_18),
.Y(n_32)
);

INVx4_ASAP7_75t_SL g33 ( 
.A(n_11),
.Y(n_33)
);

AOI22xp33_ASAP7_75t_SL g44 ( 
.A1(n_33),
.A2(n_34),
.B1(n_12),
.B2(n_20),
.Y(n_44)
);

BUFx12_ASAP7_75t_L g34 ( 
.A(n_11),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_31),
.B(n_14),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_37),
.B(n_29),
.Y(n_47)
);

CKINVDCx16_ASAP7_75t_R g52 ( 
.A(n_44),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_SL g45 ( 
.A1(n_30),
.A2(n_12),
.B1(n_20),
.B2(n_16),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g48 ( 
.A1(n_45),
.A2(n_33),
.B1(n_25),
.B2(n_26),
.Y(n_48)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_41),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_46),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_47),
.B(n_54),
.Y(n_64)
);

AOI21xp5_ASAP7_75t_L g72 ( 
.A1(n_48),
.A2(n_44),
.B(n_34),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_36),
.B(n_28),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_49),
.B(n_60),
.Y(n_61)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_40),
.Y(n_50)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_50),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g51 ( 
.A1(n_37),
.A2(n_12),
.B1(n_33),
.B2(n_26),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_51),
.A2(n_33),
.B1(n_43),
.B2(n_37),
.Y(n_69)
);

INVx11_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_53),
.A2(n_59),
.B1(n_43),
.B2(n_39),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_37),
.B(n_29),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g73 ( 
.A(n_55),
.Y(n_73)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_56),
.Y(n_79)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_45),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_57),
.B(n_58),
.Y(n_70)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_45),
.Y(n_58)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_40),
.Y(n_59)
);

INVx5_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

INVx6_ASAP7_75t_SL g62 ( 
.A(n_53),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_62),
.B(n_66),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_63),
.Y(n_97)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_46),
.Y(n_65)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_65),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_49),
.B(n_36),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_L g67 ( 
.A1(n_57),
.A2(n_36),
.B1(n_43),
.B2(n_45),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_L g90 ( 
.A1(n_67),
.A2(n_51),
.B1(n_56),
.B2(n_46),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_52),
.A2(n_45),
.B1(n_44),
.B2(n_27),
.Y(n_68)
);

OAI21xp5_ASAP7_75t_L g87 ( 
.A1(n_68),
.A2(n_48),
.B(n_22),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_69),
.A2(n_72),
.B1(n_74),
.B2(n_56),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_47),
.B(n_41),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_71),
.B(n_77),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_57),
.A2(n_43),
.B1(n_41),
.B2(n_27),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_47),
.B(n_42),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_58),
.A2(n_43),
.B1(n_39),
.B2(n_42),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_78),
.A2(n_72),
.B1(n_74),
.B2(n_63),
.Y(n_95)
);

XOR2xp5_ASAP7_75t_L g80 ( 
.A(n_64),
.B(n_54),
.Y(n_80)
);

XNOR2xp5_ASAP7_75t_L g116 ( 
.A(n_80),
.B(n_61),
.Y(n_116)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_79),
.Y(n_81)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_81),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_75),
.A2(n_52),
.B1(n_58),
.B2(n_59),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_82),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_75),
.A2(n_59),
.B1(n_60),
.B2(n_50),
.Y(n_83)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_83),
.Y(n_119)
);

AOI21xp5_ASAP7_75t_L g84 ( 
.A1(n_70),
.A2(n_48),
.B(n_54),
.Y(n_84)
);

OAI21xp5_ASAP7_75t_SL g105 ( 
.A1(n_84),
.A2(n_88),
.B(n_89),
.Y(n_105)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_79),
.Y(n_86)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_86),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_87),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_L g88 ( 
.A1(n_70),
.A2(n_23),
.B(n_19),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_75),
.A2(n_59),
.B1(n_60),
.B2(n_50),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_90),
.A2(n_93),
.B1(n_95),
.B2(n_78),
.Y(n_100)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_73),
.Y(n_94)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_94),
.Y(n_114)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_76),
.Y(n_96)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_96),
.Y(n_108)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_76),
.Y(n_98)
);

INVx1_ASAP7_75t_SL g112 ( 
.A(n_98),
.Y(n_112)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_76),
.Y(n_99)
);

CKINVDCx16_ASAP7_75t_R g115 ( 
.A(n_99),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_100),
.A2(n_101),
.B1(n_111),
.B2(n_122),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_95),
.A2(n_68),
.B1(n_72),
.B2(n_67),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_92),
.B(n_64),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_103),
.B(n_104),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_92),
.B(n_71),
.Y(n_104)
);

XOR2xp5_ASAP7_75t_L g106 ( 
.A(n_80),
.B(n_66),
.Y(n_106)
);

XNOR2xp5_ASAP7_75t_SL g160 ( 
.A(n_106),
.B(n_116),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_81),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_110),
.B(n_113),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_93),
.A2(n_68),
.B1(n_61),
.B2(n_77),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_86),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_85),
.B(n_84),
.Y(n_117)
);

CKINVDCx14_ASAP7_75t_R g145 ( 
.A(n_117),
.Y(n_145)
);

CKINVDCx16_ASAP7_75t_R g118 ( 
.A(n_96),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_118),
.B(n_120),
.Y(n_136)
);

CKINVDCx16_ASAP7_75t_R g120 ( 
.A(n_98),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_82),
.A2(n_69),
.B1(n_74),
.B2(n_55),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_87),
.A2(n_69),
.B1(n_55),
.B2(n_65),
.Y(n_123)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_123),
.Y(n_159)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_91),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_124),
.B(n_73),
.Y(n_151)
);

OR2x6_ASAP7_75t_L g125 ( 
.A(n_90),
.B(n_34),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_SL g148 ( 
.A1(n_125),
.A2(n_38),
.B(n_62),
.Y(n_148)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_111),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_126),
.B(n_132),
.Y(n_171)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_102),
.Y(n_128)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_128),
.Y(n_161)
);

AOI21xp5_ASAP7_75t_L g130 ( 
.A1(n_109),
.A2(n_97),
.B(n_85),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_L g169 ( 
.A1(n_130),
.A2(n_142),
.B(n_150),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_106),
.B(n_29),
.C(n_88),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_131),
.B(n_138),
.C(n_146),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_102),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_100),
.A2(n_125),
.B1(n_109),
.B2(n_101),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_133),
.A2(n_134),
.B1(n_119),
.B2(n_122),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_125),
.A2(n_83),
.B1(n_99),
.B2(n_91),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_107),
.Y(n_135)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_135),
.Y(n_167)
);

OAI22x1_ASAP7_75t_L g137 ( 
.A1(n_125),
.A2(n_38),
.B1(n_62),
.B2(n_34),
.Y(n_137)
);

OAI22x1_ASAP7_75t_L g181 ( 
.A1(n_137),
.A2(n_38),
.B1(n_32),
.B2(n_35),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_116),
.B(n_29),
.C(n_91),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_L g139 ( 
.A(n_103),
.B(n_34),
.Y(n_139)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_139),
.B(n_157),
.Y(n_174)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_107),
.Y(n_141)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_141),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_125),
.A2(n_94),
.B1(n_39),
.B2(n_42),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_108),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_143),
.B(n_144),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_108),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_104),
.B(n_39),
.C(n_73),
.Y(n_146)
);

HB1xp67_ASAP7_75t_L g147 ( 
.A(n_105),
.Y(n_147)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_147),
.Y(n_172)
);

AO22x1_ASAP7_75t_L g189 ( 
.A1(n_148),
.A2(n_35),
.B1(n_24),
.B2(n_14),
.Y(n_189)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_114),
.Y(n_149)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_149),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_SL g150 ( 
.A1(n_121),
.A2(n_19),
.B(n_21),
.Y(n_150)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_151),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_SL g152 ( 
.A1(n_121),
.A2(n_21),
.B(n_15),
.Y(n_152)
);

INVxp67_ASAP7_75t_L g186 ( 
.A(n_152),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_115),
.B(n_73),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_153),
.B(n_154),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_114),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_124),
.B(n_73),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_155),
.B(n_156),
.Y(n_188)
);

CKINVDCx16_ASAP7_75t_R g156 ( 
.A(n_105),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_125),
.A2(n_39),
.B1(n_20),
.B2(n_16),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_123),
.B(n_76),
.C(n_40),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_158),
.B(n_31),
.C(n_119),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_163),
.A2(n_170),
.B1(n_176),
.B2(n_185),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_164),
.B(n_167),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_160),
.B(n_40),
.C(n_112),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_165),
.B(n_183),
.C(n_184),
.Y(n_193)
);

OAI21xp33_ASAP7_75t_L g166 ( 
.A1(n_156),
.A2(n_112),
.B(n_23),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_SL g199 ( 
.A1(n_166),
.A2(n_181),
.B(n_189),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_129),
.A2(n_53),
.B1(n_31),
.B2(n_16),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_127),
.B(n_35),
.Y(n_175)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_175),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_129),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_160),
.B(n_38),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_178),
.B(n_154),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_126),
.A2(n_17),
.B1(n_32),
.B2(n_18),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_179),
.A2(n_134),
.B1(n_144),
.B2(n_143),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_140),
.B(n_17),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_182),
.B(n_17),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_138),
.B(n_14),
.C(n_38),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_131),
.B(n_14),
.C(n_38),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_133),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_185)
);

INVxp67_ASAP7_75t_SL g190 ( 
.A(n_137),
.Y(n_190)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_190),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_177),
.B(n_140),
.Y(n_191)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_191),
.Y(n_225)
);

INVxp67_ASAP7_75t_L g192 ( 
.A(n_187),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_192),
.B(n_194),
.Y(n_222)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_181),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_165),
.B(n_146),
.C(n_139),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_195),
.B(n_202),
.C(n_205),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_171),
.B(n_132),
.Y(n_197)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_197),
.Y(n_231)
);

INVxp67_ASAP7_75t_L g201 ( 
.A(n_188),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_201),
.B(n_209),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_162),
.B(n_145),
.C(n_158),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g223 ( 
.A1(n_203),
.A2(n_170),
.B1(n_185),
.B2(n_176),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_161),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_204),
.B(n_212),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_162),
.B(n_159),
.C(n_141),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_164),
.A2(n_159),
.B1(n_130),
.B2(n_135),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_206),
.B(n_210),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_178),
.B(n_128),
.C(n_142),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_207),
.B(n_211),
.C(n_169),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_180),
.B(n_136),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_208),
.Y(n_228)
);

AO22x2_ASAP7_75t_SL g209 ( 
.A1(n_163),
.A2(n_148),
.B1(n_157),
.B2(n_152),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_SL g210 ( 
.A(n_174),
.B(n_150),
.Y(n_210)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_168),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_213),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_214),
.B(n_149),
.Y(n_216)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_173),
.Y(n_215)
);

CKINVDCx16_ASAP7_75t_R g232 ( 
.A(n_215),
.Y(n_232)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_216),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_191),
.B(n_172),
.Y(n_218)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_218),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_196),
.B(n_179),
.Y(n_220)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_220),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_223),
.A2(n_227),
.B1(n_210),
.B2(n_209),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_205),
.B(n_174),
.Y(n_226)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_226),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_L g227 ( 
.A1(n_203),
.A2(n_169),
.B1(n_186),
.B2(n_184),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_229),
.B(n_193),
.Y(n_245)
);

AOI21xp5_ASAP7_75t_L g230 ( 
.A1(n_200),
.A2(n_186),
.B(n_166),
.Y(n_230)
);

CKINVDCx16_ASAP7_75t_R g254 ( 
.A(n_230),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_197),
.B(n_183),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_SL g255 ( 
.A(n_233),
.B(n_0),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_198),
.A2(n_189),
.B1(n_1),
.B2(n_2),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g248 ( 
.A1(n_234),
.A2(n_237),
.B1(n_207),
.B2(n_206),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_192),
.B(n_189),
.Y(n_235)
);

AOI21xp5_ASAP7_75t_L g246 ( 
.A1(n_235),
.A2(n_238),
.B(n_199),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_198),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_201),
.B(n_18),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_219),
.B(n_202),
.C(n_193),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_239),
.B(n_14),
.C(n_4),
.Y(n_272)
);

AND2x2_ASAP7_75t_L g242 ( 
.A(n_227),
.B(n_194),
.Y(n_242)
);

CKINVDCx14_ASAP7_75t_R g270 ( 
.A(n_242),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_243),
.A2(n_222),
.B1(n_237),
.B2(n_221),
.Y(n_262)
);

AOI21xp5_ASAP7_75t_SL g244 ( 
.A1(n_224),
.A2(n_199),
.B(n_209),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_244),
.B(n_246),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_245),
.B(n_253),
.Y(n_265)
);

BUFx6f_ASAP7_75t_L g247 ( 
.A(n_228),
.Y(n_247)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_247),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_248),
.A2(n_223),
.B1(n_236),
.B2(n_238),
.Y(n_263)
);

BUFx6f_ASAP7_75t_L g249 ( 
.A(n_228),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_249),
.B(n_251),
.Y(n_267)
);

AOI21xp5_ASAP7_75t_SL g251 ( 
.A1(n_224),
.A2(n_231),
.B(n_225),
.Y(n_251)
);

AO21x1_ASAP7_75t_L g252 ( 
.A1(n_235),
.A2(n_211),
.B(n_195),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_252),
.B(n_255),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_219),
.B(n_229),
.Y(n_253)
);

OAI21xp5_ASAP7_75t_L g256 ( 
.A1(n_230),
.A2(n_35),
.B(n_24),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_256),
.A2(n_232),
.B1(n_35),
.B2(n_14),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_239),
.B(n_221),
.C(n_231),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_259),
.B(n_261),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_L g261 ( 
.A1(n_240),
.A2(n_222),
.B1(n_225),
.B2(n_234),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_262),
.B(n_268),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_L g285 ( 
.A1(n_263),
.A2(n_271),
.B1(n_247),
.B2(n_5),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_253),
.B(n_217),
.C(n_236),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_264),
.B(n_257),
.Y(n_277)
);

XNOR2x1_ASAP7_75t_L g269 ( 
.A(n_252),
.B(n_232),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_269),
.B(n_270),
.Y(n_280)
);

AOI22xp33_ASAP7_75t_SL g271 ( 
.A1(n_242),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_SL g286 ( 
.A(n_272),
.B(n_245),
.Y(n_286)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_264),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_273),
.B(n_274),
.Y(n_287)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_267),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_263),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_275),
.B(n_276),
.Y(n_288)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_266),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_277),
.B(n_279),
.Y(n_295)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_258),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_280),
.B(n_285),
.Y(n_298)
);

AOI22xp33_ASAP7_75t_SL g281 ( 
.A1(n_269),
.A2(n_244),
.B1(n_254),
.B2(n_250),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_281),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_265),
.B(n_241),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_SL g289 ( 
.A(n_283),
.B(n_265),
.Y(n_289)
);

OAI21xp5_ASAP7_75t_SL g284 ( 
.A1(n_259),
.A2(n_251),
.B(n_249),
.Y(n_284)
);

AOI21xp5_ASAP7_75t_SL g293 ( 
.A1(n_284),
.A2(n_3),
.B(n_5),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_SL g299 ( 
.A(n_286),
.B(n_7),
.Y(n_299)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_289),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_L g290 ( 
.A1(n_282),
.A2(n_260),
.B1(n_272),
.B2(n_268),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_290),
.A2(n_294),
.B1(n_297),
.B2(n_8),
.Y(n_303)
);

INVxp33_ASAP7_75t_L g291 ( 
.A(n_281),
.Y(n_291)
);

AOI21xp33_ASAP7_75t_L g309 ( 
.A1(n_291),
.A2(n_9),
.B(n_10),
.Y(n_309)
);

INVx1_ASAP7_75t_SL g292 ( 
.A(n_284),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_292),
.B(n_296),
.Y(n_304)
);

OAI21xp5_ASAP7_75t_SL g305 ( 
.A1(n_293),
.A2(n_9),
.B(n_10),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_L g294 ( 
.A1(n_280),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_278),
.B(n_5),
.C(n_6),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_L g308 ( 
.A(n_299),
.B(n_9),
.Y(n_308)
);

OA21x2_ASAP7_75t_SL g300 ( 
.A1(n_295),
.A2(n_278),
.B(n_8),
.Y(n_300)
);

OAI21x1_ASAP7_75t_L g310 ( 
.A1(n_300),
.A2(n_308),
.B(n_309),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_287),
.B(n_7),
.C(n_8),
.Y(n_301)
);

XOR2xp5_ASAP7_75t_L g311 ( 
.A(n_301),
.B(n_302),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_SL g302 ( 
.A(n_288),
.B(n_8),
.Y(n_302)
);

CKINVDCx16_ASAP7_75t_R g312 ( 
.A(n_303),
.Y(n_312)
);

INVxp67_ASAP7_75t_L g314 ( 
.A(n_305),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_292),
.B(n_9),
.Y(n_306)
);

BUFx24_ASAP7_75t_SL g313 ( 
.A(n_306),
.Y(n_313)
);

XOR2xp5_ASAP7_75t_L g315 ( 
.A(n_311),
.B(n_304),
.Y(n_315)
);

A2O1A1O1Ixp25_ASAP7_75t_L g318 ( 
.A1(n_315),
.A2(n_316),
.B(n_317),
.C(n_291),
.D(n_310),
.Y(n_318)
);

OAI21xp5_ASAP7_75t_L g316 ( 
.A1(n_314),
.A2(n_293),
.B(n_307),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_312),
.B(n_301),
.Y(n_317)
);

BUFx24_ASAP7_75t_SL g319 ( 
.A(n_318),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_319),
.B(n_302),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_320),
.B(n_308),
.C(n_313),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_321),
.B(n_298),
.C(n_9),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_322),
.B(n_10),
.Y(n_323)
);


endmodule