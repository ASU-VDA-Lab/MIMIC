module real_aes_7732_n_104 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_104);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_104;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_319;
wire n_421;
wire n_555;
wire n_364;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_379;
wire n_374;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_744;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_178;
wire n_409;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_310;
wire n_455;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_449;
wire n_182;
wire n_363;
wire n_417;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_552;
wire n_402;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_542;
wire n_163;
wire n_645;
wire n_557;
wire n_714;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_753;
wire n_741;
wire n_283;
wire n_252;
wire n_314;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_456;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_541;
wire n_166;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_729;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_743;
wire n_105;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g266 ( .A1(n_0), .A2(n_267), .B(n_268), .C(n_271), .Y(n_266) );
NAND2xp5_ASAP7_75t_L g272 ( .A(n_1), .B(n_208), .Y(n_272) );
NAND3xp33_ASAP7_75t_SL g109 ( .A(n_2), .B(n_92), .C(n_110), .Y(n_109) );
INVx1_ASAP7_75t_L g447 ( .A(n_2), .Y(n_447) );
NAND2xp5_ASAP7_75t_SL g244 ( .A(n_3), .B(n_178), .Y(n_244) );
A2O1A1Ixp33_ASAP7_75t_L g476 ( .A1(n_4), .A2(n_148), .B(n_151), .C(n_477), .Y(n_476) );
AOI21xp5_ASAP7_75t_L g516 ( .A1(n_5), .A2(n_168), .B(n_517), .Y(n_516) );
AOI21xp5_ASAP7_75t_L g198 ( .A1(n_6), .A2(n_168), .B(n_199), .Y(n_198) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_7), .B(n_208), .Y(n_523) );
AO21x2_ASAP7_75t_L g187 ( .A1(n_8), .A2(n_135), .B(n_188), .Y(n_187) );
OAI22xp5_ASAP7_75t_SL g739 ( .A1(n_9), .A2(n_740), .B1(n_743), .B2(n_744), .Y(n_739) );
CKINVDCx20_ASAP7_75t_R g744 ( .A(n_9), .Y(n_744) );
AND2x6_ASAP7_75t_L g148 ( .A(n_10), .B(n_149), .Y(n_148) );
A2O1A1Ixp33_ASAP7_75t_L g150 ( .A1(n_11), .A2(n_148), .B(n_151), .C(n_154), .Y(n_150) );
INVx1_ASAP7_75t_L g493 ( .A(n_12), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g107 ( .A(n_13), .B(n_108), .Y(n_107) );
NOR2xp33_ASAP7_75t_L g448 ( .A(n_13), .B(n_41), .Y(n_448) );
OAI22xp5_ASAP7_75t_L g740 ( .A1(n_14), .A2(n_45), .B1(n_741), .B2(n_742), .Y(n_740) );
CKINVDCx20_ASAP7_75t_R g741 ( .A(n_14), .Y(n_741) );
NAND2xp5_ASAP7_75t_SL g479 ( .A(n_15), .B(n_158), .Y(n_479) );
INVx1_ASAP7_75t_L g140 ( .A(n_16), .Y(n_140) );
NAND2xp5_ASAP7_75t_SL g194 ( .A(n_17), .B(n_178), .Y(n_194) );
A2O1A1Ixp33_ASAP7_75t_L g500 ( .A1(n_18), .A2(n_156), .B(n_501), .C(n_503), .Y(n_500) );
NAND2xp5_ASAP7_75t_L g504 ( .A(n_19), .B(n_208), .Y(n_504) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_20), .B(n_232), .Y(n_536) );
A2O1A1Ixp33_ASAP7_75t_L g227 ( .A1(n_21), .A2(n_151), .B(n_195), .C(n_228), .Y(n_227) );
A2O1A1Ixp33_ASAP7_75t_L g509 ( .A1(n_22), .A2(n_160), .B(n_270), .C(n_510), .Y(n_509) );
NAND2xp5_ASAP7_75t_SL g555 ( .A(n_23), .B(n_158), .Y(n_555) );
NAND2xp5_ASAP7_75t_SL g544 ( .A(n_24), .B(n_158), .Y(n_544) );
CKINVDCx16_ASAP7_75t_R g551 ( .A(n_25), .Y(n_551) );
INVx1_ASAP7_75t_L g543 ( .A(n_26), .Y(n_543) );
A2O1A1Ixp33_ASAP7_75t_L g190 ( .A1(n_27), .A2(n_151), .B(n_191), .C(n_195), .Y(n_190) );
BUFx6f_ASAP7_75t_L g147 ( .A(n_28), .Y(n_147) );
CKINVDCx20_ASAP7_75t_R g475 ( .A(n_29), .Y(n_475) );
INVx1_ASAP7_75t_L g534 ( .A(n_30), .Y(n_534) );
AOI21xp5_ASAP7_75t_L g263 ( .A1(n_31), .A2(n_168), .B(n_264), .Y(n_263) );
INVx2_ASAP7_75t_L g146 ( .A(n_32), .Y(n_146) );
A2O1A1Ixp33_ASAP7_75t_L g215 ( .A1(n_33), .A2(n_170), .B(n_181), .C(n_216), .Y(n_215) );
CKINVDCx20_ASAP7_75t_R g482 ( .A(n_34), .Y(n_482) );
A2O1A1Ixp33_ASAP7_75t_L g519 ( .A1(n_35), .A2(n_270), .B(n_520), .C(n_522), .Y(n_519) );
INVxp67_ASAP7_75t_L g535 ( .A(n_36), .Y(n_535) );
OAI22xp5_ASAP7_75t_SL g449 ( .A1(n_37), .A2(n_79), .B1(n_450), .B2(n_451), .Y(n_449) );
INVx1_ASAP7_75t_L g450 ( .A(n_37), .Y(n_450) );
NAND2xp5_ASAP7_75t_L g192 ( .A(n_38), .B(n_193), .Y(n_192) );
CKINVDCx14_ASAP7_75t_R g518 ( .A(n_39), .Y(n_518) );
A2O1A1Ixp33_ASAP7_75t_L g541 ( .A1(n_40), .A2(n_151), .B(n_195), .C(n_542), .Y(n_541) );
INVx1_ASAP7_75t_L g108 ( .A(n_41), .Y(n_108) );
A2O1A1Ixp33_ASAP7_75t_L g490 ( .A1(n_42), .A2(n_271), .B(n_491), .C(n_492), .Y(n_490) );
NAND2xp5_ASAP7_75t_L g225 ( .A(n_43), .B(n_226), .Y(n_225) );
CKINVDCx20_ASAP7_75t_R g163 ( .A(n_44), .Y(n_163) );
INVx1_ASAP7_75t_L g742 ( .A(n_45), .Y(n_742) );
NAND2xp5_ASAP7_75t_L g177 ( .A(n_46), .B(n_178), .Y(n_177) );
NAND2xp5_ASAP7_75t_L g189 ( .A(n_47), .B(n_168), .Y(n_189) );
CKINVDCx20_ASAP7_75t_R g546 ( .A(n_48), .Y(n_546) );
CKINVDCx20_ASAP7_75t_R g531 ( .A(n_49), .Y(n_531) );
A2O1A1Ixp33_ASAP7_75t_L g169 ( .A1(n_50), .A2(n_170), .B(n_172), .C(n_181), .Y(n_169) );
INVx1_ASAP7_75t_L g269 ( .A(n_51), .Y(n_269) );
INVx1_ASAP7_75t_L g173 ( .A(n_52), .Y(n_173) );
AOI222xp33_ASAP7_75t_L g460 ( .A1(n_53), .A2(n_461), .B1(n_735), .B2(n_736), .C1(n_745), .C2(n_748), .Y(n_460) );
INVx1_ASAP7_75t_L g508 ( .A(n_54), .Y(n_508) );
NAND2xp5_ASAP7_75t_L g167 ( .A(n_55), .B(n_168), .Y(n_167) );
OAI22xp5_ASAP7_75t_SL g122 ( .A1(n_56), .A2(n_59), .B1(n_123), .B2(n_124), .Y(n_122) );
CKINVDCx20_ASAP7_75t_R g124 ( .A(n_56), .Y(n_124) );
CKINVDCx20_ASAP7_75t_R g235 ( .A(n_57), .Y(n_235) );
CKINVDCx14_ASAP7_75t_R g489 ( .A(n_58), .Y(n_489) );
CKINVDCx20_ASAP7_75t_R g123 ( .A(n_59), .Y(n_123) );
INVx1_ASAP7_75t_L g149 ( .A(n_60), .Y(n_149) );
NAND2xp5_ASAP7_75t_L g247 ( .A(n_61), .B(n_168), .Y(n_247) );
AOI22xp33_ASAP7_75t_L g104 ( .A1(n_62), .A2(n_105), .B1(n_113), .B2(n_753), .Y(n_104) );
NAND2xp5_ASAP7_75t_L g207 ( .A(n_63), .B(n_208), .Y(n_207) );
A2O1A1Ixp33_ASAP7_75t_L g201 ( .A1(n_64), .A2(n_202), .B(n_204), .C(n_206), .Y(n_201) );
INVx1_ASAP7_75t_L g139 ( .A(n_65), .Y(n_139) );
NAND2xp5_ASAP7_75t_L g456 ( .A(n_66), .B(n_457), .Y(n_456) );
INVx1_ASAP7_75t_SL g521 ( .A(n_67), .Y(n_521) );
CKINVDCx20_ASAP7_75t_R g118 ( .A(n_68), .Y(n_118) );
NAND2xp5_ASAP7_75t_SL g218 ( .A(n_69), .B(n_178), .Y(n_218) );
NAND2xp5_ASAP7_75t_L g512 ( .A(n_70), .B(n_208), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g155 ( .A(n_71), .B(n_156), .Y(n_155) );
INVx1_ASAP7_75t_L g554 ( .A(n_72), .Y(n_554) );
CKINVDCx16_ASAP7_75t_R g265 ( .A(n_73), .Y(n_265) );
NAND2xp5_ASAP7_75t_L g229 ( .A(n_74), .B(n_175), .Y(n_229) );
A2O1A1Ixp33_ASAP7_75t_L g241 ( .A1(n_75), .A2(n_151), .B(n_181), .C(n_242), .Y(n_241) );
CKINVDCx16_ASAP7_75t_R g200 ( .A(n_76), .Y(n_200) );
INVx1_ASAP7_75t_L g112 ( .A(n_77), .Y(n_112) );
AOI21xp5_ASAP7_75t_L g487 ( .A1(n_78), .A2(n_168), .B(n_488), .Y(n_487) );
CKINVDCx20_ASAP7_75t_R g451 ( .A(n_79), .Y(n_451) );
AOI21xp5_ASAP7_75t_L g497 ( .A1(n_80), .A2(n_168), .B(n_498), .Y(n_497) );
AOI21xp5_ASAP7_75t_L g529 ( .A1(n_81), .A2(n_226), .B(n_530), .Y(n_529) );
INVx1_ASAP7_75t_L g499 ( .A(n_82), .Y(n_499) );
CKINVDCx16_ASAP7_75t_R g540 ( .A(n_83), .Y(n_540) );
NAND2xp5_ASAP7_75t_SL g230 ( .A(n_84), .B(n_174), .Y(n_230) );
CKINVDCx20_ASAP7_75t_R g220 ( .A(n_85), .Y(n_220) );
AOI21xp5_ASAP7_75t_L g506 ( .A1(n_86), .A2(n_168), .B(n_507), .Y(n_506) );
INVx1_ASAP7_75t_L g502 ( .A(n_87), .Y(n_502) );
INVx2_ASAP7_75t_L g137 ( .A(n_88), .Y(n_137) );
INVx1_ASAP7_75t_L g478 ( .A(n_89), .Y(n_478) );
CKINVDCx20_ASAP7_75t_R g249 ( .A(n_90), .Y(n_249) );
NAND2xp5_ASAP7_75t_SL g157 ( .A(n_91), .B(n_158), .Y(n_157) );
OR2x2_ASAP7_75t_L g444 ( .A(n_92), .B(n_445), .Y(n_444) );
OR2x2_ASAP7_75t_L g464 ( .A(n_92), .B(n_446), .Y(n_464) );
INVx2_ASAP7_75t_L g734 ( .A(n_92), .Y(n_734) );
A2O1A1Ixp33_ASAP7_75t_L g552 ( .A1(n_93), .A2(n_151), .B(n_181), .C(n_553), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g214 ( .A(n_94), .B(n_168), .Y(n_214) );
AOI22xp5_ASAP7_75t_L g736 ( .A1(n_95), .A2(n_737), .B1(n_738), .B2(n_739), .Y(n_736) );
CKINVDCx20_ASAP7_75t_R g737 ( .A(n_95), .Y(n_737) );
INVx1_ASAP7_75t_L g217 ( .A(n_96), .Y(n_217) );
INVxp67_ASAP7_75t_L g205 ( .A(n_97), .Y(n_205) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_98), .B(n_135), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g111 ( .A(n_99), .B(n_112), .Y(n_111) );
INVx1_ASAP7_75t_L g142 ( .A(n_100), .Y(n_142) );
INVx1_ASAP7_75t_L g243 ( .A(n_101), .Y(n_243) );
INVx2_ASAP7_75t_L g511 ( .A(n_102), .Y(n_511) );
AND2x2_ASAP7_75t_L g184 ( .A(n_103), .B(n_183), .Y(n_184) );
INVx1_ASAP7_75t_SL g105 ( .A(n_106), .Y(n_105) );
BUFx4f_ASAP7_75t_SL g753 ( .A(n_106), .Y(n_753) );
OR2x2_ASAP7_75t_L g106 ( .A(n_107), .B(n_109), .Y(n_106) );
INVx1_ASAP7_75t_SL g110 ( .A(n_111), .Y(n_110) );
OA21x2_ASAP7_75t_L g113 ( .A1(n_114), .A2(n_119), .B(n_459), .Y(n_113) );
BUFx2_ASAP7_75t_SL g114 ( .A(n_115), .Y(n_114) );
CKINVDCx20_ASAP7_75t_R g115 ( .A(n_116), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
INVx1_ASAP7_75t_SL g752 ( .A(n_117), .Y(n_752) );
INVx2_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
OAI321xp33_ASAP7_75t_L g119 ( .A1(n_120), .A2(n_442), .A3(n_449), .B1(n_452), .B2(n_453), .C(n_456), .Y(n_119) );
NAND2xp5_ASAP7_75t_SL g453 ( .A(n_120), .B(n_454), .Y(n_453) );
AOI22xp5_ASAP7_75t_L g120 ( .A1(n_121), .A2(n_122), .B1(n_125), .B2(n_126), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
OAI22x1_ASAP7_75t_SL g461 ( .A1(n_125), .A2(n_462), .B1(n_465), .B2(n_731), .Y(n_461) );
INVx2_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
OAI22xp5_ASAP7_75t_SL g745 ( .A1(n_126), .A2(n_466), .B1(n_746), .B2(n_747), .Y(n_745) );
OR3x1_ASAP7_75t_L g126 ( .A(n_127), .B(n_340), .C(n_405), .Y(n_126) );
NAND4xp25_ASAP7_75t_SL g127 ( .A(n_128), .B(n_281), .C(n_307), .D(n_330), .Y(n_127) );
AOI221xp5_ASAP7_75t_L g128 ( .A1(n_129), .A2(n_209), .B1(n_250), .B2(n_257), .C(n_273), .Y(n_128) );
CKINVDCx14_ASAP7_75t_R g129 ( .A(n_130), .Y(n_129) );
OAI22xp5_ASAP7_75t_L g428 ( .A1(n_130), .A2(n_274), .B1(n_298), .B2(n_429), .Y(n_428) );
OR2x2_ASAP7_75t_L g130 ( .A(n_131), .B(n_185), .Y(n_130) );
INVx1_ASAP7_75t_SL g334 ( .A(n_131), .Y(n_334) );
OR2x2_ASAP7_75t_L g131 ( .A(n_132), .B(n_165), .Y(n_131) );
OR2x2_ASAP7_75t_L g255 ( .A(n_132), .B(n_256), .Y(n_255) );
AND2x2_ASAP7_75t_L g276 ( .A(n_132), .B(n_186), .Y(n_276) );
NAND2xp5_ASAP7_75t_L g289 ( .A(n_132), .B(n_196), .Y(n_289) );
AND2x2_ASAP7_75t_L g306 ( .A(n_132), .B(n_165), .Y(n_306) );
NAND2xp5_ASAP7_75t_L g328 ( .A(n_132), .B(n_253), .Y(n_328) );
NAND2xp5_ASAP7_75t_L g417 ( .A(n_132), .B(n_305), .Y(n_417) );
NOR2xp33_ASAP7_75t_L g427 ( .A(n_132), .B(n_185), .Y(n_427) );
AOI211xp5_ASAP7_75t_SL g438 ( .A1(n_132), .A2(n_344), .B(n_439), .C(n_440), .Y(n_438) );
INVx5_ASAP7_75t_SL g132 ( .A(n_133), .Y(n_132) );
NAND2xp5_ASAP7_75t_SL g310 ( .A(n_133), .B(n_186), .Y(n_310) );
AND2x2_ASAP7_75t_L g313 ( .A(n_133), .B(n_187), .Y(n_313) );
OR2x2_ASAP7_75t_L g358 ( .A(n_133), .B(n_186), .Y(n_358) );
NAND2xp5_ASAP7_75t_L g367 ( .A(n_133), .B(n_196), .Y(n_367) );
AO21x2_ASAP7_75t_L g133 ( .A1(n_134), .A2(n_141), .B(n_162), .Y(n_133) );
INVx3_ASAP7_75t_L g208 ( .A(n_134), .Y(n_208) );
NOR2xp33_ASAP7_75t_L g219 ( .A(n_134), .B(n_220), .Y(n_219) );
AO21x2_ASAP7_75t_L g239 ( .A1(n_134), .A2(n_240), .B(n_248), .Y(n_239) );
NOR2xp33_ASAP7_75t_L g248 ( .A(n_134), .B(n_249), .Y(n_248) );
NOR2xp33_ASAP7_75t_L g481 ( .A(n_134), .B(n_482), .Y(n_481) );
NOR2xp33_ASAP7_75t_L g545 ( .A(n_134), .B(n_546), .Y(n_545) );
AO21x2_ASAP7_75t_L g549 ( .A1(n_134), .A2(n_550), .B(n_556), .Y(n_549) );
INVx4_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
AOI21xp5_ASAP7_75t_L g188 ( .A1(n_135), .A2(n_189), .B(n_190), .Y(n_188) );
HB1xp67_ASAP7_75t_L g197 ( .A(n_135), .Y(n_197) );
BUFx6f_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
INVx1_ASAP7_75t_L g164 ( .A(n_136), .Y(n_164) );
AND2x2_ASAP7_75t_L g136 ( .A(n_137), .B(n_138), .Y(n_136) );
AND2x2_ASAP7_75t_SL g183 ( .A(n_137), .B(n_138), .Y(n_183) );
NAND2xp5_ASAP7_75t_L g138 ( .A(n_139), .B(n_140), .Y(n_138) );
OAI21xp5_ASAP7_75t_L g141 ( .A1(n_142), .A2(n_143), .B(n_150), .Y(n_141) );
OAI21xp5_ASAP7_75t_L g474 ( .A1(n_143), .A2(n_475), .B(n_476), .Y(n_474) );
O2A1O1Ixp33_ASAP7_75t_L g539 ( .A1(n_143), .A2(n_183), .B(n_540), .C(n_541), .Y(n_539) );
OAI21xp5_ASAP7_75t_L g550 ( .A1(n_143), .A2(n_551), .B(n_552), .Y(n_550) );
NAND2x1p5_ASAP7_75t_L g143 ( .A(n_144), .B(n_148), .Y(n_143) );
AND2x4_ASAP7_75t_L g168 ( .A(n_144), .B(n_148), .Y(n_168) );
AND2x2_ASAP7_75t_L g144 ( .A(n_145), .B(n_147), .Y(n_144) );
INVx1_ASAP7_75t_L g206 ( .A(n_145), .Y(n_206) );
INVx1_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
INVx2_ASAP7_75t_L g152 ( .A(n_146), .Y(n_152) );
INVx1_ASAP7_75t_L g161 ( .A(n_146), .Y(n_161) );
INVx1_ASAP7_75t_L g153 ( .A(n_147), .Y(n_153) );
INVx3_ASAP7_75t_L g156 ( .A(n_147), .Y(n_156) );
BUFx6f_ASAP7_75t_L g158 ( .A(n_147), .Y(n_158) );
BUFx6f_ASAP7_75t_L g176 ( .A(n_147), .Y(n_176) );
INVx1_ASAP7_75t_L g193 ( .A(n_147), .Y(n_193) );
INVx4_ASAP7_75t_SL g182 ( .A(n_148), .Y(n_182) );
BUFx3_ASAP7_75t_L g195 ( .A(n_148), .Y(n_195) );
INVx5_ASAP7_75t_L g171 ( .A(n_151), .Y(n_171) );
AND2x6_ASAP7_75t_L g151 ( .A(n_152), .B(n_153), .Y(n_151) );
BUFx3_ASAP7_75t_L g180 ( .A(n_152), .Y(n_180) );
BUFx6f_ASAP7_75t_L g246 ( .A(n_152), .Y(n_246) );
AOI21xp5_ASAP7_75t_L g154 ( .A1(n_155), .A2(n_157), .B(n_159), .Y(n_154) );
INVx5_ASAP7_75t_L g178 ( .A(n_156), .Y(n_178) );
NOR2xp33_ASAP7_75t_L g492 ( .A(n_156), .B(n_493), .Y(n_492) );
INVx4_ASAP7_75t_L g270 ( .A(n_158), .Y(n_270) );
INVx2_ASAP7_75t_L g491 ( .A(n_158), .Y(n_491) );
AOI21xp5_ASAP7_75t_L g191 ( .A1(n_159), .A2(n_192), .B(n_194), .Y(n_191) );
INVx2_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
INVx3_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
NOR2xp33_ASAP7_75t_L g162 ( .A(n_163), .B(n_164), .Y(n_162) );
INVx2_ASAP7_75t_L g528 ( .A(n_164), .Y(n_528) );
INVx5_ASAP7_75t_SL g256 ( .A(n_165), .Y(n_256) );
AND2x2_ASAP7_75t_L g275 ( .A(n_165), .B(n_276), .Y(n_275) );
NOR2xp33_ASAP7_75t_L g357 ( .A(n_165), .B(n_358), .Y(n_357) );
AND2x2_ASAP7_75t_L g361 ( .A(n_165), .B(n_362), .Y(n_361) );
AND2x2_ASAP7_75t_L g393 ( .A(n_165), .B(n_196), .Y(n_393) );
OR2x2_ASAP7_75t_L g399 ( .A(n_165), .B(n_289), .Y(n_399) );
NAND2xp5_ASAP7_75t_L g408 ( .A(n_165), .B(n_349), .Y(n_408) );
OR2x6_ASAP7_75t_L g165 ( .A(n_166), .B(n_184), .Y(n_165) );
AOI21xp5_ASAP7_75t_L g166 ( .A1(n_167), .A2(n_169), .B(n_183), .Y(n_166) );
BUFx2_ASAP7_75t_L g226 ( .A(n_168), .Y(n_226) );
INVx2_ASAP7_75t_L g170 ( .A(n_171), .Y(n_170) );
O2A1O1Ixp33_ASAP7_75t_L g199 ( .A1(n_171), .A2(n_182), .B(n_200), .C(n_201), .Y(n_199) );
O2A1O1Ixp33_ASAP7_75t_SL g264 ( .A1(n_171), .A2(n_182), .B(n_265), .C(n_266), .Y(n_264) );
O2A1O1Ixp33_ASAP7_75t_SL g488 ( .A1(n_171), .A2(n_182), .B(n_489), .C(n_490), .Y(n_488) );
O2A1O1Ixp33_ASAP7_75t_SL g498 ( .A1(n_171), .A2(n_182), .B(n_499), .C(n_500), .Y(n_498) );
O2A1O1Ixp33_ASAP7_75t_SL g507 ( .A1(n_171), .A2(n_182), .B(n_508), .C(n_509), .Y(n_507) );
O2A1O1Ixp33_ASAP7_75t_L g517 ( .A1(n_171), .A2(n_182), .B(n_518), .C(n_519), .Y(n_517) );
O2A1O1Ixp33_ASAP7_75t_SL g530 ( .A1(n_171), .A2(n_182), .B(n_531), .C(n_532), .Y(n_530) );
O2A1O1Ixp33_ASAP7_75t_L g172 ( .A1(n_173), .A2(n_174), .B(n_177), .C(n_179), .Y(n_172) );
O2A1O1Ixp33_ASAP7_75t_L g216 ( .A1(n_174), .A2(n_179), .B(n_217), .C(n_218), .Y(n_216) );
O2A1O1Ixp5_ASAP7_75t_L g477 ( .A1(n_174), .A2(n_478), .B(n_479), .C(n_480), .Y(n_477) );
O2A1O1Ixp33_ASAP7_75t_L g553 ( .A1(n_174), .A2(n_480), .B(n_554), .C(n_555), .Y(n_553) );
INVx2_ASAP7_75t_L g174 ( .A(n_175), .Y(n_174) );
INVx2_ASAP7_75t_L g175 ( .A(n_176), .Y(n_175) );
INVx4_ASAP7_75t_L g203 ( .A(n_176), .Y(n_203) );
NOR2xp33_ASAP7_75t_L g204 ( .A(n_178), .B(n_205), .Y(n_204) );
INVx2_ASAP7_75t_L g267 ( .A(n_178), .Y(n_267) );
OAI22xp33_ASAP7_75t_L g533 ( .A1(n_178), .A2(n_203), .B1(n_534), .B2(n_535), .Y(n_533) );
O2A1O1Ixp33_ASAP7_75t_L g542 ( .A1(n_178), .A2(n_231), .B(n_543), .C(n_544), .Y(n_542) );
HB1xp67_ASAP7_75t_L g179 ( .A(n_180), .Y(n_179) );
INVx2_ASAP7_75t_L g271 ( .A(n_180), .Y(n_271) );
INVx1_ASAP7_75t_L g503 ( .A(n_180), .Y(n_503) );
INVx1_ASAP7_75t_L g181 ( .A(n_182), .Y(n_181) );
AOI21xp5_ASAP7_75t_L g213 ( .A1(n_183), .A2(n_214), .B(n_215), .Y(n_213) );
INVx2_ASAP7_75t_L g233 ( .A(n_183), .Y(n_233) );
INVx1_ASAP7_75t_L g236 ( .A(n_183), .Y(n_236) );
OA21x2_ASAP7_75t_L g486 ( .A1(n_183), .A2(n_487), .B(n_494), .Y(n_486) );
NAND2xp5_ASAP7_75t_L g185 ( .A(n_186), .B(n_196), .Y(n_185) );
AND2x2_ASAP7_75t_L g290 ( .A(n_186), .B(n_256), .Y(n_290) );
INVx1_ASAP7_75t_SL g303 ( .A(n_186), .Y(n_303) );
OR2x2_ASAP7_75t_L g338 ( .A(n_186), .B(n_339), .Y(n_338) );
OR2x2_ASAP7_75t_L g344 ( .A(n_186), .B(n_196), .Y(n_344) );
AND2x2_ASAP7_75t_L g402 ( .A(n_186), .B(n_253), .Y(n_402) );
INVx2_ASAP7_75t_L g186 ( .A(n_187), .Y(n_186) );
NAND2xp5_ASAP7_75t_L g329 ( .A(n_187), .B(n_256), .Y(n_329) );
INVx3_ASAP7_75t_L g253 ( .A(n_196), .Y(n_253) );
OR2x2_ASAP7_75t_L g295 ( .A(n_196), .B(n_256), .Y(n_295) );
AND2x2_ASAP7_75t_L g305 ( .A(n_196), .B(n_303), .Y(n_305) );
HB1xp67_ASAP7_75t_L g353 ( .A(n_196), .Y(n_353) );
AND2x2_ASAP7_75t_L g362 ( .A(n_196), .B(n_276), .Y(n_362) );
OA21x2_ASAP7_75t_L g196 ( .A1(n_197), .A2(n_198), .B(n_207), .Y(n_196) );
OA21x2_ASAP7_75t_L g496 ( .A1(n_197), .A2(n_497), .B(n_504), .Y(n_496) );
OA21x2_ASAP7_75t_L g505 ( .A1(n_197), .A2(n_506), .B(n_512), .Y(n_505) );
OA21x2_ASAP7_75t_L g515 ( .A1(n_197), .A2(n_516), .B(n_523), .Y(n_515) );
O2A1O1Ixp33_ASAP7_75t_L g242 ( .A1(n_202), .A2(n_243), .B(n_244), .C(n_245), .Y(n_242) );
INVx1_ASAP7_75t_L g202 ( .A(n_203), .Y(n_202) );
NOR2xp33_ASAP7_75t_L g501 ( .A(n_203), .B(n_502), .Y(n_501) );
NOR2xp33_ASAP7_75t_L g510 ( .A(n_203), .B(n_511), .Y(n_510) );
INVx2_ASAP7_75t_L g231 ( .A(n_206), .Y(n_231) );
NAND2xp5_ASAP7_75t_SL g532 ( .A(n_206), .B(n_533), .Y(n_532) );
OA21x2_ASAP7_75t_L g262 ( .A1(n_208), .A2(n_263), .B(n_272), .Y(n_262) );
AOI221xp5_ASAP7_75t_L g378 ( .A1(n_209), .A2(n_379), .B1(n_381), .B2(n_383), .C(n_386), .Y(n_378) );
INVx2_ASAP7_75t_L g209 ( .A(n_210), .Y(n_209) );
OR2x2_ASAP7_75t_L g210 ( .A(n_211), .B(n_221), .Y(n_210) );
AND2x2_ASAP7_75t_L g352 ( .A(n_211), .B(n_333), .Y(n_352) );
NAND2xp5_ASAP7_75t_L g415 ( .A(n_211), .B(n_411), .Y(n_415) );
OR2x2_ASAP7_75t_L g436 ( .A(n_211), .B(n_437), .Y(n_436) );
NAND2xp5_ASAP7_75t_L g440 ( .A(n_211), .B(n_441), .Y(n_440) );
BUFx2_ASAP7_75t_L g211 ( .A(n_212), .Y(n_211) );
INVx5_ASAP7_75t_L g283 ( .A(n_212), .Y(n_283) );
AND2x2_ASAP7_75t_L g360 ( .A(n_212), .B(n_223), .Y(n_360) );
AND2x2_ASAP7_75t_L g421 ( .A(n_212), .B(n_300), .Y(n_421) );
AND2x2_ASAP7_75t_L g434 ( .A(n_212), .B(n_253), .Y(n_434) );
OR2x6_ASAP7_75t_L g212 ( .A(n_213), .B(n_219), .Y(n_212) );
NAND2xp5_ASAP7_75t_L g221 ( .A(n_222), .B(n_237), .Y(n_221) );
AND2x4_ASAP7_75t_L g260 ( .A(n_222), .B(n_261), .Y(n_260) );
AND2x2_ASAP7_75t_L g279 ( .A(n_222), .B(n_280), .Y(n_279) );
INVx2_ASAP7_75t_L g286 ( .A(n_222), .Y(n_286) );
AND2x2_ASAP7_75t_L g355 ( .A(n_222), .B(n_333), .Y(n_355) );
AND2x2_ASAP7_75t_L g365 ( .A(n_222), .B(n_283), .Y(n_365) );
HB1xp67_ASAP7_75t_L g373 ( .A(n_222), .Y(n_373) );
AND2x2_ASAP7_75t_L g385 ( .A(n_222), .B(n_262), .Y(n_385) );
NOR2xp33_ASAP7_75t_L g389 ( .A(n_222), .B(n_317), .Y(n_389) );
AND2x2_ASAP7_75t_L g426 ( .A(n_222), .B(n_421), .Y(n_426) );
NAND2xp5_ASAP7_75t_L g437 ( .A(n_222), .B(n_300), .Y(n_437) );
OR2x2_ASAP7_75t_L g439 ( .A(n_222), .B(n_375), .Y(n_439) );
INVx5_ASAP7_75t_L g222 ( .A(n_223), .Y(n_222) );
AND2x2_ASAP7_75t_L g325 ( .A(n_223), .B(n_326), .Y(n_325) );
AND2x2_ASAP7_75t_L g335 ( .A(n_223), .B(n_280), .Y(n_335) );
AND2x2_ASAP7_75t_L g347 ( .A(n_223), .B(n_262), .Y(n_347) );
HB1xp67_ASAP7_75t_L g377 ( .A(n_223), .Y(n_377) );
AND2x4_ASAP7_75t_L g411 ( .A(n_223), .B(n_261), .Y(n_411) );
OR2x6_ASAP7_75t_L g223 ( .A(n_224), .B(n_234), .Y(n_223) );
AOI21xp5_ASAP7_75t_SL g224 ( .A1(n_225), .A2(n_227), .B(n_232), .Y(n_224) );
AOI21xp5_ASAP7_75t_L g228 ( .A1(n_229), .A2(n_230), .B(n_231), .Y(n_228) );
INVx1_ASAP7_75t_L g232 ( .A(n_233), .Y(n_232) );
NOR2xp33_ASAP7_75t_L g556 ( .A(n_233), .B(n_451), .Y(n_556) );
NOR2xp33_ASAP7_75t_L g234 ( .A(n_235), .B(n_236), .Y(n_234) );
AO21x2_ASAP7_75t_L g473 ( .A1(n_236), .A2(n_474), .B(n_481), .Y(n_473) );
BUFx2_ASAP7_75t_L g259 ( .A(n_237), .Y(n_259) );
HB1xp67_ASAP7_75t_L g237 ( .A(n_238), .Y(n_237) );
INVx2_ASAP7_75t_L g300 ( .A(n_238), .Y(n_300) );
AND2x2_ASAP7_75t_L g333 ( .A(n_238), .B(n_262), .Y(n_333) );
INVx2_ASAP7_75t_L g238 ( .A(n_239), .Y(n_238) );
AND2x2_ASAP7_75t_L g280 ( .A(n_239), .B(n_262), .Y(n_280) );
BUFx2_ASAP7_75t_L g326 ( .A(n_239), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g240 ( .A(n_241), .B(n_247), .Y(n_240) );
HB1xp67_ASAP7_75t_L g245 ( .A(n_246), .Y(n_245) );
INVx3_ASAP7_75t_L g522 ( .A(n_246), .Y(n_522) );
INVx1_ASAP7_75t_L g250 ( .A(n_251), .Y(n_250) );
NAND2xp5_ASAP7_75t_L g251 ( .A(n_252), .B(n_254), .Y(n_251) );
NAND2xp5_ASAP7_75t_L g413 ( .A(n_252), .B(n_334), .Y(n_413) );
INVx1_ASAP7_75t_L g252 ( .A(n_253), .Y(n_252) );
NAND2xp5_ASAP7_75t_L g277 ( .A(n_253), .B(n_276), .Y(n_277) );
NAND2xp5_ASAP7_75t_L g315 ( .A(n_253), .B(n_256), .Y(n_315) );
AND2x2_ASAP7_75t_L g370 ( .A(n_253), .B(n_306), .Y(n_370) );
AOI221xp5_ASAP7_75t_SL g307 ( .A1(n_254), .A2(n_308), .B1(n_316), .B2(n_318), .C(n_322), .Y(n_307) );
INVx2_ASAP7_75t_L g254 ( .A(n_255), .Y(n_254) );
OR2x2_ASAP7_75t_L g302 ( .A(n_255), .B(n_303), .Y(n_302) );
OR2x2_ASAP7_75t_L g343 ( .A(n_255), .B(n_344), .Y(n_343) );
OAI321xp33_ASAP7_75t_L g350 ( .A1(n_255), .A2(n_309), .A3(n_351), .B1(n_353), .B2(n_354), .C(n_356), .Y(n_350) );
NAND2xp5_ASAP7_75t_L g401 ( .A(n_256), .B(n_402), .Y(n_401) );
INVx1_ASAP7_75t_L g257 ( .A(n_258), .Y(n_257) );
NAND2xp5_ASAP7_75t_L g258 ( .A(n_259), .B(n_260), .Y(n_258) );
NAND2xp5_ASAP7_75t_L g429 ( .A(n_259), .B(n_411), .Y(n_429) );
AND2x2_ASAP7_75t_L g316 ( .A(n_260), .B(n_317), .Y(n_316) );
NAND2xp5_ASAP7_75t_L g319 ( .A(n_260), .B(n_320), .Y(n_319) );
HB1xp67_ASAP7_75t_L g292 ( .A(n_261), .Y(n_292) );
AND2x2_ASAP7_75t_L g299 ( .A(n_261), .B(n_300), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g404 ( .A(n_261), .B(n_374), .Y(n_404) );
INVx1_ASAP7_75t_L g441 ( .A(n_261), .Y(n_441) );
INVx2_ASAP7_75t_L g261 ( .A(n_262), .Y(n_261) );
NOR2xp33_ASAP7_75t_L g268 ( .A(n_269), .B(n_270), .Y(n_268) );
NOR2xp33_ASAP7_75t_L g520 ( .A(n_270), .B(n_521), .Y(n_520) );
INVx2_ASAP7_75t_L g480 ( .A(n_271), .Y(n_480) );
AOI21xp5_ASAP7_75t_L g273 ( .A1(n_274), .A2(n_277), .B(n_278), .Y(n_273) );
INVx1_ASAP7_75t_SL g274 ( .A(n_275), .Y(n_274) );
A2O1A1Ixp33_ASAP7_75t_L g433 ( .A1(n_275), .A2(n_385), .B(n_434), .C(n_435), .Y(n_433) );
NAND2xp5_ASAP7_75t_L g293 ( .A(n_276), .B(n_294), .Y(n_293) );
NAND2xp5_ASAP7_75t_L g380 ( .A(n_276), .B(n_314), .Y(n_380) );
INVx1_ASAP7_75t_SL g278 ( .A(n_279), .Y(n_278) );
INVx1_ASAP7_75t_L g323 ( .A(n_280), .Y(n_323) );
NAND2xp5_ASAP7_75t_L g337 ( .A(n_280), .B(n_283), .Y(n_337) );
NOR2xp33_ASAP7_75t_L g346 ( .A(n_280), .B(n_347), .Y(n_346) );
NAND2xp5_ASAP7_75t_L g364 ( .A(n_280), .B(n_365), .Y(n_364) );
AOI22xp33_ASAP7_75t_L g281 ( .A1(n_282), .A2(n_284), .B1(n_296), .B2(n_301), .Y(n_281) );
HB1xp67_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
OR2x2_ASAP7_75t_L g297 ( .A(n_283), .B(n_298), .Y(n_297) );
AND2x2_ASAP7_75t_L g320 ( .A(n_283), .B(n_321), .Y(n_320) );
AND2x2_ASAP7_75t_L g332 ( .A(n_283), .B(n_333), .Y(n_332) );
NAND2xp5_ASAP7_75t_L g368 ( .A(n_283), .B(n_326), .Y(n_368) );
OR2x2_ASAP7_75t_L g375 ( .A(n_283), .B(n_300), .Y(n_375) );
NAND2xp5_ASAP7_75t_L g384 ( .A(n_283), .B(n_385), .Y(n_384) );
AND2x2_ASAP7_75t_L g425 ( .A(n_283), .B(n_411), .Y(n_425) );
OAI22xp33_ASAP7_75t_L g284 ( .A1(n_285), .A2(n_287), .B1(n_291), .B2(n_293), .Y(n_284) );
INVx1_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
AND2x2_ASAP7_75t_L g331 ( .A(n_286), .B(n_332), .Y(n_331) );
NAND2xp5_ASAP7_75t_L g287 ( .A(n_288), .B(n_290), .Y(n_287) );
INVx1_ASAP7_75t_SL g288 ( .A(n_289), .Y(n_288) );
OAI22xp33_ASAP7_75t_L g371 ( .A1(n_289), .A2(n_304), .B1(n_372), .B2(n_376), .Y(n_371) );
INVx1_ASAP7_75t_L g419 ( .A(n_290), .Y(n_419) );
INVx1_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
AOI221xp5_ASAP7_75t_L g330 ( .A1(n_294), .A2(n_331), .B1(n_334), .B2(n_335), .C(n_336), .Y(n_330) );
INVx1_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
OR2x2_ASAP7_75t_L g309 ( .A(n_295), .B(n_310), .Y(n_309) );
INVx1_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
INVx1_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
NAND2xp5_ASAP7_75t_L g397 ( .A(n_299), .B(n_365), .Y(n_397) );
HB1xp67_ASAP7_75t_L g317 ( .A(n_300), .Y(n_317) );
INVx1_ASAP7_75t_L g321 ( .A(n_300), .Y(n_321) );
NAND2xp33_ASAP7_75t_L g301 ( .A(n_302), .B(n_304), .Y(n_301) );
NAND2xp5_ASAP7_75t_L g304 ( .A(n_305), .B(n_306), .Y(n_304) );
INVx1_ASAP7_75t_L g339 ( .A(n_306), .Y(n_339) );
AND2x2_ASAP7_75t_L g348 ( .A(n_306), .B(n_349), .Y(n_348) );
NAND2xp33_ASAP7_75t_L g308 ( .A(n_309), .B(n_311), .Y(n_308) );
INVx2_ASAP7_75t_SL g311 ( .A(n_312), .Y(n_311) );
AND2x4_ASAP7_75t_L g312 ( .A(n_313), .B(n_314), .Y(n_312) );
AND2x2_ASAP7_75t_L g392 ( .A(n_313), .B(n_393), .Y(n_392) );
INVx2_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
AOI221xp5_ASAP7_75t_L g341 ( .A1(n_316), .A2(n_342), .B1(n_345), .B2(n_348), .C(n_350), .Y(n_341) );
INVx1_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
NAND2xp5_ASAP7_75t_L g376 ( .A(n_320), .B(n_377), .Y(n_376) );
AOI21xp33_ASAP7_75t_SL g322 ( .A1(n_323), .A2(n_324), .B(n_327), .Y(n_322) );
INVx2_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
CKINVDCx16_ASAP7_75t_R g424 ( .A(n_327), .Y(n_424) );
OR2x2_ASAP7_75t_L g327 ( .A(n_328), .B(n_329), .Y(n_327) );
OR2x2_ASAP7_75t_L g366 ( .A(n_329), .B(n_367), .Y(n_366) );
INVx1_ASAP7_75t_SL g387 ( .A(n_332), .Y(n_387) );
NAND2xp5_ASAP7_75t_L g432 ( .A(n_332), .B(n_392), .Y(n_432) );
NAND2xp5_ASAP7_75t_L g356 ( .A(n_335), .B(n_357), .Y(n_356) );
NOR2xp33_ASAP7_75t_L g336 ( .A(n_337), .B(n_338), .Y(n_336) );
NAND4xp25_ASAP7_75t_L g340 ( .A(n_341), .B(n_359), .C(n_378), .D(n_391), .Y(n_340) );
INVx1_ASAP7_75t_SL g342 ( .A(n_343), .Y(n_342) );
INVx1_ASAP7_75t_SL g349 ( .A(n_344), .Y(n_349) );
INVxp67_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
INVx1_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
OR2x2_ASAP7_75t_L g382 ( .A(n_353), .B(n_358), .Y(n_382) );
INVxp67_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
AOI211xp5_ASAP7_75t_L g359 ( .A1(n_360), .A2(n_361), .B(n_363), .C(n_371), .Y(n_359) );
AOI211xp5_ASAP7_75t_L g430 ( .A1(n_361), .A2(n_403), .B(n_431), .C(n_438), .Y(n_430) );
INVx1_ASAP7_75t_SL g390 ( .A(n_362), .Y(n_390) );
OAI22xp5_ASAP7_75t_L g363 ( .A1(n_364), .A2(n_366), .B1(n_368), .B2(n_369), .Y(n_363) );
INVx1_ASAP7_75t_L g394 ( .A(n_368), .Y(n_394) );
INVx1_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_373), .B(n_374), .Y(n_372) );
NAND2xp5_ASAP7_75t_L g410 ( .A(n_374), .B(n_411), .Y(n_410) );
NAND2xp5_ASAP7_75t_L g418 ( .A(n_374), .B(n_385), .Y(n_418) );
INVx2_ASAP7_75t_SL g374 ( .A(n_375), .Y(n_374) );
INVx1_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
INVx1_ASAP7_75t_SL g381 ( .A(n_382), .Y(n_381) );
INVx1_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
INVx1_ASAP7_75t_L g395 ( .A(n_385), .Y(n_395) );
AOI21xp33_ASAP7_75t_L g386 ( .A1(n_387), .A2(n_388), .B(n_390), .Y(n_386) );
INVxp33_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
AOI322xp5_ASAP7_75t_L g391 ( .A1(n_392), .A2(n_394), .A3(n_395), .B1(n_396), .B2(n_398), .C1(n_400), .C2(n_403), .Y(n_391) );
INVxp67_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
INVx1_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
INVx1_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
INVx1_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
NAND3xp33_ASAP7_75t_SL g405 ( .A(n_406), .B(n_423), .C(n_430), .Y(n_405) );
AOI221xp5_ASAP7_75t_L g406 ( .A1(n_407), .A2(n_409), .B1(n_412), .B2(n_414), .C(n_416), .Y(n_406) );
INVx1_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
INVx1_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
INVx1_ASAP7_75t_SL g422 ( .A(n_411), .Y(n_422) );
INVx1_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
INVxp67_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
OAI22xp33_ASAP7_75t_L g416 ( .A1(n_417), .A2(n_418), .B1(n_419), .B2(n_420), .Y(n_416) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_421), .B(n_422), .Y(n_420) );
AOI221xp5_ASAP7_75t_L g423 ( .A1(n_424), .A2(n_425), .B1(n_426), .B2(n_427), .C(n_428), .Y(n_423) );
NAND2xp33_ASAP7_75t_L g431 ( .A(n_432), .B(n_433), .Y(n_431) );
INVxp67_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
INVx1_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
HB1xp67_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
INVx1_ASAP7_75t_SL g455 ( .A(n_444), .Y(n_455) );
HB1xp67_ASAP7_75t_L g458 ( .A(n_444), .Y(n_458) );
NOR2x2_ASAP7_75t_L g750 ( .A(n_445), .B(n_734), .Y(n_750) );
INVx2_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
OR2x2_ASAP7_75t_L g733 ( .A(n_446), .B(n_734), .Y(n_733) );
AND2x2_ASAP7_75t_L g446 ( .A(n_447), .B(n_448), .Y(n_446) );
INVx1_ASAP7_75t_L g452 ( .A(n_449), .Y(n_452) );
INVx1_ASAP7_75t_SL g454 ( .A(n_455), .Y(n_454) );
NAND3xp33_ASAP7_75t_L g459 ( .A(n_456), .B(n_460), .C(n_751), .Y(n_459) );
INVx1_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
INVx2_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
INVx2_ASAP7_75t_L g746 ( .A(n_463), .Y(n_746) );
INVx1_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
INVx2_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
OR2x2_ASAP7_75t_SL g466 ( .A(n_467), .B(n_686), .Y(n_466) );
NAND5xp2_ASAP7_75t_L g467 ( .A(n_468), .B(n_598), .C(n_636), .D(n_657), .E(n_674), .Y(n_467) );
NOR3xp33_ASAP7_75t_L g468 ( .A(n_469), .B(n_570), .C(n_591), .Y(n_468) );
OAI221xp5_ASAP7_75t_SL g469 ( .A1(n_470), .A2(n_513), .B1(n_537), .B2(n_557), .C(n_561), .Y(n_469) );
NAND2xp5_ASAP7_75t_L g470 ( .A(n_471), .B(n_483), .Y(n_470) );
INVx1_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
NAND2xp5_ASAP7_75t_L g578 ( .A(n_472), .B(n_559), .Y(n_578) );
OR2x2_ASAP7_75t_L g605 ( .A(n_472), .B(n_496), .Y(n_605) );
AND2x2_ASAP7_75t_L g619 ( .A(n_472), .B(n_496), .Y(n_619) );
NOR2xp33_ASAP7_75t_L g633 ( .A(n_472), .B(n_486), .Y(n_633) );
AND2x2_ASAP7_75t_L g671 ( .A(n_472), .B(n_635), .Y(n_671) );
AND2x2_ASAP7_75t_L g700 ( .A(n_472), .B(n_610), .Y(n_700) );
NAND2xp5_ASAP7_75t_L g717 ( .A(n_472), .B(n_582), .Y(n_717) );
INVx4_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
AND2x2_ASAP7_75t_L g597 ( .A(n_473), .B(n_495), .Y(n_597) );
BUFx3_ASAP7_75t_L g622 ( .A(n_473), .Y(n_622) );
AND2x2_ASAP7_75t_L g651 ( .A(n_473), .B(n_496), .Y(n_651) );
AND3x2_ASAP7_75t_L g664 ( .A(n_473), .B(n_665), .C(n_666), .Y(n_664) );
INVx1_ASAP7_75t_L g587 ( .A(n_483), .Y(n_587) );
AND2x2_ASAP7_75t_L g483 ( .A(n_484), .B(n_495), .Y(n_483) );
AOI32xp33_ASAP7_75t_L g642 ( .A1(n_484), .A2(n_594), .A3(n_643), .B1(n_646), .B2(n_647), .Y(n_642) );
INVx1_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
AND2x2_ASAP7_75t_L g569 ( .A(n_485), .B(n_495), .Y(n_569) );
NAND2xp5_ASAP7_75t_SL g640 ( .A(n_485), .B(n_597), .Y(n_640) );
AND2x2_ASAP7_75t_L g647 ( .A(n_485), .B(n_619), .Y(n_647) );
OR2x2_ASAP7_75t_L g653 ( .A(n_485), .B(n_654), .Y(n_653) );
NAND2xp5_ASAP7_75t_L g678 ( .A(n_485), .B(n_608), .Y(n_678) );
OR2x2_ASAP7_75t_L g696 ( .A(n_485), .B(n_525), .Y(n_696) );
BUFx3_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
AND2x2_ASAP7_75t_L g560 ( .A(n_486), .B(n_505), .Y(n_560) );
INVx2_ASAP7_75t_L g582 ( .A(n_486), .Y(n_582) );
OR2x2_ASAP7_75t_L g604 ( .A(n_486), .B(n_505), .Y(n_604) );
AND2x2_ASAP7_75t_L g609 ( .A(n_486), .B(n_610), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g660 ( .A(n_486), .B(n_661), .Y(n_660) );
AND2x2_ASAP7_75t_L g665 ( .A(n_486), .B(n_559), .Y(n_665) );
INVx1_ASAP7_75t_SL g716 ( .A(n_495), .Y(n_716) );
AND2x2_ASAP7_75t_L g495 ( .A(n_496), .B(n_505), .Y(n_495) );
INVx1_ASAP7_75t_SL g559 ( .A(n_496), .Y(n_559) );
HB1xp67_ASAP7_75t_L g608 ( .A(n_496), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g644 ( .A(n_496), .B(n_645), .Y(n_644) );
NAND3xp33_ASAP7_75t_L g711 ( .A(n_496), .B(n_582), .C(n_700), .Y(n_711) );
INVx2_ASAP7_75t_L g610 ( .A(n_505), .Y(n_610) );
HB1xp67_ASAP7_75t_L g624 ( .A(n_505), .Y(n_624) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_514), .B(n_524), .Y(n_513) );
INVx1_ASAP7_75t_L g646 ( .A(n_514), .Y(n_646) );
INVx1_ASAP7_75t_L g514 ( .A(n_515), .Y(n_514) );
AND2x2_ASAP7_75t_L g564 ( .A(n_515), .B(n_548), .Y(n_564) );
INVx2_ASAP7_75t_L g581 ( .A(n_515), .Y(n_581) );
AND2x2_ASAP7_75t_L g586 ( .A(n_515), .B(n_549), .Y(n_586) );
AND2x2_ASAP7_75t_L g601 ( .A(n_515), .B(n_538), .Y(n_601) );
AND2x2_ASAP7_75t_L g613 ( .A(n_515), .B(n_585), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g628 ( .A(n_524), .B(n_629), .Y(n_628) );
NAND2x1p5_ASAP7_75t_L g685 ( .A(n_524), .B(n_586), .Y(n_685) );
NAND2xp5_ASAP7_75t_L g704 ( .A(n_524), .B(n_705), .Y(n_704) );
NAND2xp5_ASAP7_75t_L g708 ( .A(n_524), .B(n_580), .Y(n_708) );
BUFx3_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
OR2x2_ASAP7_75t_L g547 ( .A(n_525), .B(n_548), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g563 ( .A(n_525), .B(n_564), .Y(n_563) );
AND2x2_ASAP7_75t_L g590 ( .A(n_525), .B(n_538), .Y(n_590) );
AND2x2_ASAP7_75t_L g616 ( .A(n_525), .B(n_548), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g655 ( .A(n_525), .B(n_656), .Y(n_655) );
OA21x2_ASAP7_75t_L g525 ( .A1(n_526), .A2(n_529), .B(n_536), .Y(n_525) );
INVx1_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
AO21x2_ASAP7_75t_L g574 ( .A1(n_527), .A2(n_575), .B(n_576), .Y(n_574) );
INVx1_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
INVx1_ASAP7_75t_L g575 ( .A(n_529), .Y(n_575) );
INVx1_ASAP7_75t_L g576 ( .A(n_536), .Y(n_576) );
OR2x2_ASAP7_75t_L g537 ( .A(n_538), .B(n_547), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g566 ( .A(n_538), .B(n_567), .Y(n_566) );
AND2x4_ASAP7_75t_L g580 ( .A(n_538), .B(n_581), .Y(n_580) );
INVx3_ASAP7_75t_SL g585 ( .A(n_538), .Y(n_585) );
NAND2xp5_ASAP7_75t_L g638 ( .A(n_538), .B(n_572), .Y(n_638) );
OR2x2_ASAP7_75t_L g648 ( .A(n_538), .B(n_574), .Y(n_648) );
NAND2xp5_ASAP7_75t_L g676 ( .A(n_538), .B(n_616), .Y(n_676) );
OR2x2_ASAP7_75t_L g706 ( .A(n_538), .B(n_548), .Y(n_706) );
AND2x2_ASAP7_75t_L g710 ( .A(n_538), .B(n_549), .Y(n_710) );
NAND2xp5_ASAP7_75t_SL g723 ( .A(n_538), .B(n_586), .Y(n_723) );
AND2x2_ASAP7_75t_L g730 ( .A(n_538), .B(n_612), .Y(n_730) );
OR2x6_ASAP7_75t_L g538 ( .A(n_539), .B(n_545), .Y(n_538) );
INVx1_ASAP7_75t_SL g673 ( .A(n_547), .Y(n_673) );
AND2x2_ASAP7_75t_L g612 ( .A(n_548), .B(n_574), .Y(n_612) );
AND2x2_ASAP7_75t_L g626 ( .A(n_548), .B(n_581), .Y(n_626) );
AND2x2_ASAP7_75t_L g629 ( .A(n_548), .B(n_585), .Y(n_629) );
INVx1_ASAP7_75t_L g656 ( .A(n_548), .Y(n_656) );
INVx2_ASAP7_75t_SL g548 ( .A(n_549), .Y(n_548) );
BUFx2_ASAP7_75t_L g568 ( .A(n_549), .Y(n_568) );
NAND2xp5_ASAP7_75t_L g557 ( .A(n_558), .B(n_560), .Y(n_557) );
A2O1A1Ixp33_ASAP7_75t_L g727 ( .A1(n_558), .A2(n_604), .B(n_728), .C(n_729), .Y(n_727) );
HB1xp67_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
AND2x2_ASAP7_75t_L g634 ( .A(n_559), .B(n_635), .Y(n_634) );
NAND2xp5_ASAP7_75t_L g592 ( .A(n_560), .B(n_577), .Y(n_592) );
AND2x2_ASAP7_75t_L g618 ( .A(n_560), .B(n_619), .Y(n_618) );
OAI21xp5_ASAP7_75t_SL g561 ( .A1(n_562), .A2(n_565), .B(n_569), .Y(n_561) );
INVx1_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
NOR2xp33_ASAP7_75t_L g662 ( .A(n_563), .B(n_663), .Y(n_662) );
AND2x2_ASAP7_75t_L g589 ( .A(n_564), .B(n_590), .Y(n_589) );
NAND2xp5_ASAP7_75t_L g630 ( .A(n_564), .B(n_585), .Y(n_630) );
AND2x2_ASAP7_75t_L g721 ( .A(n_564), .B(n_572), .Y(n_721) );
INVxp67_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
INVx1_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
AND2x2_ASAP7_75t_L g594 ( .A(n_568), .B(n_581), .Y(n_594) );
OR2x2_ASAP7_75t_L g595 ( .A(n_568), .B(n_579), .Y(n_595) );
OAI322xp33_ASAP7_75t_L g570 ( .A1(n_571), .A2(n_578), .A3(n_579), .B1(n_582), .B2(n_583), .C1(n_587), .C2(n_588), .Y(n_570) );
NAND2xp5_ASAP7_75t_L g571 ( .A(n_572), .B(n_577), .Y(n_571) );
AND2x2_ASAP7_75t_L g682 ( .A(n_572), .B(n_594), .Y(n_682) );
NAND2xp5_ASAP7_75t_L g728 ( .A(n_572), .B(n_646), .Y(n_728) );
INVx2_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
INVx1_ASAP7_75t_SL g573 ( .A(n_574), .Y(n_573) );
AND2x2_ASAP7_75t_L g625 ( .A(n_574), .B(n_626), .Y(n_625) );
INVx1_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
OR2x2_ASAP7_75t_L g691 ( .A(n_578), .B(n_604), .Y(n_691) );
NAND2xp5_ASAP7_75t_L g672 ( .A(n_579), .B(n_673), .Y(n_672) );
INVx3_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g669 ( .A(n_580), .B(n_612), .Y(n_669) );
AND2x2_ASAP7_75t_L g615 ( .A(n_581), .B(n_585), .Y(n_615) );
AND2x2_ASAP7_75t_L g623 ( .A(n_582), .B(n_624), .Y(n_623) );
A2O1A1Ixp33_ASAP7_75t_L g720 ( .A1(n_582), .A2(n_661), .B(n_721), .C(n_722), .Y(n_720) );
AOI21xp33_ASAP7_75t_L g693 ( .A1(n_583), .A2(n_596), .B(n_694), .Y(n_693) );
INVx1_ASAP7_75t_SL g583 ( .A(n_584), .Y(n_583) );
AND2x2_ASAP7_75t_L g584 ( .A(n_585), .B(n_586), .Y(n_584) );
NAND2xp5_ASAP7_75t_L g652 ( .A(n_585), .B(n_612), .Y(n_652) );
AND2x2_ASAP7_75t_L g658 ( .A(n_585), .B(n_626), .Y(n_658) );
AND2x2_ASAP7_75t_L g692 ( .A(n_585), .B(n_594), .Y(n_692) );
NOR2xp33_ASAP7_75t_L g600 ( .A(n_586), .B(n_601), .Y(n_600) );
INVx2_ASAP7_75t_SL g702 ( .A(n_586), .Y(n_702) );
INVx1_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
AOI22xp5_ASAP7_75t_L g617 ( .A1(n_590), .A2(n_618), .B1(n_620), .B2(n_625), .Y(n_617) );
OAI22xp5_ASAP7_75t_SL g591 ( .A1(n_592), .A2(n_593), .B1(n_595), .B2(n_596), .Y(n_591) );
OAI22xp33_ASAP7_75t_L g627 ( .A1(n_592), .A2(n_628), .B1(n_630), .B2(n_631), .Y(n_627) );
INVxp67_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
INVx1_ASAP7_75t_SL g596 ( .A(n_597), .Y(n_596) );
AOI221xp5_ASAP7_75t_L g698 ( .A1(n_597), .A2(n_699), .B1(n_701), .B2(n_703), .C(n_707), .Y(n_698) );
AOI211xp5_ASAP7_75t_L g598 ( .A1(n_599), .A2(n_602), .B(n_606), .C(n_627), .Y(n_598) );
INVxp67_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
INVx1_ASAP7_75t_L g602 ( .A(n_603), .Y(n_602) );
OR2x2_ASAP7_75t_L g603 ( .A(n_604), .B(n_605), .Y(n_603) );
OR2x2_ASAP7_75t_L g668 ( .A(n_604), .B(n_621), .Y(n_668) );
INVx1_ASAP7_75t_L g719 ( .A(n_604), .Y(n_719) );
OAI221xp5_ASAP7_75t_L g606 ( .A1(n_605), .A2(n_607), .B1(n_611), .B2(n_614), .C(n_617), .Y(n_606) );
INVx2_ASAP7_75t_SL g661 ( .A(n_605), .Y(n_661) );
NAND2xp5_ASAP7_75t_L g607 ( .A(n_608), .B(n_609), .Y(n_607) );
INVx1_ASAP7_75t_L g726 ( .A(n_608), .Y(n_726) );
AND2x2_ASAP7_75t_L g650 ( .A(n_609), .B(n_651), .Y(n_650) );
INVx2_ASAP7_75t_L g635 ( .A(n_610), .Y(n_635) );
NAND2xp5_ASAP7_75t_L g611 ( .A(n_612), .B(n_613), .Y(n_611) );
INVx1_ASAP7_75t_L g697 ( .A(n_613), .Y(n_697) );
NAND2xp5_ASAP7_75t_L g614 ( .A(n_615), .B(n_616), .Y(n_614) );
AND2x2_ASAP7_75t_L g620 ( .A(n_621), .B(n_623), .Y(n_620) );
NOR2xp33_ASAP7_75t_L g722 ( .A(n_621), .B(n_723), .Y(n_722) );
CKINVDCx16_ASAP7_75t_R g621 ( .A(n_622), .Y(n_621) );
INVxp67_ASAP7_75t_L g666 ( .A(n_624), .Y(n_666) );
O2A1O1Ixp33_ASAP7_75t_L g636 ( .A1(n_625), .A2(n_637), .B(n_639), .C(n_641), .Y(n_636) );
INVx1_ASAP7_75t_L g714 ( .A(n_628), .Y(n_714) );
INVx1_ASAP7_75t_L g631 ( .A(n_632), .Y(n_631) );
NOR2xp33_ASAP7_75t_L g689 ( .A(n_632), .B(n_690), .Y(n_689) );
AND2x2_ASAP7_75t_L g632 ( .A(n_633), .B(n_634), .Y(n_632) );
INVx2_ASAP7_75t_L g645 ( .A(n_635), .Y(n_645) );
INVx1_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
INVx1_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
OAI222xp33_ASAP7_75t_L g641 ( .A1(n_642), .A2(n_648), .B1(n_649), .B2(n_652), .C1(n_653), .C2(n_655), .Y(n_641) );
INVx1_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
INVx1_ASAP7_75t_SL g681 ( .A(n_645), .Y(n_681) );
NOR2xp33_ASAP7_75t_L g701 ( .A(n_648), .B(n_702), .Y(n_701) );
NAND2xp33_ASAP7_75t_SL g679 ( .A(n_649), .B(n_680), .Y(n_679) );
INVx1_ASAP7_75t_SL g649 ( .A(n_650), .Y(n_649) );
INVx1_ASAP7_75t_SL g654 ( .A(n_651), .Y(n_654) );
AND2x2_ASAP7_75t_L g718 ( .A(n_651), .B(n_719), .Y(n_718) );
OR2x2_ASAP7_75t_L g684 ( .A(n_654), .B(n_681), .Y(n_684) );
INVx1_ASAP7_75t_L g713 ( .A(n_655), .Y(n_713) );
AOI211xp5_ASAP7_75t_L g657 ( .A1(n_658), .A2(n_659), .B(n_662), .C(n_667), .Y(n_657) );
INVx1_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
NAND2xp5_ASAP7_75t_L g680 ( .A(n_661), .B(n_681), .Y(n_680) );
INVx2_ASAP7_75t_SL g663 ( .A(n_664), .Y(n_663) );
AOI322xp5_ASAP7_75t_L g712 ( .A1(n_664), .A2(n_692), .A3(n_697), .B1(n_713), .B2(n_714), .C1(n_715), .C2(n_718), .Y(n_712) );
AND2x2_ASAP7_75t_L g699 ( .A(n_665), .B(n_700), .Y(n_699) );
OAI22xp33_ASAP7_75t_L g667 ( .A1(n_668), .A2(n_669), .B1(n_670), .B2(n_672), .Y(n_667) );
INVxp33_ASAP7_75t_L g670 ( .A(n_671), .Y(n_670) );
AOI221xp5_ASAP7_75t_L g674 ( .A1(n_675), .A2(n_677), .B1(n_679), .B2(n_682), .C(n_683), .Y(n_674) );
INVx1_ASAP7_75t_L g675 ( .A(n_676), .Y(n_675) );
INVx1_ASAP7_75t_L g677 ( .A(n_678), .Y(n_677) );
NOR2xp33_ASAP7_75t_L g683 ( .A(n_684), .B(n_685), .Y(n_683) );
NAND5xp2_ASAP7_75t_L g686 ( .A(n_687), .B(n_698), .C(n_712), .D(n_720), .E(n_724), .Y(n_686) );
AOI21xp5_ASAP7_75t_L g687 ( .A1(n_688), .A2(n_692), .B(n_693), .Y(n_687) );
INVxp67_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
INVx2_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
INVxp33_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
NOR2xp33_ASAP7_75t_L g695 ( .A(n_696), .B(n_697), .Y(n_695) );
A2O1A1Ixp33_ASAP7_75t_L g724 ( .A1(n_700), .A2(n_725), .B(n_726), .C(n_727), .Y(n_724) );
AOI31xp33_ASAP7_75t_L g707 ( .A1(n_702), .A2(n_708), .A3(n_709), .B(n_711), .Y(n_707) );
INVx1_ASAP7_75t_L g703 ( .A(n_704), .Y(n_703) );
INVx1_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
INVx1_ASAP7_75t_L g709 ( .A(n_710), .Y(n_709) );
NOR2xp33_ASAP7_75t_L g715 ( .A(n_716), .B(n_717), .Y(n_715) );
INVx1_ASAP7_75t_L g725 ( .A(n_723), .Y(n_725) );
INVx1_ASAP7_75t_L g729 ( .A(n_730), .Y(n_729) );
INVx2_ASAP7_75t_L g731 ( .A(n_732), .Y(n_731) );
INVx2_ASAP7_75t_L g747 ( .A(n_732), .Y(n_747) );
INVx1_ASAP7_75t_L g732 ( .A(n_733), .Y(n_732) );
INVx1_ASAP7_75t_L g735 ( .A(n_736), .Y(n_735) );
CKINVDCx20_ASAP7_75t_R g738 ( .A(n_739), .Y(n_738) );
INVx1_ASAP7_75t_L g743 ( .A(n_740), .Y(n_743) );
INVx1_ASAP7_75t_SL g748 ( .A(n_749), .Y(n_748) );
INVx3_ASAP7_75t_SL g749 ( .A(n_750), .Y(n_749) );
INVx1_ASAP7_75t_SL g751 ( .A(n_752), .Y(n_751) );
endmodule