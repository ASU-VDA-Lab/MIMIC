module fake_jpeg_21588_n_39 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_39);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_39;

wire n_21;
wire n_33;
wire n_23;
wire n_27;
wire n_22;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_34;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_36;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_32;

INVx1_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_12),
.Y(n_17)
);

INVx4_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_15),
.B(n_11),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

OAI22xp5_ASAP7_75t_SL g22 ( 
.A1(n_19),
.A2(n_18),
.B1(n_17),
.B2(n_16),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_22),
.B(n_23),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_SL g23 ( 
.A(n_19),
.B(n_0),
.Y(n_23)
);

AOI22xp33_ASAP7_75t_L g24 ( 
.A1(n_18),
.A2(n_6),
.B1(n_13),
.B2(n_10),
.Y(n_24)
);

OAI21xp5_ASAP7_75t_L g27 ( 
.A1(n_24),
.A2(n_25),
.B(n_26),
.Y(n_27)
);

AND2x2_ASAP7_75t_L g25 ( 
.A(n_20),
.B(n_0),
.Y(n_25)
);

AOI22xp33_ASAP7_75t_L g26 ( 
.A1(n_21),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_25),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_28),
.B(n_29),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_24),
.Y(n_29)
);

AOI21xp5_ASAP7_75t_L g31 ( 
.A1(n_27),
.A2(n_30),
.B(n_8),
.Y(n_31)
);

AOI21xp5_ASAP7_75t_L g35 ( 
.A1(n_31),
.A2(n_14),
.B(n_5),
.Y(n_35)
);

MAJIxp5_ASAP7_75t_L g32 ( 
.A(n_27),
.B(n_20),
.C(n_21),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_SL g34 ( 
.A1(n_32),
.A2(n_20),
.B1(n_4),
.B2(n_3),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_34),
.B(n_35),
.Y(n_36)
);

INVxp33_ASAP7_75t_L g37 ( 
.A(n_36),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_37),
.B(n_33),
.Y(n_38)
);

XNOR2xp5_ASAP7_75t_L g39 ( 
.A(n_38),
.B(n_7),
.Y(n_39)
);


endmodule