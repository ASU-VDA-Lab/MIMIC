module fake_jpeg_31632_n_84 (n_13, n_21, n_1, n_10, n_23, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_9, n_5, n_11, n_17, n_25, n_2, n_12, n_8, n_15, n_7, n_84);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_84;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_57;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_44;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_35;
wire n_48;
wire n_46;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_21),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_22),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_17),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_20),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_24),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_11),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_26),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_33),
.B(n_0),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_36),
.B(n_37),
.Y(n_42)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_30),
.Y(n_37)
);

BUFx2_ASAP7_75t_L g38 ( 
.A(n_26),
.Y(n_38)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_38),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_28),
.B(n_0),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_39),
.B(n_1),
.Y(n_48)
);

HB1xp67_ASAP7_75t_L g40 ( 
.A(n_27),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_40),
.B(n_31),
.Y(n_46)
);

AND2x2_ASAP7_75t_SL g41 ( 
.A(n_40),
.B(n_27),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_41),
.B(n_45),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_38),
.Y(n_44)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_44),
.Y(n_50)
);

AOI21xp5_ASAP7_75t_L g45 ( 
.A1(n_37),
.A2(n_34),
.B(n_32),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_46),
.B(n_48),
.Y(n_56)
);

INVx11_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_49),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_43),
.Y(n_52)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_52),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_41),
.A2(n_31),
.B1(n_29),
.B2(n_3),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_53),
.A2(n_55),
.B1(n_4),
.B2(n_5),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_44),
.A2(n_43),
.B1(n_47),
.B2(n_3),
.Y(n_55)
);

INVx1_ASAP7_75t_SL g57 ( 
.A(n_47),
.Y(n_57)
);

OR2x2_ASAP7_75t_L g64 ( 
.A(n_57),
.B(n_4),
.Y(n_64)
);

CKINVDCx16_ASAP7_75t_R g58 ( 
.A(n_42),
.Y(n_58)
);

INVxp67_ASAP7_75t_L g59 ( 
.A(n_58),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g60 ( 
.A(n_56),
.B(n_42),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_60),
.B(n_62),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_SL g61 ( 
.A(n_54),
.B(n_1),
.C(n_2),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_61),
.B(n_67),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_54),
.B(n_2),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_63),
.A2(n_10),
.B1(n_12),
.B2(n_13),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_64),
.Y(n_70)
);

XNOR2xp5_ASAP7_75t_L g66 ( 
.A(n_55),
.B(n_16),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_66),
.B(n_68),
.C(n_59),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_50),
.B(n_5),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_51),
.B(n_7),
.C(n_8),
.Y(n_68)
);

INVxp67_ASAP7_75t_L g75 ( 
.A(n_69),
.Y(n_75)
);

OAI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_59),
.A2(n_15),
.B1(n_18),
.B2(n_19),
.Y(n_72)
);

XNOR2xp5_ASAP7_75t_SL g76 ( 
.A(n_72),
.B(n_73),
.Y(n_76)
);

AND2x2_ASAP7_75t_SL g77 ( 
.A(n_76),
.B(n_70),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_77),
.Y(n_78)
);

OAI21xp5_ASAP7_75t_L g79 ( 
.A1(n_78),
.A2(n_71),
.B(n_74),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_79),
.A2(n_75),
.B1(n_64),
.B2(n_72),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_80),
.B(n_23),
.Y(n_81)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_81),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_82),
.B(n_65),
.Y(n_83)
);

XNOR2xp5_ASAP7_75t_L g84 ( 
.A(n_83),
.B(n_25),
.Y(n_84)
);


endmodule