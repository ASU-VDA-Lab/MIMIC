module fake_aes_12640_n_347 (n_45, n_20, n_2, n_38, n_44, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_28, n_31, n_22, n_46, n_11, n_25, n_16, n_26, n_13, n_30, n_33, n_3, n_18, n_32, n_0, n_41, n_1, n_35, n_12, n_9, n_17, n_14, n_10, n_15, n_42, n_24, n_19, n_21, n_6, n_4, n_29, n_43, n_7, n_40, n_27, n_39, n_347);
input n_45;
input n_20;
input n_2;
input n_38;
input n_44;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_28;
input n_31;
input n_22;
input n_46;
input n_11;
input n_25;
input n_16;
input n_26;
input n_13;
input n_30;
input n_33;
input n_3;
input n_18;
input n_32;
input n_0;
input n_41;
input n_1;
input n_35;
input n_12;
input n_9;
input n_17;
input n_14;
input n_10;
input n_15;
input n_42;
input n_24;
input n_19;
input n_21;
input n_6;
input n_4;
input n_29;
input n_43;
input n_7;
input n_40;
input n_27;
input n_39;
output n_347;
wire n_117;
wire n_185;
wire n_57;
wire n_284;
wire n_278;
wire n_60;
wire n_114;
wire n_94;
wire n_125;
wire n_161;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_154;
wire n_328;
wire n_229;
wire n_336;
wire n_252;
wire n_152;
wire n_113;
wire n_206;
wire n_288;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_142;
wire n_232;
wire n_316;
wire n_211;
wire n_334;
wire n_275;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_162;
wire n_163;
wire n_105;
wire n_227;
wire n_231;
wire n_298;
wire n_144;
wire n_53;
wire n_183;
wire n_199;
wire n_83;
wire n_100;
wire n_48;
wire n_305;
wire n_228;
wire n_345;
wire n_236;
wire n_340;
wire n_150;
wire n_301;
wire n_66;
wire n_222;
wire n_234;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_324;
wire n_279;
wire n_303;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_244;
wire n_50;
wire n_73;
wire n_49;
wire n_119;
wire n_141;
wire n_97;
wire n_167;
wire n_171;
wire n_65;
wire n_196;
wire n_192;
wire n_312;
wire n_137;
wire n_277;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_62;
wire n_255;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_241;
wire n_95;
wire n_238;
wire n_318;
wire n_293;
wire n_135;
wire n_247;
wire n_304;
wire n_294;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_235;
wire n_243;
wire n_331;
wire n_268;
wire n_174;
wire n_248;
wire n_72;
wire n_299;
wire n_89;
wire n_338;
wire n_256;
wire n_67;
wire n_77;
wire n_54;
wire n_172;
wire n_329;
wire n_251;
wire n_59;
wire n_218;
wire n_271;
wire n_302;
wire n_270;
wire n_153;
wire n_61;
wire n_259;
wire n_308;
wire n_93;
wire n_140;
wire n_207;
wire n_224;
wire n_96;
wire n_219;
wire n_133;
wire n_149;
wire n_81;
wire n_69;
wire n_214;
wire n_204;
wire n_88;
wire n_107;
wire n_254;
wire n_262;
wire n_239;
wire n_87;
wire n_98;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_342;
wire n_217;
wire n_139;
wire n_193;
wire n_273;
wire n_120;
wire n_70;
wire n_245;
wire n_90;
wire n_260;
wire n_78;
wire n_197;
wire n_201;
wire n_317;
wire n_111;
wire n_64;
wire n_265;
wire n_264;
wire n_200;
wire n_208;
wire n_126;
wire n_178;
wire n_118;
wire n_179;
wire n_315;
wire n_86;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_186;
wire n_75;
wire n_344;
wire n_136;
wire n_283;
wire n_76;
wire n_216;
wire n_147;
wire n_148;
wire n_212;
wire n_92;
wire n_168;
wire n_134;
wire n_233;
wire n_82;
wire n_106;
wire n_173;
wire n_327;
wire n_325;
wire n_51;
wire n_225;
wire n_220;
wire n_267;
wire n_221;
wire n_203;
wire n_52;
wire n_102;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_121;
wire n_339;
wire n_240;
wire n_346;
wire n_103;
wire n_180;
wire n_104;
wire n_74;
wire n_335;
wire n_272;
wire n_146;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_198;
wire n_169;
wire n_156;
wire n_124;
wire n_297;
wire n_128;
wire n_129;
wire n_63;
wire n_71;
wire n_56;
wire n_188;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_281;
wire n_341;
wire n_58;
wire n_122;
wire n_187;
wire n_138;
wire n_323;
wire n_258;
wire n_253;
wire n_84;
wire n_266;
wire n_55;
wire n_213;
wire n_182;
wire n_226;
wire n_159;
wire n_337;
wire n_176;
wire n_68;
wire n_123;
wire n_223;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_332;
wire n_164;
wire n_175;
wire n_145;
wire n_290;
wire n_280;
wire n_99;
wire n_109;
wire n_132;
wire n_151;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g48 ( .A(n_36), .Y(n_48) );
HB1xp67_ASAP7_75t_L g49 ( .A(n_3), .Y(n_49) );
INVx1_ASAP7_75t_L g50 ( .A(n_10), .Y(n_50) );
BUFx2_ASAP7_75t_L g51 ( .A(n_46), .Y(n_51) );
INVxp33_ASAP7_75t_L g52 ( .A(n_21), .Y(n_52) );
INVx1_ASAP7_75t_L g53 ( .A(n_33), .Y(n_53) );
INVx1_ASAP7_75t_L g54 ( .A(n_16), .Y(n_54) );
INVxp33_ASAP7_75t_SL g55 ( .A(n_5), .Y(n_55) );
INVx1_ASAP7_75t_L g56 ( .A(n_18), .Y(n_56) );
INVx1_ASAP7_75t_L g57 ( .A(n_31), .Y(n_57) );
INVxp33_ASAP7_75t_L g58 ( .A(n_40), .Y(n_58) );
CKINVDCx16_ASAP7_75t_R g59 ( .A(n_29), .Y(n_59) );
INVxp67_ASAP7_75t_L g60 ( .A(n_18), .Y(n_60) );
INVx1_ASAP7_75t_L g61 ( .A(n_7), .Y(n_61) );
CKINVDCx5p33_ASAP7_75t_R g62 ( .A(n_42), .Y(n_62) );
INVxp33_ASAP7_75t_L g63 ( .A(n_13), .Y(n_63) );
BUFx6f_ASAP7_75t_L g64 ( .A(n_5), .Y(n_64) );
INVx1_ASAP7_75t_L g65 ( .A(n_43), .Y(n_65) );
INVx1_ASAP7_75t_L g66 ( .A(n_34), .Y(n_66) );
BUFx3_ASAP7_75t_L g67 ( .A(n_35), .Y(n_67) );
CKINVDCx16_ASAP7_75t_R g68 ( .A(n_30), .Y(n_68) );
BUFx3_ASAP7_75t_L g69 ( .A(n_45), .Y(n_69) );
INVx1_ASAP7_75t_L g70 ( .A(n_19), .Y(n_70) );
INVx1_ASAP7_75t_L g71 ( .A(n_47), .Y(n_71) );
INVxp67_ASAP7_75t_L g72 ( .A(n_11), .Y(n_72) );
INVx1_ASAP7_75t_L g73 ( .A(n_1), .Y(n_73) );
INVxp67_ASAP7_75t_L g74 ( .A(n_26), .Y(n_74) );
INVx1_ASAP7_75t_L g75 ( .A(n_2), .Y(n_75) );
BUFx2_ASAP7_75t_L g76 ( .A(n_2), .Y(n_76) );
INVxp67_ASAP7_75t_L g77 ( .A(n_22), .Y(n_77) );
INVx1_ASAP7_75t_L g78 ( .A(n_25), .Y(n_78) );
CKINVDCx16_ASAP7_75t_R g79 ( .A(n_44), .Y(n_79) );
CKINVDCx5p33_ASAP7_75t_R g80 ( .A(n_32), .Y(n_80) );
INVx1_ASAP7_75t_L g81 ( .A(n_38), .Y(n_81) );
INVx2_ASAP7_75t_L g82 ( .A(n_67), .Y(n_82) );
NAND2xp5_ASAP7_75t_SL g83 ( .A(n_51), .B(n_0), .Y(n_83) );
BUFx3_ASAP7_75t_L g84 ( .A(n_67), .Y(n_84) );
CKINVDCx5p33_ASAP7_75t_R g85 ( .A(n_59), .Y(n_85) );
INVx2_ASAP7_75t_L g86 ( .A(n_67), .Y(n_86) );
CKINVDCx5p33_ASAP7_75t_R g87 ( .A(n_68), .Y(n_87) );
BUFx3_ASAP7_75t_L g88 ( .A(n_69), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_48), .Y(n_89) );
CKINVDCx5p33_ASAP7_75t_R g90 ( .A(n_68), .Y(n_90) );
INVx2_ASAP7_75t_L g91 ( .A(n_69), .Y(n_91) );
CKINVDCx5p33_ASAP7_75t_R g92 ( .A(n_79), .Y(n_92) );
CKINVDCx5p33_ASAP7_75t_R g93 ( .A(n_79), .Y(n_93) );
NOR2xp33_ASAP7_75t_L g94 ( .A(n_51), .B(n_0), .Y(n_94) );
INVxp33_ASAP7_75t_SL g95 ( .A(n_49), .Y(n_95) );
INVx2_ASAP7_75t_L g96 ( .A(n_69), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_48), .Y(n_97) );
INVx2_ASAP7_75t_L g98 ( .A(n_53), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_53), .Y(n_99) );
CKINVDCx5p33_ASAP7_75t_R g100 ( .A(n_76), .Y(n_100) );
CKINVDCx5p33_ASAP7_75t_R g101 ( .A(n_76), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_98), .Y(n_102) );
NAND2xp5_ASAP7_75t_L g103 ( .A(n_89), .B(n_57), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_98), .Y(n_104) );
BUFx3_ASAP7_75t_L g105 ( .A(n_84), .Y(n_105) );
AO22x2_ASAP7_75t_L g106 ( .A1(n_83), .A2(n_81), .B1(n_78), .B2(n_66), .Y(n_106) );
AOI22xp33_ASAP7_75t_L g107 ( .A1(n_89), .A2(n_50), .B1(n_54), .B2(n_56), .Y(n_107) );
NAND2xp5_ASAP7_75t_L g108 ( .A(n_97), .B(n_57), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_98), .Y(n_109) );
NAND2xp5_ASAP7_75t_L g110 ( .A(n_97), .B(n_65), .Y(n_110) );
AND3x4_ASAP7_75t_L g111 ( .A(n_95), .B(n_55), .C(n_63), .Y(n_111) );
AND2x2_ASAP7_75t_L g112 ( .A(n_99), .B(n_52), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_82), .Y(n_113) );
CKINVDCx5p33_ASAP7_75t_R g114 ( .A(n_85), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_82), .Y(n_115) );
BUFx3_ASAP7_75t_L g116 ( .A(n_84), .Y(n_116) );
INVx2_ASAP7_75t_L g117 ( .A(n_84), .Y(n_117) );
AND2x2_ASAP7_75t_SL g118 ( .A(n_94), .B(n_65), .Y(n_118) );
INVx2_ASAP7_75t_L g119 ( .A(n_88), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_82), .Y(n_120) );
AND2x2_ASAP7_75t_L g121 ( .A(n_99), .B(n_58), .Y(n_121) );
BUFx6f_ASAP7_75t_L g122 ( .A(n_88), .Y(n_122) );
INVx2_ASAP7_75t_L g123 ( .A(n_88), .Y(n_123) );
INVx2_ASAP7_75t_L g124 ( .A(n_86), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_86), .Y(n_125) );
AO21x2_ASAP7_75t_L g126 ( .A1(n_103), .A2(n_83), .B(n_81), .Y(n_126) );
INVx1_ASAP7_75t_L g127 ( .A(n_102), .Y(n_127) );
O2A1O1Ixp33_ASAP7_75t_L g128 ( .A1(n_103), .A2(n_94), .B(n_60), .C(n_72), .Y(n_128) );
OAI22xp5_ASAP7_75t_L g129 ( .A1(n_118), .A2(n_101), .B1(n_100), .B2(n_85), .Y(n_129) );
NOR2xp33_ASAP7_75t_R g130 ( .A(n_114), .B(n_87), .Y(n_130) );
AOI21xp5_ASAP7_75t_L g131 ( .A1(n_117), .A2(n_91), .B(n_86), .Y(n_131) );
INVx1_ASAP7_75t_L g132 ( .A(n_102), .Y(n_132) );
INVx1_ASAP7_75t_SL g133 ( .A(n_112), .Y(n_133) );
NAND2xp5_ASAP7_75t_SL g134 ( .A(n_118), .B(n_95), .Y(n_134) );
INVx2_ASAP7_75t_L g135 ( .A(n_122), .Y(n_135) );
AOI21xp5_ASAP7_75t_L g136 ( .A1(n_117), .A2(n_96), .B(n_91), .Y(n_136) );
O2A1O1Ixp33_ASAP7_75t_SL g137 ( .A1(n_108), .A2(n_110), .B(n_125), .C(n_113), .Y(n_137) );
A2O1A1Ixp33_ASAP7_75t_L g138 ( .A1(n_104), .A2(n_96), .B(n_71), .C(n_78), .Y(n_138) );
AND2x4_ASAP7_75t_L g139 ( .A(n_112), .B(n_50), .Y(n_139) );
OAI22xp5_ASAP7_75t_L g140 ( .A1(n_118), .A2(n_90), .B1(n_93), .B2(n_92), .Y(n_140) );
INVx2_ASAP7_75t_L g141 ( .A(n_122), .Y(n_141) );
AOI21xp5_ASAP7_75t_L g142 ( .A1(n_117), .A2(n_71), .B(n_74), .Y(n_142) );
INVx2_ASAP7_75t_L g143 ( .A(n_122), .Y(n_143) );
NAND2xp5_ASAP7_75t_L g144 ( .A(n_121), .B(n_80), .Y(n_144) );
OAI21xp33_ASAP7_75t_L g145 ( .A1(n_121), .A2(n_56), .B(n_75), .Y(n_145) );
NAND3xp33_ASAP7_75t_SL g146 ( .A(n_111), .B(n_62), .C(n_77), .Y(n_146) );
NAND2xp5_ASAP7_75t_SL g147 ( .A(n_118), .B(n_64), .Y(n_147) );
AND2x4_ASAP7_75t_L g148 ( .A(n_121), .B(n_75), .Y(n_148) );
NOR2xp33_ASAP7_75t_L g149 ( .A(n_110), .B(n_73), .Y(n_149) );
OAI21x1_ASAP7_75t_L g150 ( .A1(n_147), .A2(n_124), .B(n_119), .Y(n_150) );
INVx2_ASAP7_75t_L g151 ( .A(n_135), .Y(n_151) );
OAI21xp5_ASAP7_75t_L g152 ( .A1(n_147), .A2(n_123), .B(n_119), .Y(n_152) );
NOR2x1_ASAP7_75t_SL g153 ( .A(n_126), .B(n_109), .Y(n_153) );
OAI21x1_ASAP7_75t_L g154 ( .A1(n_135), .A2(n_124), .B(n_123), .Y(n_154) );
AO21x2_ASAP7_75t_L g155 ( .A1(n_137), .A2(n_115), .B(n_120), .Y(n_155) );
INVx1_ASAP7_75t_L g156 ( .A(n_127), .Y(n_156) );
AND2x2_ASAP7_75t_L g157 ( .A(n_133), .B(n_106), .Y(n_157) );
BUFx2_ASAP7_75t_L g158 ( .A(n_130), .Y(n_158) );
INVx2_ASAP7_75t_L g159 ( .A(n_141), .Y(n_159) );
INVx1_ASAP7_75t_L g160 ( .A(n_132), .Y(n_160) );
AOI21xp5_ASAP7_75t_L g161 ( .A1(n_141), .A2(n_119), .B(n_123), .Y(n_161) );
OAI21x1_ASAP7_75t_L g162 ( .A1(n_143), .A2(n_124), .B(n_120), .Y(n_162) );
INVx2_ASAP7_75t_L g163 ( .A(n_143), .Y(n_163) );
AND2x2_ASAP7_75t_SL g164 ( .A(n_139), .B(n_109), .Y(n_164) );
INVx1_ASAP7_75t_L g165 ( .A(n_138), .Y(n_165) );
OAI21x1_ASAP7_75t_L g166 ( .A1(n_131), .A2(n_107), .B(n_70), .Y(n_166) );
INVx2_ASAP7_75t_L g167 ( .A(n_126), .Y(n_167) );
AO31x2_ASAP7_75t_L g168 ( .A1(n_149), .A2(n_73), .A3(n_70), .B(n_61), .Y(n_168) );
AND2x2_ASAP7_75t_L g169 ( .A(n_134), .B(n_106), .Y(n_169) );
OAI21x1_ASAP7_75t_L g170 ( .A1(n_136), .A2(n_142), .B(n_128), .Y(n_170) );
NAND2xp5_ASAP7_75t_L g171 ( .A(n_139), .B(n_106), .Y(n_171) );
NAND2x1p5_ASAP7_75t_L g172 ( .A(n_139), .B(n_116), .Y(n_172) );
OR2x6_ASAP7_75t_L g173 ( .A(n_134), .B(n_106), .Y(n_173) );
AOI22xp5_ASAP7_75t_L g174 ( .A1(n_146), .A2(n_111), .B1(n_106), .B2(n_64), .Y(n_174) );
BUFx2_ASAP7_75t_L g175 ( .A(n_130), .Y(n_175) );
A2O1A1Ixp33_ASAP7_75t_L g176 ( .A1(n_145), .A2(n_116), .B(n_105), .C(n_64), .Y(n_176) );
BUFx6f_ASAP7_75t_L g177 ( .A(n_164), .Y(n_177) );
BUFx3_ASAP7_75t_L g178 ( .A(n_164), .Y(n_178) );
AO31x2_ASAP7_75t_L g179 ( .A1(n_153), .A2(n_129), .A3(n_144), .B(n_140), .Y(n_179) );
AND2x4_ASAP7_75t_L g180 ( .A(n_158), .B(n_148), .Y(n_180) );
INVx1_ASAP7_75t_L g181 ( .A(n_156), .Y(n_181) );
CKINVDCx16_ASAP7_75t_R g182 ( .A(n_158), .Y(n_182) );
HB1xp67_ASAP7_75t_L g183 ( .A(n_164), .Y(n_183) );
CKINVDCx11_ASAP7_75t_R g184 ( .A(n_175), .Y(n_184) );
AND2x2_ASAP7_75t_L g185 ( .A(n_164), .B(n_116), .Y(n_185) );
AND2x2_ASAP7_75t_L g186 ( .A(n_156), .B(n_105), .Y(n_186) );
INVx4_ASAP7_75t_L g187 ( .A(n_172), .Y(n_187) );
NAND2xp33_ASAP7_75t_R g188 ( .A(n_175), .B(n_1), .Y(n_188) );
NAND3xp33_ASAP7_75t_SL g189 ( .A(n_174), .B(n_64), .C(n_4), .Y(n_189) );
OR2x6_ASAP7_75t_L g190 ( .A(n_172), .B(n_64), .Y(n_190) );
INVx2_ASAP7_75t_L g191 ( .A(n_162), .Y(n_191) );
NOR3xp33_ASAP7_75t_SL g192 ( .A(n_171), .B(n_3), .C(n_6), .Y(n_192) );
INVx2_ASAP7_75t_L g193 ( .A(n_162), .Y(n_193) );
OAI21xp5_ASAP7_75t_SL g194 ( .A1(n_157), .A2(n_122), .B(n_9), .Y(n_194) );
NOR2xp33_ASAP7_75t_R g195 ( .A(n_157), .B(n_8), .Y(n_195) );
AND2x2_ASAP7_75t_L g196 ( .A(n_183), .B(n_160), .Y(n_196) );
INVx1_ASAP7_75t_L g197 ( .A(n_181), .Y(n_197) );
INVx2_ASAP7_75t_L g198 ( .A(n_191), .Y(n_198) );
INVx3_ASAP7_75t_L g199 ( .A(n_187), .Y(n_199) );
INVx1_ASAP7_75t_L g200 ( .A(n_191), .Y(n_200) );
AOI22xp33_ASAP7_75t_SL g201 ( .A1(n_195), .A2(n_157), .B1(n_169), .B2(n_173), .Y(n_201) );
OA21x2_ASAP7_75t_L g202 ( .A1(n_193), .A2(n_167), .B(n_150), .Y(n_202) );
NAND4xp25_ASAP7_75t_L g203 ( .A(n_188), .B(n_169), .C(n_165), .D(n_176), .Y(n_203) );
OA21x2_ASAP7_75t_L g204 ( .A1(n_193), .A2(n_167), .B(n_150), .Y(n_204) );
INVx1_ASAP7_75t_L g205 ( .A(n_193), .Y(n_205) );
INVx1_ASAP7_75t_L g206 ( .A(n_186), .Y(n_206) );
HB1xp67_ASAP7_75t_L g207 ( .A(n_190), .Y(n_207) );
INVx1_ASAP7_75t_SL g208 ( .A(n_190), .Y(n_208) );
AND2x4_ASAP7_75t_L g209 ( .A(n_187), .B(n_173), .Y(n_209) );
AOI211x1_ASAP7_75t_SL g210 ( .A1(n_189), .A2(n_152), .B(n_161), .C(n_168), .Y(n_210) );
AND2x4_ASAP7_75t_L g211 ( .A(n_187), .B(n_173), .Y(n_211) );
AND2x4_ASAP7_75t_L g212 ( .A(n_187), .B(n_173), .Y(n_212) );
INVx1_ASAP7_75t_L g213 ( .A(n_186), .Y(n_213) );
INVx2_ASAP7_75t_L g214 ( .A(n_198), .Y(n_214) );
INVx1_ASAP7_75t_L g215 ( .A(n_197), .Y(n_215) );
AND2x4_ASAP7_75t_L g216 ( .A(n_199), .B(n_190), .Y(n_216) );
INVx1_ASAP7_75t_L g217 ( .A(n_200), .Y(n_217) );
AND2x2_ASAP7_75t_L g218 ( .A(n_196), .B(n_183), .Y(n_218) );
INVx1_ASAP7_75t_L g219 ( .A(n_200), .Y(n_219) );
AND2x2_ASAP7_75t_L g220 ( .A(n_196), .B(n_178), .Y(n_220) );
INVx2_ASAP7_75t_L g221 ( .A(n_205), .Y(n_221) );
AND2x2_ASAP7_75t_L g222 ( .A(n_206), .B(n_178), .Y(n_222) );
INVx1_ASAP7_75t_L g223 ( .A(n_206), .Y(n_223) );
INVx1_ASAP7_75t_L g224 ( .A(n_213), .Y(n_224) );
INVx1_ASAP7_75t_L g225 ( .A(n_213), .Y(n_225) );
INVx2_ASAP7_75t_L g226 ( .A(n_202), .Y(n_226) );
INVx1_ASAP7_75t_L g227 ( .A(n_207), .Y(n_227) );
AND2x2_ASAP7_75t_L g228 ( .A(n_199), .B(n_178), .Y(n_228) );
INVx2_ASAP7_75t_L g229 ( .A(n_226), .Y(n_229) );
INVx1_ASAP7_75t_L g230 ( .A(n_217), .Y(n_230) );
INVx1_ASAP7_75t_L g231 ( .A(n_217), .Y(n_231) );
OR2x2_ASAP7_75t_L g232 ( .A(n_221), .B(n_194), .Y(n_232) );
INVx2_ASAP7_75t_L g233 ( .A(n_226), .Y(n_233) );
AND2x2_ASAP7_75t_L g234 ( .A(n_221), .B(n_202), .Y(n_234) );
INVx1_ASAP7_75t_L g235 ( .A(n_219), .Y(n_235) );
AND2x2_ASAP7_75t_L g236 ( .A(n_221), .B(n_202), .Y(n_236) );
AND2x2_ASAP7_75t_L g237 ( .A(n_214), .B(n_202), .Y(n_237) );
INVx1_ASAP7_75t_L g238 ( .A(n_219), .Y(n_238) );
NAND2xp5_ASAP7_75t_L g239 ( .A(n_215), .B(n_210), .Y(n_239) );
OR2x2_ASAP7_75t_L g240 ( .A(n_227), .B(n_207), .Y(n_240) );
INVx1_ASAP7_75t_SL g241 ( .A(n_216), .Y(n_241) );
NAND2xp5_ASAP7_75t_L g242 ( .A(n_215), .B(n_210), .Y(n_242) );
INVx2_ASAP7_75t_L g243 ( .A(n_226), .Y(n_243) );
HB1xp67_ASAP7_75t_L g244 ( .A(n_214), .Y(n_244) );
NAND2xp5_ASAP7_75t_L g245 ( .A(n_223), .B(n_179), .Y(n_245) );
BUFx3_ASAP7_75t_L g246 ( .A(n_216), .Y(n_246) );
NAND2xp5_ASAP7_75t_L g247 ( .A(n_224), .B(n_179), .Y(n_247) );
INVx1_ASAP7_75t_SL g248 ( .A(n_216), .Y(n_248) );
NAND2xp5_ASAP7_75t_SL g249 ( .A(n_216), .B(n_208), .Y(n_249) );
NAND2xp5_ASAP7_75t_L g250 ( .A(n_225), .B(n_179), .Y(n_250) );
INVx1_ASAP7_75t_L g251 ( .A(n_230), .Y(n_251) );
INVxp67_ASAP7_75t_L g252 ( .A(n_244), .Y(n_252) );
INVx2_ASAP7_75t_L g253 ( .A(n_229), .Y(n_253) );
CKINVDCx14_ASAP7_75t_R g254 ( .A(n_246), .Y(n_254) );
AND2x2_ASAP7_75t_L g255 ( .A(n_234), .B(n_227), .Y(n_255) );
INVx2_ASAP7_75t_L g256 ( .A(n_229), .Y(n_256) );
AND2x2_ASAP7_75t_L g257 ( .A(n_246), .B(n_220), .Y(n_257) );
OAI21xp5_ASAP7_75t_SL g258 ( .A1(n_232), .A2(n_201), .B(n_208), .Y(n_258) );
INVx1_ASAP7_75t_SL g259 ( .A(n_234), .Y(n_259) );
AOI22xp33_ASAP7_75t_SL g260 ( .A1(n_246), .A2(n_211), .B1(n_212), .B2(n_209), .Y(n_260) );
INVx1_ASAP7_75t_L g261 ( .A(n_231), .Y(n_261) );
AND2x2_ASAP7_75t_L g262 ( .A(n_241), .B(n_220), .Y(n_262) );
NAND2x1_ASAP7_75t_L g263 ( .A(n_235), .B(n_199), .Y(n_263) );
INVx1_ASAP7_75t_L g264 ( .A(n_235), .Y(n_264) );
HB1xp67_ASAP7_75t_L g265 ( .A(n_229), .Y(n_265) );
NAND2xp5_ASAP7_75t_L g266 ( .A(n_238), .B(n_218), .Y(n_266) );
AOI22xp5_ASAP7_75t_L g267 ( .A1(n_249), .A2(n_203), .B1(n_189), .B2(n_182), .Y(n_267) );
INVx1_ASAP7_75t_L g268 ( .A(n_238), .Y(n_268) );
NOR2x1_ASAP7_75t_L g269 ( .A(n_239), .B(n_199), .Y(n_269) );
OAI22xp5_ASAP7_75t_L g270 ( .A1(n_232), .A2(n_192), .B1(n_182), .B2(n_211), .Y(n_270) );
NOR2xp33_ASAP7_75t_L g271 ( .A(n_240), .B(n_218), .Y(n_271) );
OAI31xp33_ASAP7_75t_L g272 ( .A1(n_242), .A2(n_180), .A3(n_209), .B(n_212), .Y(n_272) );
AOI31xp33_ASAP7_75t_L g273 ( .A1(n_232), .A2(n_209), .A3(n_211), .B(n_212), .Y(n_273) );
O2A1O1Ixp33_ASAP7_75t_L g274 ( .A1(n_245), .A2(n_190), .B(n_180), .C(n_173), .Y(n_274) );
OAI22xp5_ASAP7_75t_L g275 ( .A1(n_248), .A2(n_212), .B1(n_211), .B2(n_177), .Y(n_275) );
INVx3_ASAP7_75t_L g276 ( .A(n_263), .Y(n_276) );
INVx2_ASAP7_75t_L g277 ( .A(n_265), .Y(n_277) );
INVx1_ASAP7_75t_L g278 ( .A(n_261), .Y(n_278) );
AND2x2_ASAP7_75t_L g279 ( .A(n_262), .B(n_248), .Y(n_279) );
HB1xp67_ASAP7_75t_L g280 ( .A(n_265), .Y(n_280) );
NAND2xp5_ASAP7_75t_L g281 ( .A(n_271), .B(n_236), .Y(n_281) );
INVx1_ASAP7_75t_L g282 ( .A(n_264), .Y(n_282) );
INVxp33_ASAP7_75t_L g283 ( .A(n_269), .Y(n_283) );
INVx2_ASAP7_75t_SL g284 ( .A(n_253), .Y(n_284) );
INVx1_ASAP7_75t_L g285 ( .A(n_268), .Y(n_285) );
AND2x2_ASAP7_75t_SL g286 ( .A(n_254), .B(n_237), .Y(n_286) );
NAND2xp5_ASAP7_75t_SL g287 ( .A(n_274), .B(n_272), .Y(n_287) );
NAND2xp5_ASAP7_75t_L g288 ( .A(n_255), .B(n_247), .Y(n_288) );
NAND2xp5_ASAP7_75t_L g289 ( .A(n_255), .B(n_250), .Y(n_289) );
NAND2xp5_ASAP7_75t_L g290 ( .A(n_266), .B(n_250), .Y(n_290) );
NAND2xp5_ASAP7_75t_L g291 ( .A(n_252), .B(n_237), .Y(n_291) );
OR2x2_ASAP7_75t_L g292 ( .A(n_257), .B(n_233), .Y(n_292) );
INVx1_ASAP7_75t_L g293 ( .A(n_256), .Y(n_293) );
INVx1_ASAP7_75t_L g294 ( .A(n_254), .Y(n_294) );
INVxp67_ASAP7_75t_L g295 ( .A(n_273), .Y(n_295) );
INVx1_ASAP7_75t_L g296 ( .A(n_258), .Y(n_296) );
AND2x2_ASAP7_75t_L g297 ( .A(n_260), .B(n_243), .Y(n_297) );
AOI22xp5_ASAP7_75t_L g298 ( .A1(n_270), .A2(n_228), .B1(n_222), .B2(n_184), .Y(n_298) );
INVx1_ASAP7_75t_L g299 ( .A(n_275), .Y(n_299) );
INVx2_ASAP7_75t_L g300 ( .A(n_267), .Y(n_300) );
INVx1_ASAP7_75t_L g301 ( .A(n_251), .Y(n_301) );
INVx1_ASAP7_75t_SL g302 ( .A(n_259), .Y(n_302) );
OAI22xp33_ASAP7_75t_L g303 ( .A1(n_295), .A2(n_287), .B1(n_298), .B2(n_296), .Y(n_303) );
INVx2_ASAP7_75t_L g304 ( .A(n_284), .Y(n_304) );
AOI31xp33_ASAP7_75t_SL g305 ( .A1(n_300), .A2(n_10), .A3(n_11), .B(n_12), .Y(n_305) );
A2O1A1Ixp33_ASAP7_75t_L g306 ( .A1(n_286), .A2(n_177), .B(n_185), .C(n_166), .Y(n_306) );
AOI211x1_ASAP7_75t_SL g307 ( .A1(n_290), .A2(n_14), .B(n_15), .C(n_16), .Y(n_307) );
XNOR2xp5_ASAP7_75t_L g308 ( .A(n_281), .B(n_17), .Y(n_308) );
NOR3x1_ASAP7_75t_L g309 ( .A(n_299), .B(n_20), .C(n_168), .Y(n_309) );
NOR2x1_ASAP7_75t_L g310 ( .A(n_276), .B(n_204), .Y(n_310) );
O2A1O1Ixp33_ASAP7_75t_L g311 ( .A1(n_280), .A2(n_155), .B(n_161), .C(n_163), .Y(n_311) );
INVx1_ASAP7_75t_SL g312 ( .A(n_302), .Y(n_312) );
OAI22xp33_ASAP7_75t_L g313 ( .A1(n_283), .A2(n_163), .B1(n_159), .B2(n_151), .Y(n_313) );
OAI211xp5_ASAP7_75t_L g314 ( .A1(n_297), .A2(n_170), .B(n_154), .C(n_159), .Y(n_314) );
AOI211xp5_ASAP7_75t_L g315 ( .A1(n_283), .A2(n_154), .B(n_159), .C(n_163), .Y(n_315) );
AOI221xp5_ASAP7_75t_SL g316 ( .A1(n_291), .A2(n_23), .B1(n_24), .B2(n_27), .C(n_28), .Y(n_316) );
INVx1_ASAP7_75t_SL g317 ( .A(n_292), .Y(n_317) );
O2A1O1Ixp5_ASAP7_75t_L g318 ( .A1(n_278), .A2(n_37), .B(n_39), .C(n_41), .Y(n_318) );
OAI22xp5_ASAP7_75t_L g319 ( .A1(n_303), .A2(n_289), .B1(n_288), .B2(n_279), .Y(n_319) );
AOI21xp5_ASAP7_75t_SL g320 ( .A1(n_306), .A2(n_277), .B(n_301), .Y(n_320) );
INVx2_ASAP7_75t_SL g321 ( .A(n_304), .Y(n_321) );
AOI211xp5_ASAP7_75t_L g322 ( .A1(n_305), .A2(n_285), .B(n_282), .C(n_293), .Y(n_322) );
NOR2x1_ASAP7_75t_L g323 ( .A(n_310), .B(n_313), .Y(n_323) );
NAND4xp25_ASAP7_75t_L g324 ( .A(n_309), .B(n_307), .C(n_316), .D(n_314), .Y(n_324) );
NAND3xp33_ASAP7_75t_L g325 ( .A(n_315), .B(n_318), .C(n_311), .Y(n_325) );
AOI21xp33_ASAP7_75t_SL g326 ( .A1(n_303), .A2(n_286), .B(n_308), .Y(n_326) );
AOI22xp5_ASAP7_75t_L g327 ( .A1(n_303), .A2(n_296), .B1(n_287), .B2(n_295), .Y(n_327) );
AOI22x1_ASAP7_75t_L g328 ( .A1(n_308), .A2(n_295), .B1(n_312), .B2(n_294), .Y(n_328) );
OR2x2_ASAP7_75t_L g329 ( .A(n_317), .B(n_302), .Y(n_329) );
HB1xp67_ASAP7_75t_L g330 ( .A(n_329), .Y(n_330) );
CKINVDCx20_ASAP7_75t_R g331 ( .A(n_328), .Y(n_331) );
HB1xp67_ASAP7_75t_L g332 ( .A(n_321), .Y(n_332) );
INVx1_ASAP7_75t_SL g333 ( .A(n_323), .Y(n_333) );
NAND2xp33_ASAP7_75t_R g334 ( .A(n_326), .B(n_322), .Y(n_334) );
CKINVDCx20_ASAP7_75t_R g335 ( .A(n_327), .Y(n_335) );
CKINVDCx5p33_ASAP7_75t_R g336 ( .A(n_319), .Y(n_336) );
INVx2_ASAP7_75t_L g337 ( .A(n_330), .Y(n_337) );
XNOR2x2_ASAP7_75t_L g338 ( .A(n_333), .B(n_324), .Y(n_338) );
OAI22xp5_ASAP7_75t_L g339 ( .A1(n_336), .A2(n_322), .B1(n_325), .B2(n_320), .Y(n_339) );
INVx2_ASAP7_75t_L g340 ( .A(n_332), .Y(n_340) );
INVx1_ASAP7_75t_L g341 ( .A(n_337), .Y(n_341) );
INVx2_ASAP7_75t_SL g342 ( .A(n_340), .Y(n_342) );
XNOR2xp5_ASAP7_75t_L g343 ( .A(n_338), .B(n_331), .Y(n_343) );
INVx1_ASAP7_75t_L g344 ( .A(n_341), .Y(n_344) );
INVx2_ASAP7_75t_L g345 ( .A(n_342), .Y(n_345) );
AOI22xp33_ASAP7_75t_SL g346 ( .A1(n_345), .A2(n_335), .B1(n_339), .B2(n_343), .Y(n_346) );
AOI21xp33_ASAP7_75t_L g347 ( .A1(n_346), .A2(n_344), .B(n_334), .Y(n_347) );
endmodule