module fake_aes_6106_n_537 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_6, n_4, n_40, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_537);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_6;
input n_4;
input n_40;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_537;
wire n_117;
wire n_361;
wire n_513;
wire n_185;
wire n_407;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_154;
wire n_328;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_353;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_532;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_211;
wire n_334;
wire n_389;
wire n_436;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_231;
wire n_452;
wire n_518;
wire n_298;
wire n_411;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_366;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_244;
wire n_119;
wire n_141;
wire n_517;
wire n_479;
wire n_97;
wire n_167;
wire n_447;
wire n_171;
wire n_196;
wire n_192;
wire n_502;
wire n_312;
wire n_455;
wire n_529;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_367;
wire n_250;
wire n_85;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_381;
wire n_304;
wire n_399;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_404;
wire n_369;
wire n_509;
wire n_172;
wire n_329;
wire n_251;
wire n_525;
wire n_218;
wire n_507;
wire n_271;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_133;
wire n_149;
wire n_81;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_107;
wire n_403;
wire n_516;
wire n_254;
wire n_262;
wire n_239;
wire n_439;
wire n_87;
wire n_379;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_370;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_245;
wire n_90;
wire n_357;
wire n_260;
wire n_78;
wire n_201;
wire n_197;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_126;
wire n_178;
wire n_118;
wire n_365;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_376;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_435;
wire n_216;
wire n_147;
wire n_148;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_497;
wire n_339;
wire n_240;
wire n_378;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_335;
wire n_272;
wire n_534;
wire n_531;
wire n_397;
wire n_146;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_198;
wire n_169;
wire n_424;
wire n_156;
wire n_124;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_418;
wire n_493;
wire n_380;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_258;
wire n_253;
wire n_515;
wire n_84;
wire n_266;
wire n_213;
wire n_182;
wire n_492;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_521;
wire n_469;
wire n_123;
wire n_457;
wire n_223;
wire n_494;
wire n_480;
wire n_372;
wire n_453;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_425;
wire n_332;
wire n_414;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_406;
wire n_395;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g78 ( .A(n_28), .Y(n_78) );
INVx1_ASAP7_75t_L g79 ( .A(n_31), .Y(n_79) );
INVx1_ASAP7_75t_L g80 ( .A(n_46), .Y(n_80) );
CKINVDCx5p33_ASAP7_75t_R g81 ( .A(n_4), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_2), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_55), .Y(n_83) );
INVx1_ASAP7_75t_L g84 ( .A(n_37), .Y(n_84) );
INVxp67_ASAP7_75t_SL g85 ( .A(n_5), .Y(n_85) );
INVxp67_ASAP7_75t_SL g86 ( .A(n_5), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_61), .Y(n_87) );
INVxp33_ASAP7_75t_L g88 ( .A(n_67), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_19), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_59), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_54), .Y(n_91) );
BUFx6f_ASAP7_75t_L g92 ( .A(n_33), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_16), .Y(n_93) );
CKINVDCx14_ASAP7_75t_R g94 ( .A(n_13), .Y(n_94) );
CKINVDCx5p33_ASAP7_75t_R g95 ( .A(n_4), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_2), .Y(n_96) );
CKINVDCx5p33_ASAP7_75t_R g97 ( .A(n_65), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_25), .Y(n_98) );
CKINVDCx20_ASAP7_75t_R g99 ( .A(n_11), .Y(n_99) );
CKINVDCx16_ASAP7_75t_R g100 ( .A(n_32), .Y(n_100) );
CKINVDCx20_ASAP7_75t_R g101 ( .A(n_20), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_76), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_52), .Y(n_103) );
CKINVDCx20_ASAP7_75t_R g104 ( .A(n_58), .Y(n_104) );
CKINVDCx5p33_ASAP7_75t_R g105 ( .A(n_68), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_13), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_34), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_38), .Y(n_108) );
INVx2_ASAP7_75t_L g109 ( .A(n_62), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_40), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_75), .Y(n_111) );
CKINVDCx5p33_ASAP7_75t_R g112 ( .A(n_12), .Y(n_112) );
BUFx5_ASAP7_75t_L g113 ( .A(n_71), .Y(n_113) );
INVx2_ASAP7_75t_L g114 ( .A(n_14), .Y(n_114) );
OAI21x1_ASAP7_75t_L g115 ( .A1(n_109), .A2(n_35), .B(n_74), .Y(n_115) );
BUFx6f_ASAP7_75t_L g116 ( .A(n_92), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_114), .Y(n_117) );
HB1xp67_ASAP7_75t_L g118 ( .A(n_94), .Y(n_118) );
BUFx12f_ASAP7_75t_L g119 ( .A(n_97), .Y(n_119) );
OAI21x1_ASAP7_75t_L g120 ( .A1(n_109), .A2(n_30), .B(n_73), .Y(n_120) );
INVx2_ASAP7_75t_L g121 ( .A(n_113), .Y(n_121) );
AND2x2_ASAP7_75t_L g122 ( .A(n_88), .B(n_0), .Y(n_122) );
BUFx6f_ASAP7_75t_L g123 ( .A(n_92), .Y(n_123) );
BUFx6f_ASAP7_75t_L g124 ( .A(n_92), .Y(n_124) );
INVx2_ASAP7_75t_L g125 ( .A(n_113), .Y(n_125) );
HB1xp67_ASAP7_75t_L g126 ( .A(n_81), .Y(n_126) );
INVx1_ASAP7_75t_L g127 ( .A(n_114), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_78), .Y(n_128) );
INVx1_ASAP7_75t_L g129 ( .A(n_79), .Y(n_129) );
NAND2xp5_ASAP7_75t_L g130 ( .A(n_89), .B(n_0), .Y(n_130) );
AND2x2_ASAP7_75t_L g131 ( .A(n_100), .B(n_1), .Y(n_131) );
BUFx6f_ASAP7_75t_L g132 ( .A(n_92), .Y(n_132) );
AND2x2_ASAP7_75t_SL g133 ( .A(n_80), .B(n_36), .Y(n_133) );
INVx2_ASAP7_75t_L g134 ( .A(n_113), .Y(n_134) );
NAND2xp5_ASAP7_75t_SL g135 ( .A(n_113), .B(n_1), .Y(n_135) );
HB1xp67_ASAP7_75t_L g136 ( .A(n_81), .Y(n_136) );
BUFx8_ASAP7_75t_L g137 ( .A(n_113), .Y(n_137) );
INVx2_ASAP7_75t_L g138 ( .A(n_116), .Y(n_138) );
INVx8_ASAP7_75t_L g139 ( .A(n_119), .Y(n_139) );
AND2x4_ASAP7_75t_L g140 ( .A(n_128), .B(n_89), .Y(n_140) );
AND2x6_ASAP7_75t_L g141 ( .A(n_122), .B(n_83), .Y(n_141) );
INVx1_ASAP7_75t_L g142 ( .A(n_121), .Y(n_142) );
NAND2xp5_ASAP7_75t_L g143 ( .A(n_118), .B(n_95), .Y(n_143) );
OAI221xp5_ASAP7_75t_L g144 ( .A1(n_136), .A2(n_96), .B1(n_82), .B2(n_106), .C(n_93), .Y(n_144) );
NOR2xp33_ASAP7_75t_L g145 ( .A(n_118), .B(n_84), .Y(n_145) );
INVx4_ASAP7_75t_SL g146 ( .A(n_116), .Y(n_146) );
INVx3_ASAP7_75t_L g147 ( .A(n_121), .Y(n_147) );
HB1xp67_ASAP7_75t_SL g148 ( .A(n_137), .Y(n_148) );
BUFx6f_ASAP7_75t_L g149 ( .A(n_116), .Y(n_149) );
INVx4_ASAP7_75t_L g150 ( .A(n_133), .Y(n_150) );
INVxp33_ASAP7_75t_L g151 ( .A(n_136), .Y(n_151) );
NAND2xp5_ASAP7_75t_L g152 ( .A(n_128), .B(n_95), .Y(n_152) );
INVx1_ASAP7_75t_L g153 ( .A(n_121), .Y(n_153) );
CKINVDCx5p33_ASAP7_75t_R g154 ( .A(n_119), .Y(n_154) );
INVx4_ASAP7_75t_L g155 ( .A(n_133), .Y(n_155) );
INVx1_ASAP7_75t_L g156 ( .A(n_125), .Y(n_156) );
NAND2xp5_ASAP7_75t_L g157 ( .A(n_129), .B(n_112), .Y(n_157) );
BUFx3_ASAP7_75t_L g158 ( .A(n_137), .Y(n_158) );
INVx1_ASAP7_75t_L g159 ( .A(n_125), .Y(n_159) );
NAND2x1p5_ASAP7_75t_L g160 ( .A(n_133), .B(n_87), .Y(n_160) );
NOR2xp33_ASAP7_75t_L g161 ( .A(n_129), .B(n_90), .Y(n_161) );
INVx1_ASAP7_75t_SL g162 ( .A(n_119), .Y(n_162) );
INVx1_ASAP7_75t_L g163 ( .A(n_142), .Y(n_163) );
NAND2xp5_ASAP7_75t_L g164 ( .A(n_140), .B(n_122), .Y(n_164) );
AND2x2_ASAP7_75t_L g165 ( .A(n_158), .B(n_131), .Y(n_165) );
BUFx3_ASAP7_75t_L g166 ( .A(n_158), .Y(n_166) );
BUFx6f_ASAP7_75t_L g167 ( .A(n_158), .Y(n_167) );
BUFx6f_ASAP7_75t_L g168 ( .A(n_147), .Y(n_168) );
INVx1_ASAP7_75t_L g169 ( .A(n_142), .Y(n_169) );
INVx1_ASAP7_75t_L g170 ( .A(n_153), .Y(n_170) );
INVx3_ASAP7_75t_L g171 ( .A(n_140), .Y(n_171) );
INVx1_ASAP7_75t_L g172 ( .A(n_153), .Y(n_172) );
BUFx3_ASAP7_75t_L g173 ( .A(n_141), .Y(n_173) );
NOR2xp33_ASAP7_75t_SL g174 ( .A(n_150), .B(n_104), .Y(n_174) );
INVx1_ASAP7_75t_L g175 ( .A(n_156), .Y(n_175) );
BUFx2_ASAP7_75t_L g176 ( .A(n_141), .Y(n_176) );
NAND2xp5_ASAP7_75t_L g177 ( .A(n_140), .B(n_122), .Y(n_177) );
INVx1_ASAP7_75t_L g178 ( .A(n_156), .Y(n_178) );
NOR2xp33_ASAP7_75t_L g179 ( .A(n_152), .B(n_126), .Y(n_179) );
NOR2x1p5_ASAP7_75t_L g180 ( .A(n_154), .B(n_131), .Y(n_180) );
NAND2xp5_ASAP7_75t_L g181 ( .A(n_140), .B(n_131), .Y(n_181) );
BUFx3_ASAP7_75t_L g182 ( .A(n_141), .Y(n_182) );
AND2x2_ASAP7_75t_SL g183 ( .A(n_150), .B(n_91), .Y(n_183) );
AND2x4_ASAP7_75t_L g184 ( .A(n_150), .B(n_130), .Y(n_184) );
BUFx4f_ASAP7_75t_L g185 ( .A(n_141), .Y(n_185) );
NOR2xp33_ASAP7_75t_L g186 ( .A(n_157), .B(n_130), .Y(n_186) );
NAND2xp5_ASAP7_75t_SL g187 ( .A(n_150), .B(n_137), .Y(n_187) );
INVx2_ASAP7_75t_L g188 ( .A(n_147), .Y(n_188) );
NOR2xp67_ASAP7_75t_L g189 ( .A(n_155), .B(n_161), .Y(n_189) );
INVx1_ASAP7_75t_L g190 ( .A(n_159), .Y(n_190) );
AND2x4_ASAP7_75t_L g191 ( .A(n_155), .B(n_115), .Y(n_191) );
CKINVDCx5p33_ASAP7_75t_R g192 ( .A(n_139), .Y(n_192) );
BUFx2_ASAP7_75t_L g193 ( .A(n_141), .Y(n_193) );
NAND2xp5_ASAP7_75t_SL g194 ( .A(n_155), .B(n_137), .Y(n_194) );
OAI22xp5_ASAP7_75t_L g195 ( .A1(n_155), .A2(n_160), .B1(n_144), .B2(n_104), .Y(n_195) );
INVx2_ASAP7_75t_L g196 ( .A(n_163), .Y(n_196) );
NOR2xp33_ASAP7_75t_L g197 ( .A(n_181), .B(n_160), .Y(n_197) );
OAI22xp33_ASAP7_75t_L g198 ( .A1(n_174), .A2(n_160), .B1(n_99), .B2(n_101), .Y(n_198) );
INVx4_ASAP7_75t_L g199 ( .A(n_185), .Y(n_199) );
NAND2x1p5_ASAP7_75t_L g200 ( .A(n_173), .B(n_162), .Y(n_200) );
AOI22xp33_ASAP7_75t_L g201 ( .A1(n_183), .A2(n_141), .B1(n_137), .B2(n_135), .Y(n_201) );
NOR2xp33_ASAP7_75t_L g202 ( .A(n_181), .B(n_151), .Y(n_202) );
AND2x4_ASAP7_75t_L g203 ( .A(n_173), .B(n_141), .Y(n_203) );
BUFx2_ASAP7_75t_L g204 ( .A(n_165), .Y(n_204) );
INVx2_ASAP7_75t_SL g205 ( .A(n_180), .Y(n_205) );
AOI21xp5_ASAP7_75t_L g206 ( .A1(n_191), .A2(n_159), .B(n_115), .Y(n_206) );
AND2x4_ASAP7_75t_L g207 ( .A(n_173), .B(n_141), .Y(n_207) );
INVx5_ASAP7_75t_L g208 ( .A(n_167), .Y(n_208) );
NAND2xp5_ASAP7_75t_L g209 ( .A(n_186), .B(n_139), .Y(n_209) );
OR2x6_ASAP7_75t_L g210 ( .A(n_182), .B(n_139), .Y(n_210) );
NAND2x1p5_ASAP7_75t_L g211 ( .A(n_182), .B(n_185), .Y(n_211) );
OR2x6_ASAP7_75t_L g212 ( .A(n_182), .B(n_139), .Y(n_212) );
AOI22xp5_ASAP7_75t_L g213 ( .A1(n_183), .A2(n_139), .B1(n_145), .B2(n_143), .Y(n_213) );
INVx3_ASAP7_75t_L g214 ( .A(n_166), .Y(n_214) );
INVx1_ASAP7_75t_L g215 ( .A(n_171), .Y(n_215) );
INVx3_ASAP7_75t_L g216 ( .A(n_166), .Y(n_216) );
AOI21xp5_ASAP7_75t_L g217 ( .A1(n_191), .A2(n_115), .B(n_120), .Y(n_217) );
BUFx6f_ASAP7_75t_L g218 ( .A(n_166), .Y(n_218) );
INVx2_ASAP7_75t_L g219 ( .A(n_163), .Y(n_219) );
INVx1_ASAP7_75t_L g220 ( .A(n_171), .Y(n_220) );
AOI21xp5_ASAP7_75t_L g221 ( .A1(n_191), .A2(n_194), .B(n_187), .Y(n_221) );
BUFx2_ASAP7_75t_L g222 ( .A(n_165), .Y(n_222) );
AOI21xp5_ASAP7_75t_L g223 ( .A1(n_191), .A2(n_120), .B(n_147), .Y(n_223) );
NAND2xp5_ASAP7_75t_L g224 ( .A(n_186), .B(n_112), .Y(n_224) );
AND2x4_ASAP7_75t_L g225 ( .A(n_184), .B(n_85), .Y(n_225) );
OAI22xp5_ASAP7_75t_L g226 ( .A1(n_183), .A2(n_148), .B1(n_101), .B2(n_99), .Y(n_226) );
NOR2x1_ASAP7_75t_L g227 ( .A(n_180), .B(n_98), .Y(n_227) );
AOI21xp5_ASAP7_75t_L g228 ( .A1(n_164), .A2(n_177), .B(n_189), .Y(n_228) );
OAI22xp5_ASAP7_75t_L g229 ( .A1(n_201), .A2(n_185), .B1(n_184), .B2(n_164), .Y(n_229) );
AOI22xp33_ASAP7_75t_L g230 ( .A1(n_198), .A2(n_195), .B1(n_184), .B2(n_174), .Y(n_230) );
OAI22xp5_ASAP7_75t_L g231 ( .A1(n_201), .A2(n_185), .B1(n_184), .B2(n_177), .Y(n_231) );
BUFx2_ASAP7_75t_L g232 ( .A(n_203), .Y(n_232) );
AND2x4_ASAP7_75t_L g233 ( .A(n_203), .B(n_171), .Y(n_233) );
BUFx4_ASAP7_75t_SL g234 ( .A(n_210), .Y(n_234) );
INVx1_ASAP7_75t_L g235 ( .A(n_225), .Y(n_235) );
O2A1O1Ixp33_ASAP7_75t_L g236 ( .A1(n_198), .A2(n_195), .B(n_179), .C(n_165), .Y(n_236) );
O2A1O1Ixp33_ASAP7_75t_L g237 ( .A1(n_224), .A2(n_179), .B(n_171), .C(n_189), .Y(n_237) );
BUFx2_ASAP7_75t_L g238 ( .A(n_225), .Y(n_238) );
INVx6_ASAP7_75t_L g239 ( .A(n_218), .Y(n_239) );
CKINVDCx6p67_ASAP7_75t_R g240 ( .A(n_210), .Y(n_240) );
INVx4_ASAP7_75t_L g241 ( .A(n_210), .Y(n_241) );
INVx1_ASAP7_75t_L g242 ( .A(n_225), .Y(n_242) );
NOR2x1_ASAP7_75t_SL g243 ( .A(n_212), .B(n_167), .Y(n_243) );
CKINVDCx11_ASAP7_75t_R g244 ( .A(n_212), .Y(n_244) );
AND3x4_ASAP7_75t_L g245 ( .A(n_227), .B(n_203), .C(n_207), .Y(n_245) );
OAI221xp5_ASAP7_75t_L g246 ( .A1(n_202), .A2(n_176), .B1(n_193), .B2(n_86), .C(n_192), .Y(n_246) );
AOI22xp33_ASAP7_75t_L g247 ( .A1(n_204), .A2(n_193), .B1(n_176), .B2(n_175), .Y(n_247) );
AOI22xp33_ASAP7_75t_SL g248 ( .A1(n_226), .A2(n_105), .B1(n_97), .B2(n_178), .Y(n_248) );
AOI22xp33_ASAP7_75t_SL g249 ( .A1(n_222), .A2(n_105), .B1(n_190), .B2(n_178), .Y(n_249) );
AOI22xp33_ASAP7_75t_L g250 ( .A1(n_202), .A2(n_190), .B1(n_169), .B2(n_175), .Y(n_250) );
INVx2_ASAP7_75t_SL g251 ( .A(n_212), .Y(n_251) );
AOI22xp33_ASAP7_75t_L g252 ( .A1(n_197), .A2(n_172), .B1(n_170), .B2(n_169), .Y(n_252) );
NAND2xp33_ASAP7_75t_L g253 ( .A(n_209), .B(n_167), .Y(n_253) );
INVx1_ASAP7_75t_L g254 ( .A(n_196), .Y(n_254) );
AOI22xp5_ASAP7_75t_L g255 ( .A1(n_197), .A2(n_172), .B1(n_170), .B2(n_188), .Y(n_255) );
AOI221xp5_ASAP7_75t_L g256 ( .A1(n_236), .A2(n_205), .B1(n_228), .B2(n_213), .C(n_117), .Y(n_256) );
AOI221xp5_ASAP7_75t_L g257 ( .A1(n_230), .A2(n_117), .B1(n_127), .B2(n_96), .C(n_219), .Y(n_257) );
AOI22xp33_ASAP7_75t_L g258 ( .A1(n_229), .A2(n_207), .B1(n_196), .B2(n_219), .Y(n_258) );
O2A1O1Ixp5_ASAP7_75t_L g259 ( .A1(n_241), .A2(n_221), .B(n_217), .C(n_223), .Y(n_259) );
AOI22xp33_ASAP7_75t_L g260 ( .A1(n_231), .A2(n_207), .B1(n_220), .B2(n_215), .Y(n_260) );
OAI22xp5_ASAP7_75t_L g261 ( .A1(n_252), .A2(n_200), .B1(n_206), .B2(n_211), .Y(n_261) );
AND2x2_ASAP7_75t_L g262 ( .A(n_254), .B(n_200), .Y(n_262) );
OAI22xp5_ASAP7_75t_L g263 ( .A1(n_255), .A2(n_211), .B1(n_218), .B2(n_199), .Y(n_263) );
BUFx8_ASAP7_75t_SL g264 ( .A(n_238), .Y(n_264) );
INVx1_ASAP7_75t_L g265 ( .A(n_235), .Y(n_265) );
INVx1_ASAP7_75t_L g266 ( .A(n_242), .Y(n_266) );
INVxp67_ASAP7_75t_L g267 ( .A(n_249), .Y(n_267) );
BUFx4f_ASAP7_75t_SL g268 ( .A(n_240), .Y(n_268) );
AOI21xp33_ASAP7_75t_L g269 ( .A1(n_237), .A2(n_216), .B(n_214), .Y(n_269) );
AOI22xp33_ASAP7_75t_L g270 ( .A1(n_244), .A2(n_199), .B1(n_216), .B2(n_214), .Y(n_270) );
AOI322xp5_ASAP7_75t_L g271 ( .A1(n_248), .A2(n_127), .A3(n_102), .B1(n_111), .B2(n_110), .C1(n_108), .C2(n_107), .Y(n_271) );
AO31x2_ASAP7_75t_L g272 ( .A1(n_243), .A2(n_125), .A3(n_134), .B(n_103), .Y(n_272) );
INVx1_ASAP7_75t_L g273 ( .A(n_233), .Y(n_273) );
INVx3_ASAP7_75t_L g274 ( .A(n_239), .Y(n_274) );
OAI221xp5_ASAP7_75t_L g275 ( .A1(n_250), .A2(n_199), .B1(n_188), .B2(n_218), .C(n_134), .Y(n_275) );
CKINVDCx5p33_ASAP7_75t_R g276 ( .A(n_234), .Y(n_276) );
OAI22xp33_ASAP7_75t_L g277 ( .A1(n_240), .A2(n_241), .B1(n_246), .B2(n_251), .Y(n_277) );
AND2x4_ASAP7_75t_L g278 ( .A(n_273), .B(n_241), .Y(n_278) );
AND2x2_ASAP7_75t_L g279 ( .A(n_262), .B(n_232), .Y(n_279) );
INVx1_ASAP7_75t_L g280 ( .A(n_265), .Y(n_280) );
INVx1_ASAP7_75t_L g281 ( .A(n_265), .Y(n_281) );
AOI22xp33_ASAP7_75t_SL g282 ( .A1(n_268), .A2(n_251), .B1(n_232), .B2(n_244), .Y(n_282) );
INVx2_ASAP7_75t_SL g283 ( .A(n_276), .Y(n_283) );
NAND4xp25_ASAP7_75t_SL g284 ( .A(n_271), .B(n_245), .C(n_247), .D(n_7), .Y(n_284) );
HB1xp67_ASAP7_75t_L g285 ( .A(n_262), .Y(n_285) );
AOI22xp33_ASAP7_75t_L g286 ( .A1(n_267), .A2(n_245), .B1(n_233), .B2(n_253), .Y(n_286) );
INVx1_ASAP7_75t_L g287 ( .A(n_266), .Y(n_287) );
OR2x2_ASAP7_75t_L g288 ( .A(n_266), .B(n_233), .Y(n_288) );
INVx2_ASAP7_75t_L g289 ( .A(n_259), .Y(n_289) );
INVx1_ASAP7_75t_L g290 ( .A(n_272), .Y(n_290) );
AOI222xp33_ASAP7_75t_L g291 ( .A1(n_276), .A2(n_253), .B1(n_134), .B2(n_92), .C1(n_120), .C2(n_188), .Y(n_291) );
HB1xp67_ASAP7_75t_L g292 ( .A(n_264), .Y(n_292) );
OAI211xp5_ASAP7_75t_L g293 ( .A1(n_271), .A2(n_116), .B(n_123), .C(n_124), .Y(n_293) );
OAI321xp33_ASAP7_75t_L g294 ( .A1(n_277), .A2(n_132), .A3(n_116), .B1(n_123), .B2(n_124), .C(n_168), .Y(n_294) );
NAND3xp33_ASAP7_75t_SL g295 ( .A(n_256), .B(n_138), .C(n_6), .Y(n_295) );
AND2x4_ASAP7_75t_L g296 ( .A(n_273), .B(n_208), .Y(n_296) );
AOI22xp5_ASAP7_75t_L g297 ( .A1(n_258), .A2(n_239), .B1(n_218), .B2(n_113), .Y(n_297) );
OR2x2_ASAP7_75t_L g298 ( .A(n_272), .B(n_3), .Y(n_298) );
AND2x2_ASAP7_75t_L g299 ( .A(n_272), .B(n_239), .Y(n_299) );
AND2x2_ASAP7_75t_L g300 ( .A(n_280), .B(n_272), .Y(n_300) );
NAND3xp33_ASAP7_75t_L g301 ( .A(n_298), .B(n_257), .C(n_269), .Y(n_301) );
AOI22xp5_ASAP7_75t_L g302 ( .A1(n_284), .A2(n_260), .B1(n_270), .B2(n_261), .Y(n_302) );
INVx3_ASAP7_75t_L g303 ( .A(n_299), .Y(n_303) );
AND2x4_ASAP7_75t_L g304 ( .A(n_299), .B(n_272), .Y(n_304) );
OAI31xp33_ASAP7_75t_L g305 ( .A1(n_293), .A2(n_261), .A3(n_275), .B(n_263), .Y(n_305) );
INVx1_ASAP7_75t_L g306 ( .A(n_280), .Y(n_306) );
AND2x2_ASAP7_75t_L g307 ( .A(n_281), .B(n_113), .Y(n_307) );
OR2x2_ASAP7_75t_L g308 ( .A(n_285), .B(n_274), .Y(n_308) );
NAND2xp33_ASAP7_75t_SL g309 ( .A(n_298), .B(n_274), .Y(n_309) );
NAND3xp33_ASAP7_75t_SL g310 ( .A(n_282), .B(n_3), .C(n_6), .Y(n_310) );
NOR2xp67_ASAP7_75t_L g311 ( .A(n_290), .B(n_274), .Y(n_311) );
AND2x2_ASAP7_75t_L g312 ( .A(n_281), .B(n_113), .Y(n_312) );
AND2x2_ASAP7_75t_L g313 ( .A(n_287), .B(n_7), .Y(n_313) );
INVx1_ASAP7_75t_L g314 ( .A(n_287), .Y(n_314) );
NAND2xp5_ASAP7_75t_L g315 ( .A(n_279), .B(n_239), .Y(n_315) );
NAND2xp5_ASAP7_75t_L g316 ( .A(n_279), .B(n_8), .Y(n_316) );
AOI21xp33_ASAP7_75t_L g317 ( .A1(n_289), .A2(n_291), .B(n_290), .Y(n_317) );
NOR3xp33_ASAP7_75t_L g318 ( .A(n_295), .B(n_138), .C(n_147), .Y(n_318) );
INVx1_ASAP7_75t_L g319 ( .A(n_289), .Y(n_319) );
NAND2xp5_ASAP7_75t_L g320 ( .A(n_288), .B(n_8), .Y(n_320) );
INVx1_ASAP7_75t_L g321 ( .A(n_289), .Y(n_321) );
O2A1O1Ixp5_ASAP7_75t_L g322 ( .A1(n_278), .A2(n_138), .B(n_208), .C(n_48), .Y(n_322) );
INVx1_ASAP7_75t_L g323 ( .A(n_288), .Y(n_323) );
INVx1_ASAP7_75t_L g324 ( .A(n_278), .Y(n_324) );
INVx1_ASAP7_75t_L g325 ( .A(n_278), .Y(n_325) );
INVx2_ASAP7_75t_L g326 ( .A(n_278), .Y(n_326) );
INVx1_ASAP7_75t_L g327 ( .A(n_296), .Y(n_327) );
HB1xp67_ASAP7_75t_L g328 ( .A(n_296), .Y(n_328) );
OAI33xp33_ASAP7_75t_L g329 ( .A1(n_283), .A2(n_9), .A3(n_10), .B1(n_11), .B2(n_12), .B3(n_14), .Y(n_329) );
AND2x2_ASAP7_75t_L g330 ( .A(n_303), .B(n_296), .Y(n_330) );
OR2x2_ASAP7_75t_L g331 ( .A(n_303), .B(n_286), .Y(n_331) );
BUFx2_ASAP7_75t_L g332 ( .A(n_309), .Y(n_332) );
AND2x4_ASAP7_75t_L g333 ( .A(n_303), .B(n_296), .Y(n_333) );
INVx2_ASAP7_75t_L g334 ( .A(n_319), .Y(n_334) );
INVx1_ASAP7_75t_L g335 ( .A(n_306), .Y(n_335) );
A2O1A1Ixp33_ASAP7_75t_L g336 ( .A1(n_310), .A2(n_294), .B(n_283), .C(n_292), .Y(n_336) );
OR2x2_ASAP7_75t_L g337 ( .A(n_323), .B(n_297), .Y(n_337) );
INVx2_ASAP7_75t_L g338 ( .A(n_319), .Y(n_338) );
AND2x2_ASAP7_75t_L g339 ( .A(n_321), .B(n_132), .Y(n_339) );
INVx1_ASAP7_75t_L g340 ( .A(n_306), .Y(n_340) );
OR2x2_ASAP7_75t_L g341 ( .A(n_323), .B(n_297), .Y(n_341) );
AND2x2_ASAP7_75t_L g342 ( .A(n_304), .B(n_116), .Y(n_342) );
INVx1_ASAP7_75t_L g343 ( .A(n_314), .Y(n_343) );
INVx3_ASAP7_75t_L g344 ( .A(n_304), .Y(n_344) );
NAND2xp5_ASAP7_75t_L g345 ( .A(n_314), .B(n_9), .Y(n_345) );
BUFx2_ASAP7_75t_L g346 ( .A(n_304), .Y(n_346) );
AND2x2_ASAP7_75t_L g347 ( .A(n_300), .B(n_116), .Y(n_347) );
INVx1_ASAP7_75t_L g348 ( .A(n_321), .Y(n_348) );
NAND2xp5_ASAP7_75t_L g349 ( .A(n_300), .B(n_10), .Y(n_349) );
AND2x2_ASAP7_75t_L g350 ( .A(n_324), .B(n_123), .Y(n_350) );
INVx2_ASAP7_75t_L g351 ( .A(n_307), .Y(n_351) );
INVx2_ASAP7_75t_L g352 ( .A(n_307), .Y(n_352) );
AND2x2_ASAP7_75t_L g353 ( .A(n_324), .B(n_123), .Y(n_353) );
INVx2_ASAP7_75t_SL g354 ( .A(n_328), .Y(n_354) );
INVx3_ASAP7_75t_L g355 ( .A(n_326), .Y(n_355) );
INVx1_ASAP7_75t_L g356 ( .A(n_325), .Y(n_356) );
INVx2_ASAP7_75t_L g357 ( .A(n_312), .Y(n_357) );
INVx1_ASAP7_75t_SL g358 ( .A(n_308), .Y(n_358) );
AND2x4_ASAP7_75t_L g359 ( .A(n_326), .B(n_123), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_325), .Y(n_360) );
NAND2xp5_ASAP7_75t_L g361 ( .A(n_312), .B(n_15), .Y(n_361) );
INVx1_ASAP7_75t_L g362 ( .A(n_327), .Y(n_362) );
INVx1_ASAP7_75t_L g363 ( .A(n_327), .Y(n_363) );
AND2x2_ASAP7_75t_L g364 ( .A(n_317), .B(n_123), .Y(n_364) );
OR2x2_ASAP7_75t_L g365 ( .A(n_308), .B(n_15), .Y(n_365) );
INVx1_ASAP7_75t_L g366 ( .A(n_311), .Y(n_366) );
NAND2xp5_ASAP7_75t_L g367 ( .A(n_313), .B(n_16), .Y(n_367) );
INVxp67_ASAP7_75t_SL g368 ( .A(n_311), .Y(n_368) );
AND2x4_ASAP7_75t_L g369 ( .A(n_313), .B(n_123), .Y(n_369) );
NAND3xp33_ASAP7_75t_SL g370 ( .A(n_305), .B(n_17), .C(n_18), .Y(n_370) );
AND2x2_ASAP7_75t_L g371 ( .A(n_315), .B(n_132), .Y(n_371) );
AND2x2_ASAP7_75t_L g372 ( .A(n_302), .B(n_132), .Y(n_372) );
NOR2x1_ASAP7_75t_L g373 ( .A(n_301), .B(n_124), .Y(n_373) );
INVx1_ASAP7_75t_L g374 ( .A(n_335), .Y(n_374) );
INVx1_ASAP7_75t_L g375 ( .A(n_335), .Y(n_375) );
OR2x2_ASAP7_75t_L g376 ( .A(n_358), .B(n_316), .Y(n_376) );
OR2x2_ASAP7_75t_L g377 ( .A(n_358), .B(n_320), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_340), .Y(n_378) );
NAND2xp5_ASAP7_75t_L g379 ( .A(n_349), .B(n_17), .Y(n_379) );
INVx1_ASAP7_75t_L g380 ( .A(n_340), .Y(n_380) );
AND2x2_ASAP7_75t_L g381 ( .A(n_330), .B(n_18), .Y(n_381) );
AOI21xp5_ASAP7_75t_L g382 ( .A1(n_373), .A2(n_322), .B(n_329), .Y(n_382) );
AND2x2_ASAP7_75t_L g383 ( .A(n_344), .B(n_132), .Y(n_383) );
INVx1_ASAP7_75t_SL g384 ( .A(n_365), .Y(n_384) );
AND2x2_ASAP7_75t_L g385 ( .A(n_344), .B(n_132), .Y(n_385) );
AND2x2_ASAP7_75t_L g386 ( .A(n_344), .B(n_132), .Y(n_386) );
AND2x2_ASAP7_75t_L g387 ( .A(n_344), .B(n_124), .Y(n_387) );
AOI22xp5_ASAP7_75t_L g388 ( .A1(n_370), .A2(n_318), .B1(n_208), .B2(n_124), .Y(n_388) );
NAND2xp5_ASAP7_75t_L g389 ( .A(n_349), .B(n_19), .Y(n_389) );
INVx1_ASAP7_75t_L g390 ( .A(n_343), .Y(n_390) );
AND4x1_ASAP7_75t_L g391 ( .A(n_336), .B(n_20), .C(n_21), .D(n_22), .Y(n_391) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_362), .B(n_21), .Y(n_392) );
OR2x2_ASAP7_75t_L g393 ( .A(n_346), .B(n_124), .Y(n_393) );
AND2x2_ASAP7_75t_L g394 ( .A(n_330), .B(n_124), .Y(n_394) );
OAI321xp33_ASAP7_75t_L g395 ( .A1(n_370), .A2(n_149), .A3(n_24), .B1(n_26), .B2(n_27), .C(n_29), .Y(n_395) );
NAND2xp33_ASAP7_75t_L g396 ( .A(n_373), .B(n_208), .Y(n_396) );
NAND2xp33_ASAP7_75t_SL g397 ( .A(n_332), .B(n_167), .Y(n_397) );
OR2x2_ASAP7_75t_L g398 ( .A(n_346), .B(n_23), .Y(n_398) );
O2A1O1Ixp33_ASAP7_75t_L g399 ( .A1(n_367), .A2(n_345), .B(n_365), .C(n_372), .Y(n_399) );
NOR2x1_ASAP7_75t_L g400 ( .A(n_332), .B(n_39), .Y(n_400) );
AND2x2_ASAP7_75t_L g401 ( .A(n_333), .B(n_41), .Y(n_401) );
AOI211x1_ASAP7_75t_L g402 ( .A1(n_367), .A2(n_42), .B(n_43), .C(n_44), .Y(n_402) );
INVx1_ASAP7_75t_L g403 ( .A(n_343), .Y(n_403) );
XNOR2x2_ASAP7_75t_L g404 ( .A(n_331), .B(n_45), .Y(n_404) );
NAND2xp5_ASAP7_75t_L g405 ( .A(n_362), .B(n_47), .Y(n_405) );
AND2x2_ASAP7_75t_L g406 ( .A(n_347), .B(n_49), .Y(n_406) );
INVx1_ASAP7_75t_L g407 ( .A(n_363), .Y(n_407) );
A2O1A1Ixp33_ASAP7_75t_L g408 ( .A1(n_368), .A2(n_50), .B(n_51), .C(n_53), .Y(n_408) );
AND2x2_ASAP7_75t_L g409 ( .A(n_333), .B(n_56), .Y(n_409) );
NAND2x1p5_ASAP7_75t_L g410 ( .A(n_369), .B(n_167), .Y(n_410) );
OAI31xp33_ASAP7_75t_L g411 ( .A1(n_372), .A2(n_57), .A3(n_60), .B(n_63), .Y(n_411) );
OR2x2_ASAP7_75t_L g412 ( .A(n_354), .B(n_64), .Y(n_412) );
OR2x2_ASAP7_75t_L g413 ( .A(n_354), .B(n_66), .Y(n_413) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_363), .B(n_69), .Y(n_414) );
NAND2xp5_ASAP7_75t_L g415 ( .A(n_356), .B(n_70), .Y(n_415) );
AND2x4_ASAP7_75t_L g416 ( .A(n_366), .B(n_72), .Y(n_416) );
NAND2xp5_ASAP7_75t_L g417 ( .A(n_356), .B(n_77), .Y(n_417) );
INVx2_ASAP7_75t_L g418 ( .A(n_334), .Y(n_418) );
NAND3xp33_ASAP7_75t_L g419 ( .A(n_372), .B(n_149), .C(n_168), .Y(n_419) );
NOR2x1_ASAP7_75t_L g420 ( .A(n_345), .B(n_168), .Y(n_420) );
NAND2xp5_ASAP7_75t_L g421 ( .A(n_360), .B(n_168), .Y(n_421) );
AND2x4_ASAP7_75t_L g422 ( .A(n_366), .B(n_149), .Y(n_422) );
AOI22xp33_ASAP7_75t_L g423 ( .A1(n_331), .A2(n_168), .B1(n_149), .B2(n_167), .Y(n_423) );
AND2x2_ASAP7_75t_L g424 ( .A(n_333), .B(n_168), .Y(n_424) );
INVx1_ASAP7_75t_L g425 ( .A(n_374), .Y(n_425) );
NAND2xp5_ASAP7_75t_L g426 ( .A(n_384), .B(n_347), .Y(n_426) );
INVx1_ASAP7_75t_L g427 ( .A(n_375), .Y(n_427) );
AND2x2_ASAP7_75t_L g428 ( .A(n_394), .B(n_333), .Y(n_428) );
XOR2xp5_ASAP7_75t_L g429 ( .A(n_376), .B(n_337), .Y(n_429) );
NAND2xp5_ASAP7_75t_L g430 ( .A(n_407), .B(n_360), .Y(n_430) );
XNOR2x1_ASAP7_75t_L g431 ( .A(n_381), .B(n_361), .Y(n_431) );
AOI22xp5_ASAP7_75t_L g432 ( .A1(n_379), .A2(n_342), .B1(n_364), .B2(n_354), .Y(n_432) );
NAND2xp5_ASAP7_75t_L g433 ( .A(n_378), .B(n_342), .Y(n_433) );
XNOR2xp5_ASAP7_75t_L g434 ( .A(n_391), .B(n_371), .Y(n_434) );
CKINVDCx20_ASAP7_75t_R g435 ( .A(n_377), .Y(n_435) );
INVx1_ASAP7_75t_L g436 ( .A(n_380), .Y(n_436) );
AND2x2_ASAP7_75t_L g437 ( .A(n_424), .B(n_351), .Y(n_437) );
OAI221xp5_ASAP7_75t_L g438 ( .A1(n_399), .A2(n_368), .B1(n_361), .B2(n_364), .C(n_337), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_390), .Y(n_439) );
AOI22xp5_ASAP7_75t_L g440 ( .A1(n_389), .A2(n_364), .B1(n_371), .B2(n_369), .Y(n_440) );
NAND2x1_ASAP7_75t_L g441 ( .A(n_400), .B(n_338), .Y(n_441) );
NAND3xp33_ASAP7_75t_L g442 ( .A(n_402), .B(n_353), .C(n_369), .Y(n_442) );
NAND2xp5_ASAP7_75t_L g443 ( .A(n_403), .B(n_351), .Y(n_443) );
XNOR2xp5_ASAP7_75t_L g444 ( .A(n_401), .B(n_369), .Y(n_444) );
AOI21xp5_ASAP7_75t_L g445 ( .A1(n_396), .A2(n_339), .B(n_348), .Y(n_445) );
NAND2xp5_ASAP7_75t_L g446 ( .A(n_418), .B(n_351), .Y(n_446) );
NAND3xp33_ASAP7_75t_SL g447 ( .A(n_408), .B(n_388), .C(n_411), .Y(n_447) );
NOR2xp33_ASAP7_75t_R g448 ( .A(n_397), .B(n_341), .Y(n_448) );
INVx2_ASAP7_75t_SL g449 ( .A(n_393), .Y(n_449) );
INVx3_ASAP7_75t_L g450 ( .A(n_383), .Y(n_450) );
NOR2xp33_ASAP7_75t_L g451 ( .A(n_392), .B(n_355), .Y(n_451) );
INVx1_ASAP7_75t_L g452 ( .A(n_421), .Y(n_452) );
INVx1_ASAP7_75t_L g453 ( .A(n_383), .Y(n_453) );
AND2x2_ASAP7_75t_L g454 ( .A(n_385), .B(n_352), .Y(n_454) );
INVx1_ASAP7_75t_L g455 ( .A(n_385), .Y(n_455) );
NAND2xp5_ASAP7_75t_L g456 ( .A(n_386), .B(n_357), .Y(n_456) );
NAND2xp33_ASAP7_75t_L g457 ( .A(n_398), .B(n_357), .Y(n_457) );
XNOR2xp5_ASAP7_75t_L g458 ( .A(n_409), .B(n_357), .Y(n_458) );
INVx1_ASAP7_75t_L g459 ( .A(n_386), .Y(n_459) );
INVx1_ASAP7_75t_L g460 ( .A(n_387), .Y(n_460) );
NOR2xp33_ASAP7_75t_L g461 ( .A(n_416), .B(n_355), .Y(n_461) );
HB1xp67_ASAP7_75t_L g462 ( .A(n_387), .Y(n_462) );
AND2x2_ASAP7_75t_L g463 ( .A(n_406), .B(n_352), .Y(n_463) );
AND2x2_ASAP7_75t_L g464 ( .A(n_406), .B(n_352), .Y(n_464) );
INVx1_ASAP7_75t_SL g465 ( .A(n_412), .Y(n_465) );
INVx1_ASAP7_75t_L g466 ( .A(n_420), .Y(n_466) );
NOR2x1_ASAP7_75t_SL g467 ( .A(n_413), .B(n_348), .Y(n_467) );
O2A1O1Ixp33_ASAP7_75t_L g468 ( .A1(n_408), .A2(n_353), .B(n_350), .C(n_341), .Y(n_468) );
INVx1_ASAP7_75t_L g469 ( .A(n_422), .Y(n_469) );
INVx1_ASAP7_75t_L g470 ( .A(n_422), .Y(n_470) );
OAI22xp5_ASAP7_75t_L g471 ( .A1(n_419), .A2(n_355), .B1(n_338), .B2(n_334), .Y(n_471) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_416), .B(n_353), .Y(n_472) );
AOI221x1_ASAP7_75t_SL g473 ( .A1(n_416), .A2(n_338), .B1(n_359), .B2(n_355), .C(n_339), .Y(n_473) );
NOR2xp33_ASAP7_75t_L g474 ( .A(n_405), .B(n_350), .Y(n_474) );
INVx1_ASAP7_75t_SL g475 ( .A(n_397), .Y(n_475) );
NOR2xp33_ASAP7_75t_L g476 ( .A(n_414), .B(n_339), .Y(n_476) );
INVx1_ASAP7_75t_L g477 ( .A(n_422), .Y(n_477) );
NAND2xp5_ASAP7_75t_SL g478 ( .A(n_382), .B(n_359), .Y(n_478) );
INVx2_ASAP7_75t_SL g479 ( .A(n_410), .Y(n_479) );
INVx3_ASAP7_75t_L g480 ( .A(n_404), .Y(n_480) );
NOR3xp33_ASAP7_75t_L g481 ( .A(n_395), .B(n_359), .C(n_149), .Y(n_481) );
INVx2_ASAP7_75t_L g482 ( .A(n_410), .Y(n_482) );
HB1xp67_ASAP7_75t_L g483 ( .A(n_415), .Y(n_483) );
NAND2xp5_ASAP7_75t_SL g484 ( .A(n_404), .B(n_359), .Y(n_484) );
INVx3_ASAP7_75t_L g485 ( .A(n_396), .Y(n_485) );
INVx1_ASAP7_75t_L g486 ( .A(n_417), .Y(n_486) );
INVx2_ASAP7_75t_L g487 ( .A(n_423), .Y(n_487) );
OAI321xp33_ASAP7_75t_L g488 ( .A1(n_423), .A2(n_146), .A3(n_149), .B1(n_167), .B2(n_168), .C(n_370), .Y(n_488) );
INVxp67_ASAP7_75t_SL g489 ( .A(n_393), .Y(n_489) );
HB1xp67_ASAP7_75t_L g490 ( .A(n_393), .Y(n_490) );
INVx1_ASAP7_75t_L g491 ( .A(n_407), .Y(n_491) );
INVx1_ASAP7_75t_L g492 ( .A(n_407), .Y(n_492) );
NAND2xp5_ASAP7_75t_L g493 ( .A(n_384), .B(n_146), .Y(n_493) );
XNOR2x1_ASAP7_75t_L g494 ( .A(n_384), .B(n_146), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g495 ( .A(n_384), .B(n_146), .Y(n_495) );
AOI21xp33_ASAP7_75t_L g496 ( .A1(n_480), .A2(n_486), .B(n_483), .Y(n_496) );
AND2x2_ASAP7_75t_L g497 ( .A(n_428), .B(n_462), .Y(n_497) );
XOR2x2_ASAP7_75t_L g498 ( .A(n_431), .B(n_429), .Y(n_498) );
AOI21xp5_ASAP7_75t_L g499 ( .A1(n_484), .A2(n_480), .B(n_494), .Y(n_499) );
NAND4xp25_ASAP7_75t_L g500 ( .A(n_480), .B(n_473), .C(n_447), .D(n_438), .Y(n_500) );
OAI32xp33_ASAP7_75t_L g501 ( .A1(n_475), .A2(n_435), .A3(n_485), .B1(n_462), .B2(n_442), .Y(n_501) );
AOI22xp5_ASAP7_75t_L g502 ( .A1(n_435), .A2(n_451), .B1(n_469), .B2(n_477), .Y(n_502) );
O2A1O1Ixp5_ASAP7_75t_L g503 ( .A1(n_478), .A2(n_485), .B(n_451), .C(n_489), .Y(n_503) );
NOR3xp33_ASAP7_75t_L g504 ( .A(n_488), .B(n_481), .C(n_486), .Y(n_504) );
A2O1A1Ixp33_ASAP7_75t_L g505 ( .A1(n_473), .A2(n_468), .B(n_485), .C(n_475), .Y(n_505) );
AOI21xp33_ASAP7_75t_L g506 ( .A1(n_466), .A2(n_434), .B(n_487), .Y(n_506) );
NAND2x1p5_ASAP7_75t_L g507 ( .A(n_494), .B(n_479), .Y(n_507) );
OAI22x1_ASAP7_75t_L g508 ( .A1(n_458), .A2(n_444), .B1(n_479), .B2(n_432), .Y(n_508) );
OAI32xp33_ASAP7_75t_L g509 ( .A1(n_450), .A2(n_465), .A3(n_490), .B1(n_477), .B2(n_470), .Y(n_509) );
AOI221xp5_ASAP7_75t_L g510 ( .A1(n_470), .A2(n_469), .B1(n_427), .B2(n_439), .C(n_425), .Y(n_510) );
INVx1_ASAP7_75t_L g511 ( .A(n_491), .Y(n_511) );
AOI22xp5_ASAP7_75t_L g512 ( .A1(n_431), .A2(n_440), .B1(n_457), .B2(n_449), .Y(n_512) );
O2A1O1Ixp33_ASAP7_75t_L g513 ( .A1(n_457), .A2(n_487), .B(n_441), .C(n_471), .Y(n_513) );
O2A1O1Ixp33_ASAP7_75t_L g514 ( .A1(n_500), .A2(n_495), .B(n_493), .C(n_426), .Y(n_514) );
NAND2xp5_ASAP7_75t_L g515 ( .A(n_510), .B(n_436), .Y(n_515) );
NAND4xp25_ASAP7_75t_L g516 ( .A(n_499), .B(n_461), .C(n_474), .D(n_476), .Y(n_516) );
AOI22xp33_ASAP7_75t_L g517 ( .A1(n_508), .A2(n_450), .B1(n_453), .B2(n_460), .Y(n_517) );
AO22x2_ASAP7_75t_L g518 ( .A1(n_498), .A2(n_449), .B1(n_491), .B2(n_492), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_512), .B(n_492), .Y(n_519) );
NOR3xp33_ASAP7_75t_L g520 ( .A(n_501), .B(n_450), .C(n_452), .Y(n_520) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_512), .B(n_437), .Y(n_521) );
NOR2x1_ASAP7_75t_L g522 ( .A(n_505), .B(n_482), .Y(n_522) );
AOI21xp5_ASAP7_75t_L g523 ( .A1(n_503), .A2(n_467), .B(n_445), .Y(n_523) );
OAI221xp5_ASAP7_75t_L g524 ( .A1(n_517), .A2(n_496), .B1(n_506), .B2(n_513), .C(n_507), .Y(n_524) );
AOI22xp33_ASAP7_75t_L g525 ( .A1(n_518), .A2(n_504), .B1(n_455), .B2(n_459), .Y(n_525) );
NAND4xp75_ASAP7_75t_L g526 ( .A(n_522), .B(n_502), .C(n_497), .D(n_461), .Y(n_526) );
OAI21xp33_ASAP7_75t_L g527 ( .A1(n_520), .A2(n_509), .B(n_511), .Y(n_527) );
NAND4xp25_ASAP7_75t_L g528 ( .A(n_523), .B(n_472), .C(n_482), .D(n_433), .Y(n_528) );
OAI22x1_ASAP7_75t_L g529 ( .A1(n_526), .A2(n_519), .B1(n_521), .B2(n_515), .Y(n_529) );
INVx2_ASAP7_75t_L g530 ( .A(n_524), .Y(n_530) );
AOI322xp5_ASAP7_75t_L g531 ( .A1(n_525), .A2(n_527), .A3(n_528), .B1(n_516), .B2(n_464), .C1(n_463), .C2(n_454), .Y(n_531) );
XNOR2xp5_ASAP7_75t_L g532 ( .A(n_530), .B(n_514), .Y(n_532) );
AND3x4_ASAP7_75t_L g533 ( .A(n_529), .B(n_448), .C(n_467), .Y(n_533) );
OR2x2_ASAP7_75t_L g534 ( .A(n_532), .B(n_430), .Y(n_534) );
INVx2_ASAP7_75t_L g535 ( .A(n_534), .Y(n_535) );
OAI22xp33_ASAP7_75t_L g536 ( .A1(n_535), .A2(n_533), .B1(n_531), .B2(n_443), .Y(n_536) );
AOI21xp5_ASAP7_75t_L g537 ( .A1(n_536), .A2(n_446), .B(n_456), .Y(n_537) );
endmodule