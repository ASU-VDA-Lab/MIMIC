module real_jpeg_7699_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_277, n_276, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_277;
input n_276;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_249;
wire n_166;
wire n_176;
wire n_221;
wire n_215;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_271;
wire n_163;
wire n_22;
wire n_237;
wire n_174;
wire n_87;
wire n_255;
wire n_173;
wire n_40;
wire n_105;
wire n_197;
wire n_243;
wire n_115;
wire n_98;
wire n_27;
wire n_184;
wire n_56;
wire n_48;
wire n_200;
wire n_164;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_13;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_238;
wire n_67;
wire n_79;
wire n_178;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_211;
wire n_172;
wire n_45;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_262;
wire n_148;
wire n_222;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_137;
wire n_31;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_203;
wire n_192;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_110;
wire n_61;
wire n_195;
wire n_205;
wire n_258;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_204;
wire n_158;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_225;
wire n_259;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_240;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_97;
wire n_75;
wire n_187;
wire n_34;
wire n_230;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_202;
wire n_179;
wire n_216;
wire n_213;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_210;
wire n_127;
wire n_206;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_181;
wire n_85;
wire n_101;
wire n_256;
wire n_182;
wire n_269;
wire n_96;
wire n_253;
wire n_273;
wire n_89;
wire n_16;

BUFx24_ASAP7_75t_L g86 ( 
.A(n_0),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g172 ( 
.A1(n_1),
.A2(n_25),
.B1(n_26),
.B2(n_173),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_1),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_SL g211 ( 
.A1(n_1),
.A2(n_40),
.B1(n_42),
.B2(n_173),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_L g252 ( 
.A1(n_1),
.A2(n_86),
.B1(n_87),
.B2(n_173),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_2),
.A2(n_86),
.B1(n_87),
.B2(n_114),
.Y(n_113)
);

INVx2_ASAP7_75t_SL g114 ( 
.A(n_2),
.Y(n_114)
);

AOI21xp33_ASAP7_75t_L g142 ( 
.A1(n_2),
.A2(n_9),
.B(n_86),
.Y(n_142)
);

BUFx10_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_L g44 ( 
.A1(n_5),
.A2(n_25),
.B1(n_26),
.B2(n_45),
.Y(n_44)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_5),
.Y(n_45)
);

A2O1A1Ixp33_ASAP7_75t_L g48 ( 
.A1(n_5),
.A2(n_40),
.B(n_44),
.C(n_49),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_5),
.B(n_40),
.Y(n_49)
);

AOI21xp5_ASAP7_75t_L g52 ( 
.A1(n_5),
.A2(n_9),
.B(n_26),
.Y(n_52)
);

BUFx6f_ASAP7_75t_SL g73 ( 
.A(n_6),
.Y(n_73)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_7),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_SL g24 ( 
.A1(n_8),
.A2(n_25),
.B1(n_26),
.B2(n_29),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_8),
.Y(n_29)
);

AOI22xp33_ASAP7_75t_SL g39 ( 
.A1(n_8),
.A2(n_29),
.B1(n_40),
.B2(n_42),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_8),
.A2(n_29),
.B1(n_86),
.B2(n_87),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_8),
.A2(n_11),
.B1(n_29),
.B2(n_133),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g34 ( 
.A1(n_9),
.A2(n_25),
.B1(n_26),
.B2(n_35),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_9),
.Y(n_35)
);

AOI22xp5_ASAP7_75t_SL g47 ( 
.A1(n_9),
.A2(n_35),
.B1(n_40),
.B2(n_42),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_9),
.B(n_71),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_9),
.A2(n_35),
.B1(n_86),
.B2(n_87),
.Y(n_89)
);

O2A1O1Ixp33_ASAP7_75t_L g94 ( 
.A1(n_9),
.A2(n_73),
.B(n_87),
.C(n_95),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_9),
.B(n_112),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_9),
.A2(n_11),
.B1(n_35),
.B2(n_133),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_10),
.A2(n_25),
.B1(n_26),
.B2(n_155),
.Y(n_154)
);

CKINVDCx16_ASAP7_75t_R g155 ( 
.A(n_10),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_SL g200 ( 
.A1(n_10),
.A2(n_40),
.B1(n_42),
.B2(n_155),
.Y(n_200)
);

OAI22xp33_ASAP7_75t_SL g237 ( 
.A1(n_10),
.A2(n_86),
.B1(n_87),
.B2(n_155),
.Y(n_237)
);

AOI22xp33_ASAP7_75t_SL g269 ( 
.A1(n_10),
.A2(n_11),
.B1(n_133),
.B2(n_155),
.Y(n_269)
);

INVx2_ASAP7_75t_SL g133 ( 
.A(n_11),
.Y(n_133)
);

A2O1A1Ixp33_ASAP7_75t_L g136 ( 
.A1(n_11),
.A2(n_113),
.B(n_114),
.C(n_137),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_11),
.B(n_114),
.Y(n_137)
);

A2O1A1Ixp33_ASAP7_75t_L g141 ( 
.A1(n_11),
.A2(n_35),
.B(n_114),
.C(n_142),
.Y(n_141)
);

XOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_262),
.Y(n_12)
);

OAI321xp33_ASAP7_75t_L g13 ( 
.A1(n_14),
.A2(n_230),
.A3(n_255),
.B1(n_260),
.B2(n_261),
.C(n_276),
.Y(n_13)
);

AOI321xp33_ASAP7_75t_L g14 ( 
.A1(n_15),
.A2(n_184),
.A3(n_204),
.B1(n_224),
.B2(n_229),
.C(n_277),
.Y(n_14)
);

NOR3xp33_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_147),
.C(n_181),
.Y(n_15)
);

AOI21xp5_ASAP7_75t_L g16 ( 
.A1(n_17),
.A2(n_120),
.B(n_146),
.Y(n_16)
);

OAI21xp5_ASAP7_75t_SL g17 ( 
.A1(n_18),
.A2(n_101),
.B(n_119),
.Y(n_17)
);

AOI21xp5_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_79),
.B(n_100),
.Y(n_18)
);

OAI21xp5_ASAP7_75t_SL g19 ( 
.A1(n_20),
.A2(n_64),
.B(n_78),
.Y(n_19)
);

AOI21xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_54),
.B(n_63),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_36),
.Y(n_21)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_22),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_SL g63 ( 
.A(n_22),
.B(n_36),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_22),
.A2(n_56),
.B1(n_110),
.B2(n_111),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_22),
.B(n_105),
.C(n_111),
.Y(n_143)
);

AOI21xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_30),
.B(n_31),
.Y(n_22)
);

CKINVDCx16_ASAP7_75t_R g23 ( 
.A(n_24),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_24),
.A2(n_32),
.B1(n_33),
.B2(n_34),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g57 ( 
.A(n_25),
.B(n_58),
.Y(n_57)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_26),
.B(n_33),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

BUFx24_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_30),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_30),
.B(n_98),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_30),
.A2(n_98),
.B1(n_154),
.B2(n_171),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_31),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_32),
.B(n_34),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_32),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_33),
.B(n_35),
.Y(n_58)
);

OAI21xp5_ASAP7_75t_SL g152 ( 
.A1(n_33),
.A2(n_153),
.B(n_156),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_34),
.B(n_97),
.Y(n_96)
);

A2O1A1Ixp33_ASAP7_75t_L g51 ( 
.A1(n_35),
.A2(n_42),
.B(n_45),
.C(n_52),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g60 ( 
.A(n_35),
.B(n_44),
.Y(n_60)
);

OAI21xp33_ASAP7_75t_SL g95 ( 
.A1(n_35),
.A2(n_40),
.B(n_74),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_SL g36 ( 
.A1(n_37),
.A2(n_50),
.B1(n_51),
.B2(n_53),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_37),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g65 ( 
.A(n_37),
.B(n_51),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_37),
.A2(n_53),
.B1(n_84),
.B2(n_92),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_37),
.B(n_84),
.C(n_99),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_37),
.A2(n_53),
.B1(n_151),
.B2(n_152),
.Y(n_150)
);

AOI21xp5_ASAP7_75t_L g37 ( 
.A1(n_38),
.A2(n_43),
.B(n_46),
.Y(n_37)
);

INVxp67_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_39),
.A2(n_44),
.B1(n_47),
.B2(n_48),
.Y(n_76)
);

INVx11_ASAP7_75t_L g42 ( 
.A(n_40),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_40),
.A2(n_42),
.B1(n_73),
.B2(n_74),
.Y(n_72)
);

INVx13_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVxp67_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_44),
.B(n_48),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_L g199 ( 
.A1(n_44),
.A2(n_200),
.B(n_201),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_44),
.A2(n_48),
.B1(n_200),
.B2(n_211),
.Y(n_210)
);

INVxp67_ASAP7_75t_L g201 ( 
.A(n_46),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_47),
.B(n_48),
.Y(n_46)
);

CKINVDCx14_ASAP7_75t_R g127 ( 
.A(n_47),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_51),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_53),
.B(n_152),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_L g54 ( 
.A1(n_55),
.A2(n_59),
.B(n_62),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_56),
.B(n_57),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_60),
.B(n_61),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_60),
.B(n_61),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_61),
.A2(n_67),
.B1(n_68),
.B2(n_77),
.Y(n_66)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_61),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_61),
.B(n_69),
.C(n_76),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_61),
.A2(n_77),
.B1(n_140),
.B2(n_141),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_61),
.B(n_140),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_65),
.B(n_66),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_65),
.B(n_66),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_68),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_69),
.A2(n_70),
.B1(n_75),
.B2(n_76),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_70),
.Y(n_69)
);

AOI21xp5_ASAP7_75t_L g84 ( 
.A1(n_71),
.A2(n_85),
.B(n_88),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_71),
.A2(n_85),
.B1(n_106),
.B2(n_107),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_71),
.B(n_106),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_71),
.A2(n_106),
.B1(n_237),
.B2(n_252),
.Y(n_251)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

A2O1A1Ixp33_ASAP7_75t_L g90 ( 
.A1(n_72),
.A2(n_73),
.B(n_87),
.C(n_91),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_L g235 ( 
.A1(n_72),
.A2(n_236),
.B(n_238),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_73),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_73),
.B(n_87),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_75),
.A2(n_76),
.B1(n_117),
.B2(n_118),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_75),
.A2(n_76),
.B1(n_169),
.B2(n_170),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_75),
.B(n_170),
.Y(n_191)
);

CKINVDCx16_ASAP7_75t_R g75 ( 
.A(n_76),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_76),
.B(n_104),
.C(n_118),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_80),
.B(n_81),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_80),
.B(n_81),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_82),
.A2(n_83),
.B1(n_93),
.B2(n_99),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_83),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_84),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_84),
.A2(n_92),
.B1(n_126),
.B2(n_129),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_84),
.B(n_126),
.C(n_131),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_84),
.A2(n_92),
.B1(n_160),
.B2(n_161),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_84),
.B(n_160),
.C(n_194),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_86),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g238 ( 
.A(n_88),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_90),
.Y(n_88)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_89),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g178 ( 
.A(n_89),
.B(n_179),
.Y(n_178)
);

CKINVDCx16_ASAP7_75t_R g106 ( 
.A(n_90),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_93),
.Y(n_99)
);

XOR2xp5_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_96),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_94),
.B(n_96),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_97),
.B(n_172),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_103),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_102),
.B(n_103),
.Y(n_119)
);

XOR2xp5_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_116),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_105),
.A2(n_108),
.B1(n_109),
.B2(n_115),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_105),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_105),
.A2(n_115),
.B1(n_160),
.B2(n_161),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_105),
.B(n_160),
.C(n_163),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_109),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_111),
.Y(n_110)
);

AOI21xp5_ASAP7_75t_L g131 ( 
.A1(n_112),
.A2(n_132),
.B(n_134),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_113),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_113),
.A2(n_135),
.B1(n_136),
.B2(n_162),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_113),
.B(n_136),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_L g268 ( 
.A1(n_113),
.A2(n_269),
.B(n_270),
.Y(n_268)
);

AOI21xp5_ASAP7_75t_L g209 ( 
.A1(n_115),
.A2(n_210),
.B(n_212),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_115),
.B(n_210),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_117),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_122),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g146 ( 
.A(n_121),
.B(n_122),
.Y(n_146)
);

XOR2xp5_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_138),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_123),
.B(n_139),
.C(n_145),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_124),
.A2(n_125),
.B1(n_130),
.B2(n_131),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_125),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_126),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_128),
.Y(n_126)
);

INVxp33_ASAP7_75t_L g241 ( 
.A(n_128),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_130),
.A2(n_131),
.B1(n_177),
.B2(n_178),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_130),
.A2(n_131),
.B1(n_233),
.B2(n_234),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_130),
.A2(n_131),
.B1(n_247),
.B2(n_253),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_130),
.B(n_239),
.C(n_242),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_130),
.B(n_253),
.C(n_254),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_131),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_131),
.B(n_175),
.C(n_177),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_132),
.Y(n_162)
);

INVxp67_ASAP7_75t_L g270 ( 
.A(n_134),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_136),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_135),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_139),
.A2(n_143),
.B1(n_144),
.B2(n_145),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_139),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_141),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_143),
.Y(n_145)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

AOI21xp33_ASAP7_75t_L g225 ( 
.A1(n_148),
.A2(n_226),
.B(n_227),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_164),
.Y(n_148)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_149),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_SL g227 ( 
.A(n_149),
.B(n_164),
.Y(n_227)
);

FAx1_ASAP7_75t_SL g149 ( 
.A(n_150),
.B(n_157),
.CI(n_158),
.CON(n_149),
.SN(n_149)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_152),
.Y(n_151)
);

CKINVDCx14_ASAP7_75t_R g153 ( 
.A(n_154),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_SL g158 ( 
.A(n_159),
.B(n_163),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_160),
.A2(n_161),
.B1(n_248),
.B2(n_249),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_160),
.B(n_240),
.C(n_251),
.Y(n_271)
);

CKINVDCx16_ASAP7_75t_R g160 ( 
.A(n_161),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_165),
.A2(n_166),
.B1(n_167),
.B2(n_180),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_165),
.Y(n_180)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_174),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_168),
.B(n_174),
.C(n_180),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_170),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_176),
.Y(n_174)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_179),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_183),
.Y(n_181)
);

AND2x2_ASAP7_75t_L g226 ( 
.A(n_182),
.B(n_183),
.Y(n_226)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_SL g224 ( 
.A1(n_185),
.A2(n_225),
.B(n_228),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_187),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_186),
.B(n_187),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_188),
.B(n_203),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_189),
.A2(n_190),
.B1(n_195),
.B2(n_196),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_189),
.B(n_196),
.C(n_203),
.Y(n_205)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_191),
.A2(n_192),
.B1(n_193),
.B2(n_194),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_191),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_193),
.Y(n_192)
);

CKINVDCx16_ASAP7_75t_R g195 ( 
.A(n_196),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_197),
.A2(n_198),
.B1(n_199),
.B2(n_202),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_197),
.A2(n_198),
.B1(n_216),
.B2(n_219),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_198),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_198),
.B(n_199),
.Y(n_214)
);

AOI21xp5_ASAP7_75t_L g244 ( 
.A1(n_198),
.A2(n_214),
.B(n_216),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_199),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_206),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_205),
.B(n_206),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_207),
.A2(n_208),
.B1(n_222),
.B2(n_223),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_209),
.A2(n_213),
.B1(n_220),
.B2(n_221),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_209),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_209),
.B(n_221),
.C(n_223),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_SL g240 ( 
.A(n_211),
.B(n_241),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_212),
.B(n_232),
.C(n_243),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_212),
.B(n_232),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_213),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_SL g213 ( 
.A(n_214),
.B(n_215),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_216),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_218),
.Y(n_216)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_222),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_245),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_231),
.B(n_245),
.Y(n_261)
);

CKINVDCx16_ASAP7_75t_R g233 ( 
.A(n_234),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_235),
.A2(n_239),
.B1(n_240),
.B2(n_242),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_235),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_237),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g249 ( 
.A1(n_239),
.A2(n_240),
.B1(n_250),
.B2(n_251),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_240),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_243),
.A2(n_244),
.B1(n_258),
.B2(n_259),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_244),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_254),
.Y(n_245)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_247),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_249),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_251),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_252),
.B(n_267),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_257),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_256),
.B(n_257),
.Y(n_260)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_258),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_263),
.B(n_273),
.Y(n_262)
);

INVxp67_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_272),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_265),
.B(n_272),
.Y(n_273)
);

BUFx24_ASAP7_75t_SL g274 ( 
.A(n_265),
.Y(n_274)
);

FAx1_ASAP7_75t_SL g265 ( 
.A(n_266),
.B(n_268),
.CI(n_271),
.CON(n_265),
.SN(n_265)
);


endmodule