module fake_jpeg_11533_n_580 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_580);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_580;

wire n_529;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_442;
wire n_299;
wire n_300;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_570;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_419;
wire n_378;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_260;
wire n_199;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx11_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

INVx2_ASAP7_75t_SL g20 ( 
.A(n_9),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

BUFx10_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_11),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_7),
.Y(n_28)
);

INVxp67_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

INVx6_ASAP7_75t_SL g31 ( 
.A(n_9),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

INVx5_ASAP7_75t_L g35 ( 
.A(n_1),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_11),
.Y(n_36)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_0),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_11),
.Y(n_38)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_15),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_17),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_16),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_16),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_15),
.Y(n_43)
);

OR2x2_ASAP7_75t_L g44 ( 
.A(n_16),
.B(n_6),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_0),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_2),
.Y(n_46)
);

BUFx10_ASAP7_75t_L g47 ( 
.A(n_14),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_7),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_1),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_9),
.Y(n_50)
);

BUFx5_ASAP7_75t_L g51 ( 
.A(n_5),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_7),
.Y(n_52)
);

INVxp67_ASAP7_75t_L g53 ( 
.A(n_7),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_14),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_6),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_8),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_15),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_2),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_8),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_1),
.Y(n_60)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_42),
.Y(n_61)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_61),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_20),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_62),
.A2(n_71),
.B1(n_50),
.B2(n_45),
.Y(n_198)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_22),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_63),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_22),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_64),
.Y(n_128)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_60),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_65),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_44),
.B(n_17),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_66),
.B(n_85),
.Y(n_136)
);

BUFx2_ASAP7_75t_L g67 ( 
.A(n_39),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g127 ( 
.A(n_67),
.Y(n_127)
);

BUFx12f_ASAP7_75t_L g68 ( 
.A(n_39),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g145 ( 
.A(n_68),
.Y(n_145)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_21),
.Y(n_69)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_69),
.Y(n_141)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_21),
.Y(n_70)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_70),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_L g71 ( 
.A1(n_40),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_22),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_72),
.Y(n_165)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_36),
.Y(n_73)
);

INVx3_ASAP7_75t_L g154 ( 
.A(n_73),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_41),
.B(n_17),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_74),
.B(n_83),
.Y(n_177)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_40),
.Y(n_75)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_75),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_43),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g174 ( 
.A(n_76),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_23),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_77),
.B(n_96),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_43),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g181 ( 
.A(n_78),
.Y(n_181)
);

INVx5_ASAP7_75t_L g79 ( 
.A(n_31),
.Y(n_79)
);

BUFx2_ASAP7_75t_L g142 ( 
.A(n_79),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_43),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g196 ( 
.A(n_80),
.Y(n_196)
);

BUFx12f_ASAP7_75t_L g81 ( 
.A(n_39),
.Y(n_81)
);

BUFx3_ASAP7_75t_L g199 ( 
.A(n_81),
.Y(n_199)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_42),
.Y(n_82)
);

INVx3_ASAP7_75t_L g159 ( 
.A(n_82),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_41),
.B(n_44),
.Y(n_83)
);

BUFx5_ASAP7_75t_L g84 ( 
.A(n_31),
.Y(n_84)
);

BUFx12f_ASAP7_75t_L g140 ( 
.A(n_84),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_44),
.B(n_14),
.Y(n_85)
);

INVx8_ASAP7_75t_L g86 ( 
.A(n_26),
.Y(n_86)
);

BUFx2_ASAP7_75t_L g148 ( 
.A(n_86),
.Y(n_148)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_36),
.Y(n_87)
);

INVx3_ASAP7_75t_L g187 ( 
.A(n_87),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_24),
.B(n_3),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_88),
.B(n_104),
.Y(n_162)
);

INVx8_ASAP7_75t_L g89 ( 
.A(n_26),
.Y(n_89)
);

INVx5_ASAP7_75t_L g164 ( 
.A(n_89),
.Y(n_164)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_27),
.Y(n_90)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_90),
.Y(n_147)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_27),
.Y(n_91)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_91),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_49),
.Y(n_92)
);

INVx6_ASAP7_75t_L g156 ( 
.A(n_92),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_42),
.B(n_3),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g193 ( 
.A(n_93),
.B(n_113),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_49),
.Y(n_94)
);

INVx6_ASAP7_75t_L g184 ( 
.A(n_94),
.Y(n_184)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_19),
.Y(n_95)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_95),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_23),
.Y(n_96)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_36),
.Y(n_97)
);

HB1xp67_ASAP7_75t_L g167 ( 
.A(n_97),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_23),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_98),
.B(n_107),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_49),
.Y(n_99)
);

BUFx3_ASAP7_75t_L g205 ( 
.A(n_99),
.Y(n_205)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_19),
.Y(n_100)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_100),
.Y(n_195)
);

BUFx5_ASAP7_75t_L g101 ( 
.A(n_33),
.Y(n_101)
);

INVx4_ASAP7_75t_L g157 ( 
.A(n_101),
.Y(n_157)
);

BUFx12f_ASAP7_75t_L g102 ( 
.A(n_33),
.Y(n_102)
);

INVx5_ASAP7_75t_L g178 ( 
.A(n_102),
.Y(n_178)
);

BUFx10_ASAP7_75t_L g103 ( 
.A(n_23),
.Y(n_103)
);

INVx2_ASAP7_75t_SL g168 ( 
.A(n_103),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_24),
.B(n_3),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_57),
.Y(n_105)
);

INVx4_ASAP7_75t_L g203 ( 
.A(n_105),
.Y(n_203)
);

BUFx5_ASAP7_75t_L g106 ( 
.A(n_37),
.Y(n_106)
);

INVx4_ASAP7_75t_L g158 ( 
.A(n_106),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_23),
.Y(n_107)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_36),
.Y(n_108)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_108),
.Y(n_151)
);

CKINVDCx16_ASAP7_75t_R g109 ( 
.A(n_47),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_109),
.B(n_116),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_57),
.Y(n_110)
);

INVx4_ASAP7_75t_L g161 ( 
.A(n_110),
.Y(n_161)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_25),
.Y(n_111)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_111),
.Y(n_200)
);

BUFx24_ASAP7_75t_L g112 ( 
.A(n_47),
.Y(n_112)
);

INVx13_ASAP7_75t_L g152 ( 
.A(n_112),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_28),
.B(n_4),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_28),
.B(n_13),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_114),
.B(n_125),
.Y(n_169)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_36),
.Y(n_115)
);

INVx4_ASAP7_75t_L g170 ( 
.A(n_115),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_47),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_57),
.Y(n_117)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_117),
.Y(n_153)
);

INVx8_ASAP7_75t_L g118 ( 
.A(n_37),
.Y(n_118)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_118),
.Y(n_166)
);

BUFx3_ASAP7_75t_L g119 ( 
.A(n_51),
.Y(n_119)
);

HB1xp67_ASAP7_75t_L g172 ( 
.A(n_119),
.Y(n_172)
);

INVx8_ASAP7_75t_L g120 ( 
.A(n_51),
.Y(n_120)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_120),
.Y(n_173)
);

BUFx16f_ASAP7_75t_L g121 ( 
.A(n_38),
.Y(n_121)
);

BUFx12_ASAP7_75t_L g160 ( 
.A(n_121),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_60),
.Y(n_122)
);

HB1xp67_ASAP7_75t_L g189 ( 
.A(n_122),
.Y(n_189)
);

BUFx5_ASAP7_75t_L g123 ( 
.A(n_47),
.Y(n_123)
);

BUFx10_ASAP7_75t_L g135 ( 
.A(n_123),
.Y(n_135)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_38),
.Y(n_124)
);

CKINVDCx16_ASAP7_75t_R g129 ( 
.A(n_124),
.Y(n_129)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_38),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_L g130 ( 
.A1(n_65),
.A2(n_20),
.B1(n_60),
.B2(n_47),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g251 ( 
.A1(n_130),
.A2(n_131),
.B1(n_132),
.B2(n_139),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_71),
.A2(n_59),
.B1(n_56),
.B2(n_55),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_86),
.A2(n_20),
.B1(n_29),
.B2(n_53),
.Y(n_132)
);

AOI21xp33_ASAP7_75t_SL g133 ( 
.A1(n_112),
.A2(n_18),
.B(n_38),
.Y(n_133)
);

AOI32xp33_ASAP7_75t_L g212 ( 
.A1(n_133),
.A2(n_103),
.A3(n_62),
.B1(n_115),
.B2(n_13),
.Y(n_212)
);

OA22x2_ASAP7_75t_L g138 ( 
.A1(n_112),
.A2(n_80),
.B1(n_122),
.B2(n_94),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_138),
.B(n_103),
.C(n_117),
.Y(n_213)
);

AOI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_89),
.A2(n_35),
.B1(n_18),
.B2(n_38),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_L g144 ( 
.A1(n_63),
.A2(n_34),
.B1(n_58),
.B2(n_48),
.Y(n_144)
);

OAI22xp33_ASAP7_75t_SL g248 ( 
.A1(n_144),
.A2(n_183),
.B1(n_190),
.B2(n_204),
.Y(n_248)
);

OAI22xp33_ASAP7_75t_SL g163 ( 
.A1(n_64),
.A2(n_18),
.B1(n_58),
.B2(n_48),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_163),
.A2(n_171),
.B1(n_198),
.B2(n_201),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_72),
.A2(n_78),
.B1(n_76),
.B2(n_99),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_SL g176 ( 
.A1(n_118),
.A2(n_35),
.B1(n_46),
.B2(n_34),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_SL g211 ( 
.A1(n_176),
.A2(n_180),
.B1(n_186),
.B2(n_197),
.Y(n_211)
);

AOI22xp33_ASAP7_75t_SL g180 ( 
.A1(n_120),
.A2(n_35),
.B1(n_46),
.B2(n_32),
.Y(n_180)
);

AND2x2_ASAP7_75t_SL g182 ( 
.A(n_79),
.B(n_4),
.Y(n_182)
);

AND2x2_ASAP7_75t_L g237 ( 
.A(n_182),
.B(n_140),
.Y(n_237)
);

AOI22xp33_ASAP7_75t_L g183 ( 
.A1(n_92),
.A2(n_30),
.B1(n_32),
.B2(n_25),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_121),
.B(n_59),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_185),
.B(n_188),
.Y(n_258)
);

AOI22xp33_ASAP7_75t_SL g186 ( 
.A1(n_67),
.A2(n_119),
.B1(n_102),
.B2(n_81),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_68),
.B(n_56),
.Y(n_188)
);

AOI22xp33_ASAP7_75t_L g190 ( 
.A1(n_105),
.A2(n_30),
.B1(n_55),
.B2(n_52),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_73),
.B(n_52),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_191),
.B(n_192),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_68),
.B(n_54),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_97),
.B(n_54),
.Y(n_194)
);

OR2x2_ASAP7_75t_L g225 ( 
.A(n_194),
.B(n_193),
.Y(n_225)
);

AOI22xp33_ASAP7_75t_SL g197 ( 
.A1(n_102),
.A2(n_50),
.B1(n_45),
.B2(n_6),
.Y(n_197)
);

AOI22xp33_ASAP7_75t_SL g201 ( 
.A1(n_81),
.A2(n_4),
.B1(n_5),
.B2(n_9),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_87),
.B(n_124),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_202),
.B(n_13),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_110),
.A2(n_5),
.B1(n_10),
.B2(n_12),
.Y(n_204)
);

INVx3_ASAP7_75t_L g206 ( 
.A(n_127),
.Y(n_206)
);

BUFx2_ASAP7_75t_L g278 ( 
.A(n_206),
.Y(n_278)
);

INVx6_ASAP7_75t_SL g207 ( 
.A(n_160),
.Y(n_207)
);

INVx4_ASAP7_75t_SL g332 ( 
.A(n_207),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_169),
.B(n_12),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_208),
.B(n_215),
.Y(n_301)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_134),
.Y(n_209)
);

INVx1_ASAP7_75t_SL g280 ( 
.A(n_209),
.Y(n_280)
);

O2A1O1Ixp33_ASAP7_75t_L g210 ( 
.A1(n_182),
.A2(n_138),
.B(n_163),
.C(n_179),
.Y(n_210)
);

AND2x2_ASAP7_75t_L g282 ( 
.A(n_210),
.B(n_237),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_L g298 ( 
.A1(n_212),
.A2(n_158),
.B1(n_174),
.B2(n_181),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_213),
.A2(n_266),
.B1(n_261),
.B2(n_228),
.Y(n_314)
);

CKINVDCx14_ASAP7_75t_R g289 ( 
.A(n_214),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_162),
.B(n_13),
.Y(n_215)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_153),
.Y(n_216)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_216),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_137),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_217),
.B(n_220),
.Y(n_283)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_175),
.Y(n_218)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_218),
.Y(n_287)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_195),
.Y(n_219)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_219),
.Y(n_297)
);

CKINVDCx14_ASAP7_75t_R g220 ( 
.A(n_135),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_200),
.B(n_155),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_221),
.B(n_234),
.Y(n_326)
);

INVx3_ASAP7_75t_L g222 ( 
.A(n_127),
.Y(n_222)
);

INVx4_ASAP7_75t_L g317 ( 
.A(n_222),
.Y(n_317)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_142),
.Y(n_223)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_223),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_225),
.B(n_235),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_167),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_226),
.B(n_231),
.Y(n_291)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_142),
.Y(n_227)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_227),
.Y(n_305)
);

HAxp5_ASAP7_75t_SL g228 ( 
.A(n_172),
.B(n_152),
.CON(n_228),
.SN(n_228)
);

OR2x2_ASAP7_75t_L g323 ( 
.A(n_228),
.B(n_261),
.Y(n_323)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_141),
.Y(n_229)
);

INVx2_ASAP7_75t_L g310 ( 
.A(n_229),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_136),
.B(n_149),
.C(n_147),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_230),
.B(n_275),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_160),
.Y(n_231)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_143),
.Y(n_232)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_232),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_151),
.B(n_190),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_177),
.B(n_146),
.Y(n_235)
);

CKINVDCx16_ASAP7_75t_R g236 ( 
.A(n_135),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g284 ( 
.A(n_236),
.B(n_238),
.Y(n_284)
);

CKINVDCx16_ASAP7_75t_R g238 ( 
.A(n_135),
.Y(n_238)
);

INVx3_ASAP7_75t_L g239 ( 
.A(n_170),
.Y(n_239)
);

INVx4_ASAP7_75t_L g319 ( 
.A(n_239),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_160),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_240),
.B(n_245),
.Y(n_303)
);

INVx8_ASAP7_75t_L g241 ( 
.A(n_126),
.Y(n_241)
);

INVx5_ASAP7_75t_L g295 ( 
.A(n_241),
.Y(n_295)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_187),
.Y(n_242)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_242),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_144),
.B(n_183),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_243),
.B(n_244),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_189),
.B(n_138),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_129),
.Y(n_245)
);

INVx3_ASAP7_75t_L g246 ( 
.A(n_164),
.Y(n_246)
);

INVx3_ASAP7_75t_L g318 ( 
.A(n_246),
.Y(n_318)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_203),
.Y(n_247)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_247),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_130),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_249),
.B(n_270),
.Y(n_307)
);

INVx2_ASAP7_75t_SL g250 ( 
.A(n_154),
.Y(n_250)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_250),
.Y(n_333)
);

BUFx12f_ASAP7_75t_L g252 ( 
.A(n_145),
.Y(n_252)
);

BUFx3_ASAP7_75t_L g300 ( 
.A(n_252),
.Y(n_300)
);

BUFx2_ASAP7_75t_L g253 ( 
.A(n_178),
.Y(n_253)
);

INVxp67_ASAP7_75t_L g321 ( 
.A(n_253),
.Y(n_321)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_159),
.Y(n_254)
);

INVxp67_ASAP7_75t_L g330 ( 
.A(n_254),
.Y(n_330)
);

INVx1_ASAP7_75t_SL g255 ( 
.A(n_145),
.Y(n_255)
);

AND2x2_ASAP7_75t_L g292 ( 
.A(n_255),
.B(n_265),
.Y(n_292)
);

CKINVDCx16_ASAP7_75t_R g256 ( 
.A(n_132),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g286 ( 
.A(n_256),
.B(n_263),
.Y(n_286)
);

INVx5_ASAP7_75t_L g257 ( 
.A(n_140),
.Y(n_257)
);

BUFx24_ASAP7_75t_L g315 ( 
.A(n_257),
.Y(n_315)
);

BUFx3_ASAP7_75t_L g259 ( 
.A(n_140),
.Y(n_259)
);

INVx13_ASAP7_75t_L g277 ( 
.A(n_259),
.Y(n_277)
);

BUFx2_ASAP7_75t_L g260 ( 
.A(n_203),
.Y(n_260)
);

CKINVDCx16_ASAP7_75t_R g285 ( 
.A(n_260),
.Y(n_285)
);

BUFx10_ASAP7_75t_L g261 ( 
.A(n_152),
.Y(n_261)
);

AOI22xp33_ASAP7_75t_SL g304 ( 
.A1(n_261),
.A2(n_262),
.B1(n_181),
.B2(n_196),
.Y(n_304)
);

INVx11_ASAP7_75t_L g262 ( 
.A(n_148),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_166),
.B(n_173),
.Y(n_263)
);

A2O1A1Ixp33_ASAP7_75t_L g264 ( 
.A1(n_197),
.A2(n_201),
.B(n_180),
.C(n_176),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_SL g290 ( 
.A(n_264),
.B(n_269),
.Y(n_290)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_150),
.Y(n_265)
);

OAI22xp33_ASAP7_75t_SL g266 ( 
.A1(n_139),
.A2(n_161),
.B1(n_186),
.B2(n_150),
.Y(n_266)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_156),
.Y(n_267)
);

AND2x2_ASAP7_75t_L g293 ( 
.A(n_267),
.B(n_268),
.Y(n_293)
);

INVx3_ASAP7_75t_L g268 ( 
.A(n_205),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_148),
.B(n_199),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_199),
.B(n_168),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_168),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_271),
.B(n_272),
.Y(n_311)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_205),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_156),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_273),
.B(n_274),
.Y(n_316)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_184),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_184),
.B(n_126),
.Y(n_275)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_128),
.Y(n_276)
);

AND2x2_ASAP7_75t_L g294 ( 
.A(n_276),
.B(n_165),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_233),
.A2(n_128),
.B1(n_165),
.B2(n_174),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g344 ( 
.A1(n_281),
.A2(n_329),
.B1(n_247),
.B2(n_250),
.Y(n_344)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_294),
.Y(n_334)
);

AND2x2_ASAP7_75t_L g296 ( 
.A(n_237),
.B(n_157),
.Y(n_296)
);

CKINVDCx14_ASAP7_75t_R g343 ( 
.A(n_296),
.Y(n_343)
);

AOI22xp5_ASAP7_75t_SL g377 ( 
.A1(n_298),
.A2(n_322),
.B1(n_294),
.B2(n_292),
.Y(n_377)
);

CKINVDCx16_ASAP7_75t_R g376 ( 
.A(n_304),
.Y(n_376)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_248),
.A2(n_196),
.B1(n_244),
.B2(n_210),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_L g350 ( 
.A1(n_306),
.A2(n_308),
.B1(n_313),
.B2(n_314),
.Y(n_350)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_213),
.A2(n_251),
.B1(n_243),
.B2(n_233),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_230),
.B(n_215),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g348 ( 
.A(n_312),
.B(n_206),
.C(n_222),
.Y(n_348)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_234),
.A2(n_237),
.B1(n_275),
.B2(n_208),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_258),
.B(n_224),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_320),
.B(n_325),
.Y(n_342)
);

OAI21xp33_ASAP7_75t_SL g322 ( 
.A1(n_263),
.A2(n_221),
.B(n_264),
.Y(n_322)
);

AOI21xp5_ASAP7_75t_L g346 ( 
.A1(n_323),
.A2(n_207),
.B(n_257),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_225),
.B(n_232),
.Y(n_325)
);

AOI22xp33_ASAP7_75t_SL g327 ( 
.A1(n_211),
.A2(n_261),
.B1(n_246),
.B2(n_260),
.Y(n_327)
);

AOI22xp33_ASAP7_75t_SL g361 ( 
.A1(n_327),
.A2(n_252),
.B1(n_290),
.B2(n_278),
.Y(n_361)
);

OAI22xp5_ASAP7_75t_L g329 ( 
.A1(n_265),
.A2(n_276),
.B1(n_267),
.B2(n_241),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_303),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g379 ( 
.A(n_335),
.B(n_351),
.Y(n_379)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_299),
.Y(n_336)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_336),
.Y(n_378)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_299),
.Y(n_337)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_337),
.Y(n_383)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_305),
.Y(n_338)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_338),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_288),
.B(n_229),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_339),
.B(n_340),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_288),
.B(n_216),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_312),
.B(n_242),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_341),
.B(n_355),
.Y(n_386)
);

OAI22xp5_ASAP7_75t_L g401 ( 
.A1(n_344),
.A2(n_359),
.B1(n_321),
.B2(n_285),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_279),
.B(n_239),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_SL g390 ( 
.A(n_345),
.B(n_349),
.Y(n_390)
);

OAI21xp5_ASAP7_75t_SL g407 ( 
.A1(n_346),
.A2(n_377),
.B(n_321),
.Y(n_407)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_305),
.Y(n_347)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_347),
.Y(n_408)
);

MAJIxp5_ASAP7_75t_L g380 ( 
.A(n_348),
.B(n_363),
.C(n_372),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_280),
.B(n_253),
.Y(n_349)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_333),
.Y(n_351)
);

AOI21xp5_ASAP7_75t_L g352 ( 
.A1(n_290),
.A2(n_323),
.B(n_314),
.Y(n_352)
);

AOI21xp5_ASAP7_75t_L g405 ( 
.A1(n_352),
.A2(n_361),
.B(n_365),
.Y(n_405)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_333),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_L g389 ( 
.A(n_353),
.B(n_354),
.Y(n_389)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_287),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_331),
.B(n_268),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_331),
.B(n_262),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_356),
.B(n_358),
.Y(n_388)
);

INVx3_ASAP7_75t_L g357 ( 
.A(n_295),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_L g393 ( 
.A(n_357),
.B(n_360),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_L g358 ( 
.A(n_280),
.B(n_283),
.Y(n_358)
);

AOI22xp5_ASAP7_75t_L g359 ( 
.A1(n_281),
.A2(n_255),
.B1(n_259),
.B2(n_252),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g360 ( 
.A(n_316),
.Y(n_360)
);

CKINVDCx20_ASAP7_75t_R g362 ( 
.A(n_291),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_L g403 ( 
.A(n_362),
.B(n_369),
.Y(n_403)
);

MAJIxp5_ASAP7_75t_SL g363 ( 
.A(n_282),
.B(n_296),
.C(n_301),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_301),
.B(n_326),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_364),
.B(n_366),
.Y(n_404)
);

AOI21xp5_ASAP7_75t_L g365 ( 
.A1(n_282),
.A2(n_286),
.B(n_307),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_SL g366 ( 
.A(n_326),
.B(n_313),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_308),
.B(n_282),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_367),
.B(n_368),
.Y(n_411)
);

NOR2xp33_ASAP7_75t_L g368 ( 
.A(n_289),
.B(n_287),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_297),
.Y(n_369)
);

INVx8_ASAP7_75t_L g370 ( 
.A(n_315),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_L g406 ( 
.A(n_370),
.B(n_371),
.Y(n_406)
);

CKINVDCx20_ASAP7_75t_R g371 ( 
.A(n_311),
.Y(n_371)
);

MAJIxp5_ASAP7_75t_L g372 ( 
.A(n_296),
.B(n_306),
.C(n_297),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_284),
.B(n_309),
.Y(n_373)
);

XNOR2xp5_ASAP7_75t_L g384 ( 
.A(n_373),
.B(n_293),
.Y(n_384)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_309),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_L g412 ( 
.A(n_374),
.B(n_375),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_L g375 ( 
.A(n_330),
.B(n_319),
.Y(n_375)
);

CKINVDCx16_ASAP7_75t_R g381 ( 
.A(n_373),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_L g437 ( 
.A(n_381),
.B(n_385),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_384),
.B(n_394),
.Y(n_421)
);

CKINVDCx20_ASAP7_75t_R g385 ( 
.A(n_368),
.Y(n_385)
);

MAJIxp5_ASAP7_75t_L g387 ( 
.A(n_341),
.B(n_293),
.C(n_324),
.Y(n_387)
);

XNOR2xp5_ASAP7_75t_L g423 ( 
.A(n_387),
.B(n_391),
.Y(n_423)
);

MAJIxp5_ASAP7_75t_L g391 ( 
.A(n_339),
.B(n_293),
.C(n_324),
.Y(n_391)
);

MAJIxp5_ASAP7_75t_L g392 ( 
.A(n_340),
.B(n_292),
.C(n_330),
.Y(n_392)
);

XNOR2xp5_ASAP7_75t_L g429 ( 
.A(n_392),
.B(n_396),
.Y(n_429)
);

CKINVDCx20_ASAP7_75t_R g394 ( 
.A(n_375),
.Y(n_394)
);

MAJIxp5_ASAP7_75t_L g396 ( 
.A(n_348),
.B(n_292),
.C(n_328),
.Y(n_396)
);

MAJIxp5_ASAP7_75t_L g397 ( 
.A(n_367),
.B(n_310),
.C(n_328),
.Y(n_397)
);

XOR2xp5_ASAP7_75t_L g443 ( 
.A(n_397),
.B(n_359),
.Y(n_443)
);

AOI22xp5_ASAP7_75t_L g398 ( 
.A1(n_350),
.A2(n_294),
.B1(n_318),
.B2(n_295),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_398),
.B(n_399),
.Y(n_424)
);

CKINVDCx20_ASAP7_75t_R g399 ( 
.A(n_358),
.Y(n_399)
);

XOR2xp5_ASAP7_75t_L g400 ( 
.A(n_364),
.B(n_315),
.Y(n_400)
);

XNOR2xp5_ASAP7_75t_SL g426 ( 
.A(n_400),
.B(n_363),
.Y(n_426)
);

AOI22xp5_ASAP7_75t_L g415 ( 
.A1(n_401),
.A2(n_414),
.B1(n_343),
.B2(n_334),
.Y(n_415)
);

AOI22xp5_ASAP7_75t_L g402 ( 
.A1(n_350),
.A2(n_318),
.B1(n_317),
.B2(n_319),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_402),
.B(n_410),
.Y(n_425)
);

OAI21xp5_ASAP7_75t_L g418 ( 
.A1(n_407),
.A2(n_409),
.B(n_413),
.Y(n_418)
);

AOI21xp5_ASAP7_75t_L g409 ( 
.A1(n_352),
.A2(n_332),
.B(n_315),
.Y(n_409)
);

CKINVDCx20_ASAP7_75t_R g410 ( 
.A(n_355),
.Y(n_410)
);

OAI21xp5_ASAP7_75t_L g413 ( 
.A1(n_346),
.A2(n_278),
.B(n_332),
.Y(n_413)
);

OAI22xp5_ASAP7_75t_SL g414 ( 
.A1(n_377),
.A2(n_366),
.B1(n_372),
.B2(n_356),
.Y(n_414)
);

OAI22xp5_ASAP7_75t_L g465 ( 
.A1(n_415),
.A2(n_430),
.B1(n_433),
.B2(n_434),
.Y(n_465)
);

CKINVDCx20_ASAP7_75t_R g416 ( 
.A(n_389),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_SL g464 ( 
.A(n_416),
.B(n_419),
.Y(n_464)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_389),
.Y(n_417)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_417),
.Y(n_448)
);

NOR2xp33_ASAP7_75t_SL g419 ( 
.A(n_399),
.B(n_342),
.Y(n_419)
);

OAI32xp33_ASAP7_75t_L g420 ( 
.A1(n_411),
.A2(n_342),
.A3(n_343),
.B1(n_345),
.B2(n_334),
.Y(n_420)
);

INVxp67_ASAP7_75t_L g455 ( 
.A(n_420),
.Y(n_455)
);

CKINVDCx20_ASAP7_75t_R g422 ( 
.A(n_379),
.Y(n_422)
);

CKINVDCx20_ASAP7_75t_R g462 ( 
.A(n_422),
.Y(n_462)
);

XNOR2x1_ASAP7_75t_L g461 ( 
.A(n_426),
.B(n_436),
.Y(n_461)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_378),
.Y(n_427)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_427),
.Y(n_474)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_378),
.Y(n_428)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_428),
.Y(n_458)
);

AOI22xp5_ASAP7_75t_SL g430 ( 
.A1(n_414),
.A2(n_376),
.B1(n_362),
.B2(n_335),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_383),
.Y(n_431)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_431),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_381),
.B(n_351),
.Y(n_432)
);

CKINVDCx20_ASAP7_75t_R g463 ( 
.A(n_432),
.Y(n_463)
);

AOI22xp5_ASAP7_75t_L g433 ( 
.A1(n_410),
.A2(n_376),
.B1(n_365),
.B2(n_353),
.Y(n_433)
);

AOI22xp5_ASAP7_75t_L g434 ( 
.A1(n_401),
.A2(n_354),
.B1(n_369),
.B2(n_371),
.Y(n_434)
);

HB1xp67_ASAP7_75t_L g435 ( 
.A(n_406),
.Y(n_435)
);

CKINVDCx16_ASAP7_75t_R g452 ( 
.A(n_435),
.Y(n_452)
);

AOI22xp5_ASAP7_75t_SL g436 ( 
.A1(n_385),
.A2(n_360),
.B1(n_357),
.B2(n_338),
.Y(n_436)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_393),
.Y(n_438)
);

AOI21xp33_ASAP7_75t_L g470 ( 
.A1(n_438),
.A2(n_440),
.B(n_442),
.Y(n_470)
);

AOI22xp5_ASAP7_75t_L g439 ( 
.A1(n_411),
.A2(n_394),
.B1(n_397),
.B2(n_404),
.Y(n_439)
);

OAI22xp5_ASAP7_75t_SL g456 ( 
.A1(n_439),
.A2(n_441),
.B1(n_386),
.B2(n_388),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_379),
.B(n_337),
.Y(n_440)
);

AOI22xp5_ASAP7_75t_L g441 ( 
.A1(n_404),
.A2(n_344),
.B1(n_347),
.B2(n_336),
.Y(n_441)
);

OAI21xp5_ASAP7_75t_L g442 ( 
.A1(n_405),
.A2(n_349),
.B(n_374),
.Y(n_442)
);

MAJIxp5_ASAP7_75t_L g450 ( 
.A(n_443),
.B(n_380),
.C(n_396),
.Y(n_450)
);

CKINVDCx20_ASAP7_75t_R g444 ( 
.A(n_393),
.Y(n_444)
);

AOI21xp5_ASAP7_75t_L g467 ( 
.A1(n_444),
.A2(n_412),
.B(n_384),
.Y(n_467)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_383),
.Y(n_445)
);

AOI22xp5_ASAP7_75t_SL g447 ( 
.A1(n_445),
.A2(n_395),
.B1(n_408),
.B2(n_390),
.Y(n_447)
);

NAND2xp33_ASAP7_75t_R g446 ( 
.A(n_388),
.B(n_370),
.Y(n_446)
);

XNOR2xp5_ASAP7_75t_L g453 ( 
.A(n_446),
.B(n_409),
.Y(n_453)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_447),
.Y(n_475)
);

OAI22xp33_ASAP7_75t_L g449 ( 
.A1(n_424),
.A2(n_402),
.B1(n_398),
.B2(n_407),
.Y(n_449)
);

AOI22xp5_ASAP7_75t_L g481 ( 
.A1(n_449),
.A2(n_457),
.B1(n_459),
.B2(n_472),
.Y(n_481)
);

MAJIxp5_ASAP7_75t_L g480 ( 
.A(n_450),
.B(n_451),
.C(n_423),
.Y(n_480)
);

MAJIxp5_ASAP7_75t_L g451 ( 
.A(n_429),
.B(n_380),
.C(n_400),
.Y(n_451)
);

AOI21xp5_ASAP7_75t_L g495 ( 
.A1(n_453),
.A2(n_433),
.B(n_436),
.Y(n_495)
);

XOR2xp5_ASAP7_75t_L g454 ( 
.A(n_423),
.B(n_400),
.Y(n_454)
);

XOR2xp5_ASAP7_75t_L g485 ( 
.A(n_454),
.B(n_429),
.Y(n_485)
);

NOR2xp33_ASAP7_75t_L g492 ( 
.A(n_456),
.B(n_459),
.Y(n_492)
);

OAI22xp5_ASAP7_75t_SL g457 ( 
.A1(n_430),
.A2(n_405),
.B1(n_386),
.B2(n_403),
.Y(n_457)
);

OAI22xp5_ASAP7_75t_SL g459 ( 
.A1(n_415),
.A2(n_403),
.B1(n_382),
.B2(n_406),
.Y(n_459)
);

AOI22xp5_ASAP7_75t_L g460 ( 
.A1(n_424),
.A2(n_413),
.B1(n_390),
.B2(n_387),
.Y(n_460)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_460),
.Y(n_476)
);

XNOR2x1_ASAP7_75t_L g466 ( 
.A(n_426),
.B(n_392),
.Y(n_466)
);

XNOR2xp5_ASAP7_75t_SL g494 ( 
.A(n_466),
.B(n_421),
.Y(n_494)
);

OAI21xp5_ASAP7_75t_SL g488 ( 
.A1(n_467),
.A2(n_468),
.B(n_432),
.Y(n_488)
);

A2O1A1Ixp33_ASAP7_75t_SL g468 ( 
.A1(n_418),
.A2(n_408),
.B(n_395),
.C(n_412),
.Y(n_468)
);

AOI22xp5_ASAP7_75t_L g469 ( 
.A1(n_425),
.A2(n_391),
.B1(n_382),
.B2(n_370),
.Y(n_469)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_469),
.Y(n_478)
);

OAI22xp5_ASAP7_75t_SL g472 ( 
.A1(n_439),
.A2(n_441),
.B1(n_425),
.B2(n_434),
.Y(n_472)
);

AOI22xp5_ASAP7_75t_L g473 ( 
.A1(n_443),
.A2(n_317),
.B1(n_300),
.B2(n_310),
.Y(n_473)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_473),
.Y(n_483)
);

CKINVDCx20_ASAP7_75t_R g477 ( 
.A(n_462),
.Y(n_477)
);

CKINVDCx20_ASAP7_75t_R g520 ( 
.A(n_477),
.Y(n_520)
);

CKINVDCx5p33_ASAP7_75t_R g479 ( 
.A(n_452),
.Y(n_479)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_479),
.Y(n_509)
);

MAJIxp5_ASAP7_75t_L g501 ( 
.A(n_480),
.B(n_493),
.C(n_496),
.Y(n_501)
);

AOI22xp5_ASAP7_75t_L g482 ( 
.A1(n_472),
.A2(n_442),
.B1(n_418),
.B2(n_417),
.Y(n_482)
);

OAI22xp5_ASAP7_75t_L g505 ( 
.A1(n_482),
.A2(n_498),
.B1(n_499),
.B2(n_481),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_SL g484 ( 
.A(n_464),
.B(n_437),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_SL g518 ( 
.A(n_484),
.B(n_491),
.Y(n_518)
);

XOR2xp5_ASAP7_75t_L g508 ( 
.A(n_485),
.B(n_487),
.Y(n_508)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_448),
.Y(n_486)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_486),
.Y(n_502)
);

XOR2xp5_ASAP7_75t_L g487 ( 
.A(n_451),
.B(n_420),
.Y(n_487)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_488),
.Y(n_519)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_458),
.Y(n_489)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_489),
.Y(n_506)
);

NOR2xp33_ASAP7_75t_SL g490 ( 
.A(n_467),
.B(n_440),
.Y(n_490)
);

NOR2xp33_ASAP7_75t_SL g511 ( 
.A(n_490),
.B(n_470),
.Y(n_511)
);

CKINVDCx16_ASAP7_75t_R g491 ( 
.A(n_447),
.Y(n_491)
);

XNOR2xp5_ASAP7_75t_L g504 ( 
.A(n_492),
.B(n_456),
.Y(n_504)
);

MAJIxp5_ASAP7_75t_L g493 ( 
.A(n_450),
.B(n_454),
.C(n_466),
.Y(n_493)
);

XOR2xp5_ASAP7_75t_L g516 ( 
.A(n_494),
.B(n_495),
.Y(n_516)
);

MAJIxp5_ASAP7_75t_L g496 ( 
.A(n_473),
.B(n_421),
.C(n_431),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_471),
.Y(n_497)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_497),
.Y(n_512)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_474),
.Y(n_498)
);

INVx2_ASAP7_75t_SL g499 ( 
.A(n_474),
.Y(n_499)
);

NOR2xp33_ASAP7_75t_L g500 ( 
.A(n_477),
.B(n_469),
.Y(n_500)
);

NOR2xp33_ASAP7_75t_SL g533 ( 
.A(n_500),
.B(n_515),
.Y(n_533)
);

MAJIxp5_ASAP7_75t_L g503 ( 
.A(n_480),
.B(n_460),
.C(n_461),
.Y(n_503)
);

MAJIxp5_ASAP7_75t_L g521 ( 
.A(n_503),
.B(n_510),
.C(n_513),
.Y(n_521)
);

XNOR2xp5_ASAP7_75t_L g529 ( 
.A(n_504),
.B(n_514),
.Y(n_529)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_505),
.Y(n_522)
);

FAx1_ASAP7_75t_SL g507 ( 
.A(n_488),
.B(n_455),
.CI(n_465),
.CON(n_507),
.SN(n_507)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_507),
.B(n_482),
.Y(n_524)
);

MAJIxp5_ASAP7_75t_L g510 ( 
.A(n_485),
.B(n_461),
.C(n_468),
.Y(n_510)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_511),
.Y(n_527)
);

MAJIxp5_ASAP7_75t_L g513 ( 
.A(n_493),
.B(n_468),
.C(n_457),
.Y(n_513)
);

XNOR2xp5_ASAP7_75t_L g514 ( 
.A(n_487),
.B(n_453),
.Y(n_514)
);

NOR2xp33_ASAP7_75t_L g515 ( 
.A(n_476),
.B(n_463),
.Y(n_515)
);

MAJIxp5_ASAP7_75t_L g517 ( 
.A(n_476),
.B(n_468),
.C(n_455),
.Y(n_517)
);

MAJIxp5_ASAP7_75t_L g525 ( 
.A(n_517),
.B(n_513),
.C(n_510),
.Y(n_525)
);

XOR2xp5_ASAP7_75t_L g523 ( 
.A(n_514),
.B(n_496),
.Y(n_523)
);

AND2x2_ASAP7_75t_L g543 ( 
.A(n_523),
.B(n_508),
.Y(n_543)
);

OAI21xp5_ASAP7_75t_L g546 ( 
.A1(n_524),
.A2(n_526),
.B(n_507),
.Y(n_546)
);

AOI22xp5_ASAP7_75t_SL g547 ( 
.A1(n_525),
.A2(n_503),
.B1(n_516),
.B2(n_499),
.Y(n_547)
);

AOI21xp5_ASAP7_75t_SL g526 ( 
.A1(n_519),
.A2(n_475),
.B(n_478),
.Y(n_526)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_509),
.Y(n_528)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_528),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_509),
.B(n_498),
.Y(n_530)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_530),
.Y(n_549)
);

AOI21xp5_ASAP7_75t_L g531 ( 
.A1(n_519),
.A2(n_517),
.B(n_495),
.Y(n_531)
);

OAI21x1_ASAP7_75t_SL g541 ( 
.A1(n_531),
.A2(n_530),
.B(n_479),
.Y(n_541)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_502),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_L g545 ( 
.A(n_532),
.B(n_534),
.Y(n_545)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_506),
.Y(n_534)
);

XNOR2xp5_ASAP7_75t_L g535 ( 
.A(n_501),
.B(n_481),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_L g548 ( 
.A(n_535),
.B(n_507),
.Y(n_548)
);

OAI22xp5_ASAP7_75t_SL g536 ( 
.A1(n_518),
.A2(n_478),
.B1(n_475),
.B2(n_483),
.Y(n_536)
);

AOI22xp5_ASAP7_75t_L g538 ( 
.A1(n_536),
.A2(n_483),
.B1(n_522),
.B2(n_524),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_L g556 ( 
.A(n_538),
.B(n_539),
.Y(n_556)
);

MAJIxp5_ASAP7_75t_L g539 ( 
.A(n_535),
.B(n_501),
.C(n_508),
.Y(n_539)
);

AOI22xp5_ASAP7_75t_L g540 ( 
.A1(n_536),
.A2(n_449),
.B1(n_516),
.B2(n_499),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_L g559 ( 
.A(n_540),
.B(n_542),
.Y(n_559)
);

XNOR2xp5_ASAP7_75t_L g553 ( 
.A(n_541),
.B(n_543),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_SL g542 ( 
.A(n_527),
.B(n_520),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_SL g544 ( 
.A(n_521),
.B(n_504),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_SL g551 ( 
.A(n_544),
.B(n_548),
.Y(n_551)
);

NOR2xp33_ASAP7_75t_L g550 ( 
.A(n_546),
.B(n_533),
.Y(n_550)
);

MAJIxp5_ASAP7_75t_L g555 ( 
.A(n_547),
.B(n_525),
.C(n_521),
.Y(n_555)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_550),
.Y(n_565)
);

CKINVDCx20_ASAP7_75t_R g552 ( 
.A(n_545),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_L g560 ( 
.A(n_552),
.B(n_554),
.Y(n_560)
);

NOR2xp33_ASAP7_75t_L g554 ( 
.A(n_538),
.B(n_529),
.Y(n_554)
);

MAJIxp5_ASAP7_75t_L g566 ( 
.A(n_555),
.B(n_543),
.C(n_529),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_SL g557 ( 
.A(n_539),
.B(n_523),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_L g561 ( 
.A(n_557),
.B(n_558),
.Y(n_561)
);

INVx6_ASAP7_75t_L g558 ( 
.A(n_547),
.Y(n_558)
);

NOR2xp33_ASAP7_75t_L g562 ( 
.A(n_553),
.B(n_549),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_SL g572 ( 
.A(n_562),
.B(n_566),
.Y(n_572)
);

NOR2xp33_ASAP7_75t_SL g563 ( 
.A(n_551),
.B(n_537),
.Y(n_563)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_563),
.Y(n_569)
);

INVxp67_ASAP7_75t_L g564 ( 
.A(n_556),
.Y(n_564)
);

AOI221xp5_ASAP7_75t_L g570 ( 
.A1(n_564),
.A2(n_567),
.B1(n_546),
.B2(n_553),
.C(n_558),
.Y(n_570)
);

INVxp67_ASAP7_75t_L g567 ( 
.A(n_555),
.Y(n_567)
);

NOR2xp33_ASAP7_75t_L g568 ( 
.A(n_560),
.B(n_559),
.Y(n_568)
);

AOI21xp5_ASAP7_75t_L g573 ( 
.A1(n_568),
.A2(n_561),
.B(n_564),
.Y(n_573)
);

AOI21xp5_ASAP7_75t_SL g574 ( 
.A1(n_570),
.A2(n_540),
.B(n_486),
.Y(n_574)
);

A2O1A1Ixp33_ASAP7_75t_SL g571 ( 
.A1(n_565),
.A2(n_531),
.B(n_526),
.C(n_468),
.Y(n_571)
);

MAJIxp5_ASAP7_75t_L g575 ( 
.A(n_571),
.B(n_494),
.C(n_512),
.Y(n_575)
);

OAI221xp5_ASAP7_75t_L g576 ( 
.A1(n_573),
.A2(n_574),
.B1(n_575),
.B2(n_569),
.C(n_572),
.Y(n_576)
);

AOI21xp5_ASAP7_75t_SL g578 ( 
.A1(n_576),
.A2(n_577),
.B(n_277),
.Y(n_578)
);

AOI322xp5_ASAP7_75t_L g577 ( 
.A1(n_573),
.A2(n_497),
.A3(n_489),
.B1(n_427),
.B2(n_428),
.C1(n_445),
.C2(n_277),
.Y(n_577)
);

XOR2xp5_ASAP7_75t_L g579 ( 
.A(n_578),
.B(n_300),
.Y(n_579)
);

XOR2xp5_ASAP7_75t_L g580 ( 
.A(n_579),
.B(n_302),
.Y(n_580)
);


endmodule