module fake_ibex_1194_n_190 (n_7, n_20, n_17, n_25, n_36, n_18, n_3, n_22, n_28, n_32, n_4, n_33, n_5, n_11, n_30, n_6, n_29, n_13, n_2, n_8, n_26, n_35, n_14, n_0, n_9, n_34, n_12, n_15, n_37, n_24, n_31, n_10, n_23, n_21, n_27, n_19, n_16, n_1, n_190);

input n_7;
input n_20;
input n_17;
input n_25;
input n_36;
input n_18;
input n_3;
input n_22;
input n_28;
input n_32;
input n_4;
input n_33;
input n_5;
input n_11;
input n_30;
input n_6;
input n_29;
input n_13;
input n_2;
input n_8;
input n_26;
input n_35;
input n_14;
input n_0;
input n_9;
input n_34;
input n_12;
input n_15;
input n_37;
input n_24;
input n_31;
input n_10;
input n_23;
input n_21;
input n_27;
input n_19;
input n_16;
input n_1;

output n_190;

wire n_151;
wire n_147;
wire n_85;
wire n_167;
wire n_128;
wire n_84;
wire n_64;
wire n_73;
wire n_152;
wire n_171;
wire n_145;
wire n_65;
wire n_103;
wire n_95;
wire n_139;
wire n_55;
wire n_130;
wire n_63;
wire n_98;
wire n_129;
wire n_161;
wire n_143;
wire n_106;
wire n_177;
wire n_148;
wire n_76;
wire n_118;
wire n_183;
wire n_67;
wire n_164;
wire n_38;
wire n_124;
wire n_110;
wire n_47;
wire n_169;
wire n_108;
wire n_82;
wire n_165;
wire n_78;
wire n_60;
wire n_86;
wire n_70;
wire n_109;
wire n_69;
wire n_87;
wire n_75;
wire n_127;
wire n_121;
wire n_175;
wire n_137;
wire n_48;
wire n_57;
wire n_59;
wire n_125;
wire n_39;
wire n_178;
wire n_62;
wire n_71;
wire n_153;
wire n_173;
wire n_120;
wire n_93;
wire n_168;
wire n_155;
wire n_162;
wire n_180;
wire n_122;
wire n_116;
wire n_61;
wire n_94;
wire n_134;
wire n_42;
wire n_77;
wire n_112;
wire n_150;
wire n_88;
wire n_133;
wire n_44;
wire n_142;
wire n_51;
wire n_46;
wire n_80;
wire n_172;
wire n_49;
wire n_66;
wire n_40;
wire n_90;
wire n_74;
wire n_176;
wire n_58;
wire n_43;
wire n_140;
wire n_136;
wire n_119;
wire n_100;
wire n_179;
wire n_72;
wire n_166;
wire n_163;
wire n_188;
wire n_114;
wire n_97;
wire n_102;
wire n_181;
wire n_131;
wire n_123;
wire n_52;
wire n_189;
wire n_99;
wire n_135;
wire n_105;
wire n_156;
wire n_126;
wire n_187;
wire n_154;
wire n_182;
wire n_111;
wire n_104;
wire n_41;
wire n_141;
wire n_89;
wire n_83;
wire n_53;
wire n_107;
wire n_115;
wire n_149;
wire n_54;
wire n_186;
wire n_50;
wire n_92;
wire n_144;
wire n_170;
wire n_101;
wire n_113;
wire n_138;
wire n_96;
wire n_185;
wire n_68;
wire n_117;
wire n_79;
wire n_81;
wire n_159;
wire n_158;
wire n_132;
wire n_174;
wire n_157;
wire n_160;
wire n_184;
wire n_56;
wire n_146;
wire n_91;
wire n_45;

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_12),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_21),
.Y(n_39)
);

INVxp67_ASAP7_75t_SL g40 ( 
.A(n_24),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_18),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_11),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_20),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_4),
.Y(n_44)
);

CKINVDCx5p33_ASAP7_75t_R g45 ( 
.A(n_37),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_7),
.Y(n_46)
);

CKINVDCx5p33_ASAP7_75t_R g47 ( 
.A(n_34),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_8),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_28),
.Y(n_49)
);

INVxp67_ASAP7_75t_L g50 ( 
.A(n_13),
.Y(n_50)
);

BUFx10_ASAP7_75t_L g51 ( 
.A(n_33),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_31),
.Y(n_52)
);

INVxp33_ASAP7_75t_SL g53 ( 
.A(n_26),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_25),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_5),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_27),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_10),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_4),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_22),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_5),
.B(n_16),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_15),
.Y(n_61)
);

HB1xp67_ASAP7_75t_L g62 ( 
.A(n_23),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_19),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_1),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_1),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_14),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_9),
.Y(n_67)
);

HB1xp67_ASAP7_75t_L g68 ( 
.A(n_7),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_3),
.Y(n_69)
);

BUFx2_ASAP7_75t_L g70 ( 
.A(n_35),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_30),
.Y(n_71)
);

CKINVDCx5p33_ASAP7_75t_R g72 ( 
.A(n_6),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_6),
.Y(n_73)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_41),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_42),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_38),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_41),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_62),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_39),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_70),
.B(n_0),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_42),
.Y(n_81)
);

AND2x4_ASAP7_75t_L g82 ( 
.A(n_48),
.B(n_73),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_68),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_L g84 ( 
.A1(n_57),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_38),
.A2(n_11),
.B1(n_17),
.B2(n_29),
.Y(n_85)
);

INVx1_ASAP7_75t_SL g86 ( 
.A(n_56),
.Y(n_86)
);

AND2x6_ASAP7_75t_L g87 ( 
.A(n_43),
.B(n_32),
.Y(n_87)
);

BUFx3_ASAP7_75t_L g88 ( 
.A(n_51),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_58),
.B(n_36),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_65),
.B(n_69),
.Y(n_90)
);

BUFx10_ASAP7_75t_L g91 ( 
.A(n_49),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_56),
.A2(n_59),
.B1(n_53),
.B2(n_72),
.Y(n_92)
);

BUFx3_ASAP7_75t_L g93 ( 
.A(n_51),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_50),
.B(n_66),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_54),
.Y(n_95)
);

AND2x6_ASAP7_75t_L g96 ( 
.A(n_61),
.B(n_71),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_51),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_63),
.Y(n_98)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_45),
.Y(n_99)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_47),
.Y(n_100)
);

AND2x6_ASAP7_75t_L g101 ( 
.A(n_60),
.B(n_40),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_55),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_55),
.Y(n_103)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_64),
.Y(n_104)
);

AND2x4_ASAP7_75t_L g105 ( 
.A(n_64),
.B(n_67),
.Y(n_105)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_67),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_44),
.Y(n_107)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_46),
.B(n_59),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_52),
.B(n_70),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_70),
.B(n_62),
.Y(n_110)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_62),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_97),
.B(n_93),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_110),
.B(n_111),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_88),
.B(n_91),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_91),
.B(n_110),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_78),
.B(n_100),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_99),
.B(n_83),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_94),
.B(n_98),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_94),
.B(n_82),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_79),
.B(n_95),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_79),
.B(n_95),
.Y(n_121)
);

NAND2xp33_ASAP7_75t_SL g122 ( 
.A(n_89),
.B(n_90),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_79),
.B(n_95),
.Y(n_123)
);

NAND2xp33_ASAP7_75t_SL g124 ( 
.A(n_89),
.B(n_84),
.Y(n_124)
);

AND2x4_ASAP7_75t_L g125 ( 
.A(n_74),
.B(n_80),
.Y(n_125)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_86),
.B(n_109),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_109),
.B(n_92),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_77),
.B(n_85),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_96),
.B(n_101),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_86),
.B(n_76),
.Y(n_130)
);

NAND2xp33_ASAP7_75t_SL g131 ( 
.A(n_84),
.B(n_76),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_102),
.B(n_103),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_104),
.B(n_106),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_105),
.B(n_108),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_105),
.B(n_96),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_96),
.B(n_87),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_96),
.B(n_87),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_87),
.B(n_101),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_87),
.B(n_101),
.Y(n_139)
);

NAND2xp33_ASAP7_75t_SL g140 ( 
.A(n_75),
.B(n_81),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_87),
.B(n_101),
.Y(n_141)
);

OAI21x1_ASAP7_75t_L g142 ( 
.A1(n_136),
.A2(n_101),
.B(n_107),
.Y(n_142)
);

AO21x2_ASAP7_75t_L g143 ( 
.A1(n_138),
.A2(n_141),
.B(n_139),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_L g144 ( 
.A1(n_137),
.A2(n_118),
.B(n_122),
.Y(n_144)
);

NAND2x1p5_ASAP7_75t_L g145 ( 
.A(n_135),
.B(n_128),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_113),
.B(n_119),
.Y(n_146)
);

AO31x2_ASAP7_75t_L g147 ( 
.A1(n_129),
.A2(n_124),
.A3(n_131),
.B(n_130),
.Y(n_147)
);

BUFx2_ASAP7_75t_L g148 ( 
.A(n_126),
.Y(n_148)
);

OR2x6_ASAP7_75t_L g149 ( 
.A(n_134),
.B(n_127),
.Y(n_149)
);

INVx3_ASAP7_75t_L g150 ( 
.A(n_125),
.Y(n_150)
);

AO31x2_ASAP7_75t_L g151 ( 
.A1(n_116),
.A2(n_117),
.A3(n_125),
.B(n_132),
.Y(n_151)
);

INVx1_ASAP7_75t_SL g152 ( 
.A(n_115),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_L g153 ( 
.A1(n_112),
.A2(n_125),
.B(n_120),
.Y(n_153)
);

AO21x1_ASAP7_75t_L g154 ( 
.A1(n_121),
.A2(n_123),
.B(n_133),
.Y(n_154)
);

OAI21x1_ASAP7_75t_L g155 ( 
.A1(n_114),
.A2(n_140),
.B(n_136),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_138),
.Y(n_156)
);

OR2x6_ASAP7_75t_L g157 ( 
.A(n_135),
.B(n_76),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_L g158 ( 
.A1(n_131),
.A2(n_124),
.B1(n_122),
.B2(n_128),
.Y(n_158)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_146),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_R g160 ( 
.A(n_148),
.B(n_150),
.Y(n_160)
);

BUFx3_ASAP7_75t_L g161 ( 
.A(n_156),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_150),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_150),
.Y(n_163)
);

NAND2xp33_ASAP7_75t_R g164 ( 
.A(n_148),
.B(n_157),
.Y(n_164)
);

INVx8_ASAP7_75t_L g165 ( 
.A(n_157),
.Y(n_165)
);

BUFx3_ASAP7_75t_L g166 ( 
.A(n_156),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_R g167 ( 
.A(n_152),
.B(n_158),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_147),
.Y(n_168)
);

NAND2xp33_ASAP7_75t_R g169 ( 
.A(n_157),
.B(n_149),
.Y(n_169)
);

NAND2xp33_ASAP7_75t_SL g170 ( 
.A(n_156),
.B(n_144),
.Y(n_170)
);

CKINVDCx16_ASAP7_75t_R g171 ( 
.A(n_157),
.Y(n_171)
);

OAI221xp5_ASAP7_75t_L g172 ( 
.A1(n_159),
.A2(n_149),
.B1(n_145),
.B2(n_153),
.C(n_156),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_162),
.Y(n_173)
);

AND2x2_ASAP7_75t_L g174 ( 
.A(n_171),
.B(n_147),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_163),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_R g176 ( 
.A(n_169),
.B(n_164),
.Y(n_176)
);

AND2x2_ASAP7_75t_L g177 ( 
.A(n_160),
.B(n_147),
.Y(n_177)
);

OAI33xp33_ASAP7_75t_L g178 ( 
.A1(n_168),
.A2(n_147),
.A3(n_149),
.B1(n_151),
.B2(n_155),
.B3(n_154),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_165),
.A2(n_142),
.B1(n_154),
.B2(n_143),
.Y(n_179)
);

NOR2x1_ASAP7_75t_L g180 ( 
.A(n_172),
.B(n_161),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_180),
.A2(n_165),
.B1(n_177),
.B2(n_174),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_181),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_182),
.A2(n_165),
.B1(n_174),
.B2(n_177),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_R g184 ( 
.A(n_183),
.B(n_182),
.Y(n_184)
);

AND2x4_ASAP7_75t_L g185 ( 
.A(n_184),
.B(n_179),
.Y(n_185)
);

HB1xp67_ASAP7_75t_L g186 ( 
.A(n_184),
.Y(n_186)
);

AOI22xp33_ASAP7_75t_L g187 ( 
.A1(n_186),
.A2(n_165),
.B1(n_176),
.B2(n_178),
.Y(n_187)
);

AOI22xp33_ASAP7_75t_L g188 ( 
.A1(n_185),
.A2(n_170),
.B1(n_167),
.B2(n_175),
.Y(n_188)
);

OAI22xp33_ASAP7_75t_L g189 ( 
.A1(n_187),
.A2(n_185),
.B1(n_175),
.B2(n_173),
.Y(n_189)
);

OAI221xp5_ASAP7_75t_L g190 ( 
.A1(n_189),
.A2(n_188),
.B1(n_170),
.B2(n_173),
.C(n_166),
.Y(n_190)
);


endmodule