module fake_jpeg_28797_n_142 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_142);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_142;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_15),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_23),
.Y(n_45)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_11),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_31),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_30),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_3),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_2),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_11),
.Y(n_51)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_32),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_3),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_2),
.Y(n_54)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_13),
.Y(n_55)
);

CKINVDCx14_ASAP7_75t_R g56 ( 
.A(n_43),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_33),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_16),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_22),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_27),
.Y(n_60)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_46),
.Y(n_61)
);

INVx8_ASAP7_75t_L g80 ( 
.A(n_61),
.Y(n_80)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_52),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_62),
.Y(n_70)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_52),
.Y(n_63)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_63),
.Y(n_83)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_55),
.Y(n_64)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_64),
.Y(n_76)
);

OR2x2_ASAP7_75t_L g65 ( 
.A(n_51),
.B(n_0),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_65),
.B(n_68),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_45),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_66),
.B(n_67),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_45),
.Y(n_67)
);

INVx1_ASAP7_75t_SL g68 ( 
.A(n_55),
.Y(n_68)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_60),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_69),
.B(n_60),
.Y(n_77)
);

BUFx4f_ASAP7_75t_SL g72 ( 
.A(n_62),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_72),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_68),
.A2(n_46),
.B1(n_60),
.B2(n_54),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_73),
.A2(n_79),
.B1(n_82),
.B2(n_0),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_65),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_74),
.B(n_78),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_77),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_61),
.B(n_53),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_69),
.A2(n_50),
.B1(n_49),
.B2(n_56),
.Y(n_79)
);

OA22x2_ASAP7_75t_SL g81 ( 
.A1(n_66),
.A2(n_26),
.B1(n_28),
.B2(n_42),
.Y(n_81)
);

O2A1O1Ixp33_ASAP7_75t_L g89 ( 
.A1(n_81),
.A2(n_59),
.B(n_58),
.C(n_48),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_67),
.A2(n_49),
.B1(n_50),
.B2(n_57),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_SL g84 ( 
.A1(n_71),
.A2(n_57),
.B(n_47),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_84),
.B(n_88),
.C(n_21),
.Y(n_104)
);

NOR2x1_ASAP7_75t_L g87 ( 
.A(n_81),
.B(n_44),
.Y(n_87)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_87),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_76),
.B(n_75),
.C(n_83),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_89),
.B(n_94),
.Y(n_102)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_76),
.Y(n_90)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_90),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_80),
.A2(n_63),
.B1(n_1),
.B2(n_4),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_91),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_92),
.B(n_72),
.Y(n_103)
);

AOI21xp5_ASAP7_75t_SL g93 ( 
.A1(n_81),
.A2(n_1),
.B(n_4),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_L g120 ( 
.A1(n_93),
.A2(n_13),
.B(n_14),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_83),
.B(n_5),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_80),
.A2(n_20),
.B1(n_40),
.B2(n_39),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_96),
.A2(n_9),
.B1(n_10),
.B2(n_12),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_75),
.B(n_5),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_97),
.B(n_7),
.Y(n_106)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_70),
.Y(n_98)
);

INVx13_ASAP7_75t_L g118 ( 
.A(n_98),
.Y(n_118)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_70),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_99),
.B(n_100),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_75),
.B(n_6),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_72),
.B(n_6),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_101),
.B(n_7),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_103),
.A2(n_95),
.B1(n_24),
.B2(n_25),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_104),
.B(n_111),
.C(n_113),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_89),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_105),
.B(n_106),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_88),
.B(n_19),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_107),
.B(n_109),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_85),
.B(n_8),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_110),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_98),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_112),
.A2(n_96),
.B1(n_91),
.B2(n_14),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_93),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_115),
.A2(n_120),
.B1(n_17),
.B2(n_34),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_86),
.B(n_12),
.Y(n_116)
);

INVxp33_ASAP7_75t_L g121 ( 
.A(n_116),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_87),
.B(n_29),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_117),
.B(n_95),
.C(n_18),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_122),
.B(n_123),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_124),
.A2(n_128),
.B1(n_103),
.B2(n_115),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_126),
.B(n_102),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_114),
.A2(n_35),
.B1(n_36),
.B2(n_37),
.Y(n_128)
);

A2O1A1Ixp33_ASAP7_75t_SL g135 ( 
.A1(n_131),
.A2(n_133),
.B(n_134),
.C(n_120),
.Y(n_135)
);

AO221x1_ASAP7_75t_L g134 ( 
.A1(n_129),
.A2(n_119),
.B1(n_118),
.B2(n_108),
.C(n_130),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_135),
.B(n_136),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_132),
.B(n_127),
.C(n_107),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_137),
.A2(n_131),
.B1(n_117),
.B2(n_134),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_L g139 ( 
.A1(n_138),
.A2(n_103),
.B(n_125),
.Y(n_139)
);

AOI322xp5_ASAP7_75t_L g140 ( 
.A1(n_139),
.A2(n_125),
.A3(n_118),
.B1(n_121),
.B2(n_104),
.C1(n_123),
.C2(n_106),
.Y(n_140)
);

AOI21xp33_ASAP7_75t_L g141 ( 
.A1(n_140),
.A2(n_121),
.B(n_38),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g142 ( 
.A(n_141),
.B(n_41),
.Y(n_142)
);


endmodule