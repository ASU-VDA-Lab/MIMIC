module fake_jpeg_4112_n_301 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_301);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_301;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_187;
wire n_21;
wire n_57;
wire n_288;
wire n_234;
wire n_284;
wire n_272;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_298;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_299;
wire n_211;
wire n_300;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_270;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_265;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

BUFx12_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_16),
.Y(n_18)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_16),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_16),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

INVx8_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_9),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_15),
.Y(n_28)
);

CKINVDCx14_ASAP7_75t_R g29 ( 
.A(n_15),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_8),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_11),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_19),
.B(n_7),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_SL g46 ( 
.A(n_35),
.B(n_18),
.Y(n_46)
);

HAxp5_ASAP7_75t_SL g36 ( 
.A(n_18),
.B(n_7),
.CON(n_36),
.SN(n_36)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_36),
.B(n_43),
.Y(n_65)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_33),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_37),
.B(n_42),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_33),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_33),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_39),
.Y(n_58)
);

BUFx12_ASAP7_75t_L g40 ( 
.A(n_32),
.Y(n_40)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_40),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_21),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_41),
.Y(n_64)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_21),
.Y(n_42)
);

INVx2_ASAP7_75t_R g43 ( 
.A(n_32),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g44 ( 
.A1(n_42),
.A2(n_24),
.B1(n_19),
.B2(n_30),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_44),
.A2(n_23),
.B1(n_34),
.B2(n_25),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_46),
.B(n_55),
.Y(n_72)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_43),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_48),
.B(n_50),
.Y(n_70)
);

CKINVDCx6p67_ASAP7_75t_R g49 ( 
.A(n_43),
.Y(n_49)
);

INVx1_ASAP7_75t_SL g85 ( 
.A(n_49),
.Y(n_85)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_43),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_43),
.A2(n_19),
.B1(n_24),
.B2(n_29),
.Y(n_51)
);

AOI21xp5_ASAP7_75t_L g78 ( 
.A1(n_51),
.A2(n_59),
.B(n_23),
.Y(n_78)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_42),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_52),
.B(n_57),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_35),
.B(n_29),
.Y(n_53)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_53),
.Y(n_80)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_35),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_56),
.B(n_61),
.Y(n_74)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_37),
.A2(n_24),
.B1(n_20),
.B2(n_23),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_36),
.B(n_18),
.Y(n_60)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_60),
.Y(n_90)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_39),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g62 ( 
.A(n_38),
.B(n_20),
.Y(n_62)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_62),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g63 ( 
.A(n_38),
.B(n_20),
.Y(n_63)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_63),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_41),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_66),
.Y(n_89)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_40),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_67),
.B(n_40),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g68 ( 
.A(n_49),
.B(n_30),
.Y(n_68)
);

OAI21xp5_ASAP7_75t_SL g95 ( 
.A1(n_68),
.A2(n_73),
.B(n_78),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_45),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_69),
.B(n_83),
.Y(n_98)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_49),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_71),
.B(n_75),
.Y(n_104)
);

AO22x1_ASAP7_75t_L g73 ( 
.A1(n_49),
.A2(n_41),
.B1(n_38),
.B2(n_39),
.Y(n_73)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_57),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_76),
.B(n_81),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_L g77 ( 
.A1(n_55),
.A2(n_34),
.B1(n_28),
.B2(n_25),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_77),
.A2(n_27),
.B1(n_31),
.B2(n_67),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_45),
.Y(n_81)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_54),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_82),
.B(n_84),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_46),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_49),
.B(n_40),
.C(n_39),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_86),
.B(n_58),
.C(n_61),
.Y(n_96)
);

BUFx12f_ASAP7_75t_L g87 ( 
.A(n_47),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_87),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_65),
.B(n_28),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_88),
.B(n_53),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_64),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_93),
.B(n_66),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_62),
.B(n_17),
.Y(n_94)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_94),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_96),
.B(n_97),
.C(n_117),
.Y(n_123)
);

XNOR2xp5_ASAP7_75t_L g97 ( 
.A(n_86),
.B(n_60),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_69),
.B(n_65),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_99),
.B(n_103),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_90),
.A2(n_48),
.B1(n_65),
.B2(n_50),
.Y(n_101)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_101),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_91),
.B(n_63),
.Y(n_103)
);

OR2x2_ASAP7_75t_L g105 ( 
.A(n_83),
.B(n_73),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_105),
.B(n_111),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_106),
.B(n_116),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_91),
.B(n_58),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_107),
.B(n_115),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_72),
.B(n_56),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_108),
.B(n_109),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_72),
.B(n_31),
.Y(n_109)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_73),
.Y(n_111)
);

CKINVDCx16_ASAP7_75t_R g143 ( 
.A(n_113),
.Y(n_143)
);

AND2x6_ASAP7_75t_L g114 ( 
.A(n_88),
.B(n_40),
.Y(n_114)
);

A2O1A1O1Ixp25_ASAP7_75t_L g134 ( 
.A1(n_114),
.A2(n_85),
.B(n_68),
.C(n_74),
.D(n_40),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_92),
.B(n_44),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_92),
.B(n_52),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_70),
.B(n_40),
.C(n_39),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_118),
.A2(n_120),
.B1(n_80),
.B2(n_76),
.Y(n_122)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_71),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_119),
.B(n_121),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_78),
.A2(n_47),
.B1(n_41),
.B2(n_31),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_79),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_122),
.B(n_128),
.Y(n_178)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_108),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_126),
.B(n_130),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_95),
.A2(n_90),
.B1(n_81),
.B2(n_80),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_127),
.A2(n_135),
.B1(n_141),
.B2(n_145),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_100),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_120),
.A2(n_88),
.B1(n_68),
.B2(n_85),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_129),
.A2(n_147),
.B1(n_122),
.B2(n_149),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_104),
.Y(n_130)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_98),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_133),
.B(n_137),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_134),
.B(n_26),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_114),
.A2(n_74),
.B1(n_75),
.B2(n_82),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_116),
.Y(n_137)
);

INVxp67_ASAP7_75t_L g140 ( 
.A(n_112),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_140),
.B(n_142),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_95),
.A2(n_41),
.B1(n_66),
.B2(n_64),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_SL g142 ( 
.A(n_98),
.B(n_27),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_100),
.B(n_54),
.Y(n_144)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_144),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_111),
.A2(n_64),
.B1(n_21),
.B2(n_39),
.Y(n_145)
);

CKINVDCx16_ASAP7_75t_R g146 ( 
.A(n_107),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_146),
.B(n_0),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_102),
.A2(n_101),
.B1(n_115),
.B2(n_99),
.Y(n_147)
);

BUFx5_ASAP7_75t_L g148 ( 
.A(n_100),
.Y(n_148)
);

INVx5_ASAP7_75t_L g172 ( 
.A(n_148),
.Y(n_172)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_118),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_149),
.B(n_10),
.Y(n_180)
);

INVx4_ASAP7_75t_L g150 ( 
.A(n_119),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_150),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_L g152 ( 
.A1(n_139),
.A2(n_102),
.B(n_103),
.Y(n_152)
);

AOI21xp5_ASAP7_75t_L g192 ( 
.A1(n_152),
.A2(n_157),
.B(n_158),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_123),
.B(n_96),
.C(n_117),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_153),
.B(n_154),
.C(n_161),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_123),
.B(n_106),
.C(n_110),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_126),
.B(n_110),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_155),
.B(n_156),
.Y(n_181)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_148),
.Y(n_156)
);

AND2x2_ASAP7_75t_L g157 ( 
.A(n_127),
.B(n_105),
.Y(n_157)
);

AOI21xp5_ASAP7_75t_L g158 ( 
.A1(n_132),
.A2(n_109),
.B(n_105),
.Y(n_158)
);

FAx1_ASAP7_75t_SL g203 ( 
.A(n_160),
.B(n_26),
.CI(n_22),
.CON(n_203),
.SN(n_203)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_147),
.B(n_97),
.C(n_121),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_138),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_162),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_132),
.A2(n_54),
.B1(n_21),
.B2(n_39),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_165),
.A2(n_125),
.B1(n_142),
.B2(n_89),
.Y(n_199)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_139),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_166),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_137),
.B(n_87),
.C(n_32),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_167),
.B(n_173),
.C(n_143),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_168),
.B(n_124),
.Y(n_188)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_170),
.Y(n_186)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_145),
.Y(n_171)
);

CKINVDCx14_ASAP7_75t_R g197 ( 
.A(n_171),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_124),
.B(n_87),
.C(n_32),
.Y(n_173)
);

AO22x1_ASAP7_75t_L g174 ( 
.A1(n_129),
.A2(n_32),
.B1(n_22),
.B2(n_26),
.Y(n_174)
);

OA21x2_ASAP7_75t_L g206 ( 
.A1(n_174),
.A2(n_175),
.B(n_179),
.Y(n_206)
);

OA21x2_ASAP7_75t_L g175 ( 
.A1(n_136),
.A2(n_17),
.B(n_22),
.Y(n_175)
);

INVx3_ASAP7_75t_L g177 ( 
.A(n_128),
.Y(n_177)
);

HB1xp67_ASAP7_75t_L g184 ( 
.A(n_177),
.Y(n_184)
);

AO21x2_ASAP7_75t_L g179 ( 
.A1(n_141),
.A2(n_87),
.B(n_17),
.Y(n_179)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_180),
.Y(n_191)
);

XNOR2x2_ASAP7_75t_L g183 ( 
.A(n_157),
.B(n_134),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_L g224 ( 
.A1(n_183),
.A2(n_175),
.B(n_26),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_163),
.A2(n_135),
.B1(n_146),
.B2(n_133),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_185),
.A2(n_200),
.B1(n_202),
.B2(n_179),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_187),
.B(n_188),
.C(n_198),
.Y(n_207)
);

HB1xp67_ASAP7_75t_L g189 ( 
.A(n_172),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_189),
.B(n_190),
.Y(n_215)
);

NOR4xp25_ASAP7_75t_L g190 ( 
.A(n_174),
.B(n_131),
.C(n_130),
.D(n_140),
.Y(n_190)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_176),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_193),
.B(n_194),
.Y(n_219)
);

CKINVDCx16_ASAP7_75t_R g194 ( 
.A(n_172),
.Y(n_194)
);

CKINVDCx16_ASAP7_75t_R g196 ( 
.A(n_178),
.Y(n_196)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_196),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_153),
.B(n_125),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_199),
.A2(n_179),
.B1(n_158),
.B2(n_154),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_163),
.A2(n_150),
.B1(n_93),
.B2(n_89),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_161),
.B(n_128),
.C(n_93),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_201),
.B(n_173),
.C(n_167),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_157),
.A2(n_179),
.B1(n_160),
.B2(n_168),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_203),
.B(n_175),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_152),
.A2(n_89),
.B1(n_26),
.B2(n_22),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_205),
.A2(n_151),
.B1(n_159),
.B2(n_177),
.Y(n_216)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_208),
.Y(n_237)
);

CKINVDCx14_ASAP7_75t_R g209 ( 
.A(n_181),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_209),
.B(n_211),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_193),
.B(n_169),
.Y(n_210)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_210),
.Y(n_233)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_212),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_214),
.A2(n_216),
.B1(n_191),
.B2(n_186),
.Y(n_240)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_200),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_217),
.B(n_220),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_182),
.B(n_165),
.C(n_164),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_218),
.B(n_221),
.Y(n_232)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_205),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_182),
.B(n_198),
.C(n_188),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_201),
.B(n_187),
.C(n_192),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_222),
.B(n_224),
.Y(n_234)
);

CKINVDCx14_ASAP7_75t_R g223 ( 
.A(n_199),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_223),
.B(n_229),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_204),
.B(n_156),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_225),
.B(n_226),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_195),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_192),
.B(n_22),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_227),
.B(n_228),
.Y(n_246)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_185),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_183),
.A2(n_17),
.B1(n_8),
.B2(n_9),
.Y(n_229)
);

AOI21xp5_ASAP7_75t_L g230 ( 
.A1(n_227),
.A2(n_202),
.B(n_206),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_L g249 ( 
.A1(n_230),
.A2(n_239),
.B(n_220),
.Y(n_249)
);

CKINVDCx14_ASAP7_75t_R g235 ( 
.A(n_219),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_235),
.B(n_245),
.Y(n_259)
);

OAI322xp33_ASAP7_75t_L g236 ( 
.A1(n_229),
.A2(n_203),
.A3(n_197),
.B1(n_206),
.B2(n_191),
.C1(n_186),
.C2(n_17),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_SL g252 ( 
.A(n_236),
.B(n_216),
.Y(n_252)
);

AOI21xp5_ASAP7_75t_L g239 ( 
.A1(n_228),
.A2(n_206),
.B(n_203),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_240),
.A2(n_247),
.B1(n_213),
.B2(n_215),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_226),
.B(n_184),
.Y(n_244)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_244),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_225),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_217),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_210),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_248),
.B(n_233),
.Y(n_261)
);

AOI21xp5_ASAP7_75t_L g265 ( 
.A1(n_249),
.A2(n_251),
.B(n_253),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_231),
.B(n_221),
.C(n_222),
.Y(n_251)
);

NAND3xp33_ASAP7_75t_L g273 ( 
.A(n_252),
.B(n_230),
.C(n_243),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_232),
.B(n_207),
.C(n_218),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_232),
.B(n_234),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_254),
.B(n_256),
.Y(n_264)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_242),
.Y(n_255)
);

AOI21xp5_ASAP7_75t_L g269 ( 
.A1(n_255),
.A2(n_257),
.B(n_238),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_SL g256 ( 
.A(n_246),
.B(n_212),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_242),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_234),
.B(n_207),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_258),
.B(n_254),
.Y(n_272)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_260),
.Y(n_263)
);

OAI21xp5_ASAP7_75t_L g268 ( 
.A1(n_261),
.A2(n_238),
.B(n_246),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_241),
.A2(n_208),
.B1(n_224),
.B2(n_213),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_262),
.A2(n_249),
.B1(n_237),
.B2(n_233),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_266),
.B(n_274),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_SL g267 ( 
.A(n_259),
.B(n_240),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_267),
.B(n_247),
.Y(n_275)
);

AOI21xp5_ASAP7_75t_L g278 ( 
.A1(n_268),
.A2(n_269),
.B(n_258),
.Y(n_278)
);

INVx4_ASAP7_75t_L g270 ( 
.A(n_256),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_270),
.A2(n_273),
.B1(n_9),
.B2(n_14),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_250),
.B(n_248),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_SL g279 ( 
.A(n_271),
.B(n_0),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_272),
.B(n_253),
.C(n_251),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_252),
.A2(n_241),
.B1(n_211),
.B2(n_239),
.Y(n_274)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_275),
.Y(n_289)
);

HB1xp67_ASAP7_75t_L g276 ( 
.A(n_270),
.Y(n_276)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_276),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_277),
.B(n_272),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_SL g288 ( 
.A(n_278),
.B(n_279),
.Y(n_288)
);

AOI21xp5_ASAP7_75t_L g280 ( 
.A1(n_265),
.A2(n_268),
.B(n_263),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_SL g287 ( 
.A(n_280),
.B(n_284),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_264),
.B(n_1),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_SL g285 ( 
.A(n_282),
.B(n_283),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_264),
.B(n_2),
.Y(n_284)
);

NOR2x1_ASAP7_75t_R g286 ( 
.A(n_281),
.B(n_273),
.Y(n_286)
);

NAND3xp33_ASAP7_75t_L g292 ( 
.A(n_286),
.B(n_288),
.C(n_285),
.Y(n_292)
);

OAI21xp5_ASAP7_75t_SL g295 ( 
.A1(n_290),
.A2(n_6),
.B(n_12),
.Y(n_295)
);

AOI322xp5_ASAP7_75t_L g298 ( 
.A1(n_292),
.A2(n_294),
.A3(n_296),
.B1(n_10),
.B2(n_13),
.C1(n_4),
.C2(n_2),
.Y(n_298)
);

OAI21xp5_ASAP7_75t_L g293 ( 
.A1(n_288),
.A2(n_275),
.B(n_3),
.Y(n_293)
);

AOI21xp5_ASAP7_75t_SL g297 ( 
.A1(n_293),
.A2(n_295),
.B(n_291),
.Y(n_297)
);

AOI322xp5_ASAP7_75t_L g294 ( 
.A1(n_287),
.A2(n_7),
.A3(n_14),
.B1(n_13),
.B2(n_5),
.C1(n_6),
.C2(n_15),
.Y(n_294)
);

AOI322xp5_ASAP7_75t_L g296 ( 
.A1(n_289),
.A2(n_6),
.A3(n_12),
.B1(n_10),
.B2(n_5),
.C1(n_13),
.C2(n_4),
.Y(n_296)
);

OAI31xp33_ASAP7_75t_L g299 ( 
.A1(n_297),
.A2(n_298),
.A3(n_3),
.B(n_4),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_299),
.B(n_3),
.C(n_4),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_300),
.B(n_3),
.Y(n_301)
);


endmodule