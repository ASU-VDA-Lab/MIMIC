module fake_jpeg_26558_n_337 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_337);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_337;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_9),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

BUFx16f_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

INVx8_ASAP7_75t_SL g30 ( 
.A(n_1),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_3),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_9),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_5),
.Y(n_35)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_25),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_36),
.Y(n_59)
);

INVx4_ASAP7_75t_SL g37 ( 
.A(n_30),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_37),
.B(n_29),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_38),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_39),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_40),
.Y(n_64)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_25),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_42),
.Y(n_66)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_25),
.Y(n_43)
);

HB1xp67_ASAP7_75t_L g57 ( 
.A(n_43),
.Y(n_57)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_30),
.Y(n_44)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_44),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_27),
.Y(n_45)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_45),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_29),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_46),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_46),
.Y(n_48)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_48),
.Y(n_72)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_44),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_50),
.Y(n_83)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_44),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_51),
.B(n_55),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_40),
.B(n_27),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_52),
.B(n_62),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_36),
.A2(n_27),
.B1(n_33),
.B2(n_17),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_54),
.A2(n_56),
.B1(n_43),
.B2(n_42),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g55 ( 
.A(n_45),
.B(n_21),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g56 ( 
.A1(n_36),
.A2(n_33),
.B1(n_16),
.B2(n_17),
.Y(n_56)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_46),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_58),
.Y(n_104)
);

OR2x2_ASAP7_75t_L g92 ( 
.A(n_61),
.B(n_48),
.Y(n_92)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_38),
.Y(n_62)
);

AND2x2_ASAP7_75t_SL g67 ( 
.A(n_62),
.B(n_38),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_67),
.B(n_70),
.C(n_91),
.Y(n_121)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_57),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_68),
.B(n_73),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_69),
.A2(n_105),
.B1(n_37),
.B2(n_16),
.Y(n_118)
);

AND2x2_ASAP7_75t_SL g70 ( 
.A(n_52),
.B(n_38),
.Y(n_70)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_56),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_54),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_74),
.B(n_78),
.Y(n_122)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_60),
.Y(n_75)
);

INVx1_ASAP7_75t_SL g117 ( 
.A(n_75),
.Y(n_117)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_63),
.Y(n_76)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_76),
.Y(n_133)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_63),
.Y(n_77)
);

BUFx2_ASAP7_75t_SL g123 ( 
.A(n_77),
.Y(n_123)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_65),
.Y(n_78)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_60),
.Y(n_79)
);

INVx1_ASAP7_75t_SL g119 ( 
.A(n_79),
.Y(n_119)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_65),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_80),
.B(n_81),
.Y(n_132)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_64),
.Y(n_81)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_64),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_82),
.B(n_84),
.Y(n_135)
);

INVx13_ASAP7_75t_L g84 ( 
.A(n_53),
.Y(n_84)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_59),
.Y(n_85)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_85),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_49),
.A2(n_33),
.B1(n_43),
.B2(n_42),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_86),
.A2(n_97),
.B1(n_16),
.B2(n_17),
.Y(n_128)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_47),
.Y(n_87)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_87),
.Y(n_109)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_53),
.Y(n_88)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_88),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_50),
.B(n_21),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_90),
.Y(n_111)
);

XNOR2xp5_ASAP7_75t_L g91 ( 
.A(n_47),
.B(n_45),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_92),
.B(n_46),
.Y(n_107)
);

INVx8_ASAP7_75t_L g93 ( 
.A(n_53),
.Y(n_93)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_93),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_59),
.B(n_23),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_94),
.B(n_96),
.Y(n_112)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_66),
.Y(n_95)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_95),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_L g96 ( 
.A(n_49),
.B(n_23),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_58),
.A2(n_33),
.B1(n_41),
.B2(n_31),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_66),
.B(n_31),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_98),
.Y(n_116)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_55),
.Y(n_99)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_99),
.Y(n_127)
);

INVx13_ASAP7_75t_L g100 ( 
.A(n_53),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_100),
.Y(n_120)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_63),
.Y(n_101)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_101),
.Y(n_129)
);

INVx2_ASAP7_75t_SL g102 ( 
.A(n_49),
.Y(n_102)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_102),
.Y(n_131)
);

BUFx8_ASAP7_75t_L g103 ( 
.A(n_48),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_103),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_L g105 ( 
.A1(n_52),
.A2(n_41),
.B1(n_45),
.B2(n_40),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_L g151 ( 
.A1(n_107),
.A2(n_72),
.B(n_20),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_L g110 ( 
.A1(n_89),
.A2(n_37),
.B1(n_39),
.B2(n_25),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_110),
.A2(n_130),
.B1(n_22),
.B2(n_19),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_70),
.B(n_39),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_115),
.B(n_32),
.Y(n_159)
);

AND2x2_ASAP7_75t_L g153 ( 
.A(n_118),
.B(n_83),
.Y(n_153)
);

AO22x2_ASAP7_75t_L g124 ( 
.A1(n_70),
.A2(n_39),
.B1(n_46),
.B2(n_37),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_124),
.A2(n_126),
.B1(n_97),
.B2(n_92),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_67),
.A2(n_24),
.B1(n_19),
.B2(n_20),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_128),
.A2(n_75),
.B1(n_79),
.B2(n_102),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_86),
.A2(n_19),
.B1(n_22),
.B2(n_23),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g136 ( 
.A(n_135),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_136),
.B(n_138),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_137),
.A2(n_143),
.B1(n_148),
.B2(n_153),
.Y(n_172)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_132),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_132),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_139),
.B(n_142),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g140 ( 
.A(n_121),
.B(n_91),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_140),
.B(n_146),
.C(n_131),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_SL g177 ( 
.A1(n_141),
.A2(n_150),
.B(n_161),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_135),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_118),
.A2(n_105),
.B1(n_67),
.B2(n_71),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_144),
.A2(n_156),
.B1(n_117),
.B2(n_119),
.Y(n_167)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_133),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_145),
.B(n_147),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_121),
.B(n_83),
.C(n_104),
.Y(n_146)
);

BUFx24_ASAP7_75t_SL g147 ( 
.A(n_127),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_115),
.A2(n_124),
.B1(n_122),
.B2(n_106),
.Y(n_148)
);

BUFx5_ASAP7_75t_L g149 ( 
.A(n_123),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_149),
.B(n_157),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_124),
.A2(n_22),
.B1(n_28),
.B2(n_24),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_L g169 ( 
.A1(n_151),
.A2(n_116),
.B(n_111),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_133),
.Y(n_152)
);

INVx4_ASAP7_75t_L g196 ( 
.A(n_152),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_127),
.B(n_35),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_SL g185 ( 
.A(n_154),
.B(n_155),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_106),
.B(n_35),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_SL g156 ( 
.A1(n_124),
.A2(n_88),
.B1(n_93),
.B2(n_100),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_122),
.Y(n_157)
);

INVx4_ASAP7_75t_L g158 ( 
.A(n_123),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_158),
.B(n_160),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_159),
.B(n_163),
.Y(n_187)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_126),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_L g161 ( 
.A1(n_107),
.A2(n_0),
.B(n_1),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_124),
.A2(n_84),
.B1(n_24),
.B2(n_20),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_162),
.A2(n_114),
.B1(n_109),
.B2(n_125),
.Y(n_182)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_107),
.Y(n_163)
);

CKINVDCx16_ASAP7_75t_R g164 ( 
.A(n_130),
.Y(n_164)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_164),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_112),
.B(n_104),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_165),
.B(n_166),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_112),
.B(n_29),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_SL g215 ( 
.A1(n_167),
.A2(n_176),
.B(n_181),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_L g208 ( 
.A1(n_169),
.A2(n_192),
.B(n_26),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_170),
.B(n_188),
.C(n_190),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_141),
.A2(n_129),
.B1(n_108),
.B2(n_125),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_171),
.A2(n_174),
.B1(n_103),
.B2(n_26),
.Y(n_201)
);

AO21x2_ASAP7_75t_L g174 ( 
.A1(n_153),
.A2(n_117),
.B(n_119),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_148),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_175),
.B(n_179),
.Y(n_206)
);

AOI21xp5_ASAP7_75t_SL g176 ( 
.A1(n_151),
.A2(n_109),
.B(n_28),
.Y(n_176)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_159),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_162),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_180),
.B(n_184),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_137),
.A2(n_131),
.B1(n_114),
.B2(n_28),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_182),
.A2(n_189),
.B1(n_199),
.B2(n_34),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_SL g183 ( 
.A1(n_163),
.A2(n_113),
.B(n_134),
.Y(n_183)
);

AOI21xp5_ASAP7_75t_L g226 ( 
.A1(n_183),
.A2(n_1),
.B(n_2),
.Y(n_226)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_165),
.Y(n_184)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_153),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_186),
.B(n_194),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_140),
.B(n_146),
.C(n_166),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_143),
.A2(n_108),
.B1(n_129),
.B2(n_113),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_161),
.B(n_144),
.C(n_150),
.Y(n_190)
);

BUFx2_ASAP7_75t_L g191 ( 
.A(n_152),
.Y(n_191)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_191),
.Y(n_202)
);

AOI21xp5_ASAP7_75t_SL g192 ( 
.A1(n_136),
.A2(n_142),
.B(n_120),
.Y(n_192)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_145),
.Y(n_194)
);

CKINVDCx16_ASAP7_75t_R g198 ( 
.A(n_149),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_198),
.B(n_183),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_158),
.A2(n_34),
.B1(n_32),
.B2(n_103),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_201),
.A2(n_174),
.B1(n_199),
.B2(n_186),
.Y(n_235)
);

INVx4_ASAP7_75t_L g203 ( 
.A(n_191),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_203),
.B(n_204),
.Y(n_234)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_182),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_193),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_205),
.B(n_207),
.Y(n_246)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_168),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_L g239 ( 
.A1(n_208),
.A2(n_220),
.B(n_226),
.Y(n_239)
);

CKINVDCx16_ASAP7_75t_R g209 ( 
.A(n_200),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_209),
.B(n_214),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_195),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_SL g243 ( 
.A1(n_210),
.A2(n_216),
.B(n_224),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_180),
.A2(n_32),
.B1(n_34),
.B2(n_26),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_211),
.A2(n_221),
.B1(n_225),
.B2(n_230),
.Y(n_251)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_189),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_192),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_SL g218 ( 
.A(n_176),
.B(n_169),
.Y(n_218)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_218),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_170),
.B(n_32),
.C(n_34),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_219),
.B(n_171),
.C(n_174),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_L g220 ( 
.A1(n_177),
.A2(n_26),
.B(n_2),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_185),
.B(n_173),
.Y(n_222)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_222),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_188),
.B(n_26),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_223),
.B(n_196),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_194),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_175),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_196),
.B(n_15),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_227),
.A2(n_229),
.B1(n_15),
.B2(n_14),
.Y(n_254)
);

AND2x2_ASAP7_75t_L g228 ( 
.A(n_174),
.B(n_3),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_L g248 ( 
.A1(n_228),
.A2(n_177),
.B(n_174),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_172),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_212),
.B(n_172),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_231),
.B(n_232),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_212),
.B(n_181),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_235),
.B(n_254),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_236),
.B(n_240),
.C(n_242),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_223),
.B(n_219),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_238),
.B(n_245),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_206),
.B(n_184),
.C(n_197),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_206),
.B(n_197),
.C(n_187),
.Y(n_242)
);

INVx1_ASAP7_75t_SL g244 ( 
.A(n_217),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_244),
.B(n_217),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_208),
.B(n_190),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_213),
.B(n_215),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_247),
.B(n_252),
.C(n_214),
.Y(n_271)
);

AOI21xp5_ASAP7_75t_L g269 ( 
.A1(n_248),
.A2(n_228),
.B(n_220),
.Y(n_269)
);

MAJx2_ASAP7_75t_L g249 ( 
.A(n_215),
.B(n_187),
.C(n_179),
.Y(n_249)
);

XNOR2x1_ASAP7_75t_L g261 ( 
.A(n_249),
.B(n_250),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_SL g250 ( 
.A(n_213),
.B(n_178),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_221),
.A2(n_9),
.B1(n_14),
.B2(n_13),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_253),
.A2(n_226),
.B1(n_210),
.B2(n_204),
.Y(n_272)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_246),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_257),
.B(n_258),
.Y(n_290)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_243),
.Y(n_258)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_234),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_262),
.B(n_264),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_241),
.B(n_209),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_SL g282 ( 
.A(n_263),
.B(n_265),
.Y(n_282)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_237),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_SL g265 ( 
.A(n_233),
.B(n_207),
.Y(n_265)
);

AND2x2_ASAP7_75t_L g266 ( 
.A(n_244),
.B(n_216),
.Y(n_266)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_266),
.Y(n_287)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_240),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_267),
.B(n_268),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_SL g268 ( 
.A(n_232),
.B(n_205),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_SL g276 ( 
.A1(n_269),
.A2(n_273),
.B(n_274),
.Y(n_276)
);

INVxp67_ASAP7_75t_L g270 ( 
.A(n_236),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_270),
.A2(n_272),
.B1(n_275),
.B2(n_248),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_271),
.B(n_252),
.Y(n_279)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_242),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_247),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_256),
.B(n_231),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_277),
.B(n_285),
.Y(n_301)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_278),
.Y(n_303)
);

XOR2xp5_ASAP7_75t_L g299 ( 
.A(n_279),
.B(n_281),
.Y(n_299)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_255),
.B(n_245),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_270),
.A2(n_230),
.B1(n_228),
.B2(n_218),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_L g295 ( 
.A1(n_283),
.A2(n_269),
.B1(n_261),
.B2(n_275),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_259),
.B(n_238),
.C(n_249),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_284),
.B(n_286),
.C(n_261),
.Y(n_297)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_255),
.B(n_250),
.Y(n_285)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_259),
.B(n_239),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_L g289 ( 
.A1(n_260),
.A2(n_251),
.B1(n_201),
.B2(n_239),
.Y(n_289)
);

INVxp67_ASAP7_75t_L g296 ( 
.A(n_289),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_256),
.B(n_225),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_291),
.B(n_292),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_271),
.B(n_211),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_282),
.B(n_264),
.Y(n_293)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_293),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_295),
.A2(n_292),
.B1(n_276),
.B2(n_286),
.Y(n_311)
);

XOR2xp5_ASAP7_75t_L g307 ( 
.A(n_297),
.B(n_279),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_SL g298 ( 
.A(n_288),
.B(n_272),
.Y(n_298)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_298),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_SL g300 ( 
.A(n_280),
.B(n_266),
.Y(n_300)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_300),
.Y(n_312)
);

OAI21xp5_ASAP7_75t_L g302 ( 
.A1(n_287),
.A2(n_266),
.B(n_224),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_SL g314 ( 
.A(n_302),
.B(n_306),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_L g304 ( 
.A1(n_290),
.A2(n_202),
.B1(n_203),
.B2(n_11),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_L g316 ( 
.A1(n_304),
.A2(n_15),
.B1(n_14),
.B2(n_13),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_SL g305 ( 
.A(n_291),
.B(n_202),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_305),
.B(n_306),
.Y(n_310)
);

AOI21xp5_ASAP7_75t_L g306 ( 
.A1(n_283),
.A2(n_4),
.B(n_5),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_307),
.B(n_313),
.C(n_315),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_311),
.B(n_296),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_303),
.B(n_284),
.C(n_277),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g318 ( 
.A(n_314),
.B(n_302),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_294),
.B(n_281),
.C(n_285),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_316),
.B(n_11),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_SL g326 ( 
.A(n_318),
.B(n_320),
.Y(n_326)
);

OAI21xp5_ASAP7_75t_SL g319 ( 
.A1(n_308),
.A2(n_296),
.B(n_297),
.Y(n_319)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_319),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_SL g321 ( 
.A(n_309),
.B(n_301),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_321),
.B(n_322),
.Y(n_327)
);

AOI21xp5_ASAP7_75t_L g322 ( 
.A1(n_311),
.A2(n_301),
.B(n_299),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_323),
.B(n_324),
.Y(n_325)
);

OAI321xp33_ASAP7_75t_L g324 ( 
.A1(n_310),
.A2(n_314),
.A3(n_312),
.B1(n_313),
.B2(n_315),
.C(n_307),
.Y(n_324)
);

BUFx24_ASAP7_75t_SL g328 ( 
.A(n_321),
.Y(n_328)
);

OA21x2_ASAP7_75t_L g331 ( 
.A1(n_328),
.A2(n_317),
.B(n_299),
.Y(n_331)
);

OAI21xp5_ASAP7_75t_L g330 ( 
.A1(n_325),
.A2(n_329),
.B(n_326),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_330),
.B(n_331),
.Y(n_332)
);

AOI21xp5_ASAP7_75t_L g333 ( 
.A1(n_332),
.A2(n_327),
.B(n_5),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_333),
.Y(n_334)
);

AOI21xp5_ASAP7_75t_L g335 ( 
.A1(n_334),
.A2(n_4),
.B(n_6),
.Y(n_335)
);

XNOR2xp5_ASAP7_75t_L g336 ( 
.A(n_335),
.B(n_4),
.Y(n_336)
);

AOI21xp5_ASAP7_75t_L g337 ( 
.A1(n_336),
.A2(n_8),
.B(n_6),
.Y(n_337)
);


endmodule