module real_jpeg_25757_n_6 (n_5, n_4, n_0, n_1, n_2, n_3, n_6);

input n_5;
input n_4;
input n_0;
input n_1;
input n_2;
input n_3;

output n_6;

wire n_17;
wire n_8;
wire n_37;
wire n_21;
wire n_38;
wire n_33;
wire n_35;
wire n_29;
wire n_10;
wire n_31;
wire n_9;
wire n_12;
wire n_24;
wire n_34;
wire n_28;
wire n_23;
wire n_11;
wire n_14;
wire n_25;
wire n_7;
wire n_22;
wire n_18;
wire n_36;
wire n_27;
wire n_26;
wire n_20;
wire n_19;
wire n_32;
wire n_30;
wire n_16;
wire n_15;
wire n_13;

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_0),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_1),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g9 ( 
.A(n_2),
.Y(n_9)
);

AND2x2_ASAP7_75t_L g34 ( 
.A(n_2),
.B(n_4),
.Y(n_34)
);

AND2x2_ASAP7_75t_L g15 ( 
.A(n_3),
.B(n_16),
.Y(n_15)
);

OR2x2_ASAP7_75t_SL g20 ( 
.A(n_3),
.B(n_16),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_3),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_4),
.B(n_15),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_4),
.B(n_5),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_4),
.B(n_22),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_4),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_5),
.Y(n_11)
);

AOI221xp5_ASAP7_75t_L g6 ( 
.A1(n_7),
.A2(n_18),
.B1(n_19),
.B2(n_23),
.C(n_28),
.Y(n_6)
);

OAI21xp33_ASAP7_75t_SL g7 ( 
.A1(n_8),
.A2(n_14),
.B(n_17),
.Y(n_7)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_8),
.B(n_27),
.Y(n_35)
);

AOI21xp5_ASAP7_75t_SL g8 ( 
.A1(n_9),
.A2(n_10),
.B(n_13),
.Y(n_8)
);

NAND2xp5_ASAP7_75t_SL g25 ( 
.A(n_9),
.B(n_10),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_9),
.B(n_27),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g10 ( 
.A(n_11),
.B(n_12),
.Y(n_10)
);

NOR2xp33_ASAP7_75t_L g13 ( 
.A(n_11),
.B(n_12),
.Y(n_13)
);

OAI21xp33_ASAP7_75t_SL g19 ( 
.A1(n_11),
.A2(n_20),
.B(n_21),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_13),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_15),
.Y(n_14)
);

AND2x2_ASAP7_75t_SL g30 ( 
.A(n_16),
.B(n_31),
.Y(n_30)
);

OR2x2_ASAP7_75t_L g36 ( 
.A(n_16),
.B(n_31),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_20),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_SL g37 ( 
.A(n_23),
.B(n_38),
.Y(n_37)
);

INVx1_ASAP7_75t_SL g23 ( 
.A(n_24),
.Y(n_23)
);

AOI21xp5_ASAP7_75t_SL g24 ( 
.A1(n_25),
.A2(n_26),
.B(n_27),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_L g28 ( 
.A1(n_29),
.A2(n_32),
.B1(n_36),
.B2(n_37),
.Y(n_28)
);

INVx1_ASAP7_75t_SL g29 ( 
.A(n_30),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_33),
.B(n_35),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_34),
.Y(n_33)
);


endmodule