module fake_jpeg_30724_n_265 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_265);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_265;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_182;
wire n_19;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_122;
wire n_75;
wire n_246;
wire n_37;
wire n_233;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_165;
wire n_78;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_140;
wire n_82;
wire n_155;
wire n_100;
wire n_258;
wire n_96;

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_6),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_0),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_2),
.Y(n_23)
);

INVx11_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_10),
.Y(n_26)
);

INVxp67_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_6),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_17),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

BUFx4f_ASAP7_75t_SL g31 ( 
.A(n_5),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

INVx13_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_3),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_13),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_1),
.Y(n_37)
);

INVx2_ASAP7_75t_SL g38 ( 
.A(n_8),
.Y(n_38)
);

INVx5_ASAP7_75t_L g39 ( 
.A(n_14),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_5),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_1),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_35),
.Y(n_42)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_42),
.Y(n_92)
);

BUFx12_ASAP7_75t_L g43 ( 
.A(n_39),
.Y(n_43)
);

INVx13_ASAP7_75t_L g71 ( 
.A(n_43),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_26),
.B(n_17),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_44),
.B(n_47),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_L g45 ( 
.A1(n_34),
.A2(n_37),
.B1(n_36),
.B2(n_18),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_45),
.A2(n_21),
.B1(n_25),
.B2(n_32),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_24),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_46),
.Y(n_94)
);

CKINVDCx16_ASAP7_75t_R g47 ( 
.A(n_31),
.Y(n_47)
);

OR2x2_ASAP7_75t_L g48 ( 
.A(n_18),
.B(n_0),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_48),
.B(n_49),
.Y(n_103)
);

BUFx12_ASAP7_75t_L g49 ( 
.A(n_39),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_20),
.Y(n_50)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_50),
.Y(n_70)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_20),
.Y(n_51)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_51),
.Y(n_84)
);

OR2x2_ASAP7_75t_L g52 ( 
.A(n_23),
.B(n_2),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_52),
.B(n_55),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_24),
.Y(n_53)
);

INVx6_ASAP7_75t_L g102 ( 
.A(n_53),
.Y(n_102)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_21),
.Y(n_54)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_54),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_19),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_19),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_56),
.B(n_27),
.Y(n_89)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_35),
.Y(n_57)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_57),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_26),
.B(n_9),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_58),
.B(n_63),
.Y(n_78)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_30),
.Y(n_59)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_59),
.Y(n_95)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_21),
.Y(n_60)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_60),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_38),
.B(n_3),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_61),
.B(n_68),
.Y(n_72)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_34),
.Y(n_62)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_62),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_22),
.B(n_9),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_33),
.Y(n_64)
);

INVx1_ASAP7_75t_SL g86 ( 
.A(n_64),
.Y(n_86)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_33),
.Y(n_65)
);

INVx5_ASAP7_75t_L g107 ( 
.A(n_65),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_37),
.Y(n_66)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_66),
.Y(n_83)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_30),
.Y(n_67)
);

CKINVDCx16_ASAP7_75t_R g73 ( 
.A(n_67),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_29),
.B(n_10),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_38),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_69),
.A2(n_23),
.B1(n_40),
.B2(n_28),
.Y(n_82)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_65),
.Y(n_76)
);

INVx1_ASAP7_75t_SL g132 ( 
.A(n_76),
.Y(n_132)
);

HB1xp67_ASAP7_75t_L g77 ( 
.A(n_42),
.Y(n_77)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_77),
.Y(n_139)
);

AO22x1_ASAP7_75t_SL g80 ( 
.A1(n_62),
.A2(n_36),
.B1(n_31),
.B2(n_38),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_80),
.A2(n_85),
.B1(n_90),
.B2(n_93),
.Y(n_125)
);

CKINVDCx12_ASAP7_75t_R g81 ( 
.A(n_64),
.Y(n_81)
);

INVxp67_ASAP7_75t_SL g110 ( 
.A(n_81),
.Y(n_110)
);

OR2x2_ASAP7_75t_L g121 ( 
.A(n_82),
.B(n_87),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_L g85 ( 
.A1(n_66),
.A2(n_41),
.B1(n_40),
.B2(n_28),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_50),
.A2(n_27),
.B1(n_41),
.B2(n_29),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_61),
.B(n_32),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_88),
.B(n_97),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_89),
.B(n_91),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_48),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_57),
.A2(n_21),
.B1(n_25),
.B2(n_64),
.Y(n_93)
);

BUFx3_ASAP7_75t_L g96 ( 
.A(n_54),
.Y(n_96)
);

INVx4_ASAP7_75t_L g130 ( 
.A(n_96),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_52),
.B(n_25),
.Y(n_97)
);

CKINVDCx16_ASAP7_75t_R g99 ( 
.A(n_51),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_99),
.B(n_11),
.Y(n_126)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_60),
.Y(n_101)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_101),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_59),
.B(n_25),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_104),
.B(n_16),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_67),
.A2(n_4),
.B1(n_7),
.B2(n_8),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_105),
.A2(n_16),
.B1(n_11),
.B2(n_15),
.Y(n_127)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_70),
.Y(n_108)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_108),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_96),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_109),
.B(n_112),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_72),
.B(n_31),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_111),
.B(n_115),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_76),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_84),
.A2(n_46),
.B1(n_53),
.B2(n_49),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_SL g165 ( 
.A1(n_113),
.A2(n_136),
.B(n_132),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_87),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g145 ( 
.A(n_114),
.B(n_126),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_95),
.B(n_73),
.Y(n_115)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_106),
.Y(n_117)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_117),
.Y(n_142)
);

AND2x4_ASAP7_75t_L g118 ( 
.A(n_80),
.B(n_49),
.Y(n_118)
);

AND2x2_ASAP7_75t_L g147 ( 
.A(n_118),
.B(n_122),
.Y(n_147)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_92),
.Y(n_119)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_119),
.Y(n_161)
);

BUFx2_ASAP7_75t_L g120 ( 
.A(n_101),
.Y(n_120)
);

INVx3_ASAP7_75t_L g151 ( 
.A(n_120),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_L g122 ( 
.A(n_103),
.B(n_43),
.Y(n_122)
);

OAI22xp33_ASAP7_75t_L g123 ( 
.A1(n_83),
.A2(n_43),
.B1(n_4),
.B2(n_13),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_123),
.A2(n_127),
.B1(n_135),
.B2(n_138),
.Y(n_158)
);

CKINVDCx16_ASAP7_75t_R g124 ( 
.A(n_93),
.Y(n_124)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_124),
.Y(n_148)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_92),
.Y(n_129)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_129),
.Y(n_152)
);

BUFx2_ASAP7_75t_L g131 ( 
.A(n_74),
.Y(n_131)
);

INVx3_ASAP7_75t_L g162 ( 
.A(n_131),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_94),
.Y(n_133)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_133),
.Y(n_153)
);

CKINVDCx16_ASAP7_75t_R g134 ( 
.A(n_86),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_134),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g136 ( 
.A(n_86),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_136),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_75),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g146 ( 
.A(n_137),
.B(n_140),
.Y(n_146)
);

OR2x4_ASAP7_75t_L g138 ( 
.A(n_80),
.B(n_15),
.Y(n_138)
);

OR2x4_ASAP7_75t_L g164 ( 
.A(n_138),
.B(n_123),
.Y(n_164)
);

OA21x2_ASAP7_75t_L g143 ( 
.A1(n_121),
.A2(n_90),
.B(n_105),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_SL g175 ( 
.A1(n_143),
.A2(n_164),
.B(n_155),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_L g149 ( 
.A1(n_125),
.A2(n_83),
.B1(n_102),
.B2(n_94),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_149),
.A2(n_163),
.B1(n_166),
.B2(n_164),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_121),
.A2(n_98),
.B1(n_79),
.B2(n_102),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_150),
.A2(n_157),
.B1(n_158),
.B2(n_160),
.Y(n_170)
);

AOI21xp5_ASAP7_75t_L g154 ( 
.A1(n_118),
.A2(n_107),
.B(n_74),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_L g172 ( 
.A1(n_154),
.A2(n_165),
.B(n_157),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_115),
.B(n_98),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_156),
.B(n_133),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_118),
.A2(n_100),
.B1(n_107),
.B2(n_71),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_118),
.A2(n_100),
.B1(n_71),
.B2(n_78),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_111),
.A2(n_108),
.B1(n_122),
.B2(n_116),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_117),
.A2(n_129),
.B1(n_139),
.B2(n_119),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_SL g168 ( 
.A(n_145),
.B(n_128),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_168),
.B(n_178),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_146),
.B(n_110),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_169),
.B(n_183),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_147),
.B(n_163),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_171),
.B(n_175),
.C(n_186),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_SL g203 ( 
.A1(n_172),
.A2(n_190),
.B(n_170),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_159),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_173),
.Y(n_194)
);

AND2x4_ASAP7_75t_SL g174 ( 
.A(n_154),
.B(n_128),
.Y(n_174)
);

AND2x2_ASAP7_75t_L g192 ( 
.A(n_174),
.B(n_180),
.Y(n_192)
);

AO22x1_ASAP7_75t_L g197 ( 
.A1(n_175),
.A2(n_151),
.B1(n_166),
.B2(n_189),
.Y(n_197)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_141),
.Y(n_176)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_176),
.Y(n_208)
);

INVx3_ASAP7_75t_L g177 ( 
.A(n_162),
.Y(n_177)
);

HB1xp67_ASAP7_75t_L g205 ( 
.A(n_177),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_SL g178 ( 
.A(n_155),
.B(n_130),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_141),
.Y(n_179)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_179),
.Y(n_200)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_142),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_142),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_181),
.B(n_182),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_156),
.B(n_131),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_150),
.B(n_120),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_SL g184 ( 
.A(n_158),
.B(n_130),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_184),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_185),
.B(n_186),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_147),
.B(n_132),
.Y(n_186)
);

AOI22xp33_ASAP7_75t_SL g187 ( 
.A1(n_148),
.A2(n_167),
.B1(n_165),
.B2(n_144),
.Y(n_187)
);

AOI22xp33_ASAP7_75t_SL g196 ( 
.A1(n_187),
.A2(n_153),
.B1(n_151),
.B2(n_161),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_160),
.B(n_152),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_188),
.A2(n_189),
.B1(n_190),
.B2(n_172),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_147),
.B(n_143),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_143),
.B(n_152),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_191),
.A2(n_153),
.B1(n_162),
.B2(n_161),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_193),
.A2(n_196),
.B1(n_177),
.B2(n_197),
.Y(n_225)
);

A2O1A1O1Ixp25_ASAP7_75t_L g211 ( 
.A1(n_197),
.A2(n_174),
.B(n_185),
.C(n_176),
.D(n_179),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_201),
.B(n_173),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_202),
.B(n_209),
.Y(n_220)
);

AOI21xp5_ASAP7_75t_L g221 ( 
.A1(n_203),
.A2(n_204),
.B(n_210),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_SL g204 ( 
.A1(n_184),
.A2(n_174),
.B(n_170),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_171),
.B(n_178),
.C(n_191),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_L g210 ( 
.A1(n_174),
.A2(n_182),
.B(n_168),
.Y(n_210)
);

OA21x2_ASAP7_75t_L g230 ( 
.A1(n_211),
.A2(n_204),
.B(n_192),
.Y(n_230)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_200),
.Y(n_212)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_212),
.Y(n_227)
);

CKINVDCx14_ASAP7_75t_R g213 ( 
.A(n_198),
.Y(n_213)
);

INVx13_ASAP7_75t_L g236 ( 
.A(n_213),
.Y(n_236)
);

XOR2x1_ASAP7_75t_L g214 ( 
.A(n_197),
.B(n_210),
.Y(n_214)
);

BUFx12f_ASAP7_75t_SL g234 ( 
.A(n_214),
.Y(n_234)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_200),
.Y(n_215)
);

INVxp67_ASAP7_75t_L g233 ( 
.A(n_215),
.Y(n_233)
);

CKINVDCx16_ASAP7_75t_R g216 ( 
.A(n_208),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_SL g232 ( 
.A(n_216),
.B(n_217),
.Y(n_232)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_199),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_218),
.B(n_219),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_198),
.B(n_180),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_202),
.B(n_181),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_222),
.B(n_207),
.C(n_203),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_199),
.Y(n_223)
);

BUFx12_ASAP7_75t_L g226 ( 
.A(n_223),
.Y(n_226)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_205),
.Y(n_224)
);

AOI21xp5_ASAP7_75t_L g235 ( 
.A1(n_224),
.A2(n_225),
.B(n_193),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_220),
.B(n_209),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_228),
.B(n_231),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_230),
.B(n_221),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_235),
.B(n_221),
.Y(n_243)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_232),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_238),
.A2(n_243),
.B1(n_245),
.B2(n_229),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_228),
.B(n_222),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_239),
.B(n_207),
.Y(n_249)
);

INVxp33_ASAP7_75t_SL g240 ( 
.A(n_234),
.Y(n_240)
);

XNOR2x1_ASAP7_75t_L g248 ( 
.A(n_240),
.B(n_242),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_231),
.B(n_220),
.C(n_218),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_SL g247 ( 
.A(n_241),
.B(n_244),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_SL g244 ( 
.A1(n_234),
.A2(n_219),
.B(n_206),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_229),
.B(n_194),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_246),
.B(n_249),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_237),
.B(n_211),
.Y(n_250)
);

OA21x2_ASAP7_75t_SL g253 ( 
.A1(n_250),
.A2(n_230),
.B(n_237),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_240),
.A2(n_235),
.B1(n_195),
.B2(n_227),
.Y(n_251)
);

A2O1A1Ixp33_ASAP7_75t_SL g256 ( 
.A1(n_251),
.A2(n_252),
.B(n_192),
.C(n_236),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_241),
.A2(n_192),
.B1(n_214),
.B2(n_230),
.Y(n_252)
);

AOI21x1_ASAP7_75t_L g259 ( 
.A1(n_253),
.A2(n_254),
.B(n_256),
.Y(n_259)
);

OAI21xp33_ASAP7_75t_L g254 ( 
.A1(n_247),
.A2(n_226),
.B(n_236),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_SL g257 ( 
.A1(n_248),
.A2(n_233),
.B(n_227),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_257),
.B(n_226),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_258),
.B(n_260),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_255),
.B(n_250),
.C(n_248),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_259),
.A2(n_233),
.B1(n_215),
.B2(n_212),
.Y(n_262)
);

AO21x1_ASAP7_75t_L g263 ( 
.A1(n_262),
.A2(n_226),
.B(n_224),
.Y(n_263)
);

AOI21xp5_ASAP7_75t_SL g264 ( 
.A1(n_263),
.A2(n_261),
.B(n_252),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_264),
.B(n_249),
.Y(n_265)
);


endmodule