module fake_jpeg_26755_n_324 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_324);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_324;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_14),
.Y(n_19)
);

BUFx24_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_2),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_13),
.Y(n_28)
);

INVx11_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_20),
.Y(n_35)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_29),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_36),
.Y(n_59)
);

BUFx4f_ASAP7_75t_SL g37 ( 
.A(n_20),
.Y(n_37)
);

INVx2_ASAP7_75t_SL g52 ( 
.A(n_37),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_20),
.Y(n_38)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_20),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_39),
.B(n_41),
.Y(n_45)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

INVx2_ASAP7_75t_SL g65 ( 
.A(n_40),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g41 ( 
.A(n_19),
.B(n_8),
.Y(n_41)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_29),
.Y(n_42)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_42),
.Y(n_47)
);

CKINVDCx12_ASAP7_75t_R g43 ( 
.A(n_30),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_43),
.B(n_30),
.Y(n_56)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_20),
.Y(n_44)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_44),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g48 ( 
.A1(n_40),
.A2(n_18),
.B1(n_25),
.B2(n_34),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_48),
.A2(n_68),
.B1(n_44),
.B2(n_34),
.Y(n_71)
);

OA22x2_ASAP7_75t_L g49 ( 
.A1(n_44),
.A2(n_20),
.B1(n_27),
.B2(n_30),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_49),
.B(n_35),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_41),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_51),
.B(n_61),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_41),
.B(n_18),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_53),
.B(n_57),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_43),
.A2(n_19),
.B1(n_28),
.B2(n_44),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_54),
.A2(n_64),
.B1(n_25),
.B2(n_17),
.Y(n_78)
);

OR2x2_ASAP7_75t_L g94 ( 
.A(n_56),
.B(n_63),
.Y(n_94)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_58),
.Y(n_81)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_36),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_60),
.B(n_67),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_39),
.B(n_19),
.Y(n_61)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_36),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_62),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_39),
.B(n_28),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_43),
.A2(n_27),
.B1(n_33),
.B2(n_32),
.Y(n_64)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_36),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_66),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_39),
.B(n_17),
.Y(n_67)
);

O2A1O1Ixp33_ASAP7_75t_L g68 ( 
.A1(n_44),
.A2(n_34),
.B(n_18),
.C(n_25),
.Y(n_68)
);

INVx3_ASAP7_75t_SL g70 ( 
.A(n_59),
.Y(n_70)
);

OA22x2_ASAP7_75t_L g95 ( 
.A1(n_70),
.A2(n_46),
.B1(n_55),
.B2(n_65),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_71),
.B(n_78),
.Y(n_96)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_68),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_73),
.B(n_83),
.Y(n_117)
);

HB1xp67_ASAP7_75t_L g74 ( 
.A(n_65),
.Y(n_74)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_74),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_56),
.B(n_37),
.C(n_44),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_75),
.B(n_37),
.C(n_35),
.Y(n_118)
);

INVx1_ASAP7_75t_SL g104 ( 
.A(n_76),
.Y(n_104)
);

INVx5_ASAP7_75t_L g77 ( 
.A(n_62),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_77),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_45),
.B(n_21),
.Y(n_80)
);

A2O1A1Ixp33_ASAP7_75t_L g105 ( 
.A1(n_80),
.A2(n_49),
.B(n_37),
.C(n_50),
.Y(n_105)
);

HB1xp67_ASAP7_75t_L g82 ( 
.A(n_65),
.Y(n_82)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_82),
.Y(n_103)
);

NAND3xp33_ASAP7_75t_L g83 ( 
.A(n_53),
.B(n_8),
.C(n_15),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_45),
.B(n_22),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_85),
.B(n_90),
.Y(n_112)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_68),
.Y(n_86)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_86),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_63),
.B(n_21),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_88),
.B(n_92),
.Y(n_122)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_48),
.Y(n_89)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_89),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_51),
.B(n_22),
.Y(n_90)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_67),
.Y(n_91)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_91),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_57),
.B(n_17),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_61),
.B(n_23),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_93),
.Y(n_121)
);

CKINVDCx14_ASAP7_75t_R g128 ( 
.A(n_95),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_72),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_97),
.B(n_108),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_73),
.A2(n_47),
.B1(n_58),
.B2(n_55),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_98),
.A2(n_109),
.B1(n_52),
.B2(n_60),
.Y(n_143)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_72),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_100),
.B(n_115),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_86),
.A2(n_47),
.B1(n_49),
.B2(n_42),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_101),
.A2(n_110),
.B1(n_120),
.B2(n_52),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_L g134 ( 
.A1(n_105),
.A2(n_111),
.B(n_113),
.Y(n_134)
);

INVx8_ASAP7_75t_L g107 ( 
.A(n_72),
.Y(n_107)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_107),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_87),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_76),
.A2(n_55),
.B1(n_46),
.B2(n_50),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_89),
.A2(n_49),
.B1(n_40),
.B2(n_42),
.Y(n_110)
);

AND2x2_ASAP7_75t_L g111 ( 
.A(n_90),
.B(n_49),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g113 ( 
.A(n_85),
.B(n_35),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_91),
.A2(n_52),
.B1(n_46),
.B2(n_23),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_114),
.A2(n_37),
.B1(n_35),
.B2(n_38),
.Y(n_151)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_81),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_118),
.B(n_75),
.C(n_37),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_71),
.A2(n_78),
.B1(n_76),
.B2(n_69),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_123),
.B(n_135),
.C(n_137),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_124),
.A2(n_151),
.B1(n_97),
.B2(n_108),
.Y(n_162)
);

XOR2xp5_ASAP7_75t_L g126 ( 
.A(n_120),
.B(n_69),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_126),
.B(n_130),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_96),
.A2(n_80),
.B1(n_84),
.B2(n_70),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_129),
.A2(n_135),
.B1(n_104),
.B2(n_124),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_SL g130 ( 
.A(n_112),
.B(n_79),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_106),
.A2(n_84),
.B1(n_79),
.B2(n_70),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_131),
.A2(n_143),
.B1(n_145),
.B2(n_146),
.Y(n_155)
);

CKINVDCx16_ASAP7_75t_R g133 ( 
.A(n_98),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_133),
.B(n_136),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_118),
.B(n_80),
.C(n_94),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_107),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_104),
.B(n_112),
.C(n_96),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_95),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_138),
.B(n_142),
.Y(n_157)
);

INVx5_ASAP7_75t_L g139 ( 
.A(n_99),
.Y(n_139)
);

CKINVDCx14_ASAP7_75t_R g166 ( 
.A(n_139),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_119),
.B(n_94),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g160 ( 
.A(n_140),
.B(n_141),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_119),
.B(n_94),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_95),
.Y(n_142)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_95),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_144),
.B(n_147),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_106),
.A2(n_77),
.B1(n_81),
.B2(n_40),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_116),
.A2(n_42),
.B1(n_66),
.B2(n_36),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_109),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_111),
.B(n_87),
.Y(n_148)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_148),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_116),
.A2(n_42),
.B1(n_36),
.B2(n_37),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_149),
.A2(n_110),
.B1(n_100),
.B2(n_101),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_121),
.B(n_87),
.Y(n_150)
);

OAI21xp33_ASAP7_75t_L g178 ( 
.A1(n_150),
.A2(n_23),
.B(n_26),
.Y(n_178)
);

CKINVDCx16_ASAP7_75t_R g153 ( 
.A(n_125),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_153),
.B(n_154),
.Y(n_206)
);

CKINVDCx16_ASAP7_75t_R g156 ( 
.A(n_125),
.Y(n_156)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_156),
.Y(n_187)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_127),
.Y(n_158)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_158),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_159),
.A2(n_176),
.B1(n_182),
.B2(n_136),
.Y(n_191)
);

CKINVDCx16_ASAP7_75t_R g161 ( 
.A(n_145),
.Y(n_161)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_161),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_SL g196 ( 
.A1(n_162),
.A2(n_168),
.B(n_170),
.Y(n_196)
);

AO21x2_ASAP7_75t_L g164 ( 
.A1(n_128),
.A2(n_96),
.B(n_105),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_164),
.A2(n_167),
.B1(n_38),
.B2(n_26),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_147),
.A2(n_111),
.B1(n_113),
.B2(n_117),
.Y(n_167)
);

AOI21xp5_ASAP7_75t_L g168 ( 
.A1(n_134),
.A2(n_113),
.B(n_102),
.Y(n_168)
);

OA21x2_ASAP7_75t_L g169 ( 
.A1(n_138),
.A2(n_103),
.B(n_102),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_L g203 ( 
.A1(n_169),
.A2(n_38),
.B(n_31),
.Y(n_203)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_151),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_150),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_SL g183 ( 
.A(n_171),
.B(n_131),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_126),
.B(n_121),
.C(n_103),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_173),
.B(n_177),
.C(n_134),
.Y(n_184)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_146),
.Y(n_174)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_174),
.Y(n_204)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_148),
.Y(n_175)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_175),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_142),
.A2(n_115),
.B1(n_99),
.B2(n_122),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_123),
.B(n_37),
.C(n_59),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_SL g198 ( 
.A1(n_178),
.A2(n_33),
.B(n_32),
.Y(n_198)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_149),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_179),
.B(n_132),
.Y(n_194)
);

INVx3_ASAP7_75t_L g180 ( 
.A(n_139),
.Y(n_180)
);

INVx1_ASAP7_75t_SL g199 ( 
.A(n_180),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_144),
.A2(n_32),
.B1(n_26),
.B2(n_33),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_183),
.B(n_198),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_184),
.B(n_188),
.C(n_193),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_165),
.B(n_137),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_185),
.B(n_186),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_165),
.B(n_130),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_172),
.B(n_129),
.C(n_143),
.Y(n_188)
);

FAx1_ASAP7_75t_L g189 ( 
.A(n_164),
.B(n_133),
.CI(n_35),
.CON(n_189),
.SN(n_189)
);

OAI21xp5_ASAP7_75t_SL g222 ( 
.A1(n_189),
.A2(n_191),
.B(n_200),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_172),
.B(n_132),
.C(n_59),
.Y(n_193)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_194),
.Y(n_219)
);

OAI22x1_ASAP7_75t_L g195 ( 
.A1(n_164),
.A2(n_38),
.B1(n_24),
.B2(n_22),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_195),
.A2(n_180),
.B1(n_181),
.B2(n_166),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_163),
.B(n_21),
.Y(n_197)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_197),
.Y(n_224)
);

NAND2x1_ASAP7_75t_L g200 ( 
.A(n_170),
.B(n_38),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_201),
.A2(n_182),
.B1(n_152),
.B2(n_159),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_173),
.B(n_31),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_202),
.B(n_31),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_L g210 ( 
.A1(n_203),
.A2(n_208),
.B(n_209),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_154),
.B(n_24),
.C(n_22),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_205),
.B(n_169),
.C(n_24),
.Y(n_229)
);

OAI21xp5_ASAP7_75t_L g208 ( 
.A1(n_164),
.A2(n_0),
.B(n_1),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_L g209 ( 
.A1(n_164),
.A2(n_0),
.B(n_1),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_194),
.B(n_163),
.Y(n_211)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_211),
.Y(n_240)
);

NAND3xp33_ASAP7_75t_L g212 ( 
.A(n_190),
.B(n_160),
.C(n_200),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_212),
.B(n_229),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_214),
.A2(n_218),
.B1(n_227),
.B2(n_228),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_197),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_215),
.B(n_223),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_207),
.B(n_157),
.Y(n_216)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_216),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_187),
.B(n_176),
.Y(n_217)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_217),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_192),
.A2(n_157),
.B1(n_155),
.B2(n_179),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_204),
.B(n_152),
.Y(n_223)
);

CKINVDCx16_ASAP7_75t_R g236 ( 
.A(n_225),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_198),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_226),
.B(n_231),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_189),
.A2(n_155),
.B1(n_168),
.B2(n_167),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_209),
.A2(n_169),
.B1(n_177),
.B2(n_24),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_228),
.A2(n_195),
.B1(n_206),
.B2(n_200),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_230),
.B(n_202),
.Y(n_241)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_201),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_203),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_232),
.B(n_233),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_208),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_199),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_234),
.B(n_2),
.Y(n_256)
);

AOI21xp5_ASAP7_75t_L g235 ( 
.A1(n_196),
.A2(n_1),
.B(n_2),
.Y(n_235)
);

OAI21xp5_ASAP7_75t_L g257 ( 
.A1(n_235),
.A2(n_210),
.B(n_226),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_220),
.B(n_193),
.C(n_188),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_237),
.B(n_246),
.C(n_253),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_241),
.B(n_250),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_L g272 ( 
.A1(n_243),
.A2(n_247),
.B1(n_248),
.B2(n_249),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_220),
.B(n_184),
.C(n_185),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_231),
.A2(n_189),
.B1(n_196),
.B2(n_205),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_227),
.A2(n_199),
.B1(n_186),
.B2(n_10),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_SL g250 ( 
.A(n_221),
.B(n_9),
.Y(n_250)
);

A2O1A1Ixp33_ASAP7_75t_SL g252 ( 
.A1(n_233),
.A2(n_2),
.B(n_3),
.C(n_4),
.Y(n_252)
);

AOI21xp5_ASAP7_75t_L g262 ( 
.A1(n_252),
.A2(n_222),
.B(n_4),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_221),
.B(n_9),
.C(n_15),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_230),
.B(n_219),
.C(n_224),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_254),
.B(n_255),
.C(n_8),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_219),
.B(n_9),
.C(n_15),
.Y(n_255)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_256),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_L g261 ( 
.A1(n_257),
.A2(n_210),
.B(n_235),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_244),
.B(n_215),
.Y(n_260)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_260),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_261),
.A2(n_262),
.B1(n_263),
.B2(n_3),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_236),
.A2(n_218),
.B1(n_232),
.B2(n_224),
.Y(n_263)
);

AOI322xp5_ASAP7_75t_SL g264 ( 
.A1(n_250),
.A2(n_213),
.A3(n_216),
.B1(n_223),
.B2(n_225),
.C1(n_229),
.C2(n_222),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_264),
.B(n_266),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_238),
.B(n_234),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_265),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_255),
.B(n_211),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_267),
.B(n_274),
.C(n_252),
.Y(n_279)
);

HB1xp67_ASAP7_75t_L g269 ( 
.A(n_254),
.Y(n_269)
);

INVx11_ASAP7_75t_L g287 ( 
.A(n_269),
.Y(n_287)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_239),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_270),
.B(n_242),
.Y(n_278)
);

INVxp67_ASAP7_75t_L g271 ( 
.A(n_251),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_271),
.A2(n_248),
.B1(n_247),
.B2(n_252),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_241),
.B(n_10),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_273),
.B(n_253),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_237),
.B(n_10),
.C(n_12),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_SL g294 ( 
.A(n_275),
.B(n_273),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_278),
.B(n_283),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_SL g289 ( 
.A(n_279),
.B(n_274),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_258),
.B(n_246),
.C(n_245),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_280),
.B(n_285),
.C(n_288),
.Y(n_290)
);

XNOR2x1_ASAP7_75t_L g282 ( 
.A(n_261),
.B(n_257),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_282),
.B(n_272),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_263),
.B(n_240),
.Y(n_283)
);

INVxp67_ASAP7_75t_L g299 ( 
.A(n_284),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_258),
.B(n_252),
.C(n_11),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_286),
.A2(n_259),
.B1(n_4),
.B2(n_5),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_267),
.B(n_7),
.C(n_11),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_289),
.B(n_293),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_292),
.B(n_294),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_277),
.B(n_268),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_281),
.B(n_271),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_295),
.B(n_296),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_280),
.B(n_259),
.C(n_7),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_L g303 ( 
.A1(n_297),
.A2(n_284),
.B1(n_299),
.B2(n_288),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_276),
.B(n_7),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_298),
.B(n_12),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_282),
.B(n_12),
.C(n_16),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_300),
.B(n_275),
.C(n_286),
.Y(n_305)
);

AOI21x1_ASAP7_75t_L g302 ( 
.A1(n_299),
.A2(n_285),
.B(n_279),
.Y(n_302)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_302),
.Y(n_313)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_303),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_290),
.B(n_287),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_SL g311 ( 
.A(n_304),
.B(n_305),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_290),
.B(n_287),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_306),
.B(n_309),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_301),
.B(n_307),
.C(n_308),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_310),
.B(n_316),
.Y(n_317)
);

OAI21xp5_ASAP7_75t_L g314 ( 
.A1(n_309),
.A2(n_300),
.B(n_291),
.Y(n_314)
);

INVxp67_ASAP7_75t_L g318 ( 
.A(n_314),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_301),
.B(n_16),
.C(n_3),
.Y(n_316)
);

AND2x2_ASAP7_75t_L g319 ( 
.A(n_311),
.B(n_16),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_319),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_320),
.B(n_311),
.C(n_313),
.Y(n_321)
);

AO21x1_ASAP7_75t_L g322 ( 
.A1(n_321),
.A2(n_312),
.B(n_315),
.Y(n_322)
);

XNOR2xp5_ASAP7_75t_L g323 ( 
.A(n_322),
.B(n_317),
.Y(n_323)
);

XOR2xp5_ASAP7_75t_L g324 ( 
.A(n_323),
.B(n_318),
.Y(n_324)
);


endmodule