module fake_aes_9483_n_640 (n_44, n_81, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_80, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_84, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_83, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_82, n_15, n_61, n_21, n_51, n_39, n_640);
input n_44;
input n_81;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_80;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_84;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_83;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_82;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_640;
wire n_117;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_162;
wire n_387;
wire n_163;
wire n_476;
wire n_105;
wire n_227;
wire n_434;
wire n_384;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_586;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_367;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_446;
wire n_423;
wire n_342;
wire n_420;
wire n_621;
wire n_370;
wire n_589;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_90;
wire n_357;
wire n_260;
wire n_539;
wire n_201;
wire n_197;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_573;
wire n_126;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_429;
wire n_488;
wire n_233;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_132;
wire n_99;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g85 ( .A(n_83), .Y(n_85) );
NOR2xp67_ASAP7_75t_L g86 ( .A(n_62), .B(n_31), .Y(n_86) );
INVxp67_ASAP7_75t_L g87 ( .A(n_0), .Y(n_87) );
INVxp33_ASAP7_75t_SL g88 ( .A(n_23), .Y(n_88) );
INVxp67_ASAP7_75t_SL g89 ( .A(n_60), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_44), .Y(n_90) );
INVxp67_ASAP7_75t_L g91 ( .A(n_37), .Y(n_91) );
CKINVDCx5p33_ASAP7_75t_R g92 ( .A(n_14), .Y(n_92) );
INVx2_ASAP7_75t_L g93 ( .A(n_15), .Y(n_93) );
INVx2_ASAP7_75t_L g94 ( .A(n_42), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_58), .Y(n_95) );
HB1xp67_ASAP7_75t_L g96 ( .A(n_26), .Y(n_96) );
CKINVDCx5p33_ASAP7_75t_R g97 ( .A(n_80), .Y(n_97) );
CKINVDCx16_ASAP7_75t_R g98 ( .A(n_47), .Y(n_98) );
CKINVDCx5p33_ASAP7_75t_R g99 ( .A(n_1), .Y(n_99) );
INVx2_ASAP7_75t_L g100 ( .A(n_72), .Y(n_100) );
CKINVDCx16_ASAP7_75t_R g101 ( .A(n_48), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_16), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_45), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_49), .Y(n_104) );
INVx3_ASAP7_75t_L g105 ( .A(n_35), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_33), .Y(n_106) );
BUFx6f_ASAP7_75t_L g107 ( .A(n_0), .Y(n_107) );
CKINVDCx5p33_ASAP7_75t_R g108 ( .A(n_64), .Y(n_108) );
CKINVDCx5p33_ASAP7_75t_R g109 ( .A(n_25), .Y(n_109) );
CKINVDCx5p33_ASAP7_75t_R g110 ( .A(n_65), .Y(n_110) );
CKINVDCx5p33_ASAP7_75t_R g111 ( .A(n_4), .Y(n_111) );
HB1xp67_ASAP7_75t_L g112 ( .A(n_19), .Y(n_112) );
BUFx3_ASAP7_75t_L g113 ( .A(n_2), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_67), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_40), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_69), .Y(n_116) );
INVx2_ASAP7_75t_L g117 ( .A(n_75), .Y(n_117) );
BUFx6f_ASAP7_75t_L g118 ( .A(n_21), .Y(n_118) );
INVxp67_ASAP7_75t_L g119 ( .A(n_3), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_2), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_9), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_70), .Y(n_122) );
HB1xp67_ASAP7_75t_L g123 ( .A(n_113), .Y(n_123) );
INVx3_ASAP7_75t_L g124 ( .A(n_113), .Y(n_124) );
INVx3_ASAP7_75t_L g125 ( .A(n_113), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_93), .Y(n_126) );
INVx2_ASAP7_75t_L g127 ( .A(n_105), .Y(n_127) );
NOR2xp33_ASAP7_75t_L g128 ( .A(n_96), .B(n_1), .Y(n_128) );
BUFx6f_ASAP7_75t_L g129 ( .A(n_118), .Y(n_129) );
BUFx6f_ASAP7_75t_L g130 ( .A(n_118), .Y(n_130) );
INVx5_ASAP7_75t_L g131 ( .A(n_105), .Y(n_131) );
OAI22xp5_ASAP7_75t_L g132 ( .A1(n_98), .A2(n_101), .B1(n_121), .B2(n_120), .Y(n_132) );
INVx2_ASAP7_75t_L g133 ( .A(n_105), .Y(n_133) );
AND2x6_ASAP7_75t_L g134 ( .A(n_105), .B(n_39), .Y(n_134) );
INVx1_ASAP7_75t_L g135 ( .A(n_93), .Y(n_135) );
INVx2_ASAP7_75t_L g136 ( .A(n_118), .Y(n_136) );
NAND2xp5_ASAP7_75t_L g137 ( .A(n_112), .B(n_3), .Y(n_137) );
INVx1_ASAP7_75t_L g138 ( .A(n_93), .Y(n_138) );
INVx4_ASAP7_75t_L g139 ( .A(n_118), .Y(n_139) );
INVx2_ASAP7_75t_L g140 ( .A(n_118), .Y(n_140) );
HB1xp67_ASAP7_75t_L g141 ( .A(n_87), .Y(n_141) );
AND2x2_ASAP7_75t_L g142 ( .A(n_98), .B(n_4), .Y(n_142) );
NAND2xp33_ASAP7_75t_L g143 ( .A(n_118), .B(n_84), .Y(n_143) );
AND2x2_ASAP7_75t_L g144 ( .A(n_101), .B(n_5), .Y(n_144) );
INVx2_ASAP7_75t_L g145 ( .A(n_94), .Y(n_145) );
AND2x4_ASAP7_75t_L g146 ( .A(n_102), .B(n_5), .Y(n_146) );
INVxp67_ASAP7_75t_L g147 ( .A(n_102), .Y(n_147) );
AND2x4_ASAP7_75t_L g148 ( .A(n_120), .B(n_6), .Y(n_148) );
INVx2_ASAP7_75t_L g149 ( .A(n_94), .Y(n_149) );
NAND2xp5_ASAP7_75t_L g150 ( .A(n_119), .B(n_6), .Y(n_150) );
NAND2xp5_ASAP7_75t_SL g151 ( .A(n_131), .B(n_100), .Y(n_151) );
INVx1_ASAP7_75t_L g152 ( .A(n_146), .Y(n_152) );
BUFx4f_ASAP7_75t_L g153 ( .A(n_134), .Y(n_153) );
NAND2xp5_ASAP7_75t_SL g154 ( .A(n_131), .B(n_100), .Y(n_154) );
NAND3xp33_ASAP7_75t_L g155 ( .A(n_132), .B(n_92), .C(n_99), .Y(n_155) );
AND2x4_ASAP7_75t_L g156 ( .A(n_123), .B(n_121), .Y(n_156) );
OR2x6_ASAP7_75t_L g157 ( .A(n_142), .B(n_107), .Y(n_157) );
INVx1_ASAP7_75t_L g158 ( .A(n_146), .Y(n_158) );
AOI22xp5_ASAP7_75t_L g159 ( .A1(n_141), .A2(n_111), .B1(n_88), .B2(n_107), .Y(n_159) );
OR2x2_ASAP7_75t_L g160 ( .A(n_147), .B(n_107), .Y(n_160) );
NAND2xp5_ASAP7_75t_L g161 ( .A(n_131), .B(n_97), .Y(n_161) );
INVx1_ASAP7_75t_L g162 ( .A(n_146), .Y(n_162) );
NAND2xp5_ASAP7_75t_SL g163 ( .A(n_131), .B(n_117), .Y(n_163) );
CKINVDCx5p33_ASAP7_75t_R g164 ( .A(n_142), .Y(n_164) );
INVx1_ASAP7_75t_L g165 ( .A(n_146), .Y(n_165) );
AND2x2_ASAP7_75t_L g166 ( .A(n_144), .B(n_107), .Y(n_166) );
OR2x6_ASAP7_75t_L g167 ( .A(n_144), .B(n_107), .Y(n_167) );
INVx3_ASAP7_75t_L g168 ( .A(n_148), .Y(n_168) );
INVx2_ASAP7_75t_SL g169 ( .A(n_131), .Y(n_169) );
NOR2xp33_ASAP7_75t_L g170 ( .A(n_131), .B(n_91), .Y(n_170) );
INVx1_ASAP7_75t_L g171 ( .A(n_148), .Y(n_171) );
OR2x6_ASAP7_75t_L g172 ( .A(n_148), .B(n_107), .Y(n_172) );
INVx2_ASAP7_75t_L g173 ( .A(n_139), .Y(n_173) );
BUFx2_ASAP7_75t_L g174 ( .A(n_137), .Y(n_174) );
AND2x2_ASAP7_75t_L g175 ( .A(n_124), .B(n_85), .Y(n_175) );
BUFx4f_ASAP7_75t_L g176 ( .A(n_134), .Y(n_176) );
INVx2_ASAP7_75t_L g177 ( .A(n_139), .Y(n_177) );
INVx1_ASAP7_75t_SL g178 ( .A(n_150), .Y(n_178) );
INVx1_ASAP7_75t_L g179 ( .A(n_148), .Y(n_179) );
INVx1_ASAP7_75t_SL g180 ( .A(n_127), .Y(n_180) );
AND2x2_ASAP7_75t_L g181 ( .A(n_124), .B(n_85), .Y(n_181) );
NAND2xp5_ASAP7_75t_SL g182 ( .A(n_127), .B(n_117), .Y(n_182) );
INVx1_ASAP7_75t_L g183 ( .A(n_127), .Y(n_183) );
AOI22xp5_ASAP7_75t_L g184 ( .A1(n_128), .A2(n_89), .B1(n_116), .B2(n_115), .Y(n_184) );
NAND2xp5_ASAP7_75t_L g185 ( .A(n_124), .B(n_108), .Y(n_185) );
BUFx3_ASAP7_75t_L g186 ( .A(n_153), .Y(n_186) );
NAND2xp5_ASAP7_75t_SL g187 ( .A(n_153), .B(n_133), .Y(n_187) );
INVx1_ASAP7_75t_L g188 ( .A(n_160), .Y(n_188) );
AND2x4_ASAP7_75t_L g189 ( .A(n_157), .B(n_167), .Y(n_189) );
AND2x2_ASAP7_75t_L g190 ( .A(n_174), .B(n_133), .Y(n_190) );
O2A1O1Ixp33_ASAP7_75t_L g191 ( .A1(n_152), .A2(n_149), .B(n_145), .C(n_126), .Y(n_191) );
NAND2xp5_ASAP7_75t_SL g192 ( .A(n_153), .B(n_133), .Y(n_192) );
OR2x2_ASAP7_75t_L g193 ( .A(n_178), .B(n_124), .Y(n_193) );
NOR2xp33_ASAP7_75t_L g194 ( .A(n_156), .B(n_90), .Y(n_194) );
NOR3xp33_ASAP7_75t_L g195 ( .A(n_155), .B(n_122), .C(n_90), .Y(n_195) );
OR2x2_ASAP7_75t_L g196 ( .A(n_156), .B(n_125), .Y(n_196) );
BUFx6f_ASAP7_75t_SL g197 ( .A(n_156), .Y(n_197) );
AOI22xp33_ASAP7_75t_L g198 ( .A1(n_158), .A2(n_134), .B1(n_149), .B2(n_145), .Y(n_198) );
NAND2xp5_ASAP7_75t_L g199 ( .A(n_180), .B(n_125), .Y(n_199) );
NAND2xp5_ASAP7_75t_L g200 ( .A(n_166), .B(n_125), .Y(n_200) );
INVx2_ASAP7_75t_L g201 ( .A(n_183), .Y(n_201) );
NAND2xp5_ASAP7_75t_L g202 ( .A(n_175), .B(n_125), .Y(n_202) );
INVx2_ASAP7_75t_L g203 ( .A(n_168), .Y(n_203) );
NAND2xp5_ASAP7_75t_SL g204 ( .A(n_176), .B(n_95), .Y(n_204) );
INVx2_ASAP7_75t_SL g205 ( .A(n_157), .Y(n_205) );
NAND2xp5_ASAP7_75t_L g206 ( .A(n_175), .B(n_134), .Y(n_206) );
NOR2x1p5_ASAP7_75t_L g207 ( .A(n_164), .B(n_95), .Y(n_207) );
NAND2xp5_ASAP7_75t_L g208 ( .A(n_181), .B(n_134), .Y(n_208) );
NOR2xp33_ASAP7_75t_L g209 ( .A(n_184), .B(n_103), .Y(n_209) );
INVx3_ASAP7_75t_L g210 ( .A(n_172), .Y(n_210) );
AND2x6_ASAP7_75t_SL g211 ( .A(n_157), .B(n_126), .Y(n_211) );
NAND2xp5_ASAP7_75t_L g212 ( .A(n_181), .B(n_134), .Y(n_212) );
INVxp67_ASAP7_75t_L g213 ( .A(n_164), .Y(n_213) );
BUFx6f_ASAP7_75t_L g214 ( .A(n_176), .Y(n_214) );
INVx3_ASAP7_75t_L g215 ( .A(n_172), .Y(n_215) );
INVx8_ASAP7_75t_L g216 ( .A(n_157), .Y(n_216) );
AOI21xp5_ASAP7_75t_L g217 ( .A1(n_176), .A2(n_143), .B(n_149), .Y(n_217) );
INVx1_ASAP7_75t_SL g218 ( .A(n_167), .Y(n_218) );
INVx1_ASAP7_75t_L g219 ( .A(n_167), .Y(n_219) );
INVx1_ASAP7_75t_L g220 ( .A(n_167), .Y(n_220) );
NOR2xp33_ASAP7_75t_L g221 ( .A(n_162), .B(n_103), .Y(n_221) );
OR2x6_ASAP7_75t_L g222 ( .A(n_172), .B(n_104), .Y(n_222) );
NAND2xp5_ASAP7_75t_L g223 ( .A(n_168), .B(n_134), .Y(n_223) );
INVx1_ASAP7_75t_L g224 ( .A(n_172), .Y(n_224) );
NOR2xp33_ASAP7_75t_L g225 ( .A(n_165), .B(n_104), .Y(n_225) );
NAND2xp5_ASAP7_75t_L g226 ( .A(n_168), .B(n_134), .Y(n_226) );
NAND2xp5_ASAP7_75t_L g227 ( .A(n_171), .B(n_109), .Y(n_227) );
HB1xp67_ASAP7_75t_L g228 ( .A(n_159), .Y(n_228) );
INVx3_ASAP7_75t_L g229 ( .A(n_179), .Y(n_229) );
OR2x6_ASAP7_75t_L g230 ( .A(n_182), .B(n_106), .Y(n_230) );
OAI21x1_ASAP7_75t_L g231 ( .A1(n_217), .A2(n_182), .B(n_151), .Y(n_231) );
NAND2xp5_ASAP7_75t_L g232 ( .A(n_190), .B(n_185), .Y(n_232) );
NAND2xp5_ASAP7_75t_L g233 ( .A(n_193), .B(n_194), .Y(n_233) );
OAI22xp5_ASAP7_75t_L g234 ( .A1(n_189), .A2(n_222), .B1(n_218), .B2(n_216), .Y(n_234) );
NAND2xp5_ASAP7_75t_SL g235 ( .A(n_189), .B(n_161), .Y(n_235) );
INVx2_ASAP7_75t_L g236 ( .A(n_203), .Y(n_236) );
OAI22xp5_ASAP7_75t_L g237 ( .A1(n_189), .A2(n_170), .B1(n_145), .B2(n_177), .Y(n_237) );
O2A1O1Ixp33_ASAP7_75t_L g238 ( .A1(n_209), .A2(n_163), .B(n_154), .C(n_151), .Y(n_238) );
NAND2xp5_ASAP7_75t_SL g239 ( .A(n_210), .B(n_169), .Y(n_239) );
A2O1A1Ixp33_ASAP7_75t_L g240 ( .A1(n_221), .A2(n_138), .B(n_135), .C(n_114), .Y(n_240) );
AND2x2_ASAP7_75t_L g241 ( .A(n_222), .B(n_135), .Y(n_241) );
NAND2xp5_ASAP7_75t_L g242 ( .A(n_194), .B(n_169), .Y(n_242) );
NAND2xp5_ASAP7_75t_L g243 ( .A(n_196), .B(n_138), .Y(n_243) );
NAND2xp5_ASAP7_75t_SL g244 ( .A(n_210), .B(n_110), .Y(n_244) );
NAND2xp5_ASAP7_75t_L g245 ( .A(n_209), .B(n_177), .Y(n_245) );
AOI21xp5_ASAP7_75t_L g246 ( .A1(n_223), .A2(n_226), .B(n_206), .Y(n_246) );
O2A1O1Ixp5_ASAP7_75t_L g247 ( .A1(n_204), .A2(n_163), .B(n_154), .C(n_139), .Y(n_247) );
NAND2xp5_ASAP7_75t_L g248 ( .A(n_188), .B(n_173), .Y(n_248) );
NAND2xp5_ASAP7_75t_SL g249 ( .A(n_210), .B(n_173), .Y(n_249) );
NOR2xp67_ASAP7_75t_SL g250 ( .A(n_215), .B(n_122), .Y(n_250) );
INVx3_ASAP7_75t_L g251 ( .A(n_215), .Y(n_251) );
BUFx12f_ASAP7_75t_L g252 ( .A(n_211), .Y(n_252) );
AOI21xp5_ASAP7_75t_L g253 ( .A1(n_208), .A2(n_116), .B(n_106), .Y(n_253) );
AND2x2_ASAP7_75t_L g254 ( .A(n_222), .B(n_114), .Y(n_254) );
AOI21xp5_ASAP7_75t_L g255 ( .A1(n_212), .A2(n_115), .B(n_86), .Y(n_255) );
OAI22xp5_ASAP7_75t_L g256 ( .A1(n_216), .A2(n_139), .B1(n_86), .B2(n_136), .Y(n_256) );
AND2x2_ASAP7_75t_L g257 ( .A(n_201), .B(n_7), .Y(n_257) );
O2A1O1Ixp33_ASAP7_75t_L g258 ( .A1(n_228), .A2(n_140), .B(n_136), .C(n_9), .Y(n_258) );
OAI21xp5_ASAP7_75t_L g259 ( .A1(n_198), .A2(n_140), .B(n_136), .Y(n_259) );
OAI21xp5_ASAP7_75t_L g260 ( .A1(n_198), .A2(n_140), .B(n_130), .Y(n_260) );
CKINVDCx5p33_ASAP7_75t_R g261 ( .A(n_197), .Y(n_261) );
NAND2xp5_ASAP7_75t_SL g262 ( .A(n_215), .B(n_205), .Y(n_262) );
NOR2xp33_ASAP7_75t_R g263 ( .A(n_197), .B(n_7), .Y(n_263) );
CKINVDCx14_ASAP7_75t_R g264 ( .A(n_216), .Y(n_264) );
NAND2xp5_ASAP7_75t_L g265 ( .A(n_229), .B(n_8), .Y(n_265) );
NAND2xp5_ASAP7_75t_SL g266 ( .A(n_224), .B(n_130), .Y(n_266) );
CKINVDCx16_ASAP7_75t_R g267 ( .A(n_230), .Y(n_267) );
OAI22xp5_ASAP7_75t_L g268 ( .A1(n_219), .A2(n_130), .B1(n_129), .B2(n_11), .Y(n_268) );
NOR2xp33_ASAP7_75t_L g269 ( .A(n_213), .B(n_8), .Y(n_269) );
CKINVDCx20_ASAP7_75t_R g270 ( .A(n_220), .Y(n_270) );
AOI21xp5_ASAP7_75t_L g271 ( .A1(n_187), .A2(n_130), .B(n_129), .Y(n_271) );
NAND2xp5_ASAP7_75t_SL g272 ( .A(n_214), .B(n_130), .Y(n_272) );
NOR2xp33_ASAP7_75t_R g273 ( .A(n_229), .B(n_10), .Y(n_273) );
BUFx3_ASAP7_75t_L g274 ( .A(n_186), .Y(n_274) );
NAND2xp5_ASAP7_75t_L g275 ( .A(n_233), .B(n_207), .Y(n_275) );
INVx2_ASAP7_75t_L g276 ( .A(n_236), .Y(n_276) );
INVx1_ASAP7_75t_L g277 ( .A(n_257), .Y(n_277) );
INVx2_ASAP7_75t_L g278 ( .A(n_236), .Y(n_278) );
O2A1O1Ixp33_ASAP7_75t_SL g279 ( .A1(n_240), .A2(n_187), .B(n_192), .C(n_204), .Y(n_279) );
A2O1A1Ixp33_ASAP7_75t_L g280 ( .A1(n_258), .A2(n_221), .B(n_225), .C(n_191), .Y(n_280) );
O2A1O1Ixp33_ASAP7_75t_L g281 ( .A1(n_240), .A2(n_195), .B(n_225), .C(n_202), .Y(n_281) );
OAI21x1_ASAP7_75t_L g282 ( .A1(n_271), .A2(n_192), .B(n_203), .Y(n_282) );
OAI21xp33_ASAP7_75t_L g283 ( .A1(n_232), .A2(n_199), .B(n_227), .Y(n_283) );
AO31x2_ASAP7_75t_L g284 ( .A1(n_255), .A2(n_201), .A3(n_200), .B(n_130), .Y(n_284) );
OAI22xp33_ASAP7_75t_L g285 ( .A1(n_267), .A2(n_230), .B1(n_229), .B2(n_186), .Y(n_285) );
A2O1A1Ixp33_ASAP7_75t_L g286 ( .A1(n_253), .A2(n_214), .B(n_129), .C(n_230), .Y(n_286) );
OAI22xp5_ASAP7_75t_L g287 ( .A1(n_234), .A2(n_214), .B1(n_129), .B2(n_12), .Y(n_287) );
OAI21xp5_ASAP7_75t_L g288 ( .A1(n_246), .A2(n_214), .B(n_129), .Y(n_288) );
OAI21xp5_ASAP7_75t_L g289 ( .A1(n_260), .A2(n_129), .B(n_50), .Y(n_289) );
INVx2_ASAP7_75t_L g290 ( .A(n_257), .Y(n_290) );
AOI22xp5_ASAP7_75t_L g291 ( .A1(n_270), .A2(n_10), .B1(n_11), .B2(n_12), .Y(n_291) );
OAI21xp5_ASAP7_75t_L g292 ( .A1(n_231), .A2(n_51), .B(n_81), .Y(n_292) );
O2A1O1Ixp33_ASAP7_75t_SL g293 ( .A1(n_265), .A2(n_46), .B(n_79), .C(n_78), .Y(n_293) );
CKINVDCx20_ASAP7_75t_R g294 ( .A(n_263), .Y(n_294) );
INVx3_ASAP7_75t_L g295 ( .A(n_251), .Y(n_295) );
AOI21xp5_ASAP7_75t_L g296 ( .A1(n_242), .A2(n_43), .B(n_77), .Y(n_296) );
AO21x2_ASAP7_75t_L g297 ( .A1(n_259), .A2(n_41), .B(n_76), .Y(n_297) );
O2A1O1Ixp33_ASAP7_75t_L g298 ( .A1(n_245), .A2(n_237), .B(n_243), .C(n_269), .Y(n_298) );
O2A1O1Ixp33_ASAP7_75t_L g299 ( .A1(n_238), .A2(n_13), .B(n_14), .C(n_15), .Y(n_299) );
O2A1O1Ixp33_ASAP7_75t_L g300 ( .A1(n_256), .A2(n_13), .B(n_16), .C(n_17), .Y(n_300) );
NOR2xp33_ASAP7_75t_SL g301 ( .A(n_261), .B(n_17), .Y(n_301) );
A2O1A1Ixp33_ASAP7_75t_L g302 ( .A1(n_241), .A2(n_18), .B(n_20), .C(n_22), .Y(n_302) );
O2A1O1Ixp33_ASAP7_75t_L g303 ( .A1(n_241), .A2(n_18), .B(n_24), .C(n_27), .Y(n_303) );
INVx1_ASAP7_75t_L g304 ( .A(n_248), .Y(n_304) );
NOR2xp67_ASAP7_75t_L g305 ( .A(n_261), .B(n_28), .Y(n_305) );
INVx3_ASAP7_75t_L g306 ( .A(n_251), .Y(n_306) );
AOI21xp5_ASAP7_75t_L g307 ( .A1(n_249), .A2(n_29), .B(n_30), .Y(n_307) );
AOI21xp5_ASAP7_75t_L g308 ( .A1(n_266), .A2(n_32), .B(n_34), .Y(n_308) );
INVx2_ASAP7_75t_L g309 ( .A(n_276), .Y(n_309) );
NOR2xp33_ASAP7_75t_L g310 ( .A(n_275), .B(n_270), .Y(n_310) );
AO31x2_ASAP7_75t_L g311 ( .A1(n_280), .A2(n_268), .A3(n_231), .B(n_273), .Y(n_311) );
A2O1A1Ixp33_ASAP7_75t_L g312 ( .A1(n_298), .A2(n_254), .B(n_251), .C(n_247), .Y(n_312) );
NOR2xp33_ASAP7_75t_L g313 ( .A(n_285), .B(n_252), .Y(n_313) );
INVx3_ASAP7_75t_L g314 ( .A(n_295), .Y(n_314) );
INVx1_ASAP7_75t_L g315 ( .A(n_304), .Y(n_315) );
OAI211xp5_ASAP7_75t_SL g316 ( .A1(n_291), .A2(n_300), .B(n_299), .C(n_303), .Y(n_316) );
HB1xp67_ASAP7_75t_L g317 ( .A(n_278), .Y(n_317) );
O2A1O1Ixp33_ASAP7_75t_L g318 ( .A1(n_280), .A2(n_254), .B(n_235), .C(n_244), .Y(n_318) );
AO31x2_ASAP7_75t_L g319 ( .A1(n_286), .A2(n_250), .A3(n_272), .B(n_274), .Y(n_319) );
INVx1_ASAP7_75t_L g320 ( .A(n_277), .Y(n_320) );
INVx2_ASAP7_75t_L g321 ( .A(n_282), .Y(n_321) );
NAND2xp5_ASAP7_75t_L g322 ( .A(n_290), .B(n_264), .Y(n_322) );
AOI21xp5_ASAP7_75t_L g323 ( .A1(n_288), .A2(n_239), .B(n_262), .Y(n_323) );
AOI22xp33_ASAP7_75t_L g324 ( .A1(n_285), .A2(n_252), .B1(n_283), .B2(n_287), .Y(n_324) );
INVx2_ASAP7_75t_SL g325 ( .A(n_295), .Y(n_325) );
INVxp33_ASAP7_75t_L g326 ( .A(n_301), .Y(n_326) );
INVx2_ASAP7_75t_L g327 ( .A(n_284), .Y(n_327) );
OAI22xp5_ASAP7_75t_L g328 ( .A1(n_286), .A2(n_264), .B1(n_274), .B2(n_52), .Y(n_328) );
INVx1_ASAP7_75t_L g329 ( .A(n_306), .Y(n_329) );
AOI21xp5_ASAP7_75t_L g330 ( .A1(n_279), .A2(n_36), .B(n_38), .Y(n_330) );
OAI21x1_ASAP7_75t_L g331 ( .A1(n_289), .A2(n_53), .B(n_54), .Y(n_331) );
INVx4_ASAP7_75t_L g332 ( .A(n_306), .Y(n_332) );
O2A1O1Ixp33_ASAP7_75t_L g333 ( .A1(n_281), .A2(n_55), .B(n_56), .C(n_57), .Y(n_333) );
AND2x2_ASAP7_75t_L g334 ( .A(n_302), .B(n_59), .Y(n_334) );
INVx1_ASAP7_75t_L g335 ( .A(n_284), .Y(n_335) );
NOR2xp33_ASAP7_75t_L g336 ( .A(n_322), .B(n_294), .Y(n_336) );
AO21x2_ASAP7_75t_L g337 ( .A1(n_335), .A2(n_292), .B(n_297), .Y(n_337) );
OR2x6_ASAP7_75t_L g338 ( .A(n_327), .B(n_296), .Y(n_338) );
INVx2_ASAP7_75t_L g339 ( .A(n_327), .Y(n_339) );
AND2x2_ASAP7_75t_L g340 ( .A(n_309), .B(n_284), .Y(n_340) );
NAND2xp5_ASAP7_75t_L g341 ( .A(n_320), .B(n_284), .Y(n_341) );
NAND2xp5_ASAP7_75t_SL g342 ( .A(n_327), .B(n_305), .Y(n_342) );
AO22x1_ASAP7_75t_L g343 ( .A1(n_326), .A2(n_293), .B1(n_297), .B2(n_279), .Y(n_343) );
AO21x1_ASAP7_75t_SL g344 ( .A1(n_335), .A2(n_293), .B(n_307), .Y(n_344) );
BUFx6f_ASAP7_75t_L g345 ( .A(n_321), .Y(n_345) );
INVx1_ASAP7_75t_L g346 ( .A(n_320), .Y(n_346) );
OAI21x1_ASAP7_75t_L g347 ( .A1(n_331), .A2(n_308), .B(n_63), .Y(n_347) );
OR2x6_ASAP7_75t_L g348 ( .A(n_328), .B(n_61), .Y(n_348) );
OA21x2_ASAP7_75t_L g349 ( .A1(n_321), .A2(n_66), .B(n_68), .Y(n_349) );
NAND2xp5_ASAP7_75t_L g350 ( .A(n_315), .B(n_71), .Y(n_350) );
OA21x2_ASAP7_75t_L g351 ( .A1(n_321), .A2(n_331), .B(n_330), .Y(n_351) );
AND2x2_ASAP7_75t_L g352 ( .A(n_309), .B(n_73), .Y(n_352) );
NOR2xp33_ASAP7_75t_L g353 ( .A(n_310), .B(n_74), .Y(n_353) );
OR2x2_ASAP7_75t_L g354 ( .A(n_315), .B(n_82), .Y(n_354) );
INVx1_ASAP7_75t_L g355 ( .A(n_309), .Y(n_355) );
NAND2xp5_ASAP7_75t_L g356 ( .A(n_311), .B(n_318), .Y(n_356) );
OA21x2_ASAP7_75t_L g357 ( .A1(n_312), .A2(n_323), .B(n_334), .Y(n_357) );
AND2x2_ASAP7_75t_L g358 ( .A(n_317), .B(n_311), .Y(n_358) );
AND2x2_ASAP7_75t_L g359 ( .A(n_311), .B(n_329), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_329), .Y(n_360) );
INVx2_ASAP7_75t_L g361 ( .A(n_319), .Y(n_361) );
AOI22xp33_ASAP7_75t_L g362 ( .A1(n_316), .A2(n_313), .B1(n_324), .B2(n_334), .Y(n_362) );
INVx2_ASAP7_75t_L g363 ( .A(n_339), .Y(n_363) );
INVx2_ASAP7_75t_L g364 ( .A(n_339), .Y(n_364) );
BUFx3_ASAP7_75t_L g365 ( .A(n_339), .Y(n_365) );
NOR2x1_ASAP7_75t_L g366 ( .A(n_354), .B(n_332), .Y(n_366) );
AOI211xp5_ASAP7_75t_L g367 ( .A1(n_353), .A2(n_333), .B(n_325), .C(n_314), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_341), .Y(n_368) );
INVx1_ASAP7_75t_L g369 ( .A(n_341), .Y(n_369) );
AND2x2_ASAP7_75t_L g370 ( .A(n_359), .B(n_311), .Y(n_370) );
INVx1_ASAP7_75t_L g371 ( .A(n_340), .Y(n_371) );
AND2x2_ASAP7_75t_L g372 ( .A(n_359), .B(n_311), .Y(n_372) );
AND2x2_ASAP7_75t_L g373 ( .A(n_359), .B(n_319), .Y(n_373) );
AO21x2_ASAP7_75t_L g374 ( .A1(n_356), .A2(n_319), .B(n_332), .Y(n_374) );
NAND2xp5_ASAP7_75t_L g375 ( .A(n_346), .B(n_314), .Y(n_375) );
INVx1_ASAP7_75t_L g376 ( .A(n_340), .Y(n_376) );
INVx1_ASAP7_75t_L g377 ( .A(n_340), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_346), .Y(n_378) );
INVx1_ASAP7_75t_L g379 ( .A(n_355), .Y(n_379) );
INVx2_ASAP7_75t_L g380 ( .A(n_345), .Y(n_380) );
INVx2_ASAP7_75t_L g381 ( .A(n_345), .Y(n_381) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_355), .B(n_314), .Y(n_382) );
BUFx3_ASAP7_75t_L g383 ( .A(n_352), .Y(n_383) );
INVx3_ASAP7_75t_L g384 ( .A(n_345), .Y(n_384) );
BUFx6f_ASAP7_75t_L g385 ( .A(n_345), .Y(n_385) );
OR2x2_ASAP7_75t_L g386 ( .A(n_358), .B(n_319), .Y(n_386) );
INVx2_ASAP7_75t_L g387 ( .A(n_345), .Y(n_387) );
INVx1_ASAP7_75t_L g388 ( .A(n_360), .Y(n_388) );
NAND2xp5_ASAP7_75t_L g389 ( .A(n_358), .B(n_314), .Y(n_389) );
INVx1_ASAP7_75t_L g390 ( .A(n_360), .Y(n_390) );
AND2x2_ASAP7_75t_L g391 ( .A(n_358), .B(n_319), .Y(n_391) );
INVx3_ASAP7_75t_L g392 ( .A(n_345), .Y(n_392) );
INVx1_ASAP7_75t_L g393 ( .A(n_361), .Y(n_393) );
AND2x2_ASAP7_75t_L g394 ( .A(n_361), .B(n_332), .Y(n_394) );
OR2x2_ASAP7_75t_L g395 ( .A(n_356), .B(n_332), .Y(n_395) );
INVx1_ASAP7_75t_L g396 ( .A(n_361), .Y(n_396) );
INVx2_ASAP7_75t_L g397 ( .A(n_345), .Y(n_397) );
NAND2xp5_ASAP7_75t_L g398 ( .A(n_362), .B(n_325), .Y(n_398) );
INVx1_ASAP7_75t_L g399 ( .A(n_378), .Y(n_399) );
INVx1_ASAP7_75t_L g400 ( .A(n_378), .Y(n_400) );
INVx1_ASAP7_75t_L g401 ( .A(n_379), .Y(n_401) );
AND2x2_ASAP7_75t_L g402 ( .A(n_373), .B(n_337), .Y(n_402) );
INVx1_ASAP7_75t_L g403 ( .A(n_379), .Y(n_403) );
INVx1_ASAP7_75t_SL g404 ( .A(n_365), .Y(n_404) );
NOR4xp25_ASAP7_75t_SL g405 ( .A(n_368), .B(n_342), .C(n_343), .D(n_362), .Y(n_405) );
AND2x2_ASAP7_75t_L g406 ( .A(n_373), .B(n_337), .Y(n_406) );
AND2x2_ASAP7_75t_L g407 ( .A(n_373), .B(n_337), .Y(n_407) );
NAND2x1p5_ASAP7_75t_L g408 ( .A(n_366), .B(n_354), .Y(n_408) );
AND2x2_ASAP7_75t_L g409 ( .A(n_391), .B(n_337), .Y(n_409) );
AND2x2_ASAP7_75t_L g410 ( .A(n_391), .B(n_357), .Y(n_410) );
INVx1_ASAP7_75t_L g411 ( .A(n_388), .Y(n_411) );
NOR2xp67_ASAP7_75t_L g412 ( .A(n_363), .B(n_354), .Y(n_412) );
INVx1_ASAP7_75t_L g413 ( .A(n_388), .Y(n_413) );
INVx2_ASAP7_75t_L g414 ( .A(n_393), .Y(n_414) );
NAND2x1p5_ASAP7_75t_L g415 ( .A(n_366), .B(n_352), .Y(n_415) );
INVx1_ASAP7_75t_L g416 ( .A(n_390), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_390), .Y(n_417) );
AND2x2_ASAP7_75t_L g418 ( .A(n_391), .B(n_357), .Y(n_418) );
AND2x2_ASAP7_75t_L g419 ( .A(n_371), .B(n_357), .Y(n_419) );
INVx1_ASAP7_75t_SL g420 ( .A(n_365), .Y(n_420) );
NAND2xp5_ASAP7_75t_L g421 ( .A(n_368), .B(n_357), .Y(n_421) );
INVx1_ASAP7_75t_L g422 ( .A(n_369), .Y(n_422) );
AND2x2_ASAP7_75t_L g423 ( .A(n_371), .B(n_357), .Y(n_423) );
INVx2_ASAP7_75t_L g424 ( .A(n_393), .Y(n_424) );
NAND2xp5_ASAP7_75t_L g425 ( .A(n_369), .B(n_343), .Y(n_425) );
AND2x2_ASAP7_75t_L g426 ( .A(n_376), .B(n_338), .Y(n_426) );
AND2x2_ASAP7_75t_L g427 ( .A(n_376), .B(n_338), .Y(n_427) );
INVx1_ASAP7_75t_L g428 ( .A(n_396), .Y(n_428) );
INVx1_ASAP7_75t_L g429 ( .A(n_396), .Y(n_429) );
INVx4_ASAP7_75t_L g430 ( .A(n_365), .Y(n_430) );
AND2x2_ASAP7_75t_L g431 ( .A(n_377), .B(n_338), .Y(n_431) );
OR2x2_ASAP7_75t_L g432 ( .A(n_377), .B(n_338), .Y(n_432) );
AND2x2_ASAP7_75t_L g433 ( .A(n_370), .B(n_338), .Y(n_433) );
AND2x2_ASAP7_75t_L g434 ( .A(n_370), .B(n_338), .Y(n_434) );
AND2x4_ASAP7_75t_SL g435 ( .A(n_394), .B(n_348), .Y(n_435) );
AND2x2_ASAP7_75t_L g436 ( .A(n_370), .B(n_352), .Y(n_436) );
AND2x2_ASAP7_75t_L g437 ( .A(n_372), .B(n_351), .Y(n_437) );
AND2x2_ASAP7_75t_L g438 ( .A(n_372), .B(n_351), .Y(n_438) );
AND2x2_ASAP7_75t_L g439 ( .A(n_372), .B(n_351), .Y(n_439) );
INVx1_ASAP7_75t_SL g440 ( .A(n_363), .Y(n_440) );
BUFx3_ASAP7_75t_L g441 ( .A(n_394), .Y(n_441) );
INVx1_ASAP7_75t_L g442 ( .A(n_375), .Y(n_442) );
NAND2xp5_ASAP7_75t_L g443 ( .A(n_375), .B(n_350), .Y(n_443) );
INVx2_ASAP7_75t_L g444 ( .A(n_363), .Y(n_444) );
AND2x2_ASAP7_75t_L g445 ( .A(n_386), .B(n_351), .Y(n_445) );
AND2x4_ASAP7_75t_L g446 ( .A(n_394), .B(n_342), .Y(n_446) );
INVx2_ASAP7_75t_L g447 ( .A(n_364), .Y(n_447) );
OR2x2_ASAP7_75t_L g448 ( .A(n_386), .B(n_348), .Y(n_448) );
NAND2xp5_ASAP7_75t_L g449 ( .A(n_398), .B(n_350), .Y(n_449) );
INVx1_ASAP7_75t_L g450 ( .A(n_364), .Y(n_450) );
INVx1_ASAP7_75t_L g451 ( .A(n_399), .Y(n_451) );
INVx1_ASAP7_75t_L g452 ( .A(n_399), .Y(n_452) );
INVx1_ASAP7_75t_L g453 ( .A(n_400), .Y(n_453) );
AND2x2_ASAP7_75t_L g454 ( .A(n_410), .B(n_374), .Y(n_454) );
INVx1_ASAP7_75t_L g455 ( .A(n_400), .Y(n_455) );
AND2x2_ASAP7_75t_L g456 ( .A(n_410), .B(n_374), .Y(n_456) );
HB1xp67_ASAP7_75t_L g457 ( .A(n_441), .Y(n_457) );
OAI22xp5_ASAP7_75t_L g458 ( .A1(n_435), .A2(n_348), .B1(n_383), .B2(n_398), .Y(n_458) );
INVx1_ASAP7_75t_L g459 ( .A(n_411), .Y(n_459) );
OR2x2_ASAP7_75t_L g460 ( .A(n_441), .B(n_389), .Y(n_460) );
INVx2_ASAP7_75t_L g461 ( .A(n_444), .Y(n_461) );
INVxp33_ASAP7_75t_L g462 ( .A(n_408), .Y(n_462) );
AND2x2_ASAP7_75t_L g463 ( .A(n_418), .B(n_374), .Y(n_463) );
INVx1_ASAP7_75t_L g464 ( .A(n_411), .Y(n_464) );
OR2x2_ASAP7_75t_L g465 ( .A(n_441), .B(n_389), .Y(n_465) );
INVx3_ASAP7_75t_L g466 ( .A(n_430), .Y(n_466) );
INVx1_ASAP7_75t_L g467 ( .A(n_413), .Y(n_467) );
AOI322xp5_ASAP7_75t_L g468 ( .A1(n_409), .A2(n_353), .A3(n_336), .B1(n_383), .B2(n_382), .C1(n_364), .C2(n_380), .Y(n_468) );
INVx2_ASAP7_75t_L g469 ( .A(n_444), .Y(n_469) );
INVx1_ASAP7_75t_L g470 ( .A(n_413), .Y(n_470) );
AND2x2_ASAP7_75t_L g471 ( .A(n_418), .B(n_374), .Y(n_471) );
AND2x2_ASAP7_75t_L g472 ( .A(n_402), .B(n_395), .Y(n_472) );
HB1xp67_ASAP7_75t_L g473 ( .A(n_414), .Y(n_473) );
INVx1_ASAP7_75t_L g474 ( .A(n_416), .Y(n_474) );
INVx1_ASAP7_75t_L g475 ( .A(n_416), .Y(n_475) );
AND2x2_ASAP7_75t_L g476 ( .A(n_402), .B(n_395), .Y(n_476) );
AND2x2_ASAP7_75t_L g477 ( .A(n_406), .B(n_407), .Y(n_477) );
AND2x2_ASAP7_75t_L g478 ( .A(n_406), .B(n_383), .Y(n_478) );
INVx1_ASAP7_75t_SL g479 ( .A(n_404), .Y(n_479) );
INVx1_ASAP7_75t_L g480 ( .A(n_417), .Y(n_480) );
INVxp67_ASAP7_75t_L g481 ( .A(n_422), .Y(n_481) );
INVx1_ASAP7_75t_L g482 ( .A(n_417), .Y(n_482) );
AND2x2_ASAP7_75t_L g483 ( .A(n_407), .B(n_409), .Y(n_483) );
NAND3xp33_ASAP7_75t_L g484 ( .A(n_405), .B(n_367), .C(n_382), .Y(n_484) );
NAND2xp5_ASAP7_75t_L g485 ( .A(n_442), .B(n_392), .Y(n_485) );
INVx4_ASAP7_75t_L g486 ( .A(n_435), .Y(n_486) );
NAND2x1p5_ASAP7_75t_L g487 ( .A(n_412), .B(n_349), .Y(n_487) );
INVx2_ASAP7_75t_L g488 ( .A(n_444), .Y(n_488) );
NOR2x1_ASAP7_75t_R g489 ( .A(n_430), .B(n_336), .Y(n_489) );
INVx1_ASAP7_75t_L g490 ( .A(n_401), .Y(n_490) );
AND2x2_ASAP7_75t_L g491 ( .A(n_437), .B(n_380), .Y(n_491) );
INVx2_ASAP7_75t_L g492 ( .A(n_447), .Y(n_492) );
INVx1_ASAP7_75t_L g493 ( .A(n_401), .Y(n_493) );
INVx1_ASAP7_75t_L g494 ( .A(n_403), .Y(n_494) );
OR2x2_ASAP7_75t_L g495 ( .A(n_437), .B(n_380), .Y(n_495) );
AND2x4_ASAP7_75t_L g496 ( .A(n_435), .B(n_392), .Y(n_496) );
AND2x2_ASAP7_75t_L g497 ( .A(n_438), .B(n_381), .Y(n_497) );
NAND2xp5_ASAP7_75t_L g498 ( .A(n_442), .B(n_392), .Y(n_498) );
NOR3x1_ASAP7_75t_L g499 ( .A(n_448), .B(n_347), .C(n_348), .Y(n_499) );
AND2x2_ASAP7_75t_L g500 ( .A(n_438), .B(n_381), .Y(n_500) );
AOI21xp33_ASAP7_75t_L g501 ( .A1(n_425), .A2(n_367), .B(n_348), .Y(n_501) );
INVx1_ASAP7_75t_L g502 ( .A(n_403), .Y(n_502) );
OR2x2_ASAP7_75t_L g503 ( .A(n_439), .B(n_432), .Y(n_503) );
NAND2xp5_ASAP7_75t_L g504 ( .A(n_422), .B(n_392), .Y(n_504) );
AND2x2_ASAP7_75t_L g505 ( .A(n_439), .B(n_381), .Y(n_505) );
INVx1_ASAP7_75t_L g506 ( .A(n_428), .Y(n_506) );
OAI21xp5_ASAP7_75t_L g507 ( .A1(n_412), .A2(n_348), .B(n_349), .Y(n_507) );
INVx1_ASAP7_75t_L g508 ( .A(n_428), .Y(n_508) );
OR2x2_ASAP7_75t_L g509 ( .A(n_432), .B(n_397), .Y(n_509) );
INVx2_ASAP7_75t_L g510 ( .A(n_495), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g511 ( .A(n_477), .B(n_423), .Y(n_511) );
NOR2xp33_ASAP7_75t_L g512 ( .A(n_489), .B(n_449), .Y(n_512) );
OR2x2_ASAP7_75t_L g513 ( .A(n_503), .B(n_448), .Y(n_513) );
INVx2_ASAP7_75t_L g514 ( .A(n_495), .Y(n_514) );
INVx1_ASAP7_75t_L g515 ( .A(n_451), .Y(n_515) );
AND2x2_ASAP7_75t_SL g516 ( .A(n_486), .B(n_430), .Y(n_516) );
AND2x2_ASAP7_75t_L g517 ( .A(n_477), .B(n_483), .Y(n_517) );
OR2x2_ASAP7_75t_L g518 ( .A(n_503), .B(n_436), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_483), .B(n_423), .Y(n_519) );
OR2x2_ASAP7_75t_L g520 ( .A(n_472), .B(n_436), .Y(n_520) );
OR2x2_ASAP7_75t_L g521 ( .A(n_472), .B(n_445), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_454), .B(n_419), .Y(n_522) );
INVx1_ASAP7_75t_SL g523 ( .A(n_479), .Y(n_523) );
AND2x2_ASAP7_75t_L g524 ( .A(n_476), .B(n_434), .Y(n_524) );
AND2x2_ASAP7_75t_L g525 ( .A(n_476), .B(n_434), .Y(n_525) );
OAI22xp5_ASAP7_75t_L g526 ( .A1(n_486), .A2(n_408), .B1(n_415), .B2(n_430), .Y(n_526) );
XNOR2xp5_ASAP7_75t_L g527 ( .A(n_458), .B(n_433), .Y(n_527) );
AOI21xp33_ASAP7_75t_L g528 ( .A1(n_484), .A2(n_425), .B(n_443), .Y(n_528) );
INVx1_ASAP7_75t_SL g529 ( .A(n_457), .Y(n_529) );
OR2x2_ASAP7_75t_L g530 ( .A(n_460), .B(n_445), .Y(n_530) );
AND2x4_ASAP7_75t_L g531 ( .A(n_486), .B(n_427), .Y(n_531) );
AND2x2_ASAP7_75t_L g532 ( .A(n_478), .B(n_433), .Y(n_532) );
INVxp67_ASAP7_75t_L g533 ( .A(n_466), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_454), .B(n_419), .Y(n_534) );
OR2x2_ASAP7_75t_L g535 ( .A(n_460), .B(n_465), .Y(n_535) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_456), .B(n_426), .Y(n_536) );
AOI22xp33_ASAP7_75t_SL g537 ( .A1(n_466), .A2(n_408), .B1(n_415), .B2(n_446), .Y(n_537) );
OR2x2_ASAP7_75t_L g538 ( .A(n_465), .B(n_440), .Y(n_538) );
INVx1_ASAP7_75t_L g539 ( .A(n_451), .Y(n_539) );
NOR2xp33_ASAP7_75t_L g540 ( .A(n_481), .B(n_462), .Y(n_540) );
INVx1_ASAP7_75t_L g541 ( .A(n_452), .Y(n_541) );
INVx1_ASAP7_75t_L g542 ( .A(n_453), .Y(n_542) );
INVx3_ASAP7_75t_L g543 ( .A(n_466), .Y(n_543) );
AND2x2_ASAP7_75t_L g544 ( .A(n_478), .B(n_426), .Y(n_544) );
INVx1_ASAP7_75t_L g545 ( .A(n_455), .Y(n_545) );
OAI22xp5_ASAP7_75t_L g546 ( .A1(n_462), .A2(n_415), .B1(n_404), .B2(n_420), .Y(n_546) );
OAI21xp5_ASAP7_75t_L g547 ( .A1(n_468), .A2(n_507), .B(n_501), .Y(n_547) );
OR2x2_ASAP7_75t_L g548 ( .A(n_491), .B(n_440), .Y(n_548) );
INVx1_ASAP7_75t_L g549 ( .A(n_459), .Y(n_549) );
AND2x2_ASAP7_75t_L g550 ( .A(n_491), .B(n_431), .Y(n_550) );
INVxp67_ASAP7_75t_SL g551 ( .A(n_473), .Y(n_551) );
NAND2xp33_ASAP7_75t_SL g552 ( .A(n_499), .B(n_405), .Y(n_552) );
AOI22xp33_ASAP7_75t_SL g553 ( .A1(n_456), .A2(n_446), .B1(n_427), .B2(n_431), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g554 ( .A(n_463), .B(n_429), .Y(n_554) );
AND2x2_ASAP7_75t_L g555 ( .A(n_497), .B(n_446), .Y(n_555) );
AND2x2_ASAP7_75t_L g556 ( .A(n_497), .B(n_446), .Y(n_556) );
AND2x4_ASAP7_75t_L g557 ( .A(n_496), .B(n_420), .Y(n_557) );
AND2x2_ASAP7_75t_SL g558 ( .A(n_496), .B(n_429), .Y(n_558) );
AOI322xp5_ASAP7_75t_L g559 ( .A1(n_552), .A2(n_471), .A3(n_463), .B1(n_500), .B2(n_505), .C1(n_467), .C2(n_482), .Y(n_559) );
INVx1_ASAP7_75t_SL g560 ( .A(n_523), .Y(n_560) );
OAI22xp33_ASAP7_75t_L g561 ( .A1(n_526), .A2(n_487), .B1(n_471), .B2(n_496), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g562 ( .A(n_517), .B(n_500), .Y(n_562) );
INVx1_ASAP7_75t_L g563 ( .A(n_535), .Y(n_563) );
INVx2_ASAP7_75t_L g564 ( .A(n_548), .Y(n_564) );
INVx1_ASAP7_75t_L g565 ( .A(n_554), .Y(n_565) );
INVx1_ASAP7_75t_L g566 ( .A(n_554), .Y(n_566) );
INVx1_ASAP7_75t_L g567 ( .A(n_515), .Y(n_567) );
OAI211xp5_ASAP7_75t_L g568 ( .A1(n_547), .A2(n_485), .B(n_498), .C(n_504), .Y(n_568) );
INVx2_ASAP7_75t_L g569 ( .A(n_516), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g570 ( .A(n_522), .B(n_505), .Y(n_570) );
OAI222xp33_ASAP7_75t_L g571 ( .A1(n_553), .A2(n_487), .B1(n_464), .B2(n_480), .C1(n_502), .C2(n_494), .Y(n_571) );
INVx1_ASAP7_75t_L g572 ( .A(n_539), .Y(n_572) );
INVxp67_ASAP7_75t_SL g573 ( .A(n_551), .Y(n_573) );
INVx1_ASAP7_75t_L g574 ( .A(n_541), .Y(n_574) );
OAI211xp5_ASAP7_75t_L g575 ( .A1(n_547), .A2(n_490), .B(n_493), .C(n_470), .Y(n_575) );
AOI22xp5_ASAP7_75t_L g576 ( .A1(n_512), .A2(n_474), .B1(n_475), .B2(n_506), .Y(n_576) );
AOI221xp5_ASAP7_75t_L g577 ( .A1(n_528), .A2(n_508), .B1(n_421), .B2(n_509), .C(n_488), .Y(n_577) );
INVx1_ASAP7_75t_SL g578 ( .A(n_523), .Y(n_578) );
OAI221xp5_ASAP7_75t_L g579 ( .A1(n_528), .A2(n_509), .B1(n_487), .B2(n_421), .C(n_488), .Y(n_579) );
INVxp67_ASAP7_75t_L g580 ( .A(n_529), .Y(n_580) );
INVx1_ASAP7_75t_L g581 ( .A(n_542), .Y(n_581) );
INVx1_ASAP7_75t_L g582 ( .A(n_545), .Y(n_582) );
INVx1_ASAP7_75t_SL g583 ( .A(n_529), .Y(n_583) );
NAND2x1_ASAP7_75t_L g584 ( .A(n_543), .B(n_414), .Y(n_584) );
INVx2_ASAP7_75t_L g585 ( .A(n_538), .Y(n_585) );
OAI21xp5_ASAP7_75t_L g586 ( .A1(n_526), .A2(n_424), .B(n_414), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g587 ( .A(n_522), .B(n_492), .Y(n_587) );
OAI22xp33_ASAP7_75t_L g588 ( .A1(n_543), .A2(n_424), .B1(n_450), .B2(n_492), .Y(n_588) );
INVx1_ASAP7_75t_L g589 ( .A(n_549), .Y(n_589) );
NAND2xp5_ASAP7_75t_L g590 ( .A(n_534), .B(n_469), .Y(n_590) );
INVx1_ASAP7_75t_L g591 ( .A(n_530), .Y(n_591) );
OAI22xp5_ASAP7_75t_L g592 ( .A1(n_561), .A2(n_558), .B1(n_527), .B2(n_537), .Y(n_592) );
AOI221x1_ASAP7_75t_L g593 ( .A1(n_569), .A2(n_540), .B1(n_546), .B2(n_534), .C(n_531), .Y(n_593) );
OAI321xp33_ASAP7_75t_L g594 ( .A1(n_561), .A2(n_533), .A3(n_546), .B1(n_513), .B2(n_519), .C(n_511), .Y(n_594) );
OR2x2_ASAP7_75t_L g595 ( .A(n_587), .B(n_519), .Y(n_595) );
INVx1_ASAP7_75t_SL g596 ( .A(n_560), .Y(n_596) );
INVxp67_ASAP7_75t_L g597 ( .A(n_578), .Y(n_597) );
AO32x1_ASAP7_75t_L g598 ( .A1(n_569), .A2(n_510), .A3(n_514), .B1(n_461), .B2(n_469), .Y(n_598) );
AOI22xp5_ASAP7_75t_L g599 ( .A1(n_568), .A2(n_531), .B1(n_557), .B2(n_536), .Y(n_599) );
O2A1O1Ixp33_ASAP7_75t_SL g600 ( .A1(n_571), .A2(n_518), .B(n_521), .C(n_520), .Y(n_600) );
AOI21xp5_ASAP7_75t_L g601 ( .A1(n_586), .A2(n_557), .B(n_511), .Y(n_601) );
OAI21xp33_ASAP7_75t_L g602 ( .A1(n_559), .A2(n_532), .B(n_556), .Y(n_602) );
AOI21xp5_ASAP7_75t_L g603 ( .A1(n_575), .A2(n_555), .B(n_544), .Y(n_603) );
AOI22xp5_ASAP7_75t_L g604 ( .A1(n_563), .A2(n_525), .B1(n_524), .B2(n_550), .Y(n_604) );
NAND3xp33_ASAP7_75t_L g605 ( .A(n_577), .B(n_461), .C(n_424), .Y(n_605) );
INVx2_ASAP7_75t_L g606 ( .A(n_584), .Y(n_606) );
O2A1O1Ixp33_ASAP7_75t_L g607 ( .A1(n_573), .A2(n_450), .B(n_384), .C(n_397), .Y(n_607) );
AOI221xp5_ASAP7_75t_L g608 ( .A1(n_579), .A2(n_447), .B1(n_384), .B2(n_387), .C(n_397), .Y(n_608) );
NOR3xp33_ASAP7_75t_L g609 ( .A(n_573), .B(n_384), .C(n_347), .Y(n_609) );
OAI21xp33_ASAP7_75t_SL g610 ( .A1(n_583), .A2(n_447), .B(n_384), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g611 ( .A(n_565), .B(n_387), .Y(n_611) );
OAI221xp5_ASAP7_75t_L g612 ( .A1(n_592), .A2(n_576), .B1(n_580), .B2(n_566), .C(n_582), .Y(n_612) );
NOR2xp67_ASAP7_75t_SL g613 ( .A(n_594), .B(n_349), .Y(n_613) );
NAND4xp75_ASAP7_75t_L g614 ( .A(n_593), .B(n_591), .C(n_589), .D(n_581), .Y(n_614) );
OAI311xp33_ASAP7_75t_L g615 ( .A1(n_602), .A2(n_590), .A3(n_570), .B1(n_562), .C1(n_574), .Y(n_615) );
NOR2xp33_ASAP7_75t_R g616 ( .A(n_596), .B(n_585), .Y(n_616) );
NOR4xp75_ASAP7_75t_L g617 ( .A(n_600), .B(n_597), .C(n_611), .D(n_598), .Y(n_617) );
NAND2xp5_ASAP7_75t_L g618 ( .A(n_603), .B(n_572), .Y(n_618) );
AOI221x1_ASAP7_75t_SL g619 ( .A1(n_605), .A2(n_585), .B1(n_588), .B2(n_564), .C(n_567), .Y(n_619) );
AOI21xp5_ASAP7_75t_L g620 ( .A1(n_601), .A2(n_588), .B(n_564), .Y(n_620) );
INVx3_ASAP7_75t_L g621 ( .A(n_606), .Y(n_621) );
AOI21x1_ASAP7_75t_L g622 ( .A1(n_598), .A2(n_595), .B(n_349), .Y(n_622) );
NAND4xp75_ASAP7_75t_L g623 ( .A(n_620), .B(n_610), .C(n_599), .D(n_608), .Y(n_623) );
INVx2_ASAP7_75t_SL g624 ( .A(n_616), .Y(n_624) );
OAI222xp33_ASAP7_75t_R g625 ( .A1(n_619), .A2(n_604), .B1(n_598), .B2(n_609), .C1(n_607), .C2(n_387), .Y(n_625) );
NOR3xp33_ASAP7_75t_L g626 ( .A(n_612), .B(n_347), .C(n_349), .Y(n_626) );
INVx1_ASAP7_75t_L g627 ( .A(n_618), .Y(n_627) );
NAND4xp25_ASAP7_75t_SL g628 ( .A(n_617), .B(n_344), .C(n_385), .D(n_351), .Y(n_628) );
INVx1_ASAP7_75t_L g629 ( .A(n_624), .Y(n_629) );
NAND5xp2_ASAP7_75t_L g630 ( .A(n_627), .B(n_622), .C(n_613), .D(n_615), .E(n_614), .Y(n_630) );
INVx2_ASAP7_75t_L g631 ( .A(n_623), .Y(n_631) );
NOR2xp33_ASAP7_75t_L g632 ( .A(n_629), .B(n_628), .Y(n_632) );
XNOR2xp5_ASAP7_75t_L g633 ( .A(n_631), .B(n_626), .Y(n_633) );
XOR2x1_ASAP7_75t_L g634 ( .A(n_633), .B(n_631), .Y(n_634) );
XNOR2xp5_ASAP7_75t_L g635 ( .A(n_632), .B(n_625), .Y(n_635) );
OAI22xp5_ASAP7_75t_SL g636 ( .A1(n_635), .A2(n_630), .B1(n_621), .B2(n_385), .Y(n_636) );
OAI21x1_ASAP7_75t_L g637 ( .A1(n_636), .A2(n_634), .B(n_621), .Y(n_637) );
AOI21xp5_ASAP7_75t_L g638 ( .A1(n_637), .A2(n_385), .B(n_344), .Y(n_638) );
AO21x2_ASAP7_75t_L g639 ( .A1(n_638), .A2(n_344), .B(n_385), .Y(n_639) );
AOI22xp5_ASAP7_75t_L g640 ( .A1(n_639), .A2(n_385), .B1(n_624), .B2(n_629), .Y(n_640) );
endmodule