module fake_netlist_1_3936_n_34 (n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_34);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_34;
wire n_20;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_30;
wire n_33;
wire n_18;
wire n_32;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_27;
AND2x2_ASAP7_75t_L g11 ( .A(n_0), .B(n_5), .Y(n_11) );
NOR2x1_ASAP7_75t_L g12 ( .A(n_1), .B(n_9), .Y(n_12) );
INVx3_ASAP7_75t_L g13 ( .A(n_5), .Y(n_13) );
INVx2_ASAP7_75t_L g14 ( .A(n_8), .Y(n_14) );
NOR2x1_ASAP7_75t_L g15 ( .A(n_1), .B(n_2), .Y(n_15) );
NAND2xp5_ASAP7_75t_L g16 ( .A(n_13), .B(n_0), .Y(n_16) );
INVx2_ASAP7_75t_L g17 ( .A(n_13), .Y(n_17) );
INVx2_ASAP7_75t_SL g18 ( .A(n_15), .Y(n_18) );
BUFx2_ASAP7_75t_R g19 ( .A(n_16), .Y(n_19) );
AOI22xp33_ASAP7_75t_SL g20 ( .A1(n_18), .A2(n_16), .B1(n_11), .B2(n_17), .Y(n_20) );
AND2x2_ASAP7_75t_L g21 ( .A(n_20), .B(n_12), .Y(n_21) );
BUFx6f_ASAP7_75t_L g22 ( .A(n_19), .Y(n_22) );
AND2x2_ASAP7_75t_L g23 ( .A(n_21), .B(n_19), .Y(n_23) );
INVx2_ASAP7_75t_L g24 ( .A(n_21), .Y(n_24) );
NAND2xp5_ASAP7_75t_SL g25 ( .A(n_23), .B(n_22), .Y(n_25) );
HB1xp67_ASAP7_75t_L g26 ( .A(n_24), .Y(n_26) );
AOI21xp5_ASAP7_75t_L g27 ( .A1(n_25), .A2(n_14), .B(n_12), .Y(n_27) );
OA22x2_ASAP7_75t_L g28 ( .A1(n_26), .A2(n_22), .B1(n_3), .B2(n_4), .Y(n_28) );
NAND2xp5_ASAP7_75t_L g29 ( .A(n_28), .B(n_22), .Y(n_29) );
OAI211xp5_ASAP7_75t_SL g30 ( .A1(n_27), .A2(n_22), .B(n_3), .C(n_4), .Y(n_30) );
NAND3xp33_ASAP7_75t_L g31 ( .A(n_29), .B(n_22), .C(n_6), .Y(n_31) );
INVx1_ASAP7_75t_L g32 ( .A(n_30), .Y(n_32) );
AOI211xp5_ASAP7_75t_SL g33 ( .A1(n_32), .A2(n_2), .B(n_6), .C(n_7), .Y(n_33) );
AOI22xp33_ASAP7_75t_L g34 ( .A1(n_33), .A2(n_31), .B1(n_10), .B2(n_7), .Y(n_34) );
endmodule