module fake_jpeg_14371_n_133 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_133);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_133;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_131;
wire n_56;
wire n_79;
wire n_12;
wire n_132;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_4),
.Y(n_11)
);

BUFx3_ASAP7_75t_L g12 ( 
.A(n_2),
.Y(n_12)
);

NOR2xp33_ASAP7_75t_L g13 ( 
.A(n_3),
.B(n_4),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_6),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_5),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_1),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_0),
.B(n_2),
.Y(n_17)
);

CKINVDCx14_ASAP7_75t_R g18 ( 
.A(n_7),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_0),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_10),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_6),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_3),
.Y(n_26)
);

INVx13_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_24),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_28),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_17),
.B(n_1),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_29),
.B(n_30),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_11),
.B(n_7),
.Y(n_30)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_31),
.Y(n_68)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_23),
.Y(n_32)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_32),
.Y(n_50)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_33),
.Y(n_61)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_24),
.Y(n_34)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_34),
.Y(n_71)
);

INVx1_ASAP7_75t_SL g35 ( 
.A(n_27),
.Y(n_35)
);

CKINVDCx14_ASAP7_75t_R g57 ( 
.A(n_35),
.Y(n_57)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_24),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_36),
.B(n_37),
.Y(n_51)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_20),
.Y(n_37)
);

INVxp67_ASAP7_75t_L g38 ( 
.A(n_13),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_38),
.B(n_41),
.Y(n_65)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_20),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_39),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_SL g40 ( 
.A1(n_23),
.A2(n_1),
.B1(n_8),
.B2(n_9),
.Y(n_40)
);

AOI21xp5_ASAP7_75t_L g54 ( 
.A1(n_40),
.A2(n_16),
.B(n_19),
.Y(n_54)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_21),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_11),
.B(n_8),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_42),
.B(n_43),
.Y(n_69)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_21),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_21),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_44),
.B(n_45),
.Y(n_70)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_27),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_14),
.B(n_9),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_46),
.B(n_47),
.Y(n_72)
);

BUFx4f_ASAP7_75t_SL g47 ( 
.A(n_18),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_14),
.B(n_15),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g55 ( 
.A(n_48),
.B(n_15),
.Y(n_55)
);

NOR2x1_ASAP7_75t_L g52 ( 
.A(n_47),
.B(n_16),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_52),
.B(n_55),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_54),
.B(n_63),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_L g56 ( 
.A1(n_37),
.A2(n_36),
.B1(n_39),
.B2(n_34),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_56),
.A2(n_62),
.B1(n_57),
.B2(n_49),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g58 ( 
.A(n_38),
.B(n_19),
.C(n_26),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_58),
.B(n_53),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_33),
.B(n_26),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_60),
.B(n_66),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_35),
.A2(n_22),
.B1(n_25),
.B2(n_28),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_SL g63 ( 
.A(n_47),
.B(n_22),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_43),
.B(n_25),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_64),
.B(n_67),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_29),
.B(n_32),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g67 ( 
.A(n_38),
.B(n_48),
.Y(n_67)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_59),
.Y(n_73)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_73),
.Y(n_92)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_71),
.Y(n_74)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_74),
.Y(n_103)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_59),
.Y(n_78)
);

INVx2_ASAP7_75t_SL g94 ( 
.A(n_78),
.Y(n_94)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_71),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_79),
.B(n_86),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_81),
.B(n_82),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_67),
.B(n_58),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_60),
.A2(n_66),
.B1(n_50),
.B2(n_49),
.Y(n_83)
);

OAI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_83),
.A2(n_89),
.B1(n_90),
.B2(n_79),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_55),
.B(n_63),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_84),
.B(n_85),
.Y(n_97)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_70),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_51),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_72),
.B(n_65),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_87),
.B(n_86),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_88),
.A2(n_90),
.B1(n_74),
.B2(n_91),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_50),
.A2(n_64),
.B1(n_54),
.B2(n_68),
.Y(n_89)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_61),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_69),
.A2(n_68),
.B1(n_61),
.B2(n_59),
.Y(n_91)
);

OA21x2_ASAP7_75t_L g93 ( 
.A1(n_91),
.A2(n_52),
.B(n_89),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_93),
.B(n_105),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_SL g95 ( 
.A1(n_83),
.A2(n_52),
.B(n_75),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_L g112 ( 
.A1(n_95),
.A2(n_96),
.B(n_100),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_SL g96 ( 
.A1(n_75),
.A2(n_85),
.B(n_80),
.Y(n_96)
);

OR2x2_ASAP7_75t_L g100 ( 
.A(n_76),
.B(n_77),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_100),
.B(n_102),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_101),
.A2(n_104),
.B1(n_78),
.B2(n_94),
.Y(n_111)
);

XOR2xp5_ASAP7_75t_L g105 ( 
.A(n_76),
.B(n_73),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_99),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g120 ( 
.A(n_107),
.B(n_109),
.Y(n_120)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_103),
.Y(n_108)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_108),
.Y(n_116)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_99),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_L g117 ( 
.A1(n_111),
.A2(n_113),
.B(n_114),
.Y(n_117)
);

XOR2xp5_ASAP7_75t_L g119 ( 
.A(n_112),
.B(n_94),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_98),
.B(n_102),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_97),
.B(n_96),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_110),
.A2(n_93),
.B1(n_105),
.B2(n_95),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_L g125 ( 
.A1(n_115),
.A2(n_92),
.B(n_119),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_L g118 ( 
.A(n_112),
.B(n_93),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_106),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_121),
.B(n_110),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_122),
.B(n_123),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_L g123 ( 
.A(n_118),
.B(n_111),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_120),
.A2(n_92),
.B1(n_94),
.B2(n_117),
.Y(n_124)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_124),
.Y(n_128)
);

HB1xp67_ASAP7_75t_L g126 ( 
.A(n_125),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_127),
.B(n_116),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_129),
.B(n_130),
.Y(n_131)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_128),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_131),
.B(n_126),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_132),
.B(n_123),
.Y(n_133)
);


endmodule