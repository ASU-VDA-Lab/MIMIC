module fake_netlist_1_69_n_676 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_6, n_4, n_40, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_676);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_6;
input n_4;
input n_40;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_676;
wire n_117;
wire n_663;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_85;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_77;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_90;
wire n_357;
wire n_653;
wire n_260;
wire n_78;
wire n_539;
wire n_201;
wire n_197;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_487;
wire n_451;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_84;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_132;
wire n_109;
wire n_99;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g77 ( .A(n_22), .Y(n_77) );
INVx1_ASAP7_75t_L g78 ( .A(n_25), .Y(n_78) );
INVx1_ASAP7_75t_L g79 ( .A(n_57), .Y(n_79) );
CKINVDCx5p33_ASAP7_75t_R g80 ( .A(n_53), .Y(n_80) );
INVx1_ASAP7_75t_L g81 ( .A(n_70), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_7), .Y(n_82) );
INVxp33_ASAP7_75t_L g83 ( .A(n_60), .Y(n_83) );
INVxp67_ASAP7_75t_SL g84 ( .A(n_38), .Y(n_84) );
CKINVDCx5p33_ASAP7_75t_R g85 ( .A(n_3), .Y(n_85) );
INVx1_ASAP7_75t_SL g86 ( .A(n_31), .Y(n_86) );
INVx2_ASAP7_75t_L g87 ( .A(n_64), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_5), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_59), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_14), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_42), .Y(n_91) );
CKINVDCx20_ASAP7_75t_R g92 ( .A(n_17), .Y(n_92) );
BUFx2_ASAP7_75t_L g93 ( .A(n_41), .Y(n_93) );
INVx2_ASAP7_75t_L g94 ( .A(n_26), .Y(n_94) );
CKINVDCx5p33_ASAP7_75t_R g95 ( .A(n_32), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_47), .Y(n_96) );
CKINVDCx5p33_ASAP7_75t_R g97 ( .A(n_46), .Y(n_97) );
HB1xp67_ASAP7_75t_L g98 ( .A(n_58), .Y(n_98) );
CKINVDCx20_ASAP7_75t_R g99 ( .A(n_6), .Y(n_99) );
INVx1_ASAP7_75t_SL g100 ( .A(n_5), .Y(n_100) );
CKINVDCx16_ASAP7_75t_R g101 ( .A(n_40), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_1), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_21), .Y(n_103) );
HB1xp67_ASAP7_75t_L g104 ( .A(n_69), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_71), .Y(n_105) );
CKINVDCx14_ASAP7_75t_R g106 ( .A(n_3), .Y(n_106) );
INVx2_ASAP7_75t_L g107 ( .A(n_7), .Y(n_107) );
NOR2xp33_ASAP7_75t_L g108 ( .A(n_61), .B(n_37), .Y(n_108) );
INVxp33_ASAP7_75t_L g109 ( .A(n_15), .Y(n_109) );
INVxp67_ASAP7_75t_SL g110 ( .A(n_15), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_52), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_48), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_10), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_76), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_74), .Y(n_115) );
CKINVDCx16_ASAP7_75t_R g116 ( .A(n_34), .Y(n_116) );
CKINVDCx5p33_ASAP7_75t_R g117 ( .A(n_6), .Y(n_117) );
INVxp67_ASAP7_75t_SL g118 ( .A(n_4), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_68), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_13), .Y(n_120) );
INVxp33_ASAP7_75t_SL g121 ( .A(n_43), .Y(n_121) );
CKINVDCx16_ASAP7_75t_R g122 ( .A(n_23), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_62), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_18), .Y(n_124) );
CKINVDCx20_ASAP7_75t_R g125 ( .A(n_122), .Y(n_125) );
NAND2xp5_ASAP7_75t_L g126 ( .A(n_93), .B(n_98), .Y(n_126) );
INVx3_ASAP7_75t_L g127 ( .A(n_107), .Y(n_127) );
CKINVDCx20_ASAP7_75t_R g128 ( .A(n_122), .Y(n_128) );
INVx1_ASAP7_75t_L g129 ( .A(n_107), .Y(n_129) );
INVx1_ASAP7_75t_L g130 ( .A(n_107), .Y(n_130) );
INVx1_ASAP7_75t_L g131 ( .A(n_78), .Y(n_131) );
BUFx3_ASAP7_75t_L g132 ( .A(n_93), .Y(n_132) );
NOR2xp33_ASAP7_75t_L g133 ( .A(n_104), .B(n_0), .Y(n_133) );
BUFx6f_ASAP7_75t_L g134 ( .A(n_87), .Y(n_134) );
INVx1_ASAP7_75t_L g135 ( .A(n_78), .Y(n_135) );
BUFx3_ASAP7_75t_L g136 ( .A(n_87), .Y(n_136) );
BUFx6f_ASAP7_75t_L g137 ( .A(n_87), .Y(n_137) );
OAI22xp5_ASAP7_75t_L g138 ( .A1(n_106), .A2(n_0), .B1(n_1), .B2(n_2), .Y(n_138) );
INVxp67_ASAP7_75t_L g139 ( .A(n_77), .Y(n_139) );
INVx1_ASAP7_75t_SL g140 ( .A(n_101), .Y(n_140) );
INVx1_ASAP7_75t_L g141 ( .A(n_79), .Y(n_141) );
CKINVDCx5p33_ASAP7_75t_R g142 ( .A(n_101), .Y(n_142) );
INVx1_ASAP7_75t_L g143 ( .A(n_79), .Y(n_143) );
INVx1_ASAP7_75t_L g144 ( .A(n_81), .Y(n_144) );
CKINVDCx5p33_ASAP7_75t_R g145 ( .A(n_116), .Y(n_145) );
BUFx2_ASAP7_75t_L g146 ( .A(n_116), .Y(n_146) );
AND2x6_ASAP7_75t_L g147 ( .A(n_94), .B(n_29), .Y(n_147) );
HB1xp67_ASAP7_75t_L g148 ( .A(n_77), .Y(n_148) );
CKINVDCx5p33_ASAP7_75t_R g149 ( .A(n_85), .Y(n_149) );
INVx1_ASAP7_75t_L g150 ( .A(n_81), .Y(n_150) );
HB1xp67_ASAP7_75t_L g151 ( .A(n_109), .Y(n_151) );
NAND2xp5_ASAP7_75t_L g152 ( .A(n_82), .B(n_2), .Y(n_152) );
NAND2xp5_ASAP7_75t_L g153 ( .A(n_82), .B(n_4), .Y(n_153) );
CKINVDCx5p33_ASAP7_75t_R g154 ( .A(n_117), .Y(n_154) );
INVx1_ASAP7_75t_L g155 ( .A(n_89), .Y(n_155) );
INVx1_ASAP7_75t_L g156 ( .A(n_89), .Y(n_156) );
AND2x2_ASAP7_75t_L g157 ( .A(n_83), .B(n_8), .Y(n_157) );
CKINVDCx5p33_ASAP7_75t_R g158 ( .A(n_121), .Y(n_158) );
HB1xp67_ASAP7_75t_L g159 ( .A(n_88), .Y(n_159) );
INVx2_ASAP7_75t_L g160 ( .A(n_94), .Y(n_160) );
CKINVDCx5p33_ASAP7_75t_R g161 ( .A(n_80), .Y(n_161) );
HB1xp67_ASAP7_75t_L g162 ( .A(n_88), .Y(n_162) );
INVx1_ASAP7_75t_L g163 ( .A(n_91), .Y(n_163) );
CKINVDCx5p33_ASAP7_75t_R g164 ( .A(n_95), .Y(n_164) );
INVx1_ASAP7_75t_L g165 ( .A(n_91), .Y(n_165) );
INVx1_ASAP7_75t_L g166 ( .A(n_96), .Y(n_166) );
INVx1_ASAP7_75t_L g167 ( .A(n_96), .Y(n_167) );
NOR2xp33_ASAP7_75t_L g168 ( .A(n_132), .B(n_112), .Y(n_168) );
OR2x2_ASAP7_75t_L g169 ( .A(n_151), .B(n_118), .Y(n_169) );
INVx1_ASAP7_75t_L g170 ( .A(n_136), .Y(n_170) );
AND2x4_ASAP7_75t_L g171 ( .A(n_132), .B(n_124), .Y(n_171) );
AND2x4_ASAP7_75t_L g172 ( .A(n_132), .B(n_148), .Y(n_172) );
INVx1_ASAP7_75t_L g173 ( .A(n_136), .Y(n_173) );
NOR2xp33_ASAP7_75t_SL g174 ( .A(n_146), .B(n_140), .Y(n_174) );
INVx1_ASAP7_75t_L g175 ( .A(n_136), .Y(n_175) );
INVx1_ASAP7_75t_L g176 ( .A(n_148), .Y(n_176) );
AND2x4_ASAP7_75t_L g177 ( .A(n_126), .B(n_124), .Y(n_177) );
AOI22xp5_ASAP7_75t_L g178 ( .A1(n_146), .A2(n_103), .B1(n_120), .B2(n_90), .Y(n_178) );
NAND3xp33_ASAP7_75t_L g179 ( .A(n_159), .B(n_90), .C(n_120), .Y(n_179) );
AOI22xp33_ASAP7_75t_L g180 ( .A1(n_162), .A2(n_102), .B1(n_103), .B2(n_113), .Y(n_180) );
BUFx6f_ASAP7_75t_L g181 ( .A(n_134), .Y(n_181) );
CKINVDCx5p33_ASAP7_75t_R g182 ( .A(n_142), .Y(n_182) );
AO22x2_ASAP7_75t_L g183 ( .A1(n_138), .A2(n_118), .B1(n_123), .B2(n_119), .Y(n_183) );
INVx8_ASAP7_75t_L g184 ( .A(n_147), .Y(n_184) );
INVx2_ASAP7_75t_L g185 ( .A(n_134), .Y(n_185) );
INVx1_ASAP7_75t_L g186 ( .A(n_131), .Y(n_186) );
INVx3_ASAP7_75t_L g187 ( .A(n_127), .Y(n_187) );
NOR2xp33_ASAP7_75t_L g188 ( .A(n_126), .B(n_123), .Y(n_188) );
NAND2x1p5_ASAP7_75t_L g189 ( .A(n_140), .B(n_157), .Y(n_189) );
INVx1_ASAP7_75t_L g190 ( .A(n_131), .Y(n_190) );
OAI22xp5_ASAP7_75t_L g191 ( .A1(n_145), .A2(n_102), .B1(n_113), .B2(n_110), .Y(n_191) );
INVx2_ASAP7_75t_L g192 ( .A(n_134), .Y(n_192) );
INVx6_ASAP7_75t_L g193 ( .A(n_134), .Y(n_193) );
INVx1_ASAP7_75t_L g194 ( .A(n_135), .Y(n_194) );
INVx4_ASAP7_75t_L g195 ( .A(n_147), .Y(n_195) );
BUFx6f_ASAP7_75t_L g196 ( .A(n_134), .Y(n_196) );
AOI22x1_ASAP7_75t_L g197 ( .A1(n_160), .A2(n_94), .B1(n_115), .B2(n_114), .Y(n_197) );
INVx1_ASAP7_75t_L g198 ( .A(n_135), .Y(n_198) );
INVxp33_ASAP7_75t_L g199 ( .A(n_157), .Y(n_199) );
BUFx6f_ASAP7_75t_L g200 ( .A(n_134), .Y(n_200) );
INVx2_ASAP7_75t_L g201 ( .A(n_137), .Y(n_201) );
AND2x4_ASAP7_75t_L g202 ( .A(n_139), .B(n_119), .Y(n_202) );
BUFx3_ASAP7_75t_L g203 ( .A(n_147), .Y(n_203) );
INVx1_ASAP7_75t_L g204 ( .A(n_141), .Y(n_204) );
AND2x6_ASAP7_75t_L g205 ( .A(n_141), .B(n_105), .Y(n_205) );
AND2x4_ASAP7_75t_L g206 ( .A(n_139), .B(n_115), .Y(n_206) );
AND2x2_ASAP7_75t_L g207 ( .A(n_143), .B(n_100), .Y(n_207) );
INVx1_ASAP7_75t_L g208 ( .A(n_143), .Y(n_208) );
AND2x2_ASAP7_75t_L g209 ( .A(n_144), .B(n_100), .Y(n_209) );
AND2x4_ASAP7_75t_L g210 ( .A(n_167), .B(n_114), .Y(n_210) );
OAI22xp5_ASAP7_75t_L g211 ( .A1(n_149), .A2(n_99), .B1(n_92), .B2(n_86), .Y(n_211) );
INVxp33_ASAP7_75t_L g212 ( .A(n_133), .Y(n_212) );
BUFx6f_ASAP7_75t_L g213 ( .A(n_137), .Y(n_213) );
INVx2_ASAP7_75t_L g214 ( .A(n_137), .Y(n_214) );
BUFx2_ASAP7_75t_L g215 ( .A(n_154), .Y(n_215) );
BUFx6f_ASAP7_75t_L g216 ( .A(n_137), .Y(n_216) );
INVx1_ASAP7_75t_L g217 ( .A(n_144), .Y(n_217) );
INVx2_ASAP7_75t_L g218 ( .A(n_137), .Y(n_218) );
INVx1_ASAP7_75t_L g219 ( .A(n_150), .Y(n_219) );
INVxp33_ASAP7_75t_L g220 ( .A(n_152), .Y(n_220) );
AOI22xp33_ASAP7_75t_L g221 ( .A1(n_150), .A2(n_111), .B1(n_105), .B2(n_112), .Y(n_221) );
BUFx2_ASAP7_75t_L g222 ( .A(n_161), .Y(n_222) );
INVxp67_ASAP7_75t_L g223 ( .A(n_164), .Y(n_223) );
INVx3_ASAP7_75t_L g224 ( .A(n_127), .Y(n_224) );
BUFx3_ASAP7_75t_L g225 ( .A(n_147), .Y(n_225) );
INVx1_ASAP7_75t_L g226 ( .A(n_155), .Y(n_226) );
AOI22xp33_ASAP7_75t_L g227 ( .A1(n_155), .A2(n_111), .B1(n_86), .B2(n_84), .Y(n_227) );
NAND2xp5_ASAP7_75t_SL g228 ( .A(n_156), .B(n_97), .Y(n_228) );
AND2x6_ASAP7_75t_L g229 ( .A(n_156), .B(n_108), .Y(n_229) );
CKINVDCx16_ASAP7_75t_R g230 ( .A(n_125), .Y(n_230) );
BUFx10_ASAP7_75t_L g231 ( .A(n_172), .Y(n_231) );
INVx1_ASAP7_75t_SL g232 ( .A(n_172), .Y(n_232) );
INVx1_ASAP7_75t_SL g233 ( .A(n_172), .Y(n_233) );
BUFx6f_ASAP7_75t_L g234 ( .A(n_203), .Y(n_234) );
INVx1_ASAP7_75t_L g235 ( .A(n_187), .Y(n_235) );
NAND2xp5_ASAP7_75t_SL g236 ( .A(n_195), .B(n_167), .Y(n_236) );
CKINVDCx5p33_ASAP7_75t_R g237 ( .A(n_230), .Y(n_237) );
INVx2_ASAP7_75t_L g238 ( .A(n_185), .Y(n_238) );
INVx1_ASAP7_75t_SL g239 ( .A(n_215), .Y(n_239) );
A2O1A1Ixp33_ASAP7_75t_L g240 ( .A1(n_188), .A2(n_166), .B(n_165), .C(n_163), .Y(n_240) );
BUFx4f_ASAP7_75t_SL g241 ( .A(n_215), .Y(n_241) );
AOI22xp5_ASAP7_75t_L g242 ( .A1(n_176), .A2(n_158), .B1(n_138), .B2(n_128), .Y(n_242) );
BUFx6f_ASAP7_75t_L g243 ( .A(n_203), .Y(n_243) );
NOR2xp33_ASAP7_75t_R g244 ( .A(n_182), .B(n_147), .Y(n_244) );
NAND2xp5_ASAP7_75t_L g245 ( .A(n_220), .B(n_166), .Y(n_245) );
AND2x4_ASAP7_75t_L g246 ( .A(n_171), .B(n_152), .Y(n_246) );
AOI221xp5_ASAP7_75t_L g247 ( .A1(n_183), .A2(n_165), .B1(n_163), .B2(n_153), .C(n_129), .Y(n_247) );
INVx1_ASAP7_75t_L g248 ( .A(n_187), .Y(n_248) );
CKINVDCx5p33_ASAP7_75t_R g249 ( .A(n_222), .Y(n_249) );
CKINVDCx5p33_ASAP7_75t_R g250 ( .A(n_182), .Y(n_250) );
BUFx6f_ASAP7_75t_L g251 ( .A(n_225), .Y(n_251) );
INVx3_ASAP7_75t_L g252 ( .A(n_187), .Y(n_252) );
INVx1_ASAP7_75t_L g253 ( .A(n_224), .Y(n_253) );
BUFx3_ASAP7_75t_L g254 ( .A(n_184), .Y(n_254) );
INVx1_ASAP7_75t_L g255 ( .A(n_224), .Y(n_255) );
INVx3_ASAP7_75t_L g256 ( .A(n_224), .Y(n_256) );
INVx3_ASAP7_75t_L g257 ( .A(n_210), .Y(n_257) );
INVx1_ASAP7_75t_L g258 ( .A(n_220), .Y(n_258) );
INVx1_ASAP7_75t_L g259 ( .A(n_207), .Y(n_259) );
NOR2xp67_ASAP7_75t_L g260 ( .A(n_223), .B(n_127), .Y(n_260) );
HB1xp67_ASAP7_75t_L g261 ( .A(n_189), .Y(n_261) );
INVx2_ASAP7_75t_L g262 ( .A(n_185), .Y(n_262) );
INVx8_ASAP7_75t_L g263 ( .A(n_184), .Y(n_263) );
NAND2xp5_ASAP7_75t_SL g264 ( .A(n_195), .B(n_137), .Y(n_264) );
NAND2xp5_ASAP7_75t_SL g265 ( .A(n_195), .B(n_153), .Y(n_265) );
BUFx4f_ASAP7_75t_L g266 ( .A(n_189), .Y(n_266) );
A2O1A1Ixp33_ASAP7_75t_L g267 ( .A1(n_177), .A2(n_160), .B(n_130), .C(n_129), .Y(n_267) );
INVx1_ASAP7_75t_L g268 ( .A(n_207), .Y(n_268) );
INVx1_ASAP7_75t_L g269 ( .A(n_209), .Y(n_269) );
NAND2xp33_ASAP7_75t_SL g270 ( .A(n_199), .B(n_160), .Y(n_270) );
HB1xp67_ASAP7_75t_L g271 ( .A(n_209), .Y(n_271) );
NOR3xp33_ASAP7_75t_SL g272 ( .A(n_211), .B(n_130), .C(n_9), .Y(n_272) );
OAI21xp33_ASAP7_75t_SL g273 ( .A1(n_168), .A2(n_127), .B(n_147), .Y(n_273) );
BUFx12f_ASAP7_75t_SL g274 ( .A(n_177), .Y(n_274) );
NAND2xp5_ASAP7_75t_L g275 ( .A(n_202), .B(n_147), .Y(n_275) );
INVx2_ASAP7_75t_L g276 ( .A(n_192), .Y(n_276) );
INVx1_ASAP7_75t_L g277 ( .A(n_210), .Y(n_277) );
INVx2_ASAP7_75t_L g278 ( .A(n_192), .Y(n_278) );
BUFx2_ASAP7_75t_L g279 ( .A(n_169), .Y(n_279) );
NOR2xp33_ASAP7_75t_L g280 ( .A(n_212), .B(n_147), .Y(n_280) );
AND2x2_ASAP7_75t_L g281 ( .A(n_177), .B(n_8), .Y(n_281) );
NOR2xp33_ASAP7_75t_R g282 ( .A(n_174), .B(n_9), .Y(n_282) );
INVx6_ASAP7_75t_L g283 ( .A(n_171), .Y(n_283) );
CKINVDCx5p33_ASAP7_75t_R g284 ( .A(n_191), .Y(n_284) );
NAND2x1p5_ASAP7_75t_L g285 ( .A(n_171), .B(n_10), .Y(n_285) );
BUFx2_ASAP7_75t_L g286 ( .A(n_169), .Y(n_286) );
NOR2xp33_ASAP7_75t_L g287 ( .A(n_212), .B(n_35), .Y(n_287) );
AND2x4_ASAP7_75t_L g288 ( .A(n_202), .B(n_11), .Y(n_288) );
AOI22xp5_ASAP7_75t_L g289 ( .A1(n_199), .A2(n_11), .B1(n_12), .B2(n_13), .Y(n_289) );
BUFx3_ASAP7_75t_L g290 ( .A(n_184), .Y(n_290) );
BUFx2_ASAP7_75t_L g291 ( .A(n_205), .Y(n_291) );
INVx1_ASAP7_75t_L g292 ( .A(n_210), .Y(n_292) );
INVx2_ASAP7_75t_L g293 ( .A(n_201), .Y(n_293) );
NAND2xp5_ASAP7_75t_L g294 ( .A(n_202), .B(n_12), .Y(n_294) );
AOI22xp5_ASAP7_75t_L g295 ( .A1(n_178), .A2(n_14), .B1(n_16), .B2(n_17), .Y(n_295) );
NAND2xp5_ASAP7_75t_L g296 ( .A(n_206), .B(n_16), .Y(n_296) );
AND2x4_ASAP7_75t_L g297 ( .A(n_206), .B(n_18), .Y(n_297) );
NAND2xp5_ASAP7_75t_L g298 ( .A(n_246), .B(n_206), .Y(n_298) );
HB1xp67_ASAP7_75t_L g299 ( .A(n_239), .Y(n_299) );
OR2x6_ASAP7_75t_SL g300 ( .A(n_249), .B(n_179), .Y(n_300) );
INVx1_ASAP7_75t_L g301 ( .A(n_277), .Y(n_301) );
AOI21xp33_ASAP7_75t_SL g302 ( .A1(n_249), .A2(n_183), .B(n_180), .Y(n_302) );
AOI21x1_ASAP7_75t_L g303 ( .A1(n_264), .A2(n_204), .B(n_186), .Y(n_303) );
OAI22xp5_ASAP7_75t_L g304 ( .A1(n_288), .A2(n_221), .B1(n_183), .B2(n_227), .Y(n_304) );
INVx3_ASAP7_75t_L g305 ( .A(n_252), .Y(n_305) );
BUFx6f_ASAP7_75t_L g306 ( .A(n_263), .Y(n_306) );
INVx3_ASAP7_75t_L g307 ( .A(n_252), .Y(n_307) );
AO21x1_ASAP7_75t_L g308 ( .A1(n_270), .A2(n_201), .B(n_214), .Y(n_308) );
AND2x4_ASAP7_75t_L g309 ( .A(n_288), .B(n_225), .Y(n_309) );
BUFx6f_ASAP7_75t_L g310 ( .A(n_263), .Y(n_310) );
BUFx3_ASAP7_75t_L g311 ( .A(n_231), .Y(n_311) );
AOI21xp5_ASAP7_75t_L g312 ( .A1(n_265), .A2(n_184), .B(n_228), .Y(n_312) );
BUFx3_ASAP7_75t_L g313 ( .A(n_263), .Y(n_313) );
INVx1_ASAP7_75t_L g314 ( .A(n_292), .Y(n_314) );
INVx1_ASAP7_75t_L g315 ( .A(n_257), .Y(n_315) );
AOI22xp5_ASAP7_75t_L g316 ( .A1(n_288), .A2(n_183), .B1(n_205), .B2(n_226), .Y(n_316) );
BUFx6f_ASAP7_75t_L g317 ( .A(n_234), .Y(n_317) );
INVx2_ASAP7_75t_L g318 ( .A(n_235), .Y(n_318) );
INVx1_ASAP7_75t_L g319 ( .A(n_257), .Y(n_319) );
INVx3_ASAP7_75t_L g320 ( .A(n_256), .Y(n_320) );
BUFx3_ASAP7_75t_L g321 ( .A(n_254), .Y(n_321) );
AOI21xp5_ASAP7_75t_L g322 ( .A1(n_265), .A2(n_228), .B(n_190), .Y(n_322) );
AND2x2_ASAP7_75t_L g323 ( .A(n_258), .B(n_198), .Y(n_323) );
A2O1A1Ixp33_ASAP7_75t_L g324 ( .A1(n_280), .A2(n_194), .B(n_219), .C(n_208), .Y(n_324) );
INVx1_ASAP7_75t_L g325 ( .A(n_248), .Y(n_325) );
AND2x2_ASAP7_75t_L g326 ( .A(n_271), .B(n_217), .Y(n_326) );
INVx2_ASAP7_75t_L g327 ( .A(n_253), .Y(n_327) );
BUFx3_ASAP7_75t_L g328 ( .A(n_254), .Y(n_328) );
OAI22xp5_ASAP7_75t_L g329 ( .A1(n_297), .A2(n_170), .B1(n_173), .B2(n_175), .Y(n_329) );
BUFx6f_ASAP7_75t_L g330 ( .A(n_234), .Y(n_330) );
INVx1_ASAP7_75t_L g331 ( .A(n_255), .Y(n_331) );
OAI22xp5_ASAP7_75t_L g332 ( .A1(n_297), .A2(n_197), .B1(n_205), .B2(n_193), .Y(n_332) );
AND2x4_ASAP7_75t_L g333 ( .A(n_297), .B(n_205), .Y(n_333) );
INVx3_ASAP7_75t_SL g334 ( .A(n_231), .Y(n_334) );
BUFx12f_ASAP7_75t_L g335 ( .A(n_237), .Y(n_335) );
INVx2_ASAP7_75t_L g336 ( .A(n_256), .Y(n_336) );
AOI22xp33_ASAP7_75t_L g337 ( .A1(n_274), .A2(n_205), .B1(n_229), .B2(n_193), .Y(n_337) );
OR2x6_ASAP7_75t_L g338 ( .A(n_285), .B(n_205), .Y(n_338) );
INVx1_ASAP7_75t_L g339 ( .A(n_245), .Y(n_339) );
BUFx3_ASAP7_75t_L g340 ( .A(n_290), .Y(n_340) );
INVx3_ASAP7_75t_L g341 ( .A(n_234), .Y(n_341) );
OR2x2_ASAP7_75t_L g342 ( .A(n_279), .B(n_19), .Y(n_342) );
INVx2_ASAP7_75t_SL g343 ( .A(n_231), .Y(n_343) );
INVx2_ASAP7_75t_SL g344 ( .A(n_266), .Y(n_344) );
NAND2x1_ASAP7_75t_L g345 ( .A(n_291), .B(n_193), .Y(n_345) );
NAND2xp5_ASAP7_75t_SL g346 ( .A(n_266), .B(n_213), .Y(n_346) );
AND2x4_ASAP7_75t_L g347 ( .A(n_259), .B(n_229), .Y(n_347) );
INVx3_ASAP7_75t_SL g348 ( .A(n_250), .Y(n_348) );
BUFx3_ASAP7_75t_L g349 ( .A(n_290), .Y(n_349) );
AOI221xp5_ASAP7_75t_L g350 ( .A1(n_302), .A2(n_269), .B1(n_268), .B2(n_286), .C(n_247), .Y(n_350) );
AND2x4_ASAP7_75t_L g351 ( .A(n_313), .B(n_261), .Y(n_351) );
AOI22xp33_ASAP7_75t_L g352 ( .A1(n_304), .A2(n_339), .B1(n_316), .B2(n_281), .Y(n_352) );
OAI22xp33_ASAP7_75t_L g353 ( .A1(n_316), .A2(n_285), .B1(n_289), .B2(n_295), .Y(n_353) );
NAND2x1p5_ASAP7_75t_L g354 ( .A(n_313), .B(n_232), .Y(n_354) );
NAND2xp5_ASAP7_75t_L g355 ( .A(n_339), .B(n_246), .Y(n_355) );
NAND2xp5_ASAP7_75t_L g356 ( .A(n_298), .B(n_246), .Y(n_356) );
NAND3xp33_ASAP7_75t_L g357 ( .A(n_302), .B(n_272), .C(n_287), .Y(n_357) );
OAI22xp5_ASAP7_75t_L g358 ( .A1(n_333), .A2(n_233), .B1(n_294), .B2(n_296), .Y(n_358) );
OR2x6_ASAP7_75t_L g359 ( .A(n_338), .B(n_283), .Y(n_359) );
OAI22xp5_ASAP7_75t_L g360 ( .A1(n_333), .A2(n_283), .B1(n_240), .B2(n_275), .Y(n_360) );
INVx3_ASAP7_75t_L g361 ( .A(n_306), .Y(n_361) );
OAI22xp5_ASAP7_75t_L g362 ( .A1(n_333), .A2(n_283), .B1(n_240), .B2(n_287), .Y(n_362) );
NOR2xp33_ASAP7_75t_L g363 ( .A(n_299), .B(n_274), .Y(n_363) );
HB1xp67_ASAP7_75t_L g364 ( .A(n_333), .Y(n_364) );
INVx1_ASAP7_75t_L g365 ( .A(n_323), .Y(n_365) );
AOI22xp33_ASAP7_75t_L g366 ( .A1(n_347), .A2(n_270), .B1(n_280), .B2(n_282), .Y(n_366) );
AOI22xp33_ASAP7_75t_SL g367 ( .A1(n_342), .A2(n_241), .B1(n_282), .B2(n_284), .Y(n_367) );
AOI221xp5_ASAP7_75t_L g368 ( .A1(n_326), .A2(n_242), .B1(n_267), .B2(n_273), .C(n_244), .Y(n_368) );
AOI22xp33_ASAP7_75t_SL g369 ( .A1(n_342), .A2(n_244), .B1(n_229), .B2(n_260), .Y(n_369) );
NOR2xp33_ASAP7_75t_L g370 ( .A(n_326), .B(n_267), .Y(n_370) );
OAI22xp33_ASAP7_75t_SL g371 ( .A1(n_300), .A2(n_264), .B1(n_236), .B2(n_21), .Y(n_371) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_323), .B(n_301), .Y(n_372) );
NAND2xp5_ASAP7_75t_L g373 ( .A(n_301), .B(n_229), .Y(n_373) );
OAI22xp5_ASAP7_75t_L g374 ( .A1(n_338), .A2(n_243), .B1(n_234), .B2(n_251), .Y(n_374) );
NAND2xp33_ASAP7_75t_R g375 ( .A(n_338), .B(n_19), .Y(n_375) );
AOI21xp5_ASAP7_75t_R g376 ( .A1(n_347), .A2(n_229), .B(n_22), .Y(n_376) );
INVx1_ASAP7_75t_SL g377 ( .A(n_348), .Y(n_377) );
NAND2x1p5_ASAP7_75t_L g378 ( .A(n_313), .B(n_243), .Y(n_378) );
INVx3_ASAP7_75t_L g379 ( .A(n_306), .Y(n_379) );
INVx1_ASAP7_75t_L g380 ( .A(n_314), .Y(n_380) );
BUFx3_ASAP7_75t_L g381 ( .A(n_335), .Y(n_381) );
AOI221xp5_ASAP7_75t_L g382 ( .A1(n_353), .A2(n_314), .B1(n_329), .B2(n_324), .C(n_347), .Y(n_382) );
AOI22xp5_ASAP7_75t_L g383 ( .A1(n_353), .A2(n_338), .B1(n_347), .B2(n_309), .Y(n_383) );
OAI22xp33_ASAP7_75t_L g384 ( .A1(n_375), .A2(n_338), .B1(n_348), .B2(n_300), .Y(n_384) );
AOI22xp33_ASAP7_75t_L g385 ( .A1(n_352), .A2(n_335), .B1(n_348), .B2(n_309), .Y(n_385) );
INVx1_ASAP7_75t_L g386 ( .A(n_380), .Y(n_386) );
AOI221xp5_ASAP7_75t_L g387 ( .A1(n_370), .A2(n_322), .B1(n_319), .B2(n_315), .C(n_344), .Y(n_387) );
AOI22xp33_ASAP7_75t_L g388 ( .A1(n_352), .A2(n_309), .B1(n_311), .B2(n_315), .Y(n_388) );
INVx2_ASAP7_75t_L g389 ( .A(n_365), .Y(n_389) );
AO21x2_ASAP7_75t_L g390 ( .A1(n_357), .A2(n_308), .B(n_303), .Y(n_390) );
BUFx3_ASAP7_75t_L g391 ( .A(n_354), .Y(n_391) );
BUFx2_ASAP7_75t_L g392 ( .A(n_359), .Y(n_392) );
INVx2_ASAP7_75t_SL g393 ( .A(n_359), .Y(n_393) );
OAI22xp33_ASAP7_75t_L g394 ( .A1(n_355), .A2(n_334), .B1(n_311), .B2(n_344), .Y(n_394) );
AOI22xp33_ASAP7_75t_L g395 ( .A1(n_370), .A2(n_309), .B1(n_319), .B2(n_325), .Y(n_395) );
AND2x2_ASAP7_75t_L g396 ( .A(n_372), .B(n_334), .Y(n_396) );
OAI22xp5_ASAP7_75t_L g397 ( .A1(n_376), .A2(n_337), .B1(n_332), .B2(n_343), .Y(n_397) );
AOI22xp33_ASAP7_75t_L g398 ( .A1(n_368), .A2(n_331), .B1(n_325), .B2(n_343), .Y(n_398) );
AOI22xp33_ASAP7_75t_L g399 ( .A1(n_367), .A2(n_331), .B1(n_334), .B2(n_327), .Y(n_399) );
AND2x2_ASAP7_75t_L g400 ( .A(n_356), .B(n_305), .Y(n_400) );
AOI21xp5_ASAP7_75t_L g401 ( .A1(n_373), .A2(n_308), .B(n_318), .Y(n_401) );
AND2x2_ASAP7_75t_L g402 ( .A(n_364), .B(n_320), .Y(n_402) );
AOI22xp33_ASAP7_75t_L g403 ( .A1(n_350), .A2(n_318), .B1(n_327), .B2(n_307), .Y(n_403) );
INVx2_ASAP7_75t_L g404 ( .A(n_378), .Y(n_404) );
INVx1_ASAP7_75t_L g405 ( .A(n_364), .Y(n_405) );
OR2x2_ASAP7_75t_L g406 ( .A(n_351), .B(n_336), .Y(n_406) );
AOI221xp5_ASAP7_75t_L g407 ( .A1(n_371), .A2(n_312), .B1(n_346), .B2(n_305), .C(n_307), .Y(n_407) );
OAI22xp5_ASAP7_75t_L g408 ( .A1(n_369), .A2(n_349), .B1(n_340), .B2(n_321), .Y(n_408) );
OAI22xp33_ASAP7_75t_L g409 ( .A1(n_359), .A2(n_310), .B1(n_306), .B2(n_328), .Y(n_409) );
BUFx2_ASAP7_75t_L g410 ( .A(n_391), .Y(n_410) );
NAND3xp33_ASAP7_75t_L g411 ( .A(n_407), .B(n_366), .C(n_362), .Y(n_411) );
NOR2xp33_ASAP7_75t_L g412 ( .A(n_384), .B(n_363), .Y(n_412) );
NAND2xp5_ASAP7_75t_L g413 ( .A(n_396), .B(n_351), .Y(n_413) );
AOI221xp5_ASAP7_75t_L g414 ( .A1(n_387), .A2(n_377), .B1(n_360), .B2(n_358), .C(n_366), .Y(n_414) );
AND2x2_ASAP7_75t_L g415 ( .A(n_389), .B(n_354), .Y(n_415) );
INVx2_ASAP7_75t_L g416 ( .A(n_390), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_386), .Y(n_417) );
INVx2_ASAP7_75t_L g418 ( .A(n_390), .Y(n_418) );
NAND2xp5_ASAP7_75t_SL g419 ( .A(n_394), .B(n_361), .Y(n_419) );
INVx2_ASAP7_75t_L g420 ( .A(n_390), .Y(n_420) );
OAI22xp33_ASAP7_75t_L g421 ( .A1(n_383), .A2(n_381), .B1(n_310), .B2(n_306), .Y(n_421) );
NAND2xp5_ASAP7_75t_L g422 ( .A(n_396), .B(n_379), .Y(n_422) );
OAI221xp5_ASAP7_75t_L g423 ( .A1(n_385), .A2(n_399), .B1(n_383), .B2(n_382), .C(n_395), .Y(n_423) );
OAI221xp5_ASAP7_75t_L g424 ( .A1(n_382), .A2(n_305), .B1(n_320), .B2(n_307), .C(n_336), .Y(n_424) );
AND2x2_ASAP7_75t_L g425 ( .A(n_389), .B(n_379), .Y(n_425) );
INVx1_ASAP7_75t_L g426 ( .A(n_386), .Y(n_426) );
AND2x2_ASAP7_75t_L g427 ( .A(n_389), .B(n_361), .Y(n_427) );
AOI22xp33_ASAP7_75t_L g428 ( .A1(n_388), .A2(n_229), .B1(n_320), .B2(n_305), .Y(n_428) );
NAND4xp25_ASAP7_75t_SL g429 ( .A(n_398), .B(n_20), .C(n_23), .D(n_24), .Y(n_429) );
CKINVDCx16_ASAP7_75t_R g430 ( .A(n_391), .Y(n_430) );
NAND3xp33_ASAP7_75t_L g431 ( .A(n_407), .B(n_374), .C(n_213), .Y(n_431) );
INVx1_ASAP7_75t_L g432 ( .A(n_405), .Y(n_432) );
INVx1_ASAP7_75t_L g433 ( .A(n_405), .Y(n_433) );
OAI22xp5_ASAP7_75t_L g434 ( .A1(n_403), .A2(n_378), .B1(n_310), .B2(n_306), .Y(n_434) );
INVxp67_ASAP7_75t_R g435 ( .A(n_408), .Y(n_435) );
OAI221xp5_ASAP7_75t_L g436 ( .A1(n_387), .A2(n_307), .B1(n_320), .B2(n_345), .C(n_340), .Y(n_436) );
BUFx2_ASAP7_75t_L g437 ( .A(n_391), .Y(n_437) );
AND2x2_ASAP7_75t_L g438 ( .A(n_400), .B(n_303), .Y(n_438) );
NAND3xp33_ASAP7_75t_L g439 ( .A(n_397), .B(n_196), .C(n_216), .Y(n_439) );
AND2x2_ASAP7_75t_L g440 ( .A(n_400), .B(n_341), .Y(n_440) );
INVxp67_ASAP7_75t_SL g441 ( .A(n_406), .Y(n_441) );
NAND3xp33_ASAP7_75t_L g442 ( .A(n_397), .B(n_196), .C(n_216), .Y(n_442) );
OAI22xp5_ASAP7_75t_L g443 ( .A1(n_392), .A2(n_310), .B1(n_321), .B2(n_328), .Y(n_443) );
AO21x2_ASAP7_75t_L g444 ( .A1(n_401), .A2(n_214), .B(n_218), .Y(n_444) );
A2O1A1Ixp33_ASAP7_75t_L g445 ( .A1(n_393), .A2(n_408), .B(n_392), .C(n_401), .Y(n_445) );
NAND3xp33_ASAP7_75t_L g446 ( .A(n_412), .B(n_404), .C(n_406), .Y(n_446) );
HB1xp67_ASAP7_75t_L g447 ( .A(n_415), .Y(n_447) );
NOR2x1_ASAP7_75t_L g448 ( .A(n_410), .B(n_390), .Y(n_448) );
NAND3xp33_ASAP7_75t_L g449 ( .A(n_414), .B(n_404), .C(n_393), .Y(n_449) );
INVx1_ASAP7_75t_L g450 ( .A(n_417), .Y(n_450) );
AOI22xp33_ASAP7_75t_L g451 ( .A1(n_423), .A2(n_393), .B1(n_402), .B2(n_409), .Y(n_451) );
AND2x2_ASAP7_75t_L g452 ( .A(n_417), .B(n_404), .Y(n_452) );
NAND2xp5_ASAP7_75t_L g453 ( .A(n_432), .B(n_402), .Y(n_453) );
AND2x2_ASAP7_75t_L g454 ( .A(n_426), .B(n_20), .Y(n_454) );
INVx1_ASAP7_75t_L g455 ( .A(n_426), .Y(n_455) );
HB1xp67_ASAP7_75t_L g456 ( .A(n_415), .Y(n_456) );
INVx2_ASAP7_75t_SL g457 ( .A(n_430), .Y(n_457) );
INVx1_ASAP7_75t_L g458 ( .A(n_432), .Y(n_458) );
AOI22xp5_ASAP7_75t_L g459 ( .A1(n_411), .A2(n_310), .B1(n_328), .B2(n_321), .Y(n_459) );
INVx2_ASAP7_75t_L g460 ( .A(n_416), .Y(n_460) );
AND2x4_ASAP7_75t_L g461 ( .A(n_438), .B(n_341), .Y(n_461) );
NAND2xp5_ASAP7_75t_L g462 ( .A(n_433), .B(n_341), .Y(n_462) );
OAI33xp33_ASAP7_75t_L g463 ( .A1(n_422), .A2(n_218), .A3(n_236), .B1(n_238), .B2(n_262), .B3(n_276), .Y(n_463) );
INVx1_ASAP7_75t_L g464 ( .A(n_438), .Y(n_464) );
HB1xp67_ASAP7_75t_L g465 ( .A(n_441), .Y(n_465) );
INVx1_ASAP7_75t_L g466 ( .A(n_416), .Y(n_466) );
AND2x2_ASAP7_75t_L g467 ( .A(n_425), .B(n_341), .Y(n_467) );
AND2x2_ASAP7_75t_L g468 ( .A(n_425), .B(n_27), .Y(n_468) );
AND2x2_ASAP7_75t_L g469 ( .A(n_427), .B(n_28), .Y(n_469) );
INVx1_ASAP7_75t_L g470 ( .A(n_416), .Y(n_470) );
AND2x4_ASAP7_75t_L g471 ( .A(n_445), .B(n_30), .Y(n_471) );
INVx3_ASAP7_75t_L g472 ( .A(n_418), .Y(n_472) );
AOI22xp33_ASAP7_75t_L g473 ( .A1(n_429), .A2(n_349), .B1(n_340), .B2(n_345), .Y(n_473) );
NAND3xp33_ASAP7_75t_SL g474 ( .A(n_410), .B(n_33), .C(n_36), .Y(n_474) );
NAND2xp5_ASAP7_75t_L g475 ( .A(n_430), .B(n_330), .Y(n_475) );
INVx1_ASAP7_75t_SL g476 ( .A(n_437), .Y(n_476) );
INVx2_ASAP7_75t_L g477 ( .A(n_418), .Y(n_477) );
AOI22xp33_ASAP7_75t_L g478 ( .A1(n_411), .A2(n_349), .B1(n_330), .B2(n_317), .Y(n_478) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_413), .B(n_330), .Y(n_479) );
INVx4_ASAP7_75t_L g480 ( .A(n_437), .Y(n_480) );
INVx2_ASAP7_75t_L g481 ( .A(n_418), .Y(n_481) );
AO21x2_ASAP7_75t_L g482 ( .A1(n_439), .A2(n_238), .B(n_262), .Y(n_482) );
INVx1_ASAP7_75t_L g483 ( .A(n_420), .Y(n_483) );
INVx3_ASAP7_75t_L g484 ( .A(n_420), .Y(n_484) );
NAND3xp33_ASAP7_75t_L g485 ( .A(n_439), .B(n_181), .C(n_196), .Y(n_485) );
INVx1_ASAP7_75t_L g486 ( .A(n_420), .Y(n_486) );
INVx1_ASAP7_75t_L g487 ( .A(n_427), .Y(n_487) );
HB1xp67_ASAP7_75t_L g488 ( .A(n_440), .Y(n_488) );
INVx1_ASAP7_75t_L g489 ( .A(n_444), .Y(n_489) );
INVx2_ASAP7_75t_SL g490 ( .A(n_440), .Y(n_490) );
INVx3_ASAP7_75t_L g491 ( .A(n_444), .Y(n_491) );
AOI22xp33_ASAP7_75t_L g492 ( .A1(n_421), .A2(n_317), .B1(n_330), .B2(n_181), .Y(n_492) );
INVx1_ASAP7_75t_L g493 ( .A(n_444), .Y(n_493) );
INVx2_ASAP7_75t_L g494 ( .A(n_431), .Y(n_494) );
AO31x2_ASAP7_75t_L g495 ( .A1(n_434), .A2(n_293), .A3(n_278), .B(n_276), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_465), .B(n_428), .Y(n_496) );
INVx1_ASAP7_75t_SL g497 ( .A(n_457), .Y(n_497) );
OR2x6_ASAP7_75t_L g498 ( .A(n_480), .B(n_442), .Y(n_498) );
BUFx3_ASAP7_75t_L g499 ( .A(n_457), .Y(n_499) );
INVx2_ASAP7_75t_L g500 ( .A(n_460), .Y(n_500) );
NAND2xp5_ASAP7_75t_SL g501 ( .A(n_480), .B(n_442), .Y(n_501) );
OAI33xp33_ASAP7_75t_L g502 ( .A1(n_458), .A2(n_443), .A3(n_419), .B1(n_431), .B2(n_435), .B3(n_424), .Y(n_502) );
INVx1_ASAP7_75t_L g503 ( .A(n_458), .Y(n_503) );
INVx2_ASAP7_75t_L g504 ( .A(n_460), .Y(n_504) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_487), .B(n_443), .Y(n_505) );
HB1xp67_ASAP7_75t_L g506 ( .A(n_476), .Y(n_506) );
NAND2xp5_ASAP7_75t_L g507 ( .A(n_487), .B(n_436), .Y(n_507) );
OR2x2_ASAP7_75t_SL g508 ( .A(n_446), .B(n_435), .Y(n_508) );
INVx1_ASAP7_75t_L g509 ( .A(n_450), .Y(n_509) );
HB1xp67_ASAP7_75t_L g510 ( .A(n_476), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g511 ( .A(n_453), .B(n_200), .Y(n_511) );
AND2x2_ASAP7_75t_L g512 ( .A(n_464), .B(n_216), .Y(n_512) );
NOR4xp25_ASAP7_75t_SL g513 ( .A(n_489), .B(n_39), .C(n_44), .D(n_45), .Y(n_513) );
INVx1_ASAP7_75t_L g514 ( .A(n_450), .Y(n_514) );
AND2x2_ASAP7_75t_L g515 ( .A(n_464), .B(n_216), .Y(n_515) );
NAND2xp5_ASAP7_75t_L g516 ( .A(n_488), .B(n_200), .Y(n_516) );
HB1xp67_ASAP7_75t_L g517 ( .A(n_480), .Y(n_517) );
OR2x2_ASAP7_75t_L g518 ( .A(n_447), .B(n_216), .Y(n_518) );
INVxp67_ASAP7_75t_L g519 ( .A(n_456), .Y(n_519) );
INVx2_ASAP7_75t_L g520 ( .A(n_460), .Y(n_520) );
NOR2xp67_ASAP7_75t_SL g521 ( .A(n_485), .B(n_330), .Y(n_521) );
NOR2xp33_ASAP7_75t_L g522 ( .A(n_490), .B(n_49), .Y(n_522) );
AND2x2_ASAP7_75t_L g523 ( .A(n_455), .B(n_213), .Y(n_523) );
AND2x2_ASAP7_75t_L g524 ( .A(n_455), .B(n_213), .Y(n_524) );
NAND2xp33_ASAP7_75t_SL g525 ( .A(n_480), .B(n_317), .Y(n_525) );
AND2x2_ASAP7_75t_L g526 ( .A(n_452), .B(n_213), .Y(n_526) );
INVx1_ASAP7_75t_L g527 ( .A(n_452), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g528 ( .A(n_454), .B(n_200), .Y(n_528) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_454), .B(n_196), .Y(n_529) );
INVx1_ASAP7_75t_L g530 ( .A(n_466), .Y(n_530) );
AOI221xp5_ASAP7_75t_L g531 ( .A1(n_446), .A2(n_181), .B1(n_196), .B2(n_278), .C(n_293), .Y(n_531) );
INVx1_ASAP7_75t_L g532 ( .A(n_466), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_490), .B(n_181), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_467), .B(n_181), .Y(n_534) );
AO21x1_ASAP7_75t_L g535 ( .A1(n_471), .A2(n_50), .B(n_51), .Y(n_535) );
AND2x2_ASAP7_75t_L g536 ( .A(n_472), .B(n_54), .Y(n_536) );
AND2x2_ASAP7_75t_L g537 ( .A(n_472), .B(n_55), .Y(n_537) );
NAND2xp33_ASAP7_75t_R g538 ( .A(n_471), .B(n_56), .Y(n_538) );
OR2x6_ASAP7_75t_L g539 ( .A(n_471), .B(n_317), .Y(n_539) );
BUFx2_ASAP7_75t_L g540 ( .A(n_472), .Y(n_540) );
INVx1_ASAP7_75t_L g541 ( .A(n_470), .Y(n_541) );
AND2x2_ASAP7_75t_L g542 ( .A(n_472), .B(n_63), .Y(n_542) );
INVx1_ASAP7_75t_L g543 ( .A(n_470), .Y(n_543) );
INVx1_ASAP7_75t_L g544 ( .A(n_483), .Y(n_544) );
INVx2_ASAP7_75t_L g545 ( .A(n_477), .Y(n_545) );
OR2x2_ASAP7_75t_L g546 ( .A(n_483), .B(n_65), .Y(n_546) );
AOI22xp33_ASAP7_75t_L g547 ( .A1(n_471), .A2(n_317), .B1(n_193), .B2(n_243), .Y(n_547) );
INVx2_ASAP7_75t_SL g548 ( .A(n_475), .Y(n_548) );
AND2x2_ASAP7_75t_L g549 ( .A(n_484), .B(n_461), .Y(n_549) );
AND2x2_ASAP7_75t_L g550 ( .A(n_484), .B(n_66), .Y(n_550) );
NOR2x1_ASAP7_75t_L g551 ( .A(n_474), .B(n_67), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g552 ( .A(n_467), .B(n_72), .Y(n_552) );
AOI22xp5_ASAP7_75t_L g553 ( .A1(n_538), .A2(n_451), .B1(n_473), .B2(n_449), .Y(n_553) );
NOR2xp33_ASAP7_75t_L g554 ( .A(n_497), .B(n_449), .Y(n_554) );
INVx1_ASAP7_75t_SL g555 ( .A(n_499), .Y(n_555) );
OAI32xp33_ASAP7_75t_L g556 ( .A1(n_517), .A2(n_468), .A3(n_469), .B1(n_485), .B2(n_494), .Y(n_556) );
NAND2x1_ASAP7_75t_L g557 ( .A(n_498), .B(n_539), .Y(n_557) );
INVx2_ASAP7_75t_L g558 ( .A(n_500), .Y(n_558) );
INVx1_ASAP7_75t_L g559 ( .A(n_509), .Y(n_559) );
INVx2_ASAP7_75t_L g560 ( .A(n_500), .Y(n_560) );
INVx2_ASAP7_75t_L g561 ( .A(n_504), .Y(n_561) );
AOI21xp33_ASAP7_75t_L g562 ( .A1(n_496), .A2(n_448), .B(n_493), .Y(n_562) );
OR2x2_ASAP7_75t_L g563 ( .A(n_519), .B(n_486), .Y(n_563) );
INVx2_ASAP7_75t_L g564 ( .A(n_504), .Y(n_564) );
OAI22xp5_ASAP7_75t_L g565 ( .A1(n_508), .A2(n_492), .B1(n_459), .B2(n_469), .Y(n_565) );
OAI221xp5_ASAP7_75t_L g566 ( .A1(n_547), .A2(n_448), .B1(n_459), .B2(n_494), .C(n_462), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_527), .B(n_461), .Y(n_567) );
OAI322xp33_ASAP7_75t_L g568 ( .A1(n_507), .A2(n_514), .A3(n_503), .B1(n_505), .B2(n_548), .C1(n_543), .C2(n_544), .Y(n_568) );
OAI221xp5_ASAP7_75t_L g569 ( .A1(n_499), .A2(n_494), .B1(n_462), .B2(n_493), .C(n_489), .Y(n_569) );
AOI21xp5_ASAP7_75t_L g570 ( .A1(n_525), .A2(n_463), .B(n_482), .Y(n_570) );
NOR2xp33_ASAP7_75t_L g571 ( .A(n_502), .B(n_468), .Y(n_571) );
AOI322xp5_ASAP7_75t_L g572 ( .A1(n_514), .A2(n_486), .A3(n_491), .B1(n_461), .B2(n_481), .C1(n_477), .C2(n_484), .Y(n_572) );
NAND2xp5_ASAP7_75t_SL g573 ( .A(n_525), .B(n_491), .Y(n_573) );
OAI221xp5_ASAP7_75t_SL g574 ( .A1(n_539), .A2(n_478), .B1(n_479), .B2(n_491), .C(n_481), .Y(n_574) );
OAI22xp33_ASAP7_75t_SL g575 ( .A1(n_539), .A2(n_491), .B1(n_484), .B2(n_477), .Y(n_575) );
INVx1_ASAP7_75t_L g576 ( .A(n_530), .Y(n_576) );
INVx1_ASAP7_75t_L g577 ( .A(n_530), .Y(n_577) );
INVx2_ASAP7_75t_L g578 ( .A(n_520), .Y(n_578) );
INVx1_ASAP7_75t_L g579 ( .A(n_532), .Y(n_579) );
INVx1_ASAP7_75t_L g580 ( .A(n_532), .Y(n_580) );
INVx1_ASAP7_75t_L g581 ( .A(n_541), .Y(n_581) );
NOR2xp33_ASAP7_75t_L g582 ( .A(n_548), .B(n_461), .Y(n_582) );
AND2x2_ASAP7_75t_L g583 ( .A(n_549), .B(n_481), .Y(n_583) );
AOI22xp33_ASAP7_75t_L g584 ( .A1(n_535), .A2(n_482), .B1(n_495), .B2(n_243), .Y(n_584) );
NAND2xp5_ASAP7_75t_L g585 ( .A(n_543), .B(n_544), .Y(n_585) );
INVx1_ASAP7_75t_L g586 ( .A(n_506), .Y(n_586) );
O2A1O1Ixp33_ASAP7_75t_L g587 ( .A1(n_535), .A2(n_482), .B(n_495), .C(n_73), .Y(n_587) );
OR2x2_ASAP7_75t_L g588 ( .A(n_510), .B(n_495), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g589 ( .A(n_549), .B(n_495), .Y(n_589) );
AOI31xp33_ASAP7_75t_L g590 ( .A1(n_551), .A2(n_482), .A3(n_495), .B(n_75), .Y(n_590) );
INVx1_ASAP7_75t_SL g591 ( .A(n_536), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g592 ( .A(n_520), .B(n_495), .Y(n_592) );
INVx1_ASAP7_75t_L g593 ( .A(n_545), .Y(n_593) );
AOI22xp33_ASAP7_75t_L g594 ( .A1(n_539), .A2(n_251), .B1(n_498), .B2(n_501), .Y(n_594) );
INVx2_ASAP7_75t_L g595 ( .A(n_545), .Y(n_595) );
INVx1_ASAP7_75t_SL g596 ( .A(n_536), .Y(n_596) );
NOR2xp33_ASAP7_75t_L g597 ( .A(n_508), .B(n_251), .Y(n_597) );
NAND2x1p5_ASAP7_75t_L g598 ( .A(n_546), .B(n_251), .Y(n_598) );
INVx1_ASAP7_75t_L g599 ( .A(n_523), .Y(n_599) );
INVx1_ASAP7_75t_L g600 ( .A(n_523), .Y(n_600) );
OA33x2_ASAP7_75t_L g601 ( .A1(n_567), .A2(n_552), .A3(n_511), .B1(n_528), .B2(n_529), .B3(n_534), .Y(n_601) );
INVx2_ASAP7_75t_L g602 ( .A(n_558), .Y(n_602) );
AND2x2_ASAP7_75t_L g603 ( .A(n_583), .B(n_540), .Y(n_603) );
INVx1_ASAP7_75t_L g604 ( .A(n_559), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g605 ( .A(n_586), .B(n_540), .Y(n_605) );
AND2x2_ASAP7_75t_L g606 ( .A(n_589), .B(n_498), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g607 ( .A(n_554), .B(n_512), .Y(n_607) );
INVx1_ASAP7_75t_L g608 ( .A(n_576), .Y(n_608) );
AND2x2_ASAP7_75t_L g609 ( .A(n_599), .B(n_498), .Y(n_609) );
NOR2xp33_ASAP7_75t_L g610 ( .A(n_555), .B(n_522), .Y(n_610) );
NOR2xp33_ASAP7_75t_L g611 ( .A(n_571), .B(n_518), .Y(n_611) );
NOR2x1_ASAP7_75t_L g612 ( .A(n_557), .B(n_546), .Y(n_612) );
BUFx3_ASAP7_75t_L g613 ( .A(n_558), .Y(n_613) );
OR2x2_ASAP7_75t_L g614 ( .A(n_563), .B(n_518), .Y(n_614) );
OR2x2_ASAP7_75t_L g615 ( .A(n_588), .B(n_516), .Y(n_615) );
NAND2xp5_ASAP7_75t_L g616 ( .A(n_554), .B(n_512), .Y(n_616) );
AOI21xp33_ASAP7_75t_L g617 ( .A1(n_571), .A2(n_533), .B(n_515), .Y(n_617) );
AND2x2_ASAP7_75t_L g618 ( .A(n_600), .B(n_515), .Y(n_618) );
INVx2_ASAP7_75t_L g619 ( .A(n_560), .Y(n_619) );
NAND3xp33_ASAP7_75t_SL g620 ( .A(n_587), .B(n_513), .C(n_531), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g621 ( .A(n_577), .B(n_524), .Y(n_621) );
INVx1_ASAP7_75t_L g622 ( .A(n_579), .Y(n_622) );
XNOR2xp5_ASAP7_75t_L g623 ( .A(n_553), .B(n_537), .Y(n_623) );
NOR4xp25_ASAP7_75t_SL g624 ( .A(n_574), .B(n_521), .C(n_537), .D(n_542), .Y(n_624) );
NAND2xp33_ASAP7_75t_R g625 ( .A(n_597), .B(n_542), .Y(n_625) );
INVx1_ASAP7_75t_L g626 ( .A(n_580), .Y(n_626) );
INVx1_ASAP7_75t_SL g627 ( .A(n_591), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g628 ( .A(n_581), .B(n_524), .Y(n_628) );
NOR2x1_ASAP7_75t_L g629 ( .A(n_568), .B(n_550), .Y(n_629) );
AND2x2_ASAP7_75t_L g630 ( .A(n_561), .B(n_578), .Y(n_630) );
NAND2xp5_ASAP7_75t_SL g631 ( .A(n_575), .B(n_550), .Y(n_631) );
OAI21xp5_ASAP7_75t_L g632 ( .A1(n_590), .A2(n_594), .B(n_584), .Y(n_632) );
NOR2xp33_ASAP7_75t_L g633 ( .A(n_582), .B(n_526), .Y(n_633) );
AOI22xp5_ASAP7_75t_L g634 ( .A1(n_611), .A2(n_582), .B1(n_565), .B2(n_596), .Y(n_634) );
OAI21xp5_ASAP7_75t_L g635 ( .A1(n_629), .A2(n_594), .B(n_584), .Y(n_635) );
AOI21xp5_ASAP7_75t_L g636 ( .A1(n_629), .A2(n_573), .B(n_556), .Y(n_636) );
OAI21xp33_ASAP7_75t_L g637 ( .A1(n_606), .A2(n_572), .B(n_569), .Y(n_637) );
NAND3xp33_ASAP7_75t_L g638 ( .A(n_632), .B(n_562), .C(n_566), .Y(n_638) );
XNOR2xp5_ASAP7_75t_L g639 ( .A(n_623), .B(n_585), .Y(n_639) );
OAI22xp5_ASAP7_75t_L g640 ( .A1(n_623), .A2(n_598), .B1(n_573), .B2(n_597), .Y(n_640) );
AOI32xp33_ASAP7_75t_L g641 ( .A1(n_612), .A2(n_592), .A3(n_593), .B1(n_564), .B2(n_595), .Y(n_641) );
AND4x1_ASAP7_75t_L g642 ( .A(n_610), .B(n_521), .C(n_570), .D(n_526), .Y(n_642) );
NAND3xp33_ASAP7_75t_L g643 ( .A(n_624), .B(n_617), .C(n_605), .Y(n_643) );
OR2x2_ASAP7_75t_L g644 ( .A(n_614), .B(n_615), .Y(n_644) );
AOI221x1_ASAP7_75t_L g645 ( .A1(n_620), .A2(n_616), .B1(n_607), .B2(n_622), .C(n_604), .Y(n_645) );
OAI221xp5_ASAP7_75t_L g646 ( .A1(n_601), .A2(n_631), .B1(n_625), .B2(n_627), .C(n_614), .Y(n_646) );
INVx1_ASAP7_75t_L g647 ( .A(n_608), .Y(n_647) );
NAND4xp75_ASAP7_75t_L g648 ( .A(n_609), .B(n_618), .C(n_633), .D(n_624), .Y(n_648) );
NAND2xp5_ASAP7_75t_L g649 ( .A(n_608), .B(n_626), .Y(n_649) );
INVx1_ASAP7_75t_L g650 ( .A(n_644), .Y(n_650) );
NAND2xp5_ASAP7_75t_L g651 ( .A(n_634), .B(n_637), .Y(n_651) );
CKINVDCx5p33_ASAP7_75t_R g652 ( .A(n_639), .Y(n_652) );
AOI22xp5_ASAP7_75t_L g653 ( .A1(n_638), .A2(n_609), .B1(n_618), .B2(n_603), .Y(n_653) );
OAI21xp5_ASAP7_75t_SL g654 ( .A1(n_645), .A2(n_621), .B(n_628), .Y(n_654) );
AND2x4_ASAP7_75t_L g655 ( .A(n_635), .B(n_613), .Y(n_655) );
NAND2xp33_ASAP7_75t_R g656 ( .A(n_635), .B(n_630), .Y(n_656) );
HB1xp67_ASAP7_75t_L g657 ( .A(n_649), .Y(n_657) );
INVx1_ASAP7_75t_L g658 ( .A(n_649), .Y(n_658) );
OAI221xp5_ASAP7_75t_L g659 ( .A1(n_646), .A2(n_643), .B1(n_641), .B2(n_640), .C(n_642), .Y(n_659) );
AOI22xp33_ASAP7_75t_L g660 ( .A1(n_640), .A2(n_613), .B1(n_602), .B2(n_619), .Y(n_660) );
NOR2x1_ASAP7_75t_L g661 ( .A(n_648), .B(n_619), .Y(n_661) );
O2A1O1Ixp33_ASAP7_75t_L g662 ( .A1(n_647), .A2(n_636), .B(n_638), .C(n_646), .Y(n_662) );
NAND4xp25_ASAP7_75t_L g663 ( .A(n_645), .B(n_638), .C(n_635), .D(n_643), .Y(n_663) );
INVx1_ASAP7_75t_SL g664 ( .A(n_644), .Y(n_664) );
INVx1_ASAP7_75t_L g665 ( .A(n_657), .Y(n_665) );
OR2x2_ASAP7_75t_L g666 ( .A(n_657), .B(n_658), .Y(n_666) );
HB1xp67_ASAP7_75t_L g667 ( .A(n_664), .Y(n_667) );
CKINVDCx5p33_ASAP7_75t_R g668 ( .A(n_652), .Y(n_668) );
NOR3xp33_ASAP7_75t_SL g669 ( .A(n_668), .B(n_663), .C(n_659), .Y(n_669) );
AND2x4_ASAP7_75t_L g670 ( .A(n_667), .B(n_650), .Y(n_670) );
AOI22xp5_ASAP7_75t_L g671 ( .A1(n_665), .A2(n_651), .B1(n_656), .B2(n_655), .Y(n_671) );
NOR2xp33_ASAP7_75t_R g672 ( .A(n_670), .B(n_665), .Y(n_672) );
NOR2xp33_ASAP7_75t_L g673 ( .A(n_671), .B(n_662), .Y(n_673) );
INVx2_ASAP7_75t_L g674 ( .A(n_673), .Y(n_674) );
AOI322xp5_ASAP7_75t_L g675 ( .A1(n_674), .A2(n_669), .A3(n_661), .B1(n_660), .B2(n_655), .C1(n_672), .C2(n_653), .Y(n_675) );
AO21x1_ASAP7_75t_L g676 ( .A1(n_675), .A2(n_666), .B(n_654), .Y(n_676) );
endmodule