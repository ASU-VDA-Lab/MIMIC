module real_jpeg_9961_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_316, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_316;
input n_10;
input n_9;

output n_17;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_216;
wire n_202;
wire n_127;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_215;
wire n_166;
wire n_176;
wire n_312;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_299;
wire n_243;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

A2O1A1O1Ixp25_ASAP7_75t_L g142 ( 
.A1(n_1),
.A2(n_48),
.B(n_58),
.C(n_143),
.D(n_144),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_1),
.B(n_48),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_1),
.B(n_46),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_1),
.Y(n_177)
);

OAI21xp33_ASAP7_75t_L g182 ( 
.A1(n_1),
.A2(n_82),
.B(n_162),
.Y(n_182)
);

A2O1A1O1Ixp25_ASAP7_75t_L g195 ( 
.A1(n_1),
.A2(n_31),
.B(n_42),
.C(n_196),
.D(n_197),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_1),
.B(n_31),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_1),
.B(n_130),
.Y(n_219)
);

AOI21xp33_ASAP7_75t_L g235 ( 
.A1(n_1),
.A2(n_28),
.B(n_32),
.Y(n_235)
);

OAI22xp33_ASAP7_75t_SL g252 ( 
.A1(n_1),
.A2(n_26),
.B1(n_34),
.B2(n_177),
.Y(n_252)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_2),
.A2(n_31),
.B1(n_32),
.B2(n_54),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_2),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_2),
.A2(n_47),
.B1(n_48),
.B2(n_54),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_2),
.A2(n_54),
.B1(n_63),
.B2(n_65),
.Y(n_120)
);

BUFx12_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

OAI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_4),
.A2(n_26),
.B1(n_34),
.B2(n_91),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_4),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_L g145 ( 
.A1(n_4),
.A2(n_47),
.B1(n_48),
.B2(n_91),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_4),
.A2(n_63),
.B1(n_65),
.B2(n_91),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_L g198 ( 
.A1(n_4),
.A2(n_31),
.B1(n_32),
.B2(n_91),
.Y(n_198)
);

INVx2_ASAP7_75t_SL g83 ( 
.A(n_5),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_5),
.B(n_163),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_5),
.A2(n_168),
.B1(n_170),
.B2(n_171),
.Y(n_167)
);

AOI21xp5_ASAP7_75t_L g205 ( 
.A1(n_5),
.A2(n_180),
.B(n_206),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_5),
.A2(n_170),
.B1(n_206),
.B2(n_221),
.Y(n_220)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_6),
.Y(n_64)
);

BUFx10_ASAP7_75t_L g60 ( 
.A(n_7),
.Y(n_60)
);

BUFx6f_ASAP7_75t_SL g44 ( 
.A(n_8),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_9),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g156 ( 
.A1(n_10),
.A2(n_47),
.B1(n_48),
.B2(n_157),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_10),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_SL g169 ( 
.A1(n_10),
.A2(n_63),
.B1(n_65),
.B2(n_157),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_SL g215 ( 
.A1(n_10),
.A2(n_31),
.B1(n_32),
.B2(n_157),
.Y(n_215)
);

AOI22xp33_ASAP7_75t_SL g261 ( 
.A1(n_10),
.A2(n_26),
.B1(n_34),
.B2(n_157),
.Y(n_261)
);

AOI22xp33_ASAP7_75t_SL g36 ( 
.A1(n_11),
.A2(n_26),
.B1(n_34),
.B2(n_37),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_11),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_11),
.A2(n_31),
.B1(n_32),
.B2(n_37),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_11),
.A2(n_37),
.B1(n_47),
.B2(n_48),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_11),
.A2(n_37),
.B1(n_63),
.B2(n_65),
.Y(n_221)
);

BUFx10_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_13),
.A2(n_31),
.B1(n_32),
.B2(n_51),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_13),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_L g86 ( 
.A1(n_13),
.A2(n_47),
.B1(n_48),
.B2(n_51),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_13),
.A2(n_26),
.B1(n_34),
.B2(n_51),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g239 ( 
.A1(n_13),
.A2(n_51),
.B1(n_63),
.B2(n_65),
.Y(n_239)
);

AOI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_14),
.A2(n_26),
.B1(n_34),
.B2(n_128),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_14),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_SL g161 ( 
.A1(n_14),
.A2(n_63),
.B1(n_65),
.B2(n_128),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_L g194 ( 
.A1(n_14),
.A2(n_47),
.B1(n_48),
.B2(n_128),
.Y(n_194)
);

AOI22xp33_ASAP7_75t_SL g249 ( 
.A1(n_14),
.A2(n_31),
.B1(n_32),
.B2(n_128),
.Y(n_249)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_15),
.A2(n_47),
.B1(n_48),
.B2(n_68),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_15),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_15),
.A2(n_63),
.B1(n_65),
.B2(n_68),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_15),
.A2(n_31),
.B1(n_32),
.B2(n_68),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g33 ( 
.A1(n_16),
.A2(n_26),
.B1(n_34),
.B2(n_35),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_16),
.Y(n_35)
);

OAI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_16),
.A2(n_31),
.B1(n_32),
.B2(n_35),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_16),
.A2(n_35),
.B1(n_63),
.B2(n_65),
.Y(n_206)
);

AOI22xp33_ASAP7_75t_L g246 ( 
.A1(n_16),
.A2(n_35),
.B1(n_47),
.B2(n_48),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_107),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_106),
.Y(n_18)
);

INVxp67_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_93),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_21),
.B(n_93),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_70),
.C(n_78),
.Y(n_21)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_22),
.A2(n_70),
.B1(n_71),
.B2(n_133),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_22),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_24),
.B1(n_38),
.B2(n_39),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_23),
.A2(n_24),
.B1(n_95),
.B2(n_96),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_24),
.Y(n_23)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_24),
.B(n_55),
.C(n_69),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g24 ( 
.A1(n_25),
.A2(n_30),
.B1(n_33),
.B2(n_36),
.Y(n_24)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_25),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_25),
.A2(n_30),
.B1(n_36),
.B2(n_98),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_SL g126 ( 
.A1(n_25),
.A2(n_127),
.B(n_129),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_25),
.A2(n_30),
.B1(n_127),
.B2(n_261),
.Y(n_281)
);

A2O1A1Ixp33_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_27),
.B(n_29),
.C(n_30),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_26),
.B(n_27),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_26),
.Y(n_34)
);

A2O1A1Ixp33_ASAP7_75t_L g234 ( 
.A1(n_26),
.A2(n_27),
.B(n_177),
.C(n_235),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g30 ( 
.A1(n_27),
.A2(n_28),
.B1(n_31),
.B2(n_32),
.Y(n_30)
);

CKINVDCx14_ASAP7_75t_R g27 ( 
.A(n_28),
.Y(n_27)
);

OAI21xp5_ASAP7_75t_L g88 ( 
.A1(n_30),
.A2(n_33),
.B(n_89),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_30),
.Y(n_130)
);

OAI21xp33_ASAP7_75t_L g260 ( 
.A1(n_30),
.A2(n_89),
.B(n_261),
.Y(n_260)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

O2A1O1Ixp33_ASAP7_75t_SL g42 ( 
.A1(n_32),
.A2(n_43),
.B(n_45),
.C(n_46),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_32),
.B(n_43),
.Y(n_45)
);

CKINVDCx16_ASAP7_75t_R g38 ( 
.A(n_39),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g39 ( 
.A1(n_40),
.A2(n_55),
.B1(n_56),
.B2(n_69),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_40),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g40 ( 
.A1(n_41),
.A2(n_49),
.B1(n_52),
.B2(n_53),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_41),
.A2(n_52),
.B1(n_53),
.B2(n_102),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_41),
.A2(n_52),
.B1(n_215),
.B2(n_249),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_L g263 ( 
.A1(n_41),
.A2(n_249),
.B(n_264),
.Y(n_263)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_42),
.A2(n_46),
.B1(n_50),
.B2(n_73),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_42),
.A2(n_46),
.B1(n_73),
.B2(n_124),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_42),
.B(n_217),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g46 ( 
.A1(n_43),
.A2(n_44),
.B1(n_47),
.B2(n_48),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_44),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_44),
.B(n_47),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_45),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_46),
.Y(n_52)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_47),
.Y(n_48)
);

O2A1O1Ixp33_ASAP7_75t_L g58 ( 
.A1(n_47),
.A2(n_59),
.B(n_61),
.C(n_62),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_47),
.B(n_59),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_48),
.A2(n_196),
.B1(n_203),
.B2(n_204),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_50),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_52),
.B(n_198),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_L g214 ( 
.A1(n_52),
.A2(n_215),
.B(n_216),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_L g278 ( 
.A1(n_52),
.A2(n_216),
.B(n_279),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_55),
.A2(n_56),
.B1(n_101),
.B2(n_103),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_56),
.Y(n_55)
);

AOI21xp5_ASAP7_75t_SL g56 ( 
.A1(n_57),
.A2(n_66),
.B(n_67),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_57),
.A2(n_66),
.B1(n_76),
.B2(n_86),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_57),
.A2(n_66),
.B1(n_86),
.B2(n_122),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_57),
.A2(n_66),
.B1(n_156),
.B2(n_194),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_SL g225 ( 
.A1(n_57),
.A2(n_194),
.B(n_226),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_L g269 ( 
.A1(n_57),
.A2(n_66),
.B1(n_122),
.B2(n_246),
.Y(n_269)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_58),
.A2(n_62),
.B1(n_75),
.B2(n_77),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_58),
.B(n_159),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_59),
.A2(n_60),
.B1(n_63),
.B2(n_65),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_59),
.B(n_65),
.Y(n_148)
);

CKINVDCx16_ASAP7_75t_R g59 ( 
.A(n_60),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_61),
.A2(n_63),
.B1(n_148),
.B2(n_149),
.Y(n_147)
);

CKINVDCx16_ASAP7_75t_R g66 ( 
.A(n_62),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_63),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_63),
.B(n_83),
.Y(n_82)
);

BUFx24_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g183 ( 
.A(n_65),
.B(n_184),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_66),
.B(n_145),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_L g155 ( 
.A1(n_66),
.A2(n_156),
.B(n_158),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g176 ( 
.A(n_66),
.B(n_177),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_L g245 ( 
.A1(n_66),
.A2(n_158),
.B(n_246),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_67),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_71),
.Y(n_70)
);

OAI21xp5_ASAP7_75t_L g115 ( 
.A1(n_71),
.A2(n_72),
.B(n_74),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_74),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_76),
.Y(n_75)
);

XNOR2xp5_ASAP7_75t_L g131 ( 
.A(n_78),
.B(n_132),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_L g78 ( 
.A1(n_79),
.A2(n_87),
.B(n_88),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_79),
.A2(n_80),
.B1(n_111),
.B2(n_113),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_80),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_85),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_81),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_81),
.A2(n_87),
.B1(n_88),
.B2(n_112),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g295 ( 
.A1(n_81),
.A2(n_85),
.B1(n_87),
.B2(n_296),
.Y(n_295)
);

AOI21xp5_ASAP7_75t_L g81 ( 
.A1(n_82),
.A2(n_83),
.B(n_84),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_82),
.A2(n_83),
.B1(n_84),
.B2(n_120),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_SL g160 ( 
.A1(n_82),
.A2(n_161),
.B(n_162),
.Y(n_160)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_82),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_82),
.B(n_164),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_82),
.A2(n_83),
.B1(n_238),
.B2(n_239),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_L g268 ( 
.A1(n_82),
.A2(n_83),
.B1(n_120),
.B2(n_239),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_L g178 ( 
.A1(n_83),
.A2(n_169),
.B(n_179),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_83),
.B(n_177),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_85),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_88),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_92),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_90),
.B(n_130),
.Y(n_129)
);

AOI21xp5_ASAP7_75t_L g251 ( 
.A1(n_92),
.A2(n_252),
.B(n_253),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_105),
.Y(n_93)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_97),
.A2(n_99),
.B1(n_100),
.B2(n_104),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_97),
.Y(n_104)
);

CKINVDCx16_ASAP7_75t_R g99 ( 
.A(n_100),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_101),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_L g107 ( 
.A1(n_108),
.A2(n_134),
.B(n_314),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_131),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g314 ( 
.A(n_109),
.B(n_131),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_110),
.B(n_114),
.C(n_116),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g300 ( 
.A1(n_110),
.A2(n_114),
.B1(n_115),
.B2(n_301),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_110),
.Y(n_301)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_111),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_115),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_116),
.A2(n_117),
.B1(n_299),
.B2(n_300),
.Y(n_298)
);

CKINVDCx16_ASAP7_75t_R g116 ( 
.A(n_117),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_118),
.B(n_123),
.C(n_125),
.Y(n_117)
);

XOR2xp5_ASAP7_75t_L g292 ( 
.A(n_118),
.B(n_293),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_121),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_119),
.B(n_121),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_L g293 ( 
.A1(n_123),
.A2(n_125),
.B1(n_126),
.B2(n_294),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_123),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_124),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_126),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_129),
.Y(n_253)
);

AOI321xp33_ASAP7_75t_L g134 ( 
.A1(n_135),
.A2(n_289),
.A3(n_302),
.B1(n_308),
.B2(n_313),
.C(n_316),
.Y(n_134)
);

NOR3xp33_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_255),
.C(n_285),
.Y(n_135)
);

AOI21xp5_ASAP7_75t_L g136 ( 
.A1(n_137),
.A2(n_228),
.B(n_254),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_SL g137 ( 
.A1(n_138),
.A2(n_209),
.B(n_227),
.Y(n_137)
);

AOI21xp5_ASAP7_75t_L g138 ( 
.A1(n_139),
.A2(n_188),
.B(n_208),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_SL g139 ( 
.A1(n_140),
.A2(n_165),
.B(n_187),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_150),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_141),
.B(n_150),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_SL g141 ( 
.A(n_142),
.B(n_146),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_142),
.A2(n_146),
.B1(n_147),
.B2(n_173),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_142),
.Y(n_173)
);

INVxp67_ASAP7_75t_L g149 ( 
.A(n_143),
.Y(n_149)
);

INVxp67_ASAP7_75t_L g226 ( 
.A(n_144),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_145),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_147),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_160),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_152),
.A2(n_153),
.B1(n_154),
.B2(n_155),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_152),
.B(n_155),
.C(n_160),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_153),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_155),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_161),
.Y(n_171)
);

INVxp67_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

AOI21xp5_ASAP7_75t_L g165 ( 
.A1(n_166),
.A2(n_174),
.B(n_186),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_172),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_SL g186 ( 
.A(n_167),
.B(n_172),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_169),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_SL g174 ( 
.A1(n_175),
.A2(n_181),
.B(n_185),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_178),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_176),
.B(n_178),
.Y(n_185)
);

CKINVDCx16_ASAP7_75t_R g179 ( 
.A(n_180),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_182),
.B(n_183),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_190),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_SL g208 ( 
.A(n_189),
.B(n_190),
.Y(n_208)
);

AOI22xp33_ASAP7_75t_SL g190 ( 
.A1(n_191),
.A2(n_192),
.B1(n_201),
.B2(n_207),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_193),
.A2(n_195),
.B1(n_199),
.B2(n_200),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_193),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_195),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_195),
.B(n_200),
.C(n_207),
.Y(n_210)
);

INVxp67_ASAP7_75t_L g264 ( 
.A(n_197),
.Y(n_264)
);

CKINVDCx16_ASAP7_75t_R g217 ( 
.A(n_198),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_201),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_205),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_202),
.B(n_205),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_211),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_210),
.B(n_211),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_223),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_212),
.B(n_224),
.C(n_225),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_213),
.A2(n_214),
.B1(n_218),
.B2(n_222),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_213),
.B(n_219),
.C(n_220),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_214),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_218),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_220),
.Y(n_218)
);

CKINVDCx16_ASAP7_75t_R g238 ( 
.A(n_221),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_225),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_230),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_SL g254 ( 
.A(n_229),
.B(n_230),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_243),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_232),
.A2(n_240),
.B1(n_241),
.B2(n_242),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_232),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_232),
.B(n_242),
.C(n_243),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_233),
.A2(n_234),
.B1(n_236),
.B2(n_237),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_233),
.B(n_237),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_234),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_237),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_240),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_251),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_245),
.A2(n_247),
.B1(n_248),
.B2(n_250),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_245),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_247),
.B(n_250),
.C(n_251),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_248),
.Y(n_247)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

AOI21xp33_ASAP7_75t_L g309 ( 
.A1(n_256),
.A2(n_310),
.B(n_311),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_257),
.B(n_271),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_257),
.B(n_271),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_267),
.C(n_270),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_258),
.B(n_288),
.Y(n_287)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_259),
.B(n_266),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_260),
.A2(n_262),
.B1(n_263),
.B2(n_265),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_260),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_262),
.B(n_265),
.C(n_266),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_263),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_267),
.B(n_270),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_268),
.B(n_269),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_268),
.B(n_269),
.Y(n_276)
);

AOI22xp33_ASAP7_75t_SL g271 ( 
.A1(n_272),
.A2(n_273),
.B1(n_283),
.B2(n_284),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_274),
.B(n_275),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_274),
.B(n_275),
.C(n_284),
.Y(n_304)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_276),
.B(n_277),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_276),
.B(n_280),
.C(n_282),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_278),
.A2(n_280),
.B1(n_281),
.B2(n_282),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_278),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_281),
.Y(n_280)
);

CKINVDCx16_ASAP7_75t_R g284 ( 
.A(n_283),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_286),
.B(n_287),
.Y(n_285)
);

AND2x2_ASAP7_75t_L g310 ( 
.A(n_286),
.B(n_287),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_290),
.B(n_298),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_SL g313 ( 
.A(n_290),
.B(n_298),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_291),
.B(n_295),
.C(n_297),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_291),
.A2(n_292),
.B1(n_295),
.B2(n_307),
.Y(n_306)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_295),
.Y(n_307)
);

XOR2xp5_ASAP7_75t_L g305 ( 
.A(n_297),
.B(n_306),
.Y(n_305)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

OAI21xp5_ASAP7_75t_SL g308 ( 
.A1(n_303),
.A2(n_309),
.B(n_312),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_304),
.B(n_305),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_SL g312 ( 
.A(n_304),
.B(n_305),
.Y(n_312)
);


endmodule