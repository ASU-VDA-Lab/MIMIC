module fake_jpeg_26028_n_311 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_311);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_311;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

BUFx3_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_4),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

INVx6_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

BUFx12_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_10),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_0),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_34),
.Y(n_53)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_31),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_35),
.B(n_41),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

INVx5_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_37),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_38),
.Y(n_47)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_16),
.Y(n_40)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_40),
.Y(n_63)
);

CKINVDCx16_ASAP7_75t_R g41 ( 
.A(n_27),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_42),
.Y(n_46)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_27),
.Y(n_43)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_43),
.Y(n_65)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_43),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_44),
.B(n_61),
.Y(n_78)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_42),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_48),
.Y(n_77)
);

OAI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_35),
.A2(n_25),
.B1(n_28),
.B2(n_29),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_51),
.A2(n_56),
.B1(n_59),
.B2(n_23),
.Y(n_72)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_42),
.Y(n_52)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_52),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_39),
.A2(n_25),
.B1(n_32),
.B2(n_21),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_54),
.A2(n_18),
.B1(n_33),
.B2(n_26),
.Y(n_70)
);

INVxp67_ASAP7_75t_SL g55 ( 
.A(n_41),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_55),
.B(n_62),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_37),
.A2(n_25),
.B1(n_32),
.B2(n_21),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_43),
.A2(n_28),
.B1(n_30),
.B2(n_20),
.Y(n_58)
);

INVxp67_ASAP7_75t_L g83 ( 
.A(n_58),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_37),
.A2(n_30),
.B1(n_29),
.B2(n_20),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_34),
.Y(n_60)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_60),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_34),
.B(n_31),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_34),
.B(n_31),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_38),
.A2(n_33),
.B1(n_18),
.B2(n_17),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_64),
.A2(n_33),
.B1(n_18),
.B2(n_23),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_34),
.B(n_22),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_66),
.B(n_38),
.Y(n_84)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_46),
.Y(n_68)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_68),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_49),
.B(n_17),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_69),
.B(n_76),
.Y(n_95)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_70),
.Y(n_101)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_72),
.Y(n_108)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_59),
.Y(n_73)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_73),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_74),
.Y(n_105)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_54),
.Y(n_75)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_75),
.Y(n_113)
);

INVx5_ASAP7_75t_L g76 ( 
.A(n_53),
.Y(n_76)
);

INVx8_ASAP7_75t_L g79 ( 
.A(n_46),
.Y(n_79)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_79),
.Y(n_114)
);

BUFx2_ASAP7_75t_L g80 ( 
.A(n_50),
.Y(n_80)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_80),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_58),
.A2(n_61),
.B1(n_57),
.B2(n_66),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_82),
.A2(n_88),
.B1(n_52),
.B2(n_65),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_84),
.B(n_89),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_49),
.B(n_19),
.Y(n_85)
);

FAx1_ASAP7_75t_SL g116 ( 
.A(n_85),
.B(n_27),
.CI(n_22),
.CON(n_116),
.SN(n_116)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_60),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_86),
.Y(n_93)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_57),
.Y(n_87)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_87),
.Y(n_91)
);

AO22x1_ASAP7_75t_SL g88 ( 
.A1(n_50),
.A2(n_40),
.B1(n_36),
.B2(n_23),
.Y(n_88)
);

INVx4_ASAP7_75t_SL g89 ( 
.A(n_53),
.Y(n_89)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_63),
.Y(n_90)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_90),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_78),
.B(n_40),
.C(n_36),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_96),
.B(n_88),
.C(n_70),
.Y(n_120)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_68),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_98),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_75),
.A2(n_50),
.B1(n_48),
.B2(n_63),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_99),
.A2(n_106),
.B1(n_89),
.B2(n_80),
.Y(n_134)
);

O2A1O1Ixp33_ASAP7_75t_SL g100 ( 
.A1(n_83),
.A2(n_56),
.B(n_44),
.C(n_53),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_L g122 ( 
.A1(n_100),
.A2(n_83),
.B(n_71),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_67),
.B(n_47),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_102),
.B(n_103),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_85),
.B(n_47),
.Y(n_103)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_87),
.Y(n_104)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_104),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_84),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_107),
.B(n_109),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_78),
.B(n_17),
.Y(n_109)
);

HB1xp67_ASAP7_75t_L g110 ( 
.A(n_81),
.Y(n_110)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_110),
.Y(n_128)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_79),
.Y(n_112)
);

INVxp33_ASAP7_75t_L g129 ( 
.A(n_112),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_116),
.B(n_22),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_111),
.B(n_82),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_SL g150 ( 
.A(n_117),
.B(n_130),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_96),
.B(n_73),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_118),
.B(n_123),
.Y(n_163)
);

OR2x2_ASAP7_75t_L g119 ( 
.A(n_97),
.B(n_72),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_SL g166 ( 
.A1(n_119),
.A2(n_136),
.B(n_24),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g145 ( 
.A(n_120),
.B(n_116),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_L g147 ( 
.A1(n_122),
.A2(n_126),
.B(n_101),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_107),
.B(n_88),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_105),
.A2(n_90),
.B1(n_71),
.B2(n_86),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_124),
.A2(n_133),
.B1(n_115),
.B2(n_114),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_111),
.B(n_77),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_127),
.B(n_132),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_93),
.B(n_77),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_113),
.B(n_77),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_105),
.A2(n_81),
.B1(n_65),
.B2(n_80),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_134),
.A2(n_141),
.B1(n_104),
.B2(n_92),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_98),
.A2(n_76),
.B1(n_89),
.B2(n_45),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_SL g157 ( 
.A1(n_135),
.A2(n_112),
.B1(n_94),
.B2(n_115),
.Y(n_157)
);

AOI21xp5_ASAP7_75t_L g136 ( 
.A1(n_113),
.A2(n_0),
.B(n_1),
.Y(n_136)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_99),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_138),
.B(n_140),
.Y(n_160)
);

OAI22x1_ASAP7_75t_SL g139 ( 
.A1(n_100),
.A2(n_45),
.B1(n_60),
.B2(n_26),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_L g169 ( 
.A1(n_139),
.A2(n_143),
.B1(n_138),
.B2(n_129),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g140 ( 
.A(n_95),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_108),
.A2(n_45),
.B1(n_26),
.B2(n_24),
.Y(n_141)
);

CKINVDCx16_ASAP7_75t_R g142 ( 
.A(n_106),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_142),
.B(n_92),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_L g143 ( 
.A1(n_100),
.A2(n_53),
.B(n_27),
.Y(n_143)
);

AOI21xp5_ASAP7_75t_L g168 ( 
.A1(n_143),
.A2(n_122),
.B(n_139),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_130),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_144),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_145),
.B(n_149),
.C(n_119),
.Y(n_182)
);

OAI32xp33_ASAP7_75t_L g146 ( 
.A1(n_126),
.A2(n_108),
.A3(n_101),
.B1(n_116),
.B2(n_93),
.Y(n_146)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_146),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_L g190 ( 
.A1(n_147),
.A2(n_131),
.B(n_137),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_132),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_148),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_118),
.B(n_94),
.C(n_114),
.Y(n_149)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_127),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_151),
.B(n_152),
.Y(n_174)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_124),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_121),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_153),
.B(n_155),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_154),
.A2(n_157),
.B1(n_169),
.B2(n_139),
.Y(n_173)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_121),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_123),
.Y(n_156)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_156),
.Y(n_192)
);

INVxp67_ASAP7_75t_L g158 ( 
.A(n_135),
.Y(n_158)
);

CKINVDCx14_ASAP7_75t_R g181 ( 
.A(n_158),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g159 ( 
.A(n_125),
.B(n_91),
.Y(n_159)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_159),
.B(n_162),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_137),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_161),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g162 ( 
.A(n_125),
.B(n_91),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_164),
.A2(n_134),
.B1(n_128),
.B2(n_120),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_SL g194 ( 
.A1(n_165),
.A2(n_166),
.B(n_168),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_117),
.B(n_24),
.Y(n_170)
);

CKINVDCx14_ASAP7_75t_R g197 ( 
.A(n_170),
.Y(n_197)
);

INVxp67_ASAP7_75t_L g171 ( 
.A(n_143),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_171),
.A2(n_136),
.B1(n_142),
.B2(n_119),
.Y(n_177)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_133),
.Y(n_172)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_172),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_173),
.A2(n_160),
.B1(n_153),
.B2(n_155),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g175 ( 
.A(n_145),
.B(n_120),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_175),
.B(n_189),
.Y(n_217)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_167),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_176),
.B(n_198),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_177),
.A2(n_178),
.B1(n_169),
.B2(n_170),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_156),
.A2(n_165),
.B1(n_164),
.B2(n_152),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_180),
.A2(n_183),
.B1(n_2),
.B2(n_3),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_182),
.B(n_190),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_172),
.A2(n_141),
.B1(n_128),
.B2(n_131),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g189 ( 
.A(n_149),
.B(n_137),
.Y(n_189)
);

AOI21xp5_ASAP7_75t_L g191 ( 
.A1(n_166),
.A2(n_0),
.B(n_1),
.Y(n_191)
);

AOI21xp5_ASAP7_75t_L g216 ( 
.A1(n_191),
.A2(n_194),
.B(n_190),
.Y(n_216)
);

A2O1A1O1Ixp25_ASAP7_75t_L g193 ( 
.A1(n_147),
.A2(n_146),
.B(n_150),
.C(n_163),
.D(n_168),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_SL g214 ( 
.A(n_193),
.B(n_196),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_159),
.B(n_162),
.Y(n_196)
);

INVxp67_ASAP7_75t_L g198 ( 
.A(n_160),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_175),
.B(n_163),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_201),
.B(n_219),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_202),
.A2(n_207),
.B1(n_208),
.B2(n_210),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_185),
.B(n_196),
.C(n_189),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_203),
.B(n_213),
.C(n_191),
.Y(n_227)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_188),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_204),
.B(n_206),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_181),
.A2(n_144),
.B1(n_148),
.B2(n_151),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_205),
.B(n_177),
.Y(n_224)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_188),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_187),
.A2(n_150),
.B1(n_154),
.B2(n_167),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_174),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_209),
.B(n_211),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_187),
.A2(n_161),
.B1(n_19),
.B2(n_9),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_179),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_186),
.B(n_19),
.Y(n_212)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_212),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_185),
.B(n_8),
.C(n_14),
.Y(n_213)
);

INVx4_ASAP7_75t_L g215 ( 
.A(n_178),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_215),
.B(n_216),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_197),
.Y(n_218)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_218),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_182),
.B(n_8),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_195),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_220),
.A2(n_222),
.B1(n_198),
.B2(n_195),
.Y(n_236)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_174),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_221),
.B(n_223),
.Y(n_237)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_180),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_224),
.B(n_227),
.Y(n_258)
);

INVx3_ASAP7_75t_L g226 ( 
.A(n_218),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_226),
.B(n_236),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_199),
.B(n_194),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_228),
.B(n_232),
.Y(n_249)
);

CKINVDCx16_ASAP7_75t_R g231 ( 
.A(n_200),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_231),
.B(n_239),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_199),
.B(n_193),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_202),
.B(n_184),
.Y(n_234)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_234),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_205),
.B(n_183),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_217),
.B(n_192),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_240),
.B(n_241),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_217),
.B(n_192),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_222),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_242),
.B(n_216),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_220),
.B(n_10),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_SL g250 ( 
.A(n_243),
.B(n_215),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_240),
.B(n_203),
.C(n_201),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_246),
.B(n_260),
.C(n_227),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_225),
.B(n_213),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_SL g266 ( 
.A(n_247),
.B(n_257),
.Y(n_266)
);

FAx1_ASAP7_75t_SL g248 ( 
.A(n_230),
.B(n_214),
.CI(n_219),
.CON(n_248),
.SN(n_248)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_248),
.Y(n_263)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_250),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_253),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_SL g255 ( 
.A(n_244),
.B(n_214),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_255),
.Y(n_261)
);

INVxp67_ASAP7_75t_L g256 ( 
.A(n_229),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_256),
.B(n_12),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_226),
.B(n_9),
.Y(n_257)
);

AOI21xp5_ASAP7_75t_SL g259 ( 
.A1(n_237),
.A2(n_11),
.B(n_14),
.Y(n_259)
);

OAI21xp5_ASAP7_75t_SL g267 ( 
.A1(n_259),
.A2(n_11),
.B(n_15),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_241),
.B(n_15),
.C(n_13),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_245),
.A2(n_233),
.B1(n_235),
.B2(n_236),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_262),
.A2(n_12),
.B1(n_5),
.B2(n_6),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_264),
.B(n_265),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_SL g265 ( 
.A(n_249),
.B(n_228),
.Y(n_265)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_267),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_L g268 ( 
.A1(n_251),
.A2(n_232),
.B1(n_224),
.B2(n_238),
.Y(n_268)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_268),
.Y(n_284)
);

OR2x2_ASAP7_75t_L g269 ( 
.A(n_254),
.B(n_238),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_269),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_270),
.B(n_274),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_246),
.B(n_12),
.C(n_15),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_273),
.B(n_258),
.C(n_249),
.Y(n_277)
);

HB1xp67_ASAP7_75t_L g274 ( 
.A(n_260),
.Y(n_274)
);

AOI22xp33_ASAP7_75t_SL g275 ( 
.A1(n_271),
.A2(n_259),
.B1(n_256),
.B2(n_248),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_275),
.A2(n_285),
.B1(n_3),
.B2(n_5),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_277),
.B(n_265),
.Y(n_292)
);

AOI21xp5_ASAP7_75t_L g278 ( 
.A1(n_262),
.A2(n_258),
.B(n_252),
.Y(n_278)
);

OAI21xp5_ASAP7_75t_L g288 ( 
.A1(n_278),
.A2(n_282),
.B(n_264),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_SL g280 ( 
.A(n_269),
.B(n_252),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_280),
.B(n_286),
.Y(n_289)
);

OAI21xp5_ASAP7_75t_SL g282 ( 
.A1(n_272),
.A2(n_263),
.B(n_261),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_266),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_285)
);

AOI21x1_ASAP7_75t_SL g287 ( 
.A1(n_283),
.A2(n_270),
.B(n_267),
.Y(n_287)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_287),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_SL g299 ( 
.A(n_288),
.B(n_292),
.Y(n_299)
);

BUFx24_ASAP7_75t_SL g290 ( 
.A(n_282),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_290),
.B(n_291),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_276),
.B(n_273),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_293),
.A2(n_286),
.B1(n_281),
.B2(n_285),
.Y(n_298)
);

OAI21xp5_ASAP7_75t_L g294 ( 
.A1(n_284),
.A2(n_3),
.B(n_6),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_294),
.B(n_295),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_279),
.B(n_7),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_298),
.B(n_278),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_289),
.B(n_279),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_301),
.B(n_302),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_SL g302 ( 
.A(n_287),
.B(n_277),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_299),
.B(n_296),
.C(n_300),
.Y(n_303)
);

INVxp33_ASAP7_75t_SL g306 ( 
.A(n_303),
.Y(n_306)
);

INVxp67_ASAP7_75t_L g307 ( 
.A(n_306),
.Y(n_307)
);

OAI21xp5_ASAP7_75t_SL g308 ( 
.A1(n_307),
.A2(n_304),
.B(n_305),
.Y(n_308)
);

OAI21xp5_ASAP7_75t_L g309 ( 
.A1(n_308),
.A2(n_297),
.B(n_298),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_SL g310 ( 
.A(n_309),
.B(n_7),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_310),
.B(n_7),
.C(n_233),
.Y(n_311)
);


endmodule