module fake_jpeg_29658_n_100 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_100);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_100;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_1),
.Y(n_11)
);

NAND2xp5_ASAP7_75t_L g12 ( 
.A(n_4),
.B(n_2),
.Y(n_12)
);

CKINVDCx16_ASAP7_75t_R g13 ( 
.A(n_5),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_5),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_4),
.B(n_8),
.Y(n_15)
);

AND2x2_ASAP7_75t_SL g16 ( 
.A(n_0),
.B(n_6),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_10),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_1),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_21),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_24),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_SL g25 ( 
.A(n_12),
.B(n_3),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_SL g36 ( 
.A(n_25),
.B(n_29),
.Y(n_36)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_21),
.Y(n_26)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_26),
.Y(n_41)
);

INVx11_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_27),
.Y(n_39)
);

INVx2_ASAP7_75t_SL g28 ( 
.A(n_22),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_28),
.B(n_31),
.Y(n_33)
);

HB1xp67_ASAP7_75t_L g29 ( 
.A(n_17),
.Y(n_29)
);

NOR3xp33_ASAP7_75t_L g30 ( 
.A(n_16),
.B(n_12),
.C(n_13),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_30),
.Y(n_42)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_22),
.Y(n_31)
);

INVx5_ASAP7_75t_L g32 ( 
.A(n_23),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_32),
.B(n_23),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_30),
.B(n_25),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_34),
.B(n_15),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_SL g35 ( 
.A1(n_28),
.A2(n_11),
.B1(n_20),
.B2(n_16),
.Y(n_35)
);

AOI21xp5_ASAP7_75t_L g53 ( 
.A1(n_35),
.A2(n_29),
.B(n_18),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g37 ( 
.A1(n_26),
.A2(n_16),
.B1(n_20),
.B2(n_11),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_L g55 ( 
.A1(n_37),
.A2(n_31),
.B1(n_32),
.B2(n_27),
.Y(n_55)
);

INVxp67_ASAP7_75t_L g43 ( 
.A(n_40),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g63 ( 
.A(n_44),
.B(n_46),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_34),
.B(n_19),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_45),
.B(n_51),
.Y(n_58)
);

AOI21xp33_ASAP7_75t_L g46 ( 
.A1(n_37),
.A2(n_18),
.B(n_17),
.Y(n_46)
);

AND2x4_ASAP7_75t_L g47 ( 
.A(n_35),
.B(n_28),
.Y(n_47)
);

AO21x1_ASAP7_75t_L g59 ( 
.A1(n_47),
.A2(n_53),
.B(n_55),
.Y(n_59)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_41),
.Y(n_48)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_48),
.Y(n_60)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_39),
.Y(n_49)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_49),
.Y(n_67)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_41),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_50),
.B(n_0),
.Y(n_64)
);

INVx5_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

INVx13_ASAP7_75t_L g65 ( 
.A(n_52),
.Y(n_65)
);

CKINVDCx16_ASAP7_75t_R g54 ( 
.A(n_33),
.Y(n_54)
);

INVxp67_ASAP7_75t_L g57 ( 
.A(n_54),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_42),
.A2(n_24),
.B1(n_14),
.B2(n_19),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_56),
.A2(n_42),
.B1(n_14),
.B2(n_38),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_47),
.B(n_36),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_61),
.B(n_66),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_62),
.A2(n_53),
.B1(n_47),
.B2(n_43),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_64),
.B(n_7),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_47),
.B(n_0),
.Y(n_66)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_60),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_68),
.B(n_69),
.Y(n_78)
);

INVx13_ASAP7_75t_L g69 ( 
.A(n_65),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_70),
.A2(n_71),
.B1(n_75),
.B2(n_57),
.Y(n_81)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_60),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_72),
.A2(n_74),
.B1(n_67),
.B2(n_52),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_58),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_59),
.A2(n_43),
.B1(n_50),
.B2(n_44),
.Y(n_75)
);

XOR2xp5_ASAP7_75t_L g76 ( 
.A(n_61),
.B(n_51),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_76),
.B(n_66),
.C(n_62),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_77),
.B(n_79),
.C(n_80),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_76),
.B(n_63),
.C(n_75),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_71),
.B(n_63),
.C(n_57),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_81),
.B(n_82),
.Y(n_86)
);

AOI21xp5_ASAP7_75t_L g82 ( 
.A1(n_68),
.A2(n_59),
.B(n_72),
.Y(n_82)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_83),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_77),
.B(n_73),
.C(n_67),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_85),
.B(n_87),
.Y(n_92)
);

NOR3xp33_ASAP7_75t_L g87 ( 
.A(n_78),
.B(n_59),
.C(n_73),
.Y(n_87)
);

HB1xp67_ASAP7_75t_L g89 ( 
.A(n_88),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_89),
.B(n_91),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_86),
.B(n_7),
.Y(n_90)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_90),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_84),
.B(n_8),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_92),
.B(n_9),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_95),
.B(n_9),
.Y(n_96)
);

OR2x2_ASAP7_75t_L g98 ( 
.A(n_96),
.B(n_97),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_93),
.B(n_49),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_SL g99 ( 
.A1(n_98),
.A2(n_94),
.B(n_69),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_99),
.B(n_65),
.Y(n_100)
);


endmodule