module fake_jpeg_269_n_37 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_37);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_37;

wire n_13;
wire n_21;
wire n_33;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_34;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_12;
wire n_32;
wire n_8;
wire n_15;

NOR2xp33_ASAP7_75t_L g8 ( 
.A(n_5),
.B(n_6),
.Y(n_8)
);

NAND2xp5_ASAP7_75t_L g9 ( 
.A(n_0),
.B(n_5),
.Y(n_9)
);

BUFx6f_ASAP7_75t_L g10 ( 
.A(n_7),
.Y(n_10)
);

BUFx5_ASAP7_75t_L g11 ( 
.A(n_6),
.Y(n_11)
);

INVx3_ASAP7_75t_SL g12 ( 
.A(n_0),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_7),
.B(n_2),
.Y(n_13)
);

BUFx12f_ASAP7_75t_L g14 ( 
.A(n_3),
.Y(n_14)
);

OAI22xp5_ASAP7_75t_L g15 ( 
.A1(n_3),
.A2(n_4),
.B1(n_2),
.B2(n_1),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_12),
.Y(n_16)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_16),
.Y(n_25)
);

AOI22xp5_ASAP7_75t_L g17 ( 
.A1(n_15),
.A2(n_1),
.B1(n_4),
.B2(n_9),
.Y(n_17)
);

MAJIxp5_ASAP7_75t_L g26 ( 
.A(n_17),
.B(n_19),
.C(n_11),
.Y(n_26)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_18),
.Y(n_27)
);

AND2x2_ASAP7_75t_L g19 ( 
.A(n_9),
.B(n_13),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_8),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_20),
.B(n_21),
.Y(n_23)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

INVxp67_ASAP7_75t_L g29 ( 
.A(n_22),
.Y(n_29)
);

OAI21xp5_ASAP7_75t_L g24 ( 
.A1(n_19),
.A2(n_13),
.B(n_14),
.Y(n_24)
);

AOI21x1_ASAP7_75t_L g32 ( 
.A1(n_24),
.A2(n_26),
.B(n_28),
.Y(n_32)
);

XNOR2xp5_ASAP7_75t_SL g28 ( 
.A(n_19),
.B(n_14),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_SL g30 ( 
.A1(n_28),
.A2(n_17),
.B1(n_18),
.B2(n_27),
.Y(n_30)
);

OAI31xp33_ASAP7_75t_L g35 ( 
.A1(n_30),
.A2(n_11),
.A3(n_14),
.B(n_32),
.Y(n_35)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_25),
.Y(n_31)
);

OAI21x1_ASAP7_75t_L g36 ( 
.A1(n_31),
.A2(n_33),
.B(n_30),
.Y(n_36)
);

CKINVDCx16_ASAP7_75t_R g33 ( 
.A(n_29),
.Y(n_33)
);

OAI21xp5_ASAP7_75t_SL g34 ( 
.A1(n_32),
.A2(n_23),
.B(n_29),
.Y(n_34)
);

AOI22xp5_ASAP7_75t_L g37 ( 
.A1(n_34),
.A2(n_35),
.B1(n_36),
.B2(n_31),
.Y(n_37)
);


endmodule