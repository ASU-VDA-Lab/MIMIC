module fake_jpeg_11368_n_158 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_158);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_158;

wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_93;
wire n_54;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx13_ASAP7_75t_L g43 ( 
.A(n_5),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_14),
.Y(n_44)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_40),
.Y(n_45)
);

BUFx16f_ASAP7_75t_L g46 ( 
.A(n_9),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_16),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_39),
.Y(n_49)
);

INVx1_ASAP7_75t_SL g50 ( 
.A(n_17),
.Y(n_50)
);

INVxp67_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_12),
.Y(n_52)
);

BUFx16f_ASAP7_75t_L g53 ( 
.A(n_34),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_29),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_42),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_5),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_36),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_33),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_28),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_41),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_32),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_37),
.Y(n_62)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_30),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_31),
.Y(n_64)
);

BUFx12f_ASAP7_75t_L g65 ( 
.A(n_7),
.Y(n_65)
);

BUFx5_ASAP7_75t_L g66 ( 
.A(n_25),
.Y(n_66)
);

INVx11_ASAP7_75t_L g67 ( 
.A(n_43),
.Y(n_67)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_67),
.Y(n_81)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_44),
.Y(n_68)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_68),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_65),
.B(n_0),
.Y(n_69)
);

AOI21xp33_ASAP7_75t_L g82 ( 
.A1(n_69),
.A2(n_51),
.B(n_46),
.Y(n_82)
);

INVx5_ASAP7_75t_L g70 ( 
.A(n_65),
.Y(n_70)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_70),
.Y(n_84)
);

INVx6_ASAP7_75t_SL g71 ( 
.A(n_43),
.Y(n_71)
);

INVx13_ASAP7_75t_L g90 ( 
.A(n_71),
.Y(n_90)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_66),
.Y(n_72)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_72),
.B(n_74),
.Y(n_79)
);

BUFx12f_ASAP7_75t_L g73 ( 
.A(n_52),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_73),
.B(n_76),
.Y(n_85)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_48),
.Y(n_74)
);

AOI21xp33_ASAP7_75t_L g75 ( 
.A1(n_56),
.A2(n_0),
.B(n_1),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_75),
.B(n_69),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_57),
.B(n_1),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_77),
.B(n_46),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_71),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g105 ( 
.A(n_78),
.B(n_87),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_69),
.A2(n_44),
.B1(n_47),
.B2(n_49),
.Y(n_80)
);

AOI21xp5_ASAP7_75t_L g97 ( 
.A1(n_80),
.A2(n_82),
.B(n_89),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_74),
.B(n_61),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_86),
.B(n_91),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_73),
.B(n_60),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_68),
.A2(n_58),
.B1(n_47),
.B2(n_55),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_88),
.A2(n_55),
.B1(n_63),
.B2(n_45),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_70),
.A2(n_45),
.B1(n_58),
.B2(n_49),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_73),
.B(n_64),
.Y(n_91)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_83),
.Y(n_92)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_92),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_93),
.A2(n_111),
.B1(n_24),
.B2(n_15),
.Y(n_130)
);

OR2x2_ASAP7_75t_L g94 ( 
.A(n_90),
.B(n_67),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_L g113 ( 
.A1(n_94),
.A2(n_3),
.B(n_4),
.Y(n_113)
);

AOI21xp33_ASAP7_75t_L g119 ( 
.A1(n_95),
.A2(n_99),
.B(n_101),
.Y(n_119)
);

CKINVDCx14_ASAP7_75t_R g96 ( 
.A(n_79),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_96),
.B(n_102),
.Y(n_114)
);

INVx11_ASAP7_75t_L g98 ( 
.A(n_81),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_98),
.Y(n_122)
);

AOI32xp33_ASAP7_75t_L g99 ( 
.A1(n_79),
.A2(n_51),
.A3(n_62),
.B1(n_59),
.B2(n_54),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_85),
.B(n_50),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_100),
.B(n_104),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_81),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_83),
.Y(n_103)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_103),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_84),
.B(n_2),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_90),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_106),
.B(n_107),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_84),
.B(n_2),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_77),
.B(n_53),
.Y(n_108)
);

CKINVDCx16_ASAP7_75t_R g123 ( 
.A(n_108),
.Y(n_123)
);

INVx1_ASAP7_75t_SL g109 ( 
.A(n_81),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g115 ( 
.A(n_109),
.B(n_3),
.Y(n_115)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_81),
.Y(n_110)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_110),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_L g111 ( 
.A1(n_83),
.A2(n_72),
.B1(n_53),
.B2(n_6),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_113),
.B(n_115),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_L g116 ( 
.A1(n_109),
.A2(n_4),
.B1(n_6),
.B2(n_7),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_116),
.A2(n_118),
.B1(n_121),
.B2(n_10),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_L g117 ( 
.A1(n_97),
.A2(n_8),
.B(n_9),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_117),
.B(n_119),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_111),
.A2(n_8),
.B1(n_10),
.B2(n_11),
.Y(n_118)
);

AND2x6_ASAP7_75t_L g120 ( 
.A(n_98),
.B(n_22),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_SL g140 ( 
.A1(n_120),
.A2(n_129),
.B(n_18),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_94),
.A2(n_102),
.B1(n_110),
.B2(n_105),
.Y(n_121)
);

MAJx2_ASAP7_75t_L g125 ( 
.A(n_95),
.B(n_23),
.C(n_13),
.Y(n_125)
);

CKINVDCx16_ASAP7_75t_R g129 ( 
.A(n_98),
.Y(n_129)
);

A2O1A1Ixp33_ASAP7_75t_SL g131 ( 
.A1(n_130),
.A2(n_116),
.B(n_120),
.C(n_125),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_131),
.A2(n_141),
.B1(n_142),
.B2(n_123),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_124),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_132),
.B(n_134),
.Y(n_148)
);

INVx13_ASAP7_75t_L g133 ( 
.A(n_128),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_133),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_L g135 ( 
.A1(n_114),
.A2(n_122),
.B(n_126),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_135),
.B(n_140),
.Y(n_143)
);

INVx8_ASAP7_75t_L g138 ( 
.A(n_122),
.Y(n_138)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_138),
.Y(n_144)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_112),
.Y(n_139)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_139),
.Y(n_147)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_115),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_127),
.Y(n_142)
);

NOR2x1_ASAP7_75t_L g149 ( 
.A(n_145),
.B(n_135),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_L g152 ( 
.A(n_149),
.B(n_143),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_148),
.A2(n_131),
.B1(n_137),
.B2(n_136),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_150),
.A2(n_151),
.B1(n_144),
.B2(n_146),
.Y(n_153)
);

A2O1A1Ixp33_ASAP7_75t_SL g151 ( 
.A1(n_145),
.A2(n_131),
.B(n_138),
.C(n_133),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g154 ( 
.A(n_152),
.B(n_153),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_154),
.B(n_147),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_SL g156 ( 
.A1(n_155),
.A2(n_143),
.B(n_151),
.Y(n_156)
);

OAI321xp33_ASAP7_75t_L g157 ( 
.A1(n_156),
.A2(n_131),
.A3(n_20),
.B1(n_21),
.B2(n_26),
.C(n_27),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_157),
.B(n_19),
.Y(n_158)
);


endmodule