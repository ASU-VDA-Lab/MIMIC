module fake_jpeg_2820_n_121 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_8, n_15, n_7, n_121);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_8;
input n_15;
input n_7;

output n_121;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_21),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_12),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_7),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_SL g35 ( 
.A(n_31),
.B(n_16),
.Y(n_35)
);

CKINVDCx16_ASAP7_75t_R g36 ( 
.A(n_27),
.Y(n_36)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_0),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_29),
.Y(n_39)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_3),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_0),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_10),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_8),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_34),
.B(n_1),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_44),
.B(n_50),
.Y(n_57)
);

INVx5_ASAP7_75t_L g45 ( 
.A(n_41),
.Y(n_45)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_45),
.Y(n_54)
);

AOI21xp33_ASAP7_75t_SL g46 ( 
.A1(n_38),
.A2(n_14),
.B(n_28),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g60 ( 
.A(n_46),
.B(n_17),
.Y(n_60)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_43),
.Y(n_47)
);

INVx1_ASAP7_75t_SL g58 ( 
.A(n_47),
.Y(n_58)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_41),
.Y(n_48)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_48),
.Y(n_53)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_41),
.Y(n_49)
);

INVx13_ASAP7_75t_L g55 ( 
.A(n_49),
.Y(n_55)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_47),
.B(n_42),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_51),
.B(n_59),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_L g52 ( 
.A1(n_50),
.A2(n_43),
.B1(n_39),
.B2(n_38),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_52),
.A2(n_56),
.B1(n_49),
.B2(n_40),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_48),
.A2(n_40),
.B1(n_37),
.B2(n_42),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_45),
.B(n_39),
.Y(n_59)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_60),
.Y(n_66)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_55),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_61),
.Y(n_80)
);

BUFx4f_ASAP7_75t_SL g62 ( 
.A(n_54),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_62),
.B(n_63),
.Y(n_76)
);

INVx13_ASAP7_75t_L g63 ( 
.A(n_55),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_64),
.B(n_65),
.Y(n_73)
);

A2O1A1Ixp33_ASAP7_75t_SL g65 ( 
.A1(n_51),
.A2(n_36),
.B(n_33),
.C(n_32),
.Y(n_65)
);

INVx1_ASAP7_75t_SL g67 ( 
.A(n_54),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_67),
.B(n_13),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_53),
.Y(n_68)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_68),
.Y(n_74)
);

INVx5_ASAP7_75t_L g69 ( 
.A(n_53),
.Y(n_69)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_69),
.Y(n_81)
);

INVx11_ASAP7_75t_L g70 ( 
.A(n_58),
.Y(n_70)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_70),
.Y(n_84)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_58),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_71),
.B(n_60),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_72),
.B(n_57),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_75),
.B(n_77),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_78),
.B(n_79),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_72),
.B(n_35),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_65),
.B(n_1),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_82),
.B(n_83),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_66),
.B(n_2),
.Y(n_83)
);

XNOR2xp5_ASAP7_75t_L g85 ( 
.A(n_75),
.B(n_62),
.Y(n_85)
);

XNOR2xp5_ASAP7_75t_L g104 ( 
.A(n_85),
.B(n_89),
.Y(n_104)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_81),
.Y(n_87)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_87),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_SL g89 ( 
.A1(n_73),
.A2(n_64),
.B(n_65),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_76),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_91),
.B(n_95),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_L g92 ( 
.A1(n_76),
.A2(n_2),
.B(n_3),
.Y(n_92)
);

O2A1O1Ixp33_ASAP7_75t_L g102 ( 
.A1(n_92),
.A2(n_4),
.B(n_5),
.C(n_6),
.Y(n_102)
);

XOR2xp5_ASAP7_75t_L g93 ( 
.A(n_74),
.B(n_15),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_93),
.B(n_7),
.C(n_8),
.Y(n_103)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_80),
.Y(n_94)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_94),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_84),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_95)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_81),
.Y(n_96)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_96),
.Y(n_106)
);

A2O1A1O1Ixp25_ASAP7_75t_L g97 ( 
.A1(n_88),
.A2(n_19),
.B(n_26),
.C(n_25),
.D(n_24),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_97),
.B(n_101),
.Y(n_108)
);

A2O1A1O1Ixp25_ASAP7_75t_L g101 ( 
.A1(n_90),
.A2(n_11),
.B(n_23),
.C(n_22),
.D(n_20),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_102),
.B(n_105),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_103),
.B(n_92),
.C(n_93),
.Y(n_107)
);

INVx1_ASAP7_75t_SL g105 ( 
.A(n_85),
.Y(n_105)
);

XOR2xp5_ASAP7_75t_L g114 ( 
.A(n_107),
.B(n_110),
.Y(n_114)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_98),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_109),
.A2(n_100),
.B1(n_99),
.B2(n_86),
.Y(n_113)
);

XOR2xp5_ASAP7_75t_L g110 ( 
.A(n_104),
.B(n_106),
.Y(n_110)
);

NOR3xp33_ASAP7_75t_SL g112 ( 
.A(n_111),
.B(n_99),
.C(n_102),
.Y(n_112)
);

NOR3xp33_ASAP7_75t_SL g115 ( 
.A(n_112),
.B(n_108),
.C(n_110),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_113),
.B(n_30),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_115),
.Y(n_117)
);

BUFx24_ASAP7_75t_SL g118 ( 
.A(n_117),
.Y(n_118)
);

HB1xp67_ASAP7_75t_L g119 ( 
.A(n_118),
.Y(n_119)
);

NOR3xp33_ASAP7_75t_L g120 ( 
.A(n_119),
.B(n_116),
.C(n_112),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_SL g121 ( 
.A1(n_120),
.A2(n_114),
.B(n_9),
.Y(n_121)
);


endmodule