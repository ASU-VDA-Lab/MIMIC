module real_jpeg_17062_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_271;
wire n_47;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_541;
wire n_441;
wire n_557;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_498;
wire n_369;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_553;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_574;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_562;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_332;
wire n_366;
wire n_149;
wire n_578;
wire n_456;
wire n_259;
wire n_556;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_560;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_565;
wire n_466;
wire n_353;
wire n_453;
wire n_551;
wire n_230;
wire n_417;
wire n_428;
wire n_216;
wire n_128;
wire n_202;
wire n_483;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_464;
wire n_423;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_550;
wire n_233;
wire n_73;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_288;
wire n_83;
wire n_525;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_544;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_561;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_569;
wire n_335;
wire n_214;
wire n_113;
wire n_566;
wire n_543;
wire n_251;
wire n_459;
wire n_576;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_577;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_564;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_470;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_533;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_559;
wire n_232;
wire n_582;
wire n_448;
wire n_212;
wire n_284;
wire n_579;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_583;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_25;
wire n_480;
wire n_542;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_586;
wire n_405;
wire n_412;
wire n_572;
wire n_548;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_546;
wire n_172;
wire n_285;
wire n_531;
wire n_112;
wire n_554;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_563;
wire n_558;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_575;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_584;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_537;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_585;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_581;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_358;
wire n_534;
wire n_181;
wire n_256;
wire n_520;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_545;
wire n_484;
wire n_587;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_502;
wire n_418;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_400;
wire n_174;
wire n_388;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_571;
wire n_573;
wire n_379;
wire n_141;
wire n_555;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_570;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_313;
wire n_42;
wire n_94;
wire n_547;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_588;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_368;
wire n_100;
wire n_567;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_324;
wire n_86;
wire n_261;
wire n_549;
wire n_70;
wire n_568;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_580;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_552;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_0),
.Y(n_20)
);

AND2x2_ASAP7_75t_L g21 ( 
.A(n_0),
.B(n_22),
.Y(n_21)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_1),
.A2(n_71),
.B1(n_73),
.B2(n_74),
.Y(n_70)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_1),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g182 ( 
.A1(n_1),
.A2(n_74),
.B1(n_183),
.B2(n_188),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_1),
.A2(n_74),
.B1(n_268),
.B2(n_271),
.Y(n_267)
);

AOI22xp33_ASAP7_75t_SL g345 ( 
.A1(n_1),
.A2(n_74),
.B1(n_219),
.B2(n_346),
.Y(n_345)
);

BUFx3_ASAP7_75t_L g104 ( 
.A(n_2),
.Y(n_104)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_2),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_2),
.Y(n_116)
);

AOI21xp5_ASAP7_75t_L g18 ( 
.A1(n_3),
.A2(n_19),
.B(n_21),
.Y(n_18)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_4),
.Y(n_136)
);

BUFx5_ASAP7_75t_L g139 ( 
.A(n_4),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_4),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_4),
.Y(n_150)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_4),
.Y(n_442)
);

BUFx5_ASAP7_75t_L g447 ( 
.A(n_4),
.Y(n_447)
);

AOI22xp5_ASAP7_75t_SL g312 ( 
.A1(n_5),
.A2(n_313),
.B1(n_315),
.B2(n_317),
.Y(n_312)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_5),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_L g357 ( 
.A1(n_5),
.A2(n_317),
.B1(n_358),
.B2(n_361),
.Y(n_357)
);

OAI22xp5_ASAP7_75t_SL g470 ( 
.A1(n_5),
.A2(n_154),
.B1(n_317),
.B2(n_471),
.Y(n_470)
);

OAI22xp5_ASAP7_75t_SL g479 ( 
.A1(n_5),
.A2(n_317),
.B1(n_480),
.B2(n_484),
.Y(n_479)
);

AOI22xp33_ASAP7_75t_L g78 ( 
.A1(n_6),
.A2(n_79),
.B1(n_84),
.B2(n_85),
.Y(n_78)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_6),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_6),
.A2(n_84),
.B1(n_168),
.B2(n_170),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_L g224 ( 
.A1(n_6),
.A2(n_84),
.B1(n_225),
.B2(n_229),
.Y(n_224)
);

AOI22xp33_ASAP7_75t_SL g351 ( 
.A1(n_6),
.A2(n_84),
.B1(n_352),
.B2(n_354),
.Y(n_351)
);

AOI22xp33_ASAP7_75t_L g308 ( 
.A1(n_7),
.A2(n_71),
.B1(n_309),
.B2(n_310),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_7),
.Y(n_309)
);

AOI22xp33_ASAP7_75t_SL g397 ( 
.A1(n_7),
.A2(n_309),
.B1(n_398),
.B2(n_400),
.Y(n_397)
);

OAI22xp5_ASAP7_75t_SL g457 ( 
.A1(n_7),
.A2(n_309),
.B1(n_458),
.B2(n_459),
.Y(n_457)
);

OAI22xp5_ASAP7_75t_SL g498 ( 
.A1(n_7),
.A2(n_309),
.B1(n_499),
.B2(n_502),
.Y(n_498)
);

OAI32xp33_ASAP7_75t_L g327 ( 
.A1(n_8),
.A2(n_81),
.A3(n_328),
.B1(n_332),
.B2(n_336),
.Y(n_327)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_8),
.Y(n_335)
);

AOI22xp33_ASAP7_75t_L g365 ( 
.A1(n_8),
.A2(n_335),
.B1(n_366),
.B2(n_368),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_8),
.B(n_27),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_SL g474 ( 
.A(n_8),
.B(n_114),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_8),
.B(n_208),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g513 ( 
.A(n_8),
.B(n_132),
.Y(n_513)
);

AOI22xp33_ASAP7_75t_SL g528 ( 
.A1(n_8),
.A2(n_335),
.B1(n_358),
.B2(n_529),
.Y(n_528)
);

OAI32xp33_ASAP7_75t_L g533 ( 
.A1(n_8),
.A2(n_534),
.A3(n_537),
.B1(n_541),
.B2(n_546),
.Y(n_533)
);

BUFx5_ASAP7_75t_L g209 ( 
.A(n_9),
.Y(n_209)
);

BUFx5_ASAP7_75t_L g214 ( 
.A(n_9),
.Y(n_214)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_9),
.Y(n_253)
);

BUFx3_ASAP7_75t_L g375 ( 
.A(n_9),
.Y(n_375)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_10),
.Y(n_118)
);

BUFx5_ASAP7_75t_L g119 ( 
.A(n_10),
.Y(n_119)
);

BUFx3_ASAP7_75t_L g143 ( 
.A(n_10),
.Y(n_143)
);

INVx3_ASAP7_75t_L g158 ( 
.A(n_10),
.Y(n_158)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_10),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g228 ( 
.A(n_10),
.Y(n_228)
);

BUFx3_ASAP7_75t_L g232 ( 
.A(n_10),
.Y(n_232)
);

BUFx3_ASAP7_75t_L g545 ( 
.A(n_10),
.Y(n_545)
);

OAI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_11),
.A2(n_45),
.B1(n_46),
.B2(n_48),
.Y(n_44)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_11),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_11),
.A2(n_48),
.B1(n_93),
.B2(n_95),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_11),
.A2(n_48),
.B1(n_197),
.B2(n_199),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_11),
.A2(n_48),
.B1(n_256),
.B2(n_260),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_12),
.A2(n_275),
.B1(n_276),
.B2(n_277),
.Y(n_274)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_12),
.Y(n_276)
);

AOI22xp33_ASAP7_75t_L g320 ( 
.A1(n_12),
.A2(n_276),
.B1(n_321),
.B2(n_324),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_SL g463 ( 
.A1(n_12),
.A2(n_276),
.B1(n_464),
.B2(n_465),
.Y(n_463)
);

AOI22xp33_ASAP7_75t_SL g523 ( 
.A1(n_12),
.A2(n_276),
.B1(n_524),
.B2(n_526),
.Y(n_523)
);

OAI22xp5_ASAP7_75t_L g37 ( 
.A1(n_13),
.A2(n_38),
.B1(n_39),
.B2(n_42),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_13),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_13),
.A2(n_38),
.B1(n_124),
.B2(n_127),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_13),
.A2(n_38),
.B1(n_154),
.B2(n_159),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_13),
.A2(n_38),
.B1(n_216),
.B2(n_218),
.Y(n_215)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_14),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g342 ( 
.A(n_14),
.Y(n_342)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_15),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g134 ( 
.A(n_16),
.Y(n_134)
);

BUFx4f_ASAP7_75t_L g138 ( 
.A(n_16),
.Y(n_138)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_16),
.Y(n_264)
);

BUFx6f_ASAP7_75t_L g438 ( 
.A(n_16),
.Y(n_438)
);

BUFx8_ASAP7_75t_L g41 ( 
.A(n_17),
.Y(n_41)
);

BUFx5_ASAP7_75t_L g47 ( 
.A(n_17),
.Y(n_47)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_17),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g87 ( 
.A(n_17),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_SL g22 ( 
.A(n_23),
.B(n_588),
.Y(n_22)
);

OAI221xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_61),
.B1(n_64),
.B2(n_297),
.C(n_582),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g588 ( 
.A(n_24),
.B(n_61),
.Y(n_588)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_25),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_25),
.B(n_296),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g587 ( 
.A(n_25),
.B(n_296),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_43),
.Y(n_25)
);

OAI21x1_ASAP7_75t_SL g273 ( 
.A1(n_26),
.A2(n_50),
.B(n_274),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_37),
.Y(n_26)
);

OR2x6_ASAP7_75t_L g50 ( 
.A(n_27),
.B(n_51),
.Y(n_50)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_27),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_27),
.B(n_44),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_27),
.A2(n_49),
.B1(n_307),
.B2(n_311),
.Y(n_306)
);

AO22x2_ASAP7_75t_L g27 ( 
.A1(n_28),
.A2(n_31),
.B1(n_34),
.B2(n_36),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g325 ( 
.A(n_29),
.Y(n_325)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_29),
.Y(n_363)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g94 ( 
.A(n_30),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_30),
.Y(n_97)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_30),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g187 ( 
.A(n_30),
.Y(n_187)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_33),
.Y(n_36)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_33),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g399 ( 
.A(n_34),
.Y(n_399)
);

INVx6_ASAP7_75t_L g548 ( 
.A(n_34),
.Y(n_548)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx4_ASAP7_75t_L g130 ( 
.A(n_35),
.Y(n_130)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_37),
.Y(n_63)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_41),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g314 ( 
.A(n_41),
.Y(n_314)
);

OAI21xp5_ASAP7_75t_L g69 ( 
.A1(n_43),
.A2(n_62),
.B(n_70),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_44),
.B(n_49),
.Y(n_43)
);

INVx5_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_46),
.Y(n_73)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx1_ASAP7_75t_SL g49 ( 
.A(n_50),
.Y(n_49)
);

AOI21xp5_ASAP7_75t_L g61 ( 
.A1(n_50),
.A2(n_62),
.B(n_63),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_50),
.A2(n_62),
.B1(n_70),
.B2(n_78),
.Y(n_77)
);

OAI21xp5_ASAP7_75t_L g236 ( 
.A1(n_50),
.A2(n_63),
.B(n_237),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_SL g290 ( 
.A1(n_50),
.A2(n_78),
.B(n_237),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_SL g364 ( 
.A1(n_50),
.A2(n_62),
.B1(n_308),
.B2(n_365),
.Y(n_364)
);

OAI22x1_ASAP7_75t_SL g386 ( 
.A1(n_50),
.A2(n_62),
.B1(n_274),
.B2(n_312),
.Y(n_386)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_52),
.A2(n_53),
.B1(n_56),
.B2(n_58),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_53),
.Y(n_72)
);

INVx3_ASAP7_75t_L g275 ( 
.A(n_53),
.Y(n_275)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx4_ASAP7_75t_L g310 ( 
.A(n_54),
.Y(n_310)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_55),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_57),
.Y(n_83)
);

INVx5_ASAP7_75t_L g339 ( 
.A(n_57),
.Y(n_339)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

NAND3xp33_ASAP7_75t_L g64 ( 
.A(n_65),
.B(n_286),
.C(n_295),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_66),
.B(n_238),
.Y(n_65)
);

OAI21xp5_ASAP7_75t_L g583 ( 
.A1(n_66),
.A2(n_584),
.B(n_585),
.Y(n_583)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_67),
.B(n_173),
.Y(n_66)
);

NAND2xp33_ASAP7_75t_SL g585 ( 
.A(n_67),
.B(n_173),
.Y(n_585)
);

XNOR2xp5_ASAP7_75t_L g67 ( 
.A(n_68),
.B(n_165),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_69),
.A2(n_75),
.B1(n_76),
.B2(n_164),
.Y(n_68)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_69),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_69),
.B(n_131),
.C(n_166),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_69),
.A2(n_164),
.B1(n_176),
.B2(n_177),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_69),
.B(n_165),
.C(n_288),
.Y(n_287)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx1_ASAP7_75t_SL g75 ( 
.A(n_76),
.Y(n_75)
);

HB1xp67_ASAP7_75t_L g288 ( 
.A(n_76),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g76 ( 
.A(n_77),
.B(n_88),
.Y(n_76)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_77),
.Y(n_294)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

BUFx2_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx5_ASAP7_75t_L g278 ( 
.A(n_86),
.Y(n_278)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g316 ( 
.A(n_87),
.Y(n_316)
);

BUFx12f_ASAP7_75t_L g367 ( 
.A(n_87),
.Y(n_367)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_89),
.A2(n_90),
.B1(n_131),
.B2(n_163),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_89),
.B(n_163),
.C(n_294),
.Y(n_293)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

AO21x1_ASAP7_75t_L g90 ( 
.A1(n_91),
.A2(n_98),
.B(n_121),
.Y(n_90)
);

HB1xp67_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_92),
.B(n_114),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g281 ( 
.A(n_92),
.Y(n_281)
);

HB1xp67_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_94),
.Y(n_113)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

BUFx3_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_97),
.Y(n_169)
);

INVx4_ASAP7_75t_L g323 ( 
.A(n_97),
.Y(n_323)
);

INVx2_ASAP7_75t_L g536 ( 
.A(n_97),
.Y(n_536)
);

AOI21xp5_ASAP7_75t_L g166 ( 
.A1(n_98),
.A2(n_167),
.B(n_171),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_98),
.A2(n_114),
.B1(n_167),
.B2(n_181),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_L g291 ( 
.A1(n_98),
.A2(n_114),
.B(n_292),
.Y(n_291)
);

AOI21xp5_ASAP7_75t_L g318 ( 
.A1(n_98),
.A2(n_121),
.B(n_319),
.Y(n_318)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g280 ( 
.A1(n_99),
.A2(n_122),
.B1(n_182),
.B2(n_281),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_SL g356 ( 
.A1(n_99),
.A2(n_122),
.B1(n_320),
.B2(n_357),
.Y(n_356)
);

OAI21xp5_ASAP7_75t_SL g387 ( 
.A1(n_99),
.A2(n_123),
.B(n_172),
.Y(n_387)
);

OAI22xp5_ASAP7_75t_L g396 ( 
.A1(n_99),
.A2(n_122),
.B1(n_357),
.B2(n_397),
.Y(n_396)
);

OAI22xp5_ASAP7_75t_SL g527 ( 
.A1(n_99),
.A2(n_122),
.B1(n_397),
.B2(n_528),
.Y(n_527)
);

OR2x2_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_114),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_L g100 ( 
.A1(n_101),
.A2(n_105),
.B1(n_108),
.B2(n_113),
.Y(n_100)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_104),
.Y(n_120)
);

INVx8_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx4_ASAP7_75t_L g331 ( 
.A(n_106),
.Y(n_331)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_107),
.Y(n_126)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx5_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx2_ASAP7_75t_L g551 ( 
.A(n_111),
.Y(n_551)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g170 ( 
.A(n_113),
.Y(n_170)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_114),
.Y(n_122)
);

AO22x2_ASAP7_75t_L g114 ( 
.A1(n_115),
.A2(n_117),
.B1(n_119),
.B2(n_120),
.Y(n_114)
);

BUFx5_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx2_ASAP7_75t_L g458 ( 
.A(n_117),
.Y(n_458)
);

INVx4_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

BUFx12f_ASAP7_75t_L g151 ( 
.A(n_118),
.Y(n_151)
);

INVx4_ASAP7_75t_L g198 ( 
.A(n_118),
.Y(n_198)
);

BUFx6f_ASAP7_75t_L g272 ( 
.A(n_118),
.Y(n_272)
);

BUFx3_ASAP7_75t_L g444 ( 
.A(n_118),
.Y(n_444)
);

BUFx6f_ASAP7_75t_L g433 ( 
.A(n_119),
.Y(n_433)
);

NOR2xp67_ASAP7_75t_SL g121 ( 
.A(n_122),
.B(n_123),
.Y(n_121)
);

INVxp33_ASAP7_75t_SL g292 ( 
.A(n_123),
.Y(n_292)
);

INVx2_ASAP7_75t_L g531 ( 
.A(n_124),
.Y(n_531)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g334 ( 
.A(n_126),
.Y(n_334)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_126),
.Y(n_360)
);

INVx5_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx4_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx6_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_131),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_131),
.B(n_166),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_L g131 ( 
.A1(n_132),
.A2(n_140),
.B(n_152),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_132),
.B(n_196),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g377 ( 
.A(n_132),
.B(n_267),
.Y(n_377)
);

AOI22xp5_ASAP7_75t_L g452 ( 
.A1(n_132),
.A2(n_140),
.B1(n_453),
.B2(n_457),
.Y(n_452)
);

AOI22xp5_ASAP7_75t_L g469 ( 
.A1(n_132),
.A2(n_140),
.B1(n_457),
.B2(n_470),
.Y(n_469)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

AND2x2_ASAP7_75t_L g140 ( 
.A(n_133),
.B(n_141),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_133),
.B(n_153),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g265 ( 
.A1(n_133),
.A2(n_224),
.B1(n_233),
.B2(n_266),
.Y(n_265)
);

OAI22xp33_ASAP7_75t_L g521 ( 
.A1(n_133),
.A2(n_233),
.B1(n_522),
.B2(n_523),
.Y(n_521)
);

OA22x2_ASAP7_75t_L g133 ( 
.A1(n_134),
.A2(n_135),
.B1(n_137),
.B2(n_139),
.Y(n_133)
);

INVx3_ASAP7_75t_L g212 ( 
.A(n_134),
.Y(n_212)
);

INVx3_ASAP7_75t_L g220 ( 
.A(n_134),
.Y(n_220)
);

BUFx6f_ASAP7_75t_L g464 ( 
.A(n_134),
.Y(n_464)
);

INVx2_ASAP7_75t_L g501 ( 
.A(n_134),
.Y(n_501)
);

INVx4_ASAP7_75t_L g504 ( 
.A(n_134),
.Y(n_504)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_137),
.Y(n_508)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g217 ( 
.A(n_138),
.Y(n_217)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_138),
.Y(n_259)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_138),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_140),
.B(n_196),
.Y(n_195)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_140),
.Y(n_233)
);

AOI21xp5_ASAP7_75t_L g562 ( 
.A1(n_140),
.A2(n_193),
.B(n_563),
.Y(n_562)
);

OAI22xp33_ASAP7_75t_L g141 ( 
.A1(n_142),
.A2(n_144),
.B1(n_147),
.B2(n_151),
.Y(n_141)
);

INVx5_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx8_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVx4_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVx3_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVx6_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVxp67_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_SL g369 ( 
.A1(n_153),
.A2(n_233),
.B(n_234),
.Y(n_369)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVx5_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_158),
.Y(n_201)
);

INVx2_ASAP7_75t_L g540 ( 
.A(n_158),
.Y(n_540)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

INVx3_ASAP7_75t_SL g400 ( 
.A(n_170),
.Y(n_400)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_178),
.C(n_202),
.Y(n_173)
);

HB1xp67_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_175),
.A2(n_178),
.B1(n_179),
.B2(n_285),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_175),
.Y(n_285)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_176),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

OAI21xp33_ASAP7_75t_L g244 ( 
.A1(n_179),
.A2(n_180),
.B(n_192),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_192),
.Y(n_179)
);

INVxp67_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

BUFx3_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

INVx3_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

INVx3_ASAP7_75t_L g191 ( 
.A(n_187),
.Y(n_191)
);

INVx4_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_194),
.Y(n_192)
);

INVxp33_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_195),
.B(n_377),
.Y(n_376)
);

HB1xp67_ASAP7_75t_L g526 ( 
.A(n_197),
.Y(n_526)
);

INVx3_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

BUFx3_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVx2_ASAP7_75t_L g525 ( 
.A(n_200),
.Y(n_525)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_202),
.A2(n_203),
.B1(n_283),
.B2(n_284),
.Y(n_282)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

AOI21xp33_ASAP7_75t_L g203 ( 
.A1(n_204),
.A2(n_221),
.B(n_235),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g242 ( 
.A1(n_204),
.A2(n_205),
.B1(n_235),
.B2(n_236),
.Y(n_242)
);

OAI22xp33_ASAP7_75t_SL g412 ( 
.A1(n_204),
.A2(n_205),
.B1(n_223),
.B2(n_413),
.Y(n_412)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_205),
.B(n_223),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_L g205 ( 
.A1(n_206),
.A2(n_210),
.B(n_215),
.Y(n_205)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_206),
.Y(n_489)
);

INVx4_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

INVx6_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

BUFx12f_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_210),
.B(n_255),
.Y(n_254)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_210),
.Y(n_344)
);

AOI21xp5_ASAP7_75t_L g462 ( 
.A1(n_210),
.A2(n_463),
.B(n_467),
.Y(n_462)
);

AOI22xp33_ASAP7_75t_L g494 ( 
.A1(n_210),
.A2(n_335),
.B1(n_495),
.B2(n_498),
.Y(n_494)
);

AOI22xp5_ASAP7_75t_L g510 ( 
.A1(n_210),
.A2(n_479),
.B1(n_498),
.B2(n_511),
.Y(n_510)
);

AND2x2_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_213),
.Y(n_210)
);

INVx3_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_L g404 ( 
.A1(n_213),
.A2(n_254),
.B(n_345),
.Y(n_404)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_215),
.B(n_249),
.Y(n_248)
);

INVxp67_ASAP7_75t_L g553 ( 
.A(n_215),
.Y(n_553)
);

BUFx2_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

INVx4_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

INVxp33_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_222),
.B(n_242),
.Y(n_241)
);

INVxp67_ASAP7_75t_L g413 ( 
.A(n_223),
.Y(n_413)
);

OA21x2_ASAP7_75t_L g223 ( 
.A1(n_224),
.A2(n_233),
.B(n_234),
.Y(n_223)
);

BUFx2_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

HB1xp67_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_227),
.Y(n_270)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_227),
.Y(n_460)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_227),
.Y(n_473)
);

INVx6_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

BUFx6f_ASAP7_75t_L g456 ( 
.A(n_228),
.Y(n_456)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

BUFx2_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_282),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g584 ( 
.A(n_239),
.B(n_282),
.Y(n_584)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_243),
.C(n_245),
.Y(n_239)
);

HB1xp67_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g423 ( 
.A1(n_241),
.A2(n_243),
.B1(n_244),
.B2(n_424),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_241),
.Y(n_424)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g422 ( 
.A(n_245),
.B(n_423),
.Y(n_422)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_273),
.C(n_279),
.Y(n_245)
);

XNOR2x1_ASAP7_75t_L g414 ( 
.A(n_246),
.B(n_415),
.Y(n_414)
);

AND2x2_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_265),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_SL g381 ( 
.A(n_247),
.B(n_265),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_248),
.B(n_254),
.Y(n_247)
);

INVxp67_ASAP7_75t_L g467 ( 
.A(n_248),
.Y(n_467)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

BUFx6f_ASAP7_75t_L g350 ( 
.A(n_251),
.Y(n_350)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_251),
.Y(n_512)
);

BUFx6f_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

INVx3_ASAP7_75t_L g497 ( 
.A(n_253),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_255),
.B(n_373),
.Y(n_372)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

BUFx6f_ASAP7_75t_L g354 ( 
.A(n_261),
.Y(n_354)
);

BUFx6f_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

INVx4_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

BUFx6f_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

BUFx6f_ASAP7_75t_L g348 ( 
.A(n_264),
.Y(n_348)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g415 ( 
.A(n_273),
.B(n_280),
.Y(n_415)
);

INVx2_ASAP7_75t_L g368 ( 
.A(n_275),
.Y(n_368)
);

INVx3_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

HB1xp67_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

A2O1A1O1Ixp25_ASAP7_75t_SL g582 ( 
.A1(n_286),
.A2(n_295),
.B(n_583),
.C(n_586),
.D(n_587),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_SL g286 ( 
.A(n_287),
.B(n_289),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g586 ( 
.A(n_287),
.B(n_289),
.Y(n_586)
);

BUFx24_ASAP7_75t_SL g590 ( 
.A(n_289),
.Y(n_590)
);

FAx1_ASAP7_75t_SL g289 ( 
.A(n_290),
.B(n_291),
.CI(n_293),
.CON(n_289),
.SN(n_289)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_290),
.B(n_291),
.C(n_293),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_299),
.B(n_576),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g299 ( 
.A(n_300),
.B(n_425),
.Y(n_299)
);

NOR3xp33_ASAP7_75t_L g300 ( 
.A(n_301),
.B(n_407),
.C(n_419),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_302),
.B(n_389),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_303),
.B(n_378),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g577 ( 
.A(n_303),
.B(n_378),
.C(n_578),
.Y(n_577)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_304),
.B(n_355),
.C(n_370),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g405 ( 
.A(n_304),
.B(n_406),
.Y(n_405)
);

XOR2xp5_ASAP7_75t_L g304 ( 
.A(n_305),
.B(n_326),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_306),
.B(n_318),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g379 ( 
.A(n_306),
.B(n_318),
.C(n_326),
.Y(n_379)
);

INVxp67_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);

INVx4_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

BUFx3_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

BUFx6f_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_327),
.B(n_343),
.Y(n_326)
);

XOR2xp5_ASAP7_75t_L g394 ( 
.A(n_327),
.B(n_343),
.Y(n_394)
);

HB1xp67_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

INVx3_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_331),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_SL g332 ( 
.A(n_333),
.B(n_335),
.Y(n_332)
);

BUFx2_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_335),
.B(n_444),
.Y(n_443)
);

OAI21xp33_ASAP7_75t_SL g453 ( 
.A1(n_335),
.A2(n_443),
.B(n_454),
.Y(n_453)
);

NOR2xp33_ASAP7_75t_SL g541 ( 
.A(n_335),
.B(n_542),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_337),
.B(n_340),
.Y(n_336)
);

INVx4_ASAP7_75t_L g337 ( 
.A(n_338),
.Y(n_337)
);

INVx6_ASAP7_75t_L g338 ( 
.A(n_339),
.Y(n_338)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_341),
.Y(n_340)
);

BUFx6f_ASAP7_75t_L g341 ( 
.A(n_342),
.Y(n_341)
);

OAI22xp33_ASAP7_75t_SL g343 ( 
.A1(n_344),
.A2(n_345),
.B1(n_349),
.B2(n_351),
.Y(n_343)
);

OAI21xp5_ASAP7_75t_L g371 ( 
.A1(n_344),
.A2(n_351),
.B(n_372),
.Y(n_371)
);

OAI22xp5_ASAP7_75t_SL g477 ( 
.A1(n_344),
.A2(n_478),
.B1(n_488),
.B2(n_489),
.Y(n_477)
);

OAI21xp5_ASAP7_75t_L g552 ( 
.A1(n_344),
.A2(n_372),
.B(n_553),
.Y(n_552)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_347),
.Y(n_346)
);

INVx2_ASAP7_75t_L g347 ( 
.A(n_348),
.Y(n_347)
);

INVx2_ASAP7_75t_L g353 ( 
.A(n_348),
.Y(n_353)
);

INVx3_ASAP7_75t_L g466 ( 
.A(n_348),
.Y(n_466)
);

INVx2_ASAP7_75t_L g349 ( 
.A(n_350),
.Y(n_349)
);

INVx2_ASAP7_75t_L g352 ( 
.A(n_353),
.Y(n_352)
);

XNOR2xp5_ASAP7_75t_L g406 ( 
.A(n_355),
.B(n_370),
.Y(n_406)
);

MAJx2_ASAP7_75t_L g355 ( 
.A(n_356),
.B(n_364),
.C(n_369),
.Y(n_355)
);

XNOR2xp5_ASAP7_75t_L g392 ( 
.A(n_356),
.B(n_369),
.Y(n_392)
);

INVx8_ASAP7_75t_L g358 ( 
.A(n_359),
.Y(n_358)
);

BUFx6f_ASAP7_75t_L g359 ( 
.A(n_360),
.Y(n_359)
);

BUFx3_ASAP7_75t_L g361 ( 
.A(n_362),
.Y(n_361)
);

INVx2_ASAP7_75t_L g362 ( 
.A(n_363),
.Y(n_362)
);

XOR2xp5_ASAP7_75t_L g391 ( 
.A(n_364),
.B(n_392),
.Y(n_391)
);

INVx3_ASAP7_75t_L g366 ( 
.A(n_367),
.Y(n_366)
);

XOR2xp5_ASAP7_75t_L g370 ( 
.A(n_371),
.B(n_376),
.Y(n_370)
);

AND2x2_ASAP7_75t_L g384 ( 
.A(n_371),
.B(n_376),
.Y(n_384)
);

INVx5_ASAP7_75t_L g373 ( 
.A(n_374),
.Y(n_373)
);

INVx3_ASAP7_75t_L g374 ( 
.A(n_375),
.Y(n_374)
);

XNOR2xp5_ASAP7_75t_L g378 ( 
.A(n_379),
.B(n_380),
.Y(n_378)
);

MAJIxp5_ASAP7_75t_L g409 ( 
.A(n_379),
.B(n_382),
.C(n_388),
.Y(n_409)
);

OAI22xp5_ASAP7_75t_L g380 ( 
.A1(n_381),
.A2(n_382),
.B1(n_383),
.B2(n_388),
.Y(n_380)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_381),
.Y(n_388)
);

INVx2_ASAP7_75t_L g382 ( 
.A(n_383),
.Y(n_382)
);

XOR2xp5_ASAP7_75t_L g383 ( 
.A(n_384),
.B(n_385),
.Y(n_383)
);

MAJIxp5_ASAP7_75t_L g417 ( 
.A(n_384),
.B(n_386),
.C(n_387),
.Y(n_417)
);

XNOR2xp5_ASAP7_75t_L g385 ( 
.A(n_386),
.B(n_387),
.Y(n_385)
);

OR2x2_ASAP7_75t_L g389 ( 
.A(n_390),
.B(n_405),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g578 ( 
.A(n_390),
.B(n_405),
.Y(n_578)
);

MAJIxp5_ASAP7_75t_L g390 ( 
.A(n_391),
.B(n_393),
.C(n_395),
.Y(n_390)
);

XNOR2xp5_ASAP7_75t_L g572 ( 
.A(n_391),
.B(n_573),
.Y(n_572)
);

OAI22xp5_ASAP7_75t_SL g573 ( 
.A1(n_393),
.A2(n_394),
.B1(n_395),
.B2(n_574),
.Y(n_573)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_394),
.Y(n_393)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_395),
.Y(n_574)
);

MAJIxp5_ASAP7_75t_L g395 ( 
.A(n_396),
.B(n_401),
.C(n_403),
.Y(n_395)
);

XNOR2xp5_ASAP7_75t_L g565 ( 
.A(n_396),
.B(n_566),
.Y(n_565)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_399),
.Y(n_398)
);

AOI22xp5_ASAP7_75t_L g566 ( 
.A1(n_401),
.A2(n_402),
.B1(n_404),
.B2(n_567),
.Y(n_566)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_402),
.Y(n_401)
);

HB1xp67_ASAP7_75t_L g403 ( 
.A(n_404),
.Y(n_403)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_404),
.Y(n_567)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_408),
.Y(n_407)
);

A2O1A1O1Ixp25_ASAP7_75t_SL g576 ( 
.A1(n_408),
.A2(n_577),
.B(n_579),
.C(n_580),
.D(n_581),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_409),
.B(n_410),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_L g579 ( 
.A(n_409),
.B(n_410),
.Y(n_579)
);

AOI22xp33_ASAP7_75t_SL g410 ( 
.A1(n_411),
.A2(n_416),
.B1(n_417),
.B2(n_418),
.Y(n_410)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_411),
.Y(n_418)
);

XNOR2xp5_ASAP7_75t_L g411 ( 
.A(n_412),
.B(n_414),
.Y(n_411)
);

HB1xp67_ASAP7_75t_L g421 ( 
.A(n_412),
.Y(n_421)
);

MAJIxp5_ASAP7_75t_L g420 ( 
.A(n_414),
.B(n_416),
.C(n_421),
.Y(n_420)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_417),
.Y(n_416)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_419),
.Y(n_580)
);

AND2x2_ASAP7_75t_L g419 ( 
.A(n_420),
.B(n_422),
.Y(n_419)
);

NOR2xp33_ASAP7_75t_L g581 ( 
.A(n_420),
.B(n_422),
.Y(n_581)
);

OAI21x1_ASAP7_75t_L g425 ( 
.A1(n_426),
.A2(n_570),
.B(n_575),
.Y(n_425)
);

AOI21x1_ASAP7_75t_L g426 ( 
.A1(n_427),
.A2(n_555),
.B(n_569),
.Y(n_426)
);

OAI21x1_ASAP7_75t_SL g427 ( 
.A1(n_428),
.A2(n_517),
.B(n_554),
.Y(n_427)
);

AOI21xp5_ASAP7_75t_L g428 ( 
.A1(n_429),
.A2(n_475),
.B(n_516),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_430),
.B(n_461),
.Y(n_429)
);

NOR2xp33_ASAP7_75t_L g516 ( 
.A(n_430),
.B(n_461),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_431),
.B(n_451),
.Y(n_430)
);

OAI22xp5_ASAP7_75t_SL g490 ( 
.A1(n_431),
.A2(n_451),
.B1(n_452),
.B2(n_491),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_431),
.Y(n_491)
);

OAI32xp33_ASAP7_75t_L g431 ( 
.A1(n_432),
.A2(n_434),
.A3(n_439),
.B1(n_443),
.B2(n_445),
.Y(n_431)
);

INVx4_ASAP7_75t_L g432 ( 
.A(n_433),
.Y(n_432)
);

BUFx2_ASAP7_75t_L g434 ( 
.A(n_435),
.Y(n_434)
);

BUFx6f_ASAP7_75t_L g435 ( 
.A(n_436),
.Y(n_435)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_437),
.Y(n_436)
);

INVx2_ASAP7_75t_L g487 ( 
.A(n_437),
.Y(n_487)
);

INVx3_ASAP7_75t_L g437 ( 
.A(n_438),
.Y(n_437)
);

INVx2_ASAP7_75t_L g450 ( 
.A(n_438),
.Y(n_450)
);

HB1xp67_ASAP7_75t_L g439 ( 
.A(n_440),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_441),
.Y(n_440)
);

BUFx3_ASAP7_75t_L g441 ( 
.A(n_442),
.Y(n_441)
);

NOR2xp33_ASAP7_75t_L g445 ( 
.A(n_446),
.B(n_448),
.Y(n_445)
);

INVx4_ASAP7_75t_L g446 ( 
.A(n_447),
.Y(n_446)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_449),
.Y(n_448)
);

INVx5_ASAP7_75t_L g449 ( 
.A(n_450),
.Y(n_449)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_452),
.Y(n_451)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_455),
.Y(n_454)
);

INVx4_ASAP7_75t_L g455 ( 
.A(n_456),
.Y(n_455)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_460),
.Y(n_459)
);

XNOR2xp5_ASAP7_75t_L g461 ( 
.A(n_462),
.B(n_468),
.Y(n_461)
);

MAJIxp5_ASAP7_75t_L g518 ( 
.A(n_462),
.B(n_469),
.C(n_474),
.Y(n_518)
);

INVxp67_ASAP7_75t_L g488 ( 
.A(n_463),
.Y(n_488)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_466),
.Y(n_465)
);

XNOR2xp5_ASAP7_75t_L g468 ( 
.A(n_469),
.B(n_474),
.Y(n_468)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_470),
.Y(n_522)
);

INVx2_ASAP7_75t_L g471 ( 
.A(n_472),
.Y(n_471)
);

INVx2_ASAP7_75t_L g472 ( 
.A(n_473),
.Y(n_472)
);

OAI21xp5_ASAP7_75t_SL g475 ( 
.A1(n_476),
.A2(n_492),
.B(n_515),
.Y(n_475)
);

NOR2xp33_ASAP7_75t_L g476 ( 
.A(n_477),
.B(n_490),
.Y(n_476)
);

NAND2xp33_ASAP7_75t_SL g515 ( 
.A(n_477),
.B(n_490),
.Y(n_515)
);

INVxp67_ASAP7_75t_L g478 ( 
.A(n_479),
.Y(n_478)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_481),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_482),
.Y(n_481)
);

INVx2_ASAP7_75t_L g482 ( 
.A(n_483),
.Y(n_482)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_485),
.Y(n_484)
);

INVx3_ASAP7_75t_L g485 ( 
.A(n_486),
.Y(n_485)
);

INVx2_ASAP7_75t_L g486 ( 
.A(n_487),
.Y(n_486)
);

AOI21xp5_ASAP7_75t_L g492 ( 
.A1(n_493),
.A2(n_509),
.B(n_514),
.Y(n_492)
);

NOR2xp33_ASAP7_75t_SL g493 ( 
.A(n_494),
.B(n_505),
.Y(n_493)
);

INVx6_ASAP7_75t_L g495 ( 
.A(n_496),
.Y(n_495)
);

INVx6_ASAP7_75t_L g496 ( 
.A(n_497),
.Y(n_496)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_500),
.Y(n_499)
);

HB1xp67_ASAP7_75t_L g500 ( 
.A(n_501),
.Y(n_500)
);

INVx2_ASAP7_75t_L g502 ( 
.A(n_503),
.Y(n_502)
);

INVx3_ASAP7_75t_L g503 ( 
.A(n_504),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_SL g505 ( 
.A(n_506),
.B(n_507),
.Y(n_505)
);

BUFx3_ASAP7_75t_L g507 ( 
.A(n_508),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_SL g509 ( 
.A(n_510),
.B(n_513),
.Y(n_509)
);

NOR2xp33_ASAP7_75t_L g514 ( 
.A(n_510),
.B(n_513),
.Y(n_514)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_512),
.Y(n_511)
);

NOR2xp33_ASAP7_75t_L g517 ( 
.A(n_518),
.B(n_519),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_SL g554 ( 
.A(n_518),
.B(n_519),
.Y(n_554)
);

XNOR2xp5_ASAP7_75t_L g519 ( 
.A(n_520),
.B(n_532),
.Y(n_519)
);

XNOR2xp5_ASAP7_75t_L g520 ( 
.A(n_521),
.B(n_527),
.Y(n_520)
);

HB1xp67_ASAP7_75t_L g557 ( 
.A(n_521),
.Y(n_557)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_523),
.Y(n_563)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_525),
.Y(n_524)
);

HB1xp67_ASAP7_75t_L g558 ( 
.A(n_527),
.Y(n_558)
);

INVx2_ASAP7_75t_L g529 ( 
.A(n_530),
.Y(n_529)
);

INVx2_ASAP7_75t_L g530 ( 
.A(n_531),
.Y(n_530)
);

MAJIxp5_ASAP7_75t_L g556 ( 
.A(n_532),
.B(n_557),
.C(n_558),
.Y(n_556)
);

XOR2xp5_ASAP7_75t_L g532 ( 
.A(n_533),
.B(n_552),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_L g561 ( 
.A(n_533),
.B(n_552),
.Y(n_561)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_535),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_536),
.Y(n_535)
);

INVx3_ASAP7_75t_L g537 ( 
.A(n_538),
.Y(n_537)
);

INVx2_ASAP7_75t_L g538 ( 
.A(n_539),
.Y(n_538)
);

BUFx6f_ASAP7_75t_L g539 ( 
.A(n_540),
.Y(n_539)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_543),
.Y(n_542)
);

INVx2_ASAP7_75t_L g543 ( 
.A(n_544),
.Y(n_543)
);

INVx3_ASAP7_75t_L g544 ( 
.A(n_545),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_L g546 ( 
.A(n_547),
.B(n_549),
.Y(n_546)
);

INVx6_ASAP7_75t_L g547 ( 
.A(n_548),
.Y(n_547)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_550),
.Y(n_549)
);

HB1xp67_ASAP7_75t_L g550 ( 
.A(n_551),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g555 ( 
.A(n_556),
.B(n_559),
.Y(n_555)
);

NOR2xp33_ASAP7_75t_SL g569 ( 
.A(n_556),
.B(n_559),
.Y(n_569)
);

AOI22xp5_ASAP7_75t_L g559 ( 
.A1(n_560),
.A2(n_564),
.B1(n_565),
.B2(n_568),
.Y(n_559)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_560),
.Y(n_568)
);

XOR2x1_ASAP7_75t_SL g560 ( 
.A(n_561),
.B(n_562),
.Y(n_560)
);

MAJIxp5_ASAP7_75t_L g571 ( 
.A(n_561),
.B(n_562),
.C(n_564),
.Y(n_571)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_565),
.Y(n_564)
);

NOR2xp33_ASAP7_75t_L g570 ( 
.A(n_571),
.B(n_572),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_571),
.B(n_572),
.Y(n_575)
);


endmodule