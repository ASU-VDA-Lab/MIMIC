module fake_netlist_6_857_n_800 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_68, n_28, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_144, n_127, n_125, n_153, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_157, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_800);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_68;
input n_28;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_144;
input n_127;
input n_125;
input n_153;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_157;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_800;

wire n_591;
wire n_435;
wire n_793;
wire n_326;
wire n_256;
wire n_440;
wire n_587;
wire n_695;
wire n_507;
wire n_580;
wire n_762;
wire n_209;
wire n_367;
wire n_465;
wire n_760;
wire n_741;
wire n_680;
wire n_590;
wire n_625;
wire n_661;
wire n_223;
wire n_278;
wire n_362;
wire n_341;
wire n_226;
wire n_161;
wire n_208;
wire n_462;
wire n_607;
wire n_671;
wire n_726;
wire n_316;
wire n_419;
wire n_304;
wire n_212;
wire n_700;
wire n_694;
wire n_740;
wire n_578;
wire n_703;
wire n_365;
wire n_168;
wire n_384;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_342;
wire n_783;
wire n_725;
wire n_358;
wire n_160;
wire n_751;
wire n_449;
wire n_749;
wire n_798;
wire n_188;
wire n_310;
wire n_509;
wire n_186;
wire n_245;
wire n_368;
wire n_575;
wire n_677;
wire n_396;
wire n_495;
wire n_350;
wire n_585;
wire n_732;
wire n_568;
wire n_392;
wire n_442;
wire n_480;
wire n_724;
wire n_382;
wire n_673;
wire n_180;
wire n_628;
wire n_557;
wire n_349;
wire n_643;
wire n_233;
wire n_617;
wire n_698;
wire n_255;
wire n_739;
wire n_284;
wire n_400;
wire n_337;
wire n_214;
wire n_485;
wire n_443;
wire n_246;
wire n_768;
wire n_471;
wire n_289;
wire n_421;
wire n_781;
wire n_424;
wire n_789;
wire n_615;
wire n_181;
wire n_182;
wire n_238;
wire n_573;
wire n_769;
wire n_202;
wire n_320;
wire n_639;
wire n_676;
wire n_327;
wire n_794;
wire n_727;
wire n_369;
wire n_597;
wire n_685;
wire n_280;
wire n_287;
wire n_353;
wire n_610;
wire n_555;
wire n_389;
wire n_415;
wire n_230;
wire n_605;
wire n_461;
wire n_383;
wire n_669;
wire n_200;
wire n_447;
wire n_176;
wire n_198;
wire n_300;
wire n_222;
wire n_179;
wire n_248;
wire n_517;
wire n_718;
wire n_747;
wire n_667;
wire n_229;
wire n_542;
wire n_644;
wire n_682;
wire n_621;
wire n_305;
wire n_721;
wire n_750;
wire n_532;
wire n_742;
wire n_173;
wire n_535;
wire n_691;
wire n_250;
wire n_372;
wire n_468;
wire n_544;
wire n_504;
wire n_314;
wire n_378;
wire n_413;
wire n_377;
wire n_791;
wire n_183;
wire n_510;
wire n_375;
wire n_601;
wire n_338;
wire n_522;
wire n_466;
wire n_704;
wire n_748;
wire n_506;
wire n_763;
wire n_360;
wire n_603;
wire n_235;
wire n_536;
wire n_622;
wire n_191;
wire n_340;
wire n_710;
wire n_387;
wire n_452;
wire n_616;
wire n_658;
wire n_744;
wire n_344;
wire n_581;
wire n_428;
wire n_761;
wire n_785;
wire n_746;
wire n_609;
wire n_765;
wire n_432;
wire n_641;
wire n_693;
wire n_167;
wire n_631;
wire n_174;
wire n_516;
wire n_720;
wire n_525;
wire n_758;
wire n_611;
wire n_491;
wire n_656;
wire n_772;
wire n_797;
wire n_666;
wire n_371;
wire n_795;
wire n_770;
wire n_567;
wire n_189;
wire n_738;
wire n_405;
wire n_213;
wire n_538;
wire n_294;
wire n_302;
wire n_499;
wire n_380;
wire n_705;
wire n_647;
wire n_197;
wire n_343;
wire n_448;
wire n_494;
wire n_539;
wire n_493;
wire n_397;
wire n_614;
wire n_529;
wire n_445;
wire n_425;
wire n_684;
wire n_454;
wire n_218;
wire n_638;
wire n_234;
wire n_486;
wire n_381;
wire n_236;
wire n_653;
wire n_752;
wire n_172;
wire n_713;
wire n_648;
wire n_657;
wire n_576;
wire n_472;
wire n_270;
wire n_239;
wire n_414;
wire n_563;
wire n_782;
wire n_490;
wire n_290;
wire n_220;
wire n_224;
wire n_734;
wire n_708;
wire n_196;
wire n_402;
wire n_352;
wire n_668;
wire n_478;
wire n_626;
wire n_574;
wire n_779;
wire n_460;
wire n_417;
wire n_446;
wire n_498;
wire n_662;
wire n_374;
wire n_659;
wire n_709;
wire n_366;
wire n_777;
wire n_407;
wire n_450;
wire n_272;
wire n_526;
wire n_185;
wire n_712;
wire n_348;
wire n_711;
wire n_579;
wire n_376;
wire n_390;
wire n_473;
wire n_293;
wire n_334;
wire n_559;
wire n_370;
wire n_458;
wire n_232;
wire n_650;
wire n_163;
wire n_717;
wire n_330;
wire n_771;
wire n_470;
wire n_475;
wire n_298;
wire n_492;
wire n_281;
wire n_258;
wire n_551;
wire n_699;
wire n_456;
wire n_564;
wire n_260;
wire n_265;
wire n_313;
wire n_451;
wire n_624;
wire n_279;
wire n_686;
wire n_796;
wire n_252;
wire n_757;
wire n_228;
wire n_594;
wire n_565;
wire n_719;
wire n_356;
wire n_577;
wire n_166;
wire n_184;
wire n_552;
wire n_619;
wire n_216;
wire n_455;
wire n_521;
wire n_363;
wire n_572;
wire n_395;
wire n_592;
wire n_745;
wire n_654;
wire n_323;
wire n_606;
wire n_393;
wire n_411;
wire n_503;
wire n_716;
wire n_623;
wire n_599;
wire n_513;
wire n_776;
wire n_321;
wire n_645;
wire n_331;
wire n_227;
wire n_570;
wire n_731;
wire n_406;
wire n_483;
wire n_735;
wire n_204;
wire n_482;
wire n_755;
wire n_474;
wire n_527;
wire n_261;
wire n_608;
wire n_620;
wire n_420;
wire n_683;
wire n_630;
wire n_312;
wire n_394;
wire n_519;
wire n_541;
wire n_512;
wire n_164;
wire n_292;
wire n_307;
wire n_469;
wire n_433;
wire n_500;
wire n_792;
wire n_476;
wire n_714;
wire n_291;
wire n_219;
wire n_543;
wire n_357;
wire n_264;
wire n_263;
wire n_589;
wire n_481;
wire n_788;
wire n_325;
wire n_767;
wire n_329;
wire n_464;
wire n_600;
wire n_561;
wire n_477;
wire n_549;
wire n_533;
wire n_408;
wire n_237;
wire n_584;
wire n_244;
wire n_399;
wire n_243;
wire n_548;
wire n_282;
wire n_436;
wire n_211;
wire n_523;
wire n_175;
wire n_322;
wire n_707;
wire n_345;
wire n_409;
wire n_231;
wire n_354;
wire n_689;
wire n_799;
wire n_505;
wire n_240;
wire n_756;
wire n_319;
wire n_547;
wire n_537;
wire n_273;
wire n_558;
wire n_635;
wire n_787;
wire n_311;
wire n_403;
wire n_723;
wire n_253;
wire n_634;
wire n_583;
wire n_596;
wire n_546;
wire n_562;
wire n_249;
wire n_201;
wire n_386;
wire n_764;
wire n_556;
wire n_159;
wire n_162;
wire n_692;
wire n_733;
wire n_754;
wire n_487;
wire n_550;
wire n_241;
wire n_275;
wire n_553;
wire n_652;
wire n_560;
wire n_753;
wire n_642;
wire n_276;
wire n_569;
wire n_441;
wire n_221;
wire n_444;
wire n_586;
wire n_423;
wire n_737;
wire n_318;
wire n_303;
wire n_511;
wire n_715;
wire n_467;
wire n_306;
wire n_193;
wire n_269;
wire n_359;
wire n_346;
wire n_416;
wire n_530;
wire n_277;
wire n_520;
wire n_418;
wire n_618;
wire n_790;
wire n_582;
wire n_199;
wire n_266;
wire n_296;
wire n_674;
wire n_775;
wire n_571;
wire n_268;
wire n_271;
wire n_404;
wire n_651;
wire n_439;
wire n_217;
wire n_210;
wire n_299;
wire n_518;
wire n_206;
wire n_679;
wire n_453;
wire n_612;
wire n_633;
wire n_665;
wire n_333;
wire n_588;
wire n_215;
wire n_178;
wire n_247;
wire n_225;
wire n_308;
wire n_309;
wire n_759;
wire n_355;
wire n_426;
wire n_317;
wire n_632;
wire n_702;
wire n_431;
wire n_347;
wire n_459;
wire n_502;
wire n_328;
wire n_672;
wire n_534;
wire n_488;
wire n_429;
wire n_373;
wire n_195;
wire n_285;
wire n_497;
wire n_780;
wire n_773;
wire n_675;
wire n_257;
wire n_730;
wire n_655;
wire n_706;
wire n_786;
wire n_670;
wire n_203;
wire n_286;
wire n_254;
wire n_207;
wire n_242;
wire n_690;
wire n_401;
wire n_324;
wire n_743;
wire n_766;
wire n_335;
wire n_430;
wire n_463;
wire n_545;
wire n_489;
wire n_205;
wire n_604;
wire n_251;
wire n_301;
wire n_274;
wire n_636;
wire n_728;
wire n_681;
wire n_729;
wire n_774;
wire n_412;
wire n_640;
wire n_660;
wire n_267;
wire n_438;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_515;
wire n_288;
wire n_427;
wire n_479;
wire n_496;
wire n_598;
wire n_422;
wire n_696;
wire n_688;
wire n_722;
wire n_165;
wire n_351;
wire n_437;
wire n_259;
wire n_177;
wire n_540;
wire n_593;
wire n_514;
wire n_646;
wire n_528;
wire n_391;
wire n_457;
wire n_687;
wire n_697;
wire n_364;
wire n_637;
wire n_295;
wire n_385;
wire n_701;
wire n_629;
wire n_388;
wire n_190;
wire n_262;
wire n_484;
wire n_613;
wire n_736;
wire n_187;
wire n_501;
wire n_531;
wire n_361;
wire n_508;
wire n_663;
wire n_379;
wire n_170;
wire n_778;
wire n_332;
wire n_336;
wire n_410;
wire n_398;
wire n_566;
wire n_554;
wire n_602;
wire n_194;
wire n_664;
wire n_171;
wire n_678;
wire n_192;
wire n_169;
wire n_649;
wire n_283;

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_48),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_88),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_127),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_80),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_122),
.Y(n_163)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_125),
.Y(n_164)
);

INVxp67_ASAP7_75t_L g165 ( 
.A(n_100),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_54),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_112),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_150),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_59),
.Y(n_169)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_28),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_140),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_65),
.Y(n_172)
);

INVx1_ASAP7_75t_SL g173 ( 
.A(n_18),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_3),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_119),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_73),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_155),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_51),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_85),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_87),
.Y(n_180)
);

INVx2_ASAP7_75t_SL g181 ( 
.A(n_5),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_111),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_56),
.Y(n_183)
);

INVx1_ASAP7_75t_SL g184 ( 
.A(n_75),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_70),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_49),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_21),
.Y(n_187)
);

INVx1_ASAP7_75t_SL g188 ( 
.A(n_47),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_151),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_57),
.Y(n_190)
);

CKINVDCx16_ASAP7_75t_R g191 ( 
.A(n_52),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_90),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_157),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_156),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_92),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_38),
.Y(n_196)
);

CKINVDCx14_ASAP7_75t_R g197 ( 
.A(n_25),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_148),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_98),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_67),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_23),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_123),
.Y(n_202)
);

BUFx8_ASAP7_75t_SL g203 ( 
.A(n_105),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_15),
.Y(n_204)
);

BUFx3_ASAP7_75t_L g205 ( 
.A(n_126),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_13),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_36),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_102),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_0),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_69),
.Y(n_210)
);

BUFx10_ASAP7_75t_L g211 ( 
.A(n_145),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_4),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_63),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_9),
.Y(n_214)
);

BUFx2_ASAP7_75t_L g215 ( 
.A(n_174),
.Y(n_215)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_204),
.Y(n_216)
);

OAI22x1_ASAP7_75t_SL g217 ( 
.A1(n_206),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_159),
.Y(n_218)
);

AND2x4_ASAP7_75t_L g219 ( 
.A(n_205),
.B(n_1),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_197),
.A2(n_191),
.B1(n_214),
.B2(n_209),
.Y(n_220)
);

BUFx6f_ASAP7_75t_L g221 ( 
.A(n_205),
.Y(n_221)
);

BUFx6f_ASAP7_75t_L g222 ( 
.A(n_164),
.Y(n_222)
);

OAI22x1_ASAP7_75t_SL g223 ( 
.A1(n_212),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_223)
);

HB1xp67_ASAP7_75t_L g224 ( 
.A(n_181),
.Y(n_224)
);

INVx2_ASAP7_75t_SL g225 ( 
.A(n_211),
.Y(n_225)
);

AND2x4_ASAP7_75t_L g226 ( 
.A(n_164),
.B(n_5),
.Y(n_226)
);

INVx5_ASAP7_75t_L g227 ( 
.A(n_211),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_170),
.B(n_165),
.Y(n_228)
);

BUFx6f_ASAP7_75t_L g229 ( 
.A(n_170),
.Y(n_229)
);

INVx5_ASAP7_75t_L g230 ( 
.A(n_211),
.Y(n_230)
);

AOI22x1_ASAP7_75t_SL g231 ( 
.A1(n_159),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_231)
);

BUFx6f_ASAP7_75t_L g232 ( 
.A(n_162),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_163),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_168),
.B(n_6),
.Y(n_234)
);

INVx3_ASAP7_75t_L g235 ( 
.A(n_203),
.Y(n_235)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_175),
.Y(n_236)
);

BUFx3_ASAP7_75t_L g237 ( 
.A(n_178),
.Y(n_237)
);

BUFx3_ASAP7_75t_L g238 ( 
.A(n_203),
.Y(n_238)
);

OAI22x1_ASAP7_75t_L g239 ( 
.A1(n_182),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_239)
);

BUFx6f_ASAP7_75t_L g240 ( 
.A(n_183),
.Y(n_240)
);

BUFx2_ASAP7_75t_L g241 ( 
.A(n_169),
.Y(n_241)
);

BUFx3_ASAP7_75t_L g242 ( 
.A(n_185),
.Y(n_242)
);

AND2x2_ASAP7_75t_L g243 ( 
.A(n_197),
.B(n_10),
.Y(n_243)
);

INVx5_ASAP7_75t_L g244 ( 
.A(n_160),
.Y(n_244)
);

BUFx6f_ASAP7_75t_L g245 ( 
.A(n_186),
.Y(n_245)
);

INVx5_ASAP7_75t_L g246 ( 
.A(n_161),
.Y(n_246)
);

BUFx6f_ASAP7_75t_L g247 ( 
.A(n_193),
.Y(n_247)
);

INVx4_ASAP7_75t_L g248 ( 
.A(n_166),
.Y(n_248)
);

INVx2_ASAP7_75t_SL g249 ( 
.A(n_167),
.Y(n_249)
);

OA21x2_ASAP7_75t_L g250 ( 
.A1(n_194),
.A2(n_10),
.B(n_11),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_198),
.B(n_11),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_200),
.Y(n_252)
);

AND2x2_ASAP7_75t_L g253 ( 
.A(n_173),
.B(n_12),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_207),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_184),
.B(n_12),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_171),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_L g257 ( 
.A1(n_169),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_238),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_241),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_249),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_218),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_218),
.Y(n_262)
);

NOR2xp67_ASAP7_75t_L g263 ( 
.A(n_227),
.B(n_172),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_248),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_248),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_222),
.Y(n_266)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_222),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_215),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_244),
.Y(n_269)
);

HB1xp67_ASAP7_75t_L g270 ( 
.A(n_225),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_244),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_244),
.Y(n_272)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_222),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_R g274 ( 
.A(n_235),
.B(n_176),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_244),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_222),
.Y(n_276)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_229),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_246),
.Y(n_278)
);

BUFx3_ASAP7_75t_L g279 ( 
.A(n_221),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_246),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_R g281 ( 
.A(n_235),
.B(n_176),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_246),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_246),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_229),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_256),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_R g286 ( 
.A(n_243),
.B(n_177),
.Y(n_286)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_229),
.Y(n_287)
);

HB1xp67_ASAP7_75t_L g288 ( 
.A(n_227),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_227),
.Y(n_289)
);

HB1xp67_ASAP7_75t_L g290 ( 
.A(n_227),
.Y(n_290)
);

INVx5_ASAP7_75t_L g291 ( 
.A(n_229),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_221),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_230),
.Y(n_293)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_232),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_221),
.Y(n_295)
);

HB1xp67_ASAP7_75t_L g296 ( 
.A(n_230),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_230),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_230),
.Y(n_298)
);

BUFx10_ASAP7_75t_L g299 ( 
.A(n_219),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_221),
.Y(n_300)
);

INVxp33_ASAP7_75t_L g301 ( 
.A(n_224),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_236),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_220),
.B(n_14),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_237),
.Y(n_304)
);

INVx2_ASAP7_75t_L g305 ( 
.A(n_232),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_233),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_292),
.B(n_219),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_306),
.Y(n_308)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_267),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_285),
.B(n_253),
.Y(n_310)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_267),
.Y(n_311)
);

INVx3_ASAP7_75t_L g312 ( 
.A(n_279),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_295),
.Y(n_313)
);

NOR2xp67_ASAP7_75t_L g314 ( 
.A(n_291),
.B(n_228),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_300),
.B(n_252),
.Y(n_315)
);

INVxp33_ASAP7_75t_L g316 ( 
.A(n_301),
.Y(n_316)
);

INVxp67_ASAP7_75t_L g317 ( 
.A(n_270),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_279),
.B(n_254),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_260),
.B(n_228),
.Y(n_319)
);

INVxp67_ASAP7_75t_L g320 ( 
.A(n_259),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_264),
.B(n_255),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_265),
.B(n_255),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_286),
.B(n_232),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_266),
.B(n_232),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_276),
.B(n_240),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_284),
.B(n_240),
.Y(n_326)
);

INVx2_ASAP7_75t_SL g327 ( 
.A(n_304),
.Y(n_327)
);

INVx2_ASAP7_75t_SL g328 ( 
.A(n_268),
.Y(n_328)
);

INVxp67_ASAP7_75t_L g329 ( 
.A(n_303),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_SL g330 ( 
.A(n_301),
.B(n_226),
.Y(n_330)
);

INVx2_ASAP7_75t_SL g331 ( 
.A(n_299),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_294),
.Y(n_332)
);

BUFx5_ASAP7_75t_L g333 ( 
.A(n_302),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_269),
.B(n_271),
.Y(n_334)
);

AOI22xp5_ASAP7_75t_L g335 ( 
.A1(n_299),
.A2(n_257),
.B1(n_239),
.B2(n_226),
.Y(n_335)
);

INVx2_ASAP7_75t_L g336 ( 
.A(n_273),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_294),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_272),
.B(n_240),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_SL g339 ( 
.A(n_299),
.B(n_179),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_275),
.B(n_240),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_SL g341 ( 
.A(n_274),
.B(n_180),
.Y(n_341)
);

INVx2_ASAP7_75t_L g342 ( 
.A(n_273),
.Y(n_342)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_277),
.Y(n_343)
);

BUFx6f_ASAP7_75t_L g344 ( 
.A(n_277),
.Y(n_344)
);

AOI221xp5_ASAP7_75t_L g345 ( 
.A1(n_281),
.A2(n_257),
.B1(n_223),
.B2(n_217),
.C(n_234),
.Y(n_345)
);

INVxp67_ASAP7_75t_L g346 ( 
.A(n_288),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_278),
.B(n_245),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_280),
.B(n_245),
.Y(n_348)
);

INVx2_ASAP7_75t_L g349 ( 
.A(n_287),
.Y(n_349)
);

AND2x4_ASAP7_75t_L g350 ( 
.A(n_290),
.B(n_216),
.Y(n_350)
);

INVx8_ASAP7_75t_L g351 ( 
.A(n_258),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_282),
.B(n_245),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_283),
.B(n_245),
.Y(n_353)
);

BUFx6f_ASAP7_75t_L g354 ( 
.A(n_287),
.Y(n_354)
);

BUFx8_ASAP7_75t_L g355 ( 
.A(n_261),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_305),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_305),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_291),
.Y(n_358)
);

INVx2_ASAP7_75t_L g359 ( 
.A(n_291),
.Y(n_359)
);

BUFx6f_ASAP7_75t_SL g360 ( 
.A(n_262),
.Y(n_360)
);

INVx2_ASAP7_75t_L g361 ( 
.A(n_291),
.Y(n_361)
);

INVxp67_ASAP7_75t_L g362 ( 
.A(n_296),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_263),
.B(n_247),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_289),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_298),
.Y(n_365)
);

BUFx6f_ASAP7_75t_L g366 ( 
.A(n_293),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_SL g367 ( 
.A(n_297),
.B(n_188),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_292),
.B(n_247),
.Y(n_368)
);

INVx2_ASAP7_75t_L g369 ( 
.A(n_267),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_SL g370 ( 
.A(n_304),
.B(n_187),
.Y(n_370)
);

NAND2xp33_ASAP7_75t_L g371 ( 
.A(n_285),
.B(n_189),
.Y(n_371)
);

INVx2_ASAP7_75t_SL g372 ( 
.A(n_350),
.Y(n_372)
);

INVx2_ASAP7_75t_L g373 ( 
.A(n_309),
.Y(n_373)
);

BUFx6f_ASAP7_75t_L g374 ( 
.A(n_344),
.Y(n_374)
);

BUFx4_ASAP7_75t_L g375 ( 
.A(n_355),
.Y(n_375)
);

BUFx6f_ASAP7_75t_L g376 ( 
.A(n_344),
.Y(n_376)
);

INVx3_ASAP7_75t_L g377 ( 
.A(n_344),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_308),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_319),
.B(n_250),
.Y(n_379)
);

NAND2xp33_ASAP7_75t_SL g380 ( 
.A(n_316),
.B(n_331),
.Y(n_380)
);

INVx2_ASAP7_75t_SL g381 ( 
.A(n_350),
.Y(n_381)
);

INVx2_ASAP7_75t_L g382 ( 
.A(n_311),
.Y(n_382)
);

AOI22xp5_ASAP7_75t_L g383 ( 
.A1(n_321),
.A2(n_210),
.B1(n_192),
.B2(n_195),
.Y(n_383)
);

INVx2_ASAP7_75t_SL g384 ( 
.A(n_330),
.Y(n_384)
);

AND2x2_ASAP7_75t_L g385 ( 
.A(n_310),
.B(n_224),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_307),
.Y(n_386)
);

BUFx2_ASAP7_75t_L g387 ( 
.A(n_317),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_332),
.Y(n_388)
);

AND2x4_ASAP7_75t_L g389 ( 
.A(n_312),
.B(n_237),
.Y(n_389)
);

HB1xp67_ASAP7_75t_L g390 ( 
.A(n_346),
.Y(n_390)
);

INVx3_ASAP7_75t_L g391 ( 
.A(n_354),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_SL g392 ( 
.A(n_322),
.B(n_190),
.Y(n_392)
);

INVxp67_ASAP7_75t_L g393 ( 
.A(n_367),
.Y(n_393)
);

BUFx2_ASAP7_75t_L g394 ( 
.A(n_320),
.Y(n_394)
);

OAI221xp5_ASAP7_75t_L g395 ( 
.A1(n_335),
.A2(n_251),
.B1(n_234),
.B2(n_250),
.C(n_242),
.Y(n_395)
);

AOI22xp33_ASAP7_75t_L g396 ( 
.A1(n_333),
.A2(n_250),
.B1(n_251),
.B2(n_242),
.Y(n_396)
);

AND2x4_ASAP7_75t_SL g397 ( 
.A(n_366),
.B(n_247),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_SL g398 ( 
.A(n_327),
.B(n_196),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_337),
.Y(n_399)
);

INVxp67_ASAP7_75t_L g400 ( 
.A(n_318),
.Y(n_400)
);

OAI21xp33_ASAP7_75t_L g401 ( 
.A1(n_335),
.A2(n_213),
.B(n_208),
.Y(n_401)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_336),
.Y(n_402)
);

BUFx4f_ASAP7_75t_L g403 ( 
.A(n_351),
.Y(n_403)
);

BUFx3_ASAP7_75t_L g404 ( 
.A(n_351),
.Y(n_404)
);

HB1xp67_ASAP7_75t_L g405 ( 
.A(n_362),
.Y(n_405)
);

OR2x6_ASAP7_75t_SL g406 ( 
.A(n_345),
.B(n_231),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_333),
.B(n_323),
.Y(n_407)
);

INVx3_ASAP7_75t_L g408 ( 
.A(n_354),
.Y(n_408)
);

INVx1_ASAP7_75t_SL g409 ( 
.A(n_328),
.Y(n_409)
);

BUFx3_ASAP7_75t_L g410 ( 
.A(n_351),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_SL g411 ( 
.A(n_366),
.B(n_199),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_333),
.B(n_247),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_333),
.B(n_201),
.Y(n_413)
);

BUFx6f_ASAP7_75t_L g414 ( 
.A(n_354),
.Y(n_414)
);

AND2x4_ASAP7_75t_L g415 ( 
.A(n_312),
.B(n_202),
.Y(n_415)
);

INVx3_ASAP7_75t_L g416 ( 
.A(n_342),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_SL g417 ( 
.A(n_366),
.B(n_16),
.Y(n_417)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_343),
.Y(n_418)
);

BUFx4f_ASAP7_75t_L g419 ( 
.A(n_364),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_333),
.B(n_17),
.Y(n_420)
);

AND2x2_ASAP7_75t_L g421 ( 
.A(n_365),
.B(n_16),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_356),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_357),
.B(n_19),
.Y(n_423)
);

HB1xp67_ASAP7_75t_L g424 ( 
.A(n_329),
.Y(n_424)
);

NAND3xp33_ASAP7_75t_SL g425 ( 
.A(n_339),
.B(n_20),
.C(n_22),
.Y(n_425)
);

OR2x2_ASAP7_75t_L g426 ( 
.A(n_370),
.B(n_24),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_349),
.B(n_26),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_369),
.B(n_27),
.Y(n_428)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_313),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_315),
.Y(n_430)
);

NOR2xp33_ASAP7_75t_L g431 ( 
.A(n_371),
.B(n_29),
.Y(n_431)
);

AOI21xp5_ASAP7_75t_L g432 ( 
.A1(n_338),
.A2(n_30),
.B(n_31),
.Y(n_432)
);

INVx1_ASAP7_75t_SL g433 ( 
.A(n_334),
.Y(n_433)
);

BUFx3_ASAP7_75t_L g434 ( 
.A(n_355),
.Y(n_434)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_324),
.Y(n_435)
);

AND2x2_ASAP7_75t_L g436 ( 
.A(n_341),
.B(n_32),
.Y(n_436)
);

NOR3xp33_ASAP7_75t_SL g437 ( 
.A(n_340),
.B(n_352),
.C(n_347),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_368),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_325),
.Y(n_439)
);

INVx2_ASAP7_75t_L g440 ( 
.A(n_326),
.Y(n_440)
);

BUFx6f_ASAP7_75t_SL g441 ( 
.A(n_360),
.Y(n_441)
);

A2O1A1Ixp33_ASAP7_75t_L g442 ( 
.A1(n_386),
.A2(n_348),
.B(n_353),
.C(n_314),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_400),
.B(n_314),
.Y(n_443)
);

OR2x6_ASAP7_75t_L g444 ( 
.A(n_404),
.B(n_360),
.Y(n_444)
);

OAI22x1_ASAP7_75t_L g445 ( 
.A1(n_393),
.A2(n_358),
.B1(n_363),
.B2(n_359),
.Y(n_445)
);

OAI22xp5_ASAP7_75t_L g446 ( 
.A1(n_379),
.A2(n_361),
.B1(n_34),
.B2(n_35),
.Y(n_446)
);

NOR2xp33_ASAP7_75t_L g447 ( 
.A(n_433),
.B(n_33),
.Y(n_447)
);

O2A1O1Ixp33_ASAP7_75t_L g448 ( 
.A1(n_395),
.A2(n_37),
.B(n_39),
.C(n_40),
.Y(n_448)
);

AOI21xp5_ASAP7_75t_L g449 ( 
.A1(n_407),
.A2(n_41),
.B(n_42),
.Y(n_449)
);

AOI21xp5_ASAP7_75t_L g450 ( 
.A1(n_407),
.A2(n_396),
.B(n_379),
.Y(n_450)
);

A2O1A1Ixp33_ASAP7_75t_L g451 ( 
.A1(n_431),
.A2(n_43),
.B(n_44),
.C(n_45),
.Y(n_451)
);

BUFx6f_ASAP7_75t_L g452 ( 
.A(n_410),
.Y(n_452)
);

AND2x2_ASAP7_75t_L g453 ( 
.A(n_385),
.B(n_46),
.Y(n_453)
);

O2A1O1Ixp33_ASAP7_75t_L g454 ( 
.A1(n_395),
.A2(n_50),
.B(n_53),
.C(n_55),
.Y(n_454)
);

NOR3xp33_ASAP7_75t_L g455 ( 
.A(n_424),
.B(n_58),
.C(n_60),
.Y(n_455)
);

BUFx6f_ASAP7_75t_L g456 ( 
.A(n_374),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_400),
.B(n_61),
.Y(n_457)
);

NAND2xp33_ASAP7_75t_R g458 ( 
.A(n_437),
.B(n_62),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_378),
.Y(n_459)
);

OAI21xp33_ASAP7_75t_L g460 ( 
.A1(n_401),
.A2(n_64),
.B(n_66),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_430),
.B(n_68),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_388),
.Y(n_462)
);

AOI22xp5_ASAP7_75t_L g463 ( 
.A1(n_384),
.A2(n_71),
.B1(n_72),
.B2(n_74),
.Y(n_463)
);

BUFx6f_ASAP7_75t_L g464 ( 
.A(n_403),
.Y(n_464)
);

A2O1A1Ixp33_ASAP7_75t_SL g465 ( 
.A1(n_377),
.A2(n_76),
.B(n_77),
.C(n_78),
.Y(n_465)
);

CKINVDCx16_ASAP7_75t_R g466 ( 
.A(n_441),
.Y(n_466)
);

AND2x4_ASAP7_75t_L g467 ( 
.A(n_372),
.B(n_381),
.Y(n_467)
);

A2O1A1Ixp33_ASAP7_75t_L g468 ( 
.A1(n_438),
.A2(n_79),
.B(n_81),
.C(n_82),
.Y(n_468)
);

AOI21xp5_ASAP7_75t_L g469 ( 
.A1(n_413),
.A2(n_83),
.B(n_84),
.Y(n_469)
);

AOI21xp5_ASAP7_75t_L g470 ( 
.A1(n_413),
.A2(n_86),
.B(n_89),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_399),
.Y(n_471)
);

AOI21xp5_ASAP7_75t_L g472 ( 
.A1(n_412),
.A2(n_91),
.B(n_93),
.Y(n_472)
);

INVx2_ASAP7_75t_L g473 ( 
.A(n_373),
.Y(n_473)
);

NOR2xp33_ASAP7_75t_L g474 ( 
.A(n_433),
.B(n_94),
.Y(n_474)
);

NAND2xp33_ASAP7_75t_L g475 ( 
.A(n_436),
.B(n_95),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_439),
.B(n_96),
.Y(n_476)
);

INVx2_ASAP7_75t_L g477 ( 
.A(n_382),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_435),
.B(n_97),
.Y(n_478)
);

NOR2xp33_ASAP7_75t_L g479 ( 
.A(n_393),
.B(n_99),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_422),
.Y(n_480)
);

CKINVDCx5p33_ASAP7_75t_R g481 ( 
.A(n_403),
.Y(n_481)
);

NOR2xp33_ASAP7_75t_L g482 ( 
.A(n_409),
.B(n_101),
.Y(n_482)
);

AOI22x1_ASAP7_75t_L g483 ( 
.A1(n_440),
.A2(n_103),
.B1(n_104),
.B2(n_106),
.Y(n_483)
);

NOR2xp33_ASAP7_75t_L g484 ( 
.A(n_409),
.B(n_387),
.Y(n_484)
);

AOI21xp5_ASAP7_75t_L g485 ( 
.A1(n_412),
.A2(n_107),
.B(n_108),
.Y(n_485)
);

AOI21xp5_ASAP7_75t_L g486 ( 
.A1(n_420),
.A2(n_109),
.B(n_110),
.Y(n_486)
);

NAND3xp33_ASAP7_75t_SL g487 ( 
.A(n_383),
.B(n_113),
.C(n_114),
.Y(n_487)
);

AOI21xp5_ASAP7_75t_L g488 ( 
.A1(n_420),
.A2(n_115),
.B(n_116),
.Y(n_488)
);

BUFx6f_ASAP7_75t_L g489 ( 
.A(n_434),
.Y(n_489)
);

INVx3_ASAP7_75t_SL g490 ( 
.A(n_398),
.Y(n_490)
);

INVx3_ASAP7_75t_L g491 ( 
.A(n_389),
.Y(n_491)
);

A2O1A1Ixp33_ASAP7_75t_SL g492 ( 
.A1(n_377),
.A2(n_117),
.B(n_118),
.C(n_120),
.Y(n_492)
);

BUFx2_ASAP7_75t_L g493 ( 
.A(n_394),
.Y(n_493)
);

AOI33xp33_ASAP7_75t_L g494 ( 
.A1(n_421),
.A2(n_406),
.A3(n_389),
.B1(n_429),
.B2(n_415),
.B3(n_397),
.Y(n_494)
);

HB1xp67_ASAP7_75t_L g495 ( 
.A(n_390),
.Y(n_495)
);

BUFx6f_ASAP7_75t_L g496 ( 
.A(n_374),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_392),
.B(n_415),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_416),
.B(n_121),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_SL g499 ( 
.A(n_419),
.B(n_124),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_402),
.Y(n_500)
);

AO21x2_ASAP7_75t_L g501 ( 
.A1(n_450),
.A2(n_423),
.B(n_425),
.Y(n_501)
);

BUFx2_ASAP7_75t_SL g502 ( 
.A(n_464),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_SL g503 ( 
.A(n_484),
.B(n_419),
.Y(n_503)
);

AND2x4_ASAP7_75t_L g504 ( 
.A(n_491),
.B(n_426),
.Y(n_504)
);

AOI21xp5_ASAP7_75t_L g505 ( 
.A1(n_475),
.A2(n_414),
.B(n_376),
.Y(n_505)
);

INVx3_ASAP7_75t_L g506 ( 
.A(n_456),
.Y(n_506)
);

AOI22xp33_ASAP7_75t_L g507 ( 
.A1(n_453),
.A2(n_425),
.B1(n_417),
.B2(n_418),
.Y(n_507)
);

AND2x4_ASAP7_75t_L g508 ( 
.A(n_473),
.B(n_391),
.Y(n_508)
);

OAI21xp5_ASAP7_75t_L g509 ( 
.A1(n_461),
.A2(n_423),
.B(n_428),
.Y(n_509)
);

OAI21x1_ASAP7_75t_L g510 ( 
.A1(n_498),
.A2(n_428),
.B(n_427),
.Y(n_510)
);

INVx5_ASAP7_75t_L g511 ( 
.A(n_456),
.Y(n_511)
);

AO21x2_ASAP7_75t_L g512 ( 
.A1(n_442),
.A2(n_432),
.B(n_427),
.Y(n_512)
);

OAI21x1_ASAP7_75t_L g513 ( 
.A1(n_478),
.A2(n_432),
.B(n_408),
.Y(n_513)
);

BUFx10_ASAP7_75t_L g514 ( 
.A(n_482),
.Y(n_514)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_477),
.Y(n_515)
);

AO21x2_ASAP7_75t_L g516 ( 
.A1(n_476),
.A2(n_411),
.B(n_405),
.Y(n_516)
);

INVx2_ASAP7_75t_L g517 ( 
.A(n_462),
.Y(n_517)
);

OA21x2_ASAP7_75t_L g518 ( 
.A1(n_460),
.A2(n_416),
.B(n_408),
.Y(n_518)
);

INVx3_ASAP7_75t_L g519 ( 
.A(n_456),
.Y(n_519)
);

INVx2_ASAP7_75t_L g520 ( 
.A(n_471),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_459),
.B(n_391),
.Y(n_521)
);

BUFx12f_ASAP7_75t_L g522 ( 
.A(n_489),
.Y(n_522)
);

AOI22x1_ASAP7_75t_L g523 ( 
.A1(n_445),
.A2(n_414),
.B1(n_376),
.B2(n_374),
.Y(n_523)
);

AO21x2_ASAP7_75t_L g524 ( 
.A1(n_446),
.A2(n_414),
.B(n_376),
.Y(n_524)
);

OAI21x1_ASAP7_75t_L g525 ( 
.A1(n_469),
.A2(n_128),
.B(n_129),
.Y(n_525)
);

INVx2_ASAP7_75t_L g526 ( 
.A(n_480),
.Y(n_526)
);

AOI21x1_ASAP7_75t_L g527 ( 
.A1(n_457),
.A2(n_497),
.B(n_443),
.Y(n_527)
);

OAI21x1_ASAP7_75t_L g528 ( 
.A1(n_470),
.A2(n_130),
.B(n_131),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_447),
.B(n_474),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_479),
.B(n_380),
.Y(n_530)
);

BUFx2_ASAP7_75t_L g531 ( 
.A(n_493),
.Y(n_531)
);

BUFx3_ASAP7_75t_L g532 ( 
.A(n_452),
.Y(n_532)
);

AOI22xp33_ASAP7_75t_L g533 ( 
.A1(n_487),
.A2(n_500),
.B1(n_499),
.B2(n_455),
.Y(n_533)
);

INVx2_ASAP7_75t_L g534 ( 
.A(n_496),
.Y(n_534)
);

OAI21x1_ASAP7_75t_L g535 ( 
.A1(n_448),
.A2(n_132),
.B(n_133),
.Y(n_535)
);

OAI21x1_ASAP7_75t_L g536 ( 
.A1(n_454),
.A2(n_134),
.B(n_135),
.Y(n_536)
);

NOR2xp33_ASAP7_75t_L g537 ( 
.A(n_495),
.B(n_441),
.Y(n_537)
);

INVx5_ASAP7_75t_L g538 ( 
.A(n_496),
.Y(n_538)
);

NOR2xp67_ASAP7_75t_L g539 ( 
.A(n_449),
.B(n_136),
.Y(n_539)
);

INVx2_ASAP7_75t_L g540 ( 
.A(n_496),
.Y(n_540)
);

OAI21xp5_ASAP7_75t_L g541 ( 
.A1(n_451),
.A2(n_137),
.B(n_138),
.Y(n_541)
);

OAI21x1_ASAP7_75t_L g542 ( 
.A1(n_483),
.A2(n_139),
.B(n_141),
.Y(n_542)
);

OR2x6_ASAP7_75t_L g543 ( 
.A(n_444),
.B(n_375),
.Y(n_543)
);

BUFx6f_ASAP7_75t_L g544 ( 
.A(n_464),
.Y(n_544)
);

HB1xp67_ASAP7_75t_L g545 ( 
.A(n_467),
.Y(n_545)
);

INVx2_ASAP7_75t_L g546 ( 
.A(n_463),
.Y(n_546)
);

INVx2_ASAP7_75t_L g547 ( 
.A(n_452),
.Y(n_547)
);

OAI21x1_ASAP7_75t_L g548 ( 
.A1(n_486),
.A2(n_142),
.B(n_143),
.Y(n_548)
);

INVx3_ASAP7_75t_L g549 ( 
.A(n_490),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_517),
.Y(n_550)
);

BUFx8_ASAP7_75t_L g551 ( 
.A(n_522),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_517),
.Y(n_552)
);

AOI22xp5_ASAP7_75t_SL g553 ( 
.A1(n_529),
.A2(n_481),
.B1(n_466),
.B2(n_489),
.Y(n_553)
);

AND2x2_ASAP7_75t_L g554 ( 
.A(n_531),
.B(n_494),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_520),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_520),
.Y(n_556)
);

INVx2_ASAP7_75t_SL g557 ( 
.A(n_532),
.Y(n_557)
);

INVx3_ASAP7_75t_L g558 ( 
.A(n_511),
.Y(n_558)
);

OAI22xp5_ASAP7_75t_L g559 ( 
.A1(n_530),
.A2(n_444),
.B1(n_468),
.B2(n_488),
.Y(n_559)
);

AOI22xp33_ASAP7_75t_L g560 ( 
.A1(n_546),
.A2(n_485),
.B1(n_472),
.B2(n_458),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_526),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_526),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_515),
.Y(n_563)
);

AND2x4_ASAP7_75t_L g564 ( 
.A(n_504),
.B(n_144),
.Y(n_564)
);

NOR2xp33_ASAP7_75t_L g565 ( 
.A(n_503),
.B(n_146),
.Y(n_565)
);

OA21x2_ASAP7_75t_L g566 ( 
.A1(n_509),
.A2(n_492),
.B(n_465),
.Y(n_566)
);

INVx1_ASAP7_75t_SL g567 ( 
.A(n_531),
.Y(n_567)
);

BUFx6f_ASAP7_75t_L g568 ( 
.A(n_511),
.Y(n_568)
);

INVx6_ASAP7_75t_L g569 ( 
.A(n_522),
.Y(n_569)
);

AO21x1_ASAP7_75t_SL g570 ( 
.A1(n_541),
.A2(n_147),
.B(n_149),
.Y(n_570)
);

AND2x2_ASAP7_75t_L g571 ( 
.A(n_545),
.B(n_152),
.Y(n_571)
);

OAI21x1_ASAP7_75t_L g572 ( 
.A1(n_513),
.A2(n_153),
.B(n_154),
.Y(n_572)
);

AOI22xp33_ASAP7_75t_L g573 ( 
.A1(n_546),
.A2(n_158),
.B1(n_514),
.B2(n_501),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_515),
.Y(n_574)
);

OAI21x1_ASAP7_75t_L g575 ( 
.A1(n_513),
.A2(n_505),
.B(n_510),
.Y(n_575)
);

BUFx3_ASAP7_75t_L g576 ( 
.A(n_532),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_521),
.Y(n_577)
);

HB1xp67_ASAP7_75t_L g578 ( 
.A(n_511),
.Y(n_578)
);

AOI22xp33_ASAP7_75t_SL g579 ( 
.A1(n_549),
.A2(n_514),
.B1(n_502),
.B2(n_543),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_508),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_508),
.Y(n_581)
);

INVx2_ASAP7_75t_L g582 ( 
.A(n_508),
.Y(n_582)
);

AOI21x1_ASAP7_75t_L g583 ( 
.A1(n_527),
.A2(n_518),
.B(n_510),
.Y(n_583)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_508),
.Y(n_584)
);

INVxp33_ASAP7_75t_L g585 ( 
.A(n_537),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_534),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_534),
.Y(n_587)
);

OR2x2_ASAP7_75t_L g588 ( 
.A(n_549),
.B(n_547),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_540),
.Y(n_589)
);

BUFx3_ASAP7_75t_L g590 ( 
.A(n_544),
.Y(n_590)
);

CKINVDCx11_ASAP7_75t_R g591 ( 
.A(n_543),
.Y(n_591)
);

HB1xp67_ASAP7_75t_L g592 ( 
.A(n_511),
.Y(n_592)
);

OAI22xp33_ASAP7_75t_L g593 ( 
.A1(n_549),
.A2(n_543),
.B1(n_544),
.B2(n_538),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_L g594 ( 
.A(n_504),
.B(n_514),
.Y(n_594)
);

OAI22xp5_ASAP7_75t_L g595 ( 
.A1(n_507),
.A2(n_504),
.B1(n_533),
.B2(n_538),
.Y(n_595)
);

O2A1O1Ixp33_ASAP7_75t_L g596 ( 
.A1(n_595),
.A2(n_504),
.B(n_516),
.C(n_501),
.Y(n_596)
);

AO31x2_ASAP7_75t_L g597 ( 
.A1(n_559),
.A2(n_512),
.A3(n_524),
.B(n_501),
.Y(n_597)
);

NOR2xp33_ASAP7_75t_R g598 ( 
.A(n_569),
.B(n_544),
.Y(n_598)
);

HB1xp67_ASAP7_75t_L g599 ( 
.A(n_550),
.Y(n_599)
);

NAND2xp33_ASAP7_75t_R g600 ( 
.A(n_564),
.B(n_543),
.Y(n_600)
);

CKINVDCx20_ASAP7_75t_R g601 ( 
.A(n_551),
.Y(n_601)
);

INVx4_ASAP7_75t_SL g602 ( 
.A(n_568),
.Y(n_602)
);

INVx2_ASAP7_75t_L g603 ( 
.A(n_563),
.Y(n_603)
);

AND2x2_ASAP7_75t_L g604 ( 
.A(n_554),
.B(n_547),
.Y(n_604)
);

AND2x2_ASAP7_75t_L g605 ( 
.A(n_571),
.B(n_540),
.Y(n_605)
);

AND2x2_ASAP7_75t_L g606 ( 
.A(n_588),
.B(n_567),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_552),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_555),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_L g609 ( 
.A(n_577),
.B(n_516),
.Y(n_609)
);

CKINVDCx20_ASAP7_75t_R g610 ( 
.A(n_551),
.Y(n_610)
);

NAND2xp33_ASAP7_75t_R g611 ( 
.A(n_564),
.B(n_506),
.Y(n_611)
);

BUFx8_ASAP7_75t_SL g612 ( 
.A(n_576),
.Y(n_612)
);

CKINVDCx5p33_ASAP7_75t_R g613 ( 
.A(n_591),
.Y(n_613)
);

OR2x6_ASAP7_75t_L g614 ( 
.A(n_594),
.B(n_502),
.Y(n_614)
);

HB1xp67_ASAP7_75t_L g615 ( 
.A(n_576),
.Y(n_615)
);

AND2x4_ASAP7_75t_L g616 ( 
.A(n_564),
.B(n_544),
.Y(n_616)
);

AND2x2_ASAP7_75t_SL g617 ( 
.A(n_573),
.B(n_544),
.Y(n_617)
);

CKINVDCx12_ASAP7_75t_R g618 ( 
.A(n_553),
.Y(n_618)
);

INVx2_ASAP7_75t_L g619 ( 
.A(n_574),
.Y(n_619)
);

OAI21x1_ASAP7_75t_L g620 ( 
.A1(n_575),
.A2(n_525),
.B(n_528),
.Y(n_620)
);

BUFx2_ASAP7_75t_L g621 ( 
.A(n_557),
.Y(n_621)
);

CKINVDCx5p33_ASAP7_75t_R g622 ( 
.A(n_591),
.Y(n_622)
);

BUFx10_ASAP7_75t_L g623 ( 
.A(n_569),
.Y(n_623)
);

CKINVDCx20_ASAP7_75t_R g624 ( 
.A(n_569),
.Y(n_624)
);

NOR2x1p5_ASAP7_75t_L g625 ( 
.A(n_580),
.B(n_506),
.Y(n_625)
);

CKINVDCx5p33_ASAP7_75t_R g626 ( 
.A(n_579),
.Y(n_626)
);

NAND3xp33_ASAP7_75t_L g627 ( 
.A(n_560),
.B(n_539),
.C(n_523),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_L g628 ( 
.A(n_556),
.B(n_516),
.Y(n_628)
);

AND2x2_ASAP7_75t_L g629 ( 
.A(n_582),
.B(n_519),
.Y(n_629)
);

INVx2_ASAP7_75t_L g630 ( 
.A(n_574),
.Y(n_630)
);

OAI21x1_ASAP7_75t_L g631 ( 
.A1(n_572),
.A2(n_528),
.B(n_525),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g632 ( 
.A(n_561),
.B(n_527),
.Y(n_632)
);

NAND2xp33_ASAP7_75t_SL g633 ( 
.A(n_585),
.B(n_519),
.Y(n_633)
);

AOI22xp33_ASAP7_75t_L g634 ( 
.A1(n_570),
.A2(n_565),
.B1(n_585),
.B2(n_573),
.Y(n_634)
);

CKINVDCx5p33_ASAP7_75t_R g635 ( 
.A(n_590),
.Y(n_635)
);

INVx2_ASAP7_75t_L g636 ( 
.A(n_562),
.Y(n_636)
);

AO31x2_ASAP7_75t_L g637 ( 
.A1(n_565),
.A2(n_512),
.A3(n_524),
.B(n_535),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_586),
.Y(n_638)
);

AND2x2_ASAP7_75t_L g639 ( 
.A(n_584),
.B(n_519),
.Y(n_639)
);

NAND3xp33_ASAP7_75t_SL g640 ( 
.A(n_560),
.B(n_539),
.C(n_523),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_L g641 ( 
.A(n_584),
.B(n_518),
.Y(n_641)
);

NOR3xp33_ASAP7_75t_SL g642 ( 
.A(n_593),
.B(n_548),
.C(n_535),
.Y(n_642)
);

NOR2xp33_ASAP7_75t_L g643 ( 
.A(n_581),
.B(n_511),
.Y(n_643)
);

INVxp67_ASAP7_75t_SL g644 ( 
.A(n_611),
.Y(n_644)
);

AND2x2_ASAP7_75t_SL g645 ( 
.A(n_617),
.B(n_566),
.Y(n_645)
);

AOI22xp33_ASAP7_75t_L g646 ( 
.A1(n_634),
.A2(n_593),
.B1(n_536),
.B2(n_590),
.Y(n_646)
);

INVx2_ASAP7_75t_L g647 ( 
.A(n_628),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_628),
.Y(n_648)
);

AND2x2_ASAP7_75t_L g649 ( 
.A(n_609),
.B(n_608),
.Y(n_649)
);

HB1xp67_ASAP7_75t_L g650 ( 
.A(n_606),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_L g651 ( 
.A(n_609),
.B(n_589),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_632),
.Y(n_652)
);

HB1xp67_ASAP7_75t_L g653 ( 
.A(n_615),
.Y(n_653)
);

BUFx3_ASAP7_75t_L g654 ( 
.A(n_614),
.Y(n_654)
);

INVx2_ASAP7_75t_L g655 ( 
.A(n_641),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_599),
.B(n_587),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_632),
.Y(n_657)
);

OR2x2_ASAP7_75t_L g658 ( 
.A(n_597),
.B(n_524),
.Y(n_658)
);

INVxp67_ASAP7_75t_L g659 ( 
.A(n_621),
.Y(n_659)
);

HB1xp67_ASAP7_75t_L g660 ( 
.A(n_599),
.Y(n_660)
);

INVx2_ASAP7_75t_SL g661 ( 
.A(n_623),
.Y(n_661)
);

AND2x2_ASAP7_75t_L g662 ( 
.A(n_607),
.B(n_583),
.Y(n_662)
);

AND2x2_ASAP7_75t_L g663 ( 
.A(n_636),
.B(n_638),
.Y(n_663)
);

BUFx2_ASAP7_75t_L g664 ( 
.A(n_633),
.Y(n_664)
);

HB1xp67_ASAP7_75t_L g665 ( 
.A(n_604),
.Y(n_665)
);

BUFx3_ASAP7_75t_L g666 ( 
.A(n_614),
.Y(n_666)
);

OAI21xp33_ASAP7_75t_L g667 ( 
.A1(n_626),
.A2(n_642),
.B(n_627),
.Y(n_667)
);

AND2x4_ASAP7_75t_L g668 ( 
.A(n_616),
.B(n_548),
.Y(n_668)
);

INVx2_ASAP7_75t_L g669 ( 
.A(n_641),
.Y(n_669)
);

AND2x2_ASAP7_75t_L g670 ( 
.A(n_629),
.B(n_566),
.Y(n_670)
);

AND2x2_ASAP7_75t_L g671 ( 
.A(n_639),
.B(n_512),
.Y(n_671)
);

AND2x2_ASAP7_75t_L g672 ( 
.A(n_603),
.B(n_536),
.Y(n_672)
);

INVx2_ASAP7_75t_L g673 ( 
.A(n_597),
.Y(n_673)
);

INVxp67_ASAP7_75t_L g674 ( 
.A(n_612),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_619),
.Y(n_675)
);

AO21x2_ASAP7_75t_L g676 ( 
.A1(n_640),
.A2(n_542),
.B(n_578),
.Y(n_676)
);

INVx2_ASAP7_75t_L g677 ( 
.A(n_620),
.Y(n_677)
);

BUFx2_ASAP7_75t_L g678 ( 
.A(n_614),
.Y(n_678)
);

INVx2_ASAP7_75t_L g679 ( 
.A(n_637),
.Y(n_679)
);

OA21x2_ASAP7_75t_L g680 ( 
.A1(n_642),
.A2(n_542),
.B(n_578),
.Y(n_680)
);

AOI22xp33_ASAP7_75t_L g681 ( 
.A1(n_640),
.A2(n_592),
.B1(n_568),
.B2(n_558),
.Y(n_681)
);

AO21x2_ASAP7_75t_L g682 ( 
.A1(n_631),
.A2(n_592),
.B(n_558),
.Y(n_682)
);

HB1xp67_ASAP7_75t_L g683 ( 
.A(n_653),
.Y(n_683)
);

HB1xp67_ASAP7_75t_L g684 ( 
.A(n_660),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_662),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_662),
.Y(n_686)
);

AND2x2_ASAP7_75t_L g687 ( 
.A(n_649),
.B(n_637),
.Y(n_687)
);

AND2x2_ASAP7_75t_L g688 ( 
.A(n_649),
.B(n_637),
.Y(n_688)
);

AND2x2_ASAP7_75t_L g689 ( 
.A(n_645),
.B(n_596),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_650),
.B(n_630),
.Y(n_690)
);

OAI221xp5_ASAP7_75t_SL g691 ( 
.A1(n_667),
.A2(n_596),
.B1(n_618),
.B2(n_605),
.C(n_600),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_647),
.Y(n_692)
);

HB1xp67_ASAP7_75t_L g693 ( 
.A(n_665),
.Y(n_693)
);

AND2x2_ASAP7_75t_L g694 ( 
.A(n_645),
.B(n_616),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_663),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_L g696 ( 
.A(n_663),
.B(n_635),
.Y(n_696)
);

AND2x2_ASAP7_75t_L g697 ( 
.A(n_645),
.B(n_625),
.Y(n_697)
);

AOI22xp33_ASAP7_75t_L g698 ( 
.A1(n_667),
.A2(n_622),
.B1(n_613),
.B2(n_624),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_648),
.B(n_643),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_656),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_656),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_L g702 ( 
.A(n_648),
.B(n_623),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_L g703 ( 
.A(n_647),
.B(n_598),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_651),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_SL g705 ( 
.A(n_664),
.B(n_602),
.Y(n_705)
);

OR2x2_ASAP7_75t_L g706 ( 
.A(n_655),
.B(n_568),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_647),
.Y(n_707)
);

NAND3xp33_ASAP7_75t_L g708 ( 
.A(n_646),
.B(n_601),
.C(n_610),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_652),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_L g710 ( 
.A(n_651),
.B(n_602),
.Y(n_710)
);

INVxp67_ASAP7_75t_SL g711 ( 
.A(n_652),
.Y(n_711)
);

AND2x2_ASAP7_75t_L g712 ( 
.A(n_671),
.B(n_602),
.Y(n_712)
);

AND2x2_ASAP7_75t_L g713 ( 
.A(n_671),
.B(n_568),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_L g714 ( 
.A(n_675),
.B(n_511),
.Y(n_714)
);

AND2x2_ASAP7_75t_L g715 ( 
.A(n_687),
.B(n_669),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_684),
.Y(n_716)
);

AND2x2_ASAP7_75t_L g717 ( 
.A(n_687),
.B(n_669),
.Y(n_717)
);

HB1xp67_ASAP7_75t_L g718 ( 
.A(n_686),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_709),
.Y(n_719)
);

AND2x2_ASAP7_75t_L g720 ( 
.A(n_688),
.B(n_689),
.Y(n_720)
);

BUFx2_ASAP7_75t_L g721 ( 
.A(n_686),
.Y(n_721)
);

BUFx2_ASAP7_75t_L g722 ( 
.A(n_685),
.Y(n_722)
);

HB1xp67_ASAP7_75t_L g723 ( 
.A(n_683),
.Y(n_723)
);

INVx3_ASAP7_75t_L g724 ( 
.A(n_692),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_L g725 ( 
.A(n_693),
.B(n_670),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_SL g726 ( 
.A(n_697),
.B(n_664),
.Y(n_726)
);

AND2x2_ASAP7_75t_L g727 ( 
.A(n_688),
.B(n_689),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_709),
.Y(n_728)
);

AND2x2_ASAP7_75t_L g729 ( 
.A(n_695),
.B(n_669),
.Y(n_729)
);

AND2x2_ASAP7_75t_L g730 ( 
.A(n_694),
.B(n_655),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_711),
.Y(n_731)
);

OR2x2_ASAP7_75t_L g732 ( 
.A(n_692),
.B(n_658),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_700),
.Y(n_733)
);

BUFx2_ASAP7_75t_L g734 ( 
.A(n_707),
.Y(n_734)
);

OAI322xp33_ASAP7_75t_L g735 ( 
.A1(n_716),
.A2(n_701),
.A3(n_699),
.B1(n_690),
.B2(n_704),
.C1(n_702),
.C2(n_659),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_721),
.Y(n_736)
);

OR3x2_ASAP7_75t_L g737 ( 
.A(n_731),
.B(n_706),
.C(n_658),
.Y(n_737)
);

AOI22xp5_ASAP7_75t_L g738 ( 
.A1(n_726),
.A2(n_708),
.B1(n_697),
.B2(n_644),
.Y(n_738)
);

OR2x2_ASAP7_75t_L g739 ( 
.A(n_725),
.B(n_707),
.Y(n_739)
);

OAI32xp33_ASAP7_75t_L g740 ( 
.A1(n_723),
.A2(n_710),
.A3(n_696),
.B1(n_703),
.B2(n_705),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_721),
.Y(n_741)
);

AND2x4_ASAP7_75t_L g742 ( 
.A(n_722),
.B(n_694),
.Y(n_742)
);

AOI22xp5_ASAP7_75t_L g743 ( 
.A1(n_720),
.A2(n_698),
.B1(n_678),
.B2(n_668),
.Y(n_743)
);

HB1xp67_ASAP7_75t_L g744 ( 
.A(n_718),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_734),
.Y(n_745)
);

OAI22xp5_ASAP7_75t_L g746 ( 
.A1(n_737),
.A2(n_691),
.B1(n_727),
.B2(n_720),
.Y(n_746)
);

XOR2x2_ASAP7_75t_L g747 ( 
.A(n_738),
.B(n_727),
.Y(n_747)
);

OAI21xp5_ASAP7_75t_L g748 ( 
.A1(n_743),
.A2(n_733),
.B(n_719),
.Y(n_748)
);

OAI221xp5_ASAP7_75t_L g749 ( 
.A1(n_739),
.A2(n_674),
.B1(n_661),
.B2(n_678),
.C(n_728),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_744),
.Y(n_750)
);

OAI21xp33_ASAP7_75t_L g751 ( 
.A1(n_740),
.A2(n_730),
.B(n_732),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_L g752 ( 
.A(n_742),
.B(n_730),
.Y(n_752)
);

AND2x2_ASAP7_75t_L g753 ( 
.A(n_750),
.B(n_742),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_752),
.Y(n_754)
);

OAI221xp5_ASAP7_75t_L g755 ( 
.A1(n_751),
.A2(n_745),
.B1(n_741),
.B2(n_736),
.C(n_661),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_749),
.Y(n_756)
);

AOI21xp5_ASAP7_75t_L g757 ( 
.A1(n_746),
.A2(n_735),
.B(n_732),
.Y(n_757)
);

OAI221xp5_ASAP7_75t_SL g758 ( 
.A1(n_747),
.A2(n_681),
.B1(n_722),
.B2(n_666),
.C(n_654),
.Y(n_758)
);

NOR2xp33_ASAP7_75t_L g759 ( 
.A(n_756),
.B(n_748),
.Y(n_759)
);

AOI221xp5_ASAP7_75t_L g760 ( 
.A1(n_757),
.A2(n_734),
.B1(n_729),
.B2(n_724),
.C(n_715),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_754),
.Y(n_761)
);

AOI221xp5_ASAP7_75t_L g762 ( 
.A1(n_758),
.A2(n_729),
.B1(n_724),
.B2(n_717),
.C(n_715),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_753),
.Y(n_763)
);

AOI21xp5_ASAP7_75t_SL g764 ( 
.A1(n_759),
.A2(n_755),
.B(n_753),
.Y(n_764)
);

AND4x1_ASAP7_75t_L g765 ( 
.A(n_760),
.B(n_712),
.C(n_714),
.D(n_717),
.Y(n_765)
);

INVx8_ASAP7_75t_L g766 ( 
.A(n_763),
.Y(n_766)
);

A2O1A1Ixp33_ASAP7_75t_L g767 ( 
.A1(n_764),
.A2(n_762),
.B(n_766),
.C(n_761),
.Y(n_767)
);

OAI222xp33_ASAP7_75t_L g768 ( 
.A1(n_765),
.A2(n_712),
.B1(n_654),
.B2(n_666),
.C1(n_724),
.C2(n_713),
.Y(n_768)
);

NOR2xp33_ASAP7_75t_R g769 ( 
.A(n_766),
.B(n_654),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_769),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_767),
.Y(n_771)
);

NOR2x1_ASAP7_75t_L g772 ( 
.A(n_768),
.B(n_666),
.Y(n_772)
);

AOI22xp5_ASAP7_75t_L g773 ( 
.A1(n_767),
.A2(n_713),
.B1(n_668),
.B2(n_670),
.Y(n_773)
);

INVx2_ASAP7_75t_L g774 ( 
.A(n_769),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_771),
.B(n_673),
.Y(n_775)
);

BUFx2_ASAP7_75t_L g776 ( 
.A(n_774),
.Y(n_776)
);

NAND4xp25_ASAP7_75t_L g777 ( 
.A(n_770),
.B(n_668),
.C(n_675),
.D(n_706),
.Y(n_777)
);

NOR2xp67_ASAP7_75t_L g778 ( 
.A(n_773),
.B(n_538),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_772),
.Y(n_779)
);

NOR2x1_ASAP7_75t_L g780 ( 
.A(n_771),
.B(n_682),
.Y(n_780)
);

NAND2xp33_ASAP7_75t_R g781 ( 
.A(n_776),
.B(n_680),
.Y(n_781)
);

CKINVDCx5p33_ASAP7_75t_R g782 ( 
.A(n_779),
.Y(n_782)
);

CKINVDCx5p33_ASAP7_75t_R g783 ( 
.A(n_775),
.Y(n_783)
);

CKINVDCx5p33_ASAP7_75t_R g784 ( 
.A(n_778),
.Y(n_784)
);

AND3x1_ASAP7_75t_L g785 ( 
.A(n_780),
.B(n_679),
.C(n_673),
.Y(n_785)
);

INVx2_ASAP7_75t_L g786 ( 
.A(n_782),
.Y(n_786)
);

XNOR2xp5_ASAP7_75t_L g787 ( 
.A(n_783),
.B(n_784),
.Y(n_787)
);

OAI22xp5_ASAP7_75t_L g788 ( 
.A1(n_785),
.A2(n_777),
.B1(n_781),
.B2(n_673),
.Y(n_788)
);

OA22x2_ASAP7_75t_L g789 ( 
.A1(n_782),
.A2(n_679),
.B1(n_668),
.B2(n_677),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_782),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_L g791 ( 
.A(n_790),
.B(n_679),
.Y(n_791)
);

INVx2_ASAP7_75t_L g792 ( 
.A(n_786),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_L g793 ( 
.A(n_787),
.B(n_680),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_792),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_791),
.Y(n_795)
);

OAI221xp5_ASAP7_75t_L g796 ( 
.A1(n_794),
.A2(n_793),
.B1(n_788),
.B2(n_789),
.C(n_538),
.Y(n_796)
);

NAND3xp33_ASAP7_75t_L g797 ( 
.A(n_796),
.B(n_795),
.C(n_538),
.Y(n_797)
);

AOI22xp5_ASAP7_75t_SL g798 ( 
.A1(n_797),
.A2(n_680),
.B1(n_538),
.B2(n_672),
.Y(n_798)
);

AOI221xp5_ASAP7_75t_L g799 ( 
.A1(n_798),
.A2(n_677),
.B1(n_657),
.B2(n_672),
.C(n_682),
.Y(n_799)
);

AOI22xp33_ASAP7_75t_SL g800 ( 
.A1(n_799),
.A2(n_680),
.B1(n_682),
.B2(n_676),
.Y(n_800)
);


endmodule