module fake_jpeg_15221_n_114 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_114);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_114;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

INVx1_ASAP7_75t_L g12 ( 
.A(n_7),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_7),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_11),
.Y(n_14)
);

INVx3_ASAP7_75t_L g15 ( 
.A(n_8),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_4),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_2),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

INVx13_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_19),
.Y(n_26)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_20),
.B(n_0),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_SL g43 ( 
.A(n_27),
.B(n_29),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_19),
.Y(n_28)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_20),
.B(n_0),
.Y(n_29)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_30),
.Y(n_34)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_24),
.Y(n_31)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_SL g32 ( 
.A(n_25),
.B(n_1),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_32),
.B(n_33),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_24),
.B(n_1),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_33),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_SL g56 ( 
.A(n_35),
.B(n_41),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g40 ( 
.A1(n_29),
.A2(n_23),
.B1(n_15),
.B2(n_16),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_40),
.A2(n_42),
.B1(n_23),
.B2(n_16),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_32),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_SL g42 ( 
.A1(n_30),
.A2(n_23),
.B1(n_15),
.B2(n_24),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g44 ( 
.A(n_43),
.B(n_27),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_44),
.B(n_46),
.Y(n_64)
);

INVx1_ASAP7_75t_SL g45 ( 
.A(n_39),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_45),
.B(n_49),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_35),
.B(n_43),
.Y(n_46)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_38),
.Y(n_47)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_47),
.Y(n_61)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_38),
.Y(n_48)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_48),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_41),
.B(n_21),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g62 ( 
.A1(n_50),
.A2(n_51),
.B1(n_52),
.B2(n_14),
.Y(n_62)
);

OAI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_40),
.A2(n_42),
.B1(n_31),
.B2(n_17),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g52 ( 
.A1(n_36),
.A2(n_13),
.B1(n_17),
.B2(n_22),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_34),
.B(n_13),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_53),
.B(n_59),
.Y(n_71)
);

AND2x2_ASAP7_75t_L g54 ( 
.A(n_34),
.B(n_1),
.Y(n_54)
);

XNOR2xp5_ASAP7_75t_SL g69 ( 
.A(n_54),
.B(n_19),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_39),
.B(n_37),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_55),
.B(n_26),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g57 ( 
.A(n_37),
.B(n_26),
.C(n_28),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g70 ( 
.A(n_57),
.B(n_26),
.C(n_18),
.Y(n_70)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_58),
.Y(n_67)
);

INVxp67_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_62),
.B(n_66),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_54),
.A2(n_31),
.B1(n_28),
.B2(n_14),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_65),
.A2(n_45),
.B1(n_59),
.B2(n_55),
.Y(n_74)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_47),
.Y(n_68)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_68),
.Y(n_80)
);

OAI21xp5_ASAP7_75t_SL g75 ( 
.A1(n_69),
.A2(n_54),
.B(n_56),
.Y(n_75)
);

INVxp67_ASAP7_75t_L g73 ( 
.A(n_70),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_56),
.B(n_26),
.Y(n_72)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_72),
.Y(n_81)
);

XOR2xp5_ASAP7_75t_L g92 ( 
.A(n_74),
.B(n_75),
.Y(n_92)
);

AOI21xp5_ASAP7_75t_L g76 ( 
.A1(n_72),
.A2(n_48),
.B(n_57),
.Y(n_76)
);

OAI21xp5_ASAP7_75t_SL g85 ( 
.A1(n_76),
.A2(n_82),
.B(n_67),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_SL g77 ( 
.A1(n_66),
.A2(n_58),
.B(n_25),
.Y(n_77)
);

AOI21xp5_ASAP7_75t_L g91 ( 
.A1(n_77),
.A2(n_65),
.B(n_12),
.Y(n_91)
);

OR2x2_ASAP7_75t_L g78 ( 
.A(n_62),
.B(n_18),
.Y(n_78)
);

OAI21xp5_ASAP7_75t_L g86 ( 
.A1(n_78),
.A2(n_79),
.B(n_76),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_63),
.Y(n_82)
);

INVx13_ASAP7_75t_L g83 ( 
.A(n_68),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_83),
.B(n_61),
.Y(n_87)
);

AOI21xp5_ASAP7_75t_L g84 ( 
.A1(n_73),
.A2(n_61),
.B(n_63),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_84),
.A2(n_86),
.B1(n_91),
.B2(n_82),
.Y(n_94)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_85),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_87),
.B(n_89),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_75),
.B(n_81),
.C(n_70),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_88),
.B(n_90),
.C(n_77),
.Y(n_93)
);

AOI21xp5_ASAP7_75t_SL g89 ( 
.A1(n_81),
.A2(n_60),
.B(n_69),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_L g90 ( 
.A1(n_78),
.A2(n_64),
.B(n_71),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_93),
.B(n_21),
.C(n_12),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_SL g100 ( 
.A1(n_94),
.A2(n_96),
.B(n_98),
.Y(n_100)
);

MAJx2_ASAP7_75t_L g96 ( 
.A(n_92),
.B(n_78),
.C(n_74),
.Y(n_96)
);

A2O1A1O1Ixp25_ASAP7_75t_L g98 ( 
.A1(n_84),
.A2(n_80),
.B(n_83),
.C(n_67),
.D(n_18),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_95),
.B(n_80),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_99),
.B(n_2),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_97),
.B(n_22),
.Y(n_101)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_101),
.B(n_102),
.Y(n_107)
);

AND2x6_ASAP7_75t_L g102 ( 
.A(n_98),
.B(n_96),
.Y(n_102)
);

XOR2xp5_ASAP7_75t_L g104 ( 
.A(n_103),
.B(n_8),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_104),
.B(n_105),
.C(n_99),
.Y(n_108)
);

XOR2xp5_ASAP7_75t_L g105 ( 
.A(n_100),
.B(n_83),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_106),
.B(n_3),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_108),
.B(n_109),
.Y(n_111)
);

OAI31xp33_ASAP7_75t_L g110 ( 
.A1(n_107),
.A2(n_9),
.A3(n_10),
.B(n_5),
.Y(n_110)
);

AOI21xp5_ASAP7_75t_SL g112 ( 
.A1(n_110),
.A2(n_106),
.B(n_4),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_112),
.B(n_5),
.C(n_3),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_L g114 ( 
.A(n_113),
.B(n_111),
.Y(n_114)
);


endmodule