module real_jpeg_9865_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_176;
wire n_104;
wire n_194;
wire n_153;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_126;
wire n_13;
wire n_113;
wire n_155;
wire n_120;
wire n_199;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_188;
wire n_139;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_136;
wire n_44;
wire n_28;
wire n_208;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_172;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_203;
wire n_192;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_110;
wire n_61;
wire n_195;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_30;
wire n_204;
wire n_158;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_202;
wire n_179;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_206;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;
wire n_16;

BUFx24_ASAP7_75t_L g54 ( 
.A(n_0),
.Y(n_54)
);

BUFx12_ASAP7_75t_L g52 ( 
.A(n_1),
.Y(n_52)
);

BUFx10_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

AOI22xp33_ASAP7_75t_SL g25 ( 
.A1(n_4),
.A2(n_23),
.B1(n_26),
.B2(n_27),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_4),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_L g38 ( 
.A1(n_5),
.A2(n_23),
.B1(n_26),
.B2(n_39),
.Y(n_38)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_5),
.Y(n_39)
);

O2A1O1Ixp33_ASAP7_75t_L g43 ( 
.A1(n_5),
.A2(n_37),
.B(n_38),
.C(n_44),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_SL g44 ( 
.A(n_5),
.B(n_37),
.Y(n_44)
);

AOI21xp33_ASAP7_75t_L g142 ( 
.A1(n_5),
.A2(n_7),
.B(n_23),
.Y(n_142)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_6),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_SL g41 ( 
.A1(n_7),
.A2(n_34),
.B1(n_37),
.B2(n_42),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_7),
.Y(n_42)
);

AOI21xp5_ASAP7_75t_L g59 ( 
.A1(n_7),
.A2(n_49),
.B(n_60),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_7),
.B(n_49),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_7),
.A2(n_42),
.B1(n_53),
.B2(n_54),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_7),
.B(n_84),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_7),
.A2(n_23),
.B1(n_26),
.B2(n_42),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_7),
.B(n_69),
.Y(n_163)
);

O2A1O1Ixp33_ASAP7_75t_L g176 ( 
.A1(n_7),
.A2(n_9),
.B(n_53),
.C(n_177),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g48 ( 
.A1(n_8),
.A2(n_11),
.B1(n_49),
.B2(n_50),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_8),
.Y(n_50)
);

OAI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_8),
.A2(n_50),
.B1(n_53),
.B2(n_54),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_8),
.A2(n_23),
.B1(n_26),
.B2(n_50),
.Y(n_138)
);

OAI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_8),
.A2(n_34),
.B1(n_37),
.B2(n_50),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_9),
.A2(n_34),
.B1(n_37),
.B2(n_71),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_9),
.Y(n_71)
);

A2O1A1Ixp33_ASAP7_75t_L g75 ( 
.A1(n_9),
.A2(n_53),
.B(n_70),
.C(n_76),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_9),
.B(n_53),
.Y(n_76)
);

OAI22xp33_ASAP7_75t_SL g29 ( 
.A1(n_10),
.A2(n_23),
.B1(n_26),
.B2(n_30),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_10),
.Y(n_30)
);

OAI22xp33_ASAP7_75t_SL g33 ( 
.A1(n_10),
.A2(n_30),
.B1(n_34),
.B2(n_37),
.Y(n_33)
);

AOI22xp33_ASAP7_75t_L g78 ( 
.A1(n_10),
.A2(n_30),
.B1(n_53),
.B2(n_54),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_10),
.A2(n_11),
.B1(n_30),
.B2(n_49),
.Y(n_86)
);

INVx2_ASAP7_75t_SL g49 ( 
.A(n_11),
.Y(n_49)
);

XNOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_129),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_127),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_15),
.Y(n_14)
);

AND2x2_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_110),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_16),
.B(n_110),
.Y(n_128)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_79),
.Y(n_16)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_45),
.Y(n_17)
);

XOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_31),
.Y(n_18)
);

OAI21xp5_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_25),
.B(n_28),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_20),
.B(n_103),
.Y(n_102)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_20),
.Y(n_126)
);

AOI21xp5_ASAP7_75t_L g175 ( 
.A1(n_20),
.A2(n_21),
.B(n_125),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_23),
.Y(n_20)
);

OAI21xp5_ASAP7_75t_L g100 ( 
.A1(n_21),
.A2(n_25),
.B(n_101),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_21),
.B(n_42),
.Y(n_155)
);

CKINVDCx16_ASAP7_75t_R g21 ( 
.A(n_22),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_SL g28 ( 
.A(n_22),
.B(n_29),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_22),
.B(n_138),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_22),
.B(n_124),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_23),
.Y(n_26)
);

BUFx24_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_SL g154 ( 
.A(n_26),
.B(n_155),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_28),
.B(n_123),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_28),
.B(n_151),
.Y(n_150)
);

INVxp33_ASAP7_75t_L g103 ( 
.A(n_29),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_32),
.B(n_40),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_32),
.B(n_166),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g32 ( 
.A(n_33),
.B(n_38),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_33),
.B(n_43),
.Y(n_182)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_34),
.Y(n_37)
);

A2O1A1Ixp33_ASAP7_75t_L g141 ( 
.A1(n_34),
.A2(n_39),
.B(n_42),
.C(n_142),
.Y(n_141)
);

INVx11_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx13_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

OAI21xp33_ASAP7_75t_L g177 ( 
.A1(n_37),
.A2(n_42),
.B(n_71),
.Y(n_177)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_38),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_38),
.B(n_146),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_38),
.B(n_41),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_40),
.B(n_145),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_41),
.B(n_43),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_41),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_42),
.B(n_64),
.Y(n_149)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_43),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_43),
.B(n_146),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g45 ( 
.A(n_46),
.B(n_61),
.C(n_66),
.Y(n_45)
);

XNOR2xp5_ASAP7_75t_SL g112 ( 
.A(n_46),
.B(n_113),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_47),
.B(n_56),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_48),
.B(n_51),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_48),
.Y(n_89)
);

A2O1A1Ixp33_ASAP7_75t_L g57 ( 
.A1(n_49),
.A2(n_51),
.B(n_52),
.C(n_58),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_49),
.B(n_52),
.Y(n_58)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_51),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g51 ( 
.A1(n_52),
.A2(n_53),
.B1(n_54),
.B2(n_55),
.Y(n_51)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_52),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_53),
.B(n_55),
.Y(n_106)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_54),
.A2(n_106),
.B1(n_107),
.B2(n_108),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g56 ( 
.A(n_57),
.B(n_59),
.Y(n_56)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_57),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_58),
.Y(n_108)
);

CKINVDCx14_ASAP7_75t_R g107 ( 
.A(n_60),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_61),
.A2(n_62),
.B1(n_66),
.B2(n_67),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_62),
.Y(n_61)
);

AOI21xp5_ASAP7_75t_SL g62 ( 
.A1(n_63),
.A2(n_64),
.B(n_65),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_67),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_68),
.B(n_73),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_68),
.B(n_185),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_69),
.B(n_72),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_69),
.B(n_92),
.Y(n_91)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g119 ( 
.A(n_70),
.B(n_78),
.Y(n_119)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_72),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_74),
.B(n_77),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_74),
.B(n_92),
.Y(n_185)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_75),
.B(n_95),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_78),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_80),
.A2(n_97),
.B1(n_98),
.B2(n_109),
.Y(n_79)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_80),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_81),
.A2(n_82),
.B1(n_90),
.B2(n_96),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_82),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_87),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_85),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_86),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_88),
.B(n_89),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_90),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_93),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_94),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_94),
.B(n_119),
.Y(n_118)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_99),
.B(n_104),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_99),
.A2(n_100),
.B1(n_104),
.B2(n_105),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_100),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_102),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_102),
.B(n_136),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_105),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_111),
.B(n_114),
.C(n_116),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_111),
.A2(n_112),
.B1(n_207),
.B2(n_208),
.Y(n_206)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_114),
.A2(n_115),
.B1(n_116),
.B2(n_117),
.Y(n_207)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

CKINVDCx14_ASAP7_75t_R g116 ( 
.A(n_117),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_118),
.B(n_120),
.C(n_121),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_SL g193 ( 
.A(n_118),
.B(n_194),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_120),
.A2(n_121),
.B1(n_122),
.B2(n_195),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_120),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_122),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_123),
.B(n_137),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_124),
.B(n_126),
.Y(n_123)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_126),
.B(n_138),
.Y(n_151)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

AOI21xp5_ASAP7_75t_L g129 ( 
.A1(n_130),
.A2(n_204),
.B(n_209),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_SL g130 ( 
.A1(n_131),
.A2(n_189),
.B(n_203),
.Y(n_130)
);

AOI21xp5_ASAP7_75t_L g131 ( 
.A1(n_132),
.A2(n_170),
.B(n_188),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_SL g132 ( 
.A1(n_133),
.A2(n_158),
.B(n_169),
.Y(n_132)
);

AOI21xp5_ASAP7_75t_L g133 ( 
.A1(n_134),
.A2(n_147),
.B(n_157),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_139),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_135),
.B(n_139),
.Y(n_157)
);

INVxp33_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_140),
.A2(n_141),
.B1(n_143),
.B2(n_144),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_141),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g159 ( 
.A(n_141),
.B(n_143),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_144),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_145),
.B(n_182),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_SL g147 ( 
.A1(n_148),
.A2(n_152),
.B(n_156),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_150),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_149),
.B(n_150),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_151),
.B(n_168),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_153),
.B(n_154),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_160),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_159),
.B(n_160),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_167),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_162),
.A2(n_163),
.B1(n_164),
.B2(n_165),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_162),
.B(n_165),
.C(n_167),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_163),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_165),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_166),
.B(n_199),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_172),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_171),
.B(n_172),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_173),
.A2(n_179),
.B1(n_180),
.B2(n_187),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_173),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_174),
.A2(n_175),
.B1(n_176),
.B2(n_178),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_175),
.B(n_176),
.Y(n_200)
);

CKINVDCx16_ASAP7_75t_R g178 ( 
.A(n_176),
.Y(n_178)
);

CKINVDCx16_ASAP7_75t_R g179 ( 
.A(n_180),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_181),
.A2(n_183),
.B1(n_184),
.B2(n_186),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_181),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_183),
.B(n_186),
.C(n_187),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_184),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_191),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_190),
.B(n_191),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_192),
.A2(n_193),
.B1(n_196),
.B2(n_197),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_192),
.B(n_198),
.C(n_202),
.Y(n_205)
);

CKINVDCx16_ASAP7_75t_R g192 ( 
.A(n_193),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_197),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_198),
.A2(n_200),
.B1(n_201),
.B2(n_202),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_198),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_200),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_206),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_SL g209 ( 
.A(n_205),
.B(n_206),
.Y(n_209)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_207),
.Y(n_208)
);


endmodule