module fake_jpeg_6006_n_279 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_279);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_279;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_272;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_155;
wire n_140;
wire n_258;
wire n_96;

INVx1_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

INVx2_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_1),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_11),
.Y(n_23)
);

BUFx10_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_11),
.B(n_13),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_14),
.Y(n_28)
);

INVx11_ASAP7_75t_SL g29 ( 
.A(n_0),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_3),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_6),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_29),
.Y(n_32)
);

INVx11_ASAP7_75t_L g48 ( 
.A(n_32),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_15),
.B(n_8),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_33),
.B(n_36),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_29),
.Y(n_34)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_35),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_22),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_22),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_37),
.B(n_38),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_22),
.Y(n_38)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_39),
.Y(n_45)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_24),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_40),
.B(n_35),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_SL g41 ( 
.A(n_25),
.B(n_8),
.Y(n_41)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_42),
.Y(n_71)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_44),
.B(n_50),
.Y(n_67)
);

AND2x2_ASAP7_75t_SL g46 ( 
.A(n_39),
.B(n_24),
.Y(n_46)
);

CKINVDCx14_ASAP7_75t_R g85 ( 
.A(n_46),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_33),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_47),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_L g49 ( 
.A1(n_39),
.A2(n_16),
.B1(n_18),
.B2(n_17),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_49),
.A2(n_52),
.B1(n_63),
.B2(n_20),
.Y(n_83)
);

OR2x2_ASAP7_75t_L g50 ( 
.A(n_39),
.B(n_31),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_40),
.B(n_19),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_51),
.B(n_55),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_L g52 ( 
.A1(n_40),
.A2(n_18),
.B1(n_17),
.B2(n_28),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_34),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_41),
.A2(n_19),
.B1(n_30),
.B2(n_28),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_56),
.A2(n_23),
.B1(n_26),
.B2(n_15),
.Y(n_75)
);

AND2x2_ASAP7_75t_L g57 ( 
.A(n_34),
.B(n_24),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_57),
.B(n_62),
.Y(n_70)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_32),
.Y(n_58)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_58),
.Y(n_79)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_32),
.Y(n_59)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_59),
.Y(n_86)
);

BUFx5_ASAP7_75t_L g61 ( 
.A(n_32),
.Y(n_61)
);

INVx1_ASAP7_75t_SL g87 ( 
.A(n_61),
.Y(n_87)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_32),
.Y(n_62)
);

OAI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_37),
.A2(n_31),
.B1(n_30),
.B2(n_23),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_34),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_64),
.B(n_26),
.Y(n_76)
);

INVx13_ASAP7_75t_L g66 ( 
.A(n_64),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_66),
.B(n_73),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_61),
.Y(n_68)
);

INVx3_ASAP7_75t_SL g99 ( 
.A(n_68),
.Y(n_99)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_46),
.Y(n_72)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_72),
.Y(n_92)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_50),
.Y(n_73)
);

CKINVDCx16_ASAP7_75t_R g74 ( 
.A(n_57),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_74),
.A2(n_75),
.B1(n_47),
.B2(n_21),
.Y(n_89)
);

CKINVDCx16_ASAP7_75t_R g107 ( 
.A(n_76),
.Y(n_107)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_50),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_77),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_48),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_78),
.Y(n_97)
);

INVx4_ASAP7_75t_SL g80 ( 
.A(n_46),
.Y(n_80)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_80),
.Y(n_96)
);

OA22x2_ASAP7_75t_L g82 ( 
.A1(n_46),
.A2(n_57),
.B1(n_49),
.B2(n_36),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_82),
.A2(n_60),
.B1(n_45),
.B2(n_65),
.Y(n_101)
);

OAI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_83),
.A2(n_54),
.B1(n_20),
.B2(n_21),
.Y(n_98)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_44),
.Y(n_84)
);

CKINVDCx14_ASAP7_75t_R g91 ( 
.A(n_84),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_71),
.B(n_42),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_88),
.B(n_98),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_89),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_82),
.A2(n_60),
.B1(n_51),
.B2(n_59),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_93),
.A2(n_101),
.B1(n_103),
.B2(n_108),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_85),
.B(n_55),
.C(n_57),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_94),
.B(n_81),
.C(n_72),
.Y(n_118)
);

AOI32xp33_ASAP7_75t_L g95 ( 
.A1(n_80),
.A2(n_53),
.A3(n_65),
.B1(n_60),
.B2(n_45),
.Y(n_95)
);

XOR2xp5_ASAP7_75t_L g112 ( 
.A(n_95),
.B(n_110),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_71),
.B(n_54),
.Y(n_100)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_100),
.Y(n_113)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_67),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_102),
.B(n_66),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_82),
.A2(n_62),
.B1(n_58),
.B2(n_48),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_80),
.Y(n_104)
);

INVx13_ASAP7_75t_L g133 ( 
.A(n_104),
.Y(n_133)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_82),
.B(n_53),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_SL g130 ( 
.A1(n_105),
.A2(n_86),
.B(n_79),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_69),
.B(n_34),
.Y(n_106)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_106),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_74),
.A2(n_48),
.B1(n_43),
.B2(n_37),
.Y(n_108)
);

XNOR2xp5_ASAP7_75t_L g110 ( 
.A(n_70),
.B(n_25),
.Y(n_110)
);

INVx11_ASAP7_75t_L g111 ( 
.A(n_99),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_111),
.B(n_116),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_105),
.A2(n_73),
.B1(n_77),
.B2(n_75),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_118),
.B(n_124),
.C(n_94),
.Y(n_138)
);

CKINVDCx16_ASAP7_75t_R g119 ( 
.A(n_109),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_119),
.B(n_120),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_105),
.A2(n_81),
.B1(n_83),
.B2(n_45),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_88),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_121),
.B(n_127),
.Y(n_135)
);

OA22x2_ASAP7_75t_L g122 ( 
.A1(n_103),
.A2(n_36),
.B1(n_38),
.B2(n_37),
.Y(n_122)
);

AO22x1_ASAP7_75t_SL g153 ( 
.A1(n_122),
.A2(n_99),
.B1(n_78),
.B2(n_36),
.Y(n_153)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_123),
.Y(n_141)
);

XOR2xp5_ASAP7_75t_L g124 ( 
.A(n_110),
.B(n_41),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_90),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_125),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_90),
.A2(n_43),
.B1(n_84),
.B2(n_86),
.Y(n_126)
);

INVxp67_ASAP7_75t_L g158 ( 
.A(n_126),
.Y(n_158)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_100),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_107),
.B(n_79),
.Y(n_129)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_129),
.Y(n_157)
);

AOI21xp5_ASAP7_75t_L g149 ( 
.A1(n_130),
.A2(n_96),
.B(n_92),
.Y(n_149)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_109),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_131),
.B(n_132),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_107),
.B(n_68),
.Y(n_132)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_108),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_134),
.B(n_93),
.Y(n_139)
);

AND2x6_ASAP7_75t_L g137 ( 
.A(n_112),
.B(n_96),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_137),
.B(n_151),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_138),
.B(n_147),
.C(n_155),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_SL g160 ( 
.A1(n_139),
.A2(n_145),
.B(n_149),
.Y(n_160)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_111),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_142),
.B(n_152),
.Y(n_183)
);

CKINVDCx10_ASAP7_75t_R g143 ( 
.A(n_122),
.Y(n_143)
);

INVx1_ASAP7_75t_SL g163 ( 
.A(n_143),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_125),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_SL g176 ( 
.A(n_144),
.B(n_141),
.Y(n_176)
);

AND2x2_ASAP7_75t_L g145 ( 
.A(n_116),
.B(n_95),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_121),
.B(n_106),
.Y(n_146)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_146),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g147 ( 
.A(n_112),
.B(n_101),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_SL g150 ( 
.A1(n_130),
.A2(n_92),
.B(n_102),
.Y(n_150)
);

AOI21xp5_ASAP7_75t_L g166 ( 
.A1(n_150),
.A2(n_119),
.B(n_114),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_SL g151 ( 
.A(n_120),
.B(n_24),
.Y(n_151)
);

CKINVDCx16_ASAP7_75t_R g152 ( 
.A(n_123),
.Y(n_152)
);

OA21x2_ASAP7_75t_L g173 ( 
.A1(n_153),
.A2(n_122),
.B(n_126),
.Y(n_173)
);

XOR2xp5_ASAP7_75t_L g155 ( 
.A(n_118),
.B(n_99),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_115),
.B(n_91),
.Y(n_156)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_156),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_117),
.B(n_24),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_159),
.B(n_131),
.C(n_113),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_136),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_161),
.B(n_165),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_139),
.A2(n_134),
.B1(n_122),
.B2(n_117),
.Y(n_164)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_164),
.Y(n_186)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_156),
.Y(n_165)
);

AOI21xp5_ASAP7_75t_L g192 ( 
.A1(n_166),
.A2(n_167),
.B(n_160),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_SL g167 ( 
.A1(n_149),
.A2(n_115),
.B(n_127),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_154),
.A2(n_145),
.B1(n_140),
.B2(n_158),
.Y(n_168)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_168),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_169),
.B(n_174),
.C(n_180),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_157),
.B(n_129),
.Y(n_171)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_171),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_148),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_172),
.B(n_175),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_173),
.B(n_178),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_155),
.B(n_124),
.C(n_113),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_135),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_176),
.Y(n_202)
);

INVxp67_ASAP7_75t_L g178 ( 
.A(n_150),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_146),
.B(n_128),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_179),
.B(n_34),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_147),
.B(n_128),
.C(n_122),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_137),
.A2(n_43),
.B1(n_133),
.B2(n_97),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_182),
.A2(n_158),
.B1(n_153),
.B2(n_142),
.Y(n_197)
);

INVxp67_ASAP7_75t_L g188 ( 
.A(n_183),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_188),
.B(n_196),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_162),
.B(n_174),
.C(n_138),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_189),
.B(n_191),
.C(n_193),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_162),
.B(n_151),
.C(n_145),
.Y(n_191)
);

NOR3xp33_ASAP7_75t_L g218 ( 
.A(n_192),
.B(n_194),
.C(n_0),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_SL g193 ( 
.A(n_168),
.B(n_159),
.Y(n_193)
);

XOR2x2_ASAP7_75t_SL g194 ( 
.A(n_160),
.B(n_143),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_181),
.B(n_133),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_195),
.B(n_36),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_SL g196 ( 
.A(n_169),
.B(n_133),
.Y(n_196)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_197),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_180),
.B(n_153),
.C(n_34),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_199),
.B(n_167),
.C(n_166),
.Y(n_211)
);

INVxp67_ASAP7_75t_L g200 ( 
.A(n_182),
.Y(n_200)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_200),
.Y(n_213)
);

INVxp33_ASAP7_75t_SL g201 ( 
.A(n_163),
.Y(n_201)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_201),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_204),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_184),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_SL g235 ( 
.A1(n_205),
.A2(n_219),
.B(n_222),
.Y(n_235)
);

A2O1A1Ixp33_ASAP7_75t_SL g207 ( 
.A1(n_194),
.A2(n_173),
.B(n_178),
.C(n_163),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g229 ( 
.A1(n_207),
.A2(n_197),
.B1(n_188),
.B2(n_193),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_200),
.A2(n_177),
.B1(n_170),
.B2(n_173),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_208),
.A2(n_209),
.B1(n_198),
.B2(n_187),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_186),
.A2(n_177),
.B1(n_170),
.B2(n_164),
.Y(n_209)
);

XNOR2x1_ASAP7_75t_L g210 ( 
.A(n_195),
.B(n_181),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_SL g225 ( 
.A(n_210),
.B(n_218),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_211),
.B(n_68),
.C(n_27),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_SL g215 ( 
.A(n_202),
.B(n_87),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_215),
.B(n_216),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_SL g216 ( 
.A(n_203),
.B(n_87),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_217),
.B(n_192),
.Y(n_227)
);

AND2x2_ASAP7_75t_L g219 ( 
.A(n_199),
.B(n_22),
.Y(n_219)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_190),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_211),
.B(n_185),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_223),
.B(n_227),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_206),
.B(n_189),
.C(n_185),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_SL g238 ( 
.A1(n_224),
.A2(n_231),
.B(n_232),
.Y(n_238)
);

AOI21xp5_ASAP7_75t_L g239 ( 
.A1(n_226),
.A2(n_207),
.B(n_221),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_210),
.B(n_191),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_228),
.B(n_207),
.Y(n_245)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_229),
.Y(n_244)
);

INVx5_ASAP7_75t_L g230 ( 
.A(n_214),
.Y(n_230)
);

INVxp67_ASAP7_75t_SL g247 ( 
.A(n_230),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_218),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_206),
.B(n_78),
.C(n_38),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_SL g249 ( 
.A1(n_233),
.A2(n_237),
.B(n_0),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_213),
.A2(n_27),
.B1(n_38),
.B2(n_0),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_234),
.A2(n_8),
.B1(n_13),
.B2(n_2),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_212),
.B(n_38),
.C(n_27),
.Y(n_237)
);

AOI21xp5_ASAP7_75t_L g253 ( 
.A1(n_239),
.A2(n_240),
.B(n_246),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_SL g240 ( 
.A(n_236),
.B(n_219),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_237),
.B(n_220),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_SL g257 ( 
.A(n_241),
.B(n_242),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_235),
.B(n_27),
.Y(n_242)
);

MAJx2_ASAP7_75t_L g250 ( 
.A(n_245),
.B(n_227),
.C(n_225),
.Y(n_250)
);

OAI21xp5_ASAP7_75t_L g246 ( 
.A1(n_230),
.A2(n_207),
.B(n_1),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_248),
.A2(n_9),
.B1(n_2),
.B2(n_4),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_249),
.B(n_238),
.Y(n_254)
);

MAJx2_ASAP7_75t_L g265 ( 
.A(n_250),
.B(n_255),
.C(n_9),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_247),
.B(n_246),
.Y(n_251)
);

AOI21xp5_ASAP7_75t_L g264 ( 
.A1(n_251),
.A2(n_252),
.B(n_254),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_248),
.B(n_233),
.Y(n_252)
);

NOR2x1_ASAP7_75t_R g255 ( 
.A(n_245),
.B(n_225),
.Y(n_255)
);

BUFx24_ASAP7_75t_SL g256 ( 
.A(n_243),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_256),
.B(n_259),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_244),
.B(n_224),
.Y(n_258)
);

AOI21xp5_ASAP7_75t_L g266 ( 
.A1(n_258),
.A2(n_10),
.B(n_4),
.Y(n_266)
);

OAI21xp5_ASAP7_75t_SL g261 ( 
.A1(n_253),
.A2(n_239),
.B(n_243),
.Y(n_261)
);

AOI21xp5_ASAP7_75t_L g270 ( 
.A1(n_261),
.A2(n_262),
.B(n_263),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_257),
.B(n_228),
.Y(n_262)
);

OAI21xp5_ASAP7_75t_SL g263 ( 
.A1(n_251),
.A2(n_9),
.B(n_4),
.Y(n_263)
);

OAI21x1_ASAP7_75t_SL g269 ( 
.A1(n_265),
.A2(n_6),
.B(n_7),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_SL g268 ( 
.A1(n_266),
.A2(n_11),
.B(n_5),
.Y(n_268)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_264),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_267),
.B(n_268),
.Y(n_272)
);

OAI21xp5_ASAP7_75t_SL g274 ( 
.A1(n_269),
.A2(n_12),
.B(n_13),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_260),
.B(n_6),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_271),
.B(n_7),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_273),
.B(n_274),
.C(n_270),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_275),
.B(n_276),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_272),
.B(n_12),
.C(n_14),
.Y(n_276)
);

AND2x4_ASAP7_75t_L g278 ( 
.A(n_277),
.B(n_1),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_278),
.B(n_1),
.Y(n_279)
);


endmodule