module fake_jpeg_20272_n_178 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_178);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_178;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_93;
wire n_54;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_21),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_7),
.Y(n_52)
);

INVx11_ASAP7_75t_SL g53 ( 
.A(n_35),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_14),
.Y(n_54)
);

CKINVDCx14_ASAP7_75t_R g55 ( 
.A(n_46),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_42),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_4),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_8),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_10),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_26),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_20),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_25),
.Y(n_62)
);

BUFx12_ASAP7_75t_L g63 ( 
.A(n_34),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_33),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_15),
.Y(n_65)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_30),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_11),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_9),
.Y(n_68)
);

INVx5_ASAP7_75t_L g69 ( 
.A(n_48),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_50),
.Y(n_70)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_37),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_4),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_47),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_41),
.Y(n_74)
);

BUFx10_ASAP7_75t_L g75 ( 
.A(n_7),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_28),
.Y(n_76)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_39),
.Y(n_77)
);

INVx6_ASAP7_75t_L g78 ( 
.A(n_29),
.Y(n_78)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_68),
.Y(n_79)
);

INVx6_ASAP7_75t_L g88 ( 
.A(n_79),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_61),
.Y(n_80)
);

INVx6_ASAP7_75t_L g87 ( 
.A(n_80),
.Y(n_87)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_68),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_81),
.B(n_83),
.Y(n_98)
);

BUFx3_ASAP7_75t_L g82 ( 
.A(n_59),
.Y(n_82)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_82),
.Y(n_90)
);

INVx11_ASAP7_75t_L g83 ( 
.A(n_53),
.Y(n_83)
);

BUFx2_ASAP7_75t_L g84 ( 
.A(n_59),
.Y(n_84)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_84),
.Y(n_96)
);

INVx11_ASAP7_75t_L g85 ( 
.A(n_53),
.Y(n_85)
);

CKINVDCx16_ASAP7_75t_R g97 ( 
.A(n_85),
.Y(n_97)
);

AOI21xp33_ASAP7_75t_L g86 ( 
.A1(n_55),
.A2(n_0),
.B(n_1),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_86),
.B(n_75),
.Y(n_99)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_84),
.Y(n_89)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_89),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_79),
.A2(n_78),
.B1(n_77),
.B2(n_69),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_91),
.A2(n_94),
.B1(n_63),
.B2(n_52),
.Y(n_106)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_84),
.Y(n_92)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_92),
.Y(n_102)
);

FAx1_ASAP7_75t_L g93 ( 
.A(n_81),
.B(n_63),
.CI(n_55),
.CON(n_93),
.SN(n_93)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_93),
.B(n_75),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_80),
.A2(n_66),
.B1(n_71),
.B2(n_62),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_82),
.B(n_57),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_95),
.B(n_99),
.Y(n_105)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_83),
.Y(n_100)
);

INVx2_ASAP7_75t_SL g116 ( 
.A(n_100),
.Y(n_116)
);

INVx3_ASAP7_75t_SL g103 ( 
.A(n_90),
.Y(n_103)
);

CKINVDCx16_ASAP7_75t_R g119 ( 
.A(n_103),
.Y(n_119)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_98),
.Y(n_104)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_104),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_106),
.B(n_108),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_87),
.A2(n_85),
.B1(n_51),
.B2(n_64),
.Y(n_107)
);

OAI21xp33_ASAP7_75t_L g125 ( 
.A1(n_107),
.A2(n_0),
.B(n_2),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_99),
.A2(n_65),
.B1(n_74),
.B2(n_56),
.Y(n_108)
);

OAI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_88),
.A2(n_76),
.B1(n_61),
.B2(n_70),
.Y(n_109)
);

OAI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_109),
.A2(n_87),
.B1(n_76),
.B2(n_67),
.Y(n_117)
);

AND2x2_ASAP7_75t_L g127 ( 
.A(n_110),
.B(n_2),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_93),
.B(n_72),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_111),
.B(n_112),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_98),
.B(n_58),
.Y(n_112)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_97),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_113),
.B(n_115),
.Y(n_129)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_96),
.Y(n_114)
);

INVx4_ASAP7_75t_L g118 ( 
.A(n_114),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_91),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_117),
.A2(n_129),
.B1(n_120),
.B2(n_107),
.Y(n_135)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_114),
.Y(n_121)
);

INVx1_ASAP7_75t_SL g142 ( 
.A(n_121),
.Y(n_142)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_116),
.Y(n_122)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_122),
.Y(n_130)
);

FAx1_ASAP7_75t_SL g123 ( 
.A(n_105),
.B(n_60),
.CI(n_73),
.CON(n_123),
.SN(n_123)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_123),
.B(n_124),
.Y(n_138)
);

FAx1_ASAP7_75t_SL g124 ( 
.A(n_109),
.B(n_54),
.CI(n_1),
.CON(n_124),
.SN(n_124)
);

AOI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_125),
.A2(n_119),
.B1(n_116),
.B2(n_124),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_SL g139 ( 
.A1(n_127),
.A2(n_3),
.B(n_5),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_128),
.B(n_101),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_131),
.B(n_132),
.Y(n_144)
);

AND2x2_ASAP7_75t_L g132 ( 
.A(n_127),
.B(n_102),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_123),
.B(n_103),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_133),
.B(n_137),
.Y(n_154)
);

CKINVDCx14_ASAP7_75t_R g147 ( 
.A(n_134),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_135),
.A2(n_141),
.B1(n_6),
.B2(n_8),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_126),
.B(n_23),
.C(n_45),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_136),
.B(n_19),
.C(n_40),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_117),
.B(n_22),
.Y(n_137)
);

CKINVDCx14_ASAP7_75t_R g150 ( 
.A(n_139),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_SL g140 ( 
.A1(n_125),
.A2(n_3),
.B(n_5),
.Y(n_140)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_140),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_118),
.A2(n_24),
.B1(n_44),
.B2(n_43),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_143),
.B(n_148),
.Y(n_155)
);

INVx4_ASAP7_75t_L g146 ( 
.A(n_142),
.Y(n_146)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_146),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_130),
.Y(n_148)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_141),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_149),
.B(n_151),
.Y(n_158)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_137),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_152),
.A2(n_153),
.B1(n_13),
.B2(n_16),
.Y(n_156)
);

OAI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_138),
.A2(n_6),
.B1(n_9),
.B2(n_12),
.Y(n_153)
);

INVxp33_ASAP7_75t_SL g162 ( 
.A(n_156),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_154),
.A2(n_17),
.B1(n_18),
.B2(n_27),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_159),
.B(n_160),
.C(n_152),
.Y(n_164)
);

INVxp67_ASAP7_75t_L g160 ( 
.A(n_144),
.Y(n_160)
);

XOR2xp5_ASAP7_75t_L g161 ( 
.A(n_147),
.B(n_31),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_SL g163 ( 
.A(n_161),
.B(n_143),
.Y(n_163)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_163),
.Y(n_166)
);

INVx1_ASAP7_75t_SL g165 ( 
.A(n_164),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_165),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_167),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_168),
.B(n_160),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_169),
.B(n_157),
.C(n_155),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_170),
.B(n_146),
.Y(n_171)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_171),
.Y(n_172)
);

OR2x2_ASAP7_75t_L g173 ( 
.A(n_172),
.B(n_162),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_173),
.A2(n_158),
.B1(n_153),
.B2(n_166),
.Y(n_174)
);

INVxp67_ASAP7_75t_L g175 ( 
.A(n_174),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_175),
.A2(n_145),
.B1(n_150),
.B2(n_38),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_176),
.B(n_32),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_177),
.B(n_36),
.C(n_49),
.Y(n_178)
);


endmodule