module fake_jpeg_27378_n_218 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_218);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_218;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_121;
wire n_130;
wire n_99;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_145;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_140;
wire n_82;
wire n_128;
wire n_100;
wire n_96;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_5),
.Y(n_17)
);

BUFx8_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_16),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_11),
.Y(n_21)
);

BUFx4f_ASAP7_75t_SL g22 ( 
.A(n_2),
.Y(n_22)
);

CKINVDCx16_ASAP7_75t_R g23 ( 
.A(n_16),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_2),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_10),
.Y(n_27)
);

BUFx10_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

INVx11_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

BUFx12_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_10),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_30),
.Y(n_35)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_35),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_30),
.Y(n_36)
);

INVx3_ASAP7_75t_SL g62 ( 
.A(n_36),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_17),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_37),
.B(n_39),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g38 ( 
.A(n_17),
.B(n_0),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_38),
.B(n_45),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_25),
.Y(n_39)
);

OR2x2_ASAP7_75t_L g40 ( 
.A(n_31),
.B(n_0),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_40),
.B(n_19),
.Y(n_55)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_30),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_42),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

INVx4_ASAP7_75t_SL g54 ( 
.A(n_43),
.Y(n_54)
);

INVx2_ASAP7_75t_SL g44 ( 
.A(n_22),
.Y(n_44)
);

INVx11_ASAP7_75t_L g59 ( 
.A(n_44),
.Y(n_59)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_22),
.Y(n_45)
);

HB1xp67_ASAP7_75t_L g46 ( 
.A(n_42),
.Y(n_46)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_46),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g47 ( 
.A(n_45),
.B(n_40),
.C(n_22),
.Y(n_47)
);

XNOR2xp5_ASAP7_75t_L g97 ( 
.A(n_47),
.B(n_28),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_37),
.B(n_21),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_48),
.B(n_66),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_44),
.A2(n_29),
.B1(n_25),
.B2(n_27),
.Y(n_49)
);

AOI21xp5_ASAP7_75t_L g74 ( 
.A1(n_49),
.A2(n_63),
.B(n_67),
.Y(n_74)
);

OR2x2_ASAP7_75t_L g92 ( 
.A(n_55),
.B(n_24),
.Y(n_92)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_42),
.Y(n_56)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_56),
.Y(n_91)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_58),
.Y(n_96)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_36),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_60),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_61),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_44),
.A2(n_29),
.B1(n_33),
.B2(n_27),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_40),
.B(n_28),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_64),
.B(n_22),
.Y(n_78)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_36),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_65),
.B(n_36),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_39),
.B(n_33),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_44),
.A2(n_29),
.B1(n_21),
.B2(n_34),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_38),
.A2(n_34),
.B1(n_26),
.B2(n_23),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_68),
.A2(n_34),
.B1(n_23),
.B2(n_45),
.Y(n_82)
);

INVx5_ASAP7_75t_L g69 ( 
.A(n_52),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_69),
.B(n_72),
.Y(n_107)
);

INVx13_ASAP7_75t_L g70 ( 
.A(n_52),
.Y(n_70)
);

INVx4_ASAP7_75t_L g112 ( 
.A(n_70),
.Y(n_112)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_71),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_51),
.B(n_26),
.Y(n_72)
);

INVx13_ASAP7_75t_L g73 ( 
.A(n_52),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_73),
.B(n_79),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_57),
.B(n_40),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g105 ( 
.A(n_76),
.B(n_78),
.Y(n_105)
);

INVx13_ASAP7_75t_L g79 ( 
.A(n_52),
.Y(n_79)
);

AND2x6_ASAP7_75t_L g80 ( 
.A(n_47),
.B(n_7),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_SL g102 ( 
.A(n_80),
.B(n_82),
.C(n_18),
.Y(n_102)
);

NAND3xp33_ASAP7_75t_L g81 ( 
.A(n_57),
.B(n_8),
.C(n_15),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_81),
.B(n_88),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_68),
.B(n_31),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_83),
.B(n_84),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_61),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_64),
.B(n_31),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_85),
.B(n_87),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_50),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_54),
.B(n_19),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_50),
.B(n_22),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_89),
.B(n_98),
.Y(n_103)
);

INVx13_ASAP7_75t_L g90 ( 
.A(n_54),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_90),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_92),
.B(n_19),
.Y(n_106)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_53),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_93),
.B(n_94),
.Y(n_100)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_53),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_97),
.B(n_43),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_60),
.B(n_28),
.Y(n_98)
);

HB1xp67_ASAP7_75t_L g101 ( 
.A(n_98),
.Y(n_101)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_101),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_102),
.A2(n_106),
.B1(n_111),
.B2(n_109),
.Y(n_130)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_89),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_104),
.B(n_106),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_92),
.B(n_6),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_109),
.B(n_111),
.Y(n_124)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_82),
.Y(n_111)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_75),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_113),
.B(n_114),
.Y(n_144)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_75),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_86),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_115),
.B(n_118),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_117),
.B(n_74),
.C(n_80),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_95),
.B(n_7),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_78),
.B(n_32),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_120),
.B(n_90),
.Y(n_126)
);

AND2x2_ASAP7_75t_L g122 ( 
.A(n_97),
.B(n_43),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g131 ( 
.A(n_122),
.B(n_117),
.Y(n_131)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_112),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_123),
.B(n_137),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_126),
.B(n_136),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_SL g150 ( 
.A(n_127),
.B(n_108),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_117),
.B(n_74),
.C(n_77),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_128),
.B(n_140),
.C(n_142),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_130),
.A2(n_133),
.B1(n_135),
.B2(n_138),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_L g160 ( 
.A1(n_131),
.A2(n_140),
.B(n_142),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_122),
.A2(n_94),
.B1(n_93),
.B2(n_77),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_121),
.B(n_69),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g154 ( 
.A(n_134),
.B(n_112),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_103),
.A2(n_65),
.B1(n_62),
.B2(n_96),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_100),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_100),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_122),
.A2(n_62),
.B1(n_96),
.B2(n_91),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_103),
.B(n_91),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_139),
.B(n_110),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_104),
.B(n_56),
.C(n_58),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_102),
.A2(n_62),
.B1(n_35),
.B2(n_41),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_141),
.A2(n_143),
.B1(n_73),
.B2(n_70),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_105),
.B(n_86),
.C(n_79),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_105),
.A2(n_116),
.B1(n_99),
.B2(n_114),
.Y(n_143)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_107),
.Y(n_145)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_145),
.Y(n_147)
);

CKINVDCx16_ASAP7_75t_R g148 ( 
.A(n_144),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_148),
.B(n_152),
.Y(n_173)
);

XOR2xp5_ASAP7_75t_L g149 ( 
.A(n_128),
.B(n_131),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_SL g171 ( 
.A(n_149),
.B(n_165),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_SL g176 ( 
.A(n_150),
.B(n_160),
.Y(n_176)
);

OAI32xp33_ASAP7_75t_L g151 ( 
.A1(n_129),
.A2(n_99),
.A3(n_119),
.B1(n_115),
.B2(n_113),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_151),
.A2(n_164),
.B1(n_123),
.B2(n_35),
.Y(n_169)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_139),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_153),
.B(n_154),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_138),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_156),
.B(n_158),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_131),
.B(n_110),
.Y(n_158)
);

AO21x1_ASAP7_75t_L g159 ( 
.A1(n_132),
.A2(n_118),
.B(n_18),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_159),
.B(n_161),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_127),
.B(n_59),
.C(n_32),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_163),
.B(n_32),
.C(n_28),
.Y(n_170)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_135),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_143),
.B(n_28),
.Y(n_165)
);

NAND3xp33_ASAP7_75t_L g166 ( 
.A(n_165),
.B(n_124),
.C(n_133),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_166),
.B(n_167),
.Y(n_183)
);

AOI211xp5_ASAP7_75t_L g167 ( 
.A1(n_151),
.A2(n_141),
.B(n_125),
.C(n_28),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_169),
.A2(n_175),
.B1(n_162),
.B2(n_157),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_170),
.B(n_174),
.C(n_178),
.Y(n_191)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_146),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_172),
.B(n_180),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_150),
.B(n_24),
.C(n_20),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_156),
.A2(n_18),
.B1(n_24),
.B2(n_20),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_155),
.B(n_20),
.C(n_59),
.Y(n_178)
);

BUFx24_ASAP7_75t_SL g180 ( 
.A(n_147),
.Y(n_180)
);

NAND3xp33_ASAP7_75t_L g181 ( 
.A(n_158),
.B(n_1),
.C(n_2),
.Y(n_181)
);

AOI21xp5_ASAP7_75t_L g186 ( 
.A1(n_181),
.A2(n_159),
.B(n_3),
.Y(n_186)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_173),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_182),
.B(n_185),
.Y(n_195)
);

A2O1A1Ixp33_ASAP7_75t_SL g184 ( 
.A1(n_179),
.A2(n_155),
.B(n_163),
.C(n_161),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_L g203 ( 
.A1(n_184),
.A2(n_186),
.B(n_4),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_168),
.A2(n_157),
.B1(n_160),
.B2(n_149),
.Y(n_185)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_188),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_166),
.A2(n_153),
.B1(n_18),
.B2(n_11),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_189),
.B(n_190),
.Y(n_198)
);

HB1xp67_ASAP7_75t_L g190 ( 
.A(n_177),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_172),
.A2(n_18),
.B1(n_3),
.B2(n_4),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_SL g194 ( 
.A(n_192),
.B(n_1),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_176),
.B(n_9),
.C(n_12),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_193),
.B(n_171),
.C(n_181),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_194),
.B(n_197),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_SL g206 ( 
.A(n_196),
.B(n_200),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_SL g197 ( 
.A(n_187),
.B(n_13),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_SL g200 ( 
.A(n_193),
.B(n_1),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_185),
.B(n_171),
.Y(n_201)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_201),
.Y(n_207)
);

OAI21x1_ASAP7_75t_L g202 ( 
.A1(n_183),
.A2(n_3),
.B(n_4),
.Y(n_202)
);

OAI31xp33_ASAP7_75t_L g209 ( 
.A1(n_202),
.A2(n_203),
.A3(n_184),
.B(n_198),
.Y(n_209)
);

OAI31xp33_ASAP7_75t_L g204 ( 
.A1(n_195),
.A2(n_189),
.A3(n_184),
.B(n_191),
.Y(n_204)
);

CKINVDCx16_ASAP7_75t_R g211 ( 
.A(n_204),
.Y(n_211)
);

A2O1A1Ixp33_ASAP7_75t_L g205 ( 
.A1(n_199),
.A2(n_184),
.B(n_191),
.C(n_5),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_205),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_209),
.B(n_205),
.C(n_206),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_207),
.B(n_204),
.Y(n_212)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_213),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_212),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_L g217 ( 
.A1(n_215),
.A2(n_216),
.B(n_214),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_SL g216 ( 
.A1(n_211),
.A2(n_208),
.B(n_210),
.Y(n_216)
);

BUFx24_ASAP7_75t_SL g218 ( 
.A(n_217),
.Y(n_218)
);


endmodule