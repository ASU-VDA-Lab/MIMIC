module fake_jpeg_11393_n_198 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_198);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_198;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_76;
wire n_127;
wire n_154;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g51 ( 
.A(n_46),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_24),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_42),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_49),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_16),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_22),
.Y(n_57)
);

BUFx5_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_32),
.Y(n_59)
);

INVx11_ASAP7_75t_SL g60 ( 
.A(n_30),
.Y(n_60)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_48),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_43),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_8),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_17),
.Y(n_64)
);

BUFx12f_ASAP7_75t_L g65 ( 
.A(n_35),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_38),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_14),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_0),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_27),
.Y(n_69)
);

BUFx5_ASAP7_75t_L g70 ( 
.A(n_28),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_25),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_1),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_50),
.Y(n_73)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_14),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_5),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_29),
.Y(n_76)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_44),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_21),
.Y(n_78)
);

CKINVDCx16_ASAP7_75t_R g79 ( 
.A(n_3),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_45),
.Y(n_80)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_41),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_56),
.Y(n_82)
);

INVx6_ASAP7_75t_L g96 ( 
.A(n_82),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_56),
.Y(n_83)
);

INVx6_ASAP7_75t_L g97 ( 
.A(n_83),
.Y(n_97)
);

BUFx3_ASAP7_75t_L g84 ( 
.A(n_54),
.Y(n_84)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_84),
.Y(n_94)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_74),
.Y(n_85)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_85),
.Y(n_98)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_63),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_86),
.B(n_87),
.Y(n_100)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_75),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_69),
.Y(n_88)
);

BUFx2_ASAP7_75t_L g104 ( 
.A(n_88),
.Y(n_104)
);

AND2x4_ASAP7_75t_L g89 ( 
.A(n_61),
.B(n_19),
.Y(n_89)
);

CKINVDCx16_ASAP7_75t_R g102 ( 
.A(n_89),
.Y(n_102)
);

INVx6_ASAP7_75t_SL g90 ( 
.A(n_60),
.Y(n_90)
);

BUFx2_ASAP7_75t_R g92 ( 
.A(n_90),
.Y(n_92)
);

INVx6_ASAP7_75t_L g91 ( 
.A(n_72),
.Y(n_91)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_91),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_82),
.A2(n_72),
.B1(n_65),
.B2(n_54),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_93),
.A2(n_65),
.B1(n_54),
.B2(n_77),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_89),
.B(n_68),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_95),
.B(n_99),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_89),
.B(n_67),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_83),
.B(n_52),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_101),
.B(n_65),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_88),
.A2(n_69),
.B1(n_71),
.B2(n_78),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_103),
.A2(n_60),
.B1(n_73),
.B2(n_81),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_L g106 ( 
.A1(n_91),
.A2(n_71),
.B1(n_78),
.B2(n_73),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_106),
.A2(n_59),
.B1(n_55),
.B2(n_53),
.Y(n_125)
);

NAND2xp33_ASAP7_75t_SL g107 ( 
.A(n_102),
.B(n_79),
.Y(n_107)
);

CKINVDCx16_ASAP7_75t_R g138 ( 
.A(n_107),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_108),
.B(n_111),
.Y(n_133)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_94),
.Y(n_109)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_109),
.Y(n_143)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_110),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_100),
.B(n_62),
.Y(n_111)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_105),
.Y(n_112)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_112),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_L g113 ( 
.A(n_98),
.B(n_51),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_113),
.B(n_115),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_114),
.A2(n_123),
.B1(n_129),
.B2(n_126),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_92),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_93),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_116),
.B(n_117),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_94),
.B(n_80),
.C(n_76),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_104),
.Y(n_118)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_118),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_92),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_119),
.B(n_124),
.Y(n_151)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_104),
.Y(n_120)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_120),
.Y(n_141)
);

INVx2_ASAP7_75t_SL g121 ( 
.A(n_96),
.Y(n_121)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_121),
.Y(n_146)
);

AND2x2_ASAP7_75t_L g122 ( 
.A(n_96),
.B(n_97),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_122),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_106),
.A2(n_64),
.B1(n_66),
.B2(n_57),
.Y(n_123)
);

CKINVDCx16_ASAP7_75t_R g124 ( 
.A(n_97),
.Y(n_124)
);

OA21x2_ASAP7_75t_L g139 ( 
.A1(n_125),
.A2(n_3),
.B(n_4),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_103),
.A2(n_70),
.B1(n_58),
.B2(n_2),
.Y(n_126)
);

OAI22xp33_ASAP7_75t_L g130 ( 
.A1(n_126),
.A2(n_110),
.B1(n_116),
.B2(n_107),
.Y(n_130)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_100),
.Y(n_127)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_127),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_103),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_130),
.A2(n_142),
.B1(n_6),
.B2(n_7),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_131),
.B(n_139),
.Y(n_162)
);

INVx5_ASAP7_75t_L g135 ( 
.A(n_109),
.Y(n_135)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_135),
.Y(n_155)
);

BUFx24_ASAP7_75t_SL g136 ( 
.A(n_128),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_136),
.B(n_149),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_121),
.Y(n_137)
);

BUFx5_ASAP7_75t_L g165 ( 
.A(n_137),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_122),
.Y(n_140)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_140),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_116),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_111),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_111),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_152),
.B(n_12),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_153),
.A2(n_145),
.B1(n_140),
.B2(n_143),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_L g154 ( 
.A1(n_134),
.A2(n_7),
.B(n_8),
.Y(n_154)
);

NOR3xp33_ASAP7_75t_L g179 ( 
.A(n_154),
.B(n_157),
.C(n_169),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_134),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_156),
.A2(n_161),
.B1(n_137),
.B2(n_141),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_L g157 ( 
.A1(n_150),
.A2(n_151),
.B(n_145),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_144),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_158),
.B(n_159),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_148),
.B(n_33),
.C(n_47),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_138),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_163),
.B(n_164),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_147),
.B(n_12),
.Y(n_164)
);

INVxp67_ASAP7_75t_L g166 ( 
.A(n_146),
.Y(n_166)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_166),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_133),
.B(n_13),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_167),
.B(n_139),
.Y(n_177)
);

A2O1A1Ixp33_ASAP7_75t_SL g169 ( 
.A1(n_130),
.A2(n_36),
.B(n_15),
.C(n_18),
.Y(n_169)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_155),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_170),
.B(n_176),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_166),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_173),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_174),
.A2(n_169),
.B1(n_153),
.B2(n_165),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_160),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_177),
.B(n_178),
.Y(n_182)
);

AO22x1_ASAP7_75t_SL g180 ( 
.A1(n_168),
.A2(n_132),
.B1(n_13),
.B2(n_23),
.Y(n_180)
);

AO22x1_ASAP7_75t_SL g185 ( 
.A1(n_180),
.A2(n_169),
.B1(n_165),
.B2(n_31),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_SL g183 ( 
.A(n_180),
.B(n_162),
.Y(n_183)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_183),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_184),
.Y(n_188)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_185),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_SL g190 ( 
.A1(n_189),
.A2(n_186),
.B(n_181),
.Y(n_190)
);

AOI21x1_ASAP7_75t_L g191 ( 
.A1(n_190),
.A2(n_181),
.B(n_188),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_191),
.B(n_180),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_192),
.B(n_182),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_193),
.A2(n_187),
.B1(n_172),
.B2(n_179),
.Y(n_194)
);

AO21x1_ASAP7_75t_L g195 ( 
.A1(n_194),
.A2(n_179),
.B(n_169),
.Y(n_195)
);

O2A1O1Ixp33_ASAP7_75t_SL g196 ( 
.A1(n_195),
.A2(n_175),
.B(n_26),
.C(n_34),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_L g197 ( 
.A1(n_196),
.A2(n_171),
.B(n_37),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_197),
.B(n_20),
.Y(n_198)
);


endmodule