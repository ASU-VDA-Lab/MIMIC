module real_jpeg_15688_n_8 (n_5, n_4, n_0, n_1, n_2, n_6, n_7, n_3, n_8);

input n_5;
input n_4;
input n_0;
input n_1;
input n_2;
input n_6;
input n_7;
input n_3;

output n_8;

wire n_17;
wire n_21;
wire n_10;
wire n_9;
wire n_12;
wire n_24;
wire n_23;
wire n_11;
wire n_14;
wire n_25;
wire n_22;
wire n_18;
wire n_26;
wire n_20;
wire n_19;
wire n_16;
wire n_15;
wire n_13;

OAI21xp5_ASAP7_75t_SL g16 ( 
.A1(n_0),
.A2(n_1),
.B(n_17),
.Y(n_16)
);

CKINVDCx6p67_ASAP7_75t_R g24 ( 
.A(n_0),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_1),
.Y(n_12)
);

NOR2xp33_ASAP7_75t_R g23 ( 
.A(n_1),
.B(n_24),
.Y(n_23)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_2),
.Y(n_11)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_3),
.B(n_11),
.Y(n_26)
);

INVx2_ASAP7_75t_R g19 ( 
.A(n_4),
.Y(n_19)
);

INVx2_ASAP7_75t_R g15 ( 
.A(n_5),
.Y(n_15)
);

NAND3xp33_ASAP7_75t_SL g22 ( 
.A(n_5),
.B(n_17),
.C(n_23),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g10 ( 
.A(n_6),
.B(n_11),
.Y(n_10)
);

NAND2xp5_ASAP7_75t_SL g25 ( 
.A(n_6),
.B(n_26),
.Y(n_25)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

OAI22xp5_ASAP7_75t_L g8 ( 
.A1(n_9),
.A2(n_21),
.B1(n_22),
.B2(n_25),
.Y(n_8)
);

AOI21xp5_ASAP7_75t_L g9 ( 
.A1(n_10),
.A2(n_12),
.B(n_13),
.Y(n_9)
);

AOI21xp5_ASAP7_75t_L g14 ( 
.A1(n_12),
.A2(n_15),
.B(n_16),
.Y(n_14)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_14),
.Y(n_13)
);

INVx2_ASAP7_75t_SL g17 ( 
.A(n_18),
.Y(n_17)
);

OR2x4_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_20),
.Y(n_18)
);


endmodule