module fake_jpeg_9641_n_312 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_312);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_312;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

INVx8_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_2),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_11),
.Y(n_23)
);

BUFx8_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_11),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_32),
.B(n_0),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_SL g47 ( 
.A(n_34),
.B(n_42),
.Y(n_47)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_30),
.Y(n_35)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_35),
.Y(n_60)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_33),
.Y(n_36)
);

HB1xp67_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

INVx5_ASAP7_75t_L g37 ( 
.A(n_24),
.Y(n_37)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

AND2x2_ASAP7_75t_L g38 ( 
.A(n_33),
.B(n_0),
.Y(n_38)
);

NAND2xp33_ASAP7_75t_SL g64 ( 
.A(n_38),
.B(n_19),
.Y(n_64)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_33),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_39),
.B(n_43),
.Y(n_49)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_20),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_30),
.Y(n_41)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_23),
.B(n_15),
.Y(n_42)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_20),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_23),
.B(n_15),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_SL g54 ( 
.A(n_44),
.B(n_16),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_37),
.Y(n_45)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_45),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_34),
.B(n_32),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_50),
.B(n_53),
.Y(n_92)
);

INVx6_ASAP7_75t_SL g52 ( 
.A(n_37),
.Y(n_52)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_52),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_34),
.B(n_16),
.Y(n_53)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_54),
.Y(n_80)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_42),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_55),
.B(n_56),
.Y(n_94)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_44),
.Y(n_56)
);

OR2x2_ASAP7_75t_L g57 ( 
.A(n_35),
.B(n_28),
.Y(n_57)
);

NAND2xp33_ASAP7_75t_SL g70 ( 
.A(n_57),
.B(n_64),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_40),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_58),
.Y(n_71)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_38),
.Y(n_61)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_61),
.Y(n_88)
);

INVx13_ASAP7_75t_L g62 ( 
.A(n_37),
.Y(n_62)
);

INVx5_ASAP7_75t_L g81 ( 
.A(n_62),
.Y(n_81)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_43),
.Y(n_63)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_63),
.Y(n_91)
);

INVx1_ASAP7_75t_SL g65 ( 
.A(n_35),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_65),
.A2(n_40),
.B1(n_43),
.B2(n_39),
.Y(n_68)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_38),
.Y(n_66)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_66),
.Y(n_95)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_43),
.Y(n_67)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_67),
.Y(n_73)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_68),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_55),
.A2(n_19),
.B1(n_56),
.B2(n_40),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_69),
.A2(n_85),
.B1(n_90),
.B2(n_76),
.Y(n_113)
);

O2A1O1Ixp33_ASAP7_75t_SL g72 ( 
.A1(n_64),
.A2(n_38),
.B(n_41),
.C(n_35),
.Y(n_72)
);

OAI21xp5_ASAP7_75t_SL g112 ( 
.A1(n_72),
.A2(n_83),
.B(n_54),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_L g74 ( 
.A1(n_61),
.A2(n_19),
.B1(n_39),
.B2(n_36),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_74),
.A2(n_48),
.B1(n_60),
.B2(n_51),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_66),
.A2(n_38),
.B1(n_28),
.B2(n_21),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_75),
.A2(n_79),
.B1(n_84),
.B2(n_86),
.Y(n_105)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_46),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_76),
.B(n_82),
.Y(n_103)
);

OA22x2_ASAP7_75t_L g77 ( 
.A1(n_58),
.A2(n_41),
.B1(n_36),
.B2(n_20),
.Y(n_77)
);

A2O1A1Ixp33_ASAP7_75t_SL g111 ( 
.A1(n_77),
.A2(n_51),
.B(n_45),
.C(n_24),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_50),
.A2(n_21),
.B1(n_18),
.B2(n_29),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_49),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_L g83 ( 
.A1(n_53),
.A2(n_18),
.B(n_26),
.Y(n_83)
);

OAI22xp33_ASAP7_75t_L g84 ( 
.A1(n_59),
.A2(n_52),
.B1(n_20),
.B2(n_31),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_62),
.A2(n_26),
.B1(n_29),
.B2(n_24),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_49),
.A2(n_25),
.B1(n_31),
.B2(n_22),
.Y(n_86)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_46),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_87),
.B(n_89),
.Y(n_122)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_63),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_62),
.A2(n_24),
.B1(n_12),
.B2(n_11),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_74),
.A2(n_65),
.B1(n_60),
.B2(n_59),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_96),
.A2(n_98),
.B1(n_99),
.B2(n_107),
.Y(n_125)
);

INVx8_ASAP7_75t_L g97 ( 
.A(n_81),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_97),
.B(n_104),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_88),
.A2(n_95),
.B1(n_72),
.B2(n_70),
.Y(n_98)
);

OAI22x1_ASAP7_75t_SL g99 ( 
.A1(n_72),
.A2(n_70),
.B1(n_77),
.B2(n_86),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_92),
.B(n_47),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_100),
.B(n_102),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_L g101 ( 
.A1(n_82),
.A2(n_67),
.B1(n_48),
.B2(n_59),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_101),
.A2(n_110),
.B1(n_118),
.B2(n_89),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_92),
.B(n_47),
.Y(n_102)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_81),
.Y(n_104)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_77),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_106),
.B(n_109),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_88),
.A2(n_95),
.B1(n_94),
.B2(n_71),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_108),
.A2(n_111),
.B1(n_120),
.B2(n_93),
.Y(n_135)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_81),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_75),
.A2(n_60),
.B1(n_65),
.B2(n_51),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_L g126 ( 
.A1(n_112),
.A2(n_116),
.B(n_102),
.Y(n_126)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_113),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_94),
.B(n_41),
.C(n_45),
.Y(n_114)
);

AND2x2_ASAP7_75t_L g136 ( 
.A(n_114),
.B(n_99),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_79),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_115),
.B(n_117),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_83),
.B(n_57),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_116),
.B(n_119),
.Y(n_130)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_87),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_71),
.A2(n_57),
.B1(n_27),
.B2(n_31),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_80),
.B(n_17),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_77),
.A2(n_27),
.B1(n_25),
.B2(n_22),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_80),
.B(n_13),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_123),
.B(n_15),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_126),
.B(n_137),
.Y(n_154)
);

BUFx2_ASAP7_75t_L g127 ( 
.A(n_104),
.Y(n_127)
);

CKINVDCx16_ASAP7_75t_R g166 ( 
.A(n_127),
.Y(n_166)
);

BUFx3_ASAP7_75t_L g128 ( 
.A(n_109),
.Y(n_128)
);

INVx11_ASAP7_75t_L g153 ( 
.A(n_128),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_122),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_129),
.B(n_131),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_97),
.Y(n_132)
);

CKINVDCx10_ASAP7_75t_R g157 ( 
.A(n_132),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_135),
.A2(n_138),
.B1(n_145),
.B2(n_146),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_136),
.B(n_139),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_99),
.A2(n_77),
.B1(n_73),
.B2(n_91),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_100),
.B(n_78),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_L g140 ( 
.A1(n_106),
.A2(n_78),
.B(n_91),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g160 ( 
.A(n_140),
.Y(n_160)
);

BUFx3_ASAP7_75t_L g141 ( 
.A(n_97),
.Y(n_141)
);

INVx4_ASAP7_75t_L g173 ( 
.A(n_141),
.Y(n_173)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_122),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_142),
.B(n_143),
.Y(n_165)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_117),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_98),
.A2(n_115),
.B1(n_121),
.B2(n_120),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_105),
.A2(n_73),
.B1(n_93),
.B2(n_45),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_96),
.A2(n_93),
.B1(n_45),
.B2(n_25),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_147),
.A2(n_110),
.B1(n_119),
.B2(n_103),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_108),
.B(n_27),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_148),
.B(n_101),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_127),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_150),
.B(n_151),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_127),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_133),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_152),
.B(n_155),
.Y(n_176)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_133),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_149),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_156),
.B(n_162),
.Y(n_183)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_144),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_158),
.B(n_161),
.Y(n_179)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_144),
.Y(n_161)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_128),
.Y(n_162)
);

INVx13_ASAP7_75t_L g163 ( 
.A(n_141),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_SL g199 ( 
.A1(n_163),
.A2(n_170),
.B1(n_111),
.B2(n_132),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_149),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_SL g189 ( 
.A1(n_167),
.A2(n_103),
.B(n_142),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_SL g178 ( 
.A(n_168),
.B(n_147),
.Y(n_178)
);

AND2x6_ASAP7_75t_L g169 ( 
.A(n_136),
.B(n_112),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_169),
.Y(n_186)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_140),
.Y(n_170)
);

OAI32xp33_ASAP7_75t_L g171 ( 
.A1(n_138),
.A2(n_118),
.A3(n_107),
.B1(n_105),
.B2(n_111),
.Y(n_171)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_171),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_172),
.A2(n_154),
.B1(n_158),
.B2(n_161),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_174),
.B(n_126),
.C(n_136),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_175),
.B(n_177),
.C(n_185),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_174),
.B(n_124),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_178),
.B(n_166),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_154),
.A2(n_125),
.B1(n_135),
.B2(n_145),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_180),
.A2(n_152),
.B1(n_164),
.B2(n_173),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g218 ( 
.A1(n_184),
.A2(n_192),
.B1(n_197),
.B2(n_199),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_169),
.B(n_159),
.Y(n_185)
);

INVxp67_ASAP7_75t_L g187 ( 
.A(n_157),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_187),
.B(n_188),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_165),
.Y(n_188)
);

AO21x1_ASAP7_75t_L g211 ( 
.A1(n_189),
.A2(n_190),
.B(n_163),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_SL g190 ( 
.A1(n_160),
.A2(n_134),
.B(n_125),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_170),
.B(n_114),
.C(n_124),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_191),
.B(n_196),
.C(n_155),
.Y(n_202)
);

AOI21xp5_ASAP7_75t_L g192 ( 
.A1(n_156),
.A2(n_129),
.B(n_130),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_167),
.A2(n_148),
.B1(n_146),
.B2(n_130),
.Y(n_193)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_193),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_165),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_194),
.B(n_179),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_171),
.A2(n_137),
.B1(n_139),
.B2(n_111),
.Y(n_195)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_195),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_159),
.B(n_141),
.C(n_132),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_168),
.A2(n_111),
.B1(n_143),
.B2(n_123),
.Y(n_197)
);

A2O1A1O1Ixp25_ASAP7_75t_L g198 ( 
.A1(n_164),
.A2(n_111),
.B(n_131),
.C(n_24),
.D(n_30),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_198),
.B(n_157),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_SL g200 ( 
.A(n_177),
.B(n_172),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_SL g234 ( 
.A(n_200),
.B(n_207),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_202),
.B(n_205),
.C(n_212),
.Y(n_231)
);

HB1xp67_ASAP7_75t_L g203 ( 
.A(n_187),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_203),
.B(n_216),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_204),
.A2(n_222),
.B1(n_197),
.B2(n_179),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_175),
.B(n_150),
.C(n_151),
.Y(n_205)
);

INVxp67_ASAP7_75t_L g208 ( 
.A(n_182),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_208),
.B(n_211),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_183),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_209),
.B(n_210),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_SL g210 ( 
.A(n_192),
.B(n_162),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_191),
.B(n_166),
.C(n_173),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_SL g213 ( 
.A(n_184),
.B(n_163),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_213),
.B(n_190),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_215),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_176),
.Y(n_216)
);

AND2x2_ASAP7_75t_L g217 ( 
.A(n_185),
.B(n_0),
.Y(n_217)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_217),
.Y(n_223)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_176),
.Y(n_220)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_220),
.Y(n_235)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_221),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_181),
.A2(n_153),
.B1(n_14),
.B2(n_13),
.Y(n_222)
);

AOI21x1_ASAP7_75t_L g224 ( 
.A1(n_211),
.A2(n_213),
.B(n_189),
.Y(n_224)
);

O2A1O1Ixp33_ASAP7_75t_L g246 ( 
.A1(n_224),
.A2(n_229),
.B(n_193),
.C(n_222),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_226),
.B(n_200),
.Y(n_248)
);

INVxp67_ASAP7_75t_L g228 ( 
.A(n_219),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_228),
.B(n_242),
.Y(n_245)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_204),
.Y(n_230)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_230),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_L g232 ( 
.A1(n_214),
.A2(n_181),
.B1(n_196),
.B2(n_186),
.Y(n_232)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_232),
.Y(n_249)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_218),
.Y(n_233)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_233),
.Y(n_252)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_208),
.Y(n_237)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_237),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_202),
.B(n_186),
.C(n_180),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_240),
.B(n_201),
.C(n_212),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_206),
.A2(n_194),
.B1(n_188),
.B2(n_195),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_L g253 ( 
.A1(n_241),
.A2(n_217),
.B1(n_198),
.B2(n_178),
.Y(n_253)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_205),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_231),
.B(n_201),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_243),
.B(n_248),
.Y(n_269)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_246),
.Y(n_266)
);

HB1xp67_ASAP7_75t_L g247 ( 
.A(n_224),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_247),
.B(n_251),
.Y(n_264)
);

AOI21xp5_ASAP7_75t_L g262 ( 
.A1(n_250),
.A2(n_256),
.B(n_223),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_231),
.B(n_207),
.C(n_217),
.Y(n_251)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_253),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_226),
.B(n_153),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_254),
.B(n_255),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_SL g255 ( 
.A(n_238),
.B(n_14),
.Y(n_255)
);

XNOR2x1_ASAP7_75t_L g256 ( 
.A(n_234),
.B(n_13),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_240),
.B(n_30),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_257),
.B(n_239),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_233),
.A2(n_22),
.B1(n_17),
.B2(n_30),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_259),
.A2(n_228),
.B1(n_237),
.B2(n_235),
.Y(n_263)
);

AOI21xp5_ASAP7_75t_L g260 ( 
.A1(n_252),
.A2(n_225),
.B(n_230),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_260),
.B(n_254),
.Y(n_273)
);

OAI21xp5_ASAP7_75t_L g261 ( 
.A1(n_244),
.A2(n_225),
.B(n_241),
.Y(n_261)
);

AOI21xp5_ASAP7_75t_L g274 ( 
.A1(n_261),
.A2(n_246),
.B(n_251),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_262),
.B(n_1),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_263),
.A2(n_271),
.B1(n_0),
.B2(n_1),
.Y(n_281)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_265),
.Y(n_277)
);

OAI221xp5_ASAP7_75t_L g268 ( 
.A1(n_245),
.A2(n_256),
.B1(n_223),
.B2(n_227),
.C(n_250),
.Y(n_268)
);

AND2x2_ASAP7_75t_L g275 ( 
.A(n_268),
.B(n_257),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_258),
.B(n_229),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_270),
.B(n_1),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_249),
.A2(n_236),
.B1(n_234),
.B2(n_17),
.Y(n_271)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_273),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_L g291 ( 
.A1(n_274),
.A2(n_281),
.B1(n_283),
.B2(n_2),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_275),
.B(n_279),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_269),
.B(n_243),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_276),
.B(n_278),
.C(n_280),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_269),
.B(n_248),
.C(n_1),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_SL g279 ( 
.A(n_267),
.B(n_12),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_261),
.B(n_12),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_282),
.B(n_275),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_272),
.A2(n_266),
.B1(n_271),
.B2(n_263),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_SL g286 ( 
.A(n_284),
.B(n_280),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_286),
.B(n_289),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_276),
.B(n_264),
.C(n_260),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_287),
.B(n_7),
.C(n_8),
.Y(n_298)
);

OAI21xp5_ASAP7_75t_SL g288 ( 
.A1(n_277),
.A2(n_2),
.B(n_4),
.Y(n_288)
);

AOI21xp5_ASAP7_75t_L g296 ( 
.A1(n_288),
.A2(n_291),
.B(n_294),
.Y(n_296)
);

A2O1A1Ixp33_ASAP7_75t_L g292 ( 
.A1(n_273),
.A2(n_2),
.B(n_4),
.C(n_6),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_292),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_297)
);

OAI21x1_ASAP7_75t_L g294 ( 
.A1(n_278),
.A2(n_4),
.B(n_6),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_287),
.B(n_285),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_295),
.B(n_297),
.Y(n_305)
);

OAI21xp5_ASAP7_75t_L g304 ( 
.A1(n_298),
.A2(n_9),
.B(n_10),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_285),
.B(n_7),
.Y(n_299)
);

AOI21xp5_ASAP7_75t_L g307 ( 
.A1(n_299),
.A2(n_301),
.B(n_302),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_293),
.B(n_7),
.Y(n_301)
);

OAI21xp5_ASAP7_75t_SL g302 ( 
.A1(n_290),
.A2(n_9),
.B(n_10),
.Y(n_302)
);

AOI21xp5_ASAP7_75t_SL g303 ( 
.A1(n_300),
.A2(n_292),
.B(n_9),
.Y(n_303)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_303),
.Y(n_309)
);

BUFx24_ASAP7_75t_SL g308 ( 
.A(n_304),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_298),
.A2(n_9),
.B1(n_296),
.B2(n_297),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_SL g310 ( 
.A(n_309),
.B(n_305),
.Y(n_310)
);

OAI21xp5_ASAP7_75t_L g311 ( 
.A1(n_310),
.A2(n_307),
.B(n_306),
.Y(n_311)
);

XOR2xp5_ASAP7_75t_L g312 ( 
.A(n_311),
.B(n_308),
.Y(n_312)
);


endmodule