module fake_jpeg_10314_n_233 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_233);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_233;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_187;
wire n_57;
wire n_21;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_3),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

INVxp67_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_3),
.Y(n_21)
);

BUFx12_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_5),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_2),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_10),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_4),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_28),
.Y(n_34)
);

INVx11_ASAP7_75t_L g51 ( 
.A(n_34),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_35),
.Y(n_62)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_36),
.B(n_37),
.Y(n_49)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_17),
.Y(n_37)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_38),
.B(n_39),
.Y(n_56)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_18),
.B(n_1),
.Y(n_40)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_40),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_16),
.Y(n_41)
);

INVx5_ASAP7_75t_SL g59 ( 
.A(n_41),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_16),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_25),
.Y(n_43)
);

AND2x2_ASAP7_75t_L g48 ( 
.A(n_43),
.B(n_25),
.Y(n_48)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_26),
.Y(n_44)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_44),
.Y(n_46)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_26),
.Y(n_45)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_45),
.Y(n_47)
);

HAxp5_ASAP7_75t_SL g88 ( 
.A(n_48),
.B(n_22),
.CON(n_88),
.SN(n_88)
);

AOI22xp33_ASAP7_75t_L g50 ( 
.A1(n_36),
.A2(n_19),
.B1(n_18),
.B2(n_30),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_50),
.A2(n_57),
.B1(n_61),
.B2(n_63),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_44),
.A2(n_19),
.B1(n_32),
.B2(n_27),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_52),
.A2(n_33),
.B1(n_31),
.B2(n_22),
.Y(n_78)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_45),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_53),
.B(n_55),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_40),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_54),
.B(n_60),
.Y(n_87)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_34),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_L g57 ( 
.A1(n_34),
.A2(n_21),
.B1(n_23),
.B2(n_30),
.Y(n_57)
);

INVxp67_ASAP7_75t_L g60 ( 
.A(n_42),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g61 ( 
.A1(n_38),
.A2(n_27),
.B1(n_32),
.B2(n_28),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_L g63 ( 
.A1(n_37),
.A2(n_21),
.B1(n_29),
.B2(n_24),
.Y(n_63)
);

OAI22xp33_ASAP7_75t_L g65 ( 
.A1(n_38),
.A2(n_28),
.B1(n_33),
.B2(n_29),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_65),
.A2(n_67),
.B1(n_22),
.B2(n_2),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_39),
.B(n_31),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_66),
.B(n_62),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_43),
.A2(n_24),
.B1(n_23),
.B2(n_20),
.Y(n_67)
);

INVxp67_ASAP7_75t_L g70 ( 
.A(n_49),
.Y(n_70)
);

INVx13_ASAP7_75t_L g91 ( 
.A(n_70),
.Y(n_91)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_49),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_71),
.B(n_73),
.Y(n_95)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_51),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_72),
.B(n_76),
.Y(n_98)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_56),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_56),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_74),
.B(n_75),
.Y(n_105)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_66),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_54),
.B(n_31),
.Y(n_76)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_51),
.Y(n_77)
);

INVx3_ASAP7_75t_SL g100 ( 
.A(n_77),
.Y(n_100)
);

OAI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_78),
.A2(n_82),
.B1(n_85),
.B2(n_86),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_48),
.B(n_31),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_79),
.B(n_67),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_51),
.Y(n_80)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_80),
.Y(n_106)
);

HB1xp67_ASAP7_75t_L g81 ( 
.A(n_46),
.Y(n_81)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_81),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_64),
.B(n_1),
.Y(n_83)
);

XNOR2xp5_ASAP7_75t_L g97 ( 
.A(n_83),
.B(n_5),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_61),
.A2(n_42),
.B1(n_41),
.B2(n_35),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_84),
.A2(n_59),
.B1(n_35),
.B2(n_62),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_64),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_48),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_86),
.B(n_89),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_88),
.B(n_22),
.Y(n_109)
);

XOR2xp5_ASAP7_75t_L g133 ( 
.A(n_90),
.B(n_102),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_93),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_75),
.A2(n_55),
.B1(n_53),
.B2(n_46),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_94),
.A2(n_62),
.B1(n_58),
.B2(n_8),
.Y(n_134)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_69),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_96),
.B(n_101),
.Y(n_122)
);

NOR2xp67_ASAP7_75t_R g114 ( 
.A(n_97),
.B(n_83),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_89),
.B(n_47),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_99),
.B(n_111),
.Y(n_116)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_87),
.Y(n_101)
);

XOR2xp5_ASAP7_75t_L g102 ( 
.A(n_79),
.B(n_68),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_102),
.B(n_108),
.C(n_82),
.Y(n_115)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_84),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_103),
.B(n_110),
.Y(n_127)
);

OAI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_71),
.A2(n_47),
.B1(n_59),
.B2(n_41),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_104),
.A2(n_107),
.B1(n_77),
.B2(n_72),
.Y(n_121)
);

AND2x2_ASAP7_75t_SL g108 ( 
.A(n_73),
.B(n_35),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_109),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_83),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_70),
.B(n_58),
.Y(n_111)
);

BUFx2_ASAP7_75t_SL g113 ( 
.A(n_100),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_113),
.A2(n_106),
.B1(n_91),
.B2(n_92),
.Y(n_143)
);

MAJx2_ASAP7_75t_L g145 ( 
.A(n_114),
.B(n_97),
.C(n_108),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_115),
.B(n_108),
.C(n_98),
.Y(n_142)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_99),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_117),
.B(n_120),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_112),
.B(n_74),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_118),
.B(n_119),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_112),
.B(n_68),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_95),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_121),
.A2(n_125),
.B1(n_7),
.B2(n_9),
.Y(n_153)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_95),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_123),
.B(n_126),
.Y(n_151)
);

OA21x2_ASAP7_75t_L g124 ( 
.A1(n_103),
.A2(n_80),
.B(n_59),
.Y(n_124)
);

AOI21xp5_ASAP7_75t_L g136 ( 
.A1(n_124),
.A2(n_100),
.B(n_111),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_105),
.B(n_80),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_100),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_128),
.B(n_130),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_101),
.B(n_58),
.Y(n_129)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_129),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_105),
.B(n_58),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_94),
.Y(n_131)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_131),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_133),
.B(n_92),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_134),
.A2(n_107),
.B1(n_91),
.B2(n_110),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_135),
.A2(n_143),
.B1(n_153),
.B2(n_120),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_SL g157 ( 
.A1(n_136),
.A2(n_141),
.B(n_134),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_122),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_138),
.B(n_144),
.Y(n_168)
);

AOI21xp5_ASAP7_75t_L g141 ( 
.A1(n_124),
.A2(n_109),
.B(n_90),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_142),
.B(n_133),
.C(n_115),
.Y(n_159)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_126),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_SL g161 ( 
.A(n_145),
.B(n_147),
.Y(n_161)
);

AOI32xp33_ASAP7_75t_L g146 ( 
.A1(n_127),
.A2(n_108),
.A3(n_91),
.B1(n_96),
.B2(n_106),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_L g169 ( 
.A1(n_146),
.A2(n_150),
.B(n_129),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_131),
.A2(n_15),
.B1(n_14),
.B2(n_8),
.Y(n_148)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_148),
.Y(n_163)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_113),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_149),
.B(n_154),
.Y(n_162)
);

AOI21xp5_ASAP7_75t_SL g150 ( 
.A1(n_127),
.A2(n_6),
.B(n_7),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_122),
.Y(n_154)
);

A2O1A1Ixp33_ASAP7_75t_L g156 ( 
.A1(n_141),
.A2(n_119),
.B(n_118),
.C(n_132),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_156),
.B(n_165),
.Y(n_188)
);

AOI22xp33_ASAP7_75t_L g187 ( 
.A1(n_157),
.A2(n_160),
.B1(n_169),
.B2(n_174),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_139),
.B(n_144),
.Y(n_158)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_158),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g175 ( 
.A(n_159),
.B(n_142),
.Y(n_175)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_149),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_164),
.B(n_155),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_140),
.Y(n_165)
);

MAJx2_ASAP7_75t_L g166 ( 
.A(n_145),
.B(n_114),
.C(n_116),
.Y(n_166)
);

XNOR2x1_ASAP7_75t_L g182 ( 
.A(n_166),
.B(n_124),
.Y(n_182)
);

NAND3xp33_ASAP7_75t_L g167 ( 
.A(n_135),
.B(n_130),
.C(n_123),
.Y(n_167)
);

NOR3xp33_ASAP7_75t_SL g190 ( 
.A(n_167),
.B(n_15),
.C(n_11),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_139),
.B(n_116),
.Y(n_170)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_170),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_137),
.B(n_128),
.Y(n_171)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_171),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_147),
.B(n_117),
.C(n_121),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_172),
.B(n_152),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_148),
.B(n_124),
.Y(n_173)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_173),
.Y(n_185)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_151),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_175),
.B(n_176),
.C(n_178),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_161),
.B(n_136),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g180 ( 
.A(n_161),
.B(n_150),
.Y(n_180)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_180),
.B(n_166),
.Y(n_197)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_181),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_SL g192 ( 
.A(n_182),
.B(n_169),
.Y(n_192)
);

CKINVDCx14_ASAP7_75t_R g184 ( 
.A(n_162),
.Y(n_184)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_184),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_168),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_SL g199 ( 
.A(n_186),
.B(n_163),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_159),
.B(n_153),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_189),
.B(n_172),
.C(n_174),
.Y(n_195)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_190),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_185),
.A2(n_163),
.B1(n_157),
.B2(n_165),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_191),
.A2(n_190),
.B1(n_189),
.B2(n_178),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_192),
.B(n_195),
.Y(n_208)
);

BUFx12_ASAP7_75t_L g196 ( 
.A(n_182),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_196),
.B(n_199),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_197),
.B(n_194),
.C(n_195),
.Y(n_207)
);

AOI21xp5_ASAP7_75t_L g198 ( 
.A1(n_188),
.A2(n_156),
.B(n_183),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_198),
.B(n_180),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_L g201 ( 
.A1(n_187),
.A2(n_158),
.B(n_170),
.Y(n_201)
);

AOI21xp5_ASAP7_75t_L g209 ( 
.A1(n_201),
.A2(n_164),
.B(n_175),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_192),
.A2(n_177),
.B1(n_179),
.B2(n_176),
.Y(n_203)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_203),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_204),
.B(n_206),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_207),
.B(n_194),
.C(n_197),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_209),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_SL g210 ( 
.A(n_200),
.B(n_9),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_210),
.B(n_211),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_193),
.B(n_9),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_212),
.B(n_11),
.C(n_12),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_204),
.A2(n_196),
.B1(n_201),
.B2(n_191),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_L g219 ( 
.A1(n_214),
.A2(n_203),
.B(n_207),
.Y(n_219)
);

AOI21xp5_ASAP7_75t_L g216 ( 
.A1(n_205),
.A2(n_196),
.B(n_202),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_SL g220 ( 
.A1(n_216),
.A2(n_206),
.B(n_208),
.Y(n_220)
);

MAJx2_ASAP7_75t_L g226 ( 
.A(n_219),
.B(n_223),
.C(n_213),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_220),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_215),
.A2(n_208),
.B1(n_12),
.B2(n_13),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_221),
.B(n_222),
.Y(n_224)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_218),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_SL g225 ( 
.A(n_223),
.B(n_217),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_225),
.Y(n_229)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_226),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_229),
.B(n_224),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_230),
.B(n_228),
.C(n_227),
.Y(n_231)
);

O2A1O1Ixp33_ASAP7_75t_SL g232 ( 
.A1(n_231),
.A2(n_212),
.B(n_214),
.C(n_13),
.Y(n_232)
);

AND2x2_ASAP7_75t_L g233 ( 
.A(n_232),
.B(n_13),
.Y(n_233)
);


endmodule