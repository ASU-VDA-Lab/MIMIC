module fake_jpeg_23726_n_44 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_44);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_44;

wire n_13;
wire n_21;
wire n_33;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_31;
wire n_25;
wire n_29;
wire n_37;
wire n_43;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

CKINVDCx20_ASAP7_75t_R g7 ( 
.A(n_6),
.Y(n_7)
);

NAND2xp5_ASAP7_75t_L g8 ( 
.A(n_3),
.B(n_2),
.Y(n_8)
);

INVx2_ASAP7_75t_L g9 ( 
.A(n_6),
.Y(n_9)
);

BUFx3_ASAP7_75t_L g10 ( 
.A(n_4),
.Y(n_10)
);

BUFx3_ASAP7_75t_L g11 ( 
.A(n_0),
.Y(n_11)
);

NOR2xp33_ASAP7_75t_L g12 ( 
.A(n_1),
.B(n_4),
.Y(n_12)
);

INVx2_ASAP7_75t_L g13 ( 
.A(n_2),
.Y(n_13)
);

OAI22xp5_ASAP7_75t_L g14 ( 
.A1(n_9),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_14)
);

OAI22xp5_ASAP7_75t_SL g22 ( 
.A1(n_14),
.A2(n_16),
.B1(n_12),
.B2(n_13),
.Y(n_22)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_10),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_SL g27 ( 
.A(n_15),
.B(n_19),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_SL g16 ( 
.A1(n_9),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_16)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_17),
.B(n_21),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_8),
.B(n_7),
.Y(n_18)
);

AND2x2_ASAP7_75t_L g23 ( 
.A(n_18),
.B(n_7),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_8),
.B(n_3),
.Y(n_19)
);

AOI22xp33_ASAP7_75t_SL g20 ( 
.A1(n_13),
.A2(n_0),
.B1(n_4),
.B2(n_5),
.Y(n_20)
);

OAI22xp5_ASAP7_75t_L g24 ( 
.A1(n_20),
.A2(n_10),
.B1(n_11),
.B2(n_5),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_12),
.B(n_5),
.Y(n_21)
);

OAI21xp5_ASAP7_75t_SL g29 ( 
.A1(n_22),
.A2(n_24),
.B(n_16),
.Y(n_29)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_23),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_21),
.B(n_6),
.Y(n_26)
);

INVx1_ASAP7_75t_SL g28 ( 
.A(n_26),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_L g37 ( 
.A1(n_29),
.A2(n_30),
.B1(n_20),
.B2(n_31),
.Y(n_37)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_24),
.Y(n_30)
);

MAJIxp5_ASAP7_75t_L g31 ( 
.A(n_27),
.B(n_15),
.C(n_14),
.Y(n_31)
);

MAJIxp5_ASAP7_75t_L g34 ( 
.A(n_31),
.B(n_27),
.C(n_19),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_L g33 ( 
.A1(n_30),
.A2(n_22),
.B1(n_20),
.B2(n_25),
.Y(n_33)
);

AOI21xp5_ASAP7_75t_L g40 ( 
.A1(n_33),
.A2(n_34),
.B(n_35),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_L g35 ( 
.A1(n_29),
.A2(n_17),
.B1(n_18),
.B2(n_23),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_L g36 ( 
.A1(n_31),
.A2(n_11),
.B1(n_23),
.B2(n_32),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_37),
.B(n_28),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g41 ( 
.A(n_38),
.B(n_39),
.Y(n_41)
);

INVx1_ASAP7_75t_SL g39 ( 
.A(n_36),
.Y(n_39)
);

MAJIxp5_ASAP7_75t_L g42 ( 
.A(n_40),
.B(n_34),
.C(n_39),
.Y(n_42)
);

INVxp67_ASAP7_75t_L g43 ( 
.A(n_42),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_SL g44 ( 
.A(n_43),
.B(n_41),
.Y(n_44)
);


endmodule