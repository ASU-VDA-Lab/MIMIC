module fake_jpeg_6334_n_162 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_162);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_162;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_127;
wire n_76;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_57;
wire n_21;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

NAND2xp5_ASAP7_75t_SL g13 ( 
.A(n_9),
.B(n_3),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_7),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_9),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_5),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_12),
.B(n_3),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_10),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_1),
.Y(n_21)
);

BUFx16f_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_5),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_6),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_4),
.Y(n_26)
);

HB1xp67_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_10),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_22),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_30),
.B(n_31),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_22),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_22),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_32),
.B(n_36),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_17),
.B(n_0),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_33),
.B(n_15),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g34 ( 
.A(n_17),
.B(n_0),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_34),
.B(n_35),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g35 ( 
.A(n_25),
.B(n_1),
.Y(n_35)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_18),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_37),
.B(n_40),
.Y(n_47)
);

BUFx2_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

NAND2x1_ASAP7_75t_SL g39 ( 
.A(n_25),
.B(n_2),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_39),
.A2(n_15),
.B1(n_28),
.B2(n_24),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_20),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_20),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_41),
.B(n_42),
.Y(n_54)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_20),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_16),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_43),
.Y(n_48)
);

INVx11_ASAP7_75t_L g44 ( 
.A(n_29),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_44),
.B(n_28),
.Y(n_56)
);

BUFx5_ASAP7_75t_L g49 ( 
.A(n_31),
.Y(n_49)
);

BUFx5_ASAP7_75t_L g82 ( 
.A(n_49),
.Y(n_82)
);

AO22x1_ASAP7_75t_SL g50 ( 
.A1(n_39),
.A2(n_29),
.B1(n_27),
.B2(n_13),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_50),
.A2(n_52),
.B1(n_57),
.B2(n_61),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_43),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_51),
.Y(n_89)
);

BUFx8_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

INVxp67_ASAP7_75t_L g75 ( 
.A(n_53),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_56),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_36),
.A2(n_37),
.B1(n_42),
.B2(n_41),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_58),
.B(n_69),
.Y(n_93)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_35),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_60),
.B(n_62),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_L g61 ( 
.A1(n_36),
.A2(n_14),
.B1(n_24),
.B2(n_19),
.Y(n_61)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_38),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_33),
.B(n_14),
.Y(n_63)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_63),
.Y(n_79)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_38),
.Y(n_64)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_64),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_L g65 ( 
.A1(n_44),
.A2(n_19),
.B1(n_23),
.B2(n_21),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_65),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_31),
.B(n_26),
.Y(n_66)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_66),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_34),
.B(n_26),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_67),
.B(n_72),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_32),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_68),
.Y(n_92)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_32),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_30),
.B(n_23),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_70),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g71 ( 
.A(n_30),
.Y(n_71)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_71),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_40),
.B(n_21),
.Y(n_72)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_40),
.Y(n_73)
);

BUFx2_ASAP7_75t_L g90 ( 
.A(n_73),
.Y(n_90)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_38),
.Y(n_74)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_74),
.Y(n_77)
);

A2O1A1Ixp33_ASAP7_75t_L g78 ( 
.A1(n_50),
.A2(n_16),
.B(n_8),
.C(n_11),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_78),
.B(n_86),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_84),
.A2(n_91),
.B1(n_95),
.B2(n_62),
.Y(n_105)
);

NOR2x1_ASAP7_75t_L g86 ( 
.A(n_50),
.B(n_53),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_67),
.A2(n_2),
.B1(n_4),
.B2(n_8),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_59),
.B(n_12),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_94),
.B(n_48),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_59),
.A2(n_48),
.B1(n_51),
.B2(n_60),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_SL g97 ( 
.A1(n_86),
.A2(n_53),
.B(n_72),
.Y(n_97)
);

AOI21xp5_ASAP7_75t_L g115 ( 
.A1(n_97),
.A2(n_75),
.B(n_92),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_98),
.B(n_99),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_87),
.B(n_68),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_87),
.B(n_69),
.Y(n_100)
);

XNOR2xp5_ASAP7_75t_L g120 ( 
.A(n_100),
.B(n_109),
.Y(n_120)
);

XOR2xp5_ASAP7_75t_L g101 ( 
.A(n_81),
.B(n_45),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_101),
.B(n_102),
.C(n_107),
.Y(n_122)
);

XOR2xp5_ASAP7_75t_L g102 ( 
.A(n_94),
.B(n_54),
.Y(n_102)
);

BUFx2_ASAP7_75t_L g103 ( 
.A(n_90),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_103),
.B(n_104),
.Y(n_117)
);

INVx13_ASAP7_75t_L g104 ( 
.A(n_82),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_105),
.B(n_108),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_83),
.B(n_46),
.C(n_47),
.Y(n_107)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_90),
.Y(n_108)
);

XNOR2xp5_ASAP7_75t_L g109 ( 
.A(n_75),
.B(n_49),
.Y(n_109)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_78),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_110),
.B(n_111),
.Y(n_121)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_93),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_89),
.B(n_55),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_112),
.B(n_114),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_89),
.B(n_71),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_113),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_92),
.B(n_74),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_L g139 ( 
.A1(n_115),
.A2(n_96),
.B(n_85),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_97),
.A2(n_55),
.B1(n_64),
.B2(n_73),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_116),
.A2(n_100),
.B1(n_107),
.B2(n_77),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_103),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_119),
.B(n_80),
.Y(n_130)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_108),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_123),
.B(n_126),
.Y(n_132)
);

BUFx12_ASAP7_75t_L g126 ( 
.A(n_104),
.Y(n_126)
);

CKINVDCx5p33_ASAP7_75t_R g127 ( 
.A(n_106),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_127),
.B(n_98),
.Y(n_133)
);

A2O1A1O1Ixp25_ASAP7_75t_L g129 ( 
.A1(n_118),
.A2(n_101),
.B(n_109),
.C(n_99),
.D(n_102),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_SL g142 ( 
.A1(n_129),
.A2(n_135),
.B(n_139),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_130),
.B(n_136),
.Y(n_145)
);

XOR2xp5_ASAP7_75t_L g131 ( 
.A(n_122),
.B(n_120),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_131),
.B(n_137),
.C(n_88),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_133),
.B(n_138),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_134),
.A2(n_120),
.B1(n_127),
.B2(n_88),
.Y(n_143)
);

AOI21xp5_ASAP7_75t_SL g135 ( 
.A1(n_115),
.A2(n_125),
.B(n_128),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_124),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_122),
.B(n_105),
.C(n_80),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_125),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_139),
.A2(n_116),
.B1(n_128),
.B2(n_121),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_140),
.A2(n_144),
.B1(n_96),
.B2(n_132),
.Y(n_149)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_143),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_135),
.A2(n_77),
.B1(n_117),
.B2(n_123),
.Y(n_144)
);

AND2x2_ASAP7_75t_L g150 ( 
.A(n_146),
.B(n_131),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_SL g147 ( 
.A(n_129),
.B(n_79),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_147),
.B(n_137),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_148),
.B(n_153),
.Y(n_154)
);

AOI322xp5_ASAP7_75t_L g157 ( 
.A1(n_149),
.A2(n_150),
.A3(n_146),
.B1(n_142),
.B2(n_140),
.C1(n_76),
.C2(n_79),
.Y(n_157)
);

OR2x2_ASAP7_75t_L g152 ( 
.A(n_141),
.B(n_82),
.Y(n_152)
);

OR2x2_ASAP7_75t_L g156 ( 
.A(n_152),
.B(n_145),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_144),
.B(n_126),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_152),
.B(n_126),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_155),
.B(n_76),
.Y(n_158)
);

AOI21xp5_ASAP7_75t_L g159 ( 
.A1(n_156),
.A2(n_157),
.B(n_151),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_158),
.B(n_159),
.C(n_151),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_160),
.B(n_154),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_161),
.B(n_150),
.Y(n_162)
);


endmodule