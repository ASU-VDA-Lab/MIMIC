module fake_jpeg_20604_n_253 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_253);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_253;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_11;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_12;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_140;
wire n_82;
wire n_128;
wire n_100;
wire n_96;

CKINVDCx16_ASAP7_75t_R g11 ( 
.A(n_6),
.Y(n_11)
);

BUFx5_ASAP7_75t_L g12 ( 
.A(n_4),
.Y(n_12)
);

BUFx6f_ASAP7_75t_SL g13 ( 
.A(n_3),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_5),
.Y(n_14)
);

INVx8_ASAP7_75t_L g15 ( 
.A(n_1),
.Y(n_15)
);

BUFx5_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

INVx11_ASAP7_75t_SL g17 ( 
.A(n_8),
.Y(n_17)
);

BUFx12_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

BUFx4f_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_2),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_19),
.Y(n_24)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_24),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_13),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_SL g42 ( 
.A(n_25),
.B(n_33),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_23),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_26),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_27),
.Y(n_35)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_19),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_28),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_19),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_19),
.Y(n_30)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_30),
.Y(n_39)
);

INVx5_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

AND2x2_ASAP7_75t_L g40 ( 
.A(n_31),
.B(n_32),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_11),
.B(n_5),
.Y(n_33)
);

AOI22xp33_ASAP7_75t_L g41 ( 
.A1(n_28),
.A2(n_21),
.B1(n_15),
.B2(n_17),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_41),
.A2(n_24),
.B1(n_11),
.B2(n_21),
.Y(n_49)
);

INVxp67_ASAP7_75t_L g43 ( 
.A(n_42),
.Y(n_43)
);

INVx13_ASAP7_75t_L g77 ( 
.A(n_43),
.Y(n_77)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_36),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_44),
.Y(n_78)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_45),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_42),
.B(n_33),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g62 ( 
.A(n_46),
.B(n_54),
.Y(n_62)
);

OAI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_39),
.A2(n_30),
.B1(n_24),
.B2(n_25),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_47),
.A2(n_49),
.B1(n_34),
.B2(n_35),
.Y(n_67)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_48),
.B(n_53),
.Y(n_71)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_50),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_37),
.A2(n_31),
.B1(n_22),
.B2(n_15),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_51),
.A2(n_59),
.B1(n_40),
.B2(n_37),
.Y(n_61)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_52),
.Y(n_74)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_42),
.B(n_22),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_41),
.B(n_18),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_55),
.B(n_57),
.Y(n_73)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_56),
.Y(n_68)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_39),
.A2(n_31),
.B1(n_13),
.B2(n_18),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_58),
.A2(n_40),
.B1(n_35),
.B2(n_34),
.Y(n_66)
);

OAI21xp33_ASAP7_75t_L g59 ( 
.A1(n_39),
.A2(n_10),
.B(n_9),
.Y(n_59)
);

INVxp67_ASAP7_75t_L g82 ( 
.A(n_61),
.Y(n_82)
);

XNOR2xp5_ASAP7_75t_L g63 ( 
.A(n_46),
.B(n_40),
.Y(n_63)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_63),
.B(n_65),
.C(n_48),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_55),
.A2(n_40),
.B1(n_26),
.B2(n_27),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_64),
.A2(n_66),
.B1(n_70),
.B2(n_75),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_54),
.B(n_40),
.C(n_32),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_67),
.B(n_38),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_49),
.A2(n_26),
.B1(n_32),
.B2(n_27),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_69),
.A2(n_67),
.B1(n_76),
.B2(n_61),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_L g70 ( 
.A1(n_47),
.A2(n_44),
.B1(n_53),
.B2(n_45),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_58),
.A2(n_32),
.B1(n_27),
.B2(n_34),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_50),
.B(n_34),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_76),
.B(n_35),
.Y(n_80)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_80),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_63),
.B(n_65),
.Y(n_81)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_81),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g83 ( 
.A(n_71),
.Y(n_83)
);

CKINVDCx16_ASAP7_75t_R g117 ( 
.A(n_83),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_62),
.B(n_35),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_84),
.B(n_85),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_62),
.B(n_48),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_86),
.A2(n_92),
.B1(n_74),
.B2(n_78),
.Y(n_110)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_78),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_87),
.B(n_88),
.Y(n_109)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_68),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_71),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_89),
.B(n_93),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_74),
.A2(n_52),
.B1(n_56),
.B2(n_57),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_90),
.A2(n_94),
.B1(n_72),
.B2(n_74),
.Y(n_105)
);

XNOR2xp5_ASAP7_75t_L g97 ( 
.A(n_91),
.B(n_95),
.Y(n_97)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_60),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_66),
.A2(n_52),
.B1(n_29),
.B2(n_2),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_73),
.B(n_29),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_90),
.Y(n_96)
);

CKINVDCx16_ASAP7_75t_R g129 ( 
.A(n_96),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_91),
.B(n_64),
.C(n_73),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_98),
.B(n_78),
.C(n_23),
.Y(n_133)
);

AOI21xp33_ASAP7_75t_SL g99 ( 
.A1(n_82),
.A2(n_77),
.B(n_75),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_SL g118 ( 
.A(n_99),
.B(n_79),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_L g102 ( 
.A1(n_85),
.A2(n_69),
.B1(n_72),
.B2(n_60),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_102),
.B(n_103),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_93),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_84),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_104),
.B(n_108),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_105),
.A2(n_79),
.B1(n_87),
.B2(n_68),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_L g106 ( 
.A1(n_89),
.A2(n_77),
.B(n_18),
.Y(n_106)
);

AOI21xp5_ASAP7_75t_L g120 ( 
.A1(n_106),
.A2(n_114),
.B(n_115),
.Y(n_120)
);

MAJx2_ASAP7_75t_L g107 ( 
.A(n_81),
.B(n_77),
.C(n_18),
.Y(n_107)
);

XNOR2xp5_ASAP7_75t_L g119 ( 
.A(n_107),
.B(n_92),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_95),
.Y(n_108)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_110),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_94),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_111),
.B(n_23),
.Y(n_142)
);

NAND2x1p5_ASAP7_75t_L g113 ( 
.A(n_86),
.B(n_68),
.Y(n_113)
);

NAND2x1p5_ASAP7_75t_L g131 ( 
.A(n_113),
.B(n_87),
.Y(n_131)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_94),
.B(n_91),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_L g115 ( 
.A1(n_92),
.A2(n_86),
.B(n_80),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_118),
.B(n_16),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_SL g151 ( 
.A(n_119),
.B(n_114),
.Y(n_151)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_109),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_122),
.B(n_124),
.Y(n_150)
);

AOI211xp5_ASAP7_75t_SL g123 ( 
.A1(n_113),
.A2(n_92),
.B(n_79),
.C(n_88),
.Y(n_123)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_123),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_116),
.Y(n_124)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_109),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_125),
.B(n_132),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_126),
.A2(n_117),
.B1(n_112),
.B2(n_107),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g127 ( 
.A(n_97),
.B(n_20),
.Y(n_127)
);

XOR2xp5_ASAP7_75t_L g158 ( 
.A(n_127),
.B(n_140),
.Y(n_158)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_116),
.Y(n_128)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_128),
.Y(n_156)
);

AND2x2_ASAP7_75t_L g167 ( 
.A(n_131),
.B(n_130),
.Y(n_167)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_100),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_133),
.B(n_112),
.C(n_14),
.Y(n_159)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_100),
.Y(n_134)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_134),
.Y(n_163)
);

AND2x2_ASAP7_75t_SL g135 ( 
.A(n_101),
.B(n_20),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_135),
.B(n_138),
.Y(n_148)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_101),
.Y(n_136)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_136),
.Y(n_164)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_115),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_103),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_139),
.B(n_144),
.Y(n_146)
);

XOR2xp5_ASAP7_75t_L g140 ( 
.A(n_97),
.B(n_20),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g141 ( 
.A(n_107),
.B(n_16),
.Y(n_141)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_141),
.B(n_145),
.Y(n_160)
);

CKINVDCx14_ASAP7_75t_R g147 ( 
.A(n_142),
.Y(n_147)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_110),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_143),
.B(n_113),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_106),
.Y(n_144)
);

XOR2xp5_ASAP7_75t_L g145 ( 
.A(n_98),
.B(n_16),
.Y(n_145)
);

XOR2xp5_ASAP7_75t_L g180 ( 
.A(n_151),
.B(n_162),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_128),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_152),
.B(n_135),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_153),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_137),
.B(n_117),
.Y(n_154)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_154),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_121),
.A2(n_105),
.B1(n_114),
.B2(n_99),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_155),
.A2(n_168),
.B1(n_126),
.B2(n_131),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_157),
.A2(n_123),
.B1(n_6),
.B2(n_2),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_159),
.B(n_133),
.C(n_140),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_L g162 ( 
.A1(n_120),
.A2(n_138),
.B(n_131),
.Y(n_162)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_165),
.B(n_166),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_SL g166 ( 
.A(n_145),
.B(n_12),
.Y(n_166)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_167),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_121),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_169),
.A2(n_167),
.B1(n_157),
.B2(n_153),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_SL g170 ( 
.A(n_161),
.B(n_127),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_170),
.B(n_165),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_155),
.A2(n_143),
.B1(n_120),
.B2(n_129),
.Y(n_171)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_171),
.Y(n_191)
);

XNOR2x1_ASAP7_75t_L g172 ( 
.A(n_151),
.B(n_118),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_172),
.A2(n_5),
.B1(n_9),
.B2(n_3),
.Y(n_201)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_173),
.Y(n_194)
);

AND2x2_ASAP7_75t_L g175 ( 
.A(n_146),
.B(n_119),
.Y(n_175)
);

AOI21xp5_ASAP7_75t_L g195 ( 
.A1(n_175),
.A2(n_162),
.B(n_148),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_177),
.B(n_178),
.C(n_184),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_159),
.B(n_141),
.C(n_135),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_179),
.A2(n_147),
.B1(n_168),
.B2(n_148),
.Y(n_197)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_150),
.Y(n_182)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_182),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_158),
.B(n_12),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_183),
.B(n_160),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_158),
.B(n_12),
.C(n_1),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_154),
.Y(n_185)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_185),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_187),
.B(n_195),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_179),
.A2(n_163),
.B1(n_149),
.B2(n_156),
.Y(n_188)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_188),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_189),
.B(n_169),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_177),
.B(n_160),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_190),
.B(n_200),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_192),
.B(n_186),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_197),
.B(n_174),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_178),
.B(n_166),
.C(n_167),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_199),
.B(n_186),
.C(n_184),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_180),
.B(n_164),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_201),
.B(n_180),
.Y(n_207)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_194),
.Y(n_203)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_203),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_198),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_204),
.B(n_206),
.Y(n_223)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_207),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_193),
.B(n_190),
.C(n_199),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_208),
.B(n_0),
.C(n_1),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_209),
.A2(n_212),
.B1(n_189),
.B2(n_191),
.Y(n_214)
);

AOI21xp5_ASAP7_75t_L g216 ( 
.A1(n_210),
.A2(n_187),
.B(n_183),
.Y(n_216)
);

INVx11_ASAP7_75t_L g213 ( 
.A(n_196),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_213),
.Y(n_221)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_214),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_205),
.A2(n_176),
.B1(n_181),
.B2(n_175),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_215),
.B(n_219),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_216),
.B(n_217),
.Y(n_229)
);

AOI21xp5_ASAP7_75t_L g217 ( 
.A1(n_203),
.A2(n_193),
.B(n_200),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_206),
.A2(n_172),
.B1(n_207),
.B2(n_201),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_220),
.B(n_211),
.C(n_202),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_L g226 ( 
.A1(n_223),
.A2(n_208),
.B(n_202),
.Y(n_226)
);

AOI21xp5_ASAP7_75t_L g233 ( 
.A1(n_226),
.A2(n_228),
.B(n_222),
.Y(n_233)
);

OR2x2_ASAP7_75t_L g234 ( 
.A(n_227),
.B(n_231),
.Y(n_234)
);

OAI21xp5_ASAP7_75t_L g228 ( 
.A1(n_220),
.A2(n_213),
.B(n_211),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_221),
.B(n_7),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_230),
.B(n_232),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_219),
.B(n_7),
.C(n_9),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_215),
.B(n_214),
.Y(n_232)
);

OAI21xp5_ASAP7_75t_L g244 ( 
.A1(n_233),
.A2(n_238),
.B(n_8),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_225),
.B(n_218),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_235),
.B(n_236),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_229),
.B(n_3),
.Y(n_236)
);

OR2x2_ASAP7_75t_L g238 ( 
.A(n_229),
.B(n_3),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_SL g239 ( 
.A(n_224),
.B(n_4),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_239),
.B(n_240),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_226),
.B(n_4),
.C(n_8),
.Y(n_240)
);

INVxp67_ASAP7_75t_L g241 ( 
.A(n_234),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_241),
.B(n_237),
.Y(n_246)
);

AND2x2_ASAP7_75t_L g242 ( 
.A(n_237),
.B(n_4),
.Y(n_242)
);

OAI21xp5_ASAP7_75t_L g247 ( 
.A1(n_242),
.A2(n_244),
.B(n_8),
.Y(n_247)
);

AOI21xp5_ASAP7_75t_L g248 ( 
.A1(n_246),
.A2(n_245),
.B(n_243),
.Y(n_248)
);

AO21x2_ASAP7_75t_L g249 ( 
.A1(n_247),
.A2(n_10),
.B(n_0),
.Y(n_249)
);

OAI21x1_ASAP7_75t_L g250 ( 
.A1(n_248),
.A2(n_249),
.B(n_10),
.Y(n_250)
);

BUFx24_ASAP7_75t_SL g251 ( 
.A(n_250),
.Y(n_251)
);

AOI21xp5_ASAP7_75t_L g252 ( 
.A1(n_251),
.A2(n_10),
.B(n_0),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_252),
.B(n_0),
.Y(n_253)
);


endmodule