module real_jpeg_5042_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_498;
wire n_369;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_366;
wire n_456;
wire n_259;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_21;
wire n_476;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_411;
wire n_382;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_215;
wire n_176;
wire n_166;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_502;
wire n_418;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_444;
wire n_178;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_368;
wire n_100;
wire n_51;
wire n_509;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

AOI22xp5_ASAP7_75t_L g18 ( 
.A1(n_0),
.A2(n_19),
.B1(n_22),
.B2(n_23),
.Y(n_18)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_1),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_2),
.B(n_36),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_2),
.B(n_77),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_2),
.B(n_117),
.Y(n_116)
);

AND2x2_ASAP7_75t_L g147 ( 
.A(n_2),
.B(n_148),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_2),
.B(n_187),
.Y(n_186)
);

AND2x2_ASAP7_75t_L g261 ( 
.A(n_2),
.B(n_262),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_2),
.B(n_290),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g431 ( 
.A(n_2),
.Y(n_431)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_3),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_3),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g196 ( 
.A(n_3),
.Y(n_196)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_3),
.Y(n_260)
);

BUFx6f_ASAP7_75t_L g304 ( 
.A(n_3),
.Y(n_304)
);

INVx3_ASAP7_75t_L g430 ( 
.A(n_3),
.Y(n_430)
);

BUFx5_ASAP7_75t_L g466 ( 
.A(n_3),
.Y(n_466)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_4),
.Y(n_37)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_4),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_5),
.B(n_64),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_5),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_5),
.B(n_128),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_5),
.B(n_334),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_SL g350 ( 
.A(n_5),
.B(n_351),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_5),
.B(n_152),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_6),
.B(n_43),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_6),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_6),
.B(n_133),
.Y(n_132)
);

AND2x2_ASAP7_75t_L g195 ( 
.A(n_6),
.B(n_196),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_6),
.B(n_380),
.Y(n_379)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_7),
.Y(n_41)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_7),
.Y(n_183)
);

BUFx6f_ASAP7_75t_L g349 ( 
.A(n_7),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_8),
.B(n_53),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_8),
.B(n_114),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_8),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_8),
.B(n_198),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_8),
.B(n_215),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_8),
.B(n_258),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_8),
.B(n_316),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_8),
.B(n_347),
.Y(n_346)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_9),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_10),
.B(n_39),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_10),
.Y(n_95)
);

AND2x2_ASAP7_75t_SL g175 ( 
.A(n_10),
.B(n_176),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_10),
.B(n_238),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_10),
.B(n_285),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_10),
.B(n_435),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_10),
.B(n_458),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_10),
.B(n_492),
.Y(n_491)
);

INVx3_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_12),
.Y(n_46)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_13),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_13),
.Y(n_88)
);

BUFx5_ASAP7_75t_L g104 ( 
.A(n_13),
.Y(n_104)
);

INVx3_ASAP7_75t_L g448 ( 
.A(n_13),
.Y(n_448)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_14),
.B(n_82),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_14),
.B(n_87),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_14),
.B(n_139),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_14),
.B(n_71),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_14),
.B(n_321),
.Y(n_320)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_14),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_14),
.B(n_368),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_14),
.B(n_326),
.Y(n_378)
);

INVx1_ASAP7_75t_SL g49 ( 
.A(n_15),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_15),
.B(n_109),
.Y(n_108)
);

AND2x2_ASAP7_75t_L g219 ( 
.A(n_15),
.B(n_98),
.Y(n_219)
);

AND2x2_ASAP7_75t_L g245 ( 
.A(n_15),
.B(n_246),
.Y(n_245)
);

AND2x2_ASAP7_75t_L g303 ( 
.A(n_15),
.B(n_304),
.Y(n_303)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_16),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g118 ( 
.A(n_16),
.Y(n_118)
);

INVx3_ASAP7_75t_L g154 ( 
.A(n_16),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_17),
.B(n_35),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_17),
.B(n_61),
.Y(n_60)
);

AND2x2_ASAP7_75t_L g151 ( 
.A(n_17),
.B(n_152),
.Y(n_151)
);

AND2x2_ASAP7_75t_SL g171 ( 
.A(n_17),
.B(n_172),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_17),
.B(n_71),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_17),
.B(n_277),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g444 ( 
.A(n_17),
.B(n_445),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_17),
.B(n_466),
.Y(n_465)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

INVx5_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

INVx6_ASAP7_75t_L g22 ( 
.A(n_21),
.Y(n_22)
);

XOR2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_503),
.Y(n_23)
);

OAI21xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_482),
.B(n_502),
.Y(n_24)
);

AOI21x1_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_422),
.B(n_479),
.Y(n_25)
);

AO21x1_ASAP7_75t_L g26 ( 
.A1(n_27),
.A2(n_270),
.B(n_306),
.Y(n_26)
);

OAI21xp5_ASAP7_75t_L g27 ( 
.A1(n_28),
.A2(n_227),
.B(n_269),
.Y(n_27)
);

AOI21xp5_ASAP7_75t_L g28 ( 
.A1(n_29),
.A2(n_202),
.B(n_226),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_29),
.B(n_420),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_160),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_30),
.B(n_160),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g30 ( 
.A(n_31),
.B(n_105),
.C(n_142),
.Y(n_30)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_31),
.B(n_225),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g31 ( 
.A(n_32),
.B(n_66),
.Y(n_31)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_32),
.B(n_67),
.C(n_84),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g32 ( 
.A(n_33),
.B(n_47),
.C(n_57),
.Y(n_32)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_33),
.B(n_222),
.Y(n_221)
);

BUFx24_ASAP7_75t_SL g518 ( 
.A(n_33),
.Y(n_518)
);

FAx1_ASAP7_75t_SL g33 ( 
.A(n_34),
.B(n_38),
.CI(n_42),
.CON(n_33),
.SN(n_33)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_34),
.B(n_38),
.C(n_42),
.Y(n_159)
);

BUFx2_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

BUFx8_ASAP7_75t_L g318 ( 
.A(n_37),
.Y(n_318)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_41),
.Y(n_79)
);

INVx2_ASAP7_75t_L g363 ( 
.A(n_41),
.Y(n_363)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx6_ASAP7_75t_L g130 ( 
.A(n_46),
.Y(n_130)
);

BUFx5_ASAP7_75t_L g437 ( 
.A(n_46),
.Y(n_437)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_47),
.A2(n_57),
.B1(n_58),
.B2(n_223),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_47),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g47 ( 
.A(n_48),
.B(n_52),
.C(n_56),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_48),
.A2(n_56),
.B1(n_181),
.B2(n_211),
.Y(n_210)
);

CKINVDCx16_ASAP7_75t_R g211 ( 
.A(n_48),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_48),
.A2(n_211),
.B1(n_219),
.B2(n_248),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_SL g449 ( 
.A1(n_48),
.A2(n_107),
.B1(n_108),
.B2(n_211),
.Y(n_449)
);

MAJIxp5_ASAP7_75t_L g451 ( 
.A(n_48),
.B(n_219),
.C(n_276),
.Y(n_451)
);

OR2x2_ASAP7_75t_L g48 ( 
.A(n_49),
.B(n_50),
.Y(n_48)
);

OR2x2_ASAP7_75t_SL g69 ( 
.A(n_49),
.B(n_70),
.Y(n_69)
);

OR2x2_ASAP7_75t_SL g168 ( 
.A(n_49),
.B(n_169),
.Y(n_168)
);

OR2x2_ASAP7_75t_L g182 ( 
.A(n_49),
.B(n_183),
.Y(n_182)
);

BUFx5_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g216 ( 
.A(n_51),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_SL g209 ( 
.A(n_52),
.B(n_210),
.Y(n_209)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx11_ASAP7_75t_L g111 ( 
.A(n_55),
.Y(n_111)
);

INVx3_ASAP7_75t_L g150 ( 
.A(n_55),
.Y(n_150)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_55),
.Y(n_174)
);

BUFx5_ASAP7_75t_L g352 ( 
.A(n_55),
.Y(n_352)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_56),
.A2(n_181),
.B1(n_182),
.B2(n_184),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_56),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_56),
.B(n_182),
.C(n_186),
.Y(n_233)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_59),
.B(n_62),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_59),
.A2(n_60),
.B1(n_62),
.B2(n_63),
.Y(n_220)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

XNOR2xp5_ASAP7_75t_L g66 ( 
.A(n_67),
.B(n_84),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_68),
.A2(n_69),
.B1(n_74),
.B2(n_75),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g464 ( 
.A1(n_68),
.A2(n_69),
.B1(n_107),
.B2(n_108),
.Y(n_464)
);

MAJIxp5_ASAP7_75t_L g493 ( 
.A(n_68),
.B(n_108),
.C(n_465),
.Y(n_493)
);

AOI22xp5_ASAP7_75t_L g499 ( 
.A1(n_68),
.A2(n_69),
.B1(n_167),
.B2(n_168),
.Y(n_499)
);

MAJIxp5_ASAP7_75t_L g509 ( 
.A(n_68),
.B(n_168),
.C(n_289),
.Y(n_509)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_69),
.B(n_76),
.C(n_81),
.Y(n_193)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_73),
.Y(n_114)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_73),
.Y(n_136)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_73),
.Y(n_187)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_76),
.A2(n_80),
.B1(n_81),
.B2(n_83),
.Y(n_75)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_76),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g341 ( 
.A1(n_76),
.A2(n_83),
.B1(n_126),
.B2(n_127),
.Y(n_341)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_81),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_83),
.B(n_126),
.Y(n_125)
);

XOR2xp5_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_93),
.Y(n_84)
);

OAI21xp5_ASAP7_75t_L g122 ( 
.A1(n_85),
.A2(n_86),
.B(n_89),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_85),
.B(n_94),
.C(n_101),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_86),
.B(n_89),
.Y(n_85)
);

INVx8_ASAP7_75t_L g459 ( 
.A(n_87),
.Y(n_459)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx4_ASAP7_75t_L g291 ( 
.A(n_88),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_90),
.B(n_92),
.Y(n_89)
);

INVx8_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g358 ( 
.A(n_92),
.B(n_359),
.Y(n_358)
);

XNOR2xp5_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_101),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_96),
.Y(n_94)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx3_ASAP7_75t_L g382 ( 
.A(n_98),
.Y(n_382)
);

INVx5_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g359 ( 
.A(n_99),
.Y(n_359)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_99),
.Y(n_370)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_103),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_102),
.B(n_325),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_102),
.B(n_337),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_102),
.B(n_373),
.Y(n_372)
);

INVx4_ASAP7_75t_L g246 ( 
.A(n_103),
.Y(n_246)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx6_ASAP7_75t_L g199 ( 
.A(n_104),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_105),
.B(n_142),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_106),
.B(n_121),
.C(n_123),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_106),
.A2(n_121),
.B1(n_122),
.B2(n_207),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_106),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_107),
.A2(n_108),
.B1(n_112),
.B2(n_120),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_108),
.B(n_113),
.C(n_116),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g462 ( 
.A(n_108),
.B(n_211),
.C(n_444),
.Y(n_462)
);

INVx6_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx6_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g323 ( 
.A(n_111),
.Y(n_323)
);

INVx5_ASAP7_75t_L g340 ( 
.A(n_111),
.Y(n_340)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_112),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_113),
.A2(n_115),
.B1(n_116),
.B2(n_119),
.Y(n_112)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_113),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_115),
.A2(n_116),
.B1(n_235),
.B2(n_240),
.Y(n_234)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_116),
.B(n_236),
.C(n_237),
.Y(n_280)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_SL g205 ( 
.A(n_123),
.B(n_206),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_131),
.C(n_137),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g408 ( 
.A1(n_124),
.A2(n_125),
.B1(n_409),
.B2(n_410),
.Y(n_408)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_130),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_130),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g262 ( 
.A(n_130),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g410 ( 
.A1(n_131),
.A2(n_132),
.B1(n_137),
.B2(n_138),
.Y(n_410)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVx5_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVx5_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVx4_ASAP7_75t_L g286 ( 
.A(n_136),
.Y(n_286)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx4_ASAP7_75t_SL g139 ( 
.A(n_140),
.Y(n_139)
);

INVx5_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVx3_ASAP7_75t_L g169 ( 
.A(n_141),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_159),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_145),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_144),
.B(n_145),
.C(n_159),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_SL g145 ( 
.A(n_146),
.B(n_155),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_151),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_147),
.B(n_151),
.C(n_155),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_147),
.A2(n_284),
.B1(n_287),
.B2(n_288),
.Y(n_283)
);

INVx1_ASAP7_75t_SL g288 ( 
.A(n_147),
.Y(n_288)
);

INVx5_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_150),
.Y(n_239)
);

INVx4_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

INVx4_ASAP7_75t_L g176 ( 
.A(n_154),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_157),
.Y(n_155)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

BUFx12f_ASAP7_75t_L g277 ( 
.A(n_158),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_162),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_161),
.B(n_163),
.C(n_201),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_163),
.A2(n_188),
.B1(n_200),
.B2(n_201),
.Y(n_162)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_163),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_178),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_166),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_165),
.B(n_166),
.C(n_178),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_167),
.A2(n_168),
.B1(n_170),
.B2(n_177),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g511 ( 
.A1(n_167),
.A2(n_168),
.B1(n_244),
.B2(n_245),
.Y(n_511)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_168),
.B(n_266),
.C(n_267),
.Y(n_265)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_170),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_175),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g266 ( 
.A(n_171),
.Y(n_266)
);

INVx4_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

INVx4_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_175),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_179),
.A2(n_180),
.B1(n_185),
.B2(n_186),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

CKINVDCx16_ASAP7_75t_R g184 ( 
.A(n_182),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g247 ( 
.A1(n_182),
.A2(n_184),
.B1(n_219),
.B2(n_248),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_182),
.B(n_219),
.C(n_245),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_SL g353 ( 
.A1(n_182),
.A2(n_184),
.B1(n_332),
.B2(n_333),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_SL g331 ( 
.A(n_184),
.B(n_332),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_L g433 ( 
.A1(n_185),
.A2(n_186),
.B1(n_434),
.B2(n_438),
.Y(n_433)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g460 ( 
.A(n_186),
.B(n_429),
.C(n_434),
.Y(n_460)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_188),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_SL g188 ( 
.A(n_189),
.B(n_190),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_189),
.B(n_191),
.C(n_192),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_192),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_194),
.Y(n_192)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_193),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_197),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_195),
.B(n_197),
.C(n_254),
.Y(n_253)
);

INVx4_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_224),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g420 ( 
.A(n_203),
.B(n_224),
.Y(n_420)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_208),
.C(n_221),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g414 ( 
.A1(n_204),
.A2(n_205),
.B1(n_415),
.B2(n_416),
.Y(n_414)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_SL g415 ( 
.A(n_208),
.B(n_221),
.Y(n_415)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_212),
.C(n_220),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g401 ( 
.A(n_209),
.B(n_402),
.Y(n_401)
);

XOR2xp5_ASAP7_75t_L g402 ( 
.A(n_212),
.B(n_220),
.Y(n_402)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_217),
.C(n_219),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_L g329 ( 
.A1(n_213),
.A2(n_214),
.B1(n_217),
.B2(n_218),
.Y(n_329)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

INVx3_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

INVx3_ASAP7_75t_L g326 ( 
.A(n_216),
.Y(n_326)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_219),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g327 ( 
.A1(n_219),
.A2(n_248),
.B1(n_328),
.B2(n_329),
.Y(n_327)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_228),
.B(n_270),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_230),
.Y(n_228)
);

OR2x2_ASAP7_75t_L g269 ( 
.A(n_229),
.B(n_230),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_230),
.B(n_271),
.Y(n_270)
);

OR2x2_ASAP7_75t_L g421 ( 
.A(n_230),
.B(n_271),
.Y(n_421)
);

FAx1_ASAP7_75t_SL g230 ( 
.A(n_231),
.B(n_250),
.CI(n_268),
.CON(n_230),
.SN(n_230)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_243),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_233),
.A2(n_234),
.B1(n_241),
.B2(n_242),
.Y(n_232)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_233),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_233),
.B(n_242),
.C(n_243),
.Y(n_295)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_234),
.Y(n_242)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_235),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_SL g235 ( 
.A(n_236),
.B(n_237),
.Y(n_235)
);

INVx4_ASAP7_75t_SL g238 ( 
.A(n_239),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_L g243 ( 
.A1(n_244),
.A2(n_245),
.B1(n_247),
.B2(n_249),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_247),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_SL g250 ( 
.A(n_251),
.B(n_252),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_251),
.B(n_253),
.C(n_255),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_255),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_265),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_257),
.A2(n_261),
.B1(n_263),
.B2(n_264),
.Y(n_256)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_257),
.Y(n_263)
);

BUFx6f_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_261),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_261),
.B(n_263),
.C(n_298),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_L g301 ( 
.A1(n_261),
.A2(n_264),
.B1(n_302),
.B2(n_303),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_SL g455 ( 
.A1(n_261),
.A2(n_264),
.B1(n_456),
.B2(n_457),
.Y(n_455)
);

MAJIxp5_ASAP7_75t_L g486 ( 
.A(n_261),
.B(n_456),
.C(n_460),
.Y(n_486)
);

MAJIxp5_ASAP7_75t_L g440 ( 
.A(n_264),
.B(n_300),
.C(n_303),
.Y(n_440)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_265),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_273),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g477 ( 
.A(n_272),
.B(n_274),
.C(n_293),
.Y(n_477)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_274),
.B(n_293),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_275),
.B(n_279),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g427 ( 
.A(n_275),
.B(n_280),
.C(n_281),
.Y(n_427)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_276),
.B(n_278),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_280),
.B(n_281),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_282),
.A2(n_283),
.B1(n_289),
.B2(n_292),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_284),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g450 ( 
.A(n_284),
.B(n_288),
.C(n_289),
.Y(n_450)
);

INVx6_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

INVx8_ASAP7_75t_L g334 ( 
.A(n_286),
.Y(n_334)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_289),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_SL g497 ( 
.A1(n_289),
.A2(n_292),
.B1(n_498),
.B2(n_499),
.Y(n_497)
);

INVx6_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_294),
.A2(n_295),
.B1(n_296),
.B2(n_305),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g475 ( 
.A(n_294),
.B(n_297),
.C(n_299),
.Y(n_475)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_296),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_SL g296 ( 
.A(n_297),
.B(n_299),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_300),
.B(n_301),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_303),
.Y(n_302)
);

OAI31xp33_ASAP7_75t_L g306 ( 
.A1(n_307),
.A2(n_418),
.A3(n_419),
.B(n_421),
.Y(n_306)
);

AOI21xp5_ASAP7_75t_L g307 ( 
.A1(n_308),
.A2(n_412),
.B(n_417),
.Y(n_307)
);

OAI21xp5_ASAP7_75t_SL g308 ( 
.A1(n_309),
.A2(n_397),
.B(n_411),
.Y(n_308)
);

AOI21xp5_ASAP7_75t_L g309 ( 
.A1(n_310),
.A2(n_354),
.B(n_396),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_SL g310 ( 
.A(n_311),
.B(n_342),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g396 ( 
.A(n_311),
.B(n_342),
.Y(n_396)
);

XNOR2xp5_ASAP7_75t_L g311 ( 
.A(n_312),
.B(n_330),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_313),
.B(n_327),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g398 ( 
.A(n_313),
.B(n_327),
.C(n_330),
.Y(n_398)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_314),
.B(n_319),
.C(n_324),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g344 ( 
.A1(n_314),
.A2(n_315),
.B1(n_319),
.B2(n_320),
.Y(n_344)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

INVx8_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

INVx3_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

XNOR2xp5_ASAP7_75t_SL g343 ( 
.A(n_324),
.B(n_344),
.Y(n_343)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

XNOR2xp5_ASAP7_75t_SL g330 ( 
.A(n_331),
.B(n_335),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g405 ( 
.A(n_331),
.B(n_406),
.C(n_407),
.Y(n_405)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);

XNOR2xp5_ASAP7_75t_L g335 ( 
.A(n_336),
.B(n_341),
.Y(n_335)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_336),
.Y(n_406)
);

INVx1_ASAP7_75t_SL g337 ( 
.A(n_338),
.Y(n_337)
);

BUFx3_ASAP7_75t_L g338 ( 
.A(n_339),
.Y(n_338)
);

INVx5_ASAP7_75t_L g339 ( 
.A(n_340),
.Y(n_339)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_341),
.Y(n_407)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_343),
.B(n_345),
.C(n_353),
.Y(n_342)
);

XNOR2xp5_ASAP7_75t_L g392 ( 
.A(n_343),
.B(n_393),
.Y(n_392)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_345),
.Y(n_388)
);

AOI22xp5_ASAP7_75t_L g393 ( 
.A1(n_345),
.A2(n_353),
.B1(n_388),
.B2(n_394),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_SL g345 ( 
.A(n_346),
.B(n_350),
.Y(n_345)
);

INVxp67_ASAP7_75t_L g386 ( 
.A(n_346),
.Y(n_386)
);

INVx2_ASAP7_75t_L g347 ( 
.A(n_348),
.Y(n_347)
);

INVx2_ASAP7_75t_L g348 ( 
.A(n_349),
.Y(n_348)
);

INVx3_ASAP7_75t_L g373 ( 
.A(n_349),
.Y(n_373)
);

INVxp67_ASAP7_75t_L g387 ( 
.A(n_350),
.Y(n_387)
);

INVx5_ASAP7_75t_L g351 ( 
.A(n_352),
.Y(n_351)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_353),
.Y(n_394)
);

OAI21xp5_ASAP7_75t_L g354 ( 
.A1(n_355),
.A2(n_390),
.B(n_395),
.Y(n_354)
);

AOI21xp5_ASAP7_75t_L g355 ( 
.A1(n_356),
.A2(n_375),
.B(n_389),
.Y(n_355)
);

OAI21xp5_ASAP7_75t_L g356 ( 
.A1(n_357),
.A2(n_364),
.B(n_374),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_358),
.B(n_360),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_L g360 ( 
.A(n_361),
.B(n_362),
.Y(n_360)
);

INVx4_ASAP7_75t_L g362 ( 
.A(n_363),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_SL g364 ( 
.A(n_365),
.B(n_372),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_365),
.B(n_372),
.Y(n_374)
);

AOI21xp5_ASAP7_75t_L g365 ( 
.A1(n_366),
.A2(n_367),
.B(n_371),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_L g371 ( 
.A(n_366),
.B(n_367),
.Y(n_371)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_369),
.Y(n_368)
);

INVx4_ASAP7_75t_L g369 ( 
.A(n_370),
.Y(n_369)
);

AOI22xp5_ASAP7_75t_L g376 ( 
.A1(n_371),
.A2(n_377),
.B1(n_383),
.B2(n_384),
.Y(n_376)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_371),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_SL g375 ( 
.A(n_376),
.B(n_385),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_L g389 ( 
.A(n_376),
.B(n_385),
.Y(n_389)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_377),
.Y(n_384)
);

XNOR2xp5_ASAP7_75t_SL g377 ( 
.A(n_378),
.B(n_379),
.Y(n_377)
);

OAI21xp5_ASAP7_75t_SL g391 ( 
.A1(n_378),
.A2(n_379),
.B(n_383),
.Y(n_391)
);

INVx2_ASAP7_75t_L g380 ( 
.A(n_381),
.Y(n_380)
);

HB1xp67_ASAP7_75t_L g381 ( 
.A(n_382),
.Y(n_381)
);

OAI21xp5_ASAP7_75t_SL g385 ( 
.A1(n_386),
.A2(n_387),
.B(n_388),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_L g390 ( 
.A(n_391),
.B(n_392),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_391),
.B(n_392),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_L g397 ( 
.A(n_398),
.B(n_399),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_398),
.B(n_399),
.Y(n_411)
);

OAI22xp5_ASAP7_75t_L g399 ( 
.A1(n_400),
.A2(n_401),
.B1(n_403),
.B2(n_404),
.Y(n_399)
);

MAJIxp5_ASAP7_75t_L g413 ( 
.A(n_400),
.B(n_405),
.C(n_408),
.Y(n_413)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_401),
.Y(n_400)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_404),
.Y(n_403)
);

XOR2xp5_ASAP7_75t_L g404 ( 
.A(n_405),
.B(n_408),
.Y(n_404)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_410),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_413),
.B(n_414),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_L g417 ( 
.A(n_413),
.B(n_414),
.Y(n_417)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_415),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_L g422 ( 
.A(n_423),
.B(n_476),
.Y(n_422)
);

OAI21xp5_ASAP7_75t_SL g479 ( 
.A1(n_423),
.A2(n_480),
.B(n_481),
.Y(n_479)
);

NOR2xp33_ASAP7_75t_L g423 ( 
.A(n_424),
.B(n_468),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_424),
.B(n_468),
.Y(n_481)
);

BUFx24_ASAP7_75t_SL g517 ( 
.A(n_424),
.Y(n_517)
);

FAx1_ASAP7_75t_SL g424 ( 
.A(n_425),
.B(n_441),
.CI(n_452),
.CON(n_424),
.SN(n_424)
);

MAJIxp5_ASAP7_75t_L g501 ( 
.A(n_425),
.B(n_441),
.C(n_452),
.Y(n_501)
);

MAJIxp5_ASAP7_75t_L g425 ( 
.A(n_426),
.B(n_428),
.C(n_440),
.Y(n_425)
);

AOI22xp5_ASAP7_75t_L g469 ( 
.A1(n_426),
.A2(n_427),
.B1(n_470),
.B2(n_471),
.Y(n_469)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_427),
.Y(n_426)
);

XOR2xp5_ASAP7_75t_L g470 ( 
.A(n_428),
.B(n_440),
.Y(n_470)
);

OAI22xp5_ASAP7_75t_L g428 ( 
.A1(n_429),
.A2(n_432),
.B1(n_433),
.B2(n_439),
.Y(n_428)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_429),
.Y(n_439)
);

AOI22xp5_ASAP7_75t_L g510 ( 
.A1(n_429),
.A2(n_439),
.B1(n_511),
.B2(n_512),
.Y(n_510)
);

NOR2xp33_ASAP7_75t_SL g429 ( 
.A(n_430),
.B(n_431),
.Y(n_429)
);

INVx6_ASAP7_75t_L g492 ( 
.A(n_430),
.Y(n_492)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_433),
.Y(n_432)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_434),
.Y(n_438)
);

INVx4_ASAP7_75t_L g435 ( 
.A(n_436),
.Y(n_435)
);

BUFx3_ASAP7_75t_L g436 ( 
.A(n_437),
.Y(n_436)
);

MAJIxp5_ASAP7_75t_L g441 ( 
.A(n_442),
.B(n_450),
.C(n_451),
.Y(n_441)
);

AOI22xp5_ASAP7_75t_L g472 ( 
.A1(n_442),
.A2(n_443),
.B1(n_473),
.B2(n_474),
.Y(n_472)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_443),
.Y(n_442)
);

XOR2xp5_ASAP7_75t_L g443 ( 
.A(n_444),
.B(n_449),
.Y(n_443)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_446),
.Y(n_445)
);

INVx6_ASAP7_75t_L g446 ( 
.A(n_447),
.Y(n_446)
);

INVx5_ASAP7_75t_L g447 ( 
.A(n_448),
.Y(n_447)
);

XOR2xp5_ASAP7_75t_L g474 ( 
.A(n_450),
.B(n_451),
.Y(n_474)
);

AOI22xp5_ASAP7_75t_L g452 ( 
.A1(n_453),
.A2(n_454),
.B1(n_461),
.B2(n_467),
.Y(n_452)
);

MAJIxp5_ASAP7_75t_L g500 ( 
.A(n_453),
.B(n_462),
.C(n_463),
.Y(n_500)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_454),
.Y(n_453)
);

XNOR2xp5_ASAP7_75t_SL g454 ( 
.A(n_455),
.B(n_460),
.Y(n_454)
);

CKINVDCx14_ASAP7_75t_R g456 ( 
.A(n_457),
.Y(n_456)
);

INVx3_ASAP7_75t_L g458 ( 
.A(n_459),
.Y(n_458)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_461),
.Y(n_467)
);

XNOR2xp5_ASAP7_75t_SL g461 ( 
.A(n_462),
.B(n_463),
.Y(n_461)
);

XNOR2xp5_ASAP7_75t_L g463 ( 
.A(n_464),
.B(n_465),
.Y(n_463)
);

MAJIxp5_ASAP7_75t_L g468 ( 
.A(n_469),
.B(n_472),
.C(n_475),
.Y(n_468)
);

FAx1_ASAP7_75t_SL g478 ( 
.A(n_469),
.B(n_472),
.CI(n_475),
.CON(n_478),
.SN(n_478)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_470),
.Y(n_471)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_474),
.Y(n_473)
);

NOR2xp33_ASAP7_75t_L g476 ( 
.A(n_477),
.B(n_478),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_477),
.B(n_478),
.Y(n_480)
);

BUFx24_ASAP7_75t_SL g520 ( 
.A(n_478),
.Y(n_520)
);

NOR2xp33_ASAP7_75t_L g482 ( 
.A(n_483),
.B(n_501),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_483),
.B(n_501),
.Y(n_502)
);

XOR2xp5_ASAP7_75t_L g483 ( 
.A(n_484),
.B(n_500),
.Y(n_483)
);

AOI22xp5_ASAP7_75t_L g484 ( 
.A1(n_485),
.A2(n_486),
.B1(n_487),
.B2(n_488),
.Y(n_484)
);

CKINVDCx16_ASAP7_75t_R g485 ( 
.A(n_486),
.Y(n_485)
);

MAJIxp5_ASAP7_75t_L g515 ( 
.A(n_486),
.B(n_487),
.C(n_500),
.Y(n_515)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_488),
.Y(n_487)
);

OAI22xp5_ASAP7_75t_SL g488 ( 
.A1(n_489),
.A2(n_490),
.B1(n_496),
.B2(n_497),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_490),
.Y(n_489)
);

AOI22xp5_ASAP7_75t_L g490 ( 
.A1(n_491),
.A2(n_493),
.B1(n_494),
.B2(n_495),
.Y(n_490)
);

CKINVDCx20_ASAP7_75t_R g494 ( 
.A(n_491),
.Y(n_494)
);

CKINVDCx14_ASAP7_75t_R g495 ( 
.A(n_493),
.Y(n_495)
);

MAJIxp5_ASAP7_75t_L g507 ( 
.A(n_493),
.B(n_494),
.C(n_496),
.Y(n_507)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_497),
.Y(n_496)
);

CKINVDCx16_ASAP7_75t_R g498 ( 
.A(n_499),
.Y(n_498)
);

NOR2xp33_ASAP7_75t_L g503 ( 
.A(n_504),
.B(n_516),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_505),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_506),
.B(n_515),
.Y(n_505)
);

NOR2xp33_ASAP7_75t_L g516 ( 
.A(n_506),
.B(n_515),
.Y(n_516)
);

XNOR2xp5_ASAP7_75t_L g506 ( 
.A(n_507),
.B(n_508),
.Y(n_506)
);

AOI22xp5_ASAP7_75t_L g508 ( 
.A1(n_509),
.A2(n_510),
.B1(n_513),
.B2(n_514),
.Y(n_508)
);

CKINVDCx20_ASAP7_75t_R g513 ( 
.A(n_509),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_510),
.Y(n_514)
);

CKINVDCx20_ASAP7_75t_R g512 ( 
.A(n_511),
.Y(n_512)
);


endmodule