module fake_jpeg_27872_n_164 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_164);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_164;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_11;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g11 ( 
.A(n_6),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_2),
.Y(n_12)
);

BUFx12f_ASAP7_75t_L g13 ( 
.A(n_6),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_1),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_7),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

INVx13_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_8),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_10),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_13),
.B(n_0),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_22),
.B(n_27),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_23),
.Y(n_38)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_24),
.Y(n_37)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_25),
.Y(n_36)
);

INVx11_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_26),
.Y(n_31)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_SL g30 ( 
.A(n_28),
.B(n_29),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

MAJIxp5_ASAP7_75t_L g32 ( 
.A(n_22),
.B(n_11),
.C(n_20),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_32),
.B(n_35),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g34 ( 
.A1(n_22),
.A2(n_17),
.B1(n_20),
.B2(n_19),
.Y(n_34)
);

AOI22xp5_ASAP7_75t_L g45 ( 
.A1(n_34),
.A2(n_17),
.B1(n_19),
.B2(n_15),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g35 ( 
.A(n_23),
.B(n_20),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_37),
.Y(n_39)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_38),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_40),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_L g41 ( 
.A1(n_33),
.A2(n_17),
.B1(n_27),
.B2(n_25),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_41),
.A2(n_30),
.B1(n_46),
.B2(n_26),
.Y(n_65)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_30),
.Y(n_43)
);

OAI21xp33_ASAP7_75t_L g59 ( 
.A1(n_43),
.A2(n_44),
.B(n_35),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g44 ( 
.A1(n_37),
.A2(n_17),
.B1(n_21),
.B2(n_18),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_45),
.A2(n_49),
.B1(n_36),
.B2(n_26),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_33),
.B(n_27),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_46),
.B(n_48),
.Y(n_63)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_37),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_47),
.B(n_31),
.Y(n_58)
);

CKINVDCx14_ASAP7_75t_R g48 ( 
.A(n_34),
.Y(n_48)
);

OA22x2_ASAP7_75t_L g49 ( 
.A1(n_31),
.A2(n_26),
.B1(n_25),
.B2(n_36),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_33),
.B(n_32),
.Y(n_50)
);

XNOR2xp5_ASAP7_75t_L g55 ( 
.A(n_50),
.B(n_51),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_32),
.B(n_29),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_49),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_52),
.B(n_54),
.Y(n_67)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_49),
.Y(n_54)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_49),
.Y(n_56)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_56),
.Y(n_66)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_58),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_L g76 ( 
.A1(n_59),
.A2(n_37),
.B1(n_14),
.B2(n_15),
.Y(n_76)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_49),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_60),
.B(n_28),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_43),
.B(n_35),
.Y(n_61)
);

INVxp67_ASAP7_75t_L g75 ( 
.A(n_61),
.Y(n_75)
);

XOR2xp5_ASAP7_75t_L g62 ( 
.A(n_50),
.B(n_34),
.Y(n_62)
);

MAJIxp5_ASAP7_75t_L g70 ( 
.A(n_62),
.B(n_42),
.C(n_51),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_64),
.A2(n_52),
.B1(n_60),
.B2(n_56),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_65),
.A2(n_30),
.B1(n_31),
.B2(n_25),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_64),
.A2(n_48),
.B1(n_45),
.B2(n_21),
.Y(n_68)
);

INVxp67_ASAP7_75t_L g78 ( 
.A(n_68),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_70),
.B(n_62),
.C(n_55),
.Y(n_82)
);

OR2x2_ASAP7_75t_L g71 ( 
.A(n_65),
.B(n_42),
.Y(n_71)
);

A2O1A1Ixp33_ASAP7_75t_L g89 ( 
.A1(n_71),
.A2(n_12),
.B(n_19),
.C(n_16),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_72),
.A2(n_55),
.B1(n_53),
.B2(n_36),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_73),
.A2(n_77),
.B1(n_63),
.B2(n_53),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_74),
.B(n_29),
.Y(n_80)
);

INVx1_ASAP7_75t_SL g87 ( 
.A(n_76),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_54),
.A2(n_36),
.B1(n_29),
.B2(n_28),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_79),
.B(n_68),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_80),
.B(n_74),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_67),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_81),
.B(n_86),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_82),
.B(n_70),
.C(n_71),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g83 ( 
.A(n_69),
.B(n_75),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_83),
.B(n_85),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_84),
.A2(n_88),
.B1(n_38),
.B2(n_28),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_69),
.B(n_18),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_67),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_66),
.A2(n_57),
.B1(n_47),
.B2(n_38),
.Y(n_88)
);

XOR2xp5_ASAP7_75t_L g102 ( 
.A(n_89),
.B(n_80),
.Y(n_102)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_88),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_91),
.B(n_96),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_92),
.B(n_11),
.C(n_24),
.Y(n_115)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_93),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_81),
.B(n_66),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_95),
.B(n_102),
.Y(n_105)
);

AOI21xp5_ASAP7_75t_L g97 ( 
.A1(n_86),
.A2(n_72),
.B(n_77),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_L g103 ( 
.A1(n_97),
.A2(n_95),
.B(n_78),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_84),
.B(n_75),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_98),
.B(n_99),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_79),
.B(n_57),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_100),
.A2(n_78),
.B1(n_87),
.B2(n_82),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_87),
.B(n_39),
.Y(n_101)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_101),
.Y(n_112)
);

AOI21xp5_ASAP7_75t_SL g116 ( 
.A1(n_103),
.A2(n_16),
.B(n_15),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_106),
.A2(n_23),
.B1(n_24),
.B2(n_16),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_97),
.A2(n_89),
.B1(n_38),
.B2(n_28),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_107),
.A2(n_114),
.B1(n_14),
.B2(n_12),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_94),
.B(n_39),
.Y(n_108)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_108),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_92),
.B(n_40),
.C(n_29),
.Y(n_111)
);

XOR2xp5_ASAP7_75t_L g121 ( 
.A(n_111),
.B(n_115),
.Y(n_121)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_93),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_113),
.B(n_14),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_100),
.A2(n_102),
.B1(n_90),
.B2(n_40),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_L g132 ( 
.A(n_116),
.B(n_127),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_117),
.B(n_124),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_119),
.A2(n_126),
.B1(n_112),
.B2(n_104),
.Y(n_133)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_108),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_120),
.B(n_123),
.Y(n_129)
);

XOR2xp5_ASAP7_75t_L g122 ( 
.A(n_111),
.B(n_24),
.Y(n_122)
);

XOR2xp5_ASAP7_75t_L g130 ( 
.A(n_122),
.B(n_115),
.Y(n_130)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_105),
.Y(n_123)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_105),
.Y(n_124)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_114),
.Y(n_125)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_125),
.Y(n_128)
);

A2O1A1Ixp33_ASAP7_75t_SL g126 ( 
.A1(n_103),
.A2(n_23),
.B(n_0),
.C(n_2),
.Y(n_126)
);

AND2x2_ASAP7_75t_L g141 ( 
.A(n_130),
.B(n_134),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_133),
.A2(n_136),
.B1(n_131),
.B2(n_128),
.Y(n_143)
);

XOR2xp5_ASAP7_75t_L g134 ( 
.A(n_121),
.B(n_106),
.Y(n_134)
);

XOR2xp5_ASAP7_75t_L g135 ( 
.A(n_118),
.B(n_110),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_135),
.B(n_137),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_127),
.A2(n_109),
.B1(n_107),
.B2(n_2),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_126),
.B(n_6),
.C(n_1),
.Y(n_137)
);

AOI21xp5_ASAP7_75t_L g138 ( 
.A1(n_129),
.A2(n_126),
.B(n_116),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_138),
.B(n_140),
.Y(n_151)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_135),
.Y(n_140)
);

OAI21x1_ASAP7_75t_L g142 ( 
.A1(n_130),
.A2(n_7),
.B(n_3),
.Y(n_142)
);

AND2x2_ASAP7_75t_L g149 ( 
.A(n_142),
.B(n_4),
.Y(n_149)
);

INVxp67_ASAP7_75t_L g146 ( 
.A(n_143),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_132),
.B(n_4),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g147 ( 
.A(n_144),
.Y(n_147)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_134),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_145),
.B(n_4),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_148),
.B(n_5),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_149),
.B(n_150),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_139),
.B(n_5),
.C(n_8),
.Y(n_150)
);

BUFx24_ASAP7_75t_SL g152 ( 
.A(n_146),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_152),
.B(n_153),
.Y(n_157)
);

AOI21xp5_ASAP7_75t_L g153 ( 
.A1(n_151),
.A2(n_141),
.B(n_144),
.Y(n_153)
);

NOR2x1_ASAP7_75t_SL g155 ( 
.A(n_147),
.B(n_5),
.Y(n_155)
);

AOI21x1_ASAP7_75t_L g160 ( 
.A1(n_155),
.A2(n_9),
.B(n_10),
.Y(n_160)
);

INVxp67_ASAP7_75t_L g158 ( 
.A(n_156),
.Y(n_158)
);

AOI21xp5_ASAP7_75t_L g159 ( 
.A1(n_154),
.A2(n_8),
.B(n_9),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_159),
.B(n_157),
.C(n_158),
.Y(n_162)
);

MAJx2_ASAP7_75t_L g161 ( 
.A(n_160),
.B(n_9),
.C(n_10),
.Y(n_161)
);

NAND3xp33_ASAP7_75t_SL g163 ( 
.A(n_161),
.B(n_162),
.C(n_0),
.Y(n_163)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_163),
.B(n_0),
.Y(n_164)
);


endmodule