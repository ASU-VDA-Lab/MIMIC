module fake_jpeg_32094_n_313 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_313);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_313;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_19;
wire n_182;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_8),
.Y(n_18)
);

INVxp67_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_14),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

INVx6_ASAP7_75t_SL g22 ( 
.A(n_0),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

INVx1_ASAP7_75t_SL g24 ( 
.A(n_15),
.Y(n_24)
);

BUFx10_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_15),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_15),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_17),
.Y(n_29)
);

INVx11_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_7),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_6),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_1),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_8),
.Y(n_37)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_13),
.Y(n_38)
);

INVx3_ASAP7_75t_SL g39 ( 
.A(n_38),
.Y(n_39)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_39),
.Y(n_76)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_38),
.Y(n_40)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_23),
.Y(n_41)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_30),
.Y(n_42)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_42),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_24),
.B(n_0),
.Y(n_43)
);

AND2x2_ASAP7_75t_L g51 ( 
.A(n_43),
.B(n_24),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_30),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_44),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_30),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_45),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_29),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_46),
.Y(n_69)
);

INVx5_ASAP7_75t_L g47 ( 
.A(n_38),
.Y(n_47)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_47),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_29),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_48),
.Y(n_77)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_27),
.Y(n_49)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_49),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_43),
.B(n_20),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_50),
.B(n_54),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_51),
.B(n_34),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_41),
.B(n_20),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_39),
.B(n_37),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_56),
.B(n_64),
.Y(n_105)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_46),
.Y(n_57)
);

INVx6_ASAP7_75t_L g116 ( 
.A(n_57),
.Y(n_116)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_49),
.Y(n_58)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_58),
.Y(n_98)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_44),
.Y(n_62)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_62),
.Y(n_93)
);

BUFx5_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_63),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_39),
.B(n_37),
.Y(n_64)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_40),
.Y(n_65)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_65),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_46),
.B(n_24),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_66),
.B(n_25),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_48),
.A2(n_27),
.B1(n_36),
.B2(n_29),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_67),
.A2(n_26),
.B1(n_33),
.B2(n_32),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_42),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_70),
.B(n_72),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_L g71 ( 
.A1(n_48),
.A2(n_27),
.B1(n_29),
.B2(n_36),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_71),
.A2(n_66),
.B1(n_76),
.B2(n_53),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_44),
.Y(n_72)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_40),
.Y(n_73)
);

INVx1_ASAP7_75t_SL g79 ( 
.A(n_73),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_47),
.A2(n_22),
.B1(n_35),
.B2(n_23),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_74),
.A2(n_78),
.B1(n_22),
.B2(n_36),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_45),
.B(n_28),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_75),
.B(n_18),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_45),
.A2(n_22),
.B1(n_35),
.B2(n_23),
.Y(n_78)
);

A2O1A1Ixp33_ASAP7_75t_L g80 ( 
.A1(n_51),
.A2(n_19),
.B(n_21),
.C(n_34),
.Y(n_80)
);

A2O1A1Ixp33_ASAP7_75t_L g138 ( 
.A1(n_80),
.A2(n_105),
.B(n_86),
.C(n_100),
.Y(n_138)
);

HB1xp67_ASAP7_75t_L g82 ( 
.A(n_65),
.Y(n_82)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_82),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_84),
.A2(n_4),
.B1(n_5),
.B2(n_7),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_L g85 ( 
.A1(n_67),
.A2(n_35),
.B1(n_23),
.B2(n_36),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_85),
.A2(n_77),
.B1(n_68),
.B2(n_55),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_86),
.B(n_99),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_87),
.A2(n_88),
.B1(n_102),
.B2(n_103),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_76),
.A2(n_35),
.B1(n_23),
.B2(n_21),
.Y(n_89)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_89),
.Y(n_117)
);

NAND2xp33_ASAP7_75t_SL g91 ( 
.A(n_53),
.B(n_58),
.Y(n_91)
);

NAND2xp33_ASAP7_75t_SL g148 ( 
.A(n_91),
.B(n_94),
.Y(n_148)
);

HB1xp67_ASAP7_75t_L g92 ( 
.A(n_73),
.Y(n_92)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_92),
.Y(n_139)
);

INVx1_ASAP7_75t_SL g94 ( 
.A(n_59),
.Y(n_94)
);

BUFx12f_ASAP7_75t_L g95 ( 
.A(n_59),
.Y(n_95)
);

CKINVDCx14_ASAP7_75t_R g133 ( 
.A(n_95),
.Y(n_133)
);

INVx13_ASAP7_75t_L g97 ( 
.A(n_60),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_97),
.B(n_106),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_51),
.B(n_31),
.Y(n_100)
);

FAx1_ASAP7_75t_SL g119 ( 
.A(n_100),
.B(n_113),
.CI(n_25),
.CON(n_119),
.SN(n_119)
);

OA21x2_ASAP7_75t_L g101 ( 
.A1(n_72),
.A2(n_31),
.B(n_25),
.Y(n_101)
);

OA22x2_ASAP7_75t_L g132 ( 
.A1(n_101),
.A2(n_88),
.B1(n_94),
.B2(n_79),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_57),
.A2(n_33),
.B1(n_32),
.B2(n_28),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_60),
.A2(n_35),
.B1(n_26),
.B2(n_18),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_70),
.B(n_25),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_104),
.B(n_108),
.Y(n_126)
);

INVx13_ASAP7_75t_L g106 ( 
.A(n_52),
.Y(n_106)
);

BUFx12_ASAP7_75t_L g107 ( 
.A(n_61),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_107),
.B(n_111),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_62),
.Y(n_108)
);

HB1xp67_ASAP7_75t_L g109 ( 
.A(n_61),
.Y(n_109)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_109),
.Y(n_134)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_52),
.Y(n_110)
);

INVx4_ASAP7_75t_L g141 ( 
.A(n_110),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_63),
.B(n_16),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_112),
.B(n_114),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_69),
.B(n_25),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_69),
.B(n_16),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g115 ( 
.A(n_69),
.B(n_0),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_115),
.B(n_1),
.Y(n_128)
);

AND2x2_ASAP7_75t_L g165 ( 
.A(n_119),
.B(n_132),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_83),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_121),
.B(n_138),
.Y(n_163)
);

HB1xp67_ASAP7_75t_L g123 ( 
.A(n_93),
.Y(n_123)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_123),
.Y(n_156)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_98),
.Y(n_124)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_124),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_L g127 ( 
.A(n_99),
.B(n_25),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_127),
.B(n_135),
.C(n_142),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_SL g152 ( 
.A(n_128),
.B(n_144),
.Y(n_152)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_98),
.Y(n_129)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_129),
.Y(n_168)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_96),
.Y(n_130)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_130),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_86),
.B(n_77),
.C(n_68),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_136),
.A2(n_146),
.B1(n_108),
.B2(n_101),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_SL g137 ( 
.A(n_80),
.B(n_2),
.C(n_3),
.Y(n_137)
);

AND2x2_ASAP7_75t_L g166 ( 
.A(n_137),
.B(n_9),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_110),
.A2(n_68),
.B1(n_55),
.B2(n_4),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g155 ( 
.A(n_140),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_100),
.B(n_55),
.C(n_3),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_96),
.Y(n_143)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_143),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_81),
.B(n_2),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_87),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_147),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_181)
);

AOI21xp5_ASAP7_75t_SL g149 ( 
.A1(n_104),
.A2(n_5),
.B(n_7),
.Y(n_149)
);

OR2x2_ASAP7_75t_L g151 ( 
.A(n_149),
.B(n_8),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_127),
.B(n_115),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_150),
.B(n_172),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_151),
.B(n_157),
.Y(n_184)
);

AOI21xp5_ASAP7_75t_L g153 ( 
.A1(n_117),
.A2(n_90),
.B(n_79),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_SL g197 ( 
.A1(n_153),
.A2(n_175),
.B(n_130),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_126),
.Y(n_157)
);

INVx3_ASAP7_75t_SL g158 ( 
.A(n_141),
.Y(n_158)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_158),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_159),
.A2(n_167),
.B1(n_132),
.B2(n_142),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_131),
.B(n_101),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_160),
.B(n_164),
.Y(n_192)
);

AOI22xp33_ASAP7_75t_SL g162 ( 
.A1(n_117),
.A2(n_95),
.B1(n_90),
.B2(n_93),
.Y(n_162)
);

INVxp67_ASAP7_75t_L g206 ( 
.A(n_162),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_138),
.B(n_113),
.Y(n_164)
);

INVxp67_ASAP7_75t_L g209 ( 
.A(n_166),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_120),
.A2(n_91),
.B1(n_116),
.B2(n_106),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_145),
.B(n_116),
.C(n_97),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_169),
.B(n_179),
.Y(n_191)
);

BUFx12_ASAP7_75t_L g170 ( 
.A(n_133),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_170),
.B(n_180),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_122),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_171),
.B(n_177),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_145),
.B(n_95),
.Y(n_172)
);

INVx13_ASAP7_75t_L g173 ( 
.A(n_148),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g186 ( 
.A(n_173),
.Y(n_186)
);

AND2x2_ASAP7_75t_L g175 ( 
.A(n_132),
.B(n_95),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_125),
.Y(n_177)
);

INVx4_ASAP7_75t_L g178 ( 
.A(n_141),
.Y(n_178)
);

INVx4_ASAP7_75t_L g183 ( 
.A(n_178),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_119),
.B(n_107),
.C(n_10),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_124),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_181),
.B(n_147),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_L g185 ( 
.A1(n_165),
.A2(n_137),
.B(n_149),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_L g220 ( 
.A1(n_185),
.A2(n_209),
.B(n_166),
.Y(n_220)
);

CKINVDCx14_ASAP7_75t_R g213 ( 
.A(n_187),
.Y(n_213)
);

AO32x1_ASAP7_75t_L g189 ( 
.A1(n_165),
.A2(n_132),
.A3(n_119),
.B1(n_146),
.B2(n_135),
.Y(n_189)
);

AOI21xp5_ASAP7_75t_SL g231 ( 
.A1(n_189),
.A2(n_172),
.B(n_169),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_193),
.A2(n_202),
.B1(n_208),
.B2(n_181),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_165),
.B(n_143),
.Y(n_194)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_194),
.Y(n_234)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_174),
.Y(n_195)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_195),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_171),
.B(n_134),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_196),
.B(n_198),
.Y(n_219)
);

INVx1_ASAP7_75t_SL g211 ( 
.A(n_197),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_152),
.B(n_139),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_174),
.Y(n_199)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_199),
.Y(n_222)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_176),
.Y(n_200)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_200),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_161),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_201),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_159),
.A2(n_136),
.B1(n_129),
.B2(n_139),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_176),
.Y(n_203)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_203),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_SL g205 ( 
.A(n_163),
.B(n_11),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_205),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_175),
.A2(n_118),
.B1(n_12),
.B2(n_13),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_207),
.A2(n_151),
.B1(n_155),
.B2(n_209),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_167),
.A2(n_118),
.B1(n_13),
.B2(n_14),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_161),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_210),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g239 ( 
.A1(n_212),
.A2(n_216),
.B1(n_229),
.B2(n_213),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_190),
.B(n_154),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_215),
.B(n_217),
.C(n_218),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_189),
.A2(n_175),
.B1(n_153),
.B2(n_155),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_190),
.B(n_154),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_191),
.B(n_150),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_220),
.B(n_233),
.Y(n_244)
);

NAND4xp25_ASAP7_75t_SL g221 ( 
.A(n_207),
.B(n_170),
.C(n_158),
.D(n_107),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_221),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_224),
.A2(n_206),
.B1(n_189),
.B2(n_186),
.Y(n_236)
);

INVx1_ASAP7_75t_SL g225 ( 
.A(n_186),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_225),
.B(n_188),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_206),
.A2(n_166),
.B1(n_173),
.B2(n_156),
.Y(n_229)
);

INVxp67_ASAP7_75t_L g242 ( 
.A(n_229),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_231),
.B(n_232),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_204),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_191),
.B(n_194),
.C(n_192),
.Y(n_233)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_235),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_236),
.B(n_216),
.Y(n_258)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_214),
.Y(n_238)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_238),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_239),
.A2(n_252),
.B1(n_211),
.B2(n_224),
.Y(n_260)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_222),
.Y(n_240)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_240),
.Y(n_270)
);

INVx1_ASAP7_75t_SL g241 ( 
.A(n_226),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_241),
.B(n_248),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_SL g243 ( 
.A(n_227),
.B(n_184),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g257 ( 
.A(n_243),
.B(n_249),
.Y(n_257)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_230),
.Y(n_245)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_245),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_223),
.B(n_210),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_SL g249 ( 
.A(n_219),
.B(n_205),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_212),
.A2(n_185),
.B1(n_201),
.B2(n_186),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_250),
.B(n_251),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_228),
.B(n_199),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_234),
.A2(n_197),
.B1(n_195),
.B2(n_188),
.Y(n_252)
);

INVx1_ASAP7_75t_SL g253 ( 
.A(n_221),
.Y(n_253)
);

AND2x2_ASAP7_75t_L g265 ( 
.A(n_253),
.B(n_225),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_248),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_254),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_258),
.A2(n_260),
.B1(n_261),
.B2(n_269),
.Y(n_278)
);

AOI21xp5_ASAP7_75t_L g259 ( 
.A1(n_246),
.A2(n_211),
.B(n_234),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_259),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_247),
.A2(n_217),
.B1(n_215),
.B2(n_218),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_237),
.B(n_244),
.C(n_233),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_262),
.B(n_242),
.C(n_220),
.Y(n_271)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_265),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_251),
.B(n_182),
.Y(n_266)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_266),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_237),
.B(n_244),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_267),
.B(n_236),
.Y(n_273)
);

XOR2x2_ASAP7_75t_SL g269 ( 
.A(n_242),
.B(n_231),
.Y(n_269)
);

AOI21xp33_ASAP7_75t_SL g277 ( 
.A1(n_269),
.A2(n_247),
.B(n_253),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_271),
.B(n_259),
.C(n_264),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_SL g292 ( 
.A(n_273),
.B(n_276),
.Y(n_292)
);

XOR2xp5_ASAP7_75t_L g276 ( 
.A(n_267),
.B(n_252),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_277),
.B(n_283),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_278),
.B(n_260),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_262),
.B(n_235),
.C(n_241),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_279),
.B(n_282),
.C(n_273),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_255),
.B(n_245),
.Y(n_280)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_280),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_261),
.B(n_179),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_255),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_285),
.B(n_286),
.Y(n_298)
);

OAI21xp5_ASAP7_75t_SL g287 ( 
.A1(n_271),
.A2(n_257),
.B(n_264),
.Y(n_287)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_287),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_280),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g299 ( 
.A(n_289),
.B(n_290),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_SL g290 ( 
.A(n_275),
.B(n_270),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_291),
.B(n_292),
.C(n_276),
.Y(n_293)
);

XOR2xp5_ASAP7_75t_L g300 ( 
.A(n_293),
.B(n_288),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_L g294 ( 
.A1(n_284),
.A2(n_272),
.B1(n_281),
.B2(n_256),
.Y(n_294)
);

HB1xp67_ASAP7_75t_L g303 ( 
.A(n_294),
.Y(n_303)
);

OAI21xp5_ASAP7_75t_L g295 ( 
.A1(n_291),
.A2(n_279),
.B(n_274),
.Y(n_295)
);

AOI21xp5_ASAP7_75t_SL g304 ( 
.A1(n_295),
.A2(n_240),
.B(n_238),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_292),
.B(n_278),
.C(n_282),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_SL g301 ( 
.A1(n_297),
.A2(n_265),
.B(n_268),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_300),
.B(n_293),
.C(n_297),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_SL g307 ( 
.A(n_301),
.B(n_302),
.Y(n_307)
);

OAI21xp5_ASAP7_75t_SL g302 ( 
.A1(n_296),
.A2(n_265),
.B(n_263),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_SL g305 ( 
.A(n_304),
.B(n_299),
.Y(n_305)
);

OAI21xp5_ASAP7_75t_L g308 ( 
.A1(n_305),
.A2(n_303),
.B(n_298),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_306),
.B(n_156),
.Y(n_309)
);

OAI21x1_ASAP7_75t_SL g310 ( 
.A1(n_308),
.A2(n_309),
.B(n_307),
.Y(n_310)
);

AOI322xp5_ASAP7_75t_L g311 ( 
.A1(n_310),
.A2(n_203),
.A3(n_200),
.B1(n_168),
.B2(n_183),
.C1(n_170),
.C2(n_178),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_311),
.A2(n_183),
.B1(n_168),
.B2(n_14),
.Y(n_312)
);

XOR2xp5_ASAP7_75t_L g313 ( 
.A(n_312),
.B(n_11),
.Y(n_313)
);


endmodule