module fake_jpeg_35_n_184 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_184);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_184;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_175;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g12 ( 
.A(n_2),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_6),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_0),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_2),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_8),
.Y(n_16)
);

CKINVDCx5p33_ASAP7_75t_R g17 ( 
.A(n_0),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_7),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_7),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_9),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_1),
.Y(n_30)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_29),
.Y(n_31)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_31),
.Y(n_63)
);

INVx5_ASAP7_75t_L g32 ( 
.A(n_17),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_32),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_18),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_33),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_18),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_34),
.Y(n_69)
);

INVx1_ASAP7_75t_SL g35 ( 
.A(n_29),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g82 ( 
.A(n_35),
.Y(n_82)
);

HB1xp67_ASAP7_75t_L g36 ( 
.A(n_22),
.Y(n_36)
);

CKINVDCx16_ASAP7_75t_R g78 ( 
.A(n_36),
.Y(n_78)
);

AOI21xp33_ASAP7_75t_L g37 ( 
.A1(n_12),
.A2(n_1),
.B(n_2),
.Y(n_37)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_37),
.B(n_4),
.C(n_9),
.Y(n_77)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

INVx11_ASAP7_75t_L g76 ( 
.A(n_38),
.Y(n_76)
);

INVx2_ASAP7_75t_SL g39 ( 
.A(n_29),
.Y(n_39)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_40),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g41 ( 
.A(n_14),
.B(n_30),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_41),
.B(n_47),
.Y(n_59)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_22),
.Y(n_42)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_42),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_28),
.Y(n_43)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_43),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g44 ( 
.A(n_12),
.B(n_1),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_44),
.B(n_4),
.Y(n_84)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_28),
.Y(n_45)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_45),
.Y(n_70)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_13),
.Y(n_46)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_46),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_14),
.B(n_3),
.Y(n_47)
);

BUFx12_ASAP7_75t_L g48 ( 
.A(n_17),
.Y(n_48)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_48),
.Y(n_67)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_13),
.Y(n_49)
);

BUFx2_ASAP7_75t_L g81 ( 
.A(n_49),
.Y(n_81)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_23),
.Y(n_50)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_50),
.Y(n_71)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_15),
.Y(n_51)
);

INVx5_ASAP7_75t_L g75 ( 
.A(n_51),
.Y(n_75)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_23),
.Y(n_52)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_52),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g53 ( 
.A(n_24),
.B(n_3),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_53),
.B(n_55),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_24),
.Y(n_54)
);

INVx5_ASAP7_75t_L g79 ( 
.A(n_54),
.Y(n_79)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_25),
.Y(n_55)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_25),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_56),
.B(n_16),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_L g58 ( 
.A1(n_38),
.A2(n_27),
.B1(n_26),
.B2(n_30),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_L g106 ( 
.A1(n_58),
.A2(n_64),
.B1(n_90),
.B2(n_75),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_L g64 ( 
.A1(n_32),
.A2(n_27),
.B1(n_26),
.B2(n_15),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_39),
.A2(n_21),
.B1(n_20),
.B2(n_19),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_66),
.A2(n_68),
.B1(n_74),
.B2(n_88),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_53),
.A2(n_21),
.B1(n_20),
.B2(n_19),
.Y(n_68)
);

CKINVDCx14_ASAP7_75t_R g101 ( 
.A(n_72),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_43),
.A2(n_16),
.B1(n_5),
.B2(n_7),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_77),
.B(n_83),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_51),
.B(n_50),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_80),
.B(n_86),
.Y(n_99)
);

NOR2x1_ASAP7_75t_L g83 ( 
.A(n_54),
.B(n_4),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_84),
.B(n_10),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_55),
.B(n_11),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_35),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_88)
);

OAI22xp33_ASAP7_75t_L g90 ( 
.A1(n_33),
.A2(n_10),
.B1(n_34),
.B2(n_56),
.Y(n_90)
);

MAJx2_ASAP7_75t_L g92 ( 
.A(n_85),
.B(n_60),
.C(n_81),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_92),
.B(n_105),
.Y(n_123)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_81),
.Y(n_93)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_93),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_79),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_94),
.B(n_98),
.Y(n_127)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_70),
.B(n_31),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_95),
.Y(n_119)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_62),
.Y(n_96)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_96),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_76),
.A2(n_40),
.B1(n_48),
.B2(n_73),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_100),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_59),
.B(n_48),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_102),
.B(n_106),
.Y(n_129)
);

BUFx8_ASAP7_75t_L g103 ( 
.A(n_76),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_103),
.Y(n_132)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_62),
.Y(n_104)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_104),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_73),
.A2(n_67),
.B1(n_89),
.B2(n_87),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_78),
.B(n_75),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_107),
.B(n_108),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_61),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_71),
.Y(n_109)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_109),
.Y(n_117)
);

A2O1A1Ixp33_ASAP7_75t_L g110 ( 
.A1(n_83),
.A2(n_58),
.B(n_64),
.C(n_66),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_110),
.B(n_61),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_87),
.B(n_63),
.C(n_71),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g130 ( 
.A(n_111),
.B(n_113),
.Y(n_130)
);

AO22x1_ASAP7_75t_SL g112 ( 
.A1(n_65),
.A2(n_69),
.B1(n_57),
.B2(n_88),
.Y(n_112)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_112),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_82),
.B(n_65),
.C(n_69),
.Y(n_113)
);

CKINVDCx14_ASAP7_75t_R g137 ( 
.A(n_118),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_92),
.B(n_57),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_120),
.B(n_124),
.Y(n_135)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_93),
.Y(n_122)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_122),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_99),
.B(n_82),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_101),
.B(n_91),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_125),
.B(n_111),
.Y(n_145)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_95),
.Y(n_126)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_126),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g134 ( 
.A(n_125),
.B(n_98),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_134),
.B(n_144),
.Y(n_148)
);

BUFx5_ASAP7_75t_L g138 ( 
.A(n_114),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_138),
.B(n_141),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_130),
.B(n_120),
.C(n_118),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_139),
.B(n_140),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_L g140 ( 
.A1(n_123),
.A2(n_110),
.B(n_91),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_131),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_121),
.A2(n_97),
.B1(n_112),
.B2(n_95),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_142),
.A2(n_121),
.B1(n_128),
.B2(n_129),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_114),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_143),
.B(n_94),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_124),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_145),
.B(n_126),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_130),
.B(n_113),
.Y(n_146)
);

XOR2x2_ASAP7_75t_L g147 ( 
.A(n_146),
.B(n_130),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_147),
.B(n_150),
.C(n_139),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_141),
.B(n_127),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_151),
.B(n_152),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_SL g152 ( 
.A(n_135),
.B(n_127),
.Y(n_152)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_154),
.Y(n_159)
);

INVxp67_ASAP7_75t_L g158 ( 
.A(n_155),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_135),
.B(n_117),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_156),
.B(n_133),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_153),
.B(n_145),
.C(n_146),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_160),
.B(n_119),
.C(n_133),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_161),
.B(n_163),
.Y(n_170)
);

AOI221xp5_ASAP7_75t_L g162 ( 
.A1(n_152),
.A2(n_140),
.B1(n_137),
.B2(n_142),
.C(n_136),
.Y(n_162)
);

NOR3xp33_ASAP7_75t_SL g168 ( 
.A(n_162),
.B(n_147),
.C(n_136),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_149),
.B(n_115),
.Y(n_163)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_164),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_161),
.B(n_153),
.Y(n_165)
);

AOI21xp5_ASAP7_75t_L g171 ( 
.A1(n_165),
.A2(n_166),
.B(n_169),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_158),
.A2(n_148),
.B1(n_155),
.B2(n_129),
.Y(n_166)
);

A2O1A1Ixp33_ASAP7_75t_SL g174 ( 
.A1(n_168),
.A2(n_103),
.B(n_112),
.C(n_116),
.Y(n_174)
);

AOI21xp5_ASAP7_75t_L g172 ( 
.A1(n_169),
.A2(n_159),
.B(n_158),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_172),
.A2(n_132),
.B1(n_116),
.B2(n_108),
.Y(n_176)
);

A2O1A1Ixp33_ASAP7_75t_L g173 ( 
.A1(n_168),
.A2(n_157),
.B(n_143),
.C(n_117),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_R g177 ( 
.A(n_173),
.B(n_174),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_171),
.A2(n_167),
.B1(n_165),
.B2(n_170),
.Y(n_175)
);

AO21x1_ASAP7_75t_L g179 ( 
.A1(n_175),
.A2(n_103),
.B(n_115),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_SL g178 ( 
.A(n_176),
.B(n_132),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_178),
.B(n_179),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_SL g181 ( 
.A1(n_179),
.A2(n_175),
.B(n_177),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_L g182 ( 
.A1(n_181),
.A2(n_122),
.B(n_109),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_182),
.B(n_180),
.C(n_104),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_183),
.B(n_138),
.Y(n_184)
);


endmodule