module real_jpeg_15645_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_247;
wire n_146;
wire n_78;
wire n_83;
wire n_286;
wire n_166;
wire n_176;
wire n_221;
wire n_292;
wire n_215;
wire n_249;
wire n_288;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_280;
wire n_64;
wire n_177;
wire n_291;
wire n_236;
wire n_47;
wire n_131;
wire n_271;
wire n_281;
wire n_163;
wire n_276;
wire n_22;
wire n_287;
wire n_237;
wire n_174;
wire n_87;
wire n_197;
wire n_173;
wire n_40;
wire n_243;
wire n_105;
wire n_255;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_164;
wire n_48;
wire n_200;
wire n_275;
wire n_293;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_155;
wire n_120;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_238;
wire n_67;
wire n_79;
wire n_178;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_239;
wire n_162;
wire n_290;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_285;
wire n_172;
wire n_45;
wire n_211;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_262;
wire n_222;
wire n_148;
wire n_118;
wire n_220;
wire n_294;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_298;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_296;
wire n_134;
wire n_270;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_203;
wire n_192;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_205;
wire n_258;
wire n_289;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_228;
wire n_20;
wire n_150;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_259;
wire n_103;
wire n_225;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_284;
wire n_226;
wire n_277;
wire n_125;
wire n_297;
wire n_185;
wire n_209;
wire n_55;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_240;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_279;
wire n_167;
wire n_295;
wire n_213;
wire n_179;
wire n_128;
wire n_202;
wire n_133;
wire n_216;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_206;
wire n_127;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_181;
wire n_85;
wire n_283;
wire n_101;
wire n_274;
wire n_256;
wire n_182;
wire n_253;
wire n_96;
wire n_269;
wire n_273;
wire n_89;

AND2x2_ASAP7_75t_L g41 ( 
.A(n_0),
.B(n_42),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_0),
.A2(n_5),
.B1(n_54),
.B2(n_58),
.Y(n_53)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_0),
.B(n_87),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_0),
.B(n_99),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_0),
.B(n_164),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_0),
.B(n_199),
.Y(n_198)
);

AND2x2_ASAP7_75t_L g205 ( 
.A(n_0),
.B(n_206),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_0),
.B(n_248),
.Y(n_247)
);

AND2x2_ASAP7_75t_L g28 ( 
.A(n_1),
.B(n_29),
.Y(n_28)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_1),
.B(n_68),
.Y(n_67)
);

CKINVDCx16_ASAP7_75t_R g115 ( 
.A(n_1),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_1),
.B(n_99),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_2),
.Y(n_90)
);

BUFx3_ASAP7_75t_L g123 ( 
.A(n_2),
.Y(n_123)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_2),
.Y(n_197)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_3),
.Y(n_70)
);

BUFx5_ASAP7_75t_L g84 ( 
.A(n_3),
.Y(n_84)
);

BUFx5_ASAP7_75t_L g175 ( 
.A(n_3),
.Y(n_175)
);

BUFx6f_ASAP7_75t_L g202 ( 
.A(n_3),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g230 ( 
.A(n_3),
.Y(n_230)
);

AND2x2_ASAP7_75t_L g148 ( 
.A(n_4),
.B(n_149),
.Y(n_148)
);

CKINVDCx16_ASAP7_75t_R g49 ( 
.A(n_5),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g146 ( 
.A(n_5),
.B(n_147),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_6),
.B(n_36),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_6),
.B(n_63),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_6),
.B(n_95),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_6),
.B(n_193),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_6),
.B(n_239),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_6),
.B(n_253),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_6),
.B(n_262),
.Y(n_261)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_7),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g151 ( 
.A(n_7),
.Y(n_151)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_8),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_8),
.Y(n_100)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_8),
.Y(n_242)
);

AND2x2_ASAP7_75t_L g24 ( 
.A(n_9),
.B(n_25),
.Y(n_24)
);

AND2x2_ASAP7_75t_SL g31 ( 
.A(n_9),
.B(n_32),
.Y(n_31)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_9),
.B(n_72),
.Y(n_71)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_9),
.B(n_84),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g102 ( 
.A(n_9),
.B(n_103),
.Y(n_102)
);

CKINVDCx16_ASAP7_75t_R g126 ( 
.A(n_9),
.Y(n_126)
);

NAND2x1_ASAP7_75t_L g142 ( 
.A(n_9),
.B(n_143),
.Y(n_142)
);

AND2x2_ASAP7_75t_L g214 ( 
.A(n_9),
.B(n_149),
.Y(n_214)
);

AND2x2_ASAP7_75t_SL g106 ( 
.A(n_10),
.B(n_107),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g129 ( 
.A(n_10),
.B(n_130),
.Y(n_129)
);

AND2x2_ASAP7_75t_L g172 ( 
.A(n_10),
.B(n_173),
.Y(n_172)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_11),
.B(n_79),
.Y(n_78)
);

AND2x2_ASAP7_75t_L g121 ( 
.A(n_11),
.B(n_122),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_11),
.B(n_171),
.Y(n_170)
);

AND2x2_ASAP7_75t_L g208 ( 
.A(n_11),
.B(n_209),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_11),
.B(n_213),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_11),
.B(n_228),
.Y(n_227)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_12),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_12),
.Y(n_128)
);

INVx6_ASAP7_75t_L g166 ( 
.A(n_12),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_13),
.Y(n_47)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

BUFx4f_ASAP7_75t_L g114 ( 
.A(n_14),
.Y(n_114)
);

BUFx12f_ASAP7_75t_L g132 ( 
.A(n_14),
.Y(n_132)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_15),
.Y(n_65)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

OAI22xp5_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_181),
.B1(n_297),
.B2(n_298),
.Y(n_17)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_18),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_179),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_135),
.Y(n_19)
);

NOR2xp67_ASAP7_75t_SL g180 ( 
.A(n_20),
.B(n_135),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_75),
.C(n_116),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_21),
.B(n_295),
.Y(n_294)
);

XOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_39),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_22),
.B(n_40),
.C(n_61),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_31),
.C(n_34),
.Y(n_22)
);

XNOR2xp5_ASAP7_75t_SL g284 ( 
.A(n_23),
.B(n_285),
.Y(n_284)
);

AND2x2_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_28),
.Y(n_23)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_24),
.B(n_28),
.Y(n_226)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_24),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_24),
.A2(n_246),
.B1(n_247),
.B2(n_259),
.Y(n_258)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g266 ( 
.A(n_27),
.Y(n_266)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_30),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_31),
.A2(n_34),
.B1(n_35),
.B2(n_286),
.Y(n_285)
);

INVx2_ASAP7_75t_SL g286 ( 
.A(n_31),
.Y(n_286)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_33),
.Y(n_60)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

XNOR2xp5_ASAP7_75t_L g39 ( 
.A(n_40),
.B(n_61),
.Y(n_39)
);

AOI21xp5_ASAP7_75t_L g40 ( 
.A1(n_41),
.A2(n_48),
.B(n_53),
.Y(n_40)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_47),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_49),
.B(n_50),
.Y(n_48)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_53),
.A2(n_153),
.B1(n_154),
.B2(n_155),
.Y(n_152)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_53),
.Y(n_155)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_57),
.Y(n_109)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx2_ASAP7_75t_SL g59 ( 
.A(n_60),
.Y(n_59)
);

XOR2xp5_ASAP7_75t_L g61 ( 
.A(n_62),
.B(n_66),
.Y(n_61)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_62),
.B(n_67),
.C(n_71),
.Y(n_178)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_65),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g66 ( 
.A(n_67),
.B(n_71),
.Y(n_66)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_70),
.Y(n_257)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_71),
.Y(n_190)
);

HB1xp67_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_74),
.Y(n_81)
);

HB1xp67_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_76),
.B(n_116),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_77),
.B(n_92),
.C(n_104),
.Y(n_76)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_77),
.B(n_280),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_82),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_78),
.B(n_83),
.C(n_86),
.Y(n_118)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx5_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_83),
.A2(n_85),
.B1(n_86),
.B2(n_91),
.Y(n_82)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_83),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_83),
.A2(n_91),
.B1(n_237),
.B2(n_238),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_83),
.B(n_237),
.C(n_243),
.Y(n_273)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx8_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx6_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

BUFx5_ASAP7_75t_L g103 ( 
.A(n_90),
.Y(n_103)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_93),
.B(n_105),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_98),
.C(n_101),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_94),
.A2(n_101),
.B1(n_102),
.B2(n_222),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_94),
.Y(n_222)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g171 ( 
.A(n_97),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_98),
.B(n_221),
.Y(n_220)
);

BUFx12f_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_101),
.A2(n_102),
.B1(n_163),
.B2(n_167),
.Y(n_162)
);

INVx2_ASAP7_75t_SL g101 ( 
.A(n_102),
.Y(n_101)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

XOR2xp5_ASAP7_75t_L g105 ( 
.A(n_106),
.B(n_110),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_106),
.B(n_110),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_108),
.Y(n_210)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_111),
.B(n_115),
.Y(n_110)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g207 ( 
.A(n_114),
.Y(n_207)
);

XNOR2x1_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_120),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_L g117 ( 
.A(n_118),
.B(n_119),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_118),
.B(n_119),
.C(n_158),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_120),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_124),
.Y(n_120)
);

MAJx2_ASAP7_75t_L g154 ( 
.A(n_121),
.B(n_129),
.C(n_134),
.Y(n_154)
);

BUFx3_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_125),
.A2(n_129),
.B1(n_133),
.B2(n_134),
.Y(n_124)
);

INVx1_ASAP7_75t_SL g134 ( 
.A(n_125),
.Y(n_134)
);

OR2x2_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_127),
.Y(n_125)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_129),
.Y(n_133)
);

INVx4_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g147 ( 
.A(n_132),
.Y(n_147)
);

BUFx3_ASAP7_75t_L g213 ( 
.A(n_132),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_156),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_138),
.Y(n_136)
);

XNOR2x2_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_152),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_145),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

INVx8_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_148),
.Y(n_145)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

INVx3_ASAP7_75t_L g249 ( 
.A(n_151),
.Y(n_249)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_SL g156 ( 
.A(n_157),
.B(n_159),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_168),
.Y(n_159)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_162),
.Y(n_160)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_163),
.Y(n_167)
);

HB1xp67_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_178),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_170),
.A2(n_172),
.B1(n_176),
.B2(n_177),
.Y(n_169)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_170),
.Y(n_177)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_172),
.Y(n_176)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVxp33_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_181),
.Y(n_298)
);

HB1xp67_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_SL g182 ( 
.A1(n_183),
.A2(n_292),
.B(n_296),
.Y(n_182)
);

AOI21xp5_ASAP7_75t_L g183 ( 
.A1(n_184),
.A2(n_276),
.B(n_291),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_SL g184 ( 
.A1(n_185),
.A2(n_231),
.B(n_275),
.Y(n_184)
);

AND2x2_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_217),
.Y(n_185)
);

OR2x2_ASAP7_75t_L g275 ( 
.A(n_186),
.B(n_217),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_203),
.C(n_211),
.Y(n_186)
);

HB1xp67_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_188),
.B(n_271),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_191),
.Y(n_188)
);

INVx1_ASAP7_75t_SL g189 ( 
.A(n_190),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_190),
.B(n_192),
.C(n_198),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_198),
.Y(n_191)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

BUFx6f_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

HB1xp67_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_203),
.A2(n_204),
.B1(n_211),
.B2(n_272),
.Y(n_271)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_208),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_SL g244 ( 
.A(n_205),
.B(n_208),
.Y(n_244)
);

BUFx2_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_211),
.Y(n_272)
);

AO22x1_ASAP7_75t_SL g211 ( 
.A1(n_212),
.A2(n_214),
.B1(n_215),
.B2(n_216),
.Y(n_211)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_212),
.Y(n_215)
);

INVx1_ASAP7_75t_SL g216 ( 
.A(n_214),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_214),
.B(n_215),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_216),
.B(n_261),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_223),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_220),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_219),
.B(n_223),
.C(n_290),
.Y(n_289)
);

HB1xp67_ASAP7_75t_L g290 ( 
.A(n_220),
.Y(n_290)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_225),
.Y(n_223)
);

MAJx2_ASAP7_75t_L g288 ( 
.A(n_224),
.B(n_226),
.C(n_227),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_227),
.Y(n_225)
);

INVx4_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

INVx6_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

AOI21xp5_ASAP7_75t_L g231 ( 
.A1(n_232),
.A2(n_269),
.B(n_274),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_SL g232 ( 
.A1(n_233),
.A2(n_250),
.B(n_268),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_245),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_234),
.B(n_245),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_235),
.A2(n_236),
.B1(n_243),
.B2(n_244),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

INVx3_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_SL g245 ( 
.A(n_246),
.B(n_247),
.Y(n_245)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_247),
.Y(n_259)
);

INVx5_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

AOI21x1_ASAP7_75t_SL g250 ( 
.A1(n_251),
.A2(n_260),
.B(n_267),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_258),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_252),
.B(n_258),
.Y(n_267)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

HB1xp67_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

INVx3_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g269 ( 
.A(n_270),
.B(n_273),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_270),
.B(n_273),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_277),
.B(n_289),
.Y(n_276)
);

NOR2xp67_ASAP7_75t_L g291 ( 
.A(n_277),
.B(n_289),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_278),
.A2(n_279),
.B1(n_281),
.B2(n_282),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_278),
.B(n_283),
.C(n_288),
.Y(n_293)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_283),
.A2(n_284),
.B1(n_287),
.B2(n_288),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_293),
.B(n_294),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_293),
.B(n_294),
.Y(n_296)
);


endmodule