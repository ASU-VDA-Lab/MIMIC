module fake_jpeg_31281_n_552 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_552);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_552;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx12_ASAP7_75t_L g18 ( 
.A(n_15),
.Y(n_18)
);

INVx2_ASAP7_75t_SL g19 ( 
.A(n_5),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_10),
.Y(n_20)
);

CKINVDCx14_ASAP7_75t_R g21 ( 
.A(n_10),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_14),
.Y(n_23)
);

INVx6_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_10),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_16),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_16),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_0),
.Y(n_30)
);

BUFx10_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

BUFx8_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_14),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_11),
.Y(n_35)
);

CKINVDCx11_ASAP7_75t_R g36 ( 
.A(n_15),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_9),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_11),
.Y(n_38)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_11),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_4),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_17),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_8),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_12),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_4),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_4),
.Y(n_45)
);

INVx13_ASAP7_75t_L g46 ( 
.A(n_16),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_16),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_17),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_1),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_17),
.Y(n_50)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_13),
.Y(n_51)
);

INVxp67_ASAP7_75t_L g52 ( 
.A(n_17),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_28),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_53),
.Y(n_118)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_29),
.Y(n_54)
);

INVx4_ASAP7_75t_L g128 ( 
.A(n_54),
.Y(n_128)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_32),
.Y(n_55)
);

INVx8_ASAP7_75t_L g131 ( 
.A(n_55),
.Y(n_131)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_22),
.Y(n_56)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_56),
.Y(n_117)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_29),
.Y(n_57)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_57),
.Y(n_122)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_46),
.Y(n_58)
);

BUFx5_ASAP7_75t_L g110 ( 
.A(n_58),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_52),
.B(n_7),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_59),
.B(n_72),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_28),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_60),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_28),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_61),
.Y(n_126)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_22),
.Y(n_62)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_62),
.Y(n_149)
);

INVx11_ASAP7_75t_L g63 ( 
.A(n_28),
.Y(n_63)
);

INVx6_ASAP7_75t_L g123 ( 
.A(n_63),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_34),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_64),
.Y(n_137)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_32),
.Y(n_65)
);

INVx8_ASAP7_75t_L g134 ( 
.A(n_65),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_20),
.B(n_7),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_66),
.B(n_102),
.Y(n_113)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_46),
.Y(n_67)
);

INVx5_ASAP7_75t_L g125 ( 
.A(n_67),
.Y(n_125)
);

INVx13_ASAP7_75t_L g68 ( 
.A(n_36),
.Y(n_68)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_68),
.Y(n_133)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_34),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_69),
.Y(n_153)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_29),
.Y(n_70)
);

INVx3_ASAP7_75t_L g151 ( 
.A(n_70),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_34),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_71),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_20),
.B(n_7),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_34),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_73),
.Y(n_166)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_22),
.Y(n_74)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_74),
.Y(n_111)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_44),
.Y(n_75)
);

INVx6_ASAP7_75t_L g145 ( 
.A(n_75),
.Y(n_145)
);

HAxp5_ASAP7_75t_SL g76 ( 
.A(n_36),
.B(n_7),
.CON(n_76),
.SN(n_76)
);

OR2x2_ASAP7_75t_L g127 ( 
.A(n_76),
.B(n_93),
.Y(n_127)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_39),
.Y(n_77)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_77),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_44),
.Y(n_78)
);

INVx6_ASAP7_75t_L g172 ( 
.A(n_78),
.Y(n_172)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_35),
.Y(n_79)
);

INVx3_ASAP7_75t_L g155 ( 
.A(n_79),
.Y(n_155)
);

INVx8_ASAP7_75t_L g80 ( 
.A(n_32),
.Y(n_80)
);

INVx3_ASAP7_75t_L g175 ( 
.A(n_80),
.Y(n_175)
);

INVx11_ASAP7_75t_L g81 ( 
.A(n_44),
.Y(n_81)
);

BUFx3_ASAP7_75t_L g143 ( 
.A(n_81),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_44),
.Y(n_82)
);

BUFx2_ASAP7_75t_L g114 ( 
.A(n_82),
.Y(n_114)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_39),
.Y(n_83)
);

INVx4_ASAP7_75t_L g141 ( 
.A(n_83),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_23),
.B(n_6),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_84),
.B(n_87),
.Y(n_142)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_35),
.Y(n_85)
);

INVx4_ASAP7_75t_L g174 ( 
.A(n_85),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_51),
.A2(n_6),
.B1(n_1),
.B2(n_2),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_86),
.A2(n_106),
.B1(n_19),
.B2(n_48),
.Y(n_130)
);

AND2x2_ASAP7_75t_SL g87 ( 
.A(n_39),
.B(n_6),
.Y(n_87)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_42),
.Y(n_88)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_88),
.Y(n_156)
);

BUFx5_ASAP7_75t_L g89 ( 
.A(n_38),
.Y(n_89)
);

BUFx2_ASAP7_75t_L g119 ( 
.A(n_89),
.Y(n_119)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_35),
.Y(n_90)
);

INVx4_ASAP7_75t_L g152 ( 
.A(n_90),
.Y(n_152)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_24),
.Y(n_91)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_91),
.Y(n_115)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_45),
.Y(n_92)
);

INVx4_ASAP7_75t_L g157 ( 
.A(n_92),
.Y(n_157)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_32),
.B(n_8),
.Y(n_93)
);

BUFx4f_ASAP7_75t_L g94 ( 
.A(n_32),
.Y(n_94)
);

BUFx2_ASAP7_75t_L g170 ( 
.A(n_94),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_50),
.Y(n_95)
);

INVx4_ASAP7_75t_L g158 ( 
.A(n_95),
.Y(n_158)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_24),
.Y(n_96)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_96),
.Y(n_116)
);

BUFx2_ASAP7_75t_L g97 ( 
.A(n_50),
.Y(n_97)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_97),
.Y(n_129)
);

BUFx2_ASAP7_75t_L g98 ( 
.A(n_50),
.Y(n_98)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_98),
.Y(n_136)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_45),
.Y(n_99)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_99),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_50),
.Y(n_100)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_100),
.Y(n_148)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_45),
.Y(n_101)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_101),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_23),
.B(n_8),
.Y(n_102)
);

BUFx5_ASAP7_75t_L g103 ( 
.A(n_38),
.Y(n_103)
);

CKINVDCx16_ASAP7_75t_R g144 ( 
.A(n_103),
.Y(n_144)
);

BUFx5_ASAP7_75t_L g104 ( 
.A(n_38),
.Y(n_104)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_104),
.Y(n_167)
);

BUFx5_ASAP7_75t_L g105 ( 
.A(n_38),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_105),
.B(n_107),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_L g106 ( 
.A1(n_21),
.A2(n_5),
.B1(n_1),
.B2(n_2),
.Y(n_106)
);

BUFx12_ASAP7_75t_L g107 ( 
.A(n_46),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_107),
.B(n_109),
.Y(n_160)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_24),
.Y(n_108)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_108),
.Y(n_162)
);

BUFx3_ASAP7_75t_L g109 ( 
.A(n_51),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_97),
.A2(n_21),
.B1(n_19),
.B2(n_51),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_120),
.A2(n_124),
.B1(n_132),
.B2(n_135),
.Y(n_186)
);

AOI22xp33_ASAP7_75t_L g124 ( 
.A1(n_69),
.A2(n_38),
.B1(n_48),
.B2(n_47),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_130),
.A2(n_138),
.B1(n_82),
.B2(n_78),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_87),
.A2(n_25),
.B1(n_43),
.B2(n_41),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_98),
.A2(n_19),
.B1(n_48),
.B2(n_47),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_53),
.A2(n_25),
.B1(n_43),
.B2(n_41),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_SL g146 ( 
.A(n_76),
.B(n_49),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_146),
.B(n_18),
.Y(n_203)
);

AOI22xp33_ASAP7_75t_L g147 ( 
.A1(n_75),
.A2(n_27),
.B1(n_26),
.B2(n_47),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g232 ( 
.A1(n_147),
.A2(n_159),
.B1(n_169),
.B2(n_171),
.Y(n_232)
);

AOI22xp33_ASAP7_75t_SL g159 ( 
.A1(n_55),
.A2(n_19),
.B1(n_26),
.B2(n_27),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_68),
.B(n_49),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_161),
.B(n_163),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_93),
.B(n_40),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_107),
.B(n_40),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_164),
.B(n_168),
.Y(n_178)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_83),
.Y(n_165)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_165),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_58),
.B(n_37),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_SL g169 ( 
.A1(n_65),
.A2(n_27),
.B1(n_26),
.B2(n_42),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_L g171 ( 
.A1(n_60),
.A2(n_30),
.B1(n_33),
.B2(n_37),
.Y(n_171)
);

INVxp67_ASAP7_75t_L g184 ( 
.A(n_173),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_127),
.A2(n_33),
.B1(n_30),
.B2(n_106),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g247 ( 
.A(n_176),
.Y(n_247)
);

INVx3_ASAP7_75t_L g179 ( 
.A(n_110),
.Y(n_179)
);

BUFx2_ASAP7_75t_L g253 ( 
.A(n_179),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_113),
.B(n_31),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_180),
.B(n_199),
.Y(n_242)
);

INVx3_ASAP7_75t_L g181 ( 
.A(n_143),
.Y(n_181)
);

INVx4_ASAP7_75t_L g239 ( 
.A(n_181),
.Y(n_239)
);

INVx4_ASAP7_75t_L g182 ( 
.A(n_152),
.Y(n_182)
);

INVx4_ASAP7_75t_L g246 ( 
.A(n_182),
.Y(n_246)
);

AOI22xp33_ASAP7_75t_SL g185 ( 
.A1(n_119),
.A2(n_54),
.B1(n_90),
.B2(n_58),
.Y(n_185)
);

AOI22xp33_ASAP7_75t_SL g270 ( 
.A1(n_185),
.A2(n_223),
.B1(n_227),
.B2(n_228),
.Y(n_270)
);

INVxp67_ASAP7_75t_L g187 ( 
.A(n_160),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_187),
.B(n_203),
.Y(n_250)
);

INVx6_ASAP7_75t_L g188 ( 
.A(n_118),
.Y(n_188)
);

INVx8_ASAP7_75t_L g280 ( 
.A(n_188),
.Y(n_280)
);

AND2x2_ASAP7_75t_L g189 ( 
.A(n_142),
.B(n_67),
.Y(n_189)
);

FAx1_ASAP7_75t_SL g282 ( 
.A(n_189),
.B(n_204),
.CI(n_218),
.CON(n_282),
.SN(n_282)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_111),
.Y(n_190)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_190),
.Y(n_257)
);

OAI22xp33_ASAP7_75t_SL g191 ( 
.A1(n_145),
.A2(n_108),
.B1(n_61),
.B2(n_100),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_191),
.A2(n_212),
.B1(n_157),
.B2(n_154),
.Y(n_268)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_115),
.Y(n_192)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_192),
.Y(n_262)
);

HB1xp67_ASAP7_75t_L g193 ( 
.A(n_152),
.Y(n_193)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_193),
.Y(n_255)
);

INVx4_ASAP7_75t_L g194 ( 
.A(n_128),
.Y(n_194)
);

INVx3_ASAP7_75t_L g240 ( 
.A(n_194),
.Y(n_240)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_156),
.Y(n_195)
);

CKINVDCx16_ASAP7_75t_R g272 ( 
.A(n_195),
.Y(n_272)
);

INVx3_ASAP7_75t_L g196 ( 
.A(n_143),
.Y(n_196)
);

INVx3_ASAP7_75t_L g241 ( 
.A(n_196),
.Y(n_241)
);

BUFx3_ASAP7_75t_L g197 ( 
.A(n_167),
.Y(n_197)
);

BUFx3_ASAP7_75t_L g248 ( 
.A(n_197),
.Y(n_248)
);

INVx6_ASAP7_75t_L g198 ( 
.A(n_118),
.Y(n_198)
);

INVx5_ASAP7_75t_L g254 ( 
.A(n_198),
.Y(n_254)
);

INVx6_ASAP7_75t_SL g199 ( 
.A(n_133),
.Y(n_199)
);

INVx6_ASAP7_75t_L g200 ( 
.A(n_121),
.Y(n_200)
);

INVx5_ASAP7_75t_L g259 ( 
.A(n_200),
.Y(n_259)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_117),
.Y(n_201)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_201),
.Y(n_271)
);

BUFx6f_ASAP7_75t_L g202 ( 
.A(n_121),
.Y(n_202)
);

INVx11_ASAP7_75t_L g275 ( 
.A(n_202),
.Y(n_275)
);

AND2x2_ASAP7_75t_L g204 ( 
.A(n_139),
.B(n_94),
.Y(n_204)
);

INVx3_ASAP7_75t_L g205 ( 
.A(n_125),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_205),
.B(n_206),
.Y(n_260)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_149),
.Y(n_206)
);

INVx6_ASAP7_75t_L g207 ( 
.A(n_126),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_207),
.B(n_208),
.Y(n_264)
);

INVx5_ASAP7_75t_L g208 ( 
.A(n_131),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_127),
.B(n_18),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_209),
.B(n_211),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_112),
.B(n_31),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_210),
.B(n_213),
.Y(n_263)
);

INVx3_ASAP7_75t_L g211 ( 
.A(n_123),
.Y(n_211)
);

OA22x2_ASAP7_75t_L g212 ( 
.A1(n_120),
.A2(n_80),
.B1(n_109),
.B2(n_31),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_116),
.B(n_31),
.Y(n_213)
);

INVx3_ASAP7_75t_L g214 ( 
.A(n_123),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_214),
.Y(n_251)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_162),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g284 ( 
.A(n_215),
.B(n_216),
.Y(n_284)
);

CKINVDCx16_ASAP7_75t_R g216 ( 
.A(n_159),
.Y(n_216)
);

CKINVDCx16_ASAP7_75t_R g217 ( 
.A(n_135),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_217),
.Y(n_276)
);

AND2x4_ASAP7_75t_L g218 ( 
.A(n_169),
.B(n_31),
.Y(n_218)
);

AND2x2_ASAP7_75t_L g219 ( 
.A(n_141),
.B(n_95),
.Y(n_219)
);

MAJx2_ASAP7_75t_L g285 ( 
.A(n_219),
.B(n_12),
.C(n_14),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_140),
.B(n_150),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_220),
.B(n_225),
.Y(n_243)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_129),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_221),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_L g258 ( 
.A1(n_222),
.A2(n_235),
.B1(n_137),
.B2(n_166),
.Y(n_258)
);

INVx5_ASAP7_75t_L g223 ( 
.A(n_131),
.Y(n_223)
);

HB1xp67_ASAP7_75t_L g224 ( 
.A(n_122),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_224),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_171),
.B(n_18),
.Y(n_225)
);

A2O1A1Ixp33_ASAP7_75t_L g226 ( 
.A1(n_147),
.A2(n_31),
.B(n_1),
.C(n_2),
.Y(n_226)
);

A2O1A1Ixp33_ASAP7_75t_L g278 ( 
.A1(n_226),
.A2(n_237),
.B(n_12),
.C(n_13),
.Y(n_278)
);

INVx11_ASAP7_75t_L g227 ( 
.A(n_134),
.Y(n_227)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_136),
.Y(n_228)
);

BUFx6f_ASAP7_75t_L g229 ( 
.A(n_126),
.Y(n_229)
);

AOI22xp33_ASAP7_75t_L g266 ( 
.A1(n_229),
.A2(n_154),
.B1(n_137),
.B2(n_170),
.Y(n_266)
);

AOI22xp33_ASAP7_75t_SL g230 ( 
.A1(n_119),
.A2(n_73),
.B1(n_71),
.B2(n_64),
.Y(n_230)
);

OAI22x1_ASAP7_75t_L g252 ( 
.A1(n_230),
.A2(n_234),
.B1(n_124),
.B2(n_170),
.Y(n_252)
);

INVxp67_ASAP7_75t_L g231 ( 
.A(n_151),
.Y(n_231)
);

CKINVDCx12_ASAP7_75t_R g267 ( 
.A(n_231),
.Y(n_267)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_148),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_233),
.B(n_158),
.Y(n_244)
);

AOI22xp33_ASAP7_75t_SL g234 ( 
.A1(n_114),
.A2(n_81),
.B1(n_63),
.B2(n_3),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_145),
.A2(n_9),
.B1(n_2),
.B2(n_3),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_174),
.A2(n_18),
.B1(n_3),
.B2(n_4),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_236),
.A2(n_144),
.B1(n_134),
.B2(n_175),
.Y(n_245)
);

AOI32xp33_ASAP7_75t_L g237 ( 
.A1(n_155),
.A2(n_18),
.A3(n_3),
.B1(n_5),
.B2(n_9),
.Y(n_237)
);

OAI22xp33_ASAP7_75t_SL g238 ( 
.A1(n_232),
.A2(n_114),
.B1(n_158),
.B2(n_172),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_L g288 ( 
.A1(n_238),
.A2(n_256),
.B1(n_278),
.B2(n_230),
.Y(n_288)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_244),
.Y(n_286)
);

AND2x2_ASAP7_75t_L g318 ( 
.A(n_245),
.B(n_258),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_218),
.B(n_172),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_249),
.B(n_265),
.Y(n_289)
);

AOI22xp33_ASAP7_75t_SL g310 ( 
.A1(n_252),
.A2(n_179),
.B1(n_188),
.B2(n_214),
.Y(n_310)
);

OAI22xp33_ASAP7_75t_SL g256 ( 
.A1(n_186),
.A2(n_153),
.B1(n_157),
.B2(n_166),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_189),
.B(n_187),
.C(n_204),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_261),
.B(n_274),
.C(n_285),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_218),
.B(n_153),
.Y(n_265)
);

INVxp67_ASAP7_75t_L g322 ( 
.A(n_266),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_268),
.A2(n_279),
.B1(n_234),
.B2(n_185),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_218),
.B(n_0),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_269),
.B(n_273),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_178),
.B(n_0),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_177),
.B(n_0),
.C(n_9),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_191),
.A2(n_15),
.B1(n_12),
.B2(n_13),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_SL g315 ( 
.A(n_285),
.B(n_0),
.Y(n_315)
);

AOI21xp5_ASAP7_75t_L g287 ( 
.A1(n_249),
.A2(n_212),
.B(n_231),
.Y(n_287)
);

AOI21xp5_ASAP7_75t_L g350 ( 
.A1(n_287),
.A2(n_308),
.B(n_325),
.Y(n_350)
);

AOI22xp5_ASAP7_75t_L g339 ( 
.A1(n_288),
.A2(n_294),
.B1(n_305),
.B2(n_259),
.Y(n_339)
);

BUFx5_ASAP7_75t_L g290 ( 
.A(n_248),
.Y(n_290)
);

HB1xp67_ASAP7_75t_L g359 ( 
.A(n_290),
.Y(n_359)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_244),
.Y(n_291)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_291),
.Y(n_333)
);

AOI32xp33_ASAP7_75t_L g293 ( 
.A1(n_247),
.A2(n_184),
.A3(n_212),
.B1(n_226),
.B2(n_194),
.Y(n_293)
);

OAI21xp5_ASAP7_75t_SL g326 ( 
.A1(n_293),
.A2(n_278),
.B(n_270),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_260),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_295),
.B(n_297),
.Y(n_335)
);

XNOR2xp5_ASAP7_75t_SL g349 ( 
.A(n_296),
.B(n_313),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_272),
.B(n_184),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_271),
.Y(n_298)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_298),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_SL g299 ( 
.A(n_250),
.B(n_183),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_SL g346 ( 
.A(n_299),
.B(n_324),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_273),
.B(n_182),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_300),
.B(n_303),
.Y(n_327)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_257),
.Y(n_301)
);

INVx1_ASAP7_75t_SL g345 ( 
.A(n_301),
.Y(n_345)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_271),
.Y(n_302)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_302),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_263),
.B(n_219),
.Y(n_303)
);

CKINVDCx16_ASAP7_75t_R g304 ( 
.A(n_267),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_304),
.B(n_317),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_L g305 ( 
.A1(n_265),
.A2(n_207),
.B1(n_200),
.B2(n_198),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_248),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_306),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_261),
.B(n_197),
.C(n_181),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_307),
.B(n_309),
.C(n_311),
.Y(n_336)
);

O2A1O1Ixp33_ASAP7_75t_SL g308 ( 
.A1(n_252),
.A2(n_227),
.B(n_223),
.C(n_208),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_282),
.B(n_196),
.C(n_205),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_SL g329 ( 
.A1(n_310),
.A2(n_279),
.B1(n_253),
.B2(n_275),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_282),
.B(n_211),
.C(n_229),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_253),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_312),
.Y(n_331)
);

MAJx2_ASAP7_75t_L g313 ( 
.A(n_281),
.B(n_14),
.C(n_202),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_253),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g341 ( 
.A(n_314),
.Y(n_341)
);

XNOR2xp5_ASAP7_75t_L g356 ( 
.A(n_315),
.B(n_296),
.Y(n_356)
);

XOR2xp5_ASAP7_75t_L g316 ( 
.A(n_242),
.B(n_243),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_316),
.B(n_251),
.C(n_262),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_272),
.B(n_274),
.Y(n_317)
);

NOR2x1_ASAP7_75t_L g319 ( 
.A(n_268),
.B(n_247),
.Y(n_319)
);

OAI21xp5_ASAP7_75t_L g330 ( 
.A1(n_319),
.A2(n_251),
.B(n_258),
.Y(n_330)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_255),
.Y(n_320)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_320),
.Y(n_351)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_257),
.Y(n_321)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_321),
.Y(n_355)
);

CKINVDCx16_ASAP7_75t_R g323 ( 
.A(n_284),
.Y(n_323)
);

CKINVDCx16_ASAP7_75t_R g343 ( 
.A(n_323),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_SL g324 ( 
.A(n_243),
.B(n_282),
.Y(n_324)
);

AOI21xp5_ASAP7_75t_L g325 ( 
.A1(n_269),
.A2(n_276),
.B(n_245),
.Y(n_325)
);

AOI21xp5_ASAP7_75t_L g378 ( 
.A1(n_326),
.A2(n_330),
.B(n_353),
.Y(n_378)
);

AOI21x1_ASAP7_75t_L g328 ( 
.A1(n_289),
.A2(n_276),
.B(n_264),
.Y(n_328)
);

OAI21xp5_ASAP7_75t_SL g369 ( 
.A1(n_328),
.A2(n_303),
.B(n_300),
.Y(n_369)
);

AOI22xp5_ASAP7_75t_L g388 ( 
.A1(n_329),
.A2(n_319),
.B1(n_322),
.B2(n_333),
.Y(n_388)
);

OAI21xp33_ASAP7_75t_L g338 ( 
.A1(n_324),
.A2(n_283),
.B(n_239),
.Y(n_338)
);

INVxp67_ASAP7_75t_L g361 ( 
.A(n_338),
.Y(n_361)
);

OAI22xp5_ASAP7_75t_SL g374 ( 
.A1(n_339),
.A2(n_357),
.B1(n_330),
.B2(n_358),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_286),
.B(n_283),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_340),
.B(n_342),
.Y(n_360)
);

AO22x1_ASAP7_75t_SL g342 ( 
.A1(n_286),
.A2(n_262),
.B1(n_255),
.B2(n_259),
.Y(n_342)
);

OAI21xp5_ASAP7_75t_L g347 ( 
.A1(n_325),
.A2(n_277),
.B(n_240),
.Y(n_347)
);

OAI21xp5_ASAP7_75t_L g373 ( 
.A1(n_347),
.A2(n_358),
.B(n_319),
.Y(n_373)
);

XOR2xp5_ASAP7_75t_L g348 ( 
.A(n_316),
.B(n_277),
.Y(n_348)
);

MAJIxp5_ASAP7_75t_L g362 ( 
.A(n_348),
.B(n_307),
.C(n_309),
.Y(n_362)
);

XNOR2xp5_ASAP7_75t_L g363 ( 
.A(n_352),
.B(n_356),
.Y(n_363)
);

OAI21xp5_ASAP7_75t_SL g353 ( 
.A1(n_287),
.A2(n_239),
.B(n_241),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_291),
.B(n_241),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_354),
.B(n_312),
.Y(n_376)
);

AOI22xp5_ASAP7_75t_L g357 ( 
.A1(n_288),
.A2(n_254),
.B1(n_280),
.B2(n_240),
.Y(n_357)
);

OAI21xp5_ASAP7_75t_L g358 ( 
.A1(n_289),
.A2(n_280),
.B(n_254),
.Y(n_358)
);

XNOR2xp5_ASAP7_75t_SL g408 ( 
.A(n_362),
.B(n_356),
.Y(n_408)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_337),
.Y(n_364)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_364),
.Y(n_394)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_337),
.Y(n_365)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_365),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_L g366 ( 
.A(n_334),
.B(n_299),
.Y(n_366)
);

INVxp33_ASAP7_75t_L g399 ( 
.A(n_366),
.Y(n_399)
);

NOR2xp33_ASAP7_75t_L g367 ( 
.A(n_334),
.B(n_295),
.Y(n_367)
);

CKINVDCx20_ASAP7_75t_R g405 ( 
.A(n_367),
.Y(n_405)
);

CKINVDCx16_ASAP7_75t_R g368 ( 
.A(n_335),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_L g423 ( 
.A(n_368),
.B(n_372),
.Y(n_423)
);

INVxp67_ASAP7_75t_L g416 ( 
.A(n_369),
.Y(n_416)
);

BUFx3_ASAP7_75t_L g370 ( 
.A(n_355),
.Y(n_370)
);

BUFx2_ASAP7_75t_L g418 ( 
.A(n_370),
.Y(n_418)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_344),
.Y(n_371)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_371),
.Y(n_401)
);

CKINVDCx20_ASAP7_75t_R g372 ( 
.A(n_340),
.Y(n_372)
);

AOI21xp5_ASAP7_75t_L g414 ( 
.A1(n_373),
.A2(n_385),
.B(n_386),
.Y(n_414)
);

AOI22xp5_ASAP7_75t_L g413 ( 
.A1(n_374),
.A2(n_379),
.B1(n_349),
.B2(n_346),
.Y(n_413)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_344),
.Y(n_375)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_375),
.Y(n_402)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_376),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_SL g377 ( 
.A(n_346),
.B(n_292),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_377),
.B(n_381),
.Y(n_403)
);

OAI22xp5_ASAP7_75t_SL g379 ( 
.A1(n_339),
.A2(n_294),
.B1(n_293),
.B2(n_318),
.Y(n_379)
);

MAJIxp5_ASAP7_75t_L g380 ( 
.A(n_336),
.B(n_311),
.C(n_292),
.Y(n_380)
);

MAJIxp5_ASAP7_75t_L g412 ( 
.A(n_380),
.B(n_336),
.C(n_349),
.Y(n_412)
);

INVxp67_ASAP7_75t_L g381 ( 
.A(n_332),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_351),
.Y(n_382)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_382),
.Y(n_407)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_351),
.Y(n_383)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_383),
.Y(n_421)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_354),
.Y(n_384)
);

CKINVDCx16_ASAP7_75t_R g406 ( 
.A(n_384),
.Y(n_406)
);

OAI21xp5_ASAP7_75t_SL g385 ( 
.A1(n_350),
.A2(n_318),
.B(n_308),
.Y(n_385)
);

OAI21xp5_ASAP7_75t_SL g386 ( 
.A1(n_350),
.A2(n_318),
.B(n_308),
.Y(n_386)
);

AOI21xp5_ASAP7_75t_L g387 ( 
.A1(n_353),
.A2(n_306),
.B(n_305),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_L g410 ( 
.A(n_387),
.B(n_342),
.Y(n_410)
);

OAI22xp5_ASAP7_75t_SL g398 ( 
.A1(n_388),
.A2(n_329),
.B1(n_343),
.B2(n_341),
.Y(n_398)
);

INVxp67_ASAP7_75t_L g389 ( 
.A(n_347),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_389),
.B(n_390),
.Y(n_411)
);

NOR2xp33_ASAP7_75t_L g390 ( 
.A(n_343),
.B(n_323),
.Y(n_390)
);

INVx2_ASAP7_75t_L g391 ( 
.A(n_355),
.Y(n_391)
);

AOI22xp33_ASAP7_75t_L g400 ( 
.A1(n_391),
.A2(n_314),
.B1(n_345),
.B2(n_341),
.Y(n_400)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_342),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_392),
.B(n_331),
.Y(n_417)
);

OAI22xp5_ASAP7_75t_L g393 ( 
.A1(n_392),
.A2(n_357),
.B1(n_333),
.B2(n_327),
.Y(n_393)
);

AOI22xp5_ASAP7_75t_L g436 ( 
.A1(n_393),
.A2(n_397),
.B1(n_398),
.B2(n_422),
.Y(n_436)
);

AO22x1_ASAP7_75t_SL g395 ( 
.A1(n_360),
.A2(n_328),
.B1(n_342),
.B2(n_326),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_395),
.B(n_373),
.Y(n_426)
);

OAI22xp5_ASAP7_75t_L g397 ( 
.A1(n_372),
.A2(n_327),
.B1(n_352),
.B2(n_335),
.Y(n_397)
);

INVxp67_ASAP7_75t_L g447 ( 
.A(n_400),
.Y(n_447)
);

MAJIxp5_ASAP7_75t_L g425 ( 
.A(n_408),
.B(n_412),
.C(n_363),
.Y(n_425)
);

XOR2xp5_ASAP7_75t_L g409 ( 
.A(n_363),
.B(n_348),
.Y(n_409)
);

XNOR2xp5_ASAP7_75t_SL g440 ( 
.A(n_409),
.B(n_378),
.Y(n_440)
);

AOI21xp5_ASAP7_75t_L g437 ( 
.A1(n_410),
.A2(n_361),
.B(n_387),
.Y(n_437)
);

OAI22xp5_ASAP7_75t_SL g435 ( 
.A1(n_413),
.A2(n_380),
.B1(n_362),
.B2(n_388),
.Y(n_435)
);

NOR2xp33_ASAP7_75t_L g415 ( 
.A(n_366),
.B(n_359),
.Y(n_415)
);

NOR2xp33_ASAP7_75t_L g424 ( 
.A(n_415),
.B(n_405),
.Y(n_424)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_417),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_367),
.B(n_331),
.Y(n_419)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_419),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_368),
.B(n_302),
.Y(n_420)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_420),
.Y(n_434)
);

OAI22xp5_ASAP7_75t_L g422 ( 
.A1(n_360),
.A2(n_298),
.B1(n_345),
.B2(n_320),
.Y(n_422)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_424),
.Y(n_452)
);

XOR2xp5_ASAP7_75t_L g454 ( 
.A(n_425),
.B(n_435),
.Y(n_454)
);

OAI22xp5_ASAP7_75t_SL g459 ( 
.A1(n_426),
.A2(n_404),
.B1(n_395),
.B2(n_406),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_405),
.B(n_376),
.Y(n_427)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_427),
.Y(n_453)
);

MAJIxp5_ASAP7_75t_L g428 ( 
.A(n_408),
.B(n_380),
.C(n_362),
.Y(n_428)
);

MAJIxp5_ASAP7_75t_L g457 ( 
.A(n_428),
.B(n_443),
.C(n_413),
.Y(n_457)
);

NOR2xp33_ASAP7_75t_SL g430 ( 
.A(n_399),
.B(n_390),
.Y(n_430)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_430),
.Y(n_474)
);

A2O1A1Ixp33_ASAP7_75t_L g432 ( 
.A1(n_417),
.A2(n_385),
.B(n_386),
.C(n_369),
.Y(n_432)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_432),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_419),
.B(n_384),
.Y(n_433)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_433),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_437),
.B(n_438),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_423),
.B(n_377),
.Y(n_438)
);

CKINVDCx16_ASAP7_75t_R g439 ( 
.A(n_420),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_439),
.B(n_441),
.Y(n_471)
);

XOR2xp5_ASAP7_75t_L g463 ( 
.A(n_440),
.B(n_448),
.Y(n_463)
);

CKINVDCx16_ASAP7_75t_R g441 ( 
.A(n_411),
.Y(n_441)
);

OAI21xp5_ASAP7_75t_L g442 ( 
.A1(n_414),
.A2(n_378),
.B(n_374),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_442),
.B(n_444),
.Y(n_473)
);

MAJIxp5_ASAP7_75t_L g443 ( 
.A(n_412),
.B(n_379),
.C(n_383),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_423),
.B(n_364),
.Y(n_444)
);

OAI21xp5_ASAP7_75t_L g445 ( 
.A1(n_414),
.A2(n_382),
.B(n_375),
.Y(n_445)
);

FAx1_ASAP7_75t_SL g469 ( 
.A(n_445),
.B(n_394),
.CI(n_407),
.CON(n_469),
.SN(n_469)
);

NOR2xp33_ASAP7_75t_L g446 ( 
.A(n_411),
.B(n_371),
.Y(n_446)
);

NOR2xp33_ASAP7_75t_SL g461 ( 
.A(n_446),
.B(n_449),
.Y(n_461)
);

AOI21xp5_ASAP7_75t_L g448 ( 
.A1(n_416),
.A2(n_365),
.B(n_391),
.Y(n_448)
);

CKINVDCx20_ASAP7_75t_R g449 ( 
.A(n_418),
.Y(n_449)
);

NOR2xp33_ASAP7_75t_SL g450 ( 
.A(n_403),
.B(n_313),
.Y(n_450)
);

MAJIxp5_ASAP7_75t_SL g456 ( 
.A(n_450),
.B(n_313),
.C(n_397),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_SL g451 ( 
.A(n_403),
.B(n_315),
.Y(n_451)
);

XNOR2xp5_ASAP7_75t_L g455 ( 
.A(n_451),
.B(n_409),
.Y(n_455)
);

XNOR2xp5_ASAP7_75t_L g481 ( 
.A(n_455),
.B(n_457),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_SL g480 ( 
.A(n_456),
.B(n_450),
.Y(n_480)
);

XNOR2xp5_ASAP7_75t_L g458 ( 
.A(n_443),
.B(n_393),
.Y(n_458)
);

XNOR2xp5_ASAP7_75t_L g482 ( 
.A(n_458),
.B(n_468),
.Y(n_482)
);

XOR2xp5_ASAP7_75t_L g488 ( 
.A(n_459),
.B(n_445),
.Y(n_488)
);

OAI22xp5_ASAP7_75t_SL g462 ( 
.A1(n_436),
.A2(n_404),
.B1(n_395),
.B2(n_406),
.Y(n_462)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_462),
.Y(n_476)
);

AOI22xp5_ASAP7_75t_L g464 ( 
.A1(n_447),
.A2(n_398),
.B1(n_422),
.B2(n_395),
.Y(n_464)
);

OAI22xp5_ASAP7_75t_SL g477 ( 
.A1(n_464),
.A2(n_472),
.B1(n_429),
.B2(n_439),
.Y(n_477)
);

MAJIxp5_ASAP7_75t_L g466 ( 
.A(n_428),
.B(n_425),
.C(n_443),
.Y(n_466)
);

MAJIxp5_ASAP7_75t_L g484 ( 
.A(n_466),
.B(n_470),
.C(n_425),
.Y(n_484)
);

XNOR2xp5_ASAP7_75t_L g468 ( 
.A(n_435),
.B(n_394),
.Y(n_468)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_469),
.Y(n_478)
);

MAJIxp5_ASAP7_75t_L g470 ( 
.A(n_428),
.B(n_421),
.C(n_407),
.Y(n_470)
);

AOI22xp5_ASAP7_75t_L g472 ( 
.A1(n_429),
.A2(n_421),
.B1(n_402),
.B2(n_401),
.Y(n_472)
);

HB1xp67_ASAP7_75t_L g475 ( 
.A(n_452),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_475),
.B(n_485),
.Y(n_504)
);

AOI22xp5_ASAP7_75t_L g508 ( 
.A1(n_477),
.A2(n_431),
.B1(n_434),
.B2(n_441),
.Y(n_508)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_461),
.Y(n_479)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_479),
.Y(n_498)
);

AOI21xp5_ASAP7_75t_L g494 ( 
.A1(n_480),
.A2(n_483),
.B(n_442),
.Y(n_494)
);

AOI21xp5_ASAP7_75t_L g483 ( 
.A1(n_465),
.A2(n_424),
.B(n_445),
.Y(n_483)
);

MAJIxp5_ASAP7_75t_L g499 ( 
.A(n_484),
.B(n_486),
.C(n_489),
.Y(n_499)
);

NOR2xp33_ASAP7_75t_L g485 ( 
.A(n_470),
.B(n_430),
.Y(n_485)
);

MAJIxp5_ASAP7_75t_L g486 ( 
.A(n_466),
.B(n_454),
.C(n_457),
.Y(n_486)
);

NOR2xp33_ASAP7_75t_SL g487 ( 
.A(n_460),
.B(n_438),
.Y(n_487)
);

CKINVDCx20_ASAP7_75t_R g503 ( 
.A(n_487),
.Y(n_503)
);

XNOR2xp5_ASAP7_75t_L g501 ( 
.A(n_488),
.B(n_463),
.Y(n_501)
);

MAJIxp5_ASAP7_75t_L g489 ( 
.A(n_454),
.B(n_435),
.C(n_440),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_471),
.Y(n_490)
);

CKINVDCx16_ASAP7_75t_R g496 ( 
.A(n_490),
.Y(n_496)
);

MAJIxp5_ASAP7_75t_L g491 ( 
.A(n_468),
.B(n_440),
.C(n_436),
.Y(n_491)
);

MAJIxp5_ASAP7_75t_L g500 ( 
.A(n_491),
.B(n_492),
.C(n_489),
.Y(n_500)
);

MAJIxp5_ASAP7_75t_L g492 ( 
.A(n_458),
.B(n_436),
.C(n_448),
.Y(n_492)
);

AOI21xp5_ASAP7_75t_L g493 ( 
.A1(n_478),
.A2(n_473),
.B(n_442),
.Y(n_493)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_493),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_494),
.B(n_495),
.Y(n_512)
);

OAI22xp5_ASAP7_75t_L g495 ( 
.A1(n_476),
.A2(n_474),
.B1(n_453),
.B2(n_464),
.Y(n_495)
);

OAI321xp33_ASAP7_75t_L g497 ( 
.A1(n_477),
.A2(n_427),
.A3(n_433),
.B1(n_444),
.B2(n_437),
.C(n_426),
.Y(n_497)
);

OAI22xp5_ASAP7_75t_SL g511 ( 
.A1(n_497),
.A2(n_508),
.B1(n_472),
.B2(n_469),
.Y(n_511)
);

XOR2xp5_ASAP7_75t_L g516 ( 
.A(n_500),
.B(n_501),
.Y(n_516)
);

MAJIxp5_ASAP7_75t_L g502 ( 
.A(n_486),
.B(n_463),
.C(n_462),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_502),
.B(n_505),
.Y(n_520)
);

MAJIxp5_ASAP7_75t_L g505 ( 
.A(n_484),
.B(n_459),
.C(n_455),
.Y(n_505)
);

AND2x2_ASAP7_75t_L g506 ( 
.A(n_492),
.B(n_446),
.Y(n_506)
);

AOI22xp5_ASAP7_75t_SL g509 ( 
.A1(n_506),
.A2(n_434),
.B1(n_432),
.B2(n_491),
.Y(n_509)
);

AOI21xp5_ASAP7_75t_L g507 ( 
.A1(n_488),
.A2(n_431),
.B(n_467),
.Y(n_507)
);

OAI21xp5_ASAP7_75t_SL g517 ( 
.A1(n_507),
.A2(n_432),
.B(n_469),
.Y(n_517)
);

OR2x2_ASAP7_75t_L g524 ( 
.A(n_509),
.B(n_518),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g523 ( 
.A(n_511),
.B(n_514),
.Y(n_523)
);

XNOR2xp5_ASAP7_75t_L g513 ( 
.A(n_500),
.B(n_502),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_SL g530 ( 
.A(n_513),
.B(n_515),
.Y(n_530)
);

NOR2xp33_ASAP7_75t_L g514 ( 
.A(n_503),
.B(n_482),
.Y(n_514)
);

XNOR2xp5_ASAP7_75t_L g515 ( 
.A(n_505),
.B(n_482),
.Y(n_515)
);

XNOR2xp5_ASAP7_75t_L g525 ( 
.A(n_517),
.B(n_521),
.Y(n_525)
);

OAI22xp5_ASAP7_75t_SL g518 ( 
.A1(n_498),
.A2(n_451),
.B1(n_396),
.B2(n_402),
.Y(n_518)
);

NOR2xp33_ASAP7_75t_L g519 ( 
.A(n_499),
.B(n_481),
.Y(n_519)
);

NOR2xp33_ASAP7_75t_L g528 ( 
.A(n_519),
.B(n_515),
.Y(n_528)
);

XNOR2xp5_ASAP7_75t_L g521 ( 
.A(n_506),
.B(n_481),
.Y(n_521)
);

AOI22xp5_ASAP7_75t_SL g522 ( 
.A1(n_501),
.A2(n_449),
.B1(n_401),
.B2(n_396),
.Y(n_522)
);

OAI22xp5_ASAP7_75t_L g532 ( 
.A1(n_522),
.A2(n_496),
.B1(n_418),
.B2(n_370),
.Y(n_532)
);

AOI21xp5_ASAP7_75t_L g526 ( 
.A1(n_521),
.A2(n_499),
.B(n_504),
.Y(n_526)
);

OAI21xp5_ASAP7_75t_SL g537 ( 
.A1(n_526),
.A2(n_418),
.B(n_301),
.Y(n_537)
);

OAI21xp5_ASAP7_75t_SL g527 ( 
.A1(n_520),
.A2(n_510),
.B(n_512),
.Y(n_527)
);

AOI21xp5_ASAP7_75t_L g536 ( 
.A1(n_527),
.A2(n_529),
.B(n_370),
.Y(n_536)
);

OR2x2_ASAP7_75t_L g538 ( 
.A(n_528),
.B(n_531),
.Y(n_538)
);

OAI21xp5_ASAP7_75t_SL g529 ( 
.A1(n_513),
.A2(n_493),
.B(n_507),
.Y(n_529)
);

XNOR2x2_ASAP7_75t_SL g531 ( 
.A(n_509),
.B(n_508),
.Y(n_531)
);

NOR2xp33_ASAP7_75t_L g534 ( 
.A(n_532),
.B(n_522),
.Y(n_534)
);

NOR2xp33_ASAP7_75t_SL g533 ( 
.A(n_528),
.B(n_516),
.Y(n_533)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_533),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_SL g541 ( 
.A(n_534),
.B(n_535),
.Y(n_541)
);

AND2x2_ASAP7_75t_L g535 ( 
.A(n_523),
.B(n_516),
.Y(n_535)
);

OAI21xp5_ASAP7_75t_SL g540 ( 
.A1(n_536),
.A2(n_525),
.B(n_530),
.Y(n_540)
);

NOR2xp33_ASAP7_75t_L g542 ( 
.A(n_537),
.B(n_539),
.Y(n_542)
);

NOR2xp33_ASAP7_75t_L g539 ( 
.A(n_524),
.B(n_304),
.Y(n_539)
);

AOI21xp5_ASAP7_75t_L g544 ( 
.A1(n_540),
.A2(n_530),
.B(n_533),
.Y(n_544)
);

AOI21xp5_ASAP7_75t_SL g546 ( 
.A1(n_544),
.A2(n_545),
.B(n_541),
.Y(n_546)
);

AOI21xp5_ASAP7_75t_SL g545 ( 
.A1(n_543),
.A2(n_542),
.B(n_538),
.Y(n_545)
);

INVxp67_ASAP7_75t_L g548 ( 
.A(n_546),
.Y(n_548)
);

AOI21xp5_ASAP7_75t_SL g547 ( 
.A1(n_544),
.A2(n_321),
.B(n_290),
.Y(n_547)
);

CKINVDCx20_ASAP7_75t_R g549 ( 
.A(n_548),
.Y(n_549)
);

NOR2xp67_ASAP7_75t_L g550 ( 
.A(n_549),
.B(n_547),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_SL g551 ( 
.A(n_550),
.B(n_246),
.Y(n_551)
);

XOR2xp5_ASAP7_75t_L g552 ( 
.A(n_551),
.B(n_246),
.Y(n_552)
);


endmodule