module fake_netlist_5_86_n_96 (n_16, n_0, n_12, n_9, n_18, n_22, n_1, n_8, n_10, n_21, n_4, n_11, n_17, n_19, n_7, n_15, n_20, n_5, n_14, n_2, n_13, n_3, n_6, n_96);

input n_16;
input n_0;
input n_12;
input n_9;
input n_18;
input n_22;
input n_1;
input n_8;
input n_10;
input n_21;
input n_4;
input n_11;
input n_17;
input n_19;
input n_7;
input n_15;
input n_20;
input n_5;
input n_14;
input n_2;
input n_13;
input n_3;
input n_6;

output n_96;

wire n_91;
wire n_82;
wire n_24;
wire n_86;
wire n_83;
wire n_61;
wire n_90;
wire n_75;
wire n_65;
wire n_78;
wire n_74;
wire n_57;
wire n_37;
wire n_31;
wire n_66;
wire n_60;
wire n_43;
wire n_58;
wire n_69;
wire n_42;
wire n_45;
wire n_46;
wire n_94;
wire n_38;
wire n_80;
wire n_35;
wire n_73;
wire n_92;
wire n_30;
wire n_33;
wire n_84;
wire n_23;
wire n_29;
wire n_79;
wire n_47;
wire n_25;
wire n_53;
wire n_44;
wire n_40;
wire n_34;
wire n_62;
wire n_71;
wire n_85;
wire n_95;
wire n_59;
wire n_26;
wire n_55;
wire n_49;
wire n_39;
wire n_54;
wire n_67;
wire n_36;
wire n_76;
wire n_87;
wire n_27;
wire n_77;
wire n_64;
wire n_81;
wire n_28;
wire n_89;
wire n_70;
wire n_68;
wire n_93;
wire n_72;
wire n_32;
wire n_41;
wire n_56;
wire n_51;
wire n_63;
wire n_48;
wire n_50;
wire n_52;
wire n_88;

INVx2_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

BUFx2_ASAP7_75t_L g24 ( 
.A(n_21),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_20),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_17),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_SL g31 ( 
.A(n_3),
.B(n_18),
.Y(n_31)
);

BUFx8_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_15),
.B(n_19),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_9),
.B(n_8),
.Y(n_35)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_7),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_SL g37 ( 
.A1(n_4),
.A2(n_22),
.B1(n_16),
.B2(n_1),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_11),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_0),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_13),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_24),
.B(n_1),
.Y(n_41)
);

AOI21xp5_ASAP7_75t_L g42 ( 
.A1(n_31),
.A2(n_2),
.B(n_3),
.Y(n_42)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_27),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_L g44 ( 
.A1(n_29),
.A2(n_2),
.B1(n_4),
.B2(n_39),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_29),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_36),
.B(n_23),
.Y(n_46)
);

NOR2x1p5_ASAP7_75t_L g47 ( 
.A(n_39),
.B(n_36),
.Y(n_47)
);

INVxp67_ASAP7_75t_L g48 ( 
.A(n_32),
.Y(n_48)
);

NAND3xp33_ASAP7_75t_L g49 ( 
.A(n_31),
.B(n_32),
.C(n_34),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g50 ( 
.A(n_26),
.B(n_34),
.Y(n_50)
);

INVxp67_ASAP7_75t_L g51 ( 
.A(n_45),
.Y(n_51)
);

AO31x2_ASAP7_75t_L g52 ( 
.A1(n_46),
.A2(n_23),
.A3(n_25),
.B(n_30),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_50),
.Y(n_53)
);

AOI21xp5_ASAP7_75t_L g54 ( 
.A1(n_49),
.A2(n_42),
.B(n_41),
.Y(n_54)
);

AOI21xp5_ASAP7_75t_L g55 ( 
.A1(n_44),
.A2(n_35),
.B(n_38),
.Y(n_55)
);

BUFx2_ASAP7_75t_L g56 ( 
.A(n_48),
.Y(n_56)
);

OAI21xp33_ASAP7_75t_L g57 ( 
.A1(n_47),
.A2(n_26),
.B(n_34),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_53),
.Y(n_58)
);

AO21x2_ASAP7_75t_L g59 ( 
.A1(n_55),
.A2(n_28),
.B(n_25),
.Y(n_59)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_52),
.Y(n_60)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_51),
.B(n_43),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_57),
.Y(n_62)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_52),
.Y(n_63)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_52),
.Y(n_64)
);

AO21x2_ASAP7_75t_L g65 ( 
.A1(n_54),
.A2(n_30),
.B(n_33),
.Y(n_65)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_58),
.Y(n_66)
);

BUFx2_ASAP7_75t_L g67 ( 
.A(n_62),
.Y(n_67)
);

AND2x2_ASAP7_75t_L g68 ( 
.A(n_61),
.B(n_56),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_65),
.B(n_43),
.Y(n_69)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_59),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_60),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_67),
.B(n_65),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_66),
.Y(n_73)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_71),
.Y(n_74)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_71),
.Y(n_75)
);

BUFx2_ASAP7_75t_L g76 ( 
.A(n_68),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_72),
.B(n_70),
.Y(n_77)
);

NAND3x2_ASAP7_75t_L g78 ( 
.A(n_76),
.B(n_37),
.C(n_59),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_75),
.Y(n_79)
);

OR2x2_ASAP7_75t_L g80 ( 
.A(n_73),
.B(n_69),
.Y(n_80)
);

OAI211xp5_ASAP7_75t_L g81 ( 
.A1(n_75),
.A2(n_33),
.B(n_60),
.C(n_63),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_77),
.B(n_74),
.Y(n_82)
);

AOI211xp5_ASAP7_75t_L g83 ( 
.A1(n_81),
.A2(n_34),
.B(n_40),
.C(n_63),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_80),
.B(n_74),
.Y(n_84)
);

INVxp67_ASAP7_75t_SL g85 ( 
.A(n_79),
.Y(n_85)
);

OAI21xp33_ASAP7_75t_SL g86 ( 
.A1(n_80),
.A2(n_74),
.B(n_64),
.Y(n_86)
);

NOR3x2_ASAP7_75t_L g87 ( 
.A(n_83),
.B(n_78),
.C(n_64),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_84),
.B(n_43),
.Y(n_88)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_85),
.Y(n_89)
);

HB1xp67_ASAP7_75t_L g90 ( 
.A(n_89),
.Y(n_90)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_88),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_87),
.A2(n_82),
.B1(n_40),
.B2(n_86),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_89),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_92),
.A2(n_40),
.B1(n_43),
.B2(n_93),
.Y(n_94)
);

AOI21xp5_ASAP7_75t_L g95 ( 
.A1(n_94),
.A2(n_91),
.B(n_90),
.Y(n_95)
);

OR2x6_ASAP7_75t_L g96 ( 
.A(n_95),
.B(n_40),
.Y(n_96)
);


endmodule