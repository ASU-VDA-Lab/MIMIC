module fake_jpeg_11566_n_56 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_56);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_56;

wire n_13;
wire n_21;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_23;
wire n_10;
wire n_27;
wire n_55;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_20;
wire n_18;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_25;
wire n_17;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;

CKINVDCx20_ASAP7_75t_R g8 ( 
.A(n_2),
.Y(n_8)
);

INVx2_ASAP7_75t_L g9 ( 
.A(n_6),
.Y(n_9)
);

BUFx6f_ASAP7_75t_L g10 ( 
.A(n_7),
.Y(n_10)
);

BUFx6f_ASAP7_75t_L g11 ( 
.A(n_1),
.Y(n_11)
);

BUFx3_ASAP7_75t_L g12 ( 
.A(n_3),
.Y(n_12)
);

INVx8_ASAP7_75t_L g13 ( 
.A(n_1),
.Y(n_13)
);

INVx6_ASAP7_75t_L g14 ( 
.A(n_6),
.Y(n_14)
);

INVx4_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

INVx6_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

INVx8_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

INVx8_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_19),
.Y(n_33)
);

INVx5_ASAP7_75t_L g20 ( 
.A(n_15),
.Y(n_20)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_20),
.Y(n_32)
);

INVx4_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

NAND2x1_ASAP7_75t_SL g35 ( 
.A(n_21),
.B(n_22),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_8),
.B(n_0),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_23),
.B(n_26),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_8),
.B(n_4),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_SL g36 ( 
.A(n_24),
.B(n_27),
.Y(n_36)
);

MAJIxp5_ASAP7_75t_L g25 ( 
.A(n_9),
.B(n_0),
.C(n_4),
.Y(n_25)
);

MAJIxp5_ASAP7_75t_L g34 ( 
.A(n_25),
.B(n_30),
.C(n_11),
.Y(n_34)
);

INVx4_ASAP7_75t_SL g26 ( 
.A(n_10),
.Y(n_26)
);

CKINVDCx12_ASAP7_75t_R g27 ( 
.A(n_13),
.Y(n_27)
);

AOI22xp33_ASAP7_75t_SL g28 ( 
.A1(n_12),
.A2(n_0),
.B1(n_5),
.B2(n_13),
.Y(n_28)
);

OAI32xp33_ASAP7_75t_L g37 ( 
.A1(n_28),
.A2(n_29),
.A3(n_18),
.B1(n_11),
.B2(n_16),
.Y(n_37)
);

BUFx2_ASAP7_75t_L g29 ( 
.A(n_17),
.Y(n_29)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_17),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_L g31 ( 
.A1(n_30),
.A2(n_14),
.B1(n_16),
.B2(n_10),
.Y(n_31)
);

OA21x2_ASAP7_75t_L g41 ( 
.A1(n_31),
.A2(n_37),
.B(n_28),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_34),
.B(n_22),
.Y(n_42)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_33),
.Y(n_39)
);

CKINVDCx16_ASAP7_75t_R g44 ( 
.A(n_39),
.Y(n_44)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_32),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_SL g43 ( 
.A(n_40),
.B(n_41),
.Y(n_43)
);

A2O1A1Ixp33_ASAP7_75t_L g45 ( 
.A1(n_42),
.A2(n_34),
.B(n_38),
.C(n_35),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_45),
.B(n_41),
.Y(n_47)
);

OAI21xp5_ASAP7_75t_SL g46 ( 
.A1(n_43),
.A2(n_41),
.B(n_35),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g50 ( 
.A(n_46),
.B(n_47),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_45),
.A2(n_31),
.B1(n_37),
.B2(n_29),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_48),
.B(n_36),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_49),
.B(n_46),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_50),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g53 ( 
.A(n_51),
.B(n_52),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_52),
.A2(n_44),
.B1(n_14),
.B2(n_18),
.Y(n_54)
);

AOI21xp5_ASAP7_75t_L g55 ( 
.A1(n_54),
.A2(n_20),
.B(n_21),
.Y(n_55)
);

AOI21xp5_ASAP7_75t_L g56 ( 
.A1(n_55),
.A2(n_53),
.B(n_26),
.Y(n_56)
);


endmodule