module fake_jpeg_10031_n_332 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_332);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_332;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g16 ( 
.A(n_14),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_10),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

INVx6_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_14),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_6),
.B(n_4),
.Y(n_24)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_10),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_14),
.Y(n_27)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_12),
.Y(n_30)
);

BUFx12_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_4),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

INVx8_ASAP7_75t_SL g35 ( 
.A(n_10),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_35),
.Y(n_36)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_36),
.Y(n_67)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_35),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_37),
.B(n_38),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_24),
.B(n_0),
.Y(n_38)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_25),
.Y(n_39)
);

INVx8_ASAP7_75t_L g66 ( 
.A(n_39),
.Y(n_66)
);

INVx2_ASAP7_75t_SL g40 ( 
.A(n_25),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_40),
.B(n_31),
.Y(n_50)
);

INVx4_ASAP7_75t_SL g41 ( 
.A(n_35),
.Y(n_41)
);

CKINVDCx16_ASAP7_75t_R g57 ( 
.A(n_41),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_18),
.Y(n_42)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_42),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_18),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_43),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_18),
.Y(n_44)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_44),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_18),
.Y(n_45)
);

BUFx2_ASAP7_75t_L g68 ( 
.A(n_45),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_18),
.Y(n_46)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_46),
.Y(n_56)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_49),
.B(n_52),
.Y(n_93)
);

CKINVDCx16_ASAP7_75t_R g109 ( 
.A(n_50),
.Y(n_109)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

INVx11_ASAP7_75t_L g82 ( 
.A(n_51),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_38),
.B(n_24),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_37),
.A2(n_28),
.B1(n_21),
.B2(n_19),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_53),
.A2(n_54),
.B1(n_61),
.B2(n_20),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_L g54 ( 
.A1(n_39),
.A2(n_28),
.B1(n_21),
.B2(n_25),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_37),
.B(n_24),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_55),
.B(n_58),
.Y(n_105)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_36),
.Y(n_58)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_36),
.Y(n_59)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_59),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_40),
.B(n_16),
.Y(n_60)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_60),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_L g61 ( 
.A1(n_39),
.A2(n_28),
.B1(n_21),
.B2(n_25),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_36),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_62),
.B(n_71),
.Y(n_110)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_39),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_63),
.B(n_65),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_41),
.A2(n_28),
.B1(n_21),
.B2(n_19),
.Y(n_64)
);

OAI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_64),
.A2(n_22),
.B1(n_32),
.B2(n_33),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_40),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_40),
.B(n_16),
.Y(n_70)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_70),
.Y(n_85)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_42),
.Y(n_71)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_49),
.B(n_41),
.Y(n_73)
);

AND2x2_ASAP7_75t_L g134 ( 
.A(n_73),
.B(n_102),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_47),
.B(n_19),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_75),
.B(n_77),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_47),
.A2(n_28),
.B1(n_21),
.B2(n_19),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_76),
.A2(n_87),
.B1(n_96),
.B2(n_97),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_55),
.B(n_20),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_59),
.A2(n_16),
.B1(n_23),
.B2(n_17),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_78),
.A2(n_84),
.B1(n_88),
.B2(n_89),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_52),
.B(n_22),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_79),
.B(n_86),
.Y(n_139)
);

MAJx2_ASAP7_75t_L g81 ( 
.A(n_57),
.B(n_41),
.C(n_29),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_81),
.B(n_94),
.C(n_106),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_L g83 ( 
.A1(n_67),
.A2(n_56),
.B1(n_48),
.B2(n_69),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_83),
.A2(n_56),
.B1(n_69),
.B2(n_48),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_59),
.A2(n_26),
.B1(n_17),
.B2(n_23),
.Y(n_84)
);

OR2x2_ASAP7_75t_L g86 ( 
.A(n_60),
.B(n_30),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_53),
.A2(n_46),
.B1(n_45),
.B2(n_44),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_57),
.A2(n_26),
.B1(n_17),
.B2(n_23),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_67),
.A2(n_27),
.B1(n_26),
.B2(n_30),
.Y(n_89)
);

BUFx3_ASAP7_75t_L g90 ( 
.A(n_66),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_90),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_68),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_91),
.B(n_95),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_92),
.A2(n_108),
.B1(n_67),
.B2(n_48),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_SL g94 ( 
.A(n_53),
.B(n_29),
.Y(n_94)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_70),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_54),
.A2(n_46),
.B1(n_45),
.B2(n_44),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_61),
.A2(n_46),
.B1(n_45),
.B2(n_44),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_65),
.B(n_34),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_98),
.B(n_100),
.Y(n_140)
);

AO22x1_ASAP7_75t_L g99 ( 
.A1(n_63),
.A2(n_43),
.B1(n_42),
.B2(n_29),
.Y(n_99)
);

O2A1O1Ixp33_ASAP7_75t_SL g126 ( 
.A1(n_99),
.A2(n_71),
.B(n_91),
.C(n_81),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_50),
.B(n_34),
.Y(n_100)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_56),
.Y(n_101)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_101),
.Y(n_128)
);

AND2x2_ASAP7_75t_L g102 ( 
.A(n_58),
.B(n_20),
.Y(n_102)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_51),
.Y(n_104)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_104),
.Y(n_117)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_62),
.B(n_22),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_63),
.B(n_34),
.Y(n_107)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_107),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_64),
.A2(n_43),
.B1(n_42),
.B2(n_27),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_111),
.A2(n_95),
.B1(n_80),
.B2(n_85),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_98),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_112),
.B(n_118),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_110),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_103),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_121),
.B(n_124),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_L g142 ( 
.A1(n_122),
.A2(n_101),
.B1(n_74),
.B2(n_82),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_94),
.A2(n_109),
.B1(n_87),
.B2(n_108),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_123),
.A2(n_125),
.B1(n_129),
.B2(n_132),
.Y(n_149)
);

CKINVDCx16_ASAP7_75t_R g124 ( 
.A(n_107),
.Y(n_124)
);

OA21x2_ASAP7_75t_L g156 ( 
.A1(n_126),
.A2(n_106),
.B(n_102),
.Y(n_156)
);

OAI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_127),
.A2(n_137),
.B1(n_85),
.B2(n_80),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_109),
.A2(n_92),
.B1(n_76),
.B2(n_97),
.Y(n_129)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_110),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_130),
.B(n_131),
.Y(n_152)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_105),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_96),
.A2(n_69),
.B1(n_66),
.B2(n_43),
.Y(n_132)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_105),
.Y(n_133)
);

CKINVDCx16_ASAP7_75t_R g145 ( 
.A(n_133),
.Y(n_145)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_82),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_136),
.B(n_141),
.Y(n_174)
);

OAI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_81),
.A2(n_66),
.B1(n_68),
.B2(n_72),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_L g138 ( 
.A1(n_75),
.A2(n_29),
.B1(n_32),
.B2(n_30),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_138),
.A2(n_77),
.B1(n_79),
.B2(n_100),
.Y(n_157)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_102),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_142),
.A2(n_164),
.B1(n_3),
.B2(n_4),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_143),
.B(n_146),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_SL g144 ( 
.A(n_135),
.B(n_73),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_L g181 ( 
.A1(n_144),
.A2(n_163),
.B(n_168),
.Y(n_181)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_116),
.Y(n_146)
);

NAND2xp33_ASAP7_75t_SL g147 ( 
.A(n_126),
.B(n_73),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_SL g183 ( 
.A1(n_147),
.A2(n_156),
.B(n_158),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_124),
.B(n_112),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_150),
.B(n_160),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_116),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_151),
.B(n_153),
.Y(n_182)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_132),
.Y(n_153)
);

INVxp67_ASAP7_75t_L g154 ( 
.A(n_115),
.Y(n_154)
);

INVxp67_ASAP7_75t_L g199 ( 
.A(n_154),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_138),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_155),
.B(n_162),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_157),
.A2(n_173),
.B1(n_134),
.B2(n_128),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_L g158 ( 
.A1(n_135),
.A2(n_93),
.B(n_106),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_123),
.B(n_93),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_159),
.B(n_15),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_113),
.B(n_119),
.Y(n_160)
);

CKINVDCx16_ASAP7_75t_R g162 ( 
.A(n_122),
.Y(n_162)
);

AOI21xp5_ASAP7_75t_L g163 ( 
.A1(n_115),
.A2(n_104),
.B(n_31),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_L g164 ( 
.A1(n_131),
.A2(n_74),
.B1(n_99),
.B2(n_32),
.Y(n_164)
);

INVx6_ASAP7_75t_L g165 ( 
.A(n_128),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_165),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_113),
.B(n_119),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_166),
.B(n_169),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_141),
.B(n_139),
.C(n_140),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_167),
.B(n_170),
.Y(n_205)
);

A2O1A1Ixp33_ASAP7_75t_SL g168 ( 
.A1(n_126),
.A2(n_99),
.B(n_90),
.C(n_68),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_140),
.B(n_86),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_139),
.B(n_86),
.C(n_72),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_137),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_171),
.B(n_0),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_114),
.A2(n_27),
.B1(n_72),
.B2(n_33),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_172),
.A2(n_117),
.B1(n_120),
.B2(n_114),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_125),
.A2(n_33),
.B1(n_31),
.B2(n_2),
.Y(n_173)
);

INVxp67_ASAP7_75t_L g175 ( 
.A(n_127),
.Y(n_175)
);

HB1xp67_ASAP7_75t_L g190 ( 
.A(n_175),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_154),
.A2(n_134),
.B1(n_118),
.B2(n_129),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_176),
.B(n_186),
.Y(n_209)
);

AND2x2_ASAP7_75t_SL g177 ( 
.A(n_171),
.B(n_130),
.Y(n_177)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_177),
.Y(n_213)
);

BUFx4f_ASAP7_75t_SL g178 ( 
.A(n_165),
.Y(n_178)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_178),
.Y(n_210)
);

BUFx6f_ASAP7_75t_L g179 ( 
.A(n_145),
.Y(n_179)
);

INVx13_ASAP7_75t_L g228 ( 
.A(n_179),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_185),
.A2(n_193),
.B1(n_194),
.B2(n_196),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_175),
.A2(n_134),
.B1(n_117),
.B2(n_31),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_189),
.B(n_197),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_149),
.A2(n_134),
.B1(n_136),
.B2(n_31),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_192),
.A2(n_201),
.B1(n_170),
.B2(n_158),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_153),
.A2(n_31),
.B1(n_1),
.B2(n_2),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_149),
.A2(n_31),
.B1(n_1),
.B2(n_2),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_195),
.B(n_159),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_172),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_150),
.Y(n_197)
);

OAI32xp33_ASAP7_75t_L g211 ( 
.A1(n_198),
.A2(n_169),
.A3(n_160),
.B1(n_166),
.B2(n_157),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_152),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_200),
.B(n_208),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_163),
.A2(n_0),
.B1(n_3),
.B2(n_4),
.Y(n_201)
);

CKINVDCx16_ASAP7_75t_R g202 ( 
.A(n_174),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_SL g230 ( 
.A(n_202),
.B(n_203),
.Y(n_230)
);

CKINVDCx16_ASAP7_75t_R g203 ( 
.A(n_161),
.Y(n_203)
);

INVx8_ASAP7_75t_L g204 ( 
.A(n_145),
.Y(n_204)
);

AOI22xp33_ASAP7_75t_SL g214 ( 
.A1(n_204),
.A2(n_151),
.B1(n_168),
.B2(n_155),
.Y(n_214)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_206),
.Y(n_219)
);

INVx4_ASAP7_75t_L g207 ( 
.A(n_146),
.Y(n_207)
);

INVx1_ASAP7_75t_SL g218 ( 
.A(n_207),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_148),
.Y(n_208)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_211),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_214),
.A2(n_199),
.B1(n_187),
.B2(n_204),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_215),
.B(n_220),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_216),
.B(n_195),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_205),
.B(n_144),
.C(n_167),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_217),
.B(n_225),
.Y(n_238)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_182),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_180),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_221),
.B(n_224),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_180),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_SL g250 ( 
.A(n_222),
.B(n_229),
.Y(n_250)
);

INVx1_ASAP7_75t_SL g224 ( 
.A(n_207),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_205),
.B(n_147),
.C(n_156),
.Y(n_225)
);

OA21x2_ASAP7_75t_L g226 ( 
.A1(n_177),
.A2(n_168),
.B(n_156),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_L g243 ( 
.A1(n_226),
.A2(n_186),
.B(n_181),
.Y(n_243)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_188),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_188),
.B(n_197),
.Y(n_231)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_231),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_176),
.A2(n_168),
.B1(n_173),
.B2(n_6),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_232),
.A2(n_234),
.B1(n_235),
.B2(n_198),
.Y(n_239)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_184),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_SL g257 ( 
.A(n_233),
.B(n_196),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_192),
.A2(n_168),
.B1(n_5),
.B2(n_6),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_185),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_183),
.B(n_11),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_236),
.B(n_201),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_231),
.B(n_208),
.Y(n_237)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_237),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_239),
.A2(n_245),
.B1(n_254),
.B2(n_255),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_240),
.B(n_244),
.C(n_215),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_227),
.B(n_177),
.Y(n_241)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_241),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_227),
.B(n_191),
.Y(n_242)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_242),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_SL g276 ( 
.A(n_243),
.B(n_245),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_209),
.B(n_181),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_223),
.A2(n_199),
.B1(n_189),
.B2(n_190),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_230),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_247),
.B(n_252),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_223),
.B(n_200),
.Y(n_249)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_249),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_213),
.B(n_194),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_253),
.B(n_258),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_219),
.A2(n_183),
.B1(n_187),
.B2(n_193),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_257),
.B(n_259),
.Y(n_266)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_225),
.B(n_179),
.Y(n_258)
);

BUFx5_ASAP7_75t_L g259 ( 
.A(n_228),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_258),
.B(n_217),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_260),
.B(n_261),
.C(n_265),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_256),
.A2(n_209),
.B1(n_232),
.B2(n_226),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_263),
.A2(n_212),
.B1(n_218),
.B2(n_250),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_238),
.B(n_240),
.C(n_216),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_246),
.B(n_236),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_268),
.B(n_274),
.C(n_277),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_242),
.B(n_224),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_SL g283 ( 
.A(n_269),
.B(n_278),
.Y(n_283)
);

AND2x2_ASAP7_75t_L g272 ( 
.A(n_253),
.B(n_244),
.Y(n_272)
);

AOI21xp5_ASAP7_75t_L g290 ( 
.A1(n_272),
.A2(n_261),
.B(n_274),
.Y(n_290)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_238),
.B(n_226),
.Y(n_274)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_276),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_243),
.B(n_211),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_241),
.B(n_218),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_262),
.B(n_237),
.Y(n_279)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_279),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_275),
.B(n_249),
.Y(n_280)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_280),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_L g281 ( 
.A1(n_267),
.A2(n_252),
.B1(n_212),
.B2(n_235),
.Y(n_281)
);

INVxp67_ASAP7_75t_L g294 ( 
.A(n_281),
.Y(n_294)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_266),
.Y(n_285)
);

AOI21xp5_ASAP7_75t_L g297 ( 
.A1(n_285),
.A2(n_286),
.B(n_291),
.Y(n_297)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_271),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_265),
.B(n_248),
.C(n_251),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_288),
.B(n_289),
.C(n_276),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_264),
.B(n_248),
.C(n_255),
.Y(n_289)
);

XOR2xp5_ASAP7_75t_L g301 ( 
.A(n_290),
.B(n_292),
.Y(n_301)
);

OAI21xp5_ASAP7_75t_SL g291 ( 
.A1(n_270),
.A2(n_239),
.B(n_234),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_277),
.B(n_259),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_293),
.B(n_263),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_295),
.B(n_302),
.Y(n_315)
);

BUFx24_ASAP7_75t_SL g296 ( 
.A(n_285),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_296),
.B(n_304),
.Y(n_309)
);

INVxp67_ASAP7_75t_L g298 ( 
.A(n_279),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_298),
.B(n_303),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_282),
.A2(n_272),
.B1(n_273),
.B2(n_264),
.Y(n_302)
);

HB1xp67_ASAP7_75t_L g304 ( 
.A(n_291),
.Y(n_304)
);

NAND4xp25_ASAP7_75t_SL g305 ( 
.A(n_283),
.B(n_178),
.C(n_210),
.D(n_228),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_305),
.B(n_11),
.Y(n_314)
);

AOI21xp5_ASAP7_75t_L g306 ( 
.A1(n_282),
.A2(n_178),
.B(n_210),
.Y(n_306)
);

OAI21xp5_ASAP7_75t_L g313 ( 
.A1(n_306),
.A2(n_5),
.B(n_7),
.Y(n_313)
);

AOI21xp5_ASAP7_75t_L g307 ( 
.A1(n_298),
.A2(n_288),
.B(n_289),
.Y(n_307)
);

OAI21xp5_ASAP7_75t_SL g318 ( 
.A1(n_307),
.A2(n_313),
.B(n_301),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_L g308 ( 
.A1(n_294),
.A2(n_280),
.B1(n_286),
.B2(n_292),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_308),
.B(n_312),
.Y(n_317)
);

AOI22xp33_ASAP7_75t_SL g310 ( 
.A1(n_300),
.A2(n_290),
.B1(n_287),
.B2(n_284),
.Y(n_310)
);

AO22x1_ASAP7_75t_L g316 ( 
.A1(n_310),
.A2(n_301),
.B1(n_297),
.B2(n_299),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_294),
.A2(n_287),
.B1(n_284),
.B2(n_11),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_314),
.B(n_7),
.Y(n_322)
);

XOR2xp5_ASAP7_75t_L g323 ( 
.A(n_316),
.B(n_313),
.Y(n_323)
);

XOR2xp5_ASAP7_75t_L g324 ( 
.A(n_318),
.B(n_319),
.Y(n_324)
);

OAI21x1_ASAP7_75t_L g319 ( 
.A1(n_310),
.A2(n_12),
.B(n_13),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_309),
.B(n_311),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_320),
.B(n_321),
.Y(n_325)
);

XNOR2xp5_ASAP7_75t_L g321 ( 
.A(n_315),
.B(n_13),
.Y(n_321)
);

OAI21xp5_ASAP7_75t_SL g326 ( 
.A1(n_322),
.A2(n_8),
.B(n_9),
.Y(n_326)
);

AOI21xp5_ASAP7_75t_L g327 ( 
.A1(n_323),
.A2(n_326),
.B(n_322),
.Y(n_327)
);

INVxp67_ASAP7_75t_L g329 ( 
.A(n_327),
.Y(n_329)
);

AOI21xp5_ASAP7_75t_L g328 ( 
.A1(n_325),
.A2(n_317),
.B(n_315),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_L g330 ( 
.A1(n_329),
.A2(n_328),
.B1(n_324),
.B2(n_323),
.Y(n_330)
);

AOI22xp5_ASAP7_75t_SL g331 ( 
.A1(n_330),
.A2(n_8),
.B1(n_9),
.B2(n_319),
.Y(n_331)
);

XNOR2xp5_ASAP7_75t_L g332 ( 
.A(n_331),
.B(n_8),
.Y(n_332)
);


endmodule