module fake_jpeg_22751_n_105 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_105);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_105;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_57;
wire n_21;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_1),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_7),
.Y(n_12)
);

INVx1_ASAP7_75t_SL g13 ( 
.A(n_6),
.Y(n_13)
);

INVx4_ASAP7_75t_L g14 ( 
.A(n_2),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_10),
.B(n_4),
.Y(n_17)
);

INVx11_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_9),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_23),
.B(n_24),
.Y(n_32)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_17),
.B(n_0),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_25),
.B(n_27),
.Y(n_31)
);

INVx11_ASAP7_75t_L g26 ( 
.A(n_18),
.Y(n_26)
);

BUFx10_ASAP7_75t_L g38 ( 
.A(n_26),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_11),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_11),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_28),
.B(n_29),
.Y(n_33)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_18),
.Y(n_29)
);

INVx4_ASAP7_75t_SL g30 ( 
.A(n_13),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_30),
.B(n_13),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_25),
.B(n_17),
.Y(n_34)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_SL g40 ( 
.A(n_35),
.B(n_36),
.Y(n_40)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_29),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_37),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_26),
.Y(n_39)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_39),
.Y(n_47)
);

AOI21xp5_ASAP7_75t_L g42 ( 
.A1(n_36),
.A2(n_14),
.B(n_24),
.Y(n_42)
);

AOI21xp5_ASAP7_75t_L g53 ( 
.A1(n_42),
.A2(n_51),
.B(n_44),
.Y(n_53)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_38),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_44),
.B(n_45),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g45 ( 
.A1(n_34),
.A2(n_23),
.B1(n_17),
.B2(n_18),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_31),
.B(n_16),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_46),
.B(n_43),
.Y(n_55)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_33),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_48),
.B(n_28),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_33),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_49),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g50 ( 
.A(n_31),
.B(n_30),
.Y(n_50)
);

XNOR2xp5_ASAP7_75t_L g60 ( 
.A(n_50),
.B(n_51),
.Y(n_60)
);

MAJIxp5_ASAP7_75t_L g51 ( 
.A(n_32),
.B(n_13),
.C(n_30),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_46),
.B(n_27),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_52),
.B(n_55),
.Y(n_71)
);

AOI21xp5_ASAP7_75t_L g68 ( 
.A1(n_53),
.A2(n_15),
.B(n_22),
.Y(n_68)
);

BUFx2_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_56),
.B(n_59),
.Y(n_64)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_57),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_43),
.B(n_15),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_45),
.B(n_15),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_61),
.B(n_62),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_50),
.B(n_40),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_50),
.B(n_38),
.Y(n_63)
);

XNOR2xp5_ASAP7_75t_L g72 ( 
.A(n_63),
.B(n_38),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_53),
.B(n_42),
.C(n_47),
.Y(n_65)
);

INVxp67_ASAP7_75t_L g80 ( 
.A(n_65),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_58),
.B(n_20),
.Y(n_67)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_67),
.Y(n_81)
);

OAI21xp5_ASAP7_75t_L g75 ( 
.A1(n_68),
.A2(n_69),
.B(n_70),
.Y(n_75)
);

XOR2xp5_ASAP7_75t_L g69 ( 
.A(n_60),
.B(n_38),
.Y(n_69)
);

XOR2xp5_ASAP7_75t_L g70 ( 
.A(n_60),
.B(n_38),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_72),
.B(n_56),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_65),
.A2(n_54),
.B1(n_63),
.B2(n_55),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_74),
.A2(n_82),
.B1(n_22),
.B2(n_21),
.Y(n_85)
);

XNOR2xp5_ASAP7_75t_SL g88 ( 
.A(n_76),
.B(n_39),
.Y(n_88)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_73),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_77),
.B(n_78),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_71),
.B(n_12),
.Y(n_78)
);

OAI32xp33_ASAP7_75t_L g79 ( 
.A1(n_66),
.A2(n_22),
.A3(n_21),
.B1(n_19),
.B2(n_16),
.Y(n_79)
);

XOR2xp5_ASAP7_75t_L g86 ( 
.A(n_79),
.B(n_21),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_72),
.A2(n_70),
.B1(n_69),
.B2(n_68),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_80),
.A2(n_64),
.B1(n_12),
.B2(n_20),
.Y(n_84)
);

XNOR2xp5_ASAP7_75t_L g92 ( 
.A(n_84),
.B(n_86),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_85),
.B(n_88),
.C(n_82),
.Y(n_89)
);

NAND2x1_ASAP7_75t_L g87 ( 
.A(n_75),
.B(n_39),
.Y(n_87)
);

AOI21xp5_ASAP7_75t_L g93 ( 
.A1(n_87),
.A2(n_37),
.B(n_2),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_89),
.A2(n_93),
.B1(n_83),
.B2(n_84),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_88),
.B(n_75),
.C(n_74),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_90),
.B(n_86),
.Y(n_94)
);

AOI322xp5_ASAP7_75t_L g91 ( 
.A1(n_87),
.A2(n_80),
.A3(n_81),
.B1(n_37),
.B2(n_19),
.C1(n_16),
.C2(n_7),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_91),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_L g99 ( 
.A1(n_94),
.A2(n_5),
.B(n_10),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_95),
.B(n_91),
.Y(n_98)
);

AOI21xp5_ASAP7_75t_SL g97 ( 
.A1(n_92),
.A2(n_5),
.B(n_9),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_SL g100 ( 
.A1(n_97),
.A2(n_1),
.B(n_2),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_98),
.B(n_99),
.C(n_1),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_100),
.B(n_96),
.Y(n_101)
);

AOI21x1_ASAP7_75t_L g103 ( 
.A1(n_101),
.A2(n_102),
.B(n_3),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_103),
.B(n_3),
.C(n_4),
.Y(n_104)
);

XOR2xp5_ASAP7_75t_L g105 ( 
.A(n_104),
.B(n_3),
.Y(n_105)
);


endmodule