module fake_jpeg_13981_n_52 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_52);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_52;

wire n_21;
wire n_33;
wire n_45;
wire n_23;
wire n_27;
wire n_22;
wire n_47;
wire n_51;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_44;
wire n_26;
wire n_38;
wire n_36;
wire n_31;
wire n_25;
wire n_17;
wire n_29;
wire n_43;
wire n_50;
wire n_37;
wire n_32;
wire n_15;

INVx5_ASAP7_75t_L g15 ( 
.A(n_11),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

BUFx12_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_1),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

CKINVDCx10_ASAP7_75t_R g29 ( 
.A(n_7),
.Y(n_29)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_22),
.Y(n_30)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_30),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_29),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_31),
.B(n_32),
.Y(n_42)
);

INVxp67_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

XNOR2xp5_ASAP7_75t_SL g33 ( 
.A(n_28),
.B(n_0),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_L g43 ( 
.A1(n_33),
.A2(n_34),
.B1(n_35),
.B2(n_36),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_26),
.B(n_0),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_28),
.B(n_25),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g36 ( 
.A(n_25),
.B(n_14),
.Y(n_36)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_23),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_23),
.Y(n_39)
);

OR2x2_ASAP7_75t_L g40 ( 
.A(n_24),
.B(n_21),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_43),
.B(n_36),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_44),
.B(n_40),
.Y(n_47)
);

XNOR2xp5_ASAP7_75t_L g45 ( 
.A(n_42),
.B(n_38),
.Y(n_45)
);

XNOR2xp5_ASAP7_75t_SL g46 ( 
.A(n_45),
.B(n_40),
.Y(n_46)
);

MAJIxp5_ASAP7_75t_L g48 ( 
.A(n_46),
.B(n_47),
.C(n_41),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_48),
.B(n_49),
.Y(n_50)
);

AND2x2_ASAP7_75t_L g49 ( 
.A(n_47),
.B(n_39),
.Y(n_49)
);

AOI21xp5_ASAP7_75t_L g51 ( 
.A1(n_50),
.A2(n_37),
.B(n_15),
.Y(n_51)
);

OAI221xp5_ASAP7_75t_L g52 ( 
.A1(n_51),
.A2(n_20),
.B1(n_19),
.B2(n_17),
.C(n_27),
.Y(n_52)
);


endmodule