module real_jpeg_26731_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_249;
wire n_215;
wire n_176;
wire n_166;
wire n_221;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_280;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_281;
wire n_271;
wire n_276;
wire n_163;
wire n_22;
wire n_237;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_243;
wire n_173;
wire n_255;
wire n_115;
wire n_98;
wire n_27;
wire n_184;
wire n_56;
wire n_48;
wire n_164;
wire n_200;
wire n_275;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_13;
wire n_113;
wire n_155;
wire n_120;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_211;
wire n_172;
wire n_45;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_262;
wire n_222;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_205;
wire n_258;
wire n_117;
wire n_193;
wire n_99;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_150;
wire n_32;
wire n_20;
wire n_80;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_259;
wire n_103;
wire n_225;
wire n_232;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_277;
wire n_125;
wire n_240;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_279;
wire n_59;
wire n_169;
wire n_128;
wire n_202;
wire n_167;
wire n_216;
wire n_244;
wire n_179;
wire n_133;
wire n_213;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_210;
wire n_127;
wire n_206;
wire n_224;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_181;
wire n_101;
wire n_256;
wire n_274;
wire n_182;
wire n_273;
wire n_269;
wire n_96;
wire n_253;
wire n_89;
wire n_16;

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_0),
.B(n_50),
.Y(n_81)
);

INVx11_ASAP7_75t_L g83 ( 
.A(n_0),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_0),
.B(n_98),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_0),
.B(n_211),
.Y(n_216)
);

BUFx12_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_2),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g27 ( 
.A1(n_3),
.A2(n_4),
.B1(n_28),
.B2(n_29),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_3),
.Y(n_29)
);

OAI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_3),
.A2(n_23),
.B1(n_24),
.B2(n_29),
.Y(n_67)
);

OAI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_3),
.A2(n_29),
.B1(n_42),
.B2(n_46),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_3),
.A2(n_29),
.B1(n_48),
.B2(n_50),
.Y(n_98)
);

INVx13_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_4),
.A2(n_5),
.B1(n_28),
.B2(n_113),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_5),
.Y(n_113)
);

OAI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_5),
.A2(n_23),
.B1(n_24),
.B2(n_113),
.Y(n_140)
);

OAI22xp33_ASAP7_75t_SL g184 ( 
.A1(n_5),
.A2(n_42),
.B1(n_46),
.B2(n_113),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_5),
.A2(n_48),
.B1(n_50),
.B2(n_113),
.Y(n_211)
);

AOI22xp33_ASAP7_75t_L g63 ( 
.A1(n_6),
.A2(n_23),
.B1(n_24),
.B2(n_64),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_6),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_6),
.A2(n_42),
.B1(n_46),
.B2(n_64),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_6),
.A2(n_48),
.B1(n_50),
.B2(n_64),
.Y(n_129)
);

INVx11_ASAP7_75t_L g44 ( 
.A(n_7),
.Y(n_44)
);

AOI21xp33_ASAP7_75t_L g202 ( 
.A1(n_7),
.A2(n_10),
.B(n_48),
.Y(n_202)
);

BUFx24_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_9),
.Y(n_57)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_9),
.Y(n_60)
);

AOI21xp33_ASAP7_75t_SL g177 ( 
.A1(n_9),
.A2(n_10),
.B(n_42),
.Y(n_177)
);

AOI21xp5_ASAP7_75t_L g34 ( 
.A1(n_10),
.A2(n_28),
.B(n_35),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_10),
.B(n_28),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_10),
.A2(n_42),
.B1(n_46),
.B2(n_54),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_10),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_10),
.A2(n_48),
.B1(n_50),
.B2(n_54),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_10),
.A2(n_23),
.B1(n_24),
.B2(n_54),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_10),
.B(n_20),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_10),
.B(n_59),
.Y(n_206)
);

INVx11_ASAP7_75t_SL g49 ( 
.A(n_11),
.Y(n_49)
);

XNOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_121),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_119),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_SL g14 ( 
.A(n_15),
.B(n_89),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_15),
.B(n_89),
.Y(n_120)
);

BUFx24_ASAP7_75t_SL g283 ( 
.A(n_15),
.Y(n_283)
);

FAx1_ASAP7_75t_SL g15 ( 
.A(n_16),
.B(n_68),
.CI(n_76),
.CON(n_15),
.SN(n_15)
);

AOI22xp5_ASAP7_75t_L g16 ( 
.A1(n_17),
.A2(n_18),
.B1(n_36),
.B2(n_37),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_18),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_30),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_19),
.B(n_109),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_26),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_20),
.B(n_108),
.Y(n_107)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

A2O1A1Ixp33_ASAP7_75t_L g32 ( 
.A1(n_21),
.A2(n_22),
.B(n_28),
.C(n_33),
.Y(n_32)
);

AOI21xp5_ASAP7_75t_L g88 ( 
.A1(n_21),
.A2(n_32),
.B(n_34),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_21),
.B(n_112),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_23),
.B1(n_24),
.B2(n_25),
.Y(n_21)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_22),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_22),
.B(n_28),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_23),
.B(n_25),
.Y(n_153)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

O2A1O1Ixp33_ASAP7_75t_L g56 ( 
.A1(n_24),
.A2(n_57),
.B(n_58),
.C(n_59),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_24),
.B(n_57),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_24),
.A2(n_153),
.B1(n_154),
.B2(n_155),
.Y(n_152)
);

A2O1A1Ixp33_ASAP7_75t_L g176 ( 
.A1(n_24),
.A2(n_54),
.B(n_60),
.C(n_177),
.Y(n_176)
);

CKINVDCx16_ASAP7_75t_R g26 ( 
.A(n_27),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_27),
.B(n_32),
.Y(n_256)
);

INVxp67_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_31),
.B(n_135),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g31 ( 
.A(n_32),
.B(n_34),
.Y(n_31)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_32),
.Y(n_110)
);

CKINVDCx16_ASAP7_75t_R g155 ( 
.A(n_33),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_34),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g154 ( 
.A(n_35),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_37),
.Y(n_36)
);

XNOR2xp5_ASAP7_75t_SL g37 ( 
.A(n_38),
.B(n_55),
.Y(n_37)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_38),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_38),
.A2(n_136),
.B1(n_137),
.B2(n_138),
.Y(n_161)
);

AOI21xp5_ASAP7_75t_SL g38 ( 
.A1(n_39),
.A2(n_51),
.B(n_52),
.Y(n_38)
);

OAI21xp5_ASAP7_75t_SL g85 ( 
.A1(n_39),
.A2(n_86),
.B(n_87),
.Y(n_85)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_40),
.B(n_75),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_40),
.B(n_53),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_40),
.B(n_184),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_41),
.B(n_47),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_L g41 ( 
.A1(n_42),
.A2(n_44),
.B1(n_45),
.B2(n_46),
.Y(n_41)
);

INVx4_ASAP7_75t_SL g46 ( 
.A(n_42),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_42),
.A2(n_46),
.B1(n_60),
.B2(n_61),
.Y(n_59)
);

A2O1A1Ixp33_ASAP7_75t_L g201 ( 
.A1(n_42),
.A2(n_44),
.B(n_54),
.C(n_202),
.Y(n_201)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx11_ASAP7_75t_L g45 ( 
.A(n_44),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g47 ( 
.A1(n_44),
.A2(n_45),
.B1(n_48),
.B2(n_50),
.Y(n_47)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_47),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_47),
.B(n_53),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_47),
.B(n_75),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_47),
.B(n_184),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_48),
.Y(n_50)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_50),
.B(n_226),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_L g100 ( 
.A1(n_51),
.A2(n_74),
.B(n_86),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g221 ( 
.A(n_51),
.B(n_54),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_53),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_54),
.B(n_227),
.Y(n_226)
);

AOI21xp5_ASAP7_75t_L g55 ( 
.A1(n_56),
.A2(n_62),
.B(n_65),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_56),
.B(n_67),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_56),
.B(n_104),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_56),
.B(n_140),
.Y(n_150)
);

INVxp67_ASAP7_75t_L g259 ( 
.A(n_56),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_59),
.B(n_67),
.Y(n_66)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_59),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_59),
.B(n_140),
.Y(n_139)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_60),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_63),
.Y(n_62)
);

OAI21xp5_ASAP7_75t_SL g69 ( 
.A1(n_63),
.A2(n_70),
.B(n_71),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_65),
.B(n_102),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_66),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_66),
.B(n_150),
.Y(n_165)
);

AOI21xp5_ASAP7_75t_L g114 ( 
.A1(n_68),
.A2(n_69),
.B(n_72),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_69),
.B(n_72),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_70),
.B(n_148),
.Y(n_147)
);

AOI21xp5_ASAP7_75t_L g258 ( 
.A1(n_70),
.A2(n_148),
.B(n_259),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_71),
.B(n_139),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_73),
.B(n_74),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_73),
.B(n_193),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_74),
.B(n_183),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_L g76 ( 
.A1(n_77),
.A2(n_80),
.B(n_88),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_77),
.A2(n_78),
.B1(n_116),
.B2(n_117),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_78),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_85),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_79),
.A2(n_80),
.B1(n_88),
.B2(n_118),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_79),
.A2(n_80),
.B1(n_176),
.B2(n_178),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g272 ( 
.A1(n_79),
.A2(n_80),
.B1(n_85),
.B2(n_273),
.Y(n_272)
);

CKINVDCx16_ASAP7_75t_R g79 ( 
.A(n_80),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_80),
.B(n_176),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_SL g80 ( 
.A1(n_81),
.A2(n_82),
.B(n_84),
.Y(n_80)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_81),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_81),
.B(n_84),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_81),
.B(n_211),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_82),
.B(n_84),
.Y(n_94)
);

INVx11_ASAP7_75t_L g157 ( 
.A(n_82),
.Y(n_157)
);

INVx5_ASAP7_75t_SL g227 ( 
.A(n_82),
.Y(n_227)
);

INVx11_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_85),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_87),
.B(n_132),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_87),
.B(n_193),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_88),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_114),
.C(n_115),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g278 ( 
.A1(n_90),
.A2(n_91),
.B1(n_279),
.B2(n_280),
.Y(n_278)
);

CKINVDCx16_ASAP7_75t_R g90 ( 
.A(n_91),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_101),
.C(n_105),
.Y(n_91)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_92),
.B(n_269),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_100),
.Y(n_92)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_93),
.B(n_100),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_95),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_94),
.B(n_210),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_L g156 ( 
.A1(n_95),
.A2(n_129),
.B(n_157),
.Y(n_156)
);

CKINVDCx16_ASAP7_75t_R g95 ( 
.A(n_96),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_96),
.B(n_215),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_SL g96 ( 
.A(n_97),
.B(n_99),
.Y(n_96)
);

INVxp33_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_L g128 ( 
.A1(n_99),
.A2(n_129),
.B(n_130),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_101),
.A2(n_105),
.B1(n_106),
.B2(n_270),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_101),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_103),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_103),
.B(n_139),
.Y(n_180)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_104),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_106),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_107),
.B(n_109),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_110),
.B(n_111),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_112),
.Y(n_111)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_114),
.B(n_115),
.Y(n_280)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

AOI21xp5_ASAP7_75t_L g121 ( 
.A1(n_122),
.A2(n_276),
.B(n_281),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_SL g122 ( 
.A1(n_123),
.A2(n_263),
.B(n_275),
.Y(n_122)
);

O2A1O1Ixp33_ASAP7_75t_SL g123 ( 
.A1(n_124),
.A2(n_170),
.B(n_245),
.C(n_262),
.Y(n_123)
);

AND2x2_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_158),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_125),
.B(n_158),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_141),
.Y(n_125)
);

XOR2xp5_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_133),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_127),
.B(n_133),
.C(n_141),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_131),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_128),
.B(n_131),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_130),
.B(n_169),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_130),
.B(n_210),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_132),
.B(n_183),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_136),
.C(n_137),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_134),
.B(n_161),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_135),
.B(n_256),
.Y(n_255)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_SL g141 ( 
.A(n_142),
.B(n_151),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_143),
.A2(n_144),
.B1(n_145),
.B2(n_146),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_143),
.B(n_146),
.C(n_151),
.Y(n_260)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_149),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_150),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_156),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_152),
.B(n_156),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_162),
.C(n_164),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_159),
.A2(n_160),
.B1(n_240),
.B2(n_241),
.Y(n_239)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g241 ( 
.A1(n_162),
.A2(n_163),
.B1(n_164),
.B2(n_242),
.Y(n_241)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_164),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_166),
.C(n_168),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_165),
.B(n_188),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_166),
.A2(n_167),
.B1(n_168),
.B2(n_189),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_167),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_168),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_169),
.B(n_216),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_SL g170 ( 
.A(n_171),
.B(n_244),
.Y(n_170)
);

AOI21xp5_ASAP7_75t_L g171 ( 
.A1(n_172),
.A2(n_237),
.B(n_243),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_L g172 ( 
.A1(n_173),
.A2(n_195),
.B(n_236),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_185),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_174),
.B(n_185),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_179),
.C(n_181),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_175),
.B(n_234),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_176),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_179),
.A2(n_180),
.B1(n_181),
.B2(n_182),
.Y(n_234)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_182),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_186),
.A2(n_187),
.B1(n_190),
.B2(n_191),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_186),
.B(n_192),
.C(n_194),
.Y(n_238)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_194),
.Y(n_191)
);

AOI21xp5_ASAP7_75t_L g195 ( 
.A1(n_196),
.A2(n_231),
.B(n_235),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_L g196 ( 
.A1(n_197),
.A2(n_212),
.B(n_230),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_203),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_198),
.B(n_203),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_SL g198 ( 
.A(n_199),
.B(n_201),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_199),
.A2(n_200),
.B1(n_201),
.B2(n_218),
.Y(n_217)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_201),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_209),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_205),
.A2(n_206),
.B1(n_207),
.B2(n_208),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_205),
.B(n_208),
.C(n_209),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_206),
.Y(n_205)
);

CKINVDCx16_ASAP7_75t_R g207 ( 
.A(n_208),
.Y(n_207)
);

AOI21xp5_ASAP7_75t_L g212 ( 
.A1(n_213),
.A2(n_219),
.B(n_229),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_217),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_SL g229 ( 
.A(n_214),
.B(n_217),
.Y(n_229)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_SL g219 ( 
.A1(n_220),
.A2(n_223),
.B(n_228),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_222),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_221),
.B(n_222),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_224),
.B(n_225),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_233),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_SL g235 ( 
.A(n_232),
.B(n_233),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_238),
.B(n_239),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_SL g243 ( 
.A(n_238),
.B(n_239),
.Y(n_243)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_247),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_SL g262 ( 
.A(n_246),
.B(n_247),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_248),
.A2(n_249),
.B1(n_260),
.B2(n_261),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_251),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_250),
.B(n_251),
.C(n_261),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_253),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_252),
.B(n_255),
.C(n_257),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_254),
.A2(n_255),
.B1(n_257),
.B2(n_258),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_258),
.Y(n_257)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_260),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_264),
.B(n_265),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_264),
.B(n_265),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_266),
.B(n_274),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_267),
.A2(n_268),
.B1(n_271),
.B2(n_272),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_267),
.B(n_272),
.C(n_274),
.Y(n_277)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_272),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_278),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_SL g281 ( 
.A(n_277),
.B(n_278),
.Y(n_281)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);


endmodule