module real_jpeg_27308_n_18 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_3, n_329, n_5, n_4, n_1, n_328, n_16, n_15, n_13, n_18);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_3;
input n_329;
input n_5;
input n_4;
input n_1;
input n_328;
input n_16;
input n_15;
input n_13;

output n_18;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_271;
wire n_47;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_0),
.B(n_29),
.Y(n_28)
);

INVx11_ASAP7_75t_L g35 ( 
.A(n_0),
.Y(n_35)
);

INVx5_ASAP7_75t_L g221 ( 
.A(n_0),
.Y(n_221)
);

AOI22xp33_ASAP7_75t_L g36 ( 
.A1(n_1),
.A2(n_29),
.B1(n_33),
.B2(n_37),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_1),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_1),
.A2(n_37),
.B1(n_42),
.B2(n_43),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g285 ( 
.A1(n_1),
.A2(n_37),
.B1(n_61),
.B2(n_62),
.Y(n_285)
);

AOI22xp33_ASAP7_75t_SL g320 ( 
.A1(n_1),
.A2(n_37),
.B1(n_54),
.B2(n_56),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_2),
.A2(n_54),
.B1(n_56),
.B2(n_65),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_2),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_2),
.A2(n_61),
.B1(n_62),
.B2(n_65),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_L g205 ( 
.A1(n_2),
.A2(n_29),
.B1(n_33),
.B2(n_65),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_2),
.A2(n_42),
.B1(n_43),
.B2(n_65),
.Y(n_237)
);

AOI22xp33_ASAP7_75t_L g48 ( 
.A1(n_3),
.A2(n_42),
.B1(n_43),
.B2(n_49),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_3),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_3),
.A2(n_29),
.B1(n_33),
.B2(n_49),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_3),
.A2(n_49),
.B1(n_61),
.B2(n_62),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g281 ( 
.A1(n_3),
.A2(n_49),
.B1(n_54),
.B2(n_56),
.Y(n_281)
);

BUFx12_ASAP7_75t_L g58 ( 
.A(n_4),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_5),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_6),
.Y(n_89)
);

AOI21xp33_ASAP7_75t_SL g90 ( 
.A1(n_6),
.A2(n_58),
.B(n_62),
.Y(n_90)
);

OAI22xp33_ASAP7_75t_SL g161 ( 
.A1(n_6),
.A2(n_54),
.B1(n_56),
.B2(n_89),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_6),
.B(n_60),
.Y(n_170)
);

AOI21xp5_ASAP7_75t_L g190 ( 
.A1(n_6),
.A2(n_43),
.B(n_191),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_6),
.B(n_43),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_6),
.B(n_78),
.Y(n_200)
);

OAI22xp33_ASAP7_75t_SL g220 ( 
.A1(n_6),
.A2(n_27),
.B1(n_217),
.B2(n_221),
.Y(n_220)
);

AOI21xp5_ASAP7_75t_L g232 ( 
.A1(n_6),
.A2(n_61),
.B(n_233),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_L g52 ( 
.A1(n_7),
.A2(n_53),
.B1(n_54),
.B2(n_56),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_7),
.Y(n_53)
);

OAI22xp33_ASAP7_75t_L g155 ( 
.A1(n_7),
.A2(n_53),
.B1(n_61),
.B2(n_62),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_SL g203 ( 
.A1(n_7),
.A2(n_42),
.B1(n_43),
.B2(n_53),
.Y(n_203)
);

AOI22xp33_ASAP7_75t_SL g211 ( 
.A1(n_7),
.A2(n_29),
.B1(n_33),
.B2(n_53),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g32 ( 
.A1(n_8),
.A2(n_29),
.B1(n_33),
.B2(n_34),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_8),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_L g104 ( 
.A1(n_8),
.A2(n_34),
.B1(n_42),
.B2(n_43),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_8),
.A2(n_34),
.B1(n_61),
.B2(n_62),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g296 ( 
.A1(n_8),
.A2(n_34),
.B1(n_54),
.B2(n_56),
.Y(n_296)
);

INVx13_ASAP7_75t_L g55 ( 
.A(n_9),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_10),
.A2(n_61),
.B1(n_62),
.B2(n_76),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_10),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_10),
.A2(n_54),
.B1(n_56),
.B2(n_76),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g159 ( 
.A1(n_10),
.A2(n_42),
.B1(n_43),
.B2(n_76),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_10),
.A2(n_29),
.B1(n_33),
.B2(n_76),
.Y(n_206)
);

OAI22xp33_ASAP7_75t_L g40 ( 
.A1(n_11),
.A2(n_41),
.B1(n_42),
.B2(n_43),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_11),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_11),
.A2(n_41),
.B1(n_61),
.B2(n_62),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_11),
.A2(n_41),
.B1(n_54),
.B2(n_56),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_11),
.A2(n_29),
.B1(n_33),
.B2(n_41),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g45 ( 
.A1(n_12),
.A2(n_29),
.B1(n_33),
.B2(n_46),
.Y(n_45)
);

INVx11_ASAP7_75t_L g46 ( 
.A(n_12),
.Y(n_46)
);

OAI22xp33_ASAP7_75t_L g47 ( 
.A1(n_12),
.A2(n_42),
.B1(n_43),
.B2(n_46),
.Y(n_47)
);

OAI32xp33_ASAP7_75t_L g194 ( 
.A1(n_12),
.A2(n_33),
.A3(n_43),
.B1(n_195),
.B2(n_196),
.Y(n_194)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_13),
.A2(n_29),
.B1(n_33),
.B2(n_102),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_13),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_13),
.A2(n_42),
.B1(n_43),
.B2(n_102),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g299 ( 
.A1(n_13),
.A2(n_61),
.B1(n_62),
.B2(n_102),
.Y(n_299)
);

BUFx24_ASAP7_75t_L g62 ( 
.A(n_14),
.Y(n_62)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_15),
.Y(n_70)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_15),
.Y(n_74)
);

INVx11_ASAP7_75t_SL g30 ( 
.A(n_16),
.Y(n_30)
);

OAI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_17),
.A2(n_54),
.B1(n_56),
.B2(n_84),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_17),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_L g167 ( 
.A1(n_17),
.A2(n_61),
.B1(n_62),
.B2(n_84),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_SL g192 ( 
.A1(n_17),
.A2(n_42),
.B1(n_43),
.B2(n_84),
.Y(n_192)
);

AOI22xp33_ASAP7_75t_SL g217 ( 
.A1(n_17),
.A2(n_29),
.B1(n_33),
.B2(n_84),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_308),
.Y(n_18)
);

OAI321xp33_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_276),
.A3(n_303),
.B1(n_306),
.B2(n_307),
.C(n_328),
.Y(n_19)
);

AOI321xp33_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_124),
.A3(n_147),
.B1(n_270),
.B2(n_275),
.C(n_329),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

OAI21xp5_ASAP7_75t_SL g270 ( 
.A1(n_22),
.A2(n_271),
.B(n_274),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_105),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_23),
.B(n_105),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_79),
.C(n_99),
.Y(n_23)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_24),
.B(n_99),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_SL g24 ( 
.A(n_25),
.B(n_50),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_25),
.B(n_51),
.C(n_66),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_38),
.Y(n_25)
);

XOR2xp5_ASAP7_75t_L g173 ( 
.A(n_26),
.B(n_38),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g26 ( 
.A1(n_27),
.A2(n_31),
.B1(n_35),
.B2(n_36),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_27),
.A2(n_36),
.B1(n_94),
.B2(n_101),
.Y(n_100)
);

AOI21xp5_ASAP7_75t_L g116 ( 
.A1(n_27),
.A2(n_94),
.B(n_101),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_27),
.A2(n_35),
.B1(n_205),
.B2(n_206),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_27),
.A2(n_35),
.B1(n_211),
.B2(n_217),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g244 ( 
.A1(n_27),
.A2(n_206),
.B1(n_245),
.B2(n_246),
.Y(n_244)
);

CKINVDCx14_ASAP7_75t_R g27 ( 
.A(n_28),
.Y(n_27)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_28),
.A2(n_32),
.B1(n_92),
.B2(n_93),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_28),
.A2(n_92),
.B1(n_95),
.B2(n_169),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_28),
.A2(n_95),
.B1(n_210),
.B2(n_212),
.Y(n_209)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_29),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_SL g196 ( 
.A(n_29),
.B(n_46),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_SL g222 ( 
.A(n_29),
.B(n_223),
.Y(n_222)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_32),
.Y(n_31)
);

INVx11_ASAP7_75t_L g95 ( 
.A(n_35),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_35),
.B(n_89),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_L g38 ( 
.A1(n_39),
.A2(n_44),
.B1(n_45),
.B2(n_48),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_40),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_40),
.A2(n_111),
.B1(n_114),
.B2(n_158),
.Y(n_157)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_42),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_42),
.A2(n_43),
.B1(n_70),
.B2(n_73),
.Y(n_72)
);

OAI32xp33_ASAP7_75t_L g241 ( 
.A1(n_42),
.A2(n_61),
.A3(n_73),
.B1(n_234),
.B2(n_242),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_SL g242 ( 
.A(n_43),
.B(n_243),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_44),
.A2(n_45),
.B1(n_48),
.B2(n_104),
.Y(n_103)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_44),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_44),
.A2(n_45),
.B1(n_113),
.B2(n_134),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_44),
.A2(n_45),
.B1(n_190),
.B2(n_192),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_44),
.A2(n_45),
.B1(n_192),
.B2(n_203),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_44),
.A2(n_45),
.B1(n_159),
.B2(n_260),
.Y(n_259)
);

AOI21xp5_ASAP7_75t_L g286 ( 
.A1(n_44),
.A2(n_45),
.B(n_134),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_SL g44 ( 
.A(n_45),
.B(n_47),
.Y(n_44)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_45),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g218 ( 
.A(n_45),
.B(n_89),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g50 ( 
.A(n_51),
.B(n_66),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g51 ( 
.A1(n_52),
.A2(n_57),
.B1(n_60),
.B2(n_64),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_52),
.Y(n_86)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_54),
.Y(n_56)
);

A2O1A1Ixp33_ASAP7_75t_L g88 ( 
.A1(n_54),
.A2(n_63),
.B(n_89),
.C(n_90),
.Y(n_88)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

O2A1O1Ixp33_ASAP7_75t_L g57 ( 
.A1(n_56),
.A2(n_58),
.B(n_59),
.C(n_60),
.Y(n_57)
);

NAND2xp33_ASAP7_75t_SL g59 ( 
.A(n_56),
.B(n_58),
.Y(n_59)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_57),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_57),
.A2(n_60),
.B1(n_64),
.B2(n_119),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_57),
.A2(n_60),
.B1(n_83),
.B2(n_161),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_57),
.A2(n_60),
.B1(n_295),
.B2(n_296),
.Y(n_294)
);

AO22x1_ASAP7_75t_L g60 ( 
.A1(n_58),
.A2(n_61),
.B1(n_62),
.B2(n_63),
.Y(n_60)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_58),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_60),
.Y(n_85)
);

A2O1A1Ixp33_ASAP7_75t_L g68 ( 
.A1(n_61),
.A2(n_69),
.B(n_71),
.C(n_72),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_61),
.B(n_69),
.Y(n_71)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_62),
.B(n_89),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_67),
.A2(n_75),
.B1(n_77),
.B2(n_78),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_67),
.A2(n_77),
.B1(n_78),
.B2(n_121),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_67),
.A2(n_78),
.B1(n_155),
.B2(n_166),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_67),
.A2(n_78),
.B1(n_284),
.B2(n_285),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_67),
.A2(n_78),
.B1(n_285),
.B2(n_299),
.Y(n_298)
);

CKINVDCx16_ASAP7_75t_R g67 ( 
.A(n_68),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_68),
.A2(n_72),
.B1(n_97),
.B2(n_98),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_68),
.A2(n_72),
.B1(n_131),
.B2(n_132),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_68),
.A2(n_72),
.B1(n_97),
.B2(n_154),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_68),
.A2(n_72),
.B1(n_167),
.B2(n_232),
.Y(n_231)
);

AOI21xp5_ASAP7_75t_L g315 ( 
.A1(n_68),
.A2(n_72),
.B(n_316),
.Y(n_315)
);

INVx1_ASAP7_75t_SL g69 ( 
.A(n_70),
.Y(n_69)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_72),
.Y(n_78)
);

INVx6_ASAP7_75t_L g243 ( 
.A(n_73),
.Y(n_243)
);

INVx8_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_75),
.Y(n_98)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_79),
.B(n_181),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_80),
.B(n_87),
.C(n_96),
.Y(n_79)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_80),
.B(n_96),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_81),
.A2(n_82),
.B1(n_85),
.B2(n_86),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_81),
.A2(n_85),
.B1(n_140),
.B2(n_141),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g280 ( 
.A1(n_81),
.A2(n_85),
.B1(n_141),
.B2(n_281),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_SL g318 ( 
.A1(n_81),
.A2(n_85),
.B1(n_319),
.B2(n_320),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_83),
.Y(n_82)
);

XNOR2xp5_ASAP7_75t_SL g175 ( 
.A(n_87),
.B(n_176),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_91),
.Y(n_87)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_88),
.B(n_91),
.Y(n_162)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx11_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx5_ASAP7_75t_SL g245 ( 
.A(n_95),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_103),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_100),
.B(n_103),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_104),
.Y(n_110)
);

XNOR2xp5_ASAP7_75t_L g105 ( 
.A(n_106),
.B(n_123),
.Y(n_105)
);

XNOR2xp5_ASAP7_75t_L g106 ( 
.A(n_107),
.B(n_117),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_107),
.B(n_117),
.C(n_123),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_108),
.A2(n_109),
.B1(n_115),
.B2(n_116),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_108),
.B(n_116),
.Y(n_143)
);

CKINVDCx16_ASAP7_75t_R g108 ( 
.A(n_109),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_110),
.A2(n_111),
.B1(n_112),
.B2(n_114),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_111),
.A2(n_114),
.B1(n_236),
.B2(n_237),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_113),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_115),
.A2(n_116),
.B1(n_138),
.B2(n_139),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_L g290 ( 
.A1(n_115),
.A2(n_139),
.B(n_142),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_116),
.Y(n_115)
);

BUFx24_ASAP7_75t_SL g327 ( 
.A(n_117),
.Y(n_327)
);

FAx1_ASAP7_75t_SL g117 ( 
.A(n_118),
.B(n_120),
.CI(n_122),
.CON(n_117),
.SN(n_117)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_118),
.B(n_120),
.C(n_122),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_119),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_121),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_126),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_125),
.B(n_126),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_127),
.A2(n_128),
.B1(n_145),
.B2(n_146),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

XOR2xp5_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_136),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_129),
.B(n_136),
.C(n_146),
.Y(n_304)
);

AOI21xp5_ASAP7_75t_L g129 ( 
.A1(n_130),
.A2(n_133),
.B(n_135),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_130),
.B(n_133),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_132),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_135),
.B(n_278),
.C(n_290),
.Y(n_277)
);

FAx1_ASAP7_75t_L g305 ( 
.A(n_135),
.B(n_278),
.CI(n_290),
.CON(n_305),
.SN(n_305)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_137),
.A2(n_142),
.B1(n_143),
.B2(n_144),
.Y(n_136)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_137),
.Y(n_144)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

CKINVDCx16_ASAP7_75t_R g146 ( 
.A(n_145),
.Y(n_146)
);

NOR3xp33_ASAP7_75t_SL g147 ( 
.A(n_148),
.B(n_177),
.C(n_182),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_171),
.Y(n_148)
);

AND2x2_ASAP7_75t_L g272 ( 
.A(n_149),
.B(n_171),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_162),
.C(n_163),
.Y(n_149)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_150),
.B(n_267),
.Y(n_266)
);

XOR2xp5_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_160),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_152),
.A2(n_153),
.B1(n_156),
.B2(n_157),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_152),
.B(n_157),
.C(n_160),
.Y(n_174)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_155),
.Y(n_154)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_159),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g267 ( 
.A1(n_162),
.A2(n_163),
.B1(n_164),
.B2(n_268),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_162),
.Y(n_268)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_168),
.C(n_170),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_165),
.B(n_255),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_167),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_168),
.B(n_170),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_169),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_175),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_173),
.B(n_174),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_173),
.B(n_174),
.C(n_175),
.Y(n_179)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

AOI21xp33_ASAP7_75t_L g271 ( 
.A1(n_178),
.A2(n_272),
.B(n_273),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_180),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_SL g273 ( 
.A(n_179),
.B(n_180),
.Y(n_273)
);

AOI21xp5_ASAP7_75t_L g182 ( 
.A1(n_183),
.A2(n_264),
.B(n_269),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_SL g183 ( 
.A1(n_184),
.A2(n_250),
.B(n_263),
.Y(n_183)
);

AOI21xp5_ASAP7_75t_L g184 ( 
.A1(n_185),
.A2(n_227),
.B(n_249),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_SL g185 ( 
.A1(n_186),
.A2(n_207),
.B(n_226),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_197),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_187),
.B(n_197),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_SL g187 ( 
.A(n_188),
.B(n_193),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_188),
.A2(n_189),
.B1(n_193),
.B2(n_194),
.Y(n_213)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

CKINVDCx16_ASAP7_75t_R g195 ( 
.A(n_191),
.Y(n_195)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_204),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_199),
.A2(n_200),
.B1(n_201),
.B2(n_202),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_199),
.B(n_202),
.C(n_204),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_200),
.Y(n_199)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_203),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_205),
.Y(n_212)
);

AOI21xp5_ASAP7_75t_L g207 ( 
.A1(n_208),
.A2(n_214),
.B(n_225),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_213),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_SL g225 ( 
.A(n_209),
.B(n_213),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_211),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_SL g214 ( 
.A1(n_215),
.A2(n_219),
.B(n_224),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_218),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_216),
.B(n_218),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_220),
.B(n_222),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_229),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_SL g249 ( 
.A(n_228),
.B(n_229),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_230),
.A2(n_240),
.B1(n_247),
.B2(n_248),
.Y(n_229)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_230),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_231),
.A2(n_235),
.B1(n_238),
.B2(n_239),
.Y(n_230)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_231),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_234),
.Y(n_233)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_235),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_235),
.B(n_239),
.C(n_248),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_237),
.Y(n_260)
);

CKINVDCx14_ASAP7_75t_R g248 ( 
.A(n_240),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_244),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_241),
.B(n_244),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_252),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_251),
.B(n_252),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_253),
.A2(n_254),
.B1(n_256),
.B2(n_257),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_253),
.B(n_259),
.C(n_261),
.Y(n_265)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_258),
.A2(n_259),
.B1(n_261),
.B2(n_262),
.Y(n_257)
);

CKINVDCx14_ASAP7_75t_R g261 ( 
.A(n_258),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_259),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_266),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_SL g269 ( 
.A(n_265),
.B(n_266),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_291),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_277),
.B(n_291),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_279),
.A2(n_280),
.B1(n_282),
.B2(n_289),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_279),
.A2(n_280),
.B1(n_293),
.B2(n_301),
.Y(n_292)
);

CKINVDCx14_ASAP7_75t_R g279 ( 
.A(n_280),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_280),
.B(n_283),
.C(n_288),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_280),
.B(n_301),
.C(n_302),
.Y(n_310)
);

INVxp67_ASAP7_75t_L g295 ( 
.A(n_281),
.Y(n_295)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_282),
.Y(n_289)
);

AOI22xp33_ASAP7_75t_L g282 ( 
.A1(n_283),
.A2(n_286),
.B1(n_287),
.B2(n_288),
.Y(n_282)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_283),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_286),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_286),
.A2(n_288),
.B1(n_298),
.B2(n_300),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_286),
.B(n_294),
.C(n_298),
.Y(n_322)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_292),
.B(n_302),
.Y(n_291)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_293),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_SL g293 ( 
.A(n_294),
.B(n_297),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_296),
.Y(n_319)
);

CKINVDCx16_ASAP7_75t_R g300 ( 
.A(n_298),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_299),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_304),
.B(n_305),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_SL g306 ( 
.A(n_304),
.B(n_305),
.Y(n_306)
);

BUFx24_ASAP7_75t_SL g326 ( 
.A(n_305),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_309),
.B(n_323),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_310),
.B(n_311),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_310),
.B(n_311),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_312),
.A2(n_313),
.B1(n_321),
.B2(n_322),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_314),
.A2(n_315),
.B1(n_317),
.B2(n_318),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_315),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_318),
.Y(n_317)
);

CKINVDCx16_ASAP7_75t_R g321 ( 
.A(n_322),
.Y(n_321)
);

INVxp67_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);


endmodule