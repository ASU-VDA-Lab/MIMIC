module fake_netlist_6_1208_n_1805 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_193, n_147, n_154, n_191, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_166, n_28, n_184, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_188, n_102, n_186, n_0, n_87, n_189, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_104, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_190, n_14, n_123, n_136, n_72, n_187, n_89, n_173, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_171, n_31, n_192, n_57, n_169, n_53, n_51, n_44, n_56, n_1805);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_193;
input n_147;
input n_154;
input n_191;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_184;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_188;
input n_102;
input n_186;
input n_0;
input n_87;
input n_189;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_104;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_190;
input n_14;
input n_123;
input n_136;
input n_72;
input n_187;
input n_89;
input n_173;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_171;
input n_31;
input n_192;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1805;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_1738;
wire n_798;
wire n_1575;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1688;
wire n_1691;
wire n_1009;
wire n_1743;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1803;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1704;
wire n_1078;
wire n_250;
wire n_544;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_616;
wire n_658;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1620;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1644;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1697;
wire n_243;
wire n_979;
wire n_905;
wire n_1680;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_210;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1747;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1802;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1801;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_697;
wire n_687;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_484;
wire n_1709;
wire n_1757;
wire n_1796;
wire n_1792;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_297;
wire n_595;
wire n_627;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_1788;
wire n_622;
wire n_1469;
wire n_1766;
wire n_1776;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_899;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1577;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_927;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_552;
wire n_1358;
wire n_1388;
wire n_216;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_1021;
wire n_931;
wire n_474;
wire n_527;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_211;
wire n_1483;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1769;
wire n_1220;
wire n_556;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_1286;
wire n_1773;
wire n_1775;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_1745;
wire n_914;
wire n_759;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1135;
wire n_1179;
wire n_1169;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1267;
wire n_1281;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1024;
wire n_1768;
wire n_198;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1361;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_1695;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_227;
wire n_1720;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_959;
wire n_879;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_1676;
wire n_833;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_1758;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1559;
wire n_1725;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1741;
wire n_1325;
wire n_1002;
wire n_1746;
wire n_545;
wire n_489;
wire n_1804;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1800;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1118;
wire n_1076;
wire n_194;
wire n_1007;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1631;
wire n_591;
wire n_1377;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_1729;
wire n_669;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1785;
wire n_763;
wire n_1147;
wire n_360;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_363;
wire n_1799;
wire n_1090;
wire n_592;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_271;
wire n_404;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_373;
wire n_1632;
wire n_257;
wire n_1557;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_207;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

INVx1_ASAP7_75t_L g194 ( 
.A(n_91),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_39),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_60),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_107),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_46),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_25),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_15),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_53),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_85),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_190),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_110),
.Y(n_204)
);

BUFx3_ASAP7_75t_L g205 ( 
.A(n_157),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_145),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_36),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_16),
.Y(n_208)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_60),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_192),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_193),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_33),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_168),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_45),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_129),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_56),
.Y(n_216)
);

BUFx3_ASAP7_75t_L g217 ( 
.A(n_15),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_78),
.Y(n_218)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_3),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_127),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_84),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_70),
.Y(n_222)
);

INVx1_ASAP7_75t_SL g223 ( 
.A(n_63),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_179),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_164),
.Y(n_225)
);

BUFx3_ASAP7_75t_L g226 ( 
.A(n_130),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_79),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_47),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_163),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_37),
.Y(n_230)
);

INVx2_ASAP7_75t_SL g231 ( 
.A(n_172),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_38),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_29),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_89),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_94),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_140),
.Y(n_236)
);

BUFx6f_ASAP7_75t_L g237 ( 
.A(n_161),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_62),
.Y(n_238)
);

BUFx2_ASAP7_75t_L g239 ( 
.A(n_125),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_53),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_111),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_66),
.Y(n_242)
);

BUFx6f_ASAP7_75t_L g243 ( 
.A(n_171),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_58),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_175),
.Y(n_245)
);

INVxp67_ASAP7_75t_L g246 ( 
.A(n_87),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_184),
.Y(n_247)
);

INVx2_ASAP7_75t_SL g248 ( 
.A(n_77),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_72),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_112),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_141),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_21),
.Y(n_252)
);

CKINVDCx16_ASAP7_75t_R g253 ( 
.A(n_38),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_40),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_155),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_162),
.Y(n_256)
);

INVx3_ASAP7_75t_L g257 ( 
.A(n_143),
.Y(n_257)
);

BUFx3_ASAP7_75t_L g258 ( 
.A(n_158),
.Y(n_258)
);

CKINVDCx14_ASAP7_75t_R g259 ( 
.A(n_154),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_1),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_80),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_136),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_36),
.Y(n_263)
);

BUFx6f_ASAP7_75t_L g264 ( 
.A(n_151),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_76),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_115),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_32),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_5),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_88),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_65),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_103),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_169),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_50),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_101),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_34),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_152),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_27),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_122),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_108),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_160),
.Y(n_280)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_4),
.Y(n_281)
);

INVx1_ASAP7_75t_SL g282 ( 
.A(n_58),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_55),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_86),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_186),
.Y(n_285)
);

INVx2_ASAP7_75t_SL g286 ( 
.A(n_12),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_37),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_106),
.Y(n_288)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_12),
.Y(n_289)
);

BUFx3_ASAP7_75t_L g290 ( 
.A(n_68),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_46),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_149),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_7),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_64),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_75),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_177),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_61),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_174),
.Y(n_298)
);

BUFx2_ASAP7_75t_L g299 ( 
.A(n_97),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_166),
.Y(n_300)
);

INVx1_ASAP7_75t_SL g301 ( 
.A(n_61),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_43),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_183),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_24),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_1),
.Y(n_305)
);

INVxp67_ASAP7_75t_L g306 ( 
.A(n_7),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_81),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_188),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_181),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_3),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_132),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_31),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_133),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_131),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_2),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_99),
.Y(n_316)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_134),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_43),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_180),
.Y(n_319)
);

CKINVDCx14_ASAP7_75t_R g320 ( 
.A(n_142),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_23),
.Y(n_321)
);

BUFx6f_ASAP7_75t_L g322 ( 
.A(n_51),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_173),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_144),
.Y(n_324)
);

CKINVDCx16_ASAP7_75t_R g325 ( 
.A(n_13),
.Y(n_325)
);

BUFx3_ASAP7_75t_L g326 ( 
.A(n_128),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_20),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_4),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_54),
.Y(n_329)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_6),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_73),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_123),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_26),
.Y(n_333)
);

INVx2_ASAP7_75t_L g334 ( 
.A(n_13),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_67),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_14),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_187),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_19),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g339 ( 
.A(n_21),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_153),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_30),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_147),
.Y(n_342)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_9),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_167),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_116),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_191),
.Y(n_346)
);

INVx3_ASAP7_75t_L g347 ( 
.A(n_20),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_48),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_69),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_47),
.Y(n_350)
);

BUFx5_ASAP7_75t_L g351 ( 
.A(n_182),
.Y(n_351)
);

CKINVDCx16_ASAP7_75t_R g352 ( 
.A(n_105),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_5),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_29),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_9),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_14),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_8),
.Y(n_357)
);

INVx1_ASAP7_75t_SL g358 ( 
.A(n_82),
.Y(n_358)
);

INVx2_ASAP7_75t_L g359 ( 
.A(n_124),
.Y(n_359)
);

INVx2_ASAP7_75t_SL g360 ( 
.A(n_42),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_178),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_34),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_159),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_48),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_92),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_52),
.Y(n_366)
);

CKINVDCx20_ASAP7_75t_R g367 ( 
.A(n_11),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_19),
.Y(n_368)
);

INVx2_ASAP7_75t_SL g369 ( 
.A(n_95),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_176),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_28),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_114),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_22),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_135),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_10),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_24),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_6),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_148),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_138),
.Y(n_379)
);

BUFx2_ASAP7_75t_L g380 ( 
.A(n_22),
.Y(n_380)
);

CKINVDCx16_ASAP7_75t_R g381 ( 
.A(n_44),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_49),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_57),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_146),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_L g385 ( 
.A(n_239),
.B(n_0),
.Y(n_385)
);

CKINVDCx20_ASAP7_75t_R g386 ( 
.A(n_220),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_L g387 ( 
.A(n_299),
.B(n_0),
.Y(n_387)
);

BUFx3_ASAP7_75t_L g388 ( 
.A(n_205),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_347),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_253),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_231),
.B(n_2),
.Y(n_391)
);

INVxp67_ASAP7_75t_SL g392 ( 
.A(n_347),
.Y(n_392)
);

NOR2xp67_ASAP7_75t_L g393 ( 
.A(n_347),
.B(n_8),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_325),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_217),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_217),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_322),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_322),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_381),
.Y(n_399)
);

CKINVDCx20_ASAP7_75t_R g400 ( 
.A(n_265),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_322),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_254),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_322),
.Y(n_403)
);

NOR2xp67_ASAP7_75t_L g404 ( 
.A(n_257),
.B(n_11),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_322),
.Y(n_405)
);

CKINVDCx20_ASAP7_75t_R g406 ( 
.A(n_271),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_268),
.Y(n_407)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_351),
.Y(n_408)
);

CKINVDCx20_ASAP7_75t_R g409 ( 
.A(n_272),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_198),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_209),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_209),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_200),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_212),
.Y(n_414)
);

CKINVDCx20_ASAP7_75t_R g415 ( 
.A(n_309),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_232),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_244),
.Y(n_417)
);

CKINVDCx20_ASAP7_75t_R g418 ( 
.A(n_319),
.Y(n_418)
);

CKINVDCx20_ASAP7_75t_R g419 ( 
.A(n_352),
.Y(n_419)
);

INVxp67_ASAP7_75t_L g420 ( 
.A(n_380),
.Y(n_420)
);

CKINVDCx20_ASAP7_75t_R g421 ( 
.A(n_259),
.Y(n_421)
);

CKINVDCx20_ASAP7_75t_R g422 ( 
.A(n_320),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_260),
.Y(n_423)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_351),
.Y(n_424)
);

NOR2xp67_ASAP7_75t_L g425 ( 
.A(n_257),
.B(n_16),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_263),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_275),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_277),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_267),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_287),
.Y(n_430)
);

INVxp67_ASAP7_75t_SL g431 ( 
.A(n_205),
.Y(n_431)
);

INVxp67_ASAP7_75t_L g432 ( 
.A(n_291),
.Y(n_432)
);

CKINVDCx16_ASAP7_75t_R g433 ( 
.A(n_195),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_318),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_293),
.Y(n_435)
);

CKINVDCx20_ASAP7_75t_R g436 ( 
.A(n_236),
.Y(n_436)
);

NOR2xp67_ASAP7_75t_L g437 ( 
.A(n_257),
.B(n_17),
.Y(n_437)
);

CKINVDCx20_ASAP7_75t_R g438 ( 
.A(n_238),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_302),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_327),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_304),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_328),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_305),
.Y(n_443)
);

INVxp33_ASAP7_75t_SL g444 ( 
.A(n_196),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_333),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_310),
.Y(n_446)
);

NOR2xp33_ASAP7_75t_R g447 ( 
.A(n_241),
.B(n_83),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_348),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_315),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_321),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_329),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_336),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_338),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_341),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_350),
.Y(n_455)
);

INVxp33_ASAP7_75t_SL g456 ( 
.A(n_196),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_364),
.Y(n_457)
);

INVxp67_ASAP7_75t_SL g458 ( 
.A(n_226),
.Y(n_458)
);

CKINVDCx20_ASAP7_75t_R g459 ( 
.A(n_245),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_371),
.Y(n_460)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_351),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_373),
.Y(n_462)
);

INVx4_ASAP7_75t_R g463 ( 
.A(n_226),
.Y(n_463)
);

INVxp67_ASAP7_75t_SL g464 ( 
.A(n_258),
.Y(n_464)
);

CKINVDCx5p33_ASAP7_75t_R g465 ( 
.A(n_199),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_375),
.Y(n_466)
);

NOR2xp33_ASAP7_75t_L g467 ( 
.A(n_231),
.B(n_17),
.Y(n_467)
);

NOR2xp33_ASAP7_75t_L g468 ( 
.A(n_248),
.B(n_18),
.Y(n_468)
);

CKINVDCx14_ASAP7_75t_R g469 ( 
.A(n_258),
.Y(n_469)
);

NOR2xp33_ASAP7_75t_L g470 ( 
.A(n_248),
.B(n_18),
.Y(n_470)
);

CKINVDCx20_ASAP7_75t_R g471 ( 
.A(n_247),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_382),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_290),
.Y(n_473)
);

INVxp67_ASAP7_75t_L g474 ( 
.A(n_199),
.Y(n_474)
);

CKINVDCx20_ASAP7_75t_R g475 ( 
.A(n_250),
.Y(n_475)
);

CKINVDCx5p33_ASAP7_75t_R g476 ( 
.A(n_201),
.Y(n_476)
);

CKINVDCx20_ASAP7_75t_R g477 ( 
.A(n_251),
.Y(n_477)
);

NOR2xp67_ASAP7_75t_L g478 ( 
.A(n_306),
.B(n_25),
.Y(n_478)
);

INVxp67_ASAP7_75t_SL g479 ( 
.A(n_290),
.Y(n_479)
);

XOR2xp5_ASAP7_75t_L g480 ( 
.A(n_240),
.B(n_26),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_326),
.Y(n_481)
);

CKINVDCx5p33_ASAP7_75t_R g482 ( 
.A(n_201),
.Y(n_482)
);

CKINVDCx5p33_ASAP7_75t_R g483 ( 
.A(n_207),
.Y(n_483)
);

AND2x4_ASAP7_75t_L g484 ( 
.A(n_392),
.B(n_326),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_397),
.Y(n_485)
);

INVx2_ASAP7_75t_L g486 ( 
.A(n_398),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_SL g487 ( 
.A(n_421),
.B(n_369),
.Y(n_487)
);

BUFx6f_ASAP7_75t_L g488 ( 
.A(n_401),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_403),
.Y(n_489)
);

CKINVDCx5p33_ASAP7_75t_R g490 ( 
.A(n_436),
.Y(n_490)
);

XNOR2xp5_ASAP7_75t_L g491 ( 
.A(n_480),
.B(n_252),
.Y(n_491)
);

NOR2xp33_ASAP7_75t_R g492 ( 
.A(n_469),
.B(n_256),
.Y(n_492)
);

NOR2xp33_ASAP7_75t_R g493 ( 
.A(n_422),
.B(n_262),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_405),
.Y(n_494)
);

CKINVDCx20_ASAP7_75t_R g495 ( 
.A(n_386),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_389),
.Y(n_496)
);

INVxp67_ASAP7_75t_L g497 ( 
.A(n_390),
.Y(n_497)
);

CKINVDCx5p33_ASAP7_75t_R g498 ( 
.A(n_438),
.Y(n_498)
);

CKINVDCx8_ASAP7_75t_R g499 ( 
.A(n_433),
.Y(n_499)
);

INVx3_ASAP7_75t_L g500 ( 
.A(n_408),
.Y(n_500)
);

BUFx2_ASAP7_75t_L g501 ( 
.A(n_394),
.Y(n_501)
);

CKINVDCx5p33_ASAP7_75t_R g502 ( 
.A(n_459),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_410),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_413),
.Y(n_504)
);

CKINVDCx5p33_ASAP7_75t_R g505 ( 
.A(n_471),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_414),
.Y(n_506)
);

INVx2_ASAP7_75t_L g507 ( 
.A(n_408),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_424),
.Y(n_508)
);

CKINVDCx5p33_ASAP7_75t_R g509 ( 
.A(n_475),
.Y(n_509)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_424),
.Y(n_510)
);

AOI22x1_ASAP7_75t_SL g511 ( 
.A1(n_400),
.A2(n_297),
.B1(n_312),
.B2(n_339),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_416),
.Y(n_512)
);

AND2x2_ASAP7_75t_L g513 ( 
.A(n_431),
.B(n_286),
.Y(n_513)
);

BUFx6f_ASAP7_75t_L g514 ( 
.A(n_461),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_417),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_458),
.B(n_464),
.Y(n_516)
);

NOR2xp33_ASAP7_75t_L g517 ( 
.A(n_391),
.B(n_369),
.Y(n_517)
);

HB1xp67_ASAP7_75t_L g518 ( 
.A(n_394),
.Y(n_518)
);

CKINVDCx5p33_ASAP7_75t_R g519 ( 
.A(n_477),
.Y(n_519)
);

HB1xp67_ASAP7_75t_L g520 ( 
.A(n_399),
.Y(n_520)
);

CKINVDCx5p33_ASAP7_75t_R g521 ( 
.A(n_419),
.Y(n_521)
);

NOR2xp33_ASAP7_75t_R g522 ( 
.A(n_402),
.B(n_266),
.Y(n_522)
);

INVx2_ASAP7_75t_L g523 ( 
.A(n_461),
.Y(n_523)
);

NOR2xp67_ASAP7_75t_L g524 ( 
.A(n_474),
.B(n_246),
.Y(n_524)
);

CKINVDCx5p33_ASAP7_75t_R g525 ( 
.A(n_406),
.Y(n_525)
);

CKINVDCx5p33_ASAP7_75t_R g526 ( 
.A(n_409),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_423),
.Y(n_527)
);

CKINVDCx20_ASAP7_75t_R g528 ( 
.A(n_415),
.Y(n_528)
);

CKINVDCx5p33_ASAP7_75t_R g529 ( 
.A(n_418),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_479),
.B(n_317),
.Y(n_530)
);

CKINVDCx5p33_ASAP7_75t_R g531 ( 
.A(n_402),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_388),
.B(n_317),
.Y(n_532)
);

CKINVDCx5p33_ASAP7_75t_R g533 ( 
.A(n_407),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_426),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_429),
.Y(n_535)
);

AND2x4_ASAP7_75t_L g536 ( 
.A(n_393),
.B(n_359),
.Y(n_536)
);

CKINVDCx5p33_ASAP7_75t_R g537 ( 
.A(n_407),
.Y(n_537)
);

INVx2_ASAP7_75t_L g538 ( 
.A(n_411),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_430),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_434),
.Y(n_540)
);

CKINVDCx5p33_ASAP7_75t_R g541 ( 
.A(n_427),
.Y(n_541)
);

BUFx6f_ASAP7_75t_L g542 ( 
.A(n_411),
.Y(n_542)
);

BUFx6f_ASAP7_75t_L g543 ( 
.A(n_412),
.Y(n_543)
);

INVx2_ASAP7_75t_L g544 ( 
.A(n_412),
.Y(n_544)
);

CKINVDCx5p33_ASAP7_75t_R g545 ( 
.A(n_427),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_L g546 ( 
.A(n_388),
.B(n_359),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_440),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_442),
.Y(n_548)
);

AND2x4_ASAP7_75t_L g549 ( 
.A(n_404),
.B(n_425),
.Y(n_549)
);

CKINVDCx5p33_ASAP7_75t_R g550 ( 
.A(n_428),
.Y(n_550)
);

HB1xp67_ASAP7_75t_L g551 ( 
.A(n_399),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_L g552 ( 
.A(n_473),
.B(n_194),
.Y(n_552)
);

OAI22xp5_ASAP7_75t_L g553 ( 
.A1(n_420),
.A2(n_456),
.B1(n_444),
.B2(n_465),
.Y(n_553)
);

NOR2xp33_ASAP7_75t_SL g554 ( 
.A(n_385),
.B(n_223),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_L g555 ( 
.A(n_481),
.B(n_202),
.Y(n_555)
);

BUFx6f_ASAP7_75t_L g556 ( 
.A(n_445),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_L g557 ( 
.A(n_395),
.B(n_210),
.Y(n_557)
);

BUFx6f_ASAP7_75t_L g558 ( 
.A(n_448),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_SL g559 ( 
.A(n_428),
.B(n_197),
.Y(n_559)
);

BUFx6f_ASAP7_75t_L g560 ( 
.A(n_455),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_457),
.Y(n_561)
);

CKINVDCx5p33_ASAP7_75t_R g562 ( 
.A(n_435),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_SL g563 ( 
.A(n_554),
.B(n_437),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_503),
.Y(n_564)
);

NOR2xp33_ASAP7_75t_L g565 ( 
.A(n_516),
.B(n_517),
.Y(n_565)
);

NOR2xp33_ASAP7_75t_L g566 ( 
.A(n_484),
.B(n_444),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_486),
.Y(n_567)
);

INVx2_ASAP7_75t_SL g568 ( 
.A(n_522),
.Y(n_568)
);

AND2x4_ASAP7_75t_L g569 ( 
.A(n_484),
.B(n_460),
.Y(n_569)
);

AOI22xp5_ASAP7_75t_L g570 ( 
.A1(n_553),
.A2(n_387),
.B1(n_452),
.B2(n_451),
.Y(n_570)
);

BUFx6f_ASAP7_75t_L g571 ( 
.A(n_514),
.Y(n_571)
);

INVxp67_ASAP7_75t_L g572 ( 
.A(n_501),
.Y(n_572)
);

INVx5_ASAP7_75t_L g573 ( 
.A(n_514),
.Y(n_573)
);

AND2x2_ASAP7_75t_L g574 ( 
.A(n_513),
.B(n_435),
.Y(n_574)
);

INVx2_ASAP7_75t_L g575 ( 
.A(n_486),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_504),
.Y(n_576)
);

AOI22xp33_ASAP7_75t_L g577 ( 
.A1(n_536),
.A2(n_468),
.B1(n_467),
.B2(n_470),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_507),
.Y(n_578)
);

INVx3_ASAP7_75t_L g579 ( 
.A(n_500),
.Y(n_579)
);

OR2x2_ASAP7_75t_L g580 ( 
.A(n_484),
.B(n_465),
.Y(n_580)
);

INVx2_ASAP7_75t_SL g581 ( 
.A(n_549),
.Y(n_581)
);

HB1xp67_ASAP7_75t_L g582 ( 
.A(n_524),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_506),
.Y(n_583)
);

NOR2xp33_ASAP7_75t_L g584 ( 
.A(n_530),
.B(n_456),
.Y(n_584)
);

HB1xp67_ASAP7_75t_L g585 ( 
.A(n_518),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_SL g586 ( 
.A(n_536),
.B(n_237),
.Y(n_586)
);

INVx6_ASAP7_75t_L g587 ( 
.A(n_536),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_SL g588 ( 
.A(n_556),
.B(n_237),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_SL g589 ( 
.A(n_556),
.B(n_237),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_512),
.Y(n_590)
);

AND2x4_ASAP7_75t_L g591 ( 
.A(n_496),
.B(n_462),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_515),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_527),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_534),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_507),
.Y(n_595)
);

INVx2_ASAP7_75t_L g596 ( 
.A(n_508),
.Y(n_596)
);

INVx4_ASAP7_75t_L g597 ( 
.A(n_514),
.Y(n_597)
);

AND2x2_ASAP7_75t_L g598 ( 
.A(n_497),
.B(n_439),
.Y(n_598)
);

NOR2xp33_ASAP7_75t_L g599 ( 
.A(n_559),
.B(n_441),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_SL g600 ( 
.A(n_556),
.B(n_237),
.Y(n_600)
);

CKINVDCx5p33_ASAP7_75t_R g601 ( 
.A(n_493),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_535),
.Y(n_602)
);

BUFx3_ASAP7_75t_L g603 ( 
.A(n_539),
.Y(n_603)
);

CKINVDCx6p67_ASAP7_75t_R g604 ( 
.A(n_495),
.Y(n_604)
);

NOR2x1p5_ASAP7_75t_L g605 ( 
.A(n_531),
.B(n_476),
.Y(n_605)
);

INVx4_ASAP7_75t_L g606 ( 
.A(n_514),
.Y(n_606)
);

INVx4_ASAP7_75t_L g607 ( 
.A(n_514),
.Y(n_607)
);

NOR2xp33_ASAP7_75t_L g608 ( 
.A(n_532),
.B(n_441),
.Y(n_608)
);

AOI22xp5_ASAP7_75t_L g609 ( 
.A1(n_487),
.A2(n_452),
.B1(n_446),
.B2(n_449),
.Y(n_609)
);

INVx4_ASAP7_75t_L g610 ( 
.A(n_488),
.Y(n_610)
);

BUFx2_ASAP7_75t_L g611 ( 
.A(n_501),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_SL g612 ( 
.A(n_556),
.B(n_237),
.Y(n_612)
);

AND2x4_ASAP7_75t_L g613 ( 
.A(n_540),
.B(n_466),
.Y(n_613)
);

NAND3xp33_ASAP7_75t_L g614 ( 
.A(n_546),
.B(n_446),
.C(n_443),
.Y(n_614)
);

AND2x2_ASAP7_75t_L g615 ( 
.A(n_492),
.B(n_443),
.Y(n_615)
);

BUFx4f_ASAP7_75t_L g616 ( 
.A(n_556),
.Y(n_616)
);

BUFx6f_ASAP7_75t_L g617 ( 
.A(n_558),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_547),
.Y(n_618)
);

INVx4_ASAP7_75t_L g619 ( 
.A(n_488),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_548),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_L g621 ( 
.A(n_485),
.B(n_489),
.Y(n_621)
);

BUFx3_ASAP7_75t_L g622 ( 
.A(n_561),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_494),
.Y(n_623)
);

INVx5_ASAP7_75t_L g624 ( 
.A(n_488),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_558),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_L g626 ( 
.A(n_500),
.B(n_510),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_SL g627 ( 
.A(n_558),
.B(n_243),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_558),
.Y(n_628)
);

BUFx6f_ASAP7_75t_L g629 ( 
.A(n_558),
.Y(n_629)
);

CKINVDCx16_ASAP7_75t_R g630 ( 
.A(n_528),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_L g631 ( 
.A(n_510),
.B(n_449),
.Y(n_631)
);

BUFx4f_ASAP7_75t_L g632 ( 
.A(n_560),
.Y(n_632)
);

AND2x2_ASAP7_75t_L g633 ( 
.A(n_531),
.B(n_450),
.Y(n_633)
);

INVx3_ASAP7_75t_L g634 ( 
.A(n_488),
.Y(n_634)
);

INVx2_ASAP7_75t_L g635 ( 
.A(n_523),
.Y(n_635)
);

BUFx3_ASAP7_75t_L g636 ( 
.A(n_560),
.Y(n_636)
);

NOR2xp33_ASAP7_75t_L g637 ( 
.A(n_552),
.B(n_450),
.Y(n_637)
);

AOI22xp5_ASAP7_75t_L g638 ( 
.A1(n_533),
.A2(n_454),
.B1(n_453),
.B2(n_451),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_560),
.Y(n_639)
);

BUFx6f_ASAP7_75t_L g640 ( 
.A(n_560),
.Y(n_640)
);

INVx2_ASAP7_75t_SL g641 ( 
.A(n_520),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_560),
.Y(n_642)
);

OR2x2_ASAP7_75t_SL g643 ( 
.A(n_551),
.B(n_219),
.Y(n_643)
);

OAI21xp33_ASAP7_75t_SL g644 ( 
.A1(n_555),
.A2(n_478),
.B(n_360),
.Y(n_644)
);

INVx2_ASAP7_75t_SL g645 ( 
.A(n_533),
.Y(n_645)
);

AOI22xp33_ASAP7_75t_L g646 ( 
.A1(n_557),
.A2(n_219),
.B1(n_343),
.B2(n_334),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_SL g647 ( 
.A(n_537),
.B(n_243),
.Y(n_647)
);

INVx2_ASAP7_75t_SL g648 ( 
.A(n_537),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_523),
.B(n_453),
.Y(n_649)
);

INVx3_ASAP7_75t_L g650 ( 
.A(n_488),
.Y(n_650)
);

INVx2_ASAP7_75t_L g651 ( 
.A(n_542),
.Y(n_651)
);

NAND2xp33_ASAP7_75t_R g652 ( 
.A(n_541),
.B(n_476),
.Y(n_652)
);

AND2x6_ASAP7_75t_L g653 ( 
.A(n_538),
.B(n_243),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_542),
.Y(n_654)
);

INVx3_ASAP7_75t_L g655 ( 
.A(n_542),
.Y(n_655)
);

BUFx6f_ASAP7_75t_L g656 ( 
.A(n_542),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_SL g657 ( 
.A(n_541),
.B(n_243),
.Y(n_657)
);

AOI22xp5_ASAP7_75t_L g658 ( 
.A1(n_545),
.A2(n_454),
.B1(n_483),
.B2(n_482),
.Y(n_658)
);

BUFx4f_ASAP7_75t_L g659 ( 
.A(n_542),
.Y(n_659)
);

NAND3xp33_ASAP7_75t_L g660 ( 
.A(n_545),
.B(n_483),
.C(n_482),
.Y(n_660)
);

NOR2xp33_ASAP7_75t_L g661 ( 
.A(n_550),
.B(n_396),
.Y(n_661)
);

AOI22xp33_ASAP7_75t_L g662 ( 
.A1(n_538),
.A2(n_289),
.B1(n_343),
.B2(n_281),
.Y(n_662)
);

NOR2xp33_ASAP7_75t_L g663 ( 
.A(n_550),
.B(n_432),
.Y(n_663)
);

AND2x4_ASAP7_75t_L g664 ( 
.A(n_544),
.B(n_472),
.Y(n_664)
);

AOI22xp33_ASAP7_75t_L g665 ( 
.A1(n_544),
.A2(n_289),
.B1(n_334),
.B2(n_330),
.Y(n_665)
);

BUFx6f_ASAP7_75t_L g666 ( 
.A(n_543),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_L g667 ( 
.A(n_543),
.B(n_358),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_SL g668 ( 
.A(n_562),
.B(n_243),
.Y(n_668)
);

INVx4_ASAP7_75t_L g669 ( 
.A(n_543),
.Y(n_669)
);

BUFx3_ASAP7_75t_L g670 ( 
.A(n_543),
.Y(n_670)
);

INVx2_ASAP7_75t_L g671 ( 
.A(n_543),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_SL g672 ( 
.A(n_562),
.B(n_264),
.Y(n_672)
);

AOI22xp33_ASAP7_75t_L g673 ( 
.A1(n_491),
.A2(n_281),
.B1(n_330),
.B2(n_286),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_SL g674 ( 
.A(n_499),
.B(n_264),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_499),
.Y(n_675)
);

INVx4_ASAP7_75t_L g676 ( 
.A(n_490),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_490),
.B(n_269),
.Y(n_677)
);

BUFx10_ASAP7_75t_L g678 ( 
.A(n_521),
.Y(n_678)
);

AND2x2_ASAP7_75t_L g679 ( 
.A(n_498),
.B(n_282),
.Y(n_679)
);

INVx2_ASAP7_75t_L g680 ( 
.A(n_498),
.Y(n_680)
);

NOR2xp33_ASAP7_75t_L g681 ( 
.A(n_502),
.B(n_360),
.Y(n_681)
);

INVx2_ASAP7_75t_L g682 ( 
.A(n_502),
.Y(n_682)
);

AOI22xp33_ASAP7_75t_L g683 ( 
.A1(n_491),
.A2(n_264),
.B1(n_384),
.B2(n_235),
.Y(n_683)
);

AND2x2_ASAP7_75t_L g684 ( 
.A(n_505),
.B(n_301),
.Y(n_684)
);

AND2x2_ASAP7_75t_L g685 ( 
.A(n_509),
.B(n_208),
.Y(n_685)
);

INVx2_ASAP7_75t_L g686 ( 
.A(n_509),
.Y(n_686)
);

AOI22xp33_ASAP7_75t_L g687 ( 
.A1(n_519),
.A2(n_264),
.B1(n_300),
.B2(n_276),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_519),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_525),
.Y(n_689)
);

INVx5_ASAP7_75t_L g690 ( 
.A(n_511),
.Y(n_690)
);

NOR2xp33_ASAP7_75t_L g691 ( 
.A(n_525),
.B(n_197),
.Y(n_691)
);

INVx3_ASAP7_75t_L g692 ( 
.A(n_526),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_526),
.Y(n_693)
);

NOR2xp33_ASAP7_75t_L g694 ( 
.A(n_529),
.B(n_203),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_529),
.Y(n_695)
);

INVx5_ASAP7_75t_L g696 ( 
.A(n_511),
.Y(n_696)
);

INVx6_ASAP7_75t_L g697 ( 
.A(n_484),
.Y(n_697)
);

AND2x6_ASAP7_75t_L g698 ( 
.A(n_517),
.B(n_264),
.Y(n_698)
);

CKINVDCx5p33_ASAP7_75t_R g699 ( 
.A(n_493),
.Y(n_699)
);

BUFx8_ASAP7_75t_SL g700 ( 
.A(n_495),
.Y(n_700)
);

INVx4_ASAP7_75t_L g701 ( 
.A(n_514),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_503),
.Y(n_702)
);

INVxp33_ASAP7_75t_L g703 ( 
.A(n_513),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_L g704 ( 
.A(n_565),
.B(n_211),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_L g705 ( 
.A(n_565),
.B(n_225),
.Y(n_705)
);

AOI22xp5_ASAP7_75t_L g706 ( 
.A1(n_566),
.A2(n_584),
.B1(n_697),
.B2(n_637),
.Y(n_706)
);

BUFx3_ASAP7_75t_L g707 ( 
.A(n_697),
.Y(n_707)
);

NAND2xp33_ASAP7_75t_L g708 ( 
.A(n_698),
.B(n_351),
.Y(n_708)
);

OAI21xp5_ASAP7_75t_L g709 ( 
.A1(n_703),
.A2(n_249),
.B(n_242),
.Y(n_709)
);

NOR2xp33_ASAP7_75t_L g710 ( 
.A(n_703),
.B(n_203),
.Y(n_710)
);

AND2x2_ASAP7_75t_L g711 ( 
.A(n_574),
.B(n_480),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_L g712 ( 
.A(n_697),
.B(n_255),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_564),
.Y(n_713)
);

INVx2_ASAP7_75t_L g714 ( 
.A(n_579),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_SL g715 ( 
.A(n_637),
.B(n_204),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_576),
.Y(n_716)
);

NOR2xp33_ASAP7_75t_L g717 ( 
.A(n_584),
.B(n_204),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_L g718 ( 
.A(n_608),
.B(n_261),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_583),
.Y(n_719)
);

INVx2_ASAP7_75t_L g720 ( 
.A(n_579),
.Y(n_720)
);

BUFx6f_ASAP7_75t_SL g721 ( 
.A(n_678),
.Y(n_721)
);

AOI21xp5_ASAP7_75t_L g722 ( 
.A1(n_616),
.A2(n_270),
.B(n_280),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_L g723 ( 
.A(n_608),
.B(n_284),
.Y(n_723)
);

INVxp67_ASAP7_75t_L g724 ( 
.A(n_663),
.Y(n_724)
);

NOR2xp33_ASAP7_75t_L g725 ( 
.A(n_566),
.B(n_206),
.Y(n_725)
);

INVxp67_ASAP7_75t_L g726 ( 
.A(n_663),
.Y(n_726)
);

A2O1A1Ixp33_ASAP7_75t_L g727 ( 
.A1(n_577),
.A2(n_285),
.B(n_292),
.C(n_295),
.Y(n_727)
);

CKINVDCx5p33_ASAP7_75t_R g728 ( 
.A(n_601),
.Y(n_728)
);

BUFx3_ASAP7_75t_L g729 ( 
.A(n_587),
.Y(n_729)
);

AOI22xp33_ASAP7_75t_L g730 ( 
.A1(n_683),
.A2(n_367),
.B1(n_283),
.B2(n_273),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_590),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_581),
.B(n_307),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_L g733 ( 
.A(n_587),
.B(n_308),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_592),
.Y(n_734)
);

INVx8_ASAP7_75t_L g735 ( 
.A(n_569),
.Y(n_735)
);

AOI22xp33_ASAP7_75t_SL g736 ( 
.A1(n_599),
.A2(n_233),
.B1(n_208),
.B2(n_383),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_L g737 ( 
.A(n_587),
.B(n_311),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_SL g738 ( 
.A(n_569),
.B(n_599),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_SL g739 ( 
.A(n_569),
.B(n_351),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_SL g740 ( 
.A(n_683),
.B(n_351),
.Y(n_740)
);

NOR2xp33_ASAP7_75t_L g741 ( 
.A(n_580),
.B(n_206),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_593),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_SL g743 ( 
.A(n_563),
.B(n_351),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_SL g744 ( 
.A(n_568),
.B(n_213),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_L g745 ( 
.A(n_631),
.B(n_331),
.Y(n_745)
);

NOR2xp33_ASAP7_75t_L g746 ( 
.A(n_661),
.B(n_213),
.Y(n_746)
);

NOR2xp33_ASAP7_75t_L g747 ( 
.A(n_661),
.B(n_215),
.Y(n_747)
);

A2O1A1Ixp33_ASAP7_75t_L g748 ( 
.A1(n_577),
.A2(n_342),
.B(n_344),
.C(n_349),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_649),
.B(n_370),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_SL g750 ( 
.A(n_687),
.B(n_215),
.Y(n_750)
);

AND2x2_ASAP7_75t_SL g751 ( 
.A(n_687),
.B(n_378),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_594),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_L g753 ( 
.A(n_602),
.B(n_274),
.Y(n_753)
);

INVx2_ASAP7_75t_L g754 ( 
.A(n_578),
.Y(n_754)
);

INVxp67_ASAP7_75t_SL g755 ( 
.A(n_571),
.Y(n_755)
);

INVxp67_ASAP7_75t_L g756 ( 
.A(n_679),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_618),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_SL g758 ( 
.A(n_667),
.B(n_351),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_620),
.B(n_278),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_702),
.Y(n_760)
);

OR2x6_ASAP7_75t_L g761 ( 
.A(n_676),
.B(n_463),
.Y(n_761)
);

INVx2_ASAP7_75t_SL g762 ( 
.A(n_684),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_623),
.B(n_279),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_SL g764 ( 
.A(n_598),
.B(n_614),
.Y(n_764)
);

AND2x2_ASAP7_75t_L g765 ( 
.A(n_633),
.B(n_214),
.Y(n_765)
);

NOR2xp33_ASAP7_75t_L g766 ( 
.A(n_582),
.B(n_218),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_SL g767 ( 
.A(n_651),
.B(n_294),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_591),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_L g769 ( 
.A(n_636),
.B(n_296),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_L g770 ( 
.A(n_571),
.B(n_298),
.Y(n_770)
);

A2O1A1Ixp33_ASAP7_75t_L g771 ( 
.A1(n_681),
.A2(n_335),
.B(n_323),
.C(n_324),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_SL g772 ( 
.A(n_651),
.B(n_303),
.Y(n_772)
);

OAI21xp5_ASAP7_75t_L g773 ( 
.A1(n_626),
.A2(n_345),
.B(n_340),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_L g774 ( 
.A(n_571),
.B(n_313),
.Y(n_774)
);

NAND2x1p5_ASAP7_75t_L g775 ( 
.A(n_616),
.B(n_71),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_591),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_L g777 ( 
.A(n_670),
.B(n_314),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_591),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_SL g779 ( 
.A(n_671),
.B(n_316),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_670),
.B(n_655),
.Y(n_780)
);

BUFx6f_ASAP7_75t_L g781 ( 
.A(n_603),
.Y(n_781)
);

INVx3_ASAP7_75t_L g782 ( 
.A(n_664),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_L g783 ( 
.A(n_655),
.B(n_332),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_625),
.B(n_337),
.Y(n_784)
);

NOR2xp33_ASAP7_75t_L g785 ( 
.A(n_647),
.B(n_218),
.Y(n_785)
);

INVx2_ASAP7_75t_L g786 ( 
.A(n_595),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_SL g787 ( 
.A(n_671),
.B(n_346),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_SL g788 ( 
.A(n_609),
.B(n_221),
.Y(n_788)
);

NOR2xp33_ASAP7_75t_L g789 ( 
.A(n_657),
.B(n_222),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_603),
.Y(n_790)
);

NOR2xp33_ASAP7_75t_L g791 ( 
.A(n_657),
.B(n_222),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_628),
.B(n_224),
.Y(n_792)
);

NOR2xp33_ASAP7_75t_L g793 ( 
.A(n_668),
.B(n_672),
.Y(n_793)
);

AND2x2_ASAP7_75t_L g794 ( 
.A(n_615),
.B(n_214),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_L g795 ( 
.A(n_639),
.B(n_224),
.Y(n_795)
);

AND2x2_ASAP7_75t_L g796 ( 
.A(n_611),
.B(n_216),
.Y(n_796)
);

AOI22xp33_ASAP7_75t_L g797 ( 
.A1(n_673),
.A2(n_646),
.B1(n_698),
.B2(n_665),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_622),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_622),
.Y(n_799)
);

NOR2xp33_ASAP7_75t_SL g800 ( 
.A(n_601),
.B(n_227),
.Y(n_800)
);

INVx2_ASAP7_75t_SL g801 ( 
.A(n_685),
.Y(n_801)
);

INVx2_ASAP7_75t_L g802 ( 
.A(n_595),
.Y(n_802)
);

INVx2_ASAP7_75t_L g803 ( 
.A(n_596),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_SL g804 ( 
.A(n_642),
.B(n_227),
.Y(n_804)
);

INVx2_ASAP7_75t_L g805 ( 
.A(n_596),
.Y(n_805)
);

AOI22xp5_ASAP7_75t_L g806 ( 
.A1(n_570),
.A2(n_361),
.B1(n_229),
.B2(n_379),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_L g807 ( 
.A(n_621),
.B(n_701),
.Y(n_807)
);

INVx3_ASAP7_75t_L g808 ( 
.A(n_664),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_L g809 ( 
.A(n_701),
.B(n_229),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_701),
.B(n_234),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_L g811 ( 
.A(n_698),
.B(n_234),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_664),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_SL g813 ( 
.A(n_638),
.B(n_288),
.Y(n_813)
);

INVx4_ASAP7_75t_L g814 ( 
.A(n_617),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_L g815 ( 
.A(n_698),
.B(n_288),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_698),
.B(n_361),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_L g817 ( 
.A(n_597),
.B(n_363),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_L g818 ( 
.A(n_597),
.B(n_363),
.Y(n_818)
);

AND2x2_ASAP7_75t_L g819 ( 
.A(n_641),
.B(n_216),
.Y(n_819)
);

AOI21xp5_ASAP7_75t_L g820 ( 
.A1(n_632),
.A2(n_365),
.B(n_372),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_L g821 ( 
.A(n_606),
.B(n_607),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_L g822 ( 
.A(n_606),
.B(n_365),
.Y(n_822)
);

INVx8_ASAP7_75t_L g823 ( 
.A(n_700),
.Y(n_823)
);

OR2x6_ASAP7_75t_L g824 ( 
.A(n_676),
.B(n_27),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_613),
.Y(n_825)
);

AOI22xp5_ASAP7_75t_L g826 ( 
.A1(n_660),
.A2(n_372),
.B1(n_374),
.B2(n_379),
.Y(n_826)
);

AND2x2_ASAP7_75t_L g827 ( 
.A(n_645),
.B(n_357),
.Y(n_827)
);

O2A1O1Ixp33_ASAP7_75t_L g828 ( 
.A1(n_586),
.A2(n_668),
.B(n_672),
.C(n_644),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_SL g829 ( 
.A(n_632),
.B(n_658),
.Y(n_829)
);

AND2x2_ASAP7_75t_L g830 ( 
.A(n_648),
.B(n_681),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_613),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_L g832 ( 
.A(n_607),
.B(n_617),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_SL g833 ( 
.A(n_617),
.B(n_374),
.Y(n_833)
);

INVxp33_ASAP7_75t_L g834 ( 
.A(n_691),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_L g835 ( 
.A(n_629),
.B(n_447),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_L g836 ( 
.A(n_629),
.B(n_383),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_L g837 ( 
.A(n_629),
.B(n_377),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_613),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_567),
.Y(n_839)
);

NOR2xp33_ASAP7_75t_L g840 ( 
.A(n_677),
.B(n_377),
.Y(n_840)
);

BUFx3_ASAP7_75t_L g841 ( 
.A(n_604),
.Y(n_841)
);

HB1xp67_ASAP7_75t_L g842 ( 
.A(n_643),
.Y(n_842)
);

INVx2_ASAP7_75t_SL g843 ( 
.A(n_585),
.Y(n_843)
);

OAI21xp5_ASAP7_75t_L g844 ( 
.A1(n_635),
.A2(n_376),
.B(n_368),
.Y(n_844)
);

BUFx3_ASAP7_75t_L g845 ( 
.A(n_700),
.Y(n_845)
);

BUFx6f_ASAP7_75t_L g846 ( 
.A(n_640),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_567),
.Y(n_847)
);

BUFx8_ASAP7_75t_L g848 ( 
.A(n_680),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_575),
.Y(n_849)
);

NOR2xp67_ASAP7_75t_SL g850 ( 
.A(n_586),
.B(n_368),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_575),
.Y(n_851)
);

NOR2xp33_ASAP7_75t_L g852 ( 
.A(n_674),
.B(n_366),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_L g853 ( 
.A(n_640),
.B(n_366),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_640),
.B(n_362),
.Y(n_854)
);

AOI22xp5_ASAP7_75t_L g855 ( 
.A1(n_691),
.A2(n_362),
.B1(n_357),
.B2(n_356),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_SL g856 ( 
.A(n_640),
.B(n_356),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_SL g857 ( 
.A(n_699),
.B(n_355),
.Y(n_857)
);

BUFx3_ASAP7_75t_L g858 ( 
.A(n_699),
.Y(n_858)
);

AND2x2_ASAP7_75t_L g859 ( 
.A(n_762),
.B(n_692),
.Y(n_859)
);

O2A1O1Ixp33_ASAP7_75t_L g860 ( 
.A1(n_727),
.A2(n_674),
.B(n_673),
.C(n_589),
.Y(n_860)
);

NAND3x1_ASAP7_75t_L g861 ( 
.A(n_711),
.B(n_692),
.C(n_688),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_717),
.B(n_694),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_L g863 ( 
.A(n_717),
.B(n_694),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_SL g864 ( 
.A(n_706),
.B(n_680),
.Y(n_864)
);

BUFx4f_ASAP7_75t_L g865 ( 
.A(n_761),
.Y(n_865)
);

AOI21xp5_ASAP7_75t_L g866 ( 
.A1(n_807),
.A2(n_738),
.B(n_739),
.Y(n_866)
);

AND2x2_ASAP7_75t_L g867 ( 
.A(n_756),
.B(n_572),
.Y(n_867)
);

AOI22xp5_ASAP7_75t_L g868 ( 
.A1(n_738),
.A2(n_652),
.B1(n_605),
.B2(n_675),
.Y(n_868)
);

BUFx6f_ASAP7_75t_L g869 ( 
.A(n_735),
.Y(n_869)
);

HB1xp67_ASAP7_75t_L g870 ( 
.A(n_842),
.Y(n_870)
);

AOI21xp5_ASAP7_75t_L g871 ( 
.A1(n_739),
.A2(n_659),
.B(n_654),
.Y(n_871)
);

AOI221xp5_ASAP7_75t_L g872 ( 
.A1(n_704),
.A2(n_646),
.B1(n_665),
.B2(n_662),
.C(n_230),
.Y(n_872)
);

AOI21xp5_ASAP7_75t_L g873 ( 
.A1(n_780),
.A2(n_659),
.B(n_612),
.Y(n_873)
);

BUFx4f_ASAP7_75t_L g874 ( 
.A(n_761),
.Y(n_874)
);

AOI21xp5_ASAP7_75t_L g875 ( 
.A1(n_758),
.A2(n_612),
.B(n_589),
.Y(n_875)
);

OAI22xp5_ASAP7_75t_L g876 ( 
.A1(n_793),
.A2(n_682),
.B1(n_686),
.B2(n_662),
.Y(n_876)
);

OAI22xp5_ASAP7_75t_L g877 ( 
.A1(n_793),
.A2(n_682),
.B1(n_686),
.B2(n_693),
.Y(n_877)
);

A2O1A1Ixp33_ASAP7_75t_L g878 ( 
.A1(n_709),
.A2(n_695),
.B(n_689),
.C(n_588),
.Y(n_878)
);

AOI21xp5_ASAP7_75t_L g879 ( 
.A1(n_755),
.A2(n_814),
.B(n_769),
.Y(n_879)
);

AND2x6_ASAP7_75t_SL g880 ( 
.A(n_824),
.B(n_630),
.Y(n_880)
);

AOI21xp5_ASAP7_75t_L g881 ( 
.A1(n_814),
.A2(n_669),
.B(n_573),
.Y(n_881)
);

OAI22xp5_ASAP7_75t_L g882 ( 
.A1(n_797),
.A2(n_588),
.B1(n_600),
.B2(n_627),
.Y(n_882)
);

AOI21xp5_ASAP7_75t_L g883 ( 
.A1(n_777),
.A2(n_573),
.B(n_610),
.Y(n_883)
);

AND2x2_ASAP7_75t_L g884 ( 
.A(n_724),
.B(n_678),
.Y(n_884)
);

AOI21x1_ASAP7_75t_L g885 ( 
.A1(n_758),
.A2(n_600),
.B(n_627),
.Y(n_885)
);

AND2x2_ASAP7_75t_L g886 ( 
.A(n_726),
.B(n_678),
.Y(n_886)
);

NOR2xp33_ASAP7_75t_L g887 ( 
.A(n_834),
.B(n_696),
.Y(n_887)
);

AOI21xp5_ASAP7_75t_L g888 ( 
.A1(n_770),
.A2(n_573),
.B(n_610),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_L g889 ( 
.A(n_718),
.B(n_650),
.Y(n_889)
);

NOR2xp33_ASAP7_75t_L g890 ( 
.A(n_746),
.B(n_696),
.Y(n_890)
);

AOI21x1_ASAP7_75t_L g891 ( 
.A1(n_839),
.A2(n_619),
.B(n_634),
.Y(n_891)
);

INVx4_ASAP7_75t_L g892 ( 
.A(n_735),
.Y(n_892)
);

A2O1A1Ixp33_ASAP7_75t_L g893 ( 
.A1(n_746),
.A2(n_650),
.B(n_230),
.C(n_233),
.Y(n_893)
);

INVx1_ASAP7_75t_SL g894 ( 
.A(n_843),
.Y(n_894)
);

AND2x2_ASAP7_75t_L g895 ( 
.A(n_830),
.B(n_696),
.Y(n_895)
);

INVx2_ASAP7_75t_L g896 ( 
.A(n_808),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_L g897 ( 
.A(n_723),
.B(n_747),
.Y(n_897)
);

OAI21xp33_ASAP7_75t_L g898 ( 
.A1(n_747),
.A2(n_228),
.B(n_353),
.Y(n_898)
);

AND2x2_ASAP7_75t_L g899 ( 
.A(n_765),
.B(n_696),
.Y(n_899)
);

AND2x6_ASAP7_75t_L g900 ( 
.A(n_768),
.B(n_666),
.Y(n_900)
);

AOI21xp5_ASAP7_75t_L g901 ( 
.A1(n_743),
.A2(n_666),
.B(n_656),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_L g902 ( 
.A(n_840),
.B(n_666),
.Y(n_902)
);

OAI321xp33_ASAP7_75t_L g903 ( 
.A1(n_852),
.A2(n_652),
.A3(n_353),
.B1(n_354),
.B2(n_355),
.C(n_228),
.Y(n_903)
);

AND3x2_ASAP7_75t_L g904 ( 
.A(n_852),
.B(n_690),
.C(n_354),
.Y(n_904)
);

AOI21x1_ASAP7_75t_L g905 ( 
.A1(n_847),
.A2(n_666),
.B(n_656),
.Y(n_905)
);

AOI21xp5_ASAP7_75t_L g906 ( 
.A1(n_774),
.A2(n_712),
.B(n_783),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_L g907 ( 
.A(n_840),
.B(n_656),
.Y(n_907)
);

O2A1O1Ixp33_ASAP7_75t_SL g908 ( 
.A1(n_748),
.A2(n_653),
.B(n_31),
.C(n_32),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_849),
.Y(n_909)
);

NOR3xp33_ASAP7_75t_L g910 ( 
.A(n_857),
.B(n_690),
.C(n_33),
.Y(n_910)
);

BUFx4f_ASAP7_75t_L g911 ( 
.A(n_761),
.Y(n_911)
);

INVxp33_ASAP7_75t_L g912 ( 
.A(n_796),
.Y(n_912)
);

BUFx6f_ASAP7_75t_L g913 ( 
.A(n_735),
.Y(n_913)
);

AOI22xp33_ASAP7_75t_L g914 ( 
.A1(n_751),
.A2(n_653),
.B1(n_690),
.B2(n_624),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_L g915 ( 
.A(n_725),
.B(n_624),
.Y(n_915)
);

AOI21xp5_ASAP7_75t_L g916 ( 
.A1(n_733),
.A2(n_653),
.B(n_100),
.Y(n_916)
);

OAI22xp5_ASAP7_75t_L g917 ( 
.A1(n_751),
.A2(n_690),
.B1(n_98),
.B2(n_102),
.Y(n_917)
);

A2O1A1Ixp33_ASAP7_75t_L g918 ( 
.A1(n_828),
.A2(n_28),
.B(n_35),
.C(n_40),
.Y(n_918)
);

AOI21xp5_ASAP7_75t_L g919 ( 
.A1(n_737),
.A2(n_653),
.B(n_104),
.Y(n_919)
);

NOR2x1_ASAP7_75t_L g920 ( 
.A(n_858),
.B(n_96),
.Y(n_920)
);

NOR2xp33_ASAP7_75t_L g921 ( 
.A(n_715),
.B(n_35),
.Y(n_921)
);

O2A1O1Ixp5_ASAP7_75t_L g922 ( 
.A1(n_764),
.A2(n_653),
.B(n_109),
.C(n_113),
.Y(n_922)
);

OAI22xp33_ASAP7_75t_L g923 ( 
.A1(n_842),
.A2(n_41),
.B1(n_42),
.B2(n_44),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_L g924 ( 
.A(n_725),
.B(n_710),
.Y(n_924)
);

AOI21xp5_ASAP7_75t_L g925 ( 
.A1(n_784),
.A2(n_117),
.B(n_185),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_SL g926 ( 
.A(n_781),
.B(n_93),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_851),
.Y(n_927)
);

CKINVDCx20_ASAP7_75t_R g928 ( 
.A(n_728),
.Y(n_928)
);

HB1xp67_ASAP7_75t_L g929 ( 
.A(n_801),
.Y(n_929)
);

INVxp67_ASAP7_75t_L g930 ( 
.A(n_827),
.Y(n_930)
);

NOR2xp33_ASAP7_75t_L g931 ( 
.A(n_800),
.B(n_41),
.Y(n_931)
);

OAI21xp5_ASAP7_75t_L g932 ( 
.A1(n_745),
.A2(n_118),
.B(n_170),
.Y(n_932)
);

AOI21xp5_ASAP7_75t_L g933 ( 
.A1(n_749),
.A2(n_90),
.B(n_165),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_L g934 ( 
.A(n_710),
.B(n_785),
.Y(n_934)
);

INVx2_ASAP7_75t_L g935 ( 
.A(n_754),
.Y(n_935)
);

NOR2xp33_ASAP7_75t_L g936 ( 
.A(n_857),
.B(n_45),
.Y(n_936)
);

AOI21xp5_ASAP7_75t_L g937 ( 
.A1(n_767),
.A2(n_119),
.B(n_156),
.Y(n_937)
);

AOI21xp5_ASAP7_75t_L g938 ( 
.A1(n_767),
.A2(n_74),
.B(n_150),
.Y(n_938)
);

NOR2xp33_ASAP7_75t_R g939 ( 
.A(n_823),
.B(n_189),
.Y(n_939)
);

OAI22xp5_ASAP7_75t_L g940 ( 
.A1(n_829),
.A2(n_139),
.B1(n_137),
.B2(n_126),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_L g941 ( 
.A(n_789),
.B(n_52),
.Y(n_941)
);

NOR2x1_ASAP7_75t_L g942 ( 
.A(n_858),
.B(n_120),
.Y(n_942)
);

AOI21xp5_ASAP7_75t_L g943 ( 
.A1(n_772),
.A2(n_787),
.B(n_779),
.Y(n_943)
);

AOI21xp5_ASAP7_75t_L g944 ( 
.A1(n_772),
.A2(n_121),
.B(n_55),
.Y(n_944)
);

AOI21xp5_ASAP7_75t_L g945 ( 
.A1(n_779),
.A2(n_54),
.B(n_56),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_L g946 ( 
.A(n_789),
.B(n_57),
.Y(n_946)
);

OAI21x1_ASAP7_75t_L g947 ( 
.A1(n_786),
.A2(n_59),
.B(n_802),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_L g948 ( 
.A(n_791),
.B(n_713),
.Y(n_948)
);

BUFx6f_ASAP7_75t_L g949 ( 
.A(n_707),
.Y(n_949)
);

OAI22x1_ASAP7_75t_L g950 ( 
.A1(n_855),
.A2(n_788),
.B1(n_764),
.B2(n_806),
.Y(n_950)
);

CKINVDCx10_ASAP7_75t_R g951 ( 
.A(n_721),
.Y(n_951)
);

AOI22xp33_ASAP7_75t_L g952 ( 
.A1(n_740),
.A2(n_750),
.B1(n_791),
.B2(n_788),
.Y(n_952)
);

NOR2xp33_ASAP7_75t_L g953 ( 
.A(n_766),
.B(n_794),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_L g954 ( 
.A(n_716),
.B(n_719),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_L g955 ( 
.A(n_731),
.B(n_734),
.Y(n_955)
);

AOI21x1_ASAP7_75t_L g956 ( 
.A1(n_787),
.A2(n_810),
.B(n_809),
.Y(n_956)
);

NOR2x1p5_ASAP7_75t_SL g957 ( 
.A(n_803),
.B(n_805),
.Y(n_957)
);

INVx1_ASAP7_75t_L g958 ( 
.A(n_742),
.Y(n_958)
);

HB1xp67_ASAP7_75t_L g959 ( 
.A(n_836),
.Y(n_959)
);

INVx5_ASAP7_75t_L g960 ( 
.A(n_846),
.Y(n_960)
);

HB1xp67_ASAP7_75t_L g961 ( 
.A(n_837),
.Y(n_961)
);

AOI21xp5_ASAP7_75t_L g962 ( 
.A1(n_846),
.A2(n_835),
.B(n_822),
.Y(n_962)
);

AOI21xp5_ASAP7_75t_L g963 ( 
.A1(n_846),
.A2(n_818),
.B(n_817),
.Y(n_963)
);

INVx1_ASAP7_75t_L g964 ( 
.A(n_752),
.Y(n_964)
);

BUFx2_ASAP7_75t_L g965 ( 
.A(n_848),
.Y(n_965)
);

AND2x2_ASAP7_75t_L g966 ( 
.A(n_819),
.B(n_730),
.Y(n_966)
);

A2O1A1Ixp33_ASAP7_75t_L g967 ( 
.A1(n_844),
.A2(n_741),
.B(n_838),
.C(n_831),
.Y(n_967)
);

AOI21xp5_ASAP7_75t_L g968 ( 
.A1(n_714),
.A2(n_720),
.B(n_732),
.Y(n_968)
);

NAND3xp33_ASAP7_75t_L g969 ( 
.A(n_730),
.B(n_736),
.C(n_766),
.Y(n_969)
);

AOI22xp5_ASAP7_75t_L g970 ( 
.A1(n_776),
.A2(n_778),
.B1(n_825),
.B2(n_741),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_L g971 ( 
.A(n_757),
.B(n_760),
.Y(n_971)
);

BUFx4f_ASAP7_75t_L g972 ( 
.A(n_823),
.Y(n_972)
);

AOI21xp5_ASAP7_75t_L g973 ( 
.A1(n_792),
.A2(n_795),
.B(n_854),
.Y(n_973)
);

NOR2xp33_ASAP7_75t_L g974 ( 
.A(n_813),
.B(n_744),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_L g975 ( 
.A(n_790),
.B(n_798),
.Y(n_975)
);

A2O1A1Ixp33_ASAP7_75t_L g976 ( 
.A1(n_771),
.A2(n_799),
.B(n_856),
.C(n_729),
.Y(n_976)
);

NOR2xp33_ASAP7_75t_L g977 ( 
.A(n_826),
.B(n_763),
.Y(n_977)
);

INVx2_ASAP7_75t_L g978 ( 
.A(n_781),
.Y(n_978)
);

NAND2xp5_ASAP7_75t_L g979 ( 
.A(n_853),
.B(n_773),
.Y(n_979)
);

INVxp67_ASAP7_75t_SL g980 ( 
.A(n_775),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_L g981 ( 
.A(n_804),
.B(n_753),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_L g982 ( 
.A(n_804),
.B(n_759),
.Y(n_982)
);

AOI21xp5_ASAP7_75t_L g983 ( 
.A1(n_833),
.A2(n_708),
.B(n_856),
.Y(n_983)
);

INVx3_ASAP7_75t_L g984 ( 
.A(n_775),
.Y(n_984)
);

AND2x4_ASAP7_75t_L g985 ( 
.A(n_841),
.B(n_833),
.Y(n_985)
);

OAI21xp5_ASAP7_75t_L g986 ( 
.A1(n_811),
.A2(n_815),
.B(n_816),
.Y(n_986)
);

NAND2xp5_ASAP7_75t_L g987 ( 
.A(n_850),
.B(n_820),
.Y(n_987)
);

INVx2_ASAP7_75t_L g988 ( 
.A(n_824),
.Y(n_988)
);

INVx1_ASAP7_75t_L g989 ( 
.A(n_824),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_L g990 ( 
.A(n_722),
.B(n_848),
.Y(n_990)
);

OAI21xp5_ASAP7_75t_L g991 ( 
.A1(n_841),
.A2(n_845),
.B(n_721),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_L g992 ( 
.A(n_845),
.B(n_823),
.Y(n_992)
);

AOI21xp5_ASAP7_75t_L g993 ( 
.A1(n_807),
.A2(n_738),
.B(n_739),
.Y(n_993)
);

BUFx3_ASAP7_75t_L g994 ( 
.A(n_841),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_SL g995 ( 
.A(n_706),
.B(n_781),
.Y(n_995)
);

O2A1O1Ixp33_ASAP7_75t_L g996 ( 
.A1(n_727),
.A2(n_748),
.B(n_740),
.C(n_705),
.Y(n_996)
);

AOI21xp5_ASAP7_75t_L g997 ( 
.A1(n_807),
.A2(n_632),
.B(n_616),
.Y(n_997)
);

AO22x1_ASAP7_75t_L g998 ( 
.A1(n_717),
.A2(n_834),
.B1(n_747),
.B2(n_746),
.Y(n_998)
);

AOI21xp5_ASAP7_75t_L g999 ( 
.A1(n_807),
.A2(n_632),
.B(n_616),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_SL g1000 ( 
.A(n_706),
.B(n_781),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_L g1001 ( 
.A(n_717),
.B(n_565),
.Y(n_1001)
);

BUFx12f_ASAP7_75t_L g1002 ( 
.A(n_848),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_L g1003 ( 
.A(n_717),
.B(n_565),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_812),
.Y(n_1004)
);

INVx3_ASAP7_75t_L g1005 ( 
.A(n_729),
.Y(n_1005)
);

INVx2_ASAP7_75t_L g1006 ( 
.A(n_782),
.Y(n_1006)
);

NOR2xp33_ASAP7_75t_L g1007 ( 
.A(n_724),
.B(n_726),
.Y(n_1007)
);

AOI22xp5_ASAP7_75t_L g1008 ( 
.A1(n_738),
.A2(n_717),
.B1(n_793),
.B2(n_706),
.Y(n_1008)
);

AOI21xp5_ASAP7_75t_L g1009 ( 
.A1(n_807),
.A2(n_738),
.B(n_739),
.Y(n_1009)
);

INVx1_ASAP7_75t_L g1010 ( 
.A(n_812),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_SL g1011 ( 
.A(n_706),
.B(n_781),
.Y(n_1011)
);

INVx11_ASAP7_75t_L g1012 ( 
.A(n_848),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_L g1013 ( 
.A(n_717),
.B(n_565),
.Y(n_1013)
);

INVx1_ASAP7_75t_L g1014 ( 
.A(n_812),
.Y(n_1014)
);

AOI21xp5_ASAP7_75t_L g1015 ( 
.A1(n_807),
.A2(n_738),
.B(n_739),
.Y(n_1015)
);

OAI21x1_ASAP7_75t_L g1016 ( 
.A1(n_832),
.A2(n_821),
.B(n_780),
.Y(n_1016)
);

INVx3_ASAP7_75t_L g1017 ( 
.A(n_729),
.Y(n_1017)
);

INVx1_ASAP7_75t_L g1018 ( 
.A(n_812),
.Y(n_1018)
);

OAI22xp5_ASAP7_75t_L g1019 ( 
.A1(n_706),
.A2(n_793),
.B1(n_717),
.B2(n_705),
.Y(n_1019)
);

A2O1A1Ixp33_ASAP7_75t_L g1020 ( 
.A1(n_717),
.A2(n_793),
.B(n_565),
.C(n_709),
.Y(n_1020)
);

NAND2xp5_ASAP7_75t_L g1021 ( 
.A(n_717),
.B(n_565),
.Y(n_1021)
);

O2A1O1Ixp33_ASAP7_75t_L g1022 ( 
.A1(n_727),
.A2(n_748),
.B(n_740),
.C(n_705),
.Y(n_1022)
);

AOI21xp5_ASAP7_75t_L g1023 ( 
.A1(n_807),
.A2(n_738),
.B(n_739),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_L g1024 ( 
.A(n_717),
.B(n_565),
.Y(n_1024)
);

NAND2xp5_ASAP7_75t_L g1025 ( 
.A(n_717),
.B(n_565),
.Y(n_1025)
);

AOI21xp5_ASAP7_75t_L g1026 ( 
.A1(n_807),
.A2(n_738),
.B(n_739),
.Y(n_1026)
);

NAND2xp5_ASAP7_75t_L g1027 ( 
.A(n_717),
.B(n_565),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_L g1028 ( 
.A(n_1001),
.B(n_1003),
.Y(n_1028)
);

BUFx3_ASAP7_75t_L g1029 ( 
.A(n_928),
.Y(n_1029)
);

OAI21x1_ASAP7_75t_L g1030 ( 
.A1(n_1016),
.A2(n_901),
.B(n_962),
.Y(n_1030)
);

NAND2x1p5_ASAP7_75t_L g1031 ( 
.A(n_892),
.B(n_869),
.Y(n_1031)
);

OAI21x1_ASAP7_75t_L g1032 ( 
.A1(n_901),
.A2(n_963),
.B(n_885),
.Y(n_1032)
);

NAND2x1_ASAP7_75t_L g1033 ( 
.A(n_900),
.B(n_892),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_SL g1034 ( 
.A(n_953),
.B(n_862),
.Y(n_1034)
);

BUFx3_ASAP7_75t_L g1035 ( 
.A(n_994),
.Y(n_1035)
);

AO31x2_ASAP7_75t_L g1036 ( 
.A1(n_1020),
.A2(n_1019),
.A3(n_918),
.B(n_878),
.Y(n_1036)
);

NAND2xp5_ASAP7_75t_L g1037 ( 
.A(n_1013),
.B(n_1021),
.Y(n_1037)
);

OAI21x1_ASAP7_75t_SL g1038 ( 
.A1(n_932),
.A2(n_1022),
.B(n_996),
.Y(n_1038)
);

INVx6_ASAP7_75t_L g1039 ( 
.A(n_1002),
.Y(n_1039)
);

OAI22xp33_ASAP7_75t_L g1040 ( 
.A1(n_1024),
.A2(n_1027),
.B1(n_1025),
.B2(n_863),
.Y(n_1040)
);

BUFx3_ASAP7_75t_L g1041 ( 
.A(n_972),
.Y(n_1041)
);

BUFx3_ASAP7_75t_L g1042 ( 
.A(n_972),
.Y(n_1042)
);

BUFx3_ASAP7_75t_L g1043 ( 
.A(n_894),
.Y(n_1043)
);

NOR2xp33_ASAP7_75t_L g1044 ( 
.A(n_1007),
.B(n_924),
.Y(n_1044)
);

OAI21xp33_ASAP7_75t_L g1045 ( 
.A1(n_898),
.A2(n_969),
.B(n_897),
.Y(n_1045)
);

OR2x2_ASAP7_75t_L g1046 ( 
.A(n_966),
.B(n_870),
.Y(n_1046)
);

AOI221xp5_ASAP7_75t_L g1047 ( 
.A1(n_903),
.A2(n_936),
.B1(n_921),
.B2(n_998),
.C(n_923),
.Y(n_1047)
);

OR2x2_ASAP7_75t_L g1048 ( 
.A(n_948),
.B(n_867),
.Y(n_1048)
);

OR2x6_ASAP7_75t_L g1049 ( 
.A(n_869),
.B(n_913),
.Y(n_1049)
);

AND2x2_ASAP7_75t_L g1050 ( 
.A(n_912),
.B(n_884),
.Y(n_1050)
);

A2O1A1Ixp33_ASAP7_75t_SL g1051 ( 
.A1(n_890),
.A2(n_974),
.B(n_977),
.C(n_887),
.Y(n_1051)
);

OAI21xp5_ASAP7_75t_L g1052 ( 
.A1(n_1008),
.A2(n_993),
.B(n_866),
.Y(n_1052)
);

NOR2x1_ASAP7_75t_SL g1053 ( 
.A(n_960),
.B(n_869),
.Y(n_1053)
);

NOR2xp33_ASAP7_75t_L g1054 ( 
.A(n_934),
.B(n_959),
.Y(n_1054)
);

AOI221x1_ASAP7_75t_L g1055 ( 
.A1(n_950),
.A2(n_946),
.B1(n_941),
.B2(n_943),
.C(n_979),
.Y(n_1055)
);

OAI21xp5_ASAP7_75t_L g1056 ( 
.A1(n_1026),
.A2(n_1015),
.B(n_1009),
.Y(n_1056)
);

AND2x4_ASAP7_75t_L g1057 ( 
.A(n_913),
.B(n_949),
.Y(n_1057)
);

O2A1O1Ixp5_ASAP7_75t_L g1058 ( 
.A1(n_915),
.A2(n_864),
.B(n_987),
.C(n_997),
.Y(n_1058)
);

AOI21xp5_ASAP7_75t_L g1059 ( 
.A1(n_1009),
.A2(n_1026),
.B(n_1015),
.Y(n_1059)
);

NAND2xp5_ASAP7_75t_L g1060 ( 
.A(n_961),
.B(n_876),
.Y(n_1060)
);

INVx4_ASAP7_75t_L g1061 ( 
.A(n_913),
.Y(n_1061)
);

AND2x2_ASAP7_75t_L g1062 ( 
.A(n_886),
.B(n_859),
.Y(n_1062)
);

AOI21xp5_ASAP7_75t_L g1063 ( 
.A1(n_1023),
.A2(n_960),
.B(n_906),
.Y(n_1063)
);

INVx1_ASAP7_75t_L g1064 ( 
.A(n_958),
.Y(n_1064)
);

NAND2xp5_ASAP7_75t_L g1065 ( 
.A(n_981),
.B(n_982),
.Y(n_1065)
);

AOI21xp5_ASAP7_75t_L g1066 ( 
.A1(n_960),
.A2(n_999),
.B(n_973),
.Y(n_1066)
);

INVx1_ASAP7_75t_L g1067 ( 
.A(n_964),
.Y(n_1067)
);

AOI21xp5_ASAP7_75t_L g1068 ( 
.A1(n_973),
.A2(n_879),
.B(n_902),
.Y(n_1068)
);

OAI21x1_ASAP7_75t_L g1069 ( 
.A1(n_871),
.A2(n_883),
.B(n_888),
.Y(n_1069)
);

INVx3_ASAP7_75t_SL g1070 ( 
.A(n_985),
.Y(n_1070)
);

BUFx4_ASAP7_75t_SL g1071 ( 
.A(n_880),
.Y(n_1071)
);

A2O1A1Ixp33_ASAP7_75t_L g1072 ( 
.A1(n_860),
.A2(n_952),
.B(n_967),
.C(n_983),
.Y(n_1072)
);

AND3x4_ASAP7_75t_L g1073 ( 
.A(n_910),
.B(n_985),
.C(n_988),
.Y(n_1073)
);

CKINVDCx5p33_ASAP7_75t_R g1074 ( 
.A(n_951),
.Y(n_1074)
);

AND2x6_ASAP7_75t_L g1075 ( 
.A(n_984),
.B(n_920),
.Y(n_1075)
);

INVx1_ASAP7_75t_L g1076 ( 
.A(n_1004),
.Y(n_1076)
);

OAI21xp5_ASAP7_75t_L g1077 ( 
.A1(n_882),
.A2(n_986),
.B(n_983),
.Y(n_1077)
);

AOI21x1_ASAP7_75t_L g1078 ( 
.A1(n_956),
.A2(n_907),
.B(n_873),
.Y(n_1078)
);

AO31x2_ASAP7_75t_L g1079 ( 
.A1(n_943),
.A2(n_976),
.A3(n_893),
.B(n_873),
.Y(n_1079)
);

NAND2xp5_ASAP7_75t_SL g1080 ( 
.A(n_868),
.B(n_949),
.Y(n_1080)
);

CKINVDCx5p33_ASAP7_75t_R g1081 ( 
.A(n_1012),
.Y(n_1081)
);

NAND2xp5_ASAP7_75t_L g1082 ( 
.A(n_995),
.B(n_1000),
.Y(n_1082)
);

NAND2xp5_ASAP7_75t_L g1083 ( 
.A(n_1011),
.B(n_889),
.Y(n_1083)
);

NAND2xp5_ASAP7_75t_L g1084 ( 
.A(n_954),
.B(n_955),
.Y(n_1084)
);

BUFx3_ASAP7_75t_L g1085 ( 
.A(n_992),
.Y(n_1085)
);

OAI21x1_ASAP7_75t_L g1086 ( 
.A1(n_968),
.A2(n_875),
.B(n_947),
.Y(n_1086)
);

AOI21xp33_ASAP7_75t_L g1087 ( 
.A1(n_931),
.A2(n_877),
.B(n_971),
.Y(n_1087)
);

AO21x1_ASAP7_75t_L g1088 ( 
.A1(n_940),
.A2(n_944),
.B(n_945),
.Y(n_1088)
);

NAND2xp5_ASAP7_75t_L g1089 ( 
.A(n_1010),
.B(n_1018),
.Y(n_1089)
);

AOI21x1_ASAP7_75t_L g1090 ( 
.A1(n_881),
.A2(n_927),
.B(n_909),
.Y(n_1090)
);

INVx1_ASAP7_75t_SL g1091 ( 
.A(n_895),
.Y(n_1091)
);

INVx5_ASAP7_75t_L g1092 ( 
.A(n_900),
.Y(n_1092)
);

OAI21xp5_ASAP7_75t_L g1093 ( 
.A1(n_922),
.A2(n_970),
.B(n_1014),
.Y(n_1093)
);

AO21x1_ASAP7_75t_L g1094 ( 
.A1(n_980),
.A2(n_933),
.B(n_938),
.Y(n_1094)
);

OAI21xp33_ASAP7_75t_L g1095 ( 
.A1(n_930),
.A2(n_975),
.B(n_899),
.Y(n_1095)
);

NOR2x1_ASAP7_75t_R g1096 ( 
.A(n_965),
.B(n_990),
.Y(n_1096)
);

NAND2xp5_ASAP7_75t_L g1097 ( 
.A(n_1005),
.B(n_1017),
.Y(n_1097)
);

A2O1A1Ixp33_ASAP7_75t_L g1098 ( 
.A1(n_984),
.A2(n_872),
.B(n_896),
.C(n_1006),
.Y(n_1098)
);

BUFx3_ASAP7_75t_L g1099 ( 
.A(n_929),
.Y(n_1099)
);

AOI21xp5_ASAP7_75t_L g1100 ( 
.A1(n_1005),
.A2(n_1017),
.B(n_978),
.Y(n_1100)
);

A2O1A1Ixp33_ASAP7_75t_L g1101 ( 
.A1(n_872),
.A2(n_937),
.B(n_957),
.C(n_935),
.Y(n_1101)
);

AND2x4_ASAP7_75t_L g1102 ( 
.A(n_949),
.B(n_989),
.Y(n_1102)
);

NAND2xp5_ASAP7_75t_L g1103 ( 
.A(n_900),
.B(n_942),
.Y(n_1103)
);

NAND2xp5_ASAP7_75t_L g1104 ( 
.A(n_900),
.B(n_914),
.Y(n_1104)
);

INVx1_ASAP7_75t_SL g1105 ( 
.A(n_861),
.Y(n_1105)
);

NAND2xp5_ASAP7_75t_SL g1106 ( 
.A(n_865),
.B(n_874),
.Y(n_1106)
);

BUFx3_ASAP7_75t_L g1107 ( 
.A(n_865),
.Y(n_1107)
);

AOI21xp33_ASAP7_75t_L g1108 ( 
.A1(n_917),
.A2(n_926),
.B(n_874),
.Y(n_1108)
);

AND3x4_ASAP7_75t_L g1109 ( 
.A(n_904),
.B(n_991),
.C(n_911),
.Y(n_1109)
);

INVx1_ASAP7_75t_L g1110 ( 
.A(n_900),
.Y(n_1110)
);

NOR2xp67_ASAP7_75t_L g1111 ( 
.A(n_925),
.B(n_916),
.Y(n_1111)
);

NAND2xp5_ASAP7_75t_SL g1112 ( 
.A(n_911),
.B(n_939),
.Y(n_1112)
);

AOI21xp33_ASAP7_75t_L g1113 ( 
.A1(n_919),
.A2(n_1003),
.B(n_1001),
.Y(n_1113)
);

NAND2xp5_ASAP7_75t_L g1114 ( 
.A(n_908),
.B(n_1001),
.Y(n_1114)
);

AOI21xp33_ASAP7_75t_L g1115 ( 
.A1(n_1001),
.A2(n_1013),
.B(n_1003),
.Y(n_1115)
);

AOI221xp5_ASAP7_75t_SL g1116 ( 
.A1(n_1020),
.A2(n_1013),
.B1(n_1021),
.B2(n_1003),
.C(n_1001),
.Y(n_1116)
);

AO21x1_ASAP7_75t_L g1117 ( 
.A1(n_1019),
.A2(n_924),
.B(n_934),
.Y(n_1117)
);

NAND2xp5_ASAP7_75t_SL g1118 ( 
.A(n_953),
.B(n_706),
.Y(n_1118)
);

BUFx3_ASAP7_75t_L g1119 ( 
.A(n_928),
.Y(n_1119)
);

NAND2xp5_ASAP7_75t_L g1120 ( 
.A(n_1001),
.B(n_1003),
.Y(n_1120)
);

OAI21xp5_ASAP7_75t_L g1121 ( 
.A1(n_1020),
.A2(n_1008),
.B(n_1019),
.Y(n_1121)
);

A2O1A1Ixp33_ASAP7_75t_L g1122 ( 
.A1(n_1020),
.A2(n_1001),
.B(n_1013),
.C(n_1003),
.Y(n_1122)
);

NAND2xp5_ASAP7_75t_L g1123 ( 
.A(n_1001),
.B(n_1003),
.Y(n_1123)
);

OAI21xp33_ASAP7_75t_L g1124 ( 
.A1(n_1001),
.A2(n_730),
.B(n_717),
.Y(n_1124)
);

INVx1_ASAP7_75t_L g1125 ( 
.A(n_958),
.Y(n_1125)
);

NOR2xp33_ASAP7_75t_L g1126 ( 
.A(n_1001),
.B(n_724),
.Y(n_1126)
);

CKINVDCx5p33_ASAP7_75t_R g1127 ( 
.A(n_928),
.Y(n_1127)
);

AOI21xp33_ASAP7_75t_L g1128 ( 
.A1(n_1001),
.A2(n_1013),
.B(n_1003),
.Y(n_1128)
);

A2O1A1Ixp33_ASAP7_75t_L g1129 ( 
.A1(n_1020),
.A2(n_1001),
.B(n_1013),
.C(n_1003),
.Y(n_1129)
);

AND2x2_ASAP7_75t_L g1130 ( 
.A(n_966),
.B(n_756),
.Y(n_1130)
);

INVx2_ASAP7_75t_SL g1131 ( 
.A(n_894),
.Y(n_1131)
);

OR2x6_ASAP7_75t_L g1132 ( 
.A(n_869),
.B(n_823),
.Y(n_1132)
);

INVx1_ASAP7_75t_L g1133 ( 
.A(n_958),
.Y(n_1133)
);

BUFx6f_ASAP7_75t_L g1134 ( 
.A(n_869),
.Y(n_1134)
);

AOI22x1_ASAP7_75t_L g1135 ( 
.A1(n_950),
.A2(n_943),
.B1(n_973),
.B2(n_983),
.Y(n_1135)
);

A2O1A1Ixp33_ASAP7_75t_L g1136 ( 
.A1(n_1020),
.A2(n_1001),
.B(n_1013),
.C(n_1003),
.Y(n_1136)
);

AOI221x1_ASAP7_75t_L g1137 ( 
.A1(n_1020),
.A2(n_1019),
.B1(n_924),
.B2(n_1025),
.C(n_1024),
.Y(n_1137)
);

AOI22xp5_ASAP7_75t_L g1138 ( 
.A1(n_1001),
.A2(n_1013),
.B1(n_1021),
.B2(n_1003),
.Y(n_1138)
);

OAI21xp5_ASAP7_75t_L g1139 ( 
.A1(n_1020),
.A2(n_1008),
.B(n_1019),
.Y(n_1139)
);

AND2x4_ASAP7_75t_L g1140 ( 
.A(n_892),
.B(n_869),
.Y(n_1140)
);

CKINVDCx8_ASAP7_75t_R g1141 ( 
.A(n_951),
.Y(n_1141)
);

NOR2x1_ASAP7_75t_SL g1142 ( 
.A(n_960),
.B(n_869),
.Y(n_1142)
);

OR2x6_ASAP7_75t_L g1143 ( 
.A(n_869),
.B(n_823),
.Y(n_1143)
);

INVx1_ASAP7_75t_L g1144 ( 
.A(n_958),
.Y(n_1144)
);

OAI21x1_ASAP7_75t_SL g1145 ( 
.A1(n_932),
.A2(n_1022),
.B(n_996),
.Y(n_1145)
);

NAND2xp5_ASAP7_75t_SL g1146 ( 
.A(n_953),
.B(n_706),
.Y(n_1146)
);

AND2x2_ASAP7_75t_L g1147 ( 
.A(n_966),
.B(n_756),
.Y(n_1147)
);

A2O1A1Ixp33_ASAP7_75t_L g1148 ( 
.A1(n_1020),
.A2(n_1001),
.B(n_1013),
.C(n_1003),
.Y(n_1148)
);

AND2x2_ASAP7_75t_L g1149 ( 
.A(n_966),
.B(n_756),
.Y(n_1149)
);

OAI21x1_ASAP7_75t_L g1150 ( 
.A1(n_1016),
.A2(n_905),
.B(n_891),
.Y(n_1150)
);

NOR2xp33_ASAP7_75t_L g1151 ( 
.A(n_1001),
.B(n_724),
.Y(n_1151)
);

AO31x2_ASAP7_75t_L g1152 ( 
.A1(n_1020),
.A2(n_1019),
.A3(n_918),
.B(n_878),
.Y(n_1152)
);

INVx1_ASAP7_75t_SL g1153 ( 
.A(n_894),
.Y(n_1153)
);

AOI221xp5_ASAP7_75t_L g1154 ( 
.A1(n_969),
.A2(n_673),
.B1(n_683),
.B2(n_1003),
.C(n_1001),
.Y(n_1154)
);

NAND2xp5_ASAP7_75t_SL g1155 ( 
.A(n_953),
.B(n_706),
.Y(n_1155)
);

OAI21x1_ASAP7_75t_L g1156 ( 
.A1(n_1016),
.A2(n_905),
.B(n_891),
.Y(n_1156)
);

NAND2xp5_ASAP7_75t_L g1157 ( 
.A(n_1001),
.B(n_1003),
.Y(n_1157)
);

INVx3_ASAP7_75t_L g1158 ( 
.A(n_1033),
.Y(n_1158)
);

CKINVDCx16_ASAP7_75t_R g1159 ( 
.A(n_1029),
.Y(n_1159)
);

AND2x4_ASAP7_75t_L g1160 ( 
.A(n_1057),
.B(n_1102),
.Y(n_1160)
);

INVx2_ASAP7_75t_SL g1161 ( 
.A(n_1043),
.Y(n_1161)
);

INVx2_ASAP7_75t_SL g1162 ( 
.A(n_1035),
.Y(n_1162)
);

AND2x2_ASAP7_75t_L g1163 ( 
.A(n_1149),
.B(n_1054),
.Y(n_1163)
);

NAND2xp5_ASAP7_75t_L g1164 ( 
.A(n_1044),
.B(n_1138),
.Y(n_1164)
);

AOI21xp5_ASAP7_75t_L g1165 ( 
.A1(n_1063),
.A2(n_1077),
.B(n_1068),
.Y(n_1165)
);

NAND2xp5_ASAP7_75t_L g1166 ( 
.A(n_1028),
.B(n_1037),
.Y(n_1166)
);

INVx3_ASAP7_75t_L g1167 ( 
.A(n_1092),
.Y(n_1167)
);

AND2x2_ASAP7_75t_L g1168 ( 
.A(n_1126),
.B(n_1151),
.Y(n_1168)
);

AND2x2_ASAP7_75t_L g1169 ( 
.A(n_1062),
.B(n_1050),
.Y(n_1169)
);

AND2x4_ASAP7_75t_L g1170 ( 
.A(n_1057),
.B(n_1102),
.Y(n_1170)
);

AND2x4_ASAP7_75t_L g1171 ( 
.A(n_1140),
.B(n_1107),
.Y(n_1171)
);

AOI22xp33_ASAP7_75t_L g1172 ( 
.A1(n_1124),
.A2(n_1047),
.B1(n_1154),
.B2(n_1121),
.Y(n_1172)
);

OAI22xp5_ASAP7_75t_L g1173 ( 
.A1(n_1028),
.A2(n_1157),
.B1(n_1037),
.B2(n_1123),
.Y(n_1173)
);

INVx5_ASAP7_75t_L g1174 ( 
.A(n_1049),
.Y(n_1174)
);

AND2x4_ASAP7_75t_L g1175 ( 
.A(n_1140),
.B(n_1049),
.Y(n_1175)
);

NAND2xp5_ASAP7_75t_L g1176 ( 
.A(n_1123),
.B(n_1157),
.Y(n_1176)
);

AND2x4_ASAP7_75t_L g1177 ( 
.A(n_1049),
.B(n_1106),
.Y(n_1177)
);

AOI21xp5_ASAP7_75t_L g1178 ( 
.A1(n_1077),
.A2(n_1145),
.B(n_1038),
.Y(n_1178)
);

O2A1O1Ixp5_ASAP7_75t_L g1179 ( 
.A1(n_1088),
.A2(n_1121),
.B(n_1139),
.C(n_1117),
.Y(n_1179)
);

AND2x2_ASAP7_75t_L g1180 ( 
.A(n_1091),
.B(n_1034),
.Y(n_1180)
);

NAND2xp5_ASAP7_75t_SL g1181 ( 
.A(n_1040),
.B(n_1153),
.Y(n_1181)
);

INVx1_ASAP7_75t_L g1182 ( 
.A(n_1067),
.Y(n_1182)
);

NOR2xp33_ASAP7_75t_L g1183 ( 
.A(n_1120),
.B(n_1115),
.Y(n_1183)
);

AOI22xp33_ASAP7_75t_L g1184 ( 
.A1(n_1139),
.A2(n_1146),
.B1(n_1155),
.B2(n_1118),
.Y(n_1184)
);

OR2x2_ASAP7_75t_L g1185 ( 
.A(n_1065),
.B(n_1153),
.Y(n_1185)
);

AND2x4_ASAP7_75t_L g1186 ( 
.A(n_1041),
.B(n_1042),
.Y(n_1186)
);

A2O1A1Ixp33_ASAP7_75t_L g1187 ( 
.A1(n_1045),
.A2(n_1128),
.B(n_1115),
.C(n_1136),
.Y(n_1187)
);

BUFx6f_ASAP7_75t_L g1188 ( 
.A(n_1134),
.Y(n_1188)
);

NAND2xp5_ASAP7_75t_L g1189 ( 
.A(n_1128),
.B(n_1084),
.Y(n_1189)
);

AOI21xp5_ASAP7_75t_SL g1190 ( 
.A1(n_1122),
.A2(n_1129),
.B(n_1148),
.Y(n_1190)
);

A2O1A1Ixp33_ASAP7_75t_SL g1191 ( 
.A1(n_1113),
.A2(n_1052),
.B(n_1056),
.C(n_1093),
.Y(n_1191)
);

BUFx6f_ASAP7_75t_L g1192 ( 
.A(n_1134),
.Y(n_1192)
);

INVx3_ASAP7_75t_SL g1193 ( 
.A(n_1127),
.Y(n_1193)
);

NAND2xp5_ASAP7_75t_L g1194 ( 
.A(n_1084),
.B(n_1065),
.Y(n_1194)
);

BUFx6f_ASAP7_75t_L g1195 ( 
.A(n_1134),
.Y(n_1195)
);

OAI22xp5_ASAP7_75t_L g1196 ( 
.A1(n_1060),
.A2(n_1073),
.B1(n_1072),
.B2(n_1092),
.Y(n_1196)
);

NAND2xp5_ASAP7_75t_L g1197 ( 
.A(n_1137),
.B(n_1116),
.Y(n_1197)
);

AND2x4_ASAP7_75t_L g1198 ( 
.A(n_1132),
.B(n_1143),
.Y(n_1198)
);

O2A1O1Ixp5_ASAP7_75t_L g1199 ( 
.A1(n_1094),
.A2(n_1058),
.B(n_1066),
.C(n_1113),
.Y(n_1199)
);

OAI22xp5_ASAP7_75t_L g1200 ( 
.A1(n_1089),
.A2(n_1114),
.B1(n_1104),
.B2(n_1133),
.Y(n_1200)
);

INVx2_ASAP7_75t_L g1201 ( 
.A(n_1125),
.Y(n_1201)
);

NAND2xp5_ASAP7_75t_L g1202 ( 
.A(n_1116),
.B(n_1082),
.Y(n_1202)
);

NAND2xp5_ASAP7_75t_L g1203 ( 
.A(n_1082),
.B(n_1095),
.Y(n_1203)
);

INVx1_ASAP7_75t_SL g1204 ( 
.A(n_1099),
.Y(n_1204)
);

NOR2xp33_ASAP7_75t_SL g1205 ( 
.A(n_1108),
.B(n_1132),
.Y(n_1205)
);

CKINVDCx6p67_ASAP7_75t_R g1206 ( 
.A(n_1119),
.Y(n_1206)
);

INVx1_ASAP7_75t_L g1207 ( 
.A(n_1144),
.Y(n_1207)
);

INVx1_ASAP7_75t_L g1208 ( 
.A(n_1076),
.Y(n_1208)
);

OAI21xp33_ASAP7_75t_L g1209 ( 
.A1(n_1087),
.A2(n_1105),
.B(n_1083),
.Y(n_1209)
);

OAI22xp5_ASAP7_75t_L g1210 ( 
.A1(n_1104),
.A2(n_1105),
.B1(n_1052),
.B2(n_1087),
.Y(n_1210)
);

NOR2xp67_ASAP7_75t_L g1211 ( 
.A(n_1112),
.B(n_1061),
.Y(n_1211)
);

OAI21xp5_ASAP7_75t_L g1212 ( 
.A1(n_1059),
.A2(n_1056),
.B(n_1055),
.Y(n_1212)
);

INVx2_ASAP7_75t_SL g1213 ( 
.A(n_1085),
.Y(n_1213)
);

NOR2xp33_ASAP7_75t_L g1214 ( 
.A(n_1070),
.B(n_1080),
.Y(n_1214)
);

BUFx2_ASAP7_75t_SL g1215 ( 
.A(n_1061),
.Y(n_1215)
);

BUFx6f_ASAP7_75t_L g1216 ( 
.A(n_1143),
.Y(n_1216)
);

HB1xp67_ASAP7_75t_L g1217 ( 
.A(n_1097),
.Y(n_1217)
);

BUFx3_ASAP7_75t_L g1218 ( 
.A(n_1143),
.Y(n_1218)
);

INVx3_ASAP7_75t_L g1219 ( 
.A(n_1031),
.Y(n_1219)
);

NAND2xp5_ASAP7_75t_L g1220 ( 
.A(n_1051),
.B(n_1152),
.Y(n_1220)
);

AOI21xp5_ASAP7_75t_L g1221 ( 
.A1(n_1101),
.A2(n_1135),
.B(n_1111),
.Y(n_1221)
);

NAND2xp5_ASAP7_75t_L g1222 ( 
.A(n_1036),
.B(n_1152),
.Y(n_1222)
);

A2O1A1Ixp33_ASAP7_75t_L g1223 ( 
.A1(n_1108),
.A2(n_1093),
.B(n_1098),
.C(n_1103),
.Y(n_1223)
);

CKINVDCx6p67_ASAP7_75t_R g1224 ( 
.A(n_1075),
.Y(n_1224)
);

INVx3_ASAP7_75t_L g1225 ( 
.A(n_1031),
.Y(n_1225)
);

NAND2xp5_ASAP7_75t_L g1226 ( 
.A(n_1036),
.B(n_1152),
.Y(n_1226)
);

NOR2xp33_ASAP7_75t_L g1227 ( 
.A(n_1096),
.B(n_1109),
.Y(n_1227)
);

AOI21xp5_ASAP7_75t_L g1228 ( 
.A1(n_1030),
.A2(n_1069),
.B(n_1032),
.Y(n_1228)
);

AND2x2_ASAP7_75t_L g1229 ( 
.A(n_1036),
.B(n_1081),
.Y(n_1229)
);

OAI22xp5_ASAP7_75t_L g1230 ( 
.A1(n_1103),
.A2(n_1110),
.B1(n_1100),
.B2(n_1090),
.Y(n_1230)
);

NAND2xp5_ASAP7_75t_L g1231 ( 
.A(n_1075),
.B(n_1079),
.Y(n_1231)
);

HB1xp67_ASAP7_75t_L g1232 ( 
.A(n_1079),
.Y(n_1232)
);

AOI22xp33_ASAP7_75t_L g1233 ( 
.A1(n_1075),
.A2(n_1086),
.B1(n_1039),
.B2(n_1156),
.Y(n_1233)
);

CKINVDCx5p33_ASAP7_75t_R g1234 ( 
.A(n_1141),
.Y(n_1234)
);

NAND2xp5_ASAP7_75t_L g1235 ( 
.A(n_1075),
.B(n_1079),
.Y(n_1235)
);

INVx2_ASAP7_75t_SL g1236 ( 
.A(n_1039),
.Y(n_1236)
);

INVx2_ASAP7_75t_L g1237 ( 
.A(n_1053),
.Y(n_1237)
);

NOR2xp33_ASAP7_75t_L g1238 ( 
.A(n_1078),
.B(n_1142),
.Y(n_1238)
);

NOR2xp33_ASAP7_75t_L g1239 ( 
.A(n_1074),
.B(n_1150),
.Y(n_1239)
);

NOR2xp67_ASAP7_75t_L g1240 ( 
.A(n_1071),
.B(n_568),
.Y(n_1240)
);

AND2x4_ASAP7_75t_L g1241 ( 
.A(n_1057),
.B(n_1102),
.Y(n_1241)
);

OAI22xp5_ASAP7_75t_L g1242 ( 
.A1(n_1138),
.A2(n_1003),
.B1(n_1013),
.B2(n_1001),
.Y(n_1242)
);

INVx2_ASAP7_75t_SL g1243 ( 
.A(n_1043),
.Y(n_1243)
);

NAND2xp5_ASAP7_75t_L g1244 ( 
.A(n_1044),
.B(n_1138),
.Y(n_1244)
);

AOI21xp5_ASAP7_75t_L g1245 ( 
.A1(n_1063),
.A2(n_1077),
.B(n_1068),
.Y(n_1245)
);

INVx4_ASAP7_75t_L g1246 ( 
.A(n_1134),
.Y(n_1246)
);

NAND2xp5_ASAP7_75t_L g1247 ( 
.A(n_1044),
.B(n_1138),
.Y(n_1247)
);

BUFx3_ASAP7_75t_L g1248 ( 
.A(n_1043),
.Y(n_1248)
);

NAND2xp5_ASAP7_75t_L g1249 ( 
.A(n_1044),
.B(n_1138),
.Y(n_1249)
);

CKINVDCx20_ASAP7_75t_R g1250 ( 
.A(n_1127),
.Y(n_1250)
);

NAND2xp5_ASAP7_75t_L g1251 ( 
.A(n_1044),
.B(n_1138),
.Y(n_1251)
);

AOI22xp33_ASAP7_75t_L g1252 ( 
.A1(n_1124),
.A2(n_969),
.B1(n_1047),
.B2(n_717),
.Y(n_1252)
);

BUFx4f_ASAP7_75t_SL g1253 ( 
.A(n_1043),
.Y(n_1253)
);

AOI21xp5_ASAP7_75t_L g1254 ( 
.A1(n_1063),
.A2(n_1077),
.B(n_1068),
.Y(n_1254)
);

OR2x6_ASAP7_75t_L g1255 ( 
.A(n_1132),
.B(n_1143),
.Y(n_1255)
);

OAI22xp5_ASAP7_75t_L g1256 ( 
.A1(n_1138),
.A2(n_1003),
.B1(n_1013),
.B2(n_1001),
.Y(n_1256)
);

NAND2xp5_ASAP7_75t_L g1257 ( 
.A(n_1138),
.B(n_1028),
.Y(n_1257)
);

BUFx12f_ASAP7_75t_L g1258 ( 
.A(n_1081),
.Y(n_1258)
);

NOR2xp67_ASAP7_75t_L g1259 ( 
.A(n_1131),
.B(n_568),
.Y(n_1259)
);

INVx2_ASAP7_75t_SL g1260 ( 
.A(n_1043),
.Y(n_1260)
);

NAND2xp5_ASAP7_75t_L g1261 ( 
.A(n_1138),
.B(n_1028),
.Y(n_1261)
);

AOI22xp5_ASAP7_75t_L g1262 ( 
.A1(n_1124),
.A2(n_969),
.B1(n_1003),
.B2(n_1001),
.Y(n_1262)
);

CKINVDCx20_ASAP7_75t_R g1263 ( 
.A(n_1127),
.Y(n_1263)
);

AOI21xp5_ASAP7_75t_L g1264 ( 
.A1(n_1063),
.A2(n_1077),
.B(n_1068),
.Y(n_1264)
);

NAND2xp33_ASAP7_75t_L g1265 ( 
.A(n_1124),
.B(n_1020),
.Y(n_1265)
);

AO21x2_ASAP7_75t_L g1266 ( 
.A1(n_1077),
.A2(n_1145),
.B(n_1038),
.Y(n_1266)
);

NAND2xp5_ASAP7_75t_L g1267 ( 
.A(n_1138),
.B(n_1028),
.Y(n_1267)
);

NAND2xp5_ASAP7_75t_L g1268 ( 
.A(n_1138),
.B(n_1028),
.Y(n_1268)
);

CKINVDCx6p67_ASAP7_75t_R g1269 ( 
.A(n_1043),
.Y(n_1269)
);

INVxp67_ASAP7_75t_SL g1270 ( 
.A(n_1043),
.Y(n_1270)
);

BUFx6f_ASAP7_75t_L g1271 ( 
.A(n_1134),
.Y(n_1271)
);

AND2x4_ASAP7_75t_L g1272 ( 
.A(n_1057),
.B(n_1102),
.Y(n_1272)
);

NAND2x1p5_ASAP7_75t_L g1273 ( 
.A(n_1092),
.B(n_892),
.Y(n_1273)
);

INVx2_ASAP7_75t_SL g1274 ( 
.A(n_1043),
.Y(n_1274)
);

AND2x4_ASAP7_75t_L g1275 ( 
.A(n_1057),
.B(n_1102),
.Y(n_1275)
);

NAND2x1p5_ASAP7_75t_L g1276 ( 
.A(n_1092),
.B(n_892),
.Y(n_1276)
);

BUFx3_ASAP7_75t_L g1277 ( 
.A(n_1043),
.Y(n_1277)
);

HB1xp67_ASAP7_75t_L g1278 ( 
.A(n_1153),
.Y(n_1278)
);

NAND2xp5_ASAP7_75t_L g1279 ( 
.A(n_1044),
.B(n_1138),
.Y(n_1279)
);

BUFx6f_ASAP7_75t_L g1280 ( 
.A(n_1134),
.Y(n_1280)
);

AOI21xp5_ASAP7_75t_SL g1281 ( 
.A1(n_1121),
.A2(n_1020),
.B(n_1139),
.Y(n_1281)
);

INVxp67_ASAP7_75t_SL g1282 ( 
.A(n_1043),
.Y(n_1282)
);

INVx3_ASAP7_75t_L g1283 ( 
.A(n_1033),
.Y(n_1283)
);

INVx3_ASAP7_75t_L g1284 ( 
.A(n_1033),
.Y(n_1284)
);

AND2x2_ASAP7_75t_L g1285 ( 
.A(n_1130),
.B(n_1147),
.Y(n_1285)
);

INVx1_ASAP7_75t_L g1286 ( 
.A(n_1064),
.Y(n_1286)
);

OR2x2_ASAP7_75t_L g1287 ( 
.A(n_1048),
.B(n_1046),
.Y(n_1287)
);

INVx1_ASAP7_75t_L g1288 ( 
.A(n_1064),
.Y(n_1288)
);

AND2x4_ASAP7_75t_L g1289 ( 
.A(n_1057),
.B(n_1102),
.Y(n_1289)
);

NAND2xp5_ASAP7_75t_L g1290 ( 
.A(n_1044),
.B(n_1138),
.Y(n_1290)
);

AND2x4_ASAP7_75t_L g1291 ( 
.A(n_1057),
.B(n_1102),
.Y(n_1291)
);

AOI22xp5_ASAP7_75t_L g1292 ( 
.A1(n_1124),
.A2(n_969),
.B1(n_1003),
.B2(n_1001),
.Y(n_1292)
);

OAI22xp33_ASAP7_75t_L g1293 ( 
.A1(n_1138),
.A2(n_1003),
.B1(n_1013),
.B2(n_1001),
.Y(n_1293)
);

AO21x2_ASAP7_75t_L g1294 ( 
.A1(n_1221),
.A2(n_1228),
.B(n_1165),
.Y(n_1294)
);

AOI22xp33_ASAP7_75t_SL g1295 ( 
.A1(n_1164),
.A2(n_1251),
.B1(n_1249),
.B2(n_1279),
.Y(n_1295)
);

INVx2_ASAP7_75t_SL g1296 ( 
.A(n_1174),
.Y(n_1296)
);

CKINVDCx5p33_ASAP7_75t_R g1297 ( 
.A(n_1234),
.Y(n_1297)
);

AO21x2_ASAP7_75t_L g1298 ( 
.A1(n_1245),
.A2(n_1264),
.B(n_1254),
.Y(n_1298)
);

AO21x1_ASAP7_75t_SL g1299 ( 
.A1(n_1172),
.A2(n_1220),
.B(n_1231),
.Y(n_1299)
);

HB1xp67_ASAP7_75t_L g1300 ( 
.A(n_1278),
.Y(n_1300)
);

AOI22xp33_ASAP7_75t_L g1301 ( 
.A1(n_1252),
.A2(n_1184),
.B1(n_1290),
.B2(n_1247),
.Y(n_1301)
);

BUFx6f_ASAP7_75t_L g1302 ( 
.A(n_1175),
.Y(n_1302)
);

NAND2x1p5_ASAP7_75t_L g1303 ( 
.A(n_1174),
.B(n_1167),
.Y(n_1303)
);

INVx1_ASAP7_75t_L g1304 ( 
.A(n_1182),
.Y(n_1304)
);

INVx1_ASAP7_75t_L g1305 ( 
.A(n_1207),
.Y(n_1305)
);

BUFx4f_ASAP7_75t_L g1306 ( 
.A(n_1175),
.Y(n_1306)
);

INVx2_ASAP7_75t_L g1307 ( 
.A(n_1208),
.Y(n_1307)
);

BUFx6f_ASAP7_75t_L g1308 ( 
.A(n_1174),
.Y(n_1308)
);

BUFx3_ASAP7_75t_L g1309 ( 
.A(n_1248),
.Y(n_1309)
);

AND2x2_ASAP7_75t_L g1310 ( 
.A(n_1183),
.B(n_1166),
.Y(n_1310)
);

BUFx6f_ASAP7_75t_L g1311 ( 
.A(n_1188),
.Y(n_1311)
);

OR2x2_ASAP7_75t_L g1312 ( 
.A(n_1266),
.B(n_1222),
.Y(n_1312)
);

INVxp67_ASAP7_75t_SL g1313 ( 
.A(n_1194),
.Y(n_1313)
);

AND2x4_ASAP7_75t_L g1314 ( 
.A(n_1177),
.B(n_1198),
.Y(n_1314)
);

INVx2_ASAP7_75t_L g1315 ( 
.A(n_1286),
.Y(n_1315)
);

AND2x2_ASAP7_75t_L g1316 ( 
.A(n_1166),
.B(n_1176),
.Y(n_1316)
);

INVx1_ASAP7_75t_L g1317 ( 
.A(n_1288),
.Y(n_1317)
);

AO21x1_ASAP7_75t_SL g1318 ( 
.A1(n_1235),
.A2(n_1197),
.B(n_1226),
.Y(n_1318)
);

HB1xp67_ASAP7_75t_L g1319 ( 
.A(n_1185),
.Y(n_1319)
);

OA21x2_ASAP7_75t_L g1320 ( 
.A1(n_1199),
.A2(n_1179),
.B(n_1212),
.Y(n_1320)
);

AND2x4_ASAP7_75t_L g1321 ( 
.A(n_1177),
.B(n_1198),
.Y(n_1321)
);

BUFx2_ASAP7_75t_R g1322 ( 
.A(n_1193),
.Y(n_1322)
);

AOI22xp33_ASAP7_75t_L g1323 ( 
.A1(n_1244),
.A2(n_1265),
.B1(n_1196),
.B2(n_1168),
.Y(n_1323)
);

OAI22xp33_ASAP7_75t_L g1324 ( 
.A1(n_1205),
.A2(n_1261),
.B1(n_1257),
.B2(n_1268),
.Y(n_1324)
);

OAI22xp5_ASAP7_75t_L g1325 ( 
.A1(n_1176),
.A2(n_1257),
.B1(n_1268),
.B2(n_1267),
.Y(n_1325)
);

CKINVDCx8_ASAP7_75t_R g1326 ( 
.A(n_1215),
.Y(n_1326)
);

INVx1_ASAP7_75t_SL g1327 ( 
.A(n_1204),
.Y(n_1327)
);

BUFx10_ASAP7_75t_L g1328 ( 
.A(n_1186),
.Y(n_1328)
);

NAND2x1p5_ASAP7_75t_L g1329 ( 
.A(n_1158),
.B(n_1283),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_1285),
.Y(n_1330)
);

INVx1_ASAP7_75t_L g1331 ( 
.A(n_1217),
.Y(n_1331)
);

INVx1_ASAP7_75t_SL g1332 ( 
.A(n_1204),
.Y(n_1332)
);

NOR2x1_ASAP7_75t_R g1333 ( 
.A(n_1258),
.B(n_1277),
.Y(n_1333)
);

INVx3_ASAP7_75t_L g1334 ( 
.A(n_1273),
.Y(n_1334)
);

NOR2xp33_ASAP7_75t_L g1335 ( 
.A(n_1163),
.B(n_1169),
.Y(n_1335)
);

OAI22xp33_ASAP7_75t_L g1336 ( 
.A1(n_1205),
.A2(n_1262),
.B1(n_1292),
.B2(n_1189),
.Y(n_1336)
);

AO21x1_ASAP7_75t_SL g1337 ( 
.A1(n_1226),
.A2(n_1202),
.B(n_1232),
.Y(n_1337)
);

INVx1_ASAP7_75t_L g1338 ( 
.A(n_1180),
.Y(n_1338)
);

OAI21x1_ASAP7_75t_L g1339 ( 
.A1(n_1230),
.A2(n_1178),
.B(n_1233),
.Y(n_1339)
);

NAND2xp5_ASAP7_75t_L g1340 ( 
.A(n_1173),
.B(n_1293),
.Y(n_1340)
);

INVx1_ASAP7_75t_L g1341 ( 
.A(n_1287),
.Y(n_1341)
);

INVx2_ASAP7_75t_L g1342 ( 
.A(n_1202),
.Y(n_1342)
);

INVx11_ASAP7_75t_L g1343 ( 
.A(n_1253),
.Y(n_1343)
);

INVxp67_ASAP7_75t_L g1344 ( 
.A(n_1270),
.Y(n_1344)
);

AND2x2_ASAP7_75t_L g1345 ( 
.A(n_1262),
.B(n_1292),
.Y(n_1345)
);

OAI21xp5_ASAP7_75t_L g1346 ( 
.A1(n_1187),
.A2(n_1256),
.B(n_1242),
.Y(n_1346)
);

AOI22xp33_ASAP7_75t_L g1347 ( 
.A1(n_1181),
.A2(n_1242),
.B1(n_1256),
.B2(n_1209),
.Y(n_1347)
);

OAI21xp5_ASAP7_75t_L g1348 ( 
.A1(n_1281),
.A2(n_1223),
.B(n_1209),
.Y(n_1348)
);

INVx1_ASAP7_75t_L g1349 ( 
.A(n_1203),
.Y(n_1349)
);

OA21x2_ASAP7_75t_L g1350 ( 
.A1(n_1200),
.A2(n_1210),
.B(n_1238),
.Y(n_1350)
);

HB1xp67_ASAP7_75t_L g1351 ( 
.A(n_1282),
.Y(n_1351)
);

INVx1_ASAP7_75t_L g1352 ( 
.A(n_1200),
.Y(n_1352)
);

AOI22xp33_ASAP7_75t_L g1353 ( 
.A1(n_1214),
.A2(n_1210),
.B1(n_1229),
.B2(n_1227),
.Y(n_1353)
);

INVx1_ASAP7_75t_L g1354 ( 
.A(n_1237),
.Y(n_1354)
);

AOI22xp33_ASAP7_75t_SL g1355 ( 
.A1(n_1239),
.A2(n_1216),
.B1(n_1159),
.B2(n_1218),
.Y(n_1355)
);

INVx2_ASAP7_75t_L g1356 ( 
.A(n_1190),
.Y(n_1356)
);

AOI22xp5_ASAP7_75t_L g1357 ( 
.A1(n_1240),
.A2(n_1259),
.B1(n_1269),
.B2(n_1250),
.Y(n_1357)
);

NAND2x1p5_ASAP7_75t_L g1358 ( 
.A(n_1219),
.B(n_1225),
.Y(n_1358)
);

HB1xp67_ASAP7_75t_L g1359 ( 
.A(n_1161),
.Y(n_1359)
);

AOI22xp33_ASAP7_75t_L g1360 ( 
.A1(n_1224),
.A2(n_1206),
.B1(n_1213),
.B2(n_1255),
.Y(n_1360)
);

INVx6_ASAP7_75t_L g1361 ( 
.A(n_1171),
.Y(n_1361)
);

BUFx3_ASAP7_75t_L g1362 ( 
.A(n_1186),
.Y(n_1362)
);

INVx2_ASAP7_75t_L g1363 ( 
.A(n_1158),
.Y(n_1363)
);

OA21x2_ASAP7_75t_L g1364 ( 
.A1(n_1191),
.A2(n_1211),
.B(n_1291),
.Y(n_1364)
);

INVx1_ASAP7_75t_L g1365 ( 
.A(n_1160),
.Y(n_1365)
);

INVx1_ASAP7_75t_L g1366 ( 
.A(n_1160),
.Y(n_1366)
);

BUFx12f_ASAP7_75t_L g1367 ( 
.A(n_1243),
.Y(n_1367)
);

INVx1_ASAP7_75t_L g1368 ( 
.A(n_1170),
.Y(n_1368)
);

INVx1_ASAP7_75t_L g1369 ( 
.A(n_1170),
.Y(n_1369)
);

INVx1_ASAP7_75t_SL g1370 ( 
.A(n_1260),
.Y(n_1370)
);

INVx1_ASAP7_75t_L g1371 ( 
.A(n_1241),
.Y(n_1371)
);

INVx1_ASAP7_75t_L g1372 ( 
.A(n_1241),
.Y(n_1372)
);

CKINVDCx20_ASAP7_75t_R g1373 ( 
.A(n_1263),
.Y(n_1373)
);

AOI22xp33_ASAP7_75t_L g1374 ( 
.A1(n_1255),
.A2(n_1272),
.B1(n_1289),
.B2(n_1275),
.Y(n_1374)
);

HB1xp67_ASAP7_75t_L g1375 ( 
.A(n_1274),
.Y(n_1375)
);

OAI21x1_ASAP7_75t_L g1376 ( 
.A1(n_1284),
.A2(n_1273),
.B(n_1276),
.Y(n_1376)
);

OAI21xp5_ASAP7_75t_L g1377 ( 
.A1(n_1284),
.A2(n_1276),
.B(n_1171),
.Y(n_1377)
);

AOI21x1_ASAP7_75t_L g1378 ( 
.A1(n_1255),
.A2(n_1291),
.B(n_1289),
.Y(n_1378)
);

HB1xp67_ASAP7_75t_L g1379 ( 
.A(n_1272),
.Y(n_1379)
);

INVx2_ASAP7_75t_L g1380 ( 
.A(n_1275),
.Y(n_1380)
);

OAI22xp5_ASAP7_75t_L g1381 ( 
.A1(n_1216),
.A2(n_1162),
.B1(n_1236),
.B2(n_1246),
.Y(n_1381)
);

AND2x4_ASAP7_75t_L g1382 ( 
.A(n_1216),
.B(n_1246),
.Y(n_1382)
);

CKINVDCx20_ASAP7_75t_R g1383 ( 
.A(n_1192),
.Y(n_1383)
);

BUFx8_ASAP7_75t_SL g1384 ( 
.A(n_1195),
.Y(n_1384)
);

AND2x2_ASAP7_75t_L g1385 ( 
.A(n_1280),
.B(n_1195),
.Y(n_1385)
);

AND2x2_ASAP7_75t_L g1386 ( 
.A(n_1271),
.B(n_1280),
.Y(n_1386)
);

AOI22xp33_ASAP7_75t_L g1387 ( 
.A1(n_1271),
.A2(n_1124),
.B1(n_969),
.B2(n_1047),
.Y(n_1387)
);

CKINVDCx5p33_ASAP7_75t_R g1388 ( 
.A(n_1280),
.Y(n_1388)
);

AOI22xp33_ASAP7_75t_L g1389 ( 
.A1(n_1252),
.A2(n_1124),
.B1(n_969),
.B2(n_1047),
.Y(n_1389)
);

CKINVDCx11_ASAP7_75t_R g1390 ( 
.A(n_1250),
.Y(n_1390)
);

INVx1_ASAP7_75t_L g1391 ( 
.A(n_1201),
.Y(n_1391)
);

AND2x2_ASAP7_75t_L g1392 ( 
.A(n_1183),
.B(n_1184),
.Y(n_1392)
);

BUFx3_ASAP7_75t_L g1393 ( 
.A(n_1248),
.Y(n_1393)
);

AOI22xp33_ASAP7_75t_SL g1394 ( 
.A1(n_1164),
.A2(n_969),
.B1(n_386),
.B2(n_406),
.Y(n_1394)
);

AOI21xp5_ASAP7_75t_SL g1395 ( 
.A1(n_1223),
.A2(n_1020),
.B(n_1121),
.Y(n_1395)
);

INVx1_ASAP7_75t_L g1396 ( 
.A(n_1201),
.Y(n_1396)
);

INVx2_ASAP7_75t_SL g1397 ( 
.A(n_1174),
.Y(n_1397)
);

BUFx3_ASAP7_75t_L g1398 ( 
.A(n_1248),
.Y(n_1398)
);

INVx1_ASAP7_75t_L g1399 ( 
.A(n_1201),
.Y(n_1399)
);

HB1xp67_ASAP7_75t_L g1400 ( 
.A(n_1278),
.Y(n_1400)
);

BUFx4f_ASAP7_75t_SL g1401 ( 
.A(n_1258),
.Y(n_1401)
);

OAI22xp5_ASAP7_75t_L g1402 ( 
.A1(n_1164),
.A2(n_1003),
.B1(n_1013),
.B2(n_1001),
.Y(n_1402)
);

BUFx3_ASAP7_75t_L g1403 ( 
.A(n_1248),
.Y(n_1403)
);

AND2x4_ASAP7_75t_L g1404 ( 
.A(n_1177),
.B(n_1198),
.Y(n_1404)
);

INVxp67_ASAP7_75t_L g1405 ( 
.A(n_1278),
.Y(n_1405)
);

INVx2_ASAP7_75t_L g1406 ( 
.A(n_1201),
.Y(n_1406)
);

INVx4_ASAP7_75t_SL g1407 ( 
.A(n_1255),
.Y(n_1407)
);

INVx2_ASAP7_75t_L g1408 ( 
.A(n_1201),
.Y(n_1408)
);

INVx4_ASAP7_75t_L g1409 ( 
.A(n_1174),
.Y(n_1409)
);

HB1xp67_ASAP7_75t_L g1410 ( 
.A(n_1278),
.Y(n_1410)
);

AOI22xp33_ASAP7_75t_L g1411 ( 
.A1(n_1252),
.A2(n_1124),
.B1(n_969),
.B2(n_1047),
.Y(n_1411)
);

HB1xp67_ASAP7_75t_L g1412 ( 
.A(n_1351),
.Y(n_1412)
);

BUFx12f_ASAP7_75t_L g1413 ( 
.A(n_1390),
.Y(n_1413)
);

BUFx2_ASAP7_75t_L g1414 ( 
.A(n_1312),
.Y(n_1414)
);

AND2x2_ASAP7_75t_L g1415 ( 
.A(n_1310),
.B(n_1392),
.Y(n_1415)
);

INVx1_ASAP7_75t_L g1416 ( 
.A(n_1312),
.Y(n_1416)
);

NAND2xp5_ASAP7_75t_L g1417 ( 
.A(n_1295),
.B(n_1313),
.Y(n_1417)
);

BUFx3_ASAP7_75t_L g1418 ( 
.A(n_1384),
.Y(n_1418)
);

AND2x2_ASAP7_75t_L g1419 ( 
.A(n_1345),
.B(n_1316),
.Y(n_1419)
);

AND2x4_ASAP7_75t_L g1420 ( 
.A(n_1407),
.B(n_1378),
.Y(n_1420)
);

OA21x2_ASAP7_75t_L g1421 ( 
.A1(n_1339),
.A2(n_1346),
.B(n_1348),
.Y(n_1421)
);

OR2x2_ASAP7_75t_L g1422 ( 
.A(n_1350),
.B(n_1340),
.Y(n_1422)
);

INVx1_ASAP7_75t_L g1423 ( 
.A(n_1352),
.Y(n_1423)
);

INVx4_ASAP7_75t_L g1424 ( 
.A(n_1407),
.Y(n_1424)
);

CKINVDCx5p33_ASAP7_75t_R g1425 ( 
.A(n_1390),
.Y(n_1425)
);

HB1xp67_ASAP7_75t_L g1426 ( 
.A(n_1319),
.Y(n_1426)
);

INVx1_ASAP7_75t_L g1427 ( 
.A(n_1307),
.Y(n_1427)
);

OAI21xp5_ASAP7_75t_L g1428 ( 
.A1(n_1389),
.A2(n_1411),
.B(n_1402),
.Y(n_1428)
);

CKINVDCx20_ASAP7_75t_R g1429 ( 
.A(n_1373),
.Y(n_1429)
);

INVx1_ASAP7_75t_L g1430 ( 
.A(n_1315),
.Y(n_1430)
);

AO21x2_ASAP7_75t_L g1431 ( 
.A1(n_1294),
.A2(n_1395),
.B(n_1298),
.Y(n_1431)
);

AND2x2_ASAP7_75t_L g1432 ( 
.A(n_1345),
.B(n_1316),
.Y(n_1432)
);

INVx1_ASAP7_75t_SL g1433 ( 
.A(n_1327),
.Y(n_1433)
);

HB1xp67_ASAP7_75t_L g1434 ( 
.A(n_1300),
.Y(n_1434)
);

BUFx2_ASAP7_75t_L g1435 ( 
.A(n_1364),
.Y(n_1435)
);

OR2x2_ASAP7_75t_L g1436 ( 
.A(n_1350),
.B(n_1325),
.Y(n_1436)
);

OA21x2_ASAP7_75t_L g1437 ( 
.A1(n_1347),
.A2(n_1342),
.B(n_1323),
.Y(n_1437)
);

BUFx3_ASAP7_75t_L g1438 ( 
.A(n_1384),
.Y(n_1438)
);

AND2x2_ASAP7_75t_L g1439 ( 
.A(n_1318),
.B(n_1299),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_1320),
.Y(n_1440)
);

INVx1_ASAP7_75t_L g1441 ( 
.A(n_1320),
.Y(n_1441)
);

OA21x2_ASAP7_75t_L g1442 ( 
.A1(n_1387),
.A2(n_1301),
.B(n_1349),
.Y(n_1442)
);

OA21x2_ASAP7_75t_L g1443 ( 
.A1(n_1356),
.A2(n_1353),
.B(n_1305),
.Y(n_1443)
);

HB1xp67_ASAP7_75t_L g1444 ( 
.A(n_1400),
.Y(n_1444)
);

INVx1_ASAP7_75t_L g1445 ( 
.A(n_1304),
.Y(n_1445)
);

AND2x4_ASAP7_75t_L g1446 ( 
.A(n_1407),
.B(n_1378),
.Y(n_1446)
);

OAI21xp5_ASAP7_75t_L g1447 ( 
.A1(n_1395),
.A2(n_1394),
.B(n_1324),
.Y(n_1447)
);

AO21x2_ASAP7_75t_L g1448 ( 
.A1(n_1294),
.A2(n_1298),
.B(n_1336),
.Y(n_1448)
);

INVx2_ASAP7_75t_SL g1449 ( 
.A(n_1328),
.Y(n_1449)
);

OA21x2_ASAP7_75t_L g1450 ( 
.A1(n_1356),
.A2(n_1317),
.B(n_1408),
.Y(n_1450)
);

BUFx2_ASAP7_75t_R g1451 ( 
.A(n_1297),
.Y(n_1451)
);

NAND3xp33_ASAP7_75t_L g1452 ( 
.A(n_1355),
.B(n_1335),
.C(n_1344),
.Y(n_1452)
);

AND2x2_ASAP7_75t_L g1453 ( 
.A(n_1318),
.B(n_1299),
.Y(n_1453)
);

HB1xp67_ASAP7_75t_L g1454 ( 
.A(n_1410),
.Y(n_1454)
);

OR2x2_ASAP7_75t_L g1455 ( 
.A(n_1338),
.B(n_1298),
.Y(n_1455)
);

OR2x2_ASAP7_75t_L g1456 ( 
.A(n_1331),
.B(n_1341),
.Y(n_1456)
);

AND2x4_ASAP7_75t_L g1457 ( 
.A(n_1407),
.B(n_1377),
.Y(n_1457)
);

AND2x2_ASAP7_75t_L g1458 ( 
.A(n_1337),
.B(n_1406),
.Y(n_1458)
);

BUFx4f_ASAP7_75t_SL g1459 ( 
.A(n_1373),
.Y(n_1459)
);

INVx1_ASAP7_75t_L g1460 ( 
.A(n_1391),
.Y(n_1460)
);

OAI21xp5_ASAP7_75t_L g1461 ( 
.A1(n_1405),
.A2(n_1354),
.B(n_1303),
.Y(n_1461)
);

INVx1_ASAP7_75t_L g1462 ( 
.A(n_1396),
.Y(n_1462)
);

INVx1_ASAP7_75t_L g1463 ( 
.A(n_1399),
.Y(n_1463)
);

OR2x6_ASAP7_75t_L g1464 ( 
.A(n_1376),
.B(n_1409),
.Y(n_1464)
);

OAI21x1_ASAP7_75t_L g1465 ( 
.A1(n_1376),
.A2(n_1329),
.B(n_1363),
.Y(n_1465)
);

BUFx3_ASAP7_75t_L g1466 ( 
.A(n_1309),
.Y(n_1466)
);

INVx1_ASAP7_75t_SL g1467 ( 
.A(n_1332),
.Y(n_1467)
);

AND2x2_ASAP7_75t_L g1468 ( 
.A(n_1330),
.B(n_1314),
.Y(n_1468)
);

AND2x2_ASAP7_75t_L g1469 ( 
.A(n_1314),
.B(n_1404),
.Y(n_1469)
);

NAND2xp5_ASAP7_75t_SL g1470 ( 
.A(n_1306),
.B(n_1314),
.Y(n_1470)
);

OR2x2_ASAP7_75t_L g1471 ( 
.A(n_1321),
.B(n_1404),
.Y(n_1471)
);

AND2x2_ASAP7_75t_L g1472 ( 
.A(n_1321),
.B(n_1404),
.Y(n_1472)
);

INVx1_ASAP7_75t_L g1473 ( 
.A(n_1296),
.Y(n_1473)
);

NAND2xp5_ASAP7_75t_L g1474 ( 
.A(n_1380),
.B(n_1379),
.Y(n_1474)
);

INVx1_ASAP7_75t_L g1475 ( 
.A(n_1296),
.Y(n_1475)
);

OR2x2_ASAP7_75t_L g1476 ( 
.A(n_1321),
.B(n_1380),
.Y(n_1476)
);

CKINVDCx6p67_ASAP7_75t_R g1477 ( 
.A(n_1309),
.Y(n_1477)
);

AND2x2_ASAP7_75t_L g1478 ( 
.A(n_1365),
.B(n_1369),
.Y(n_1478)
);

INVx1_ASAP7_75t_L g1479 ( 
.A(n_1397),
.Y(n_1479)
);

OAI21x1_ASAP7_75t_L g1480 ( 
.A1(n_1334),
.A2(n_1358),
.B(n_1360),
.Y(n_1480)
);

NAND2xp5_ASAP7_75t_L g1481 ( 
.A(n_1366),
.B(n_1372),
.Y(n_1481)
);

OR2x2_ASAP7_75t_L g1482 ( 
.A(n_1368),
.B(n_1371),
.Y(n_1482)
);

AND2x4_ASAP7_75t_L g1483 ( 
.A(n_1420),
.B(n_1409),
.Y(n_1483)
);

AND2x2_ASAP7_75t_L g1484 ( 
.A(n_1419),
.B(n_1385),
.Y(n_1484)
);

BUFx2_ASAP7_75t_L g1485 ( 
.A(n_1414),
.Y(n_1485)
);

INVx3_ASAP7_75t_L g1486 ( 
.A(n_1465),
.Y(n_1486)
);

AND2x2_ASAP7_75t_L g1487 ( 
.A(n_1419),
.B(n_1385),
.Y(n_1487)
);

AND2x2_ASAP7_75t_L g1488 ( 
.A(n_1432),
.B(n_1386),
.Y(n_1488)
);

INVx2_ASAP7_75t_L g1489 ( 
.A(n_1450),
.Y(n_1489)
);

INVx2_ASAP7_75t_L g1490 ( 
.A(n_1450),
.Y(n_1490)
);

INVx2_ASAP7_75t_L g1491 ( 
.A(n_1450),
.Y(n_1491)
);

NOR2xp33_ASAP7_75t_L g1492 ( 
.A(n_1459),
.B(n_1297),
.Y(n_1492)
);

NAND2xp5_ASAP7_75t_L g1493 ( 
.A(n_1416),
.B(n_1308),
.Y(n_1493)
);

AND2x4_ASAP7_75t_L g1494 ( 
.A(n_1420),
.B(n_1409),
.Y(n_1494)
);

OR2x6_ASAP7_75t_L g1495 ( 
.A(n_1420),
.B(n_1302),
.Y(n_1495)
);

BUFx2_ASAP7_75t_L g1496 ( 
.A(n_1458),
.Y(n_1496)
);

NOR2x1_ASAP7_75t_SL g1497 ( 
.A(n_1464),
.B(n_1367),
.Y(n_1497)
);

NAND2xp5_ASAP7_75t_L g1498 ( 
.A(n_1416),
.B(n_1375),
.Y(n_1498)
);

BUFx3_ASAP7_75t_L g1499 ( 
.A(n_1420),
.Y(n_1499)
);

NAND2xp5_ASAP7_75t_L g1500 ( 
.A(n_1415),
.B(n_1359),
.Y(n_1500)
);

NAND2xp5_ASAP7_75t_L g1501 ( 
.A(n_1423),
.B(n_1362),
.Y(n_1501)
);

INVx2_ASAP7_75t_SL g1502 ( 
.A(n_1412),
.Y(n_1502)
);

NOR2xp33_ASAP7_75t_L g1503 ( 
.A(n_1429),
.B(n_1370),
.Y(n_1503)
);

AND2x2_ASAP7_75t_L g1504 ( 
.A(n_1421),
.B(n_1306),
.Y(n_1504)
);

AND2x2_ASAP7_75t_L g1505 ( 
.A(n_1421),
.B(n_1306),
.Y(n_1505)
);

BUFx3_ASAP7_75t_L g1506 ( 
.A(n_1446),
.Y(n_1506)
);

AND2x2_ASAP7_75t_L g1507 ( 
.A(n_1421),
.B(n_1382),
.Y(n_1507)
);

AOI221xp5_ASAP7_75t_L g1508 ( 
.A1(n_1428),
.A2(n_1381),
.B1(n_1374),
.B2(n_1403),
.C(n_1398),
.Y(n_1508)
);

BUFx3_ASAP7_75t_L g1509 ( 
.A(n_1446),
.Y(n_1509)
);

OR2x2_ASAP7_75t_L g1510 ( 
.A(n_1455),
.B(n_1403),
.Y(n_1510)
);

AND2x4_ASAP7_75t_L g1511 ( 
.A(n_1464),
.B(n_1382),
.Y(n_1511)
);

AND2x2_ASAP7_75t_L g1512 ( 
.A(n_1455),
.B(n_1311),
.Y(n_1512)
);

AOI22xp5_ASAP7_75t_L g1513 ( 
.A1(n_1447),
.A2(n_1361),
.B1(n_1357),
.B2(n_1383),
.Y(n_1513)
);

HB1xp67_ASAP7_75t_L g1514 ( 
.A(n_1426),
.Y(n_1514)
);

OR2x2_ASAP7_75t_L g1515 ( 
.A(n_1422),
.B(n_1398),
.Y(n_1515)
);

OAI221xp5_ASAP7_75t_L g1516 ( 
.A1(n_1417),
.A2(n_1326),
.B1(n_1361),
.B2(n_1393),
.C(n_1388),
.Y(n_1516)
);

OAI22xp33_ASAP7_75t_L g1517 ( 
.A1(n_1452),
.A2(n_1326),
.B1(n_1361),
.B2(n_1393),
.Y(n_1517)
);

INVxp67_ASAP7_75t_SL g1518 ( 
.A(n_1434),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_1445),
.Y(n_1519)
);

INVx2_ASAP7_75t_L g1520 ( 
.A(n_1440),
.Y(n_1520)
);

NOR2xp33_ASAP7_75t_L g1521 ( 
.A(n_1433),
.B(n_1322),
.Y(n_1521)
);

INVx2_ASAP7_75t_L g1522 ( 
.A(n_1440),
.Y(n_1522)
);

HB1xp67_ASAP7_75t_L g1523 ( 
.A(n_1444),
.Y(n_1523)
);

NOR2xp33_ASAP7_75t_L g1524 ( 
.A(n_1467),
.B(n_1361),
.Y(n_1524)
);

BUFx3_ASAP7_75t_L g1525 ( 
.A(n_1480),
.Y(n_1525)
);

INVx2_ASAP7_75t_L g1526 ( 
.A(n_1441),
.Y(n_1526)
);

INVxp67_ASAP7_75t_L g1527 ( 
.A(n_1454),
.Y(n_1527)
);

BUFx2_ASAP7_75t_L g1528 ( 
.A(n_1464),
.Y(n_1528)
);

BUFx4f_ASAP7_75t_SL g1529 ( 
.A(n_1413),
.Y(n_1529)
);

AND2x2_ASAP7_75t_L g1530 ( 
.A(n_1496),
.B(n_1435),
.Y(n_1530)
);

NAND2xp5_ASAP7_75t_L g1531 ( 
.A(n_1514),
.B(n_1442),
.Y(n_1531)
);

NAND3xp33_ASAP7_75t_L g1532 ( 
.A(n_1508),
.B(n_1452),
.C(n_1461),
.Y(n_1532)
);

NAND2xp5_ASAP7_75t_L g1533 ( 
.A(n_1518),
.B(n_1442),
.Y(n_1533)
);

AND2x2_ASAP7_75t_L g1534 ( 
.A(n_1512),
.B(n_1507),
.Y(n_1534)
);

AOI22xp33_ASAP7_75t_L g1535 ( 
.A1(n_1517),
.A2(n_1442),
.B1(n_1439),
.B2(n_1453),
.Y(n_1535)
);

NOR2xp67_ASAP7_75t_L g1536 ( 
.A(n_1520),
.B(n_1441),
.Y(n_1536)
);

NAND3xp33_ASAP7_75t_L g1537 ( 
.A(n_1508),
.B(n_1442),
.C(n_1481),
.Y(n_1537)
);

AND2x2_ASAP7_75t_SL g1538 ( 
.A(n_1504),
.B(n_1505),
.Y(n_1538)
);

AOI22xp33_ASAP7_75t_L g1539 ( 
.A1(n_1516),
.A2(n_1439),
.B1(n_1453),
.B2(n_1457),
.Y(n_1539)
);

NAND2xp5_ASAP7_75t_L g1540 ( 
.A(n_1523),
.B(n_1456),
.Y(n_1540)
);

NAND2xp5_ASAP7_75t_L g1541 ( 
.A(n_1527),
.B(n_1502),
.Y(n_1541)
);

OAI21xp5_ASAP7_75t_SL g1542 ( 
.A1(n_1513),
.A2(n_1457),
.B(n_1470),
.Y(n_1542)
);

NAND2xp5_ASAP7_75t_L g1543 ( 
.A(n_1502),
.B(n_1456),
.Y(n_1543)
);

INVx1_ASAP7_75t_L g1544 ( 
.A(n_1519),
.Y(n_1544)
);

AOI22xp33_ASAP7_75t_L g1545 ( 
.A1(n_1516),
.A2(n_1457),
.B1(n_1413),
.B2(n_1437),
.Y(n_1545)
);

AOI22xp33_ASAP7_75t_L g1546 ( 
.A1(n_1513),
.A2(n_1457),
.B1(n_1437),
.B2(n_1468),
.Y(n_1546)
);

NAND3xp33_ASAP7_75t_L g1547 ( 
.A(n_1515),
.B(n_1443),
.C(n_1475),
.Y(n_1547)
);

NOR3xp33_ASAP7_75t_L g1548 ( 
.A(n_1524),
.B(n_1480),
.C(n_1449),
.Y(n_1548)
);

AND2x2_ASAP7_75t_L g1549 ( 
.A(n_1499),
.B(n_1431),
.Y(n_1549)
);

NOR2xp33_ASAP7_75t_L g1550 ( 
.A(n_1521),
.B(n_1425),
.Y(n_1550)
);

NAND3xp33_ASAP7_75t_L g1551 ( 
.A(n_1515),
.B(n_1510),
.C(n_1498),
.Y(n_1551)
);

NAND3xp33_ASAP7_75t_L g1552 ( 
.A(n_1510),
.B(n_1443),
.C(n_1479),
.Y(n_1552)
);

NAND2xp5_ASAP7_75t_L g1553 ( 
.A(n_1500),
.B(n_1427),
.Y(n_1553)
);

OAI22xp5_ASAP7_75t_L g1554 ( 
.A1(n_1529),
.A2(n_1477),
.B1(n_1425),
.B2(n_1471),
.Y(n_1554)
);

NAND3xp33_ASAP7_75t_L g1555 ( 
.A(n_1501),
.B(n_1482),
.C(n_1474),
.Y(n_1555)
);

OAI221xp5_ASAP7_75t_SL g1556 ( 
.A1(n_1525),
.A2(n_1436),
.B1(n_1422),
.B2(n_1471),
.C(n_1477),
.Y(n_1556)
);

OAI21xp33_ASAP7_75t_L g1557 ( 
.A1(n_1501),
.A2(n_1436),
.B(n_1468),
.Y(n_1557)
);

AOI22xp33_ASAP7_75t_L g1558 ( 
.A1(n_1504),
.A2(n_1437),
.B1(n_1472),
.B2(n_1469),
.Y(n_1558)
);

NAND2xp5_ASAP7_75t_L g1559 ( 
.A(n_1484),
.B(n_1487),
.Y(n_1559)
);

OAI21xp5_ASAP7_75t_SL g1560 ( 
.A1(n_1492),
.A2(n_1469),
.B(n_1472),
.Y(n_1560)
);

NAND2xp5_ASAP7_75t_L g1561 ( 
.A(n_1484),
.B(n_1430),
.Y(n_1561)
);

AOI22xp33_ASAP7_75t_L g1562 ( 
.A1(n_1505),
.A2(n_1437),
.B1(n_1476),
.B2(n_1443),
.Y(n_1562)
);

NAND3xp33_ASAP7_75t_L g1563 ( 
.A(n_1493),
.B(n_1443),
.C(n_1479),
.Y(n_1563)
);

OAI22xp5_ASAP7_75t_L g1564 ( 
.A1(n_1503),
.A2(n_1466),
.B1(n_1418),
.B2(n_1438),
.Y(n_1564)
);

NAND2xp5_ASAP7_75t_L g1565 ( 
.A(n_1487),
.B(n_1488),
.Y(n_1565)
);

OAI21xp5_ASAP7_75t_SL g1566 ( 
.A1(n_1483),
.A2(n_1494),
.B(n_1511),
.Y(n_1566)
);

INVx1_ASAP7_75t_L g1567 ( 
.A(n_1519),
.Y(n_1567)
);

AND2x2_ASAP7_75t_L g1568 ( 
.A(n_1499),
.B(n_1448),
.Y(n_1568)
);

AND2x2_ASAP7_75t_L g1569 ( 
.A(n_1506),
.B(n_1448),
.Y(n_1569)
);

OAI21xp33_ASAP7_75t_L g1570 ( 
.A1(n_1525),
.A2(n_1451),
.B(n_1478),
.Y(n_1570)
);

NAND4xp25_ASAP7_75t_L g1571 ( 
.A(n_1493),
.B(n_1462),
.C(n_1460),
.D(n_1463),
.Y(n_1571)
);

OAI22xp5_ASAP7_75t_L g1572 ( 
.A1(n_1495),
.A2(n_1418),
.B1(n_1438),
.B2(n_1424),
.Y(n_1572)
);

NAND3xp33_ASAP7_75t_L g1573 ( 
.A(n_1525),
.B(n_1473),
.C(n_1475),
.Y(n_1573)
);

AND2x2_ASAP7_75t_L g1574 ( 
.A(n_1534),
.B(n_1528),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_1544),
.Y(n_1575)
);

NAND2xp5_ASAP7_75t_L g1576 ( 
.A(n_1531),
.B(n_1533),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_1544),
.Y(n_1577)
);

AND2x2_ASAP7_75t_L g1578 ( 
.A(n_1534),
.B(n_1528),
.Y(n_1578)
);

INVx1_ASAP7_75t_L g1579 ( 
.A(n_1567),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_1536),
.Y(n_1580)
);

AND2x2_ASAP7_75t_L g1581 ( 
.A(n_1568),
.B(n_1509),
.Y(n_1581)
);

OR2x2_ASAP7_75t_L g1582 ( 
.A(n_1551),
.B(n_1485),
.Y(n_1582)
);

AND2x2_ASAP7_75t_L g1583 ( 
.A(n_1569),
.B(n_1538),
.Y(n_1583)
);

AND2x2_ASAP7_75t_L g1584 ( 
.A(n_1538),
.B(n_1489),
.Y(n_1584)
);

NAND2xp5_ASAP7_75t_L g1585 ( 
.A(n_1553),
.B(n_1555),
.Y(n_1585)
);

OR2x2_ASAP7_75t_L g1586 ( 
.A(n_1547),
.B(n_1520),
.Y(n_1586)
);

NAND2xp5_ASAP7_75t_L g1587 ( 
.A(n_1555),
.B(n_1522),
.Y(n_1587)
);

AND2x2_ASAP7_75t_L g1588 ( 
.A(n_1549),
.B(n_1489),
.Y(n_1588)
);

BUFx2_ASAP7_75t_L g1589 ( 
.A(n_1530),
.Y(n_1589)
);

INVx3_ASAP7_75t_L g1590 ( 
.A(n_1549),
.Y(n_1590)
);

OR2x2_ASAP7_75t_L g1591 ( 
.A(n_1540),
.B(n_1526),
.Y(n_1591)
);

OR2x2_ASAP7_75t_L g1592 ( 
.A(n_1552),
.B(n_1490),
.Y(n_1592)
);

INVxp67_ASAP7_75t_L g1593 ( 
.A(n_1573),
.Y(n_1593)
);

INVx3_ASAP7_75t_L g1594 ( 
.A(n_1561),
.Y(n_1594)
);

INVx1_ASAP7_75t_L g1595 ( 
.A(n_1543),
.Y(n_1595)
);

AND2x2_ASAP7_75t_L g1596 ( 
.A(n_1562),
.B(n_1491),
.Y(n_1596)
);

HB1xp67_ASAP7_75t_L g1597 ( 
.A(n_1541),
.Y(n_1597)
);

AND2x4_ASAP7_75t_L g1598 ( 
.A(n_1548),
.B(n_1497),
.Y(n_1598)
);

AND2x2_ASAP7_75t_L g1599 ( 
.A(n_1590),
.B(n_1566),
.Y(n_1599)
);

OAI21xp33_ASAP7_75t_L g1600 ( 
.A1(n_1593),
.A2(n_1532),
.B(n_1537),
.Y(n_1600)
);

OR2x2_ASAP7_75t_L g1601 ( 
.A(n_1592),
.B(n_1563),
.Y(n_1601)
);

INVx1_ASAP7_75t_L g1602 ( 
.A(n_1575),
.Y(n_1602)
);

OR2x2_ASAP7_75t_L g1603 ( 
.A(n_1592),
.B(n_1571),
.Y(n_1603)
);

INVxp67_ASAP7_75t_L g1604 ( 
.A(n_1585),
.Y(n_1604)
);

INVx1_ASAP7_75t_L g1605 ( 
.A(n_1575),
.Y(n_1605)
);

INVx1_ASAP7_75t_L g1606 ( 
.A(n_1577),
.Y(n_1606)
);

AND2x4_ASAP7_75t_L g1607 ( 
.A(n_1590),
.B(n_1497),
.Y(n_1607)
);

INVx2_ASAP7_75t_L g1608 ( 
.A(n_1586),
.Y(n_1608)
);

INVx2_ASAP7_75t_L g1609 ( 
.A(n_1586),
.Y(n_1609)
);

AND2x2_ASAP7_75t_L g1610 ( 
.A(n_1590),
.B(n_1558),
.Y(n_1610)
);

NOR2xp33_ASAP7_75t_L g1611 ( 
.A(n_1585),
.B(n_1560),
.Y(n_1611)
);

NAND2xp5_ASAP7_75t_L g1612 ( 
.A(n_1593),
.B(n_1557),
.Y(n_1612)
);

NAND2xp5_ASAP7_75t_L g1613 ( 
.A(n_1576),
.B(n_1559),
.Y(n_1613)
);

INVx1_ASAP7_75t_L g1614 ( 
.A(n_1579),
.Y(n_1614)
);

AND2x2_ASAP7_75t_L g1615 ( 
.A(n_1583),
.B(n_1565),
.Y(n_1615)
);

AND2x2_ASAP7_75t_L g1616 ( 
.A(n_1583),
.B(n_1584),
.Y(n_1616)
);

AND2x2_ASAP7_75t_L g1617 ( 
.A(n_1583),
.B(n_1486),
.Y(n_1617)
);

HB1xp67_ASAP7_75t_L g1618 ( 
.A(n_1586),
.Y(n_1618)
);

INVx1_ASAP7_75t_L g1619 ( 
.A(n_1579),
.Y(n_1619)
);

HB1xp67_ASAP7_75t_L g1620 ( 
.A(n_1587),
.Y(n_1620)
);

INVx4_ASAP7_75t_L g1621 ( 
.A(n_1598),
.Y(n_1621)
);

INVxp67_ASAP7_75t_SL g1622 ( 
.A(n_1587),
.Y(n_1622)
);

O2A1O1Ixp33_ASAP7_75t_L g1623 ( 
.A1(n_1582),
.A2(n_1537),
.B(n_1556),
.C(n_1554),
.Y(n_1623)
);

INVx1_ASAP7_75t_L g1624 ( 
.A(n_1591),
.Y(n_1624)
);

INVx2_ASAP7_75t_L g1625 ( 
.A(n_1588),
.Y(n_1625)
);

AOI22xp5_ASAP7_75t_L g1626 ( 
.A1(n_1600),
.A2(n_1570),
.B1(n_1542),
.B2(n_1598),
.Y(n_1626)
);

AND2x2_ASAP7_75t_L g1627 ( 
.A(n_1616),
.B(n_1574),
.Y(n_1627)
);

INVx1_ASAP7_75t_L g1628 ( 
.A(n_1602),
.Y(n_1628)
);

NAND2xp5_ASAP7_75t_L g1629 ( 
.A(n_1600),
.B(n_1597),
.Y(n_1629)
);

OR2x2_ASAP7_75t_L g1630 ( 
.A(n_1603),
.B(n_1582),
.Y(n_1630)
);

INVx2_ASAP7_75t_L g1631 ( 
.A(n_1625),
.Y(n_1631)
);

OR2x2_ASAP7_75t_L g1632 ( 
.A(n_1603),
.B(n_1591),
.Y(n_1632)
);

NAND2xp5_ASAP7_75t_L g1633 ( 
.A(n_1604),
.B(n_1597),
.Y(n_1633)
);

A2O1A1Ixp33_ASAP7_75t_L g1634 ( 
.A1(n_1623),
.A2(n_1570),
.B(n_1598),
.C(n_1596),
.Y(n_1634)
);

INVx1_ASAP7_75t_L g1635 ( 
.A(n_1605),
.Y(n_1635)
);

AND2x2_ASAP7_75t_L g1636 ( 
.A(n_1616),
.B(n_1574),
.Y(n_1636)
);

NAND2xp5_ASAP7_75t_L g1637 ( 
.A(n_1604),
.B(n_1595),
.Y(n_1637)
);

INVx2_ASAP7_75t_SL g1638 ( 
.A(n_1621),
.Y(n_1638)
);

NOR3xp33_ASAP7_75t_L g1639 ( 
.A(n_1623),
.B(n_1611),
.C(n_1612),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_1606),
.Y(n_1640)
);

NAND2xp5_ASAP7_75t_L g1641 ( 
.A(n_1611),
.B(n_1595),
.Y(n_1641)
);

AND2x2_ASAP7_75t_L g1642 ( 
.A(n_1616),
.B(n_1574),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1606),
.Y(n_1643)
);

NAND2xp5_ASAP7_75t_L g1644 ( 
.A(n_1612),
.B(n_1594),
.Y(n_1644)
);

AND2x4_ASAP7_75t_L g1645 ( 
.A(n_1621),
.B(n_1598),
.Y(n_1645)
);

NAND2xp5_ASAP7_75t_L g1646 ( 
.A(n_1613),
.B(n_1594),
.Y(n_1646)
);

AOI31xp33_ASAP7_75t_L g1647 ( 
.A1(n_1603),
.A2(n_1564),
.A3(n_1598),
.B(n_1539),
.Y(n_1647)
);

AND2x2_ASAP7_75t_L g1648 ( 
.A(n_1599),
.B(n_1578),
.Y(n_1648)
);

INVx2_ASAP7_75t_L g1649 ( 
.A(n_1625),
.Y(n_1649)
);

NAND2xp5_ASAP7_75t_L g1650 ( 
.A(n_1613),
.B(n_1594),
.Y(n_1650)
);

AND2x2_ASAP7_75t_L g1651 ( 
.A(n_1599),
.B(n_1578),
.Y(n_1651)
);

NAND2x1_ASAP7_75t_L g1652 ( 
.A(n_1621),
.B(n_1589),
.Y(n_1652)
);

AND2x2_ASAP7_75t_L g1653 ( 
.A(n_1599),
.B(n_1578),
.Y(n_1653)
);

INVx1_ASAP7_75t_L g1654 ( 
.A(n_1614),
.Y(n_1654)
);

AND2x2_ASAP7_75t_L g1655 ( 
.A(n_1621),
.B(n_1581),
.Y(n_1655)
);

INVxp33_ASAP7_75t_L g1656 ( 
.A(n_1615),
.Y(n_1656)
);

AND2x4_ASAP7_75t_L g1657 ( 
.A(n_1621),
.B(n_1580),
.Y(n_1657)
);

NOR2xp33_ASAP7_75t_SL g1658 ( 
.A(n_1601),
.B(n_1572),
.Y(n_1658)
);

INVx1_ASAP7_75t_L g1659 ( 
.A(n_1619),
.Y(n_1659)
);

INVx2_ASAP7_75t_L g1660 ( 
.A(n_1625),
.Y(n_1660)
);

AND2x2_ASAP7_75t_L g1661 ( 
.A(n_1610),
.B(n_1581),
.Y(n_1661)
);

AND2x4_ASAP7_75t_L g1662 ( 
.A(n_1607),
.B(n_1580),
.Y(n_1662)
);

INVx2_ASAP7_75t_L g1663 ( 
.A(n_1631),
.Y(n_1663)
);

INVx4_ASAP7_75t_L g1664 ( 
.A(n_1645),
.Y(n_1664)
);

OR2x2_ASAP7_75t_L g1665 ( 
.A(n_1632),
.B(n_1601),
.Y(n_1665)
);

INVx1_ASAP7_75t_L g1666 ( 
.A(n_1628),
.Y(n_1666)
);

INVx2_ASAP7_75t_L g1667 ( 
.A(n_1649),
.Y(n_1667)
);

INVxp67_ASAP7_75t_L g1668 ( 
.A(n_1629),
.Y(n_1668)
);

AOI21xp5_ASAP7_75t_L g1669 ( 
.A1(n_1634),
.A2(n_1622),
.B(n_1601),
.Y(n_1669)
);

NAND2x1_ASAP7_75t_SL g1670 ( 
.A(n_1626),
.B(n_1618),
.Y(n_1670)
);

INVx2_ASAP7_75t_L g1671 ( 
.A(n_1649),
.Y(n_1671)
);

INVx1_ASAP7_75t_L g1672 ( 
.A(n_1628),
.Y(n_1672)
);

HB1xp67_ASAP7_75t_L g1673 ( 
.A(n_1635),
.Y(n_1673)
);

NAND2xp5_ASAP7_75t_L g1674 ( 
.A(n_1639),
.B(n_1641),
.Y(n_1674)
);

AND2x2_ASAP7_75t_L g1675 ( 
.A(n_1648),
.B(n_1622),
.Y(n_1675)
);

AND2x2_ASAP7_75t_L g1676 ( 
.A(n_1648),
.B(n_1618),
.Y(n_1676)
);

INVx1_ASAP7_75t_L g1677 ( 
.A(n_1635),
.Y(n_1677)
);

NAND2xp5_ASAP7_75t_L g1678 ( 
.A(n_1637),
.B(n_1620),
.Y(n_1678)
);

BUFx3_ASAP7_75t_L g1679 ( 
.A(n_1652),
.Y(n_1679)
);

AND2x2_ASAP7_75t_L g1680 ( 
.A(n_1651),
.B(n_1617),
.Y(n_1680)
);

INVx1_ASAP7_75t_L g1681 ( 
.A(n_1640),
.Y(n_1681)
);

INVx2_ASAP7_75t_L g1682 ( 
.A(n_1660),
.Y(n_1682)
);

OR2x2_ASAP7_75t_L g1683 ( 
.A(n_1632),
.B(n_1620),
.Y(n_1683)
);

HB1xp67_ASAP7_75t_L g1684 ( 
.A(n_1640),
.Y(n_1684)
);

HB1xp67_ASAP7_75t_L g1685 ( 
.A(n_1643),
.Y(n_1685)
);

OAI22xp33_ASAP7_75t_L g1686 ( 
.A1(n_1647),
.A2(n_1609),
.B1(n_1610),
.B2(n_1608),
.Y(n_1686)
);

INVx1_ASAP7_75t_L g1687 ( 
.A(n_1643),
.Y(n_1687)
);

INVx3_ASAP7_75t_L g1688 ( 
.A(n_1652),
.Y(n_1688)
);

AND2x2_ASAP7_75t_L g1689 ( 
.A(n_1653),
.B(n_1655),
.Y(n_1689)
);

BUFx3_ASAP7_75t_L g1690 ( 
.A(n_1638),
.Y(n_1690)
);

INVx2_ASAP7_75t_L g1691 ( 
.A(n_1660),
.Y(n_1691)
);

INVx1_ASAP7_75t_L g1692 ( 
.A(n_1654),
.Y(n_1692)
);

INVxp67_ASAP7_75t_L g1693 ( 
.A(n_1658),
.Y(n_1693)
);

AOI22xp33_ASAP7_75t_L g1694 ( 
.A1(n_1656),
.A2(n_1535),
.B1(n_1545),
.B2(n_1546),
.Y(n_1694)
);

INVx1_ASAP7_75t_SL g1695 ( 
.A(n_1638),
.Y(n_1695)
);

INVx1_ASAP7_75t_L g1696 ( 
.A(n_1654),
.Y(n_1696)
);

INVxp67_ASAP7_75t_L g1697 ( 
.A(n_1693),
.Y(n_1697)
);

NAND2xp5_ASAP7_75t_L g1698 ( 
.A(n_1674),
.B(n_1661),
.Y(n_1698)
);

AND2x2_ASAP7_75t_L g1699 ( 
.A(n_1689),
.B(n_1661),
.Y(n_1699)
);

OAI22xp5_ASAP7_75t_L g1700 ( 
.A1(n_1686),
.A2(n_1630),
.B1(n_1653),
.B2(n_1644),
.Y(n_1700)
);

INVx2_ASAP7_75t_L g1701 ( 
.A(n_1690),
.Y(n_1701)
);

INVx1_ASAP7_75t_L g1702 ( 
.A(n_1673),
.Y(n_1702)
);

AOI21xp33_ASAP7_75t_L g1703 ( 
.A1(n_1686),
.A2(n_1630),
.B(n_1633),
.Y(n_1703)
);

AND2x2_ASAP7_75t_L g1704 ( 
.A(n_1689),
.B(n_1627),
.Y(n_1704)
);

INVx1_ASAP7_75t_L g1705 ( 
.A(n_1673),
.Y(n_1705)
);

INVx1_ASAP7_75t_SL g1706 ( 
.A(n_1670),
.Y(n_1706)
);

INVx1_ASAP7_75t_L g1707 ( 
.A(n_1684),
.Y(n_1707)
);

INVx2_ASAP7_75t_L g1708 ( 
.A(n_1690),
.Y(n_1708)
);

NAND2xp33_ASAP7_75t_L g1709 ( 
.A(n_1674),
.B(n_1610),
.Y(n_1709)
);

NAND2xp5_ASAP7_75t_L g1710 ( 
.A(n_1668),
.B(n_1627),
.Y(n_1710)
);

AND2x2_ASAP7_75t_L g1711 ( 
.A(n_1689),
.B(n_1636),
.Y(n_1711)
);

INVx2_ASAP7_75t_L g1712 ( 
.A(n_1690),
.Y(n_1712)
);

AND2x2_ASAP7_75t_L g1713 ( 
.A(n_1664),
.B(n_1636),
.Y(n_1713)
);

OAI221xp5_ASAP7_75t_L g1714 ( 
.A1(n_1670),
.A2(n_1646),
.B1(n_1650),
.B2(n_1655),
.C(n_1608),
.Y(n_1714)
);

INVx1_ASAP7_75t_L g1715 ( 
.A(n_1684),
.Y(n_1715)
);

INVx1_ASAP7_75t_L g1716 ( 
.A(n_1685),
.Y(n_1716)
);

NAND5xp2_ASAP7_75t_L g1717 ( 
.A(n_1669),
.B(n_1550),
.C(n_1642),
.D(n_1615),
.E(n_1659),
.Y(n_1717)
);

NAND2xp5_ASAP7_75t_L g1718 ( 
.A(n_1668),
.B(n_1642),
.Y(n_1718)
);

AOI22xp5_ASAP7_75t_L g1719 ( 
.A1(n_1693),
.A2(n_1645),
.B1(n_1662),
.B2(n_1607),
.Y(n_1719)
);

AOI221xp5_ASAP7_75t_L g1720 ( 
.A1(n_1669),
.A2(n_1609),
.B1(n_1608),
.B2(n_1657),
.C(n_1645),
.Y(n_1720)
);

NOR2xp33_ASAP7_75t_L g1721 ( 
.A(n_1664),
.B(n_1401),
.Y(n_1721)
);

INVx1_ASAP7_75t_L g1722 ( 
.A(n_1685),
.Y(n_1722)
);

NAND2xp5_ASAP7_75t_L g1723 ( 
.A(n_1676),
.B(n_1615),
.Y(n_1723)
);

NAND2xp5_ASAP7_75t_L g1724 ( 
.A(n_1676),
.B(n_1624),
.Y(n_1724)
);

INVx1_ASAP7_75t_L g1725 ( 
.A(n_1666),
.Y(n_1725)
);

INVx1_ASAP7_75t_L g1726 ( 
.A(n_1702),
.Y(n_1726)
);

INVx1_ASAP7_75t_L g1727 ( 
.A(n_1702),
.Y(n_1727)
);

AND2x2_ASAP7_75t_L g1728 ( 
.A(n_1699),
.B(n_1664),
.Y(n_1728)
);

AND2x2_ASAP7_75t_L g1729 ( 
.A(n_1699),
.B(n_1664),
.Y(n_1729)
);

INVx1_ASAP7_75t_L g1730 ( 
.A(n_1716),
.Y(n_1730)
);

OR2x2_ASAP7_75t_L g1731 ( 
.A(n_1723),
.B(n_1698),
.Y(n_1731)
);

NOR2xp33_ASAP7_75t_L g1732 ( 
.A(n_1697),
.B(n_1664),
.Y(n_1732)
);

INVx1_ASAP7_75t_L g1733 ( 
.A(n_1716),
.Y(n_1733)
);

INVx1_ASAP7_75t_SL g1734 ( 
.A(n_1706),
.Y(n_1734)
);

NAND2xp5_ASAP7_75t_L g1735 ( 
.A(n_1709),
.B(n_1676),
.Y(n_1735)
);

AND2x2_ASAP7_75t_L g1736 ( 
.A(n_1713),
.B(n_1704),
.Y(n_1736)
);

INVx1_ASAP7_75t_L g1737 ( 
.A(n_1705),
.Y(n_1737)
);

INVx1_ASAP7_75t_L g1738 ( 
.A(n_1725),
.Y(n_1738)
);

INVx1_ASAP7_75t_SL g1739 ( 
.A(n_1709),
.Y(n_1739)
);

AND2x2_ASAP7_75t_L g1740 ( 
.A(n_1713),
.B(n_1675),
.Y(n_1740)
);

OAI21xp5_ASAP7_75t_SL g1741 ( 
.A1(n_1700),
.A2(n_1694),
.B(n_1675),
.Y(n_1741)
);

INVx2_ASAP7_75t_SL g1742 ( 
.A(n_1701),
.Y(n_1742)
);

AND2x2_ASAP7_75t_L g1743 ( 
.A(n_1704),
.B(n_1675),
.Y(n_1743)
);

NAND2xp5_ASAP7_75t_L g1744 ( 
.A(n_1701),
.B(n_1708),
.Y(n_1744)
);

NAND2xp5_ASAP7_75t_L g1745 ( 
.A(n_1708),
.B(n_1695),
.Y(n_1745)
);

AND2x2_ASAP7_75t_L g1746 ( 
.A(n_1711),
.B(n_1695),
.Y(n_1746)
);

NAND3xp33_ASAP7_75t_L g1747 ( 
.A(n_1741),
.B(n_1720),
.C(n_1703),
.Y(n_1747)
);

NAND2xp5_ASAP7_75t_L g1748 ( 
.A(n_1734),
.B(n_1712),
.Y(n_1748)
);

OAI21xp33_ASAP7_75t_L g1749 ( 
.A1(n_1732),
.A2(n_1717),
.B(n_1710),
.Y(n_1749)
);

NAND2xp5_ASAP7_75t_L g1750 ( 
.A(n_1739),
.B(n_1712),
.Y(n_1750)
);

AND2x2_ASAP7_75t_L g1751 ( 
.A(n_1736),
.B(n_1746),
.Y(n_1751)
);

NOR2xp33_ASAP7_75t_L g1752 ( 
.A(n_1731),
.B(n_1721),
.Y(n_1752)
);

NAND2xp5_ASAP7_75t_L g1753 ( 
.A(n_1746),
.B(n_1707),
.Y(n_1753)
);

AOI21xp5_ASAP7_75t_L g1754 ( 
.A1(n_1735),
.A2(n_1714),
.B(n_1718),
.Y(n_1754)
);

NOR3xp33_ASAP7_75t_L g1755 ( 
.A(n_1745),
.B(n_1722),
.C(n_1715),
.Y(n_1755)
);

O2A1O1Ixp33_ASAP7_75t_L g1756 ( 
.A1(n_1737),
.A2(n_1725),
.B(n_1678),
.C(n_1665),
.Y(n_1756)
);

OR2x2_ASAP7_75t_L g1757 ( 
.A(n_1731),
.B(n_1724),
.Y(n_1757)
);

NAND3xp33_ASAP7_75t_L g1758 ( 
.A(n_1744),
.B(n_1719),
.C(n_1665),
.Y(n_1758)
);

AOI21xp33_ASAP7_75t_SL g1759 ( 
.A1(n_1742),
.A2(n_1665),
.B(n_1683),
.Y(n_1759)
);

NAND4xp75_ASAP7_75t_L g1760 ( 
.A(n_1748),
.B(n_1742),
.C(n_1727),
.D(n_1726),
.Y(n_1760)
);

AOI22xp5_ASAP7_75t_L g1761 ( 
.A1(n_1747),
.A2(n_1736),
.B1(n_1740),
.B2(n_1743),
.Y(n_1761)
);

AOI211xp5_ASAP7_75t_L g1762 ( 
.A1(n_1759),
.A2(n_1737),
.B(n_1733),
.C(n_1730),
.Y(n_1762)
);

INVx1_ASAP7_75t_L g1763 ( 
.A(n_1751),
.Y(n_1763)
);

AND2x4_ASAP7_75t_L g1764 ( 
.A(n_1750),
.B(n_1728),
.Y(n_1764)
);

OAI211xp5_ASAP7_75t_SL g1765 ( 
.A1(n_1749),
.A2(n_1727),
.B(n_1726),
.C(n_1738),
.Y(n_1765)
);

AND2x2_ASAP7_75t_L g1766 ( 
.A(n_1752),
.B(n_1740),
.Y(n_1766)
);

NAND3xp33_ASAP7_75t_L g1767 ( 
.A(n_1755),
.B(n_1729),
.C(n_1728),
.Y(n_1767)
);

NOR2xp33_ASAP7_75t_L g1768 ( 
.A(n_1753),
.B(n_1729),
.Y(n_1768)
);

AND4x1_ASAP7_75t_L g1769 ( 
.A(n_1758),
.B(n_1743),
.C(n_1694),
.D(n_1711),
.Y(n_1769)
);

NOR4xp25_ASAP7_75t_L g1770 ( 
.A(n_1756),
.B(n_1696),
.C(n_1666),
.D(n_1677),
.Y(n_1770)
);

NAND2xp5_ASAP7_75t_L g1771 ( 
.A(n_1764),
.B(n_1754),
.Y(n_1771)
);

AND2x2_ASAP7_75t_L g1772 ( 
.A(n_1766),
.B(n_1757),
.Y(n_1772)
);

AND2x2_ASAP7_75t_L g1773 ( 
.A(n_1763),
.B(n_1680),
.Y(n_1773)
);

NOR3xp33_ASAP7_75t_L g1774 ( 
.A(n_1765),
.B(n_1333),
.C(n_1688),
.Y(n_1774)
);

AOI221xp5_ASAP7_75t_L g1775 ( 
.A1(n_1770),
.A2(n_1678),
.B1(n_1679),
.B2(n_1690),
.C(n_1696),
.Y(n_1775)
);

AND2x2_ASAP7_75t_L g1776 ( 
.A(n_1764),
.B(n_1680),
.Y(n_1776)
);

INVx1_ASAP7_75t_L g1777 ( 
.A(n_1776),
.Y(n_1777)
);

AOI22xp5_ASAP7_75t_L g1778 ( 
.A1(n_1774),
.A2(n_1768),
.B1(n_1761),
.B2(n_1767),
.Y(n_1778)
);

AND2x2_ASAP7_75t_L g1779 ( 
.A(n_1773),
.B(n_1772),
.Y(n_1779)
);

NAND3xp33_ASAP7_75t_L g1780 ( 
.A(n_1771),
.B(n_1769),
.C(n_1762),
.Y(n_1780)
);

NAND2xp5_ASAP7_75t_L g1781 ( 
.A(n_1775),
.B(n_1760),
.Y(n_1781)
);

INVx1_ASAP7_75t_L g1782 ( 
.A(n_1776),
.Y(n_1782)
);

INVx1_ASAP7_75t_L g1783 ( 
.A(n_1776),
.Y(n_1783)
);

NOR3xp33_ASAP7_75t_L g1784 ( 
.A(n_1780),
.B(n_1688),
.C(n_1343),
.Y(n_1784)
);

NOR2x1_ASAP7_75t_L g1785 ( 
.A(n_1779),
.B(n_1679),
.Y(n_1785)
);

AND2x4_ASAP7_75t_L g1786 ( 
.A(n_1777),
.B(n_1679),
.Y(n_1786)
);

NAND4xp25_ASAP7_75t_L g1787 ( 
.A(n_1778),
.B(n_1781),
.C(n_1783),
.D(n_1782),
.Y(n_1787)
);

OAI22xp33_ASAP7_75t_L g1788 ( 
.A1(n_1781),
.A2(n_1679),
.B1(n_1688),
.B2(n_1683),
.Y(n_1788)
);

NAND2xp5_ASAP7_75t_L g1789 ( 
.A(n_1779),
.B(n_1683),
.Y(n_1789)
);

NOR3xp33_ASAP7_75t_L g1790 ( 
.A(n_1787),
.B(n_1343),
.C(n_1688),
.Y(n_1790)
);

OAI21xp5_ASAP7_75t_L g1791 ( 
.A1(n_1785),
.A2(n_1688),
.B(n_1677),
.Y(n_1791)
);

INVx1_ASAP7_75t_L g1792 ( 
.A(n_1789),
.Y(n_1792)
);

INVx1_ASAP7_75t_L g1793 ( 
.A(n_1786),
.Y(n_1793)
);

NOR2xp33_ASAP7_75t_L g1794 ( 
.A(n_1793),
.B(n_1788),
.Y(n_1794)
);

XNOR2xp5_ASAP7_75t_L g1795 ( 
.A(n_1790),
.B(n_1784),
.Y(n_1795)
);

NAND3xp33_ASAP7_75t_SL g1796 ( 
.A(n_1794),
.B(n_1792),
.C(n_1791),
.Y(n_1796)
);

XOR2xp5_ASAP7_75t_L g1797 ( 
.A(n_1796),
.B(n_1795),
.Y(n_1797)
);

INVx1_ASAP7_75t_L g1798 ( 
.A(n_1796),
.Y(n_1798)
);

OAI22xp5_ASAP7_75t_L g1799 ( 
.A1(n_1798),
.A2(n_1692),
.B1(n_1672),
.B2(n_1687),
.Y(n_1799)
);

AOI21xp5_ASAP7_75t_L g1800 ( 
.A1(n_1797),
.A2(n_1681),
.B(n_1672),
.Y(n_1800)
);

AOI21xp5_ASAP7_75t_L g1801 ( 
.A1(n_1800),
.A2(n_1687),
.B(n_1681),
.Y(n_1801)
);

INVx1_ASAP7_75t_L g1802 ( 
.A(n_1801),
.Y(n_1802)
);

HB1xp67_ASAP7_75t_L g1803 ( 
.A(n_1802),
.Y(n_1803)
);

AOI221xp5_ASAP7_75t_L g1804 ( 
.A1(n_1803),
.A2(n_1799),
.B1(n_1692),
.B2(n_1682),
.C(n_1691),
.Y(n_1804)
);

AOI211xp5_ASAP7_75t_L g1805 ( 
.A1(n_1804),
.A2(n_1663),
.B(n_1671),
.C(n_1667),
.Y(n_1805)
);


endmodule