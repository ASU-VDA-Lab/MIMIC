module fake_jpeg_15380_n_229 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_229);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_229;

wire n_159;
wire n_117;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_212;
wire n_131;
wire n_56;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g15 ( 
.A(n_9),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_14),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_14),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

INVx11_ASAP7_75t_SL g23 ( 
.A(n_14),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_5),
.Y(n_24)
);

BUFx2_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

BUFx10_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_6),
.B(n_9),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_10),
.B(n_12),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_17),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_31),
.Y(n_43)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_17),
.Y(n_32)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_32),
.Y(n_47)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_17),
.Y(n_33)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_33),
.Y(n_52)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

HB1xp67_ASAP7_75t_L g49 ( 
.A(n_34),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_27),
.B(n_7),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_35),
.B(n_40),
.Y(n_44)
);

AND2x2_ASAP7_75t_L g36 ( 
.A(n_27),
.B(n_0),
.Y(n_36)
);

AND2x2_ASAP7_75t_L g56 ( 
.A(n_36),
.B(n_0),
.Y(n_56)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_17),
.Y(n_37)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_37),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_22),
.Y(n_38)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_38),
.Y(n_41)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_22),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_39),
.B(n_22),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_27),
.B(n_7),
.Y(n_40)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_33),
.Y(n_45)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_45),
.Y(n_64)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_46),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_39),
.A2(n_23),
.B1(n_21),
.B2(n_24),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_L g80 ( 
.A1(n_48),
.A2(n_57),
.B1(n_19),
.B2(n_30),
.Y(n_80)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_31),
.Y(n_50)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_50),
.Y(n_70)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_31),
.Y(n_51)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_51),
.Y(n_79)
);

CKINVDCx14_ASAP7_75t_R g72 ( 
.A(n_53),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_36),
.A2(n_16),
.B1(n_21),
.B2(n_24),
.Y(n_54)
);

CKINVDCx16_ASAP7_75t_R g75 ( 
.A(n_54),
.Y(n_75)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_55),
.B(n_38),
.Y(n_58)
);

OR2x2_ASAP7_75t_SL g59 ( 
.A(n_56),
.B(n_36),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_35),
.A2(n_16),
.B1(n_20),
.B2(n_15),
.Y(n_57)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_58),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_59),
.B(n_1),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_56),
.B(n_36),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_60),
.B(n_44),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_55),
.A2(n_23),
.B1(n_20),
.B2(n_15),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_62),
.A2(n_69),
.B1(n_74),
.B2(n_30),
.Y(n_89)
);

BUFx4f_ASAP7_75t_L g63 ( 
.A(n_43),
.Y(n_63)
);

HB1xp67_ASAP7_75t_L g100 ( 
.A(n_63),
.Y(n_100)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_43),
.Y(n_65)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_65),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_43),
.Y(n_66)
);

INVx13_ASAP7_75t_L g84 ( 
.A(n_66),
.Y(n_84)
);

NOR2x1_ASAP7_75t_L g67 ( 
.A(n_54),
.B(n_40),
.Y(n_67)
);

OR2x2_ASAP7_75t_L g86 ( 
.A(n_67),
.B(n_34),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_49),
.B(n_29),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_68),
.B(n_77),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_41),
.A2(n_20),
.B1(n_32),
.B2(n_28),
.Y(n_69)
);

CKINVDCx12_ASAP7_75t_R g71 ( 
.A(n_42),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_71),
.B(n_73),
.Y(n_102)
);

INVx13_ASAP7_75t_L g73 ( 
.A(n_41),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_50),
.A2(n_32),
.B1(n_28),
.B2(n_19),
.Y(n_74)
);

INVx4_ASAP7_75t_SL g76 ( 
.A(n_47),
.Y(n_76)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_76),
.Y(n_87)
);

INVx1_ASAP7_75t_SL g77 ( 
.A(n_56),
.Y(n_77)
);

INVx6_ASAP7_75t_L g78 ( 
.A(n_51),
.Y(n_78)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_78),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_80),
.B(n_48),
.Y(n_91)
);

AO22x1_ASAP7_75t_SL g81 ( 
.A1(n_67),
.A2(n_46),
.B1(n_45),
.B2(n_42),
.Y(n_81)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_81),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_82),
.B(n_86),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_75),
.A2(n_47),
.B1(n_52),
.B2(n_44),
.Y(n_85)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_85),
.Y(n_111)
);

AND2x6_ASAP7_75t_L g88 ( 
.A(n_75),
.B(n_1),
.Y(n_88)
);

A2O1A1O1Ixp25_ASAP7_75t_L g117 ( 
.A1(n_88),
.A2(n_25),
.B(n_2),
.C(n_3),
.D(n_4),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_89),
.B(n_25),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_60),
.B(n_52),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_90),
.B(n_92),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_91),
.B(n_93),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_77),
.B(n_26),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_59),
.B(n_29),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_72),
.B(n_26),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_95),
.B(n_96),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_64),
.B(n_26),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_SL g108 ( 
.A1(n_99),
.A2(n_25),
.B(n_18),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_64),
.B(n_26),
.C(n_18),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_101),
.B(n_103),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_61),
.B(n_26),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_105),
.A2(n_87),
.B1(n_65),
.B2(n_78),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_SL g138 ( 
.A1(n_108),
.A2(n_117),
.B(n_121),
.Y(n_138)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_96),
.Y(n_112)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_112),
.Y(n_133)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_94),
.Y(n_113)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_113),
.Y(n_148)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_94),
.Y(n_114)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_114),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_83),
.B(n_61),
.Y(n_115)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_115),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_90),
.B(n_79),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_116),
.B(n_120),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_L g118 ( 
.A1(n_86),
.A2(n_76),
.B(n_25),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_L g132 ( 
.A1(n_118),
.A2(n_86),
.B(n_87),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_83),
.B(n_73),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_SL g121 ( 
.A1(n_92),
.A2(n_76),
.B(n_63),
.Y(n_121)
);

INVx2_ASAP7_75t_SL g122 ( 
.A(n_100),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_L g146 ( 
.A1(n_122),
.A2(n_63),
.B1(n_84),
.B2(n_70),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_95),
.B(n_18),
.Y(n_123)
);

CKINVDCx16_ASAP7_75t_R g134 ( 
.A(n_123),
.Y(n_134)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_98),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_124),
.Y(n_130)
);

BUFx2_ASAP7_75t_L g125 ( 
.A(n_98),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_125),
.Y(n_136)
);

XOR2x2_ASAP7_75t_L g126 ( 
.A(n_81),
.B(n_82),
.Y(n_126)
);

XOR2x2_ASAP7_75t_SL g127 ( 
.A(n_126),
.B(n_81),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_SL g166 ( 
.A(n_127),
.B(n_132),
.C(n_139),
.Y(n_166)
);

OAI32xp33_ASAP7_75t_L g128 ( 
.A1(n_126),
.A2(n_91),
.A3(n_97),
.B1(n_81),
.B2(n_89),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_SL g161 ( 
.A(n_128),
.B(n_129),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_L g129 ( 
.A(n_126),
.B(n_97),
.Y(n_129)
);

XOR2xp5_ASAP7_75t_L g131 ( 
.A(n_110),
.B(n_85),
.Y(n_131)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_131),
.B(n_142),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g137 ( 
.A(n_122),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_137),
.B(n_140),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_113),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_106),
.A2(n_99),
.B1(n_88),
.B2(n_103),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_141),
.A2(n_144),
.B1(n_117),
.B2(n_112),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g142 ( 
.A(n_104),
.B(n_101),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_106),
.A2(n_99),
.B1(n_79),
.B2(n_70),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_146),
.Y(n_151)
);

AOI21xp5_ASAP7_75t_L g147 ( 
.A1(n_121),
.A2(n_102),
.B(n_93),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_SL g158 ( 
.A1(n_147),
.A2(n_149),
.B(n_111),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_L g149 ( 
.A1(n_118),
.A2(n_111),
.B(n_119),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_133),
.B(n_109),
.Y(n_150)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_150),
.Y(n_171)
);

INVx13_ASAP7_75t_L g152 ( 
.A(n_137),
.Y(n_152)
);

CKINVDCx14_ASAP7_75t_R g169 ( 
.A(n_152),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_133),
.B(n_109),
.Y(n_153)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_153),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_SL g154 ( 
.A(n_143),
.B(n_107),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_SL g174 ( 
.A(n_154),
.B(n_155),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_134),
.B(n_107),
.Y(n_155)
);

BUFx12f_ASAP7_75t_SL g156 ( 
.A(n_127),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_156),
.A2(n_144),
.B1(n_141),
.B2(n_147),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_SL g176 ( 
.A(n_158),
.B(n_108),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_148),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_159),
.B(n_163),
.Y(n_182)
);

HB1xp67_ASAP7_75t_L g160 ( 
.A(n_135),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_160),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_SL g162 ( 
.A(n_145),
.B(n_116),
.Y(n_162)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_162),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_136),
.B(n_122),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_SL g164 ( 
.A1(n_138),
.A2(n_110),
.B(n_104),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_164),
.B(n_161),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_167),
.A2(n_168),
.B1(n_148),
.B2(n_138),
.Y(n_172)
);

AOI22x1_ASAP7_75t_L g168 ( 
.A1(n_128),
.A2(n_125),
.B1(n_114),
.B2(n_84),
.Y(n_168)
);

AOI21xp5_ASAP7_75t_L g189 ( 
.A1(n_170),
.A2(n_158),
.B(n_164),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_172),
.A2(n_173),
.B1(n_175),
.B2(n_178),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_168),
.A2(n_149),
.B1(n_132),
.B2(n_131),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_168),
.A2(n_129),
.B1(n_142),
.B2(n_130),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_176),
.B(n_180),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_156),
.A2(n_124),
.B1(n_84),
.B2(n_125),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g179 ( 
.A(n_151),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_179),
.B(n_152),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_171),
.A2(n_150),
.B1(n_153),
.B2(n_166),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_184),
.B(n_191),
.Y(n_204)
);

CKINVDCx14_ASAP7_75t_R g185 ( 
.A(n_182),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_185),
.B(n_188),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_174),
.B(n_157),
.Y(n_186)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_186),
.Y(n_202)
);

INVxp67_ASAP7_75t_L g188 ( 
.A(n_182),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_189),
.B(n_195),
.C(n_165),
.Y(n_198)
);

INVxp67_ASAP7_75t_L g191 ( 
.A(n_178),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_171),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_192),
.A2(n_193),
.B1(n_194),
.B2(n_159),
.Y(n_196)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_177),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_180),
.B(n_165),
.C(n_161),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_196),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_198),
.B(n_199),
.C(n_200),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_195),
.B(n_175),
.C(n_181),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_187),
.B(n_172),
.C(n_173),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_187),
.B(n_183),
.C(n_176),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_SL g206 ( 
.A(n_201),
.B(n_203),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_190),
.B(n_169),
.C(n_179),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_190),
.B(n_166),
.C(n_22),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_L g210 ( 
.A1(n_205),
.A2(n_191),
.B(n_151),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_197),
.B(n_188),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_208),
.B(n_66),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_210),
.B(n_1),
.Y(n_214)
);

XNOR2x1_ASAP7_75t_L g211 ( 
.A(n_204),
.B(n_197),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_211),
.B(n_212),
.Y(n_216)
);

AOI21xp5_ASAP7_75t_L g212 ( 
.A1(n_202),
.A2(n_184),
.B(n_2),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_213),
.Y(n_220)
);

AOI21xp5_ASAP7_75t_L g218 ( 
.A1(n_214),
.A2(n_6),
.B(n_8),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_209),
.A2(n_3),
.B1(n_4),
.B2(n_6),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_215),
.B(n_217),
.C(n_216),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_207),
.B(n_4),
.Y(n_217)
);

AOI322xp5_ASAP7_75t_L g223 ( 
.A1(n_218),
.A2(n_8),
.A3(n_10),
.B1(n_11),
.B2(n_12),
.C1(n_13),
.C2(n_66),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_219),
.B(n_221),
.C(n_217),
.Y(n_222)
);

AOI21xp5_ASAP7_75t_L g221 ( 
.A1(n_216),
.A2(n_206),
.B(n_208),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_222),
.B(n_224),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_SL g225 ( 
.A(n_223),
.B(n_11),
.Y(n_225)
);

AOI322xp5_ASAP7_75t_L g224 ( 
.A1(n_220),
.A2(n_8),
.A3(n_11),
.B1(n_12),
.B2(n_13),
.C1(n_26),
.C2(n_206),
.Y(n_224)
);

INVxp33_ASAP7_75t_SL g227 ( 
.A(n_225),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_227),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_228),
.B(n_226),
.Y(n_229)
);


endmodule