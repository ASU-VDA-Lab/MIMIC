module fake_jpeg_8804_n_204 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_204);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_204;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_155;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_5),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_7),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_12),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

INVx11_ASAP7_75t_SL g21 ( 
.A(n_0),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

BUFx10_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_12),
.B(n_5),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_10),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

INVx11_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_29),
.Y(n_42)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_24),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_30),
.B(n_31),
.Y(n_43)
);

INVx5_ASAP7_75t_L g31 ( 
.A(n_21),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_24),
.Y(n_32)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_32),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_23),
.Y(n_33)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_24),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_34),
.B(n_35),
.Y(n_52)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_24),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_26),
.B(n_0),
.Y(n_36)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

INVx11_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

INVx4_ASAP7_75t_SL g38 ( 
.A(n_14),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_38),
.A2(n_34),
.B1(n_35),
.B2(n_29),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_L g40 ( 
.A1(n_30),
.A2(n_15),
.B1(n_27),
.B2(n_22),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_40),
.A2(n_41),
.B1(n_46),
.B2(n_17),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_L g41 ( 
.A1(n_30),
.A2(n_15),
.B1(n_27),
.B2(n_22),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_L g46 ( 
.A1(n_34),
.A2(n_25),
.B1(n_17),
.B2(n_18),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_33),
.Y(n_47)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_47),
.Y(n_57)
);

INVxp67_ASAP7_75t_L g61 ( 
.A(n_48),
.Y(n_61)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_32),
.Y(n_50)
);

INVx3_ASAP7_75t_SL g65 ( 
.A(n_50),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_36),
.B(n_19),
.Y(n_51)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_51),
.B(n_18),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_53),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_33),
.Y(n_54)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_54),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_31),
.B(n_16),
.Y(n_55)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_55),
.Y(n_62)
);

CKINVDCx14_ASAP7_75t_R g56 ( 
.A(n_43),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_56),
.B(n_58),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_45),
.B(n_16),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_59),
.B(n_66),
.Y(n_78)
);

OAI21xp5_ASAP7_75t_SL g60 ( 
.A1(n_52),
.A2(n_19),
.B(n_25),
.Y(n_60)
);

AOI21xp5_ASAP7_75t_L g81 ( 
.A1(n_60),
.A2(n_50),
.B(n_29),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_63),
.A2(n_38),
.B1(n_37),
.B2(n_14),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_51),
.B(n_35),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_64),
.B(n_75),
.Y(n_96)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_42),
.Y(n_66)
);

NAND2xp33_ASAP7_75t_SL g67 ( 
.A(n_45),
.B(n_23),
.Y(n_67)
);

OAI21xp5_ASAP7_75t_SL g80 ( 
.A1(n_67),
.A2(n_68),
.B(n_73),
.Y(n_80)
);

AO21x1_ASAP7_75t_L g68 ( 
.A1(n_39),
.A2(n_26),
.B(n_38),
.Y(n_68)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_42),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_70),
.B(n_71),
.Y(n_85)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_47),
.Y(n_71)
);

INVx2_ASAP7_75t_SL g72 ( 
.A(n_54),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_72),
.B(n_76),
.Y(n_92)
);

AND2x4_ASAP7_75t_SL g73 ( 
.A(n_39),
.B(n_38),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_44),
.B(n_28),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_44),
.B(n_31),
.Y(n_76)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_65),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_77),
.B(n_79),
.Y(n_115)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_75),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_81),
.B(n_82),
.Y(n_116)
);

INVx1_ASAP7_75t_SL g82 ( 
.A(n_73),
.Y(n_82)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_72),
.Y(n_83)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_83),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_65),
.Y(n_86)
);

INVx1_ASAP7_75t_SL g106 ( 
.A(n_86),
.Y(n_106)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_65),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_87),
.B(n_91),
.Y(n_119)
);

A2O1A1Ixp33_ASAP7_75t_SL g118 ( 
.A1(n_88),
.A2(n_70),
.B(n_28),
.C(n_20),
.Y(n_118)
);

BUFx2_ASAP7_75t_L g89 ( 
.A(n_73),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_89),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_61),
.A2(n_37),
.B1(n_32),
.B2(n_42),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_90),
.A2(n_93),
.B1(n_95),
.B2(n_97),
.Y(n_109)
);

INVx1_ASAP7_75t_SL g91 ( 
.A(n_64),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_61),
.A2(n_32),
.B1(n_49),
.B2(n_53),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_72),
.B(n_21),
.Y(n_94)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_94),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_68),
.A2(n_53),
.B1(n_49),
.B2(n_33),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_66),
.A2(n_49),
.B1(n_28),
.B2(n_20),
.Y(n_97)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_71),
.Y(n_98)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_98),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_58),
.B(n_28),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_99),
.B(n_58),
.Y(n_102)
);

OAI32xp33_ASAP7_75t_L g100 ( 
.A1(n_96),
.A2(n_99),
.A3(n_89),
.B1(n_82),
.B2(n_80),
.Y(n_100)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_100),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_84),
.B(n_62),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_101),
.B(n_102),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_96),
.B(n_60),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_103),
.B(n_108),
.Y(n_123)
);

OR2x2_ASAP7_75t_L g104 ( 
.A(n_92),
.B(n_0),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_104),
.B(n_112),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_L g105 ( 
.A(n_80),
.B(n_89),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_105),
.B(n_110),
.C(n_23),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_91),
.B(n_62),
.Y(n_108)
);

XOR2xp5_ASAP7_75t_L g110 ( 
.A(n_81),
.B(n_23),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_78),
.B(n_11),
.Y(n_112)
);

NOR2x1_ASAP7_75t_L g113 ( 
.A(n_95),
.B(n_93),
.Y(n_113)
);

NOR2x1_ASAP7_75t_L g132 ( 
.A(n_113),
.B(n_90),
.Y(n_132)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_85),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_114),
.B(n_97),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_118),
.A2(n_87),
.B1(n_77),
.B2(n_86),
.Y(n_129)
);

XOR2xp5_ASAP7_75t_L g121 ( 
.A(n_105),
.B(n_79),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_121),
.B(n_138),
.C(n_109),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_103),
.B(n_98),
.Y(n_124)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_124),
.Y(n_154)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_115),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_126),
.B(n_127),
.Y(n_141)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_119),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_129),
.B(n_135),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_120),
.B(n_74),
.Y(n_130)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_130),
.Y(n_140)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_131),
.Y(n_149)
);

AND2x2_ASAP7_75t_L g142 ( 
.A(n_132),
.B(n_110),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_SL g133 ( 
.A1(n_116),
.A2(n_83),
.B(n_23),
.Y(n_133)
);

AOI21xp5_ASAP7_75t_L g155 ( 
.A1(n_133),
.A2(n_136),
.B(n_107),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_108),
.B(n_20),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g143 ( 
.A(n_134),
.B(n_114),
.Y(n_143)
);

BUFx3_ASAP7_75t_L g135 ( 
.A(n_111),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_SL g136 ( 
.A1(n_117),
.A2(n_23),
.B(n_57),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_113),
.A2(n_69),
.B1(n_74),
.B2(n_57),
.Y(n_137)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_137),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_109),
.A2(n_69),
.B1(n_20),
.B2(n_13),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_139),
.B(n_104),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_SL g162 ( 
.A1(n_142),
.A2(n_155),
.B(n_127),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_143),
.B(n_146),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g144 ( 
.A(n_121),
.B(n_102),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_144),
.B(n_148),
.C(n_150),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_123),
.B(n_111),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_126),
.B(n_106),
.Y(n_147)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_147),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_138),
.B(n_100),
.C(n_107),
.Y(n_150)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_151),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_123),
.B(n_124),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_153),
.B(n_122),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_150),
.B(n_125),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_156),
.B(n_142),
.C(n_118),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_149),
.B(n_140),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_159),
.B(n_163),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_152),
.A2(n_125),
.B1(n_132),
.B2(n_137),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_160),
.A2(n_164),
.B1(n_165),
.B2(n_145),
.Y(n_170)
);

AND2x2_ASAP7_75t_L g173 ( 
.A(n_162),
.B(n_1),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_154),
.A2(n_129),
.B1(n_139),
.B2(n_136),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_154),
.A2(n_106),
.B1(n_118),
.B2(n_133),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_SL g166 ( 
.A(n_141),
.B(n_128),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_166),
.B(n_1),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_158),
.B(n_151),
.Y(n_168)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_168),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_170),
.Y(n_185)
);

OAI322xp33_ASAP7_75t_L g171 ( 
.A1(n_163),
.A2(n_153),
.A3(n_155),
.B1(n_144),
.B2(n_142),
.C1(n_148),
.C2(n_118),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_L g179 ( 
.A1(n_171),
.A2(n_167),
.B(n_162),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_172),
.B(n_176),
.C(n_177),
.Y(n_183)
);

AND2x2_ASAP7_75t_L g182 ( 
.A(n_173),
.B(n_2),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_157),
.B(n_11),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_174),
.B(n_175),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_161),
.B(n_135),
.C(n_2),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_161),
.B(n_1),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_179),
.B(n_176),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_SL g180 ( 
.A(n_169),
.B(n_156),
.Y(n_180)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_180),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_172),
.B(n_160),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_181),
.B(n_182),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_185),
.A2(n_164),
.B1(n_165),
.B2(n_173),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_187),
.B(n_192),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_188),
.B(n_190),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_181),
.B(n_2),
.C(n_3),
.Y(n_190)
);

O2A1O1Ixp33_ASAP7_75t_SL g191 ( 
.A1(n_184),
.A2(n_3),
.B(n_4),
.C(n_5),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_SL g194 ( 
.A1(n_191),
.A2(n_6),
.B(n_7),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_183),
.A2(n_4),
.B1(n_6),
.B2(n_7),
.Y(n_192)
);

NAND3xp33_ASAP7_75t_SL g193 ( 
.A(n_186),
.B(n_182),
.C(n_178),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_193),
.B(n_196),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_194),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_SL g196 ( 
.A(n_189),
.B(n_8),
.Y(n_196)
);

INVxp67_ASAP7_75t_L g198 ( 
.A(n_197),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_L g203 ( 
.A1(n_198),
.A2(n_199),
.B(n_10),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_195),
.B(n_190),
.C(n_188),
.Y(n_199)
);

AOI22xp33_ASAP7_75t_SL g202 ( 
.A1(n_201),
.A2(n_10),
.B1(n_191),
.B2(n_200),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_202),
.B(n_203),
.Y(n_204)
);


endmodule