module fake_jpeg_22140_n_327 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_327);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_327;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx2_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_16),
.Y(n_18)
);

BUFx10_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

INVx13_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_3),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_16),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_4),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_11),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_1),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_2),
.Y(n_35)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_1),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_15),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_21),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_38),
.B(n_43),
.Y(n_69)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_20),
.Y(n_39)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_39),
.Y(n_65)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_21),
.Y(n_40)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_23),
.Y(n_41)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

INVx11_ASAP7_75t_L g42 ( 
.A(n_19),
.Y(n_42)
);

BUFx10_ASAP7_75t_L g55 ( 
.A(n_42),
.Y(n_55)
);

CKINVDCx16_ASAP7_75t_R g43 ( 
.A(n_20),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_21),
.Y(n_44)
);

INVx2_ASAP7_75t_SL g63 ( 
.A(n_44),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_21),
.Y(n_45)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_45),
.Y(n_73)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_24),
.Y(n_46)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_46),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_24),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_47),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_24),
.Y(n_48)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_48),
.Y(n_53)
);

INVx13_ASAP7_75t_L g49 ( 
.A(n_19),
.Y(n_49)
);

BUFx4f_ASAP7_75t_SL g60 ( 
.A(n_49),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_39),
.A2(n_28),
.B1(n_17),
.B2(n_35),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_50),
.A2(n_77),
.B1(n_38),
.B2(n_31),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_39),
.A2(n_28),
.B1(n_17),
.B2(n_35),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_51),
.A2(n_62),
.B1(n_64),
.B2(n_41),
.Y(n_94)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_42),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_56),
.B(n_57),
.Y(n_84)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_40),
.B(n_27),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_58),
.B(n_19),
.Y(n_83)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_46),
.Y(n_59)
);

INVx6_ASAP7_75t_L g107 ( 
.A(n_59),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_39),
.A2(n_23),
.B1(n_36),
.B2(n_24),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_42),
.A2(n_36),
.B1(n_37),
.B2(n_34),
.Y(n_64)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_42),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_66),
.B(n_67),
.Y(n_116)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_41),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_44),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_68),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_43),
.A2(n_18),
.B1(n_34),
.B2(n_37),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_70),
.A2(n_29),
.B1(n_25),
.B2(n_65),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_46),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_71),
.Y(n_91)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_46),
.Y(n_72)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_72),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_44),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_74),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_48),
.Y(n_76)
);

HB1xp67_ASAP7_75t_L g97 ( 
.A(n_76),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_43),
.A2(n_25),
.B1(n_27),
.B2(n_30),
.Y(n_77)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_48),
.Y(n_78)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_78),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_69),
.B(n_77),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_79),
.B(n_100),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_65),
.A2(n_18),
.B1(n_49),
.B2(n_30),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_82),
.A2(n_89),
.B1(n_103),
.B2(n_78),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_83),
.B(n_87),
.Y(n_131)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_75),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_85),
.B(n_88),
.Y(n_120)
);

BUFx12f_ASAP7_75t_L g86 ( 
.A(n_60),
.Y(n_86)
);

BUFx3_ASAP7_75t_L g145 ( 
.A(n_86),
.Y(n_145)
);

A2O1A1Ixp33_ASAP7_75t_L g87 ( 
.A1(n_50),
.A2(n_19),
.B(n_44),
.C(n_47),
.Y(n_87)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_60),
.Y(n_88)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_60),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_90),
.B(n_95),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_61),
.B(n_29),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_93),
.B(n_102),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_94),
.A2(n_109),
.B1(n_113),
.B2(n_22),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_55),
.Y(n_95)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_54),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_96),
.B(n_98),
.Y(n_138)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_54),
.Y(n_98)
);

CKINVDCx14_ASAP7_75t_R g99 ( 
.A(n_53),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_99),
.B(n_104),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_55),
.B(n_45),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_59),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_101),
.Y(n_150)
);

A2O1A1Ixp33_ASAP7_75t_L g102 ( 
.A1(n_55),
.A2(n_44),
.B(n_47),
.C(n_45),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_73),
.A2(n_49),
.B1(n_40),
.B2(n_44),
.Y(n_103)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_52),
.Y(n_104)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_52),
.Y(n_105)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_105),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_61),
.B(n_38),
.C(n_48),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_108),
.B(n_63),
.C(n_76),
.Y(n_121)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_56),
.B(n_49),
.Y(n_110)
);

AND2x2_ASAP7_75t_L g128 ( 
.A(n_110),
.B(n_0),
.Y(n_128)
);

INVx1_ASAP7_75t_SL g111 ( 
.A(n_55),
.Y(n_111)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_111),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_66),
.Y(n_112)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_112),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_73),
.A2(n_20),
.B1(n_33),
.B2(n_31),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_53),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_114),
.B(n_117),
.Y(n_125)
);

INVx1_ASAP7_75t_SL g115 ( 
.A(n_63),
.Y(n_115)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_115),
.Y(n_139)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_75),
.Y(n_117)
);

AO21x1_ASAP7_75t_L g155 ( 
.A1(n_118),
.A2(n_128),
.B(n_80),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_87),
.A2(n_72),
.B1(n_45),
.B2(n_47),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_119),
.A2(n_123),
.B1(n_140),
.B2(n_144),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_121),
.B(n_129),
.C(n_130),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_79),
.A2(n_33),
.B1(n_31),
.B2(n_26),
.Y(n_123)
);

INVx2_ASAP7_75t_SL g124 ( 
.A(n_97),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_124),
.B(n_127),
.Y(n_156)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_86),
.Y(n_127)
);

XOR2xp5_ASAP7_75t_L g129 ( 
.A(n_109),
.B(n_33),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_108),
.B(n_71),
.C(n_26),
.Y(n_130)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_86),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_132),
.B(n_143),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g133 ( 
.A(n_89),
.B(n_26),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_133),
.B(n_135),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_81),
.B(n_22),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_102),
.A2(n_22),
.B1(n_32),
.B2(n_0),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_141),
.A2(n_148),
.B1(n_105),
.B2(n_104),
.Y(n_153)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_84),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_100),
.A2(n_32),
.B1(n_0),
.B2(n_3),
.Y(n_144)
);

BUFx24_ASAP7_75t_SL g146 ( 
.A(n_92),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_146),
.B(n_88),
.Y(n_177)
);

AOI21xp33_ASAP7_75t_L g147 ( 
.A1(n_116),
.A2(n_9),
.B(n_1),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_SL g171 ( 
.A1(n_147),
.A2(n_95),
.B(n_106),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_112),
.A2(n_0),
.B1(n_3),
.B2(n_5),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_110),
.B(n_5),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_149),
.B(n_152),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_110),
.B(n_6),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_153),
.B(n_155),
.Y(n_186)
);

INVxp67_ASAP7_75t_L g154 ( 
.A(n_134),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_154),
.B(n_157),
.Y(n_190)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_138),
.Y(n_157)
);

INVx4_ASAP7_75t_L g158 ( 
.A(n_145),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_158),
.B(n_161),
.Y(n_189)
);

AO21x2_ASAP7_75t_L g159 ( 
.A1(n_140),
.A2(n_111),
.B(n_96),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_SL g212 ( 
.A1(n_159),
.A2(n_182),
.B(n_128),
.Y(n_212)
);

INVx5_ASAP7_75t_L g161 ( 
.A(n_145),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_SL g162 ( 
.A(n_125),
.B(n_90),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_SL g198 ( 
.A(n_162),
.B(n_152),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_126),
.B(n_106),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_163),
.B(n_169),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_150),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_167),
.Y(n_193)
);

BUFx2_ASAP7_75t_L g168 ( 
.A(n_124),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_168),
.Y(n_195)
);

INVx8_ASAP7_75t_L g169 ( 
.A(n_124),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_120),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_170),
.Y(n_208)
);

CKINVDCx14_ASAP7_75t_R g213 ( 
.A(n_171),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_126),
.B(n_80),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_172),
.B(n_133),
.Y(n_191)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_151),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_173),
.B(n_174),
.Y(n_202)
);

CKINVDCx16_ASAP7_75t_R g174 ( 
.A(n_135),
.Y(n_174)
);

INVx3_ASAP7_75t_L g176 ( 
.A(n_127),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_176),
.B(n_177),
.Y(n_210)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_119),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_178),
.B(n_179),
.Y(n_211)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_148),
.Y(n_179)
);

INVx6_ASAP7_75t_SL g180 ( 
.A(n_132),
.Y(n_180)
);

INVx13_ASAP7_75t_L g206 ( 
.A(n_180),
.Y(n_206)
);

INVx3_ASAP7_75t_L g181 ( 
.A(n_122),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_181),
.Y(n_214)
);

AND2x2_ASAP7_75t_L g182 ( 
.A(n_121),
.B(n_6),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_144),
.Y(n_183)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_183),
.Y(n_192)
);

BUFx6f_ASAP7_75t_L g184 ( 
.A(n_137),
.Y(n_184)
);

BUFx5_ASAP7_75t_L g188 ( 
.A(n_184),
.Y(n_188)
);

INVx4_ASAP7_75t_L g185 ( 
.A(n_137),
.Y(n_185)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_185),
.Y(n_194)
);

MAJx2_ASAP7_75t_L g187 ( 
.A(n_160),
.B(n_129),
.C(n_142),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_SL g242 ( 
.A(n_187),
.B(n_9),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_191),
.B(n_196),
.Y(n_226)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_168),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_SL g197 ( 
.A(n_160),
.B(n_141),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_197),
.B(n_184),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_198),
.B(n_205),
.Y(n_227)
);

AND2x2_ASAP7_75t_L g199 ( 
.A(n_172),
.B(n_149),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_SL g220 ( 
.A1(n_199),
.A2(n_212),
.B(n_205),
.Y(n_220)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_156),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_201),
.B(n_203),
.Y(n_228)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_185),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_164),
.B(n_130),
.C(n_131),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_204),
.B(n_207),
.C(n_182),
.Y(n_221)
);

NOR2x1_ASAP7_75t_L g205 ( 
.A(n_159),
.B(n_128),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_164),
.B(n_123),
.Y(n_207)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_165),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_209),
.B(n_215),
.Y(n_232)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_159),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_SL g216 ( 
.A(n_166),
.B(n_139),
.Y(n_216)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_216),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_215),
.A2(n_175),
.B1(n_159),
.B2(n_155),
.Y(n_217)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_217),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_186),
.A2(n_159),
.B1(n_175),
.B2(n_166),
.Y(n_218)
);

CKINVDCx14_ASAP7_75t_R g255 ( 
.A(n_218),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_186),
.A2(n_171),
.B1(n_154),
.B2(n_182),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_219),
.B(n_238),
.Y(n_245)
);

AO21x1_ASAP7_75t_L g251 ( 
.A1(n_220),
.A2(n_235),
.B(n_198),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_221),
.B(n_222),
.C(n_237),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_197),
.B(n_136),
.C(n_115),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_213),
.A2(n_169),
.B1(n_180),
.B2(n_176),
.Y(n_223)
);

INVxp67_ASAP7_75t_L g259 ( 
.A(n_223),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_193),
.B(n_158),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_224),
.B(n_225),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_193),
.B(n_181),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_229),
.B(n_240),
.Y(n_252)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_202),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_231),
.B(n_233),
.Y(n_260)
);

INVxp67_ASAP7_75t_L g233 ( 
.A(n_189),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_200),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_234),
.B(n_239),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_211),
.A2(n_136),
.B1(n_107),
.B2(n_98),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_L g236 ( 
.A1(n_192),
.A2(n_107),
.B1(n_161),
.B2(n_91),
.Y(n_236)
);

A2O1A1Ixp33_ASAP7_75t_SL g250 ( 
.A1(n_236),
.A2(n_188),
.B(n_195),
.C(n_214),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_204),
.B(n_91),
.C(n_7),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_192),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_238)
);

INVxp67_ASAP7_75t_L g239 ( 
.A(n_188),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_191),
.B(n_8),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_187),
.B(n_16),
.C(n_10),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_241),
.B(n_242),
.C(n_207),
.Y(n_262)
);

OAI21xp5_ASAP7_75t_L g243 ( 
.A1(n_227),
.A2(n_212),
.B(n_216),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_243),
.B(n_217),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_235),
.B(n_214),
.Y(n_246)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_246),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_226),
.B(n_232),
.Y(n_247)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_247),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_230),
.B(n_199),
.Y(n_248)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_248),
.Y(n_271)
);

NOR4xp25_ASAP7_75t_L g249 ( 
.A(n_228),
.B(n_210),
.C(n_208),
.D(n_199),
.Y(n_249)
);

FAx1_ASAP7_75t_SL g266 ( 
.A(n_249),
.B(n_263),
.CI(n_237),
.CON(n_266),
.SN(n_266)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_250),
.A2(n_251),
.B1(n_256),
.B2(n_194),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_238),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_254),
.B(n_257),
.Y(n_281)
);

HAxp5_ASAP7_75t_SL g256 ( 
.A(n_223),
.B(n_208),
.CON(n_256),
.SN(n_256)
);

NOR3xp33_ASAP7_75t_L g257 ( 
.A(n_241),
.B(n_209),
.C(n_201),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_262),
.B(n_222),
.C(n_221),
.Y(n_267)
);

XNOR2x2_ASAP7_75t_L g263 ( 
.A(n_242),
.B(n_190),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_SL g285 ( 
.A(n_265),
.B(n_266),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_267),
.B(n_270),
.C(n_274),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_252),
.B(n_229),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_268),
.B(n_243),
.Y(n_291)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_252),
.B(n_240),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_L g272 ( 
.A1(n_259),
.A2(n_233),
.B1(n_206),
.B2(n_239),
.Y(n_272)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_272),
.Y(n_294)
);

O2A1O1Ixp33_ASAP7_75t_L g288 ( 
.A1(n_273),
.A2(n_256),
.B(n_251),
.C(n_247),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_244),
.B(n_194),
.C(n_203),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_L g275 ( 
.A1(n_259),
.A2(n_206),
.B1(n_195),
.B2(n_196),
.Y(n_275)
);

CKINVDCx16_ASAP7_75t_R g289 ( 
.A(n_275),
.Y(n_289)
);

XOR2xp5_ASAP7_75t_L g276 ( 
.A(n_244),
.B(n_10),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_276),
.B(n_279),
.C(n_267),
.Y(n_283)
);

BUFx2_ASAP7_75t_L g277 ( 
.A(n_250),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_277),
.B(n_280),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_L g278 ( 
.A1(n_253),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_L g287 ( 
.A1(n_278),
.A2(n_254),
.B1(n_245),
.B2(n_248),
.Y(n_287)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_262),
.B(n_263),
.Y(n_279)
);

INVx1_ASAP7_75t_SL g280 ( 
.A(n_258),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_283),
.B(n_292),
.C(n_295),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_269),
.B(n_261),
.Y(n_286)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_286),
.Y(n_300)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_287),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_288),
.A2(n_276),
.B1(n_13),
.B2(n_14),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_280),
.B(n_260),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_290),
.B(n_291),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_274),
.B(n_255),
.C(n_253),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_264),
.A2(n_250),
.B1(n_13),
.B2(n_14),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_SL g302 ( 
.A(n_293),
.B(n_12),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_270),
.B(n_250),
.C(n_13),
.Y(n_295)
);

OAI21xp5_ASAP7_75t_SL g296 ( 
.A1(n_284),
.A2(n_281),
.B(n_277),
.Y(n_296)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_296),
.Y(n_313)
);

OAI21xp5_ASAP7_75t_L g298 ( 
.A1(n_289),
.A2(n_271),
.B(n_265),
.Y(n_298)
);

AOI21xp5_ASAP7_75t_SL g308 ( 
.A1(n_298),
.A2(n_285),
.B(n_283),
.Y(n_308)
);

AO21x1_ASAP7_75t_L g299 ( 
.A1(n_288),
.A2(n_266),
.B(n_279),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_299),
.B(n_304),
.Y(n_312)
);

AOI21xp5_ASAP7_75t_L g301 ( 
.A1(n_294),
.A2(n_266),
.B(n_268),
.Y(n_301)
);

XOR2xp5_ASAP7_75t_L g311 ( 
.A(n_301),
.B(n_282),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_302),
.B(n_12),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_L g307 ( 
.A1(n_303),
.A2(n_295),
.B1(n_292),
.B2(n_285),
.Y(n_307)
);

INVx11_ASAP7_75t_L g306 ( 
.A(n_298),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_SL g315 ( 
.A(n_306),
.B(n_307),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_SL g314 ( 
.A(n_308),
.B(n_309),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_297),
.B(n_282),
.C(n_305),
.Y(n_310)
);

AND2x2_ASAP7_75t_L g318 ( 
.A(n_310),
.B(n_311),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_L g317 ( 
.A1(n_312),
.A2(n_303),
.B1(n_300),
.B2(n_297),
.Y(n_317)
);

INVxp33_ASAP7_75t_SL g316 ( 
.A(n_306),
.Y(n_316)
);

OR2x2_ASAP7_75t_L g321 ( 
.A(n_316),
.B(n_312),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_SL g319 ( 
.A(n_317),
.B(n_308),
.Y(n_319)
);

AOI21xp5_ASAP7_75t_L g322 ( 
.A1(n_319),
.A2(n_320),
.B(n_321),
.Y(n_322)
);

OAI21xp5_ASAP7_75t_L g320 ( 
.A1(n_315),
.A2(n_310),
.B(n_313),
.Y(n_320)
);

INVxp67_ASAP7_75t_L g323 ( 
.A(n_319),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_323),
.B(n_318),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_324),
.Y(n_325)
);

OAI21xp33_ASAP7_75t_R g326 ( 
.A1(n_325),
.A2(n_322),
.B(n_314),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_326),
.B(n_311),
.Y(n_327)
);


endmodule