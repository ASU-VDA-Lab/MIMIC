module real_jpeg_23541_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_286;
wire n_288;
wire n_166;
wire n_176;
wire n_292;
wire n_215;
wire n_221;
wire n_249;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_280;
wire n_64;
wire n_177;
wire n_291;
wire n_236;
wire n_47;
wire n_131;
wire n_271;
wire n_281;
wire n_163;
wire n_276;
wire n_22;
wire n_287;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_243;
wire n_173;
wire n_255;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_293;
wire n_48;
wire n_164;
wire n_200;
wire n_184;
wire n_275;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_155;
wire n_120;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_238;
wire n_76;
wire n_67;
wire n_79;
wire n_178;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_239;
wire n_162;
wire n_290;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_285;
wire n_172;
wire n_45;
wire n_211;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_148;
wire n_19;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_205;
wire n_195;
wire n_258;
wire n_289;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_103;
wire n_225;
wire n_259;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_284;
wire n_226;
wire n_277;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_279;
wire n_167;
wire n_128;
wire n_213;
wire n_179;
wire n_216;
wire n_202;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_210;
wire n_53;
wire n_127;
wire n_206;
wire n_224;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_181;
wire n_283;
wire n_101;
wire n_256;
wire n_274;
wire n_182;
wire n_273;
wire n_96;
wire n_269;
wire n_253;
wire n_89;

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_0),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g35 ( 
.A1(n_1),
.A2(n_27),
.B1(n_28),
.B2(n_36),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_1),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_1),
.A2(n_36),
.B1(n_42),
.B2(n_43),
.Y(n_96)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_2),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_3),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_3),
.B(n_82),
.Y(n_172)
);

O2A1O1Ixp33_ASAP7_75t_L g209 ( 
.A1(n_3),
.A2(n_58),
.B(n_61),
.C(n_210),
.Y(n_209)
);

AOI22xp33_ASAP7_75t_L g223 ( 
.A1(n_3),
.A2(n_61),
.B1(n_62),
.B2(n_157),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_3),
.B(n_28),
.C(n_48),
.Y(n_231)
);

AOI22xp33_ASAP7_75t_L g234 ( 
.A1(n_3),
.A2(n_42),
.B1(n_43),
.B2(n_157),
.Y(n_234)
);

OAI21xp5_ASAP7_75t_SL g244 ( 
.A1(n_3),
.A2(n_31),
.B(n_245),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_3),
.B(n_148),
.Y(n_256)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_5),
.A2(n_61),
.B1(n_62),
.B2(n_65),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_5),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_5),
.A2(n_65),
.B1(n_71),
.B2(n_111),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_5),
.A2(n_42),
.B1(n_43),
.B2(n_65),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_L g174 ( 
.A1(n_5),
.A2(n_27),
.B1(n_28),
.B2(n_65),
.Y(n_174)
);

INVx8_ASAP7_75t_SL g79 ( 
.A(n_6),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_7),
.A2(n_70),
.B1(n_71),
.B2(n_73),
.Y(n_69)
);

CKINVDCx16_ASAP7_75t_R g70 ( 
.A(n_7),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_7),
.A2(n_61),
.B1(n_62),
.B2(n_70),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_7),
.A2(n_42),
.B1(n_43),
.B2(n_70),
.Y(n_205)
);

AOI22xp33_ASAP7_75t_L g239 ( 
.A1(n_7),
.A2(n_27),
.B1(n_28),
.B2(n_70),
.Y(n_239)
);

BUFx5_ASAP7_75t_L g58 ( 
.A(n_8),
.Y(n_58)
);

INVx13_ASAP7_75t_L g72 ( 
.A(n_9),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_L g41 ( 
.A1(n_10),
.A2(n_42),
.B1(n_43),
.B2(n_45),
.Y(n_41)
);

CKINVDCx14_ASAP7_75t_R g45 ( 
.A(n_10),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_10),
.A2(n_45),
.B1(n_61),
.B2(n_62),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_10),
.A2(n_27),
.B1(n_28),
.B2(n_45),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_SL g26 ( 
.A1(n_11),
.A2(n_27),
.B1(n_28),
.B2(n_30),
.Y(n_26)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_11),
.A2(n_30),
.B1(n_42),
.B2(n_43),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_L g85 ( 
.A1(n_12),
.A2(n_73),
.B1(n_80),
.B2(n_86),
.Y(n_85)
);

CKINVDCx14_ASAP7_75t_R g86 ( 
.A(n_12),
.Y(n_86)
);

OAI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_12),
.A2(n_61),
.B1(n_62),
.B2(n_86),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_12),
.A2(n_42),
.B1(n_43),
.B2(n_86),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_12),
.A2(n_27),
.B1(n_28),
.B2(n_86),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_13),
.A2(n_71),
.B1(n_72),
.B2(n_135),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_13),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_13),
.A2(n_61),
.B1(n_62),
.B2(n_135),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_L g220 ( 
.A1(n_13),
.A2(n_42),
.B1(n_43),
.B2(n_135),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_13),
.A2(n_27),
.B1(n_28),
.B2(n_135),
.Y(n_237)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_14),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g52 ( 
.A1(n_15),
.A2(n_42),
.B1(n_43),
.B2(n_53),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_15),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_15),
.A2(n_53),
.B1(n_61),
.B2(n_62),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_15),
.A2(n_27),
.B1(n_28),
.B2(n_53),
.Y(n_125)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_16),
.A2(n_32),
.B1(n_125),
.B2(n_163),
.Y(n_162)
);

INVx6_ASAP7_75t_L g177 ( 
.A(n_16),
.Y(n_177)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_16),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_16),
.A2(n_32),
.B1(n_236),
.B2(n_238),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_138),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_136),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_116),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_20),
.B(n_116),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_22),
.B1(n_87),
.B2(n_115),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_55),
.C(n_67),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_23),
.A2(n_24),
.B1(n_118),
.B2(n_119),
.Y(n_117)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_38),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_25),
.A2(n_38),
.B1(n_39),
.B2(n_282),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_25),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_SL g25 ( 
.A1(n_26),
.A2(n_31),
.B1(n_35),
.B2(n_37),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_26),
.A2(n_31),
.B1(n_34),
.B2(n_124),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_27),
.B(n_33),
.Y(n_32)
);

OA22x2_ASAP7_75t_L g51 ( 
.A1(n_27),
.A2(n_28),
.B1(n_48),
.B2(n_50),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_27),
.B(n_243),
.Y(n_242)
);

INVx6_ASAP7_75t_SL g27 ( 
.A(n_28),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

AOI21xp5_ASAP7_75t_L g101 ( 
.A1(n_31),
.A2(n_35),
.B(n_102),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_31),
.A2(n_164),
.B1(n_174),
.B2(n_175),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_L g259 ( 
.A1(n_31),
.A2(n_239),
.B(n_245),
.Y(n_259)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_32),
.B(n_214),
.Y(n_213)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx5_ASAP7_75t_L g103 ( 
.A(n_34),
.Y(n_103)
);

INVx3_ASAP7_75t_L g246 ( 
.A(n_37),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_L g248 ( 
.A1(n_37),
.A2(n_213),
.B(n_237),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_39),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g39 ( 
.A1(n_40),
.A2(n_46),
.B1(n_52),
.B2(n_54),
.Y(n_39)
);

INVxp67_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_41),
.A2(n_51),
.B1(n_93),
.B2(n_127),
.Y(n_126)
);

OAI22xp33_ASAP7_75t_L g47 ( 
.A1(n_42),
.A2(n_43),
.B1(n_48),
.B2(n_50),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_42),
.A2(n_43),
.B1(n_58),
.B2(n_59),
.Y(n_57)
);

OAI21xp33_ASAP7_75t_L g210 ( 
.A1(n_42),
.A2(n_59),
.B(n_157),
.Y(n_210)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_43),
.B(n_231),
.Y(n_230)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_46),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_46),
.A2(n_52),
.B1(n_54),
.B2(n_95),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_46),
.B(n_153),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_46),
.A2(n_54),
.B1(n_205),
.B2(n_219),
.Y(n_218)
);

AND2x2_ASAP7_75t_L g46 ( 
.A(n_47),
.B(n_51),
.Y(n_46)
);

INVx13_ASAP7_75t_L g50 ( 
.A(n_48),
.Y(n_50)
);

BUFx24_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_51),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_51),
.A2(n_93),
.B1(n_94),
.B2(n_96),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_L g151 ( 
.A1(n_51),
.A2(n_127),
.B(n_152),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_51),
.B(n_157),
.Y(n_249)
);

OAI21xp5_ASAP7_75t_L g258 ( 
.A1(n_51),
.A2(n_152),
.B(n_220),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_54),
.B(n_153),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_SL g119 ( 
.A(n_55),
.B(n_67),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_56),
.A2(n_57),
.B1(n_64),
.B2(n_66),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_56),
.A2(n_57),
.B1(n_66),
.B2(n_91),
.Y(n_90)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_56),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_SL g181 ( 
.A1(n_56),
.A2(n_182),
.B(n_183),
.Y(n_181)
);

OAI21xp33_ASAP7_75t_L g222 ( 
.A1(n_56),
.A2(n_183),
.B(n_223),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_57),
.B(n_60),
.Y(n_56)
);

OAI21xp5_ASAP7_75t_L g129 ( 
.A1(n_57),
.A2(n_64),
.B(n_130),
.Y(n_129)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_57),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_SL g169 ( 
.A1(n_57),
.A2(n_130),
.B(n_170),
.Y(n_169)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_58),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_58),
.A2(n_59),
.B1(n_61),
.B2(n_62),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_61),
.A2(n_62),
.B1(n_78),
.B2(n_79),
.Y(n_82)
);

NAND3xp33_ASAP7_75t_SL g167 ( 
.A(n_61),
.B(n_79),
.C(n_112),
.Y(n_167)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

A2O1A1Ixp33_ASAP7_75t_L g166 ( 
.A1(n_62),
.A2(n_78),
.B(n_158),
.C(n_167),
.Y(n_166)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

OAI21xp5_ASAP7_75t_L g67 ( 
.A1(n_68),
.A2(n_75),
.B(n_83),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_69),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_69),
.A2(n_76),
.B1(n_82),
.B2(n_134),
.Y(n_133)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx11_ASAP7_75t_L g74 ( 
.A(n_72),
.Y(n_74)
);

INVx8_ASAP7_75t_L g80 ( 
.A(n_72),
.Y(n_80)
);

INVx6_ASAP7_75t_L g112 ( 
.A(n_72),
.Y(n_112)
);

OAI22xp33_ASAP7_75t_L g77 ( 
.A1(n_73),
.A2(n_78),
.B1(n_79),
.B2(n_80),
.Y(n_77)
);

INVx8_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_74),
.B(n_157),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_76),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_76),
.B(n_114),
.Y(n_113)
);

AOI21xp5_ASAP7_75t_L g154 ( 
.A1(n_76),
.A2(n_84),
.B(n_155),
.Y(n_154)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_77),
.B(n_81),
.Y(n_76)
);

INVx8_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_81),
.B(n_85),
.Y(n_84)
);

OAI21xp5_ASAP7_75t_L g109 ( 
.A1(n_81),
.A2(n_110),
.B(n_113),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_L g184 ( 
.A1(n_81),
.A2(n_113),
.B(n_185),
.Y(n_184)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVxp67_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_85),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_87),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_88),
.A2(n_89),
.B1(n_98),
.B2(n_99),
.Y(n_87)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

AOI21xp5_ASAP7_75t_L g89 ( 
.A1(n_90),
.A2(n_92),
.B(n_97),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_90),
.B(n_92),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_SL g203 ( 
.A1(n_93),
.A2(n_204),
.B(n_206),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_SL g233 ( 
.A1(n_93),
.A2(n_206),
.B(n_234),
.Y(n_233)
);

CKINVDCx14_ASAP7_75t_R g94 ( 
.A(n_95),
.Y(n_94)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

XOR2xp5_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_106),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_104),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_101),
.A2(n_107),
.B1(n_108),
.B2(n_109),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_101),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_101),
.A2(n_104),
.B1(n_105),
.B2(n_107),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g243 ( 
.A(n_102),
.B(n_157),
.Y(n_243)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_105),
.Y(n_104)
);

CKINVDCx14_ASAP7_75t_R g108 ( 
.A(n_109),
.Y(n_108)
);

INVx8_ASAP7_75t_L g156 ( 
.A(n_111),
.Y(n_156)
);

INVx8_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_120),
.C(n_121),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_117),
.B(n_120),
.Y(n_292)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_121),
.B(n_292),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_128),
.C(n_133),
.Y(n_121)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_122),
.B(n_285),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_126),
.Y(n_122)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_123),
.B(n_126),
.Y(n_188)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_128),
.A2(n_129),
.B1(n_133),
.B2(n_286),
.Y(n_285)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_132),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_131),
.B(n_148),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_132),
.A2(n_147),
.B1(n_148),
.B2(n_149),
.Y(n_146)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_133),
.Y(n_286)
);

INVxp67_ASAP7_75t_L g185 ( 
.A(n_134),
.Y(n_185)
);

INVxp67_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_SL g138 ( 
.A1(n_139),
.A2(n_289),
.B(n_293),
.Y(n_138)
);

O2A1O1Ixp33_ASAP7_75t_SL g139 ( 
.A1(n_140),
.A2(n_191),
.B(n_276),
.C(n_288),
.Y(n_139)
);

AND2x2_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_178),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g192 ( 
.A(n_141),
.B(n_178),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_159),
.C(n_168),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_142),
.A2(n_143),
.B1(n_271),
.B2(n_272),
.Y(n_270)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

XOR2xp5_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_154),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_145),
.A2(n_146),
.B1(n_150),
.B2(n_151),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_146),
.B(n_150),
.C(n_154),
.Y(n_189)
);

CKINVDCx16_ASAP7_75t_R g170 ( 
.A(n_147),
.Y(n_170)
);

CKINVDCx14_ASAP7_75t_R g182 ( 
.A(n_149),
.Y(n_182)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

OAI21xp33_ASAP7_75t_L g155 ( 
.A1(n_156),
.A2(n_157),
.B(n_158),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_159),
.A2(n_160),
.B1(n_168),
.B2(n_273),
.Y(n_272)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_161),
.A2(n_162),
.B1(n_165),
.B2(n_166),
.Y(n_160)
);

CKINVDCx14_ASAP7_75t_R g161 ( 
.A(n_162),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_162),
.B(n_165),
.Y(n_180)
);

INVxp67_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

CKINVDCx14_ASAP7_75t_R g165 ( 
.A(n_166),
.Y(n_165)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_168),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_171),
.C(n_173),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_169),
.B(n_199),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_171),
.A2(n_172),
.B1(n_173),
.B2(n_200),
.Y(n_199)
);

CKINVDCx16_ASAP7_75t_R g171 ( 
.A(n_172),
.Y(n_171)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_173),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_L g211 ( 
.A1(n_174),
.A2(n_212),
.B(n_213),
.Y(n_211)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_179),
.A2(n_186),
.B1(n_187),
.B2(n_190),
.Y(n_178)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_179),
.Y(n_190)
);

BUFx24_ASAP7_75t_SL g294 ( 
.A(n_179),
.Y(n_294)
);

FAx1_ASAP7_75t_SL g179 ( 
.A(n_180),
.B(n_181),
.CI(n_184),
.CON(n_179),
.SN(n_179)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_180),
.B(n_181),
.C(n_184),
.Y(n_278)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_SL g187 ( 
.A(n_188),
.B(n_189),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_188),
.B(n_189),
.C(n_190),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_193),
.Y(n_191)
);

AOI21xp5_ASAP7_75t_SL g193 ( 
.A1(n_194),
.A2(n_269),
.B(n_275),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_L g194 ( 
.A1(n_195),
.A2(n_224),
.B(n_268),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_SL g195 ( 
.A(n_196),
.B(n_216),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_196),
.B(n_216),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_197),
.A2(n_198),
.B1(n_201),
.B2(n_215),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_197),
.B(n_203),
.C(n_207),
.Y(n_274)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_201),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_202),
.A2(n_203),
.B1(n_207),
.B2(n_208),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_205),
.Y(n_204)
);

CKINVDCx16_ASAP7_75t_R g207 ( 
.A(n_208),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_211),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_SL g217 ( 
.A(n_209),
.B(n_211),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_214),
.B(n_246),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_218),
.C(n_221),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_217),
.B(n_264),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_218),
.A2(n_221),
.B1(n_222),
.B2(n_265),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_218),
.Y(n_265)
);

INVxp67_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

AOI21xp5_ASAP7_75t_L g224 ( 
.A1(n_225),
.A2(n_262),
.B(n_267),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_L g225 ( 
.A1(n_226),
.A2(n_252),
.B(n_261),
.Y(n_225)
);

AOI21xp5_ASAP7_75t_L g226 ( 
.A1(n_227),
.A2(n_240),
.B(n_251),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_228),
.B(n_235),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_228),
.B(n_235),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_229),
.A2(n_230),
.B1(n_232),
.B2(n_233),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_230),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_230),
.B(n_232),
.Y(n_260)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

CKINVDCx16_ASAP7_75t_R g236 ( 
.A(n_237),
.Y(n_236)
);

INVxp67_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

OAI21xp5_ASAP7_75t_L g240 ( 
.A1(n_241),
.A2(n_247),
.B(n_250),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_244),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_SL g247 ( 
.A(n_248),
.B(n_249),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_248),
.B(n_249),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_SL g252 ( 
.A(n_253),
.B(n_260),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_253),
.B(n_260),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_259),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_255),
.A2(n_256),
.B1(n_257),
.B2(n_258),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_255),
.B(n_258),
.C(n_259),
.Y(n_266)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_263),
.B(n_266),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_263),
.B(n_266),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_SL g269 ( 
.A(n_270),
.B(n_274),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_270),
.B(n_274),
.Y(n_275)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_277),
.B(n_287),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_277),
.B(n_287),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_278),
.B(n_279),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_278),
.B(n_281),
.C(n_283),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_280),
.A2(n_281),
.B1(n_283),
.B2(n_284),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_290),
.B(n_291),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_290),
.B(n_291),
.Y(n_293)
);


endmodule