module fake_jpeg_11283_n_481 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_481);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_481;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_419;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_1),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_16),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_4),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_3),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_16),
.Y(n_25)
);

INVx5_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_16),
.Y(n_29)
);

BUFx4f_ASAP7_75t_SL g30 ( 
.A(n_10),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

CKINVDCx16_ASAP7_75t_R g34 ( 
.A(n_12),
.Y(n_34)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_9),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_14),
.Y(n_36)
);

BUFx10_ASAP7_75t_L g37 ( 
.A(n_15),
.Y(n_37)
);

BUFx24_ASAP7_75t_L g38 ( 
.A(n_11),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_7),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_14),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_3),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_13),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_9),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_2),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_13),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_11),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_6),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_2),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_10),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_18),
.B(n_15),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_50),
.B(n_51),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_24),
.B(n_0),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_30),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_52),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_24),
.B(n_0),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_53),
.B(n_62),
.Y(n_117)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

INVx5_ASAP7_75t_L g103 ( 
.A(n_54),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_30),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_55),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_37),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_56),
.B(n_60),
.Y(n_102)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

HB1xp67_ASAP7_75t_L g108 ( 
.A(n_57),
.Y(n_108)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g144 ( 
.A(n_58),
.Y(n_144)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_39),
.Y(n_59)
);

BUFx2_ASAP7_75t_L g129 ( 
.A(n_59),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_37),
.Y(n_60)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_38),
.Y(n_61)
);

INVx5_ASAP7_75t_L g132 ( 
.A(n_61),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_17),
.B(n_0),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_30),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_63),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_30),
.Y(n_64)
);

INVx6_ASAP7_75t_L g126 ( 
.A(n_64),
.Y(n_126)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_25),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_65),
.B(n_87),
.Y(n_111)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_35),
.Y(n_66)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_66),
.Y(n_133)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_38),
.Y(n_67)
);

INVx5_ASAP7_75t_L g135 ( 
.A(n_67),
.Y(n_135)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_42),
.Y(n_68)
);

INVx6_ASAP7_75t_L g140 ( 
.A(n_68),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_25),
.B(n_0),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_69),
.B(n_84),
.Y(n_128)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_35),
.Y(n_70)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_70),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_30),
.Y(n_71)
);

INVx6_ASAP7_75t_L g150 ( 
.A(n_71),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_42),
.Y(n_72)
);

INVx8_ASAP7_75t_L g151 ( 
.A(n_72),
.Y(n_151)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_39),
.Y(n_73)
);

BUFx3_ASAP7_75t_L g147 ( 
.A(n_73),
.Y(n_147)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_39),
.Y(n_74)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_74),
.Y(n_124)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_28),
.Y(n_75)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_75),
.Y(n_143)
);

INVx1_ASAP7_75t_SL g76 ( 
.A(n_38),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_76),
.B(n_83),
.Y(n_100)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_41),
.Y(n_77)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_77),
.Y(n_113)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_29),
.Y(n_78)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_78),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_42),
.Y(n_79)
);

INVx4_ASAP7_75t_L g138 ( 
.A(n_79),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_42),
.Y(n_80)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_80),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_19),
.Y(n_81)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_81),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_37),
.B(n_1),
.C(n_2),
.Y(n_82)
);

AOI21xp5_ASAP7_75t_L g120 ( 
.A1(n_82),
.A2(n_26),
.B(n_43),
.Y(n_120)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_29),
.Y(n_83)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_35),
.Y(n_84)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_29),
.Y(n_85)
);

INVx4_ASAP7_75t_SL g123 ( 
.A(n_85),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_19),
.Y(n_86)
);

INVx11_ASAP7_75t_L g116 ( 
.A(n_86),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_27),
.B(n_36),
.Y(n_87)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_28),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_88),
.B(n_92),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_19),
.Y(n_89)
);

INVx11_ASAP7_75t_L g137 ( 
.A(n_89),
.Y(n_137)
);

BUFx24_ASAP7_75t_L g90 ( 
.A(n_38),
.Y(n_90)
);

OR2x2_ASAP7_75t_L g99 ( 
.A(n_90),
.B(n_91),
.Y(n_99)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_41),
.Y(n_91)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_28),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_27),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_93),
.B(n_94),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_22),
.Y(n_94)
);

INVx8_ASAP7_75t_L g95 ( 
.A(n_22),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_95),
.Y(n_106)
);

INVx6_ASAP7_75t_SL g96 ( 
.A(n_37),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_96),
.B(n_97),
.Y(n_134)
);

BUFx12f_ASAP7_75t_L g97 ( 
.A(n_48),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_81),
.A2(n_40),
.B1(n_37),
.B2(n_36),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_98),
.A2(n_22),
.B1(n_31),
.B2(n_33),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_68),
.B(n_49),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_101),
.B(n_115),
.Y(n_159)
);

AOI21xp33_ASAP7_75t_SL g107 ( 
.A1(n_90),
.A2(n_41),
.B(n_26),
.Y(n_107)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_107),
.B(n_41),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_90),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_110),
.B(n_142),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_76),
.A2(n_26),
.B1(n_48),
.B2(n_54),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g154 ( 
.A1(n_114),
.A2(n_125),
.B1(n_71),
.B2(n_77),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_57),
.B(n_49),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g161 ( 
.A(n_120),
.B(n_41),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_59),
.B(n_21),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_121),
.B(n_122),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_74),
.B(n_21),
.Y(n_122)
);

OA22x2_ASAP7_75t_L g125 ( 
.A1(n_75),
.A2(n_95),
.B1(n_61),
.B2(n_67),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_97),
.B(n_17),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_136),
.B(n_139),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_97),
.B(n_20),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g142 ( 
.A(n_52),
.B(n_20),
.Y(n_142)
);

OR2x2_ASAP7_75t_L g145 ( 
.A(n_55),
.B(n_45),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_145),
.B(n_148),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_86),
.B(n_45),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_146),
.B(n_6),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_63),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g149 ( 
.A(n_64),
.B(n_47),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_149),
.B(n_1),
.Y(n_185)
);

BUFx3_ASAP7_75t_L g152 ( 
.A(n_144),
.Y(n_152)
);

INVx5_ASAP7_75t_L g225 ( 
.A(n_152),
.Y(n_225)
);

AOI22xp33_ASAP7_75t_L g153 ( 
.A1(n_141),
.A2(n_94),
.B1(n_89),
.B2(n_34),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_153),
.A2(n_166),
.B1(n_173),
.B2(n_179),
.Y(n_216)
);

AOI21xp5_ASAP7_75t_L g247 ( 
.A1(n_154),
.A2(n_171),
.B(n_103),
.Y(n_247)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_143),
.Y(n_155)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_155),
.Y(n_208)
);

AND2x2_ASAP7_75t_L g227 ( 
.A(n_156),
.B(n_161),
.Y(n_227)
);

INVx5_ASAP7_75t_L g157 ( 
.A(n_126),
.Y(n_157)
);

INVx3_ASAP7_75t_L g205 ( 
.A(n_157),
.Y(n_205)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_143),
.Y(n_158)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_158),
.Y(n_235)
);

INVx6_ASAP7_75t_L g160 ( 
.A(n_151),
.Y(n_160)
);

INVx6_ASAP7_75t_L g212 ( 
.A(n_160),
.Y(n_212)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_130),
.Y(n_163)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_163),
.Y(n_204)
);

AOI22xp33_ASAP7_75t_SL g164 ( 
.A1(n_107),
.A2(n_32),
.B1(n_48),
.B2(n_125),
.Y(n_164)
);

INVxp67_ASAP7_75t_L g209 ( 
.A(n_164),
.Y(n_209)
);

INVx3_ASAP7_75t_L g165 ( 
.A(n_126),
.Y(n_165)
);

INVx4_ASAP7_75t_L g218 ( 
.A(n_165),
.Y(n_218)
);

AOI22xp33_ASAP7_75t_L g166 ( 
.A1(n_141),
.A2(n_34),
.B1(n_79),
.B2(n_72),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_102),
.Y(n_167)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_167),
.Y(n_214)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_104),
.Y(n_168)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_168),
.Y(n_229)
);

AOI21xp33_ASAP7_75t_L g169 ( 
.A1(n_128),
.A2(n_43),
.B(n_47),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_SL g210 ( 
.A(n_169),
.B(n_185),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_120),
.B(n_32),
.C(n_80),
.Y(n_170)
);

AND2x2_ASAP7_75t_L g248 ( 
.A(n_170),
.B(n_178),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_SL g171 ( 
.A1(n_115),
.A2(n_23),
.B(n_73),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_101),
.A2(n_40),
.B1(n_46),
.B2(n_44),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_L g223 ( 
.A1(n_172),
.A2(n_176),
.B1(n_106),
.B2(n_138),
.Y(n_223)
);

OAI22xp33_ASAP7_75t_L g173 ( 
.A1(n_146),
.A2(n_58),
.B1(n_46),
.B2(n_44),
.Y(n_173)
);

FAx1_ASAP7_75t_SL g174 ( 
.A(n_121),
.B(n_122),
.CI(n_117),
.CON(n_174),
.SN(n_174)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_174),
.B(n_195),
.Y(n_206)
);

BUFx6f_ASAP7_75t_L g175 ( 
.A(n_151),
.Y(n_175)
);

INVx3_ASAP7_75t_L g221 ( 
.A(n_175),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_145),
.A2(n_112),
.B1(n_99),
.B2(n_104),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_131),
.Y(n_177)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_177),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_133),
.B(n_40),
.C(n_46),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_SL g181 ( 
.A1(n_125),
.A2(n_23),
.B1(n_33),
.B2(n_31),
.Y(n_181)
);

INVxp67_ASAP7_75t_L g239 ( 
.A(n_181),
.Y(n_239)
);

AOI22xp33_ASAP7_75t_L g182 ( 
.A1(n_131),
.A2(n_33),
.B1(n_31),
.B2(n_44),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_182),
.A2(n_184),
.B1(n_186),
.B2(n_188),
.Y(n_217)
);

AOI22xp33_ASAP7_75t_L g184 ( 
.A1(n_116),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_184)
);

OAI22xp33_ASAP7_75t_SL g186 ( 
.A1(n_99),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_186)
);

AND2x2_ASAP7_75t_L g187 ( 
.A(n_100),
.B(n_13),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_187),
.B(n_192),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_140),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_188)
);

INVx13_ASAP7_75t_L g189 ( 
.A(n_123),
.Y(n_189)
);

BUFx10_ASAP7_75t_L g231 ( 
.A(n_189),
.Y(n_231)
);

BUFx6f_ASAP7_75t_L g190 ( 
.A(n_109),
.Y(n_190)
);

INVx3_ASAP7_75t_L g246 ( 
.A(n_190),
.Y(n_246)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_124),
.Y(n_191)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_191),
.Y(n_226)
);

OAI22xp33_ASAP7_75t_L g193 ( 
.A1(n_125),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_193),
.A2(n_138),
.B1(n_137),
.B2(n_116),
.Y(n_233)
);

INVx8_ASAP7_75t_L g194 ( 
.A(n_109),
.Y(n_194)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_194),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_108),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_105),
.B(n_8),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_196),
.B(n_10),
.Y(n_215)
);

HB1xp67_ASAP7_75t_L g197 ( 
.A(n_119),
.Y(n_197)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_197),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_111),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_198),
.B(n_201),
.Y(n_219)
);

INVx1_ASAP7_75t_SL g199 ( 
.A(n_100),
.Y(n_199)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_199),
.Y(n_249)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_124),
.Y(n_200)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_200),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_100),
.B(n_8),
.Y(n_201)
);

INVxp67_ASAP7_75t_L g203 ( 
.A(n_134),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_SL g228 ( 
.A(n_203),
.B(n_123),
.Y(n_228)
);

AOI22xp33_ASAP7_75t_SL g211 ( 
.A1(n_199),
.A2(n_129),
.B1(n_150),
.B2(n_135),
.Y(n_211)
);

INVxp67_ASAP7_75t_L g250 ( 
.A(n_211),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_SL g254 ( 
.A(n_215),
.B(n_228),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_159),
.B(n_133),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_220),
.B(n_222),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_159),
.B(n_106),
.Y(n_222)
);

OAI21xp33_ASAP7_75t_SL g252 ( 
.A1(n_223),
.A2(n_244),
.B(n_177),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_174),
.B(n_140),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_224),
.B(n_230),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_174),
.B(n_119),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_162),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_232),
.B(n_204),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_233),
.A2(n_245),
.B1(n_173),
.B2(n_193),
.Y(n_266)
);

AOI22xp33_ASAP7_75t_SL g236 ( 
.A1(n_176),
.A2(n_129),
.B1(n_150),
.B2(n_135),
.Y(n_236)
);

INVxp67_ASAP7_75t_L g283 ( 
.A(n_236),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_SL g237 ( 
.A(n_203),
.B(n_144),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_SL g285 ( 
.A(n_237),
.B(n_242),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_180),
.B(n_113),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_240),
.B(n_243),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_SL g242 ( 
.A(n_202),
.B(n_144),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_180),
.B(n_113),
.Y(n_243)
);

AOI22xp33_ASAP7_75t_L g244 ( 
.A1(n_172),
.A2(n_137),
.B1(n_118),
.B2(n_127),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_170),
.A2(n_179),
.B1(n_192),
.B2(n_156),
.Y(n_245)
);

OAI21xp5_ASAP7_75t_SL g253 ( 
.A1(n_247),
.A2(n_161),
.B(n_183),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_231),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_251),
.B(n_260),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_252),
.A2(n_277),
.B1(n_286),
.B2(n_205),
.Y(n_321)
);

AOI21xp5_ASAP7_75t_L g292 ( 
.A1(n_253),
.A2(n_255),
.B(n_258),
.Y(n_292)
);

AOI21xp5_ASAP7_75t_L g255 ( 
.A1(n_247),
.A2(n_209),
.B(n_239),
.Y(n_255)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_207),
.Y(n_257)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_257),
.Y(n_293)
);

AOI21xp5_ASAP7_75t_L g258 ( 
.A1(n_209),
.A2(n_239),
.B(n_230),
.Y(n_258)
);

BUFx8_ASAP7_75t_L g259 ( 
.A(n_231),
.Y(n_259)
);

INVx13_ASAP7_75t_L g301 ( 
.A(n_259),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_231),
.Y(n_260)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_207),
.Y(n_263)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_263),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_227),
.B(n_161),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_264),
.B(n_268),
.C(n_275),
.Y(n_303)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_226),
.Y(n_265)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_265),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_SL g312 ( 
.A1(n_266),
.A2(n_267),
.B1(n_271),
.B2(n_290),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_245),
.A2(n_216),
.B1(n_248),
.B2(n_217),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_227),
.B(n_224),
.Y(n_268)
);

CKINVDCx14_ASAP7_75t_R g316 ( 
.A(n_269),
.Y(n_316)
);

OAI21xp5_ASAP7_75t_SL g270 ( 
.A1(n_227),
.A2(n_171),
.B(n_187),
.Y(n_270)
);

OAI21xp5_ASAP7_75t_L g322 ( 
.A1(n_270),
.A2(n_274),
.B(n_289),
.Y(n_322)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_216),
.A2(n_163),
.B1(n_187),
.B2(n_178),
.Y(n_271)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_226),
.Y(n_272)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_272),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_222),
.B(n_201),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_273),
.B(n_278),
.Y(n_300)
);

NAND2x1p5_ASAP7_75t_L g274 ( 
.A(n_248),
.B(n_189),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_248),
.B(n_196),
.C(n_191),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_204),
.B(n_214),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_SL g294 ( 
.A(n_276),
.B(n_279),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_206),
.A2(n_188),
.B1(n_165),
.B2(n_160),
.Y(n_277)
);

A2O1A1Ixp33_ASAP7_75t_L g278 ( 
.A1(n_240),
.A2(n_158),
.B(n_155),
.C(n_200),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_210),
.B(n_152),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_229),
.Y(n_280)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_280),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_249),
.B(n_175),
.C(n_127),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_281),
.B(n_205),
.C(n_238),
.Y(n_310)
);

AO22x1_ASAP7_75t_SL g282 ( 
.A1(n_249),
.A2(n_194),
.B1(n_157),
.B2(n_190),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_282),
.B(n_241),
.Y(n_309)
);

CKINVDCx14_ASAP7_75t_R g284 ( 
.A(n_231),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_284),
.B(n_288),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_243),
.A2(n_118),
.B1(n_103),
.B2(n_132),
.Y(n_286)
);

INVx13_ASAP7_75t_L g287 ( 
.A(n_225),
.Y(n_287)
);

CKINVDCx16_ASAP7_75t_R g304 ( 
.A(n_287),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_220),
.Y(n_288)
);

OAI21xp5_ASAP7_75t_SL g289 ( 
.A1(n_213),
.A2(n_147),
.B(n_132),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_217),
.A2(n_147),
.B1(n_11),
.B2(n_12),
.Y(n_290)
);

INVxp33_ASAP7_75t_L g291 ( 
.A(n_212),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_291),
.B(n_221),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_268),
.B(n_213),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_SL g335 ( 
.A(n_296),
.B(n_307),
.Y(n_335)
);

OAI21xp5_ASAP7_75t_SL g298 ( 
.A1(n_258),
.A2(n_215),
.B(n_219),
.Y(n_298)
);

INVxp67_ASAP7_75t_L g331 ( 
.A(n_298),
.Y(n_331)
);

AND2x2_ASAP7_75t_L g299 ( 
.A(n_289),
.B(n_233),
.Y(n_299)
);

INVxp67_ASAP7_75t_L g332 ( 
.A(n_299),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_251),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_305),
.B(n_313),
.Y(n_351)
);

XNOR2xp5_ASAP7_75t_L g307 ( 
.A(n_256),
.B(n_234),
.Y(n_307)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_309),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g357 ( 
.A(n_310),
.B(n_282),
.C(n_246),
.Y(n_357)
);

BUFx3_ASAP7_75t_L g311 ( 
.A(n_259),
.Y(n_311)
);

INVx2_ASAP7_75t_L g360 ( 
.A(n_311),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_288),
.B(n_212),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_256),
.B(n_218),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_314),
.B(n_319),
.Y(n_359)
);

INVxp67_ASAP7_75t_L g333 ( 
.A(n_317),
.Y(n_333)
);

AOI21xp33_ASAP7_75t_L g318 ( 
.A1(n_285),
.A2(n_225),
.B(n_218),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_SL g350 ( 
.A(n_318),
.B(n_323),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_SL g319 ( 
.A(n_262),
.B(n_208),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_257),
.Y(n_320)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_320),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_L g334 ( 
.A1(n_321),
.A2(n_324),
.B1(n_250),
.B2(n_283),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_SL g323 ( 
.A(n_254),
.B(n_208),
.Y(n_323)
);

AOI22xp33_ASAP7_75t_SL g324 ( 
.A1(n_250),
.A2(n_283),
.B1(n_286),
.B2(n_260),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_SL g325 ( 
.A(n_262),
.B(n_235),
.Y(n_325)
);

XNOR2xp5_ASAP7_75t_SL g342 ( 
.A(n_325),
.B(n_261),
.Y(n_342)
);

AND2x6_ASAP7_75t_L g326 ( 
.A(n_253),
.B(n_221),
.Y(n_326)
);

OAI21xp5_ASAP7_75t_SL g338 ( 
.A1(n_326),
.A2(n_255),
.B(n_271),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_265),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_327),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_267),
.B(n_235),
.Y(n_328)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_328),
.Y(n_337)
);

XOR2xp5_ASAP7_75t_L g330 ( 
.A(n_303),
.B(n_296),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g365 ( 
.A(n_330),
.B(n_343),
.C(n_347),
.Y(n_365)
);

AOI22xp5_ASAP7_75t_L g387 ( 
.A1(n_334),
.A2(n_346),
.B1(n_356),
.B2(n_337),
.Y(n_387)
);

AO22x1_ASAP7_75t_L g336 ( 
.A1(n_322),
.A2(n_292),
.B1(n_299),
.B2(n_300),
.Y(n_336)
);

OAI21xp5_ASAP7_75t_SL g366 ( 
.A1(n_336),
.A2(n_309),
.B(n_314),
.Y(n_366)
);

INVxp67_ASAP7_75t_L g376 ( 
.A(n_338),
.Y(n_376)
);

OAI22xp5_ASAP7_75t_L g339 ( 
.A1(n_321),
.A2(n_266),
.B1(n_290),
.B2(n_254),
.Y(n_339)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_339),
.Y(n_361)
);

OAI22xp5_ASAP7_75t_L g341 ( 
.A1(n_316),
.A2(n_285),
.B1(n_261),
.B2(n_275),
.Y(n_341)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_341),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_L g382 ( 
.A(n_342),
.B(n_358),
.Y(n_382)
);

XNOR2xp5_ASAP7_75t_L g343 ( 
.A(n_303),
.B(n_264),
.Y(n_343)
);

AOI22xp5_ASAP7_75t_L g345 ( 
.A1(n_312),
.A2(n_277),
.B1(n_263),
.B2(n_274),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_L g368 ( 
.A1(n_345),
.A2(n_325),
.B1(n_319),
.B2(n_327),
.Y(n_368)
);

OAI22xp5_ASAP7_75t_SL g346 ( 
.A1(n_328),
.A2(n_270),
.B1(n_274),
.B2(n_273),
.Y(n_346)
);

XNOR2xp5_ASAP7_75t_L g347 ( 
.A(n_307),
.B(n_281),
.Y(n_347)
);

CKINVDCx20_ASAP7_75t_R g348 ( 
.A(n_308),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_348),
.B(n_353),
.Y(n_363)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_313),
.Y(n_349)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_349),
.Y(n_378)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_293),
.Y(n_352)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_352),
.Y(n_381)
);

CKINVDCx20_ASAP7_75t_R g353 ( 
.A(n_315),
.Y(n_353)
);

OAI21xp5_ASAP7_75t_SL g354 ( 
.A1(n_292),
.A2(n_278),
.B(n_272),
.Y(n_354)
);

AOI21xp5_ASAP7_75t_SL g374 ( 
.A1(n_354),
.A2(n_355),
.B(n_295),
.Y(n_374)
);

OAI21xp5_ASAP7_75t_SL g355 ( 
.A1(n_299),
.A2(n_282),
.B(n_280),
.Y(n_355)
);

OAI22xp5_ASAP7_75t_SL g356 ( 
.A1(n_300),
.A2(n_282),
.B1(n_238),
.B2(n_246),
.Y(n_356)
);

MAJIxp5_ASAP7_75t_L g372 ( 
.A(n_357),
.B(n_302),
.C(n_320),
.Y(n_372)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_293),
.Y(n_358)
);

XOR2xp5_ASAP7_75t_L g362 ( 
.A(n_330),
.B(n_322),
.Y(n_362)
);

XOR2xp5_ASAP7_75t_L g394 ( 
.A(n_362),
.B(n_331),
.Y(n_394)
);

NOR3xp33_ASAP7_75t_SL g364 ( 
.A(n_350),
.B(n_294),
.C(n_326),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_364),
.B(n_366),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_L g367 ( 
.A(n_340),
.B(n_294),
.Y(n_367)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_367),
.Y(n_388)
);

AOI22xp5_ASAP7_75t_L g402 ( 
.A1(n_368),
.A2(n_359),
.B1(n_358),
.B2(n_333),
.Y(n_402)
);

OAI22xp5_ASAP7_75t_L g369 ( 
.A1(n_329),
.A2(n_312),
.B1(n_305),
.B2(n_310),
.Y(n_369)
);

AOI22xp5_ASAP7_75t_L g397 ( 
.A1(n_369),
.A2(n_356),
.B1(n_349),
.B2(n_357),
.Y(n_397)
);

AOI21xp5_ASAP7_75t_L g370 ( 
.A1(n_332),
.A2(n_298),
.B(n_323),
.Y(n_370)
);

INVxp33_ASAP7_75t_L g389 ( 
.A(n_370),
.Y(n_389)
);

MAJIxp5_ASAP7_75t_L g391 ( 
.A(n_372),
.B(n_373),
.C(n_377),
.Y(n_391)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_343),
.B(n_347),
.C(n_335),
.Y(n_373)
);

OAI21xp33_ASAP7_75t_L g390 ( 
.A1(n_374),
.A2(n_351),
.B(n_336),
.Y(n_390)
);

OAI21xp5_ASAP7_75t_L g375 ( 
.A1(n_332),
.A2(n_295),
.B(n_297),
.Y(n_375)
);

XNOR2x2_ASAP7_75t_SL g398 ( 
.A(n_375),
.B(n_386),
.Y(n_398)
);

MAJIxp5_ASAP7_75t_L g377 ( 
.A(n_335),
.B(n_297),
.C(n_302),
.Y(n_377)
);

MAJIxp5_ASAP7_75t_L g379 ( 
.A(n_346),
.B(n_306),
.C(n_304),
.Y(n_379)
);

XNOR2xp5_ASAP7_75t_L g392 ( 
.A(n_379),
.B(n_336),
.Y(n_392)
);

NOR2xp33_ASAP7_75t_L g380 ( 
.A(n_342),
.B(n_306),
.Y(n_380)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_380),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_L g383 ( 
.A(n_329),
.B(n_344),
.Y(n_383)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_383),
.Y(n_395)
);

INVxp67_ASAP7_75t_L g384 ( 
.A(n_354),
.Y(n_384)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_384),
.Y(n_400)
);

CKINVDCx20_ASAP7_75t_R g385 ( 
.A(n_351),
.Y(n_385)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_385),
.Y(n_406)
);

OAI21xp5_ASAP7_75t_L g386 ( 
.A1(n_331),
.A2(n_311),
.B(n_301),
.Y(n_386)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_387),
.Y(n_407)
);

O2A1O1Ixp33_ASAP7_75t_L g422 ( 
.A1(n_390),
.A2(n_370),
.B(n_376),
.C(n_366),
.Y(n_422)
);

XOR2xp5_ASAP7_75t_L g412 ( 
.A(n_392),
.B(n_394),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_397),
.B(n_403),
.Y(n_413)
);

XOR2xp5_ASAP7_75t_L g399 ( 
.A(n_365),
.B(n_338),
.Y(n_399)
);

NOR2xp67_ASAP7_75t_SL g428 ( 
.A(n_399),
.B(n_405),
.Y(n_428)
);

AOI22xp5_ASAP7_75t_L g401 ( 
.A1(n_361),
.A2(n_337),
.B1(n_359),
.B2(n_345),
.Y(n_401)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_401),
.Y(n_415)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_402),
.Y(n_418)
);

AOI22xp5_ASAP7_75t_L g403 ( 
.A1(n_361),
.A2(n_355),
.B1(n_333),
.B2(n_360),
.Y(n_403)
);

AOI22xp5_ASAP7_75t_L g404 ( 
.A1(n_369),
.A2(n_360),
.B1(n_304),
.B2(n_301),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_404),
.B(n_386),
.Y(n_421)
);

XOR2xp5_ASAP7_75t_L g405 ( 
.A(n_365),
.B(n_287),
.Y(n_405)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_383),
.Y(n_408)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_408),
.Y(n_417)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_363),
.Y(n_409)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_409),
.Y(n_426)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_381),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_L g420 ( 
.A(n_410),
.B(n_395),
.Y(n_420)
);

AOI22xp5_ASAP7_75t_L g411 ( 
.A1(n_407),
.A2(n_368),
.B1(n_371),
.B2(n_385),
.Y(n_411)
);

INVxp33_ASAP7_75t_L g437 ( 
.A(n_411),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_SL g414 ( 
.A(n_388),
.B(n_371),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_414),
.B(n_416),
.Y(n_436)
);

MAJIxp5_ASAP7_75t_L g416 ( 
.A(n_391),
.B(n_372),
.C(n_373),
.Y(n_416)
);

AOI21xp5_ASAP7_75t_L g419 ( 
.A1(n_389),
.A2(n_384),
.B(n_376),
.Y(n_419)
);

OAI21xp5_ASAP7_75t_SL g435 ( 
.A1(n_419),
.A2(n_374),
.B(n_404),
.Y(n_435)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_420),
.Y(n_432)
);

OAI321xp33_ASAP7_75t_L g431 ( 
.A1(n_421),
.A2(n_425),
.A3(n_400),
.B1(n_398),
.B2(n_393),
.C(n_382),
.Y(n_431)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_422),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_406),
.B(n_378),
.Y(n_423)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_423),
.Y(n_442)
);

AOI22xp5_ASAP7_75t_SL g424 ( 
.A1(n_389),
.A2(n_379),
.B1(n_377),
.B2(n_378),
.Y(n_424)
);

XOR2xp5_ASAP7_75t_L g434 ( 
.A(n_424),
.B(n_392),
.Y(n_434)
);

FAx1_ASAP7_75t_SL g425 ( 
.A(n_396),
.B(n_390),
.CI(n_382),
.CON(n_425),
.SN(n_425)
);

BUFx24_ASAP7_75t_SL g427 ( 
.A(n_399),
.Y(n_427)
);

NOR2xp33_ASAP7_75t_SL g429 ( 
.A(n_427),
.B(n_428),
.Y(n_429)
);

NOR2xp33_ASAP7_75t_L g445 ( 
.A(n_429),
.B(n_417),
.Y(n_445)
);

MAJIxp5_ASAP7_75t_L g430 ( 
.A(n_416),
.B(n_391),
.C(n_405),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_430),
.B(n_438),
.Y(n_449)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_431),
.Y(n_453)
);

NOR2xp67_ASAP7_75t_SL g447 ( 
.A(n_434),
.B(n_418),
.Y(n_447)
);

OR2x2_ASAP7_75t_L g454 ( 
.A(n_435),
.B(n_425),
.Y(n_454)
);

MAJIxp5_ASAP7_75t_L g438 ( 
.A(n_412),
.B(n_362),
.C(n_397),
.Y(n_438)
);

MAJIxp5_ASAP7_75t_L g439 ( 
.A(n_412),
.B(n_398),
.C(n_394),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_439),
.B(n_440),
.Y(n_450)
);

MAJIxp5_ASAP7_75t_L g440 ( 
.A(n_424),
.B(n_375),
.C(n_403),
.Y(n_440)
);

AOI22xp5_ASAP7_75t_L g441 ( 
.A1(n_418),
.A2(n_364),
.B1(n_387),
.B2(n_401),
.Y(n_441)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_441),
.Y(n_456)
);

NOR2xp33_ASAP7_75t_SL g443 ( 
.A(n_426),
.B(n_381),
.Y(n_443)
);

NOR2xp33_ASAP7_75t_SL g452 ( 
.A(n_443),
.B(n_423),
.Y(n_452)
);

XOR2xp5_ASAP7_75t_L g444 ( 
.A(n_438),
.B(n_413),
.Y(n_444)
);

XNOR2xp5_ASAP7_75t_L g465 ( 
.A(n_444),
.B(n_455),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_SL g457 ( 
.A(n_445),
.B(n_446),
.Y(n_457)
);

MAJIxp5_ASAP7_75t_L g446 ( 
.A(n_430),
.B(n_413),
.C(n_421),
.Y(n_446)
);

XOR2xp5_ASAP7_75t_L g460 ( 
.A(n_447),
.B(n_435),
.Y(n_460)
);

AOI21xp5_ASAP7_75t_L g448 ( 
.A1(n_433),
.A2(n_419),
.B(n_411),
.Y(n_448)
);

OAI21xp5_ASAP7_75t_SL g459 ( 
.A1(n_448),
.A2(n_454),
.B(n_437),
.Y(n_459)
);

NOR2xp67_ASAP7_75t_SL g451 ( 
.A(n_434),
.B(n_415),
.Y(n_451)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_451),
.Y(n_458)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_452),
.Y(n_461)
);

MAJIxp5_ASAP7_75t_L g455 ( 
.A(n_440),
.B(n_415),
.C(n_422),
.Y(n_455)
);

HB1xp67_ASAP7_75t_L g462 ( 
.A(n_455),
.Y(n_462)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_459),
.Y(n_469)
);

NOR2xp67_ASAP7_75t_SL g471 ( 
.A(n_460),
.B(n_465),
.Y(n_471)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_453),
.Y(n_463)
);

AOI22xp5_ASAP7_75t_L g467 ( 
.A1(n_463),
.A2(n_464),
.B1(n_466),
.B2(n_437),
.Y(n_467)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_446),
.Y(n_464)
);

AOI322xp5_ASAP7_75t_L g466 ( 
.A1(n_456),
.A2(n_442),
.A3(n_432),
.B1(n_441),
.B2(n_454),
.C1(n_425),
.C2(n_448),
.Y(n_466)
);

AOI21xp5_ASAP7_75t_L g475 ( 
.A1(n_467),
.A2(n_468),
.B(n_460),
.Y(n_475)
);

OAI21xp5_ASAP7_75t_L g468 ( 
.A1(n_457),
.A2(n_436),
.B(n_449),
.Y(n_468)
);

AOI22xp5_ASAP7_75t_L g470 ( 
.A1(n_461),
.A2(n_444),
.B1(n_450),
.B2(n_439),
.Y(n_470)
);

NOR2xp33_ASAP7_75t_L g473 ( 
.A(n_470),
.B(n_458),
.Y(n_473)
);

MAJx2_ASAP7_75t_L g472 ( 
.A(n_462),
.B(n_301),
.C(n_287),
.Y(n_472)
);

OAI21xp5_ASAP7_75t_L g476 ( 
.A1(n_472),
.A2(n_259),
.B(n_11),
.Y(n_476)
);

NAND3xp33_ASAP7_75t_L g477 ( 
.A(n_473),
.B(n_474),
.C(n_475),
.Y(n_477)
);

OAI21xp5_ASAP7_75t_SL g474 ( 
.A1(n_471),
.A2(n_465),
.B(n_459),
.Y(n_474)
);

OAI21xp5_ASAP7_75t_SL g478 ( 
.A1(n_476),
.A2(n_469),
.B(n_259),
.Y(n_478)
);

OAI22xp5_ASAP7_75t_L g479 ( 
.A1(n_478),
.A2(n_13),
.B1(n_10),
.B2(n_12),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_479),
.B(n_477),
.Y(n_480)
);

XNOR2xp5_ASAP7_75t_L g481 ( 
.A(n_480),
.B(n_12),
.Y(n_481)
);


endmodule