module fake_jpeg_31876_n_59 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_59);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_59;

wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_23;
wire n_27;
wire n_55;
wire n_47;
wire n_22;
wire n_51;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_44;
wire n_28;
wire n_38;
wire n_26;
wire n_24;
wire n_36;
wire n_31;
wire n_25;
wire n_56;
wire n_37;
wire n_29;
wire n_43;
wire n_50;
wire n_32;

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_6),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_16),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_17),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_3),
.Y(n_23)
);

INVx5_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

BUFx2_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

INVx11_ASAP7_75t_L g35 ( 
.A(n_1),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_10),
.Y(n_36)
);

INVx5_ASAP7_75t_L g37 ( 
.A(n_35),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_37),
.B(n_38),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_L g38 ( 
.A1(n_27),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_29),
.B(n_5),
.Y(n_39)
);

MAJIxp5_ASAP7_75t_L g46 ( 
.A(n_39),
.B(n_40),
.C(n_41),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g40 ( 
.A1(n_21),
.A2(n_11),
.B1(n_12),
.B2(n_7),
.Y(n_40)
);

OA22x2_ASAP7_75t_L g41 ( 
.A1(n_30),
.A2(n_33),
.B1(n_31),
.B2(n_26),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_21),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_25),
.B(n_7),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_SL g44 ( 
.A1(n_27),
.A2(n_8),
.B1(n_29),
.B2(n_34),
.Y(n_44)
);

OAI32xp33_ASAP7_75t_L g47 ( 
.A1(n_45),
.A2(n_43),
.A3(n_40),
.B1(n_41),
.B2(n_39),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_47),
.A2(n_43),
.B1(n_44),
.B2(n_41),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g48 ( 
.A(n_46),
.B(n_18),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_L g50 ( 
.A1(n_48),
.A2(n_23),
.B1(n_36),
.B2(n_29),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_49),
.B(n_50),
.Y(n_52)
);

AOI322xp5_ASAP7_75t_L g51 ( 
.A1(n_49),
.A2(n_41),
.A3(n_22),
.B1(n_25),
.B2(n_42),
.C1(n_28),
.C2(n_32),
.Y(n_51)
);

MAJIxp5_ASAP7_75t_L g53 ( 
.A(n_51),
.B(n_52),
.C(n_22),
.Y(n_53)
);

MAJIxp5_ASAP7_75t_L g56 ( 
.A(n_53),
.B(n_54),
.C(n_42),
.Y(n_56)
);

XOR2xp5_ASAP7_75t_L g54 ( 
.A(n_52),
.B(n_19),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_54),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_55),
.B(n_56),
.Y(n_57)
);

AOI322xp5_ASAP7_75t_L g58 ( 
.A1(n_57),
.A2(n_20),
.A3(n_34),
.B1(n_32),
.B2(n_28),
.C1(n_25),
.C2(n_42),
.Y(n_58)
);

OAI221xp5_ASAP7_75t_L g59 ( 
.A1(n_58),
.A2(n_57),
.B1(n_20),
.B2(n_35),
.C(n_24),
.Y(n_59)
);


endmodule