module fake_jpeg_5057_n_9 (n_0, n_3, n_2, n_1, n_9);

input n_0;
input n_3;
input n_2;
input n_1;

output n_9;

wire n_4;
wire n_8;
wire n_6;
wire n_5;
wire n_7;

INVx2_ASAP7_75t_L g4 ( 
.A(n_1),
.Y(n_4)
);

INVx3_ASAP7_75t_L g5 ( 
.A(n_2),
.Y(n_5)
);

NAND2xp5_ASAP7_75t_L g6 ( 
.A(n_4),
.B(n_0),
.Y(n_6)
);

OAI22xp5_ASAP7_75t_SL g8 ( 
.A1(n_6),
.A2(n_7),
.B1(n_5),
.B2(n_2),
.Y(n_8)
);

MAJIxp5_ASAP7_75t_L g7 ( 
.A(n_5),
.B(n_0),
.C(n_1),
.Y(n_7)
);

NAND4xp25_ASAP7_75t_L g9 ( 
.A(n_8),
.B(n_0),
.C(n_3),
.D(n_6),
.Y(n_9)
);


endmodule