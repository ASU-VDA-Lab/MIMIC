module fake_jpeg_7305_n_75 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_75);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_75;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_23;
wire n_10;
wire n_69;
wire n_27;
wire n_55;
wire n_64;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_73;
wire n_19;
wire n_20;
wire n_18;
wire n_59;
wire n_35;
wire n_48;
wire n_68;
wire n_52;
wire n_71;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_65;
wire n_63;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_72;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_74;
wire n_11;
wire n_62;
wire n_17;
wire n_25;
wire n_31;
wire n_56;
wire n_67;
wire n_43;
wire n_37;
wire n_50;
wire n_29;
wire n_12;
wire n_32;
wire n_70;
wire n_15;
wire n_66;

CKINVDCx20_ASAP7_75t_R g9 ( 
.A(n_1),
.Y(n_9)
);

INVx1_ASAP7_75t_L g10 ( 
.A(n_6),
.Y(n_10)
);

INVx13_ASAP7_75t_L g11 ( 
.A(n_2),
.Y(n_11)
);

BUFx10_ASAP7_75t_L g12 ( 
.A(n_5),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_7),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_2),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_SL g15 ( 
.A(n_2),
.B(n_7),
.Y(n_15)
);

AND2x2_ASAP7_75t_L g16 ( 
.A(n_5),
.B(n_1),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_3),
.B(n_8),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_5),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_20),
.B(n_21),
.Y(n_34)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_17),
.Y(n_21)
);

AOI22xp33_ASAP7_75t_SL g22 ( 
.A1(n_11),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_22)
);

OAI21xp33_ASAP7_75t_L g36 ( 
.A1(n_22),
.A2(n_0),
.B(n_3),
.Y(n_36)
);

INVxp67_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_23),
.Y(n_28)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_24),
.B(n_25),
.Y(n_37)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

INVx13_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

HB1xp67_ASAP7_75t_L g29 ( 
.A(n_26),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_SL g27 ( 
.A(n_15),
.B(n_6),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_27),
.B(n_15),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_30),
.B(n_31),
.Y(n_41)
);

A2O1A1Ixp33_ASAP7_75t_L g31 ( 
.A1(n_23),
.A2(n_17),
.B(n_16),
.C(n_19),
.Y(n_31)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_20),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_32),
.B(n_33),
.Y(n_39)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_24),
.Y(n_33)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_25),
.Y(n_35)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

NAND3xp33_ASAP7_75t_L g46 ( 
.A(n_36),
.B(n_0),
.C(n_4),
.Y(n_46)
);

XOR2xp5_ASAP7_75t_L g38 ( 
.A(n_34),
.B(n_17),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_38),
.B(n_40),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g40 ( 
.A(n_30),
.B(n_16),
.Y(n_40)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_35),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_42),
.B(n_47),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g43 ( 
.A1(n_32),
.A2(n_26),
.B1(n_11),
.B2(n_18),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g49 ( 
.A1(n_43),
.A2(n_11),
.B1(n_33),
.B2(n_37),
.Y(n_49)
);

MAJIxp5_ASAP7_75t_L g44 ( 
.A(n_28),
.B(n_10),
.C(n_18),
.Y(n_44)
);

AOI21xp5_ASAP7_75t_L g53 ( 
.A1(n_44),
.A2(n_16),
.B(n_10),
.Y(n_53)
);

NOR2xp67_ASAP7_75t_SL g50 ( 
.A(n_46),
.B(n_16),
.Y(n_50)
);

INVxp67_ASAP7_75t_L g47 ( 
.A(n_37),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g60 ( 
.A1(n_49),
.A2(n_42),
.B1(n_14),
.B2(n_9),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_50),
.B(n_53),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_44),
.B(n_39),
.Y(n_52)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_52),
.Y(n_59)
);

AOI21xp5_ASAP7_75t_L g54 ( 
.A1(n_47),
.A2(n_31),
.B(n_28),
.Y(n_54)
);

O2A1O1Ixp33_ASAP7_75t_L g56 ( 
.A1(n_54),
.A2(n_41),
.B(n_38),
.C(n_14),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_43),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_55),
.B(n_45),
.Y(n_58)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_56),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_58),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g65 ( 
.A(n_60),
.B(n_9),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g61 ( 
.A1(n_54),
.A2(n_48),
.B1(n_49),
.B2(n_51),
.Y(n_61)
);

MAJIxp5_ASAP7_75t_L g64 ( 
.A(n_61),
.B(n_53),
.C(n_13),
.Y(n_64)
);

XNOR2xp5_ASAP7_75t_SL g68 ( 
.A(n_64),
.B(n_61),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g67 ( 
.A(n_65),
.B(n_60),
.Y(n_67)
);

HB1xp67_ASAP7_75t_SL g66 ( 
.A(n_62),
.Y(n_66)
);

OAI21xp5_ASAP7_75t_L g69 ( 
.A1(n_66),
.A2(n_68),
.B(n_64),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_67),
.B(n_63),
.Y(n_70)
);

A2O1A1Ixp33_ASAP7_75t_SL g72 ( 
.A1(n_69),
.A2(n_56),
.B(n_57),
.C(n_19),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_70),
.B(n_59),
.Y(n_71)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_71),
.Y(n_73)
);

OAI21xp5_ASAP7_75t_L g74 ( 
.A1(n_73),
.A2(n_72),
.B(n_8),
.Y(n_74)
);

AOI322xp5_ASAP7_75t_L g75 ( 
.A1(n_74),
.A2(n_4),
.A3(n_12),
.B1(n_29),
.B2(n_73),
.C1(n_66),
.C2(n_63),
.Y(n_75)
);


endmodule