module fake_jpeg_27279_n_273 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_273);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_273;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_272;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_212;
wire n_131;
wire n_56;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_258;
wire n_96;

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_14),
.B(n_3),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_16),
.Y(n_20)
);

BUFx4f_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_12),
.Y(n_23)
);

INVx6_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_4),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_5),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_16),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

INVxp67_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_12),
.Y(n_33)
);

BUFx16f_ASAP7_75t_L g34 ( 
.A(n_4),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_36),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_17),
.Y(n_37)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_29),
.B(n_1),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_38),
.B(n_41),
.Y(n_47)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

INVx11_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

INVx5_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_19),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_18),
.B(n_1),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_42),
.B(n_32),
.Y(n_46)
);

INVx11_ASAP7_75t_L g43 ( 
.A(n_18),
.Y(n_43)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_43),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_18),
.Y(n_44)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_44),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_39),
.A2(n_24),
.B1(n_33),
.B2(n_23),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_45),
.A2(n_49),
.B1(n_55),
.B2(n_57),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_46),
.B(n_66),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_39),
.A2(n_24),
.B1(n_33),
.B2(n_23),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_52),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_42),
.A2(n_29),
.B1(n_21),
.B2(n_31),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_54),
.A2(n_43),
.B1(n_40),
.B2(n_28),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_39),
.A2(n_26),
.B1(n_25),
.B2(n_30),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_41),
.B(n_25),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_SL g72 ( 
.A(n_56),
.B(n_27),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_39),
.A2(n_26),
.B1(n_31),
.B2(n_30),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_58),
.B(n_61),
.Y(n_68)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_42),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_41),
.B(n_32),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_62),
.B(n_38),
.Y(n_69)
);

BUFx8_ASAP7_75t_L g63 ( 
.A(n_40),
.Y(n_63)
);

INVx13_ASAP7_75t_L g91 ( 
.A(n_63),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_40),
.A2(n_21),
.B1(n_20),
.B2(n_22),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_64),
.A2(n_40),
.B1(n_43),
.B2(n_35),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_38),
.B(n_21),
.Y(n_66)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_63),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_67),
.A2(n_60),
.B1(n_50),
.B2(n_48),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_69),
.B(n_70),
.Y(n_102)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_51),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_64),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_71),
.B(n_72),
.Y(n_110)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_51),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_74),
.B(n_75),
.Y(n_116)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_51),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_47),
.B(n_61),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_76),
.B(n_88),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_77),
.A2(n_87),
.B1(n_65),
.B2(n_44),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_47),
.B(n_41),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_78),
.B(n_79),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_58),
.B(n_36),
.Y(n_79)
);

OR2x2_ASAP7_75t_L g81 ( 
.A(n_54),
.B(n_36),
.Y(n_81)
);

OAI21xp5_ASAP7_75t_SL g109 ( 
.A1(n_81),
.A2(n_44),
.B(n_37),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_56),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_82),
.Y(n_112)
);

BUFx12_ASAP7_75t_L g83 ( 
.A(n_63),
.Y(n_83)
);

INVx13_ASAP7_75t_L g107 ( 
.A(n_83),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_84),
.A2(n_90),
.B1(n_50),
.B2(n_53),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_46),
.B(n_32),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_85),
.B(n_36),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_48),
.A2(n_43),
.B1(n_20),
.B2(n_37),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_59),
.Y(n_88)
);

BUFx3_ASAP7_75t_L g89 ( 
.A(n_59),
.Y(n_89)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_89),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_L g90 ( 
.A1(n_66),
.A2(n_43),
.B1(n_20),
.B2(n_28),
.Y(n_90)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_63),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_92),
.B(n_52),
.Y(n_103)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_87),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_95),
.B(n_100),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_84),
.A2(n_50),
.B1(n_48),
.B2(n_53),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_SL g142 ( 
.A1(n_97),
.A2(n_109),
.B(n_37),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_98),
.A2(n_99),
.B1(n_104),
.B2(n_73),
.Y(n_120)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_77),
.Y(n_100)
);

A2O1A1Ixp33_ASAP7_75t_L g101 ( 
.A1(n_80),
.A2(n_34),
.B(n_32),
.C(n_28),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_L g119 ( 
.A(n_101),
.B(n_106),
.Y(n_119)
);

AND2x2_ASAP7_75t_L g123 ( 
.A(n_103),
.B(n_91),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_71),
.A2(n_60),
.B1(n_65),
.B2(n_27),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_105),
.B(n_115),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_L g106 ( 
.A(n_80),
.B(n_34),
.Y(n_106)
);

AND2x6_ASAP7_75t_L g108 ( 
.A(n_76),
.B(n_81),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_108),
.B(n_111),
.Y(n_126)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_79),
.Y(n_111)
);

AND2x6_ASAP7_75t_L g113 ( 
.A(n_81),
.B(n_1),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_113),
.B(n_114),
.Y(n_129)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_88),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_68),
.B(n_44),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_117),
.A2(n_70),
.B1(n_75),
.B2(n_74),
.Y(n_127)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_116),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_118),
.B(n_135),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_120),
.A2(n_121),
.B1(n_131),
.B2(n_133),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_100),
.A2(n_85),
.B1(n_68),
.B2(n_82),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_SL g167 ( 
.A1(n_123),
.A2(n_140),
.B(n_142),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g124 ( 
.A(n_106),
.B(n_93),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_124),
.B(n_115),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_127),
.A2(n_107),
.B1(n_113),
.B2(n_35),
.Y(n_163)
);

XOR2xp5_ASAP7_75t_L g128 ( 
.A(n_105),
.B(n_69),
.Y(n_128)
);

XOR2xp5_ASAP7_75t_L g149 ( 
.A(n_128),
.B(n_119),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_112),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_130),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_95),
.A2(n_78),
.B1(n_92),
.B2(n_86),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_94),
.B(n_72),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_132),
.B(n_136),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_99),
.A2(n_86),
.B1(n_67),
.B2(n_44),
.Y(n_133)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_96),
.Y(n_134)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_134),
.Y(n_150)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_116),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_94),
.B(n_89),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_102),
.B(n_28),
.Y(n_137)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_137),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_112),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_138),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_93),
.B(n_44),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_139),
.B(n_102),
.Y(n_158)
);

AOI21xp5_ASAP7_75t_L g140 ( 
.A1(n_109),
.A2(n_91),
.B(n_83),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_97),
.A2(n_91),
.B1(n_37),
.B2(n_35),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_141),
.A2(n_117),
.B1(n_103),
.B2(n_111),
.Y(n_154)
);

INVx8_ASAP7_75t_L g143 ( 
.A(n_107),
.Y(n_143)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_143),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_130),
.B(n_138),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_SL g177 ( 
.A(n_145),
.B(n_160),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g147 ( 
.A(n_140),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_147),
.B(n_151),
.Y(n_175)
);

NOR2x1_ASAP7_75t_L g148 ( 
.A(n_127),
.B(n_110),
.Y(n_148)
);

OR2x2_ASAP7_75t_L g181 ( 
.A(n_148),
.B(n_129),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_149),
.B(n_161),
.C(n_169),
.Y(n_178)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_143),
.Y(n_151)
);

CKINVDCx14_ASAP7_75t_R g174 ( 
.A(n_154),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_L g155 ( 
.A1(n_126),
.A2(n_110),
.B(n_101),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_155),
.B(n_156),
.Y(n_182)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_134),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_157),
.B(n_164),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_158),
.B(n_139),
.Y(n_184)
);

BUFx12_ASAP7_75t_L g159 ( 
.A(n_118),
.Y(n_159)
);

INVx13_ASAP7_75t_L g193 ( 
.A(n_159),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_131),
.B(n_114),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_128),
.B(n_108),
.C(n_37),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_163),
.A2(n_166),
.B1(n_141),
.B2(n_133),
.Y(n_176)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_122),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_121),
.A2(n_107),
.B1(n_35),
.B2(n_34),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_132),
.B(n_83),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_168),
.B(n_2),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_124),
.B(n_119),
.Y(n_169)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_158),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_171),
.B(n_172),
.Y(n_215)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_152),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_153),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_173),
.B(n_179),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_176),
.A2(n_180),
.B1(n_144),
.B2(n_166),
.Y(n_196)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_153),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_147),
.A2(n_146),
.B1(n_148),
.B2(n_162),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_L g212 ( 
.A1(n_181),
.A2(n_183),
.B(n_190),
.Y(n_212)
);

AND2x2_ASAP7_75t_L g183 ( 
.A(n_165),
.B(n_136),
.Y(n_183)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_184),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_150),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_185),
.Y(n_197)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_154),
.Y(n_187)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_187),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_144),
.A2(n_142),
.B1(n_135),
.B2(n_125),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_188),
.A2(n_174),
.B1(n_176),
.B2(n_180),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_149),
.B(n_125),
.C(n_123),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_189),
.B(n_191),
.C(n_167),
.Y(n_195)
);

AND2x2_ASAP7_75t_L g190 ( 
.A(n_167),
.B(n_123),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_169),
.B(n_35),
.C(n_83),
.Y(n_191)
);

A2O1A1O1Ixp25_ASAP7_75t_L g192 ( 
.A1(n_161),
.A2(n_22),
.B(n_3),
.C(n_4),
.D(n_5),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_192),
.B(n_2),
.Y(n_206)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_194),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_195),
.B(n_207),
.Y(n_231)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_196),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_187),
.A2(n_170),
.B1(n_155),
.B2(n_157),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_198),
.A2(n_211),
.B1(n_213),
.B2(n_172),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_178),
.B(n_156),
.C(n_159),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_200),
.B(n_191),
.C(n_182),
.Y(n_219)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_186),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_202),
.B(n_203),
.Y(n_228)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_183),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_205),
.B(n_209),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_206),
.B(n_208),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_178),
.B(n_159),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_183),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_177),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_184),
.Y(n_210)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_210),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_188),
.A2(n_181),
.B1(n_179),
.B2(n_171),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_189),
.A2(n_170),
.B1(n_150),
.B2(n_6),
.Y(n_213)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_216),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_219),
.B(n_215),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_200),
.B(n_182),
.C(n_190),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_220),
.B(n_224),
.Y(n_236)
);

AOI21xp5_ASAP7_75t_L g223 ( 
.A1(n_212),
.A2(n_175),
.B(n_190),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_223),
.B(n_227),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_207),
.B(n_193),
.C(n_192),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_195),
.B(n_193),
.C(n_3),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_225),
.B(n_226),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_211),
.B(n_2),
.C(n_6),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_SL g227 ( 
.A(n_201),
.B(n_7),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_213),
.B(n_7),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_229),
.B(n_230),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_SL g230 ( 
.A(n_215),
.B(n_8),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_217),
.A2(n_205),
.B1(n_199),
.B2(n_214),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_232),
.A2(n_237),
.B1(n_240),
.B2(n_8),
.Y(n_249)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_228),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_235),
.B(n_242),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_222),
.A2(n_198),
.B1(n_197),
.B2(n_212),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_238),
.B(n_219),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_218),
.A2(n_204),
.B1(n_206),
.B2(n_10),
.Y(n_240)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_226),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_225),
.B(n_204),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_243),
.B(n_224),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_244),
.B(n_250),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_245),
.B(n_238),
.Y(n_259)
);

OAI21xp5_ASAP7_75t_SL g247 ( 
.A1(n_236),
.A2(n_221),
.B(n_220),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_SL g260 ( 
.A1(n_247),
.A2(n_251),
.B(n_233),
.Y(n_260)
);

NAND3xp33_ASAP7_75t_L g248 ( 
.A(n_240),
.B(n_231),
.C(n_9),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_SL g257 ( 
.A(n_248),
.B(n_249),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_242),
.B(n_231),
.Y(n_250)
);

NOR2x1_ASAP7_75t_SL g251 ( 
.A(n_239),
.B(n_8),
.Y(n_251)
);

AO21x1_ASAP7_75t_L g252 ( 
.A1(n_234),
.A2(n_9),
.B(n_10),
.Y(n_252)
);

AOI21xp5_ASAP7_75t_L g255 ( 
.A1(n_252),
.A2(n_10),
.B(n_11),
.Y(n_255)
);

INVxp67_ASAP7_75t_L g253 ( 
.A(n_237),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_253),
.B(n_232),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_255),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_256),
.B(n_258),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_253),
.B(n_241),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_259),
.B(n_246),
.Y(n_263)
);

OAI21xp5_ASAP7_75t_SL g265 ( 
.A1(n_260),
.A2(n_11),
.B(n_12),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_263),
.B(n_265),
.Y(n_267)
);

OAI21x1_ASAP7_75t_L g264 ( 
.A1(n_254),
.A2(n_248),
.B(n_252),
.Y(n_264)
);

OAI211xp5_ASAP7_75t_L g266 ( 
.A1(n_264),
.A2(n_257),
.B(n_255),
.C(n_259),
.Y(n_266)
);

INVxp67_ASAP7_75t_L g269 ( 
.A(n_266),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_261),
.A2(n_11),
.B1(n_13),
.B2(n_14),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_SL g270 ( 
.A1(n_268),
.A2(n_262),
.B(n_15),
.Y(n_270)
);

HB1xp67_ASAP7_75t_L g271 ( 
.A(n_270),
.Y(n_271)
);

AOI21xp5_ASAP7_75t_L g272 ( 
.A1(n_271),
.A2(n_269),
.B(n_267),
.Y(n_272)
);

AOI21xp5_ASAP7_75t_L g273 ( 
.A1(n_272),
.A2(n_15),
.B(n_260),
.Y(n_273)
);


endmodule