module fake_jpeg_8708_n_275 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_275);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_275;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_272;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_122;
wire n_75;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_258;
wire n_96;

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_2),
.Y(n_19)
);

BUFx12_ASAP7_75t_L g20 ( 
.A(n_15),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_15),
.B(n_3),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_1),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_6),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

INVx13_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_12),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_10),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_18),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_SL g61 ( 
.A(n_36),
.B(n_20),
.Y(n_61)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_21),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_37),
.B(n_39),
.Y(n_69)
);

BUFx16f_ASAP7_75t_L g38 ( 
.A(n_21),
.Y(n_38)
);

INVx2_ASAP7_75t_SL g50 ( 
.A(n_38),
.Y(n_50)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_21),
.Y(n_39)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_26),
.Y(n_40)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_40),
.Y(n_65)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_18),
.Y(n_41)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_41),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_18),
.Y(n_42)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_23),
.Y(n_43)
);

AND2x2_ASAP7_75t_L g47 ( 
.A(n_43),
.B(n_29),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_18),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_44),
.Y(n_70)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_18),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_45),
.Y(n_67)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_38),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_46),
.B(n_49),
.Y(n_72)
);

NAND3xp33_ASAP7_75t_L g77 ( 
.A(n_47),
.B(n_0),
.C(n_2),
.Y(n_77)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_38),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_48),
.B(n_55),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_36),
.B(n_28),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g51 ( 
.A1(n_43),
.A2(n_29),
.B1(n_19),
.B2(n_24),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_51),
.A2(n_57),
.B1(n_59),
.B2(n_60),
.Y(n_86)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_52),
.B(n_54),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_42),
.B(n_28),
.Y(n_54)
);

INVx2_ASAP7_75t_SL g55 ( 
.A(n_39),
.Y(n_55)
);

OA22x2_ASAP7_75t_L g56 ( 
.A1(n_40),
.A2(n_35),
.B1(n_19),
.B2(n_31),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_L g95 ( 
.A1(n_56),
.A2(n_30),
.B1(n_17),
.B2(n_34),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g57 ( 
.A1(n_37),
.A2(n_29),
.B1(n_33),
.B2(n_32),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_58),
.B(n_61),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_45),
.A2(n_27),
.B1(n_22),
.B2(n_33),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g60 ( 
.A1(n_44),
.A2(n_32),
.B1(n_27),
.B2(n_22),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_45),
.A2(n_35),
.B1(n_24),
.B2(n_31),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_62),
.A2(n_64),
.B1(n_34),
.B2(n_30),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_44),
.A2(n_25),
.B1(n_23),
.B2(n_26),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_41),
.B(n_25),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_66),
.B(n_26),
.Y(n_74)
);

INVx5_ASAP7_75t_L g68 ( 
.A(n_41),
.Y(n_68)
);

INVx5_ASAP7_75t_L g75 ( 
.A(n_68),
.Y(n_75)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_65),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_71),
.B(n_73),
.Y(n_132)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_65),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_74),
.B(n_84),
.Y(n_129)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_70),
.Y(n_76)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_76),
.Y(n_110)
);

NOR2x1_ASAP7_75t_L g108 ( 
.A(n_77),
.B(n_99),
.Y(n_108)
);

AOI21xp5_ASAP7_75t_L g78 ( 
.A1(n_49),
.A2(n_20),
.B(n_28),
.Y(n_78)
);

OAI21xp5_ASAP7_75t_L g128 ( 
.A1(n_78),
.A2(n_91),
.B(n_0),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_53),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_80),
.B(n_87),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_54),
.B(n_45),
.C(n_41),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_81),
.B(n_105),
.Y(n_112)
);

BUFx2_ASAP7_75t_L g82 ( 
.A(n_70),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_82),
.Y(n_109)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_63),
.Y(n_83)
);

INVx2_ASAP7_75t_SL g106 ( 
.A(n_83),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g84 ( 
.A(n_69),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_53),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_61),
.Y(n_88)
);

INVx13_ASAP7_75t_L g124 ( 
.A(n_88),
.Y(n_124)
);

INVx13_ASAP7_75t_L g89 ( 
.A(n_50),
.Y(n_89)
);

INVx13_ASAP7_75t_L g127 ( 
.A(n_89),
.Y(n_127)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_47),
.B(n_45),
.Y(n_91)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_60),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_92),
.B(n_93),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_57),
.Y(n_93)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_68),
.Y(n_94)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_94),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_95),
.A2(n_102),
.B1(n_17),
.B2(n_52),
.Y(n_120)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_58),
.Y(n_96)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_96),
.Y(n_126)
);

BUFx12f_ASAP7_75t_L g97 ( 
.A(n_50),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_97),
.Y(n_130)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_56),
.Y(n_98)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_98),
.Y(n_114)
);

NOR2x1_ASAP7_75t_L g99 ( 
.A(n_47),
.B(n_41),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_100),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_48),
.B(n_20),
.Y(n_101)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_101),
.Y(n_116)
);

OAI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_56),
.A2(n_55),
.B1(n_30),
.B2(n_17),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_55),
.B(n_20),
.Y(n_103)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_103),
.Y(n_119)
);

BUFx8_ASAP7_75t_L g104 ( 
.A(n_50),
.Y(n_104)
);

BUFx4f_ASAP7_75t_SL g111 ( 
.A(n_104),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_67),
.B(n_28),
.Y(n_105)
);

AND2x6_ASAP7_75t_L g107 ( 
.A(n_99),
.B(n_56),
.Y(n_107)
);

NAND3xp33_ASAP7_75t_L g136 ( 
.A(n_107),
.B(n_91),
.C(n_86),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_72),
.B(n_67),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_113),
.B(n_117),
.Y(n_146)
);

A2O1A1Ixp33_ASAP7_75t_L g117 ( 
.A1(n_88),
.A2(n_63),
.B(n_34),
.C(n_28),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_120),
.B(n_82),
.Y(n_139)
);

BUFx8_ASAP7_75t_L g121 ( 
.A(n_104),
.Y(n_121)
);

INVx3_ASAP7_75t_L g147 ( 
.A(n_121),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_72),
.B(n_46),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_122),
.B(n_79),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_SL g154 ( 
.A1(n_128),
.A2(n_2),
.B(n_3),
.Y(n_154)
);

BUFx8_ASAP7_75t_L g131 ( 
.A(n_104),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_131),
.B(n_97),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_124),
.A2(n_75),
.B1(n_73),
.B2(n_71),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g181 ( 
.A(n_133),
.Y(n_181)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_132),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_134),
.B(n_137),
.Y(n_170)
);

AOI21xp5_ASAP7_75t_L g135 ( 
.A1(n_128),
.A2(n_98),
.B(n_91),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_L g163 ( 
.A1(n_135),
.A2(n_154),
.B(n_161),
.Y(n_163)
);

XOR2xp5_ASAP7_75t_SL g184 ( 
.A(n_136),
.B(n_150),
.Y(n_184)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_123),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_115),
.A2(n_81),
.B1(n_85),
.B2(n_90),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_138),
.A2(n_145),
.B1(n_160),
.B2(n_119),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_L g164 ( 
.A1(n_139),
.A2(n_156),
.B1(n_110),
.B2(n_127),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_126),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_140),
.B(n_141),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_106),
.B(n_85),
.Y(n_142)
);

CKINVDCx16_ASAP7_75t_R g165 ( 
.A(n_142),
.Y(n_165)
);

AND2x2_ASAP7_75t_L g143 ( 
.A(n_114),
.B(n_78),
.Y(n_143)
);

AOI21xp5_ASAP7_75t_L g162 ( 
.A1(n_143),
.A2(n_149),
.B(n_117),
.Y(n_162)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_113),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_144),
.B(n_151),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_115),
.A2(n_84),
.B1(n_76),
.B2(n_75),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_SL g167 ( 
.A(n_148),
.B(n_157),
.Y(n_167)
);

AND2x2_ASAP7_75t_L g149 ( 
.A(n_114),
.B(n_89),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_SL g150 ( 
.A(n_112),
.B(n_16),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_106),
.B(n_94),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_L g152 ( 
.A(n_112),
.B(n_122),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_152),
.B(n_153),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_106),
.B(n_83),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_125),
.B(n_96),
.Y(n_155)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_155),
.Y(n_168)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_129),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_126),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_118),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_SL g183 ( 
.A(n_158),
.B(n_111),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_118),
.B(n_97),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_159),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_107),
.A2(n_120),
.B1(n_108),
.B2(n_124),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_108),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_L g198 ( 
.A1(n_162),
.A2(n_166),
.B(n_172),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_164),
.A2(n_175),
.B1(n_187),
.B2(n_5),
.Y(n_203)
);

AOI21xp5_ASAP7_75t_L g166 ( 
.A1(n_143),
.A2(n_111),
.B(n_130),
.Y(n_166)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_155),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_169),
.B(n_173),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_L g172 ( 
.A1(n_135),
.A2(n_119),
.B(n_116),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_148),
.Y(n_173)
);

INVx1_ASAP7_75t_SL g174 ( 
.A(n_146),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_174),
.B(n_180),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_L g176 ( 
.A1(n_146),
.A2(n_116),
.B(n_109),
.Y(n_176)
);

AOI21xp5_ASAP7_75t_L g194 ( 
.A1(n_176),
.A2(n_180),
.B(n_186),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_160),
.A2(n_110),
.B1(n_127),
.B2(n_111),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_177),
.A2(n_134),
.B1(n_150),
.B2(n_156),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_149),
.Y(n_180)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_183),
.Y(n_191)
);

INVx1_ASAP7_75t_SL g185 ( 
.A(n_147),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_185),
.B(n_147),
.Y(n_190)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_149),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_186),
.B(n_157),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_138),
.A2(n_145),
.B1(n_144),
.B2(n_143),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g189 ( 
.A(n_187),
.B(n_152),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_189),
.B(n_208),
.C(n_163),
.Y(n_214)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_190),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_192),
.A2(n_196),
.B1(n_203),
.B2(n_163),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_170),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_193),
.B(n_199),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_L g224 ( 
.A1(n_194),
.A2(n_195),
.B(n_197),
.Y(n_224)
);

AOI21xp5_ASAP7_75t_L g195 ( 
.A1(n_181),
.A2(n_184),
.B(n_176),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_177),
.A2(n_137),
.B1(n_154),
.B2(n_161),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_SL g199 ( 
.A(n_165),
.B(n_16),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_185),
.B(n_14),
.Y(n_200)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_200),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_182),
.B(n_131),
.C(n_121),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_201),
.B(n_202),
.C(n_171),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_184),
.B(n_131),
.C(n_121),
.Y(n_202)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_179),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_204),
.B(n_205),
.Y(n_217)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_178),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_183),
.B(n_14),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_206),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_162),
.B(n_5),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_195),
.A2(n_181),
.B1(n_175),
.B2(n_166),
.Y(n_210)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_210),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_191),
.A2(n_174),
.B1(n_165),
.B2(n_169),
.Y(n_213)
);

INVxp67_ASAP7_75t_L g235 ( 
.A(n_213),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_214),
.B(n_216),
.C(n_218),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_189),
.B(n_172),
.C(n_173),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_198),
.B(n_168),
.C(n_167),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_219),
.B(n_6),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_198),
.B(n_168),
.C(n_167),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_220),
.B(n_221),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_197),
.B(n_194),
.C(n_202),
.Y(n_221)
);

AOI321xp33_ASAP7_75t_L g222 ( 
.A1(n_191),
.A2(n_192),
.A3(n_207),
.B1(n_188),
.B2(n_208),
.C(n_196),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_222),
.B(n_225),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_201),
.B(n_171),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_223),
.B(n_216),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_209),
.B(n_193),
.Y(n_227)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_227),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_211),
.B(n_205),
.Y(n_229)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_229),
.Y(n_246)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_217),
.Y(n_230)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_230),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_221),
.B(n_204),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_231),
.B(n_236),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_232),
.A2(n_212),
.B1(n_224),
.B2(n_225),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_215),
.B(n_7),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_233),
.A2(n_234),
.B1(n_7),
.B2(n_8),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_218),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_226),
.B(n_223),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_239),
.B(n_241),
.C(n_244),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_226),
.B(n_220),
.Y(n_241)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_242),
.Y(n_250)
);

HB1xp67_ASAP7_75t_L g243 ( 
.A(n_235),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_243),
.B(n_247),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_236),
.B(n_214),
.C(n_224),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_238),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_248),
.A2(n_235),
.B1(n_10),
.B2(n_11),
.Y(n_252)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_252),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_239),
.B(n_231),
.C(n_237),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_253),
.B(n_257),
.C(n_12),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_244),
.B(n_228),
.Y(n_254)
);

AND2x2_ASAP7_75t_L g262 ( 
.A(n_254),
.B(n_251),
.Y(n_262)
);

OAI21xp5_ASAP7_75t_L g256 ( 
.A1(n_245),
.A2(n_249),
.B(n_246),
.Y(n_256)
);

AOI21xp5_ASAP7_75t_SL g258 ( 
.A1(n_256),
.A2(n_240),
.B(n_9),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_241),
.B(n_228),
.Y(n_257)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_258),
.Y(n_265)
);

OAI21xp5_ASAP7_75t_SL g260 ( 
.A1(n_250),
.A2(n_240),
.B(n_9),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_260),
.B(n_262),
.Y(n_264)
);

OR2x2_ASAP7_75t_L g261 ( 
.A(n_255),
.B(n_12),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_261),
.B(n_263),
.Y(n_267)
);

BUFx2_ASAP7_75t_L g266 ( 
.A(n_259),
.Y(n_266)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_266),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_264),
.B(n_251),
.C(n_253),
.Y(n_268)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_268),
.Y(n_271)
);

AOI21xp5_ASAP7_75t_L g269 ( 
.A1(n_265),
.A2(n_254),
.B(n_257),
.Y(n_269)
);

OAI21x1_ASAP7_75t_SL g272 ( 
.A1(n_269),
.A2(n_267),
.B(n_270),
.Y(n_272)
);

HB1xp67_ASAP7_75t_L g273 ( 
.A(n_272),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_273),
.B(n_267),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_274),
.B(n_271),
.Y(n_275)
);


endmodule