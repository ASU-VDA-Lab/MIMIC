module fake_jpeg_26322_n_170 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_170);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_170;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx5_ASAP7_75t_L g47 ( 
.A(n_2),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_15),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_20),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_3),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_5),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_21),
.Y(n_52)
);

BUFx10_ASAP7_75t_L g53 ( 
.A(n_9),
.Y(n_53)
);

BUFx5_ASAP7_75t_L g54 ( 
.A(n_46),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_44),
.Y(n_55)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_13),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_1),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_37),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_27),
.Y(n_59)
);

INVx11_ASAP7_75t_L g60 ( 
.A(n_45),
.Y(n_60)
);

BUFx16f_ASAP7_75t_L g61 ( 
.A(n_7),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_34),
.Y(n_62)
);

BUFx12_ASAP7_75t_L g63 ( 
.A(n_35),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_1),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_12),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_38),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_36),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_18),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_40),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_8),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_10),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_14),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_50),
.B(n_0),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_73),
.B(n_74),
.Y(n_84)
);

CKINVDCx16_ASAP7_75t_R g74 ( 
.A(n_53),
.Y(n_74)
);

INVx8_ASAP7_75t_L g75 ( 
.A(n_49),
.Y(n_75)
);

INVx8_ASAP7_75t_L g91 ( 
.A(n_75),
.Y(n_91)
);

BUFx12f_ASAP7_75t_L g76 ( 
.A(n_49),
.Y(n_76)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_76),
.Y(n_89)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_49),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_77),
.Y(n_85)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_60),
.Y(n_78)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_78),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_60),
.Y(n_79)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_79),
.Y(n_86)
);

HAxp5_ASAP7_75t_SL g81 ( 
.A(n_76),
.B(n_64),
.CON(n_81),
.SN(n_81)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_81),
.B(n_83),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_75),
.A2(n_47),
.B1(n_56),
.B2(n_55),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_82),
.A2(n_90),
.B1(n_74),
.B2(n_53),
.Y(n_94)
);

INVx11_ASAP7_75t_L g83 ( 
.A(n_76),
.Y(n_83)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_77),
.Y(n_87)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_87),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_76),
.B(n_62),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_88),
.B(n_53),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_L g90 ( 
.A1(n_78),
.A2(n_47),
.B1(n_56),
.B2(n_67),
.Y(n_90)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_79),
.Y(n_92)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_92),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_94),
.A2(n_96),
.B1(n_65),
.B2(n_57),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_88),
.A2(n_72),
.B1(n_59),
.B2(n_48),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_97),
.B(n_98),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_80),
.B(n_68),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_85),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_99),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_80),
.B(n_68),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_100),
.B(n_102),
.Y(n_109)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_91),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_85),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_103),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_84),
.Y(n_104)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_104),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_86),
.B(n_67),
.Y(n_105)
);

XOR2xp5_ASAP7_75t_L g110 ( 
.A(n_105),
.B(n_92),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_81),
.B(n_71),
.Y(n_106)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_106),
.Y(n_115)
);

AOI32xp33_ASAP7_75t_L g108 ( 
.A1(n_95),
.A2(n_52),
.A3(n_58),
.B1(n_91),
.B2(n_63),
.Y(n_108)
);

A2O1A1O1Ixp25_ASAP7_75t_L g128 ( 
.A1(n_108),
.A2(n_54),
.B(n_61),
.C(n_51),
.D(n_25),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_110),
.B(n_119),
.Y(n_123)
);

AND2x2_ASAP7_75t_SL g111 ( 
.A(n_97),
.B(n_62),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_111),
.B(n_105),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_114),
.A2(n_70),
.B1(n_94),
.B2(n_83),
.Y(n_125)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_101),
.Y(n_116)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_116),
.Y(n_127)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_98),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_117),
.B(n_0),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_100),
.A2(n_86),
.B1(n_66),
.B2(n_69),
.Y(n_119)
);

OR2x2_ASAP7_75t_L g120 ( 
.A(n_109),
.B(n_96),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_120),
.B(n_124),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_112),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_121),
.B(n_122),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_113),
.B(n_93),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_125),
.A2(n_126),
.B1(n_129),
.B2(n_120),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_114),
.A2(n_89),
.B1(n_51),
.B2(n_63),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_126),
.A2(n_129),
.B1(n_2),
.B2(n_3),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_128),
.A2(n_22),
.B1(n_43),
.B2(n_42),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_107),
.A2(n_89),
.B1(n_61),
.B2(n_24),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_130),
.B(n_131),
.Y(n_139)
);

CKINVDCx16_ASAP7_75t_R g131 ( 
.A(n_111),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_123),
.A2(n_111),
.B1(n_118),
.B2(n_110),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_134),
.A2(n_137),
.B1(n_145),
.B2(n_7),
.Y(n_150)
);

AOI21x1_ASAP7_75t_SL g135 ( 
.A1(n_125),
.A2(n_115),
.B(n_23),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_L g147 ( 
.A1(n_135),
.A2(n_143),
.B(n_6),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_SL g154 ( 
.A(n_136),
.B(n_142),
.C(n_8),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_127),
.B(n_19),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_SL g149 ( 
.A(n_138),
.B(n_28),
.Y(n_149)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_122),
.Y(n_140)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_140),
.Y(n_146)
);

HB1xp67_ASAP7_75t_L g141 ( 
.A(n_128),
.Y(n_141)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_141),
.Y(n_151)
);

NAND2xp33_ASAP7_75t_SL g143 ( 
.A(n_131),
.B(n_4),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_121),
.Y(n_144)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_144),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_123),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_147),
.B(n_149),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_132),
.B(n_29),
.C(n_41),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_148),
.B(n_150),
.C(n_153),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_L g153 ( 
.A1(n_133),
.A2(n_30),
.B(n_39),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_154),
.B(n_155),
.C(n_139),
.Y(n_157)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_142),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_157),
.B(n_148),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_159),
.B(n_160),
.C(n_158),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_156),
.B(n_151),
.C(n_152),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_161),
.A2(n_147),
.B1(n_146),
.B2(n_135),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_162),
.B(n_143),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_163),
.B(n_9),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_164),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_165),
.B(n_11),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_SL g167 ( 
.A1(n_166),
.A2(n_16),
.B(n_17),
.Y(n_167)
);

AOI311xp33_ASAP7_75t_L g168 ( 
.A1(n_167),
.A2(n_26),
.A3(n_31),
.B(n_32),
.C(n_33),
.Y(n_168)
);

BUFx24_ASAP7_75t_SL g169 ( 
.A(n_168),
.Y(n_169)
);

BUFx24_ASAP7_75t_SL g170 ( 
.A(n_169),
.Y(n_170)
);


endmodule