module real_jpeg_18334_n_10 (n_5, n_4, n_8, n_0, n_1, n_2, n_6, n_7, n_3, n_9, n_10);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_2;
input n_6;
input n_7;
input n_3;
input n_9;

output n_10;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_176;
wire n_104;
wire n_153;
wire n_161;
wire n_64;
wire n_177;
wire n_11;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_140;
wire n_126;
wire n_13;
wire n_113;
wire n_155;
wire n_120;
wire n_93;
wire n_95;
wire n_141;
wire n_139;
wire n_33;
wire n_65;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_170;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_172;
wire n_45;
wire n_112;
wire n_42;
wire n_145;
wire n_18;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_100;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_30;
wire n_158;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_185;
wire n_55;
wire n_180;
wire n_58;
wire n_52;
wire n_63;
wire n_12;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_179;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_181;
wire n_85;
wire n_101;
wire n_182;
wire n_96;
wire n_89;
wire n_16;

BUFx3_ASAP7_75t_L g167 ( 
.A(n_0),
.Y(n_167)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_0),
.Y(n_175)
);

BUFx5_ASAP7_75t_L g60 ( 
.A(n_1),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_1),
.Y(n_71)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_1),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_1),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g21 ( 
.A1(n_2),
.A2(n_22),
.B1(n_25),
.B2(n_28),
.Y(n_21)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_2),
.A2(n_28),
.B1(n_179),
.B2(n_181),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_3),
.A2(n_51),
.B1(n_155),
.B2(n_156),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_3),
.Y(n_155)
);

BUFx3_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g142 ( 
.A(n_4),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g33 ( 
.A1(n_5),
.A2(n_34),
.B1(n_38),
.B2(n_39),
.Y(n_33)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_5),
.Y(n_38)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_6),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_6),
.Y(n_66)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_6),
.Y(n_82)
);

BUFx3_ASAP7_75t_L g102 ( 
.A(n_6),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_6),
.Y(n_111)
);

BUFx3_ASAP7_75t_L g169 ( 
.A(n_6),
.Y(n_169)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_7),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_7),
.A2(n_15),
.B1(n_126),
.B2(n_132),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_7),
.B(n_162),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_8),
.A2(n_104),
.B1(n_108),
.B2(n_109),
.Y(n_103)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_8),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_8),
.A2(n_108),
.B1(n_127),
.B2(n_129),
.Y(n_126)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

BUFx4f_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_9),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_9),
.Y(n_56)
);

XNOR2xp5_ASAP7_75t_L g10 ( 
.A(n_11),
.B(n_146),
.Y(n_10)
);

AOI21xp5_ASAP7_75t_L g11 ( 
.A1(n_12),
.A2(n_116),
.B(n_145),
.Y(n_11)
);

NAND2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_45),
.Y(n_12)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_13),
.B(n_45),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g13 ( 
.A1(n_14),
.A2(n_20),
.B1(n_29),
.B2(n_32),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_15),
.Y(n_14)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_15),
.A2(n_21),
.B1(n_126),
.B2(n_139),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_15),
.A2(n_33),
.B1(n_152),
.B2(n_153),
.Y(n_151)
);

OR2x2_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_18),
.Y(n_15)
);

BUFx3_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_17),
.Y(n_124)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

INVx5_ASAP7_75t_L g37 ( 
.A(n_19),
.Y(n_37)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_19),
.Y(n_76)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_19),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_24),
.Y(n_27)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_24),
.Y(n_131)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_31),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

HB1xp67_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_42),
.Y(n_88)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_43),
.Y(n_120)
);

INVx4_ASAP7_75t_L g159 ( 
.A(n_43),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g45 ( 
.A1(n_46),
.A2(n_77),
.B1(n_114),
.B2(n_115),
.Y(n_45)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_46),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_46),
.B(n_115),
.Y(n_149)
);

OAI32xp33_ASAP7_75t_L g46 ( 
.A1(n_47),
.A2(n_51),
.A3(n_57),
.B1(n_61),
.B2(n_67),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_50),
.Y(n_107)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

BUFx2_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g89 ( 
.A(n_56),
.Y(n_89)
);

BUFx2_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_60),
.Y(n_99)
);

OAI21xp33_ASAP7_75t_SL g78 ( 
.A1(n_61),
.A2(n_62),
.B(n_79),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_62),
.B(n_63),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g121 ( 
.A(n_62),
.B(n_122),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_62),
.B(n_113),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx6_ASAP7_75t_L g95 ( 
.A(n_66),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_68),
.B(n_72),
.Y(n_67)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_71),
.Y(n_98)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_77),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_78),
.A2(n_83),
.B1(n_103),
.B2(n_112),
.Y(n_77)
);

BUFx2_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

BUFx3_ASAP7_75t_L g171 ( 
.A(n_82),
.Y(n_171)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_82),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_83),
.A2(n_103),
.B1(n_112),
.B2(n_178),
.Y(n_177)
);

AND2x2_ASAP7_75t_SL g83 ( 
.A(n_84),
.B(n_92),
.Y(n_83)
);

BUFx2_ASAP7_75t_L g113 ( 
.A(n_84),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_85),
.A2(n_88),
.B1(n_89),
.B2(n_90),
.Y(n_84)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

BUFx3_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx6_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

OAI22xp33_ASAP7_75t_L g92 ( 
.A1(n_93),
.A2(n_96),
.B1(n_99),
.B2(n_100),
.Y(n_92)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx5_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx4_ASAP7_75t_L g180 ( 
.A(n_111),
.Y(n_180)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_L g116 ( 
.A1(n_117),
.A2(n_137),
.B(n_144),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_118),
.B(n_125),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_121),
.Y(n_118)
);

BUFx3_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx6_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx5_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

BUFx2_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

HB1xp67_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx4_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVx4_ASAP7_75t_SL g134 ( 
.A(n_135),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_143),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_138),
.B(n_143),
.Y(n_144)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_142),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_186),
.Y(n_146)
);

INVxp67_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

AND2x2_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_150),
.Y(n_148)
);

OR2x2_ASAP7_75t_L g186 ( 
.A(n_149),
.B(n_150),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_160),
.Y(n_150)
);

INVxp67_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_161),
.A2(n_176),
.B1(n_177),
.B2(n_185),
.Y(n_160)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_161),
.Y(n_185)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

BUFx2_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_165),
.A2(n_168),
.B1(n_170),
.B2(n_172),
.Y(n_164)
);

INVx3_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

INVx3_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

INVx4_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

BUFx2_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);


endmodule