module real_aes_8052_n_104 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_104);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_104;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_766;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_666;
wire n_537;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_310;
wire n_455;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_527;
wire n_434;
wire n_502;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_552;
wire n_402;
wire n_733;
wire n_602;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_768;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_756;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_765;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_456;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_762;
wire n_210;
wire n_212;
wire n_325;
wire n_575;
wire n_479;
wire n_338;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_687;
wire n_729;
wire n_646;
wire n_710;
wire n_650;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
NAND3xp33_ASAP7_75t_SL g112 ( .A(n_0), .B(n_88), .C(n_113), .Y(n_112) );
INVx1_ASAP7_75t_L g463 ( .A(n_0), .Y(n_463) );
INVx1_ASAP7_75t_L g514 ( .A(n_1), .Y(n_514) );
INVx1_ASAP7_75t_L g210 ( .A(n_2), .Y(n_210) );
AOI22xp5_ASAP7_75t_L g127 ( .A1(n_3), .A2(n_81), .B1(n_128), .B2(n_129), .Y(n_127) );
CKINVDCx20_ASAP7_75t_R g129 ( .A(n_3), .Y(n_129) );
AOI22xp33_ASAP7_75t_L g540 ( .A1(n_4), .A2(n_37), .B1(n_166), .B2(n_530), .Y(n_540) );
AOI21xp33_ASAP7_75t_L g190 ( .A1(n_5), .A2(n_147), .B(n_191), .Y(n_190) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_6), .B(n_140), .Y(n_505) );
AND2x6_ASAP7_75t_L g152 ( .A(n_7), .B(n_153), .Y(n_152) );
AOI21xp5_ASAP7_75t_L g248 ( .A1(n_8), .A2(n_249), .B(n_250), .Y(n_248) );
INVx1_ASAP7_75t_L g111 ( .A(n_9), .Y(n_111) );
NOR2xp33_ASAP7_75t_L g464 ( .A(n_9), .B(n_38), .Y(n_464) );
INVx1_ASAP7_75t_L g197 ( .A(n_10), .Y(n_197) );
NAND2xp5_ASAP7_75t_L g240 ( .A(n_11), .B(n_241), .Y(n_240) );
INVx1_ASAP7_75t_L g145 ( .A(n_12), .Y(n_145) );
INVx1_ASAP7_75t_L g509 ( .A(n_13), .Y(n_509) );
INVx1_ASAP7_75t_L g255 ( .A(n_14), .Y(n_255) );
NAND2xp5_ASAP7_75t_L g525 ( .A(n_15), .B(n_178), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g486 ( .A(n_16), .B(n_141), .Y(n_486) );
AO32x2_ASAP7_75t_L g538 ( .A1(n_17), .A2(n_140), .A3(n_175), .B1(n_492), .B2(n_539), .Y(n_538) );
NAND2xp5_ASAP7_75t_SL g528 ( .A(n_18), .B(n_166), .Y(n_528) );
NAND2xp5_ASAP7_75t_L g266 ( .A(n_19), .B(n_161), .Y(n_266) );
NAND2xp5_ASAP7_75t_L g516 ( .A(n_20), .B(n_141), .Y(n_516) );
AOI22xp33_ASAP7_75t_L g541 ( .A1(n_21), .A2(n_52), .B1(n_166), .B2(n_530), .Y(n_541) );
NAND2xp5_ASAP7_75t_SL g221 ( .A(n_22), .B(n_147), .Y(n_221) );
AOI22xp33_ASAP7_75t_SL g536 ( .A1(n_23), .A2(n_77), .B1(n_166), .B2(n_178), .Y(n_536) );
NAND2xp5_ASAP7_75t_SL g551 ( .A(n_24), .B(n_166), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g168 ( .A(n_25), .B(n_169), .Y(n_168) );
A2O1A1Ixp33_ASAP7_75t_L g252 ( .A1(n_26), .A2(n_253), .B(n_254), .C(n_256), .Y(n_252) );
BUFx6f_ASAP7_75t_L g151 ( .A(n_27), .Y(n_151) );
XNOR2xp5_ASAP7_75t_L g122 ( .A(n_28), .B(n_123), .Y(n_122) );
NAND2xp5_ASAP7_75t_L g574 ( .A(n_28), .B(n_199), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g212 ( .A(n_29), .B(n_195), .Y(n_212) );
OAI22xp5_ASAP7_75t_L g761 ( .A1(n_30), .A2(n_41), .B1(n_762), .B2(n_763), .Y(n_761) );
CKINVDCx20_ASAP7_75t_R g762 ( .A(n_30), .Y(n_762) );
INVx1_ASAP7_75t_L g184 ( .A(n_31), .Y(n_184) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_32), .B(n_199), .Y(n_553) );
INVx2_ASAP7_75t_L g150 ( .A(n_33), .Y(n_150) );
NAND2xp5_ASAP7_75t_SL g569 ( .A(n_34), .B(n_166), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_35), .B(n_199), .Y(n_531) );
A2O1A1Ixp33_ASAP7_75t_L g222 ( .A1(n_36), .A2(n_152), .B(n_156), .C(n_223), .Y(n_222) );
NAND2xp5_ASAP7_75t_L g110 ( .A(n_38), .B(n_111), .Y(n_110) );
INVx1_ASAP7_75t_L g182 ( .A(n_39), .Y(n_182) );
NAND2xp5_ASAP7_75t_SL g265 ( .A(n_40), .B(n_195), .Y(n_265) );
CKINVDCx14_ASAP7_75t_R g763 ( .A(n_41), .Y(n_763) );
AOI22xp5_ASAP7_75t_L g104 ( .A1(n_42), .A2(n_105), .B1(n_116), .B2(n_771), .Y(n_104) );
NAND2xp5_ASAP7_75t_SL g499 ( .A(n_43), .B(n_166), .Y(n_499) );
AOI222xp33_ASAP7_75t_L g469 ( .A1(n_44), .A2(n_470), .B1(n_756), .B2(n_757), .C1(n_766), .C2(n_768), .Y(n_469) );
OAI22xp5_ASAP7_75t_SL g760 ( .A1(n_45), .A2(n_761), .B1(n_764), .B2(n_765), .Y(n_760) );
CKINVDCx20_ASAP7_75t_R g765 ( .A(n_45), .Y(n_765) );
AOI22xp33_ASAP7_75t_L g535 ( .A1(n_46), .A2(n_89), .B1(n_228), .B2(n_530), .Y(n_535) );
NAND2xp5_ASAP7_75t_SL g502 ( .A(n_47), .B(n_166), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_48), .B(n_166), .Y(n_510) );
CKINVDCx16_ASAP7_75t_R g185 ( .A(n_49), .Y(n_185) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_50), .B(n_504), .Y(n_503) );
NAND2xp5_ASAP7_75t_L g243 ( .A(n_51), .B(n_147), .Y(n_243) );
AOI22xp33_ASAP7_75t_SL g491 ( .A1(n_53), .A2(n_62), .B1(n_166), .B2(n_178), .Y(n_491) );
AOI22xp5_ASAP7_75t_L g177 ( .A1(n_54), .A2(n_156), .B1(n_178), .B2(n_180), .Y(n_177) );
CKINVDCx20_ASAP7_75t_R g231 ( .A(n_55), .Y(n_231) );
NAND2xp5_ASAP7_75t_SL g524 ( .A(n_56), .B(n_166), .Y(n_524) );
CKINVDCx16_ASAP7_75t_R g207 ( .A(n_57), .Y(n_207) );
NAND2xp5_ASAP7_75t_SL g573 ( .A(n_58), .B(n_166), .Y(n_573) );
A2O1A1Ixp33_ASAP7_75t_L g193 ( .A1(n_59), .A2(n_165), .B(n_194), .C(n_196), .Y(n_193) );
CKINVDCx20_ASAP7_75t_R g269 ( .A(n_60), .Y(n_269) );
INVx1_ASAP7_75t_L g192 ( .A(n_61), .Y(n_192) );
INVx1_ASAP7_75t_L g153 ( .A(n_63), .Y(n_153) );
NAND2xp5_ASAP7_75t_L g515 ( .A(n_64), .B(n_166), .Y(n_515) );
INVx1_ASAP7_75t_L g144 ( .A(n_65), .Y(n_144) );
CKINVDCx20_ASAP7_75t_R g120 ( .A(n_66), .Y(n_120) );
AO32x2_ASAP7_75t_L g533 ( .A1(n_67), .A2(n_140), .A3(n_235), .B1(n_492), .B2(n_534), .Y(n_533) );
INVx1_ASAP7_75t_L g572 ( .A(n_68), .Y(n_572) );
INVx1_ASAP7_75t_L g548 ( .A(n_69), .Y(n_548) );
AOI22xp5_ASAP7_75t_L g757 ( .A1(n_70), .A2(n_758), .B1(n_759), .B2(n_760), .Y(n_757) );
CKINVDCx20_ASAP7_75t_R g758 ( .A(n_70), .Y(n_758) );
A2O1A1Ixp33_ASAP7_75t_SL g160 ( .A1(n_71), .A2(n_161), .B(n_162), .C(n_165), .Y(n_160) );
INVxp67_ASAP7_75t_L g163 ( .A(n_72), .Y(n_163) );
NAND2xp5_ASAP7_75t_SL g549 ( .A(n_73), .B(n_178), .Y(n_549) );
INVx1_ASAP7_75t_L g115 ( .A(n_74), .Y(n_115) );
CKINVDCx20_ASAP7_75t_R g188 ( .A(n_75), .Y(n_188) );
INVx1_ASAP7_75t_L g262 ( .A(n_76), .Y(n_262) );
NAND2xp5_ASAP7_75t_SL g465 ( .A(n_78), .B(n_466), .Y(n_465) );
A2O1A1Ixp33_ASAP7_75t_L g263 ( .A1(n_79), .A2(n_152), .B(n_156), .C(n_264), .Y(n_263) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_80), .B(n_530), .Y(n_529) );
CKINVDCx20_ASAP7_75t_R g128 ( .A(n_81), .Y(n_128) );
NAND2xp5_ASAP7_75t_SL g552 ( .A(n_82), .B(n_178), .Y(n_552) );
NAND2xp5_ASAP7_75t_SL g224 ( .A(n_83), .B(n_211), .Y(n_224) );
INVx2_ASAP7_75t_L g142 ( .A(n_84), .Y(n_142) );
NAND2xp5_ASAP7_75t_L g225 ( .A(n_85), .B(n_161), .Y(n_225) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_86), .B(n_178), .Y(n_500) );
A2O1A1Ixp33_ASAP7_75t_L g208 ( .A1(n_87), .A2(n_152), .B(n_156), .C(n_209), .Y(n_208) );
OR2x2_ASAP7_75t_L g460 ( .A(n_88), .B(n_461), .Y(n_460) );
OR2x2_ASAP7_75t_L g473 ( .A(n_88), .B(n_462), .Y(n_473) );
INVx2_ASAP7_75t_L g477 ( .A(n_88), .Y(n_477) );
AOI22xp33_ASAP7_75t_L g489 ( .A1(n_90), .A2(n_103), .B1(n_178), .B2(n_179), .Y(n_489) );
NAND2xp5_ASAP7_75t_L g198 ( .A(n_91), .B(n_199), .Y(n_198) );
CKINVDCx20_ASAP7_75t_R g215 ( .A(n_92), .Y(n_215) );
A2O1A1Ixp33_ASAP7_75t_L g237 ( .A1(n_93), .A2(n_152), .B(n_156), .C(n_238), .Y(n_237) );
CKINVDCx20_ASAP7_75t_R g245 ( .A(n_94), .Y(n_245) );
INVx1_ASAP7_75t_L g159 ( .A(n_95), .Y(n_159) );
CKINVDCx16_ASAP7_75t_R g251 ( .A(n_96), .Y(n_251) );
NAND2xp5_ASAP7_75t_SL g239 ( .A(n_97), .B(n_211), .Y(n_239) );
NAND2xp5_ASAP7_75t_L g570 ( .A(n_98), .B(n_178), .Y(n_570) );
NAND2xp5_ASAP7_75t_L g257 ( .A(n_99), .B(n_140), .Y(n_257) );
NAND2xp5_ASAP7_75t_L g114 ( .A(n_100), .B(n_115), .Y(n_114) );
AOI21xp5_ASAP7_75t_L g146 ( .A1(n_101), .A2(n_147), .B(n_154), .Y(n_146) );
OAI22xp5_ASAP7_75t_SL g125 ( .A1(n_102), .A2(n_126), .B1(n_127), .B2(n_130), .Y(n_125) );
CKINVDCx20_ASAP7_75t_R g130 ( .A(n_102), .Y(n_130) );
CKINVDCx20_ASAP7_75t_R g105 ( .A(n_106), .Y(n_105) );
CKINVDCx20_ASAP7_75t_R g106 ( .A(n_107), .Y(n_106) );
CKINVDCx9p33_ASAP7_75t_R g107 ( .A(n_108), .Y(n_107) );
CKINVDCx6p67_ASAP7_75t_R g772 ( .A(n_108), .Y(n_772) );
CKINVDCx9p33_ASAP7_75t_R g108 ( .A(n_109), .Y(n_108) );
NOR2xp33_ASAP7_75t_L g109 ( .A(n_110), .B(n_112), .Y(n_109) );
INVx1_ASAP7_75t_SL g113 ( .A(n_114), .Y(n_113) );
OA21x2_ASAP7_75t_L g116 ( .A1(n_117), .A2(n_121), .B(n_468), .Y(n_116) );
NAND3xp33_ASAP7_75t_L g468 ( .A(n_117), .B(n_465), .C(n_469), .Y(n_468) );
INVx2_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
INVx2_ASAP7_75t_SL g118 ( .A(n_119), .Y(n_118) );
INVx2_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
OAI21xp5_ASAP7_75t_L g121 ( .A1(n_122), .A2(n_457), .B(n_465), .Y(n_121) );
OAI22xp5_ASAP7_75t_L g123 ( .A1(n_124), .A2(n_125), .B1(n_131), .B2(n_132), .Y(n_123) );
CKINVDCx20_ASAP7_75t_R g124 ( .A(n_125), .Y(n_124) );
CKINVDCx20_ASAP7_75t_R g126 ( .A(n_127), .Y(n_126) );
OAI22x1_ASAP7_75t_SL g766 ( .A1(n_131), .A2(n_476), .B1(n_479), .B2(n_767), .Y(n_766) );
INVx1_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
OAI22xp5_ASAP7_75t_L g470 ( .A1(n_132), .A2(n_471), .B1(n_474), .B2(n_478), .Y(n_470) );
AND2x2_ASAP7_75t_SL g132 ( .A(n_133), .B(n_394), .Y(n_132) );
NOR4xp25_ASAP7_75t_L g133 ( .A(n_134), .B(n_324), .C(n_355), .D(n_374), .Y(n_133) );
NAND4xp25_ASAP7_75t_L g134 ( .A(n_135), .B(n_282), .C(n_297), .D(n_315), .Y(n_134) );
AOI222xp33_ASAP7_75t_L g135 ( .A1(n_136), .A2(n_217), .B1(n_258), .B2(n_270), .C1(n_275), .C2(n_277), .Y(n_135) );
NAND2xp5_ASAP7_75t_L g136 ( .A(n_137), .B(n_200), .Y(n_136) );
INVx1_ASAP7_75t_L g338 ( .A(n_137), .Y(n_338) );
NAND2xp5_ASAP7_75t_L g137 ( .A(n_138), .B(n_171), .Y(n_137) );
AND2x2_ASAP7_75t_L g201 ( .A(n_138), .B(n_189), .Y(n_201) );
NAND2xp5_ASAP7_75t_L g367 ( .A(n_138), .B(n_204), .Y(n_367) );
INVx3_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
OR2x2_ASAP7_75t_L g274 ( .A(n_139), .B(n_173), .Y(n_274) );
AND2x2_ASAP7_75t_L g283 ( .A(n_139), .B(n_284), .Y(n_283) );
INVx1_ASAP7_75t_L g309 ( .A(n_139), .Y(n_309) );
AND2x2_ASAP7_75t_L g330 ( .A(n_139), .B(n_173), .Y(n_330) );
BUFx2_ASAP7_75t_L g353 ( .A(n_139), .Y(n_353) );
AND2x2_ASAP7_75t_L g377 ( .A(n_139), .B(n_174), .Y(n_377) );
AND2x2_ASAP7_75t_L g441 ( .A(n_139), .B(n_189), .Y(n_441) );
OA21x2_ASAP7_75t_L g139 ( .A1(n_140), .A2(n_146), .B(n_168), .Y(n_139) );
INVx4_ASAP7_75t_L g170 ( .A(n_140), .Y(n_170) );
OA21x2_ASAP7_75t_L g496 ( .A1(n_140), .A2(n_497), .B(n_505), .Y(n_496) );
BUFx6f_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
INVx1_ASAP7_75t_L g175 ( .A(n_141), .Y(n_175) );
AND2x2_ASAP7_75t_L g141 ( .A(n_142), .B(n_143), .Y(n_141) );
AND2x2_ASAP7_75t_SL g199 ( .A(n_142), .B(n_143), .Y(n_199) );
NAND2xp5_ASAP7_75t_L g143 ( .A(n_144), .B(n_145), .Y(n_143) );
BUFx2_ASAP7_75t_L g249 ( .A(n_147), .Y(n_249) );
AND2x4_ASAP7_75t_L g147 ( .A(n_148), .B(n_152), .Y(n_147) );
NAND2x1p5_ASAP7_75t_L g186 ( .A(n_148), .B(n_152), .Y(n_186) );
AND2x2_ASAP7_75t_L g148 ( .A(n_149), .B(n_151), .Y(n_148) );
INVx1_ASAP7_75t_L g504 ( .A(n_149), .Y(n_504) );
INVx1_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
INVx2_ASAP7_75t_L g157 ( .A(n_150), .Y(n_157) );
INVx1_ASAP7_75t_L g179 ( .A(n_150), .Y(n_179) );
INVx1_ASAP7_75t_L g158 ( .A(n_151), .Y(n_158) );
INVx1_ASAP7_75t_L g161 ( .A(n_151), .Y(n_161) );
INVx3_ASAP7_75t_L g164 ( .A(n_151), .Y(n_164) );
BUFx6f_ASAP7_75t_L g181 ( .A(n_151), .Y(n_181) );
BUFx6f_ASAP7_75t_L g195 ( .A(n_151), .Y(n_195) );
INVx4_ASAP7_75t_SL g167 ( .A(n_152), .Y(n_167) );
BUFx3_ASAP7_75t_L g492 ( .A(n_152), .Y(n_492) );
OAI21xp5_ASAP7_75t_L g497 ( .A1(n_152), .A2(n_498), .B(n_501), .Y(n_497) );
OAI21xp5_ASAP7_75t_L g507 ( .A1(n_152), .A2(n_508), .B(n_512), .Y(n_507) );
OAI21xp5_ASAP7_75t_L g522 ( .A1(n_152), .A2(n_523), .B(n_527), .Y(n_522) );
OAI21xp5_ASAP7_75t_L g546 ( .A1(n_152), .A2(n_547), .B(n_550), .Y(n_546) );
O2A1O1Ixp33_ASAP7_75t_L g154 ( .A1(n_155), .A2(n_159), .B(n_160), .C(n_167), .Y(n_154) );
O2A1O1Ixp33_ASAP7_75t_L g191 ( .A1(n_155), .A2(n_167), .B(n_192), .C(n_193), .Y(n_191) );
O2A1O1Ixp33_ASAP7_75t_L g250 ( .A1(n_155), .A2(n_167), .B(n_251), .C(n_252), .Y(n_250) );
INVx5_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
AND2x6_ASAP7_75t_L g156 ( .A(n_157), .B(n_158), .Y(n_156) );
BUFx6f_ASAP7_75t_L g166 ( .A(n_157), .Y(n_166) );
BUFx3_ASAP7_75t_L g228 ( .A(n_157), .Y(n_228) );
INVx1_ASAP7_75t_L g530 ( .A(n_157), .Y(n_530) );
INVx1_ASAP7_75t_L g526 ( .A(n_161), .Y(n_526) );
NOR2xp33_ASAP7_75t_L g162 ( .A(n_163), .B(n_164), .Y(n_162) );
NOR2xp33_ASAP7_75t_L g196 ( .A(n_164), .B(n_197), .Y(n_196) );
INVx5_ASAP7_75t_L g211 ( .A(n_164), .Y(n_211) );
OAI22xp5_ASAP7_75t_SL g534 ( .A1(n_164), .A2(n_195), .B1(n_535), .B2(n_536), .Y(n_534) );
O2A1O1Ixp5_ASAP7_75t_SL g547 ( .A1(n_165), .A2(n_211), .B(n_548), .C(n_549), .Y(n_547) );
INVx3_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
HB1xp67_ASAP7_75t_L g242 ( .A(n_166), .Y(n_242) );
OAI22xp33_ASAP7_75t_L g176 ( .A1(n_167), .A2(n_177), .B1(n_185), .B2(n_186), .Y(n_176) );
OA21x2_ASAP7_75t_L g189 ( .A1(n_169), .A2(n_190), .B(n_198), .Y(n_189) );
INVx3_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
NOR2xp33_ASAP7_75t_SL g230 ( .A(n_170), .B(n_231), .Y(n_230) );
NAND3xp33_ASAP7_75t_L g487 ( .A(n_170), .B(n_488), .C(n_492), .Y(n_487) );
AO21x1_ASAP7_75t_L g580 ( .A1(n_170), .A2(n_488), .B(n_581), .Y(n_580) );
AND2x2_ASAP7_75t_L g342 ( .A(n_171), .B(n_273), .Y(n_342) );
INVx1_ASAP7_75t_L g171 ( .A(n_172), .Y(n_171) );
NOR2xp33_ASAP7_75t_L g366 ( .A(n_172), .B(n_367), .Y(n_366) );
OR2x2_ASAP7_75t_L g172 ( .A(n_173), .B(n_189), .Y(n_172) );
OR2x2_ASAP7_75t_L g302 ( .A(n_173), .B(n_205), .Y(n_302) );
AND2x2_ASAP7_75t_L g314 ( .A(n_173), .B(n_273), .Y(n_314) );
BUFx2_ASAP7_75t_L g446 ( .A(n_173), .Y(n_446) );
INVx3_ASAP7_75t_L g173 ( .A(n_174), .Y(n_173) );
OR2x2_ASAP7_75t_L g203 ( .A(n_174), .B(n_204), .Y(n_203) );
AND2x2_ASAP7_75t_L g296 ( .A(n_174), .B(n_205), .Y(n_296) );
AND2x2_ASAP7_75t_L g349 ( .A(n_174), .B(n_189), .Y(n_349) );
HB1xp67_ASAP7_75t_L g385 ( .A(n_174), .Y(n_385) );
AO21x2_ASAP7_75t_L g174 ( .A1(n_175), .A2(n_176), .B(n_187), .Y(n_174) );
NOR2xp33_ASAP7_75t_L g187 ( .A(n_175), .B(n_188), .Y(n_187) );
AO21x2_ASAP7_75t_L g205 ( .A1(n_175), .A2(n_206), .B(n_214), .Y(n_205) );
INVx2_ASAP7_75t_L g229 ( .A(n_175), .Y(n_229) );
INVx2_ASAP7_75t_L g213 ( .A(n_178), .Y(n_213) );
INVx3_ASAP7_75t_L g178 ( .A(n_179), .Y(n_178) );
OAI22xp5_ASAP7_75t_SL g180 ( .A1(n_181), .A2(n_182), .B1(n_183), .B2(n_184), .Y(n_180) );
INVx2_ASAP7_75t_L g183 ( .A(n_181), .Y(n_183) );
INVx4_ASAP7_75t_L g253 ( .A(n_181), .Y(n_253) );
OAI21xp5_ASAP7_75t_L g206 ( .A1(n_186), .A2(n_207), .B(n_208), .Y(n_206) );
OAI21xp5_ASAP7_75t_L g261 ( .A1(n_186), .A2(n_262), .B(n_263), .Y(n_261) );
AND2x2_ASAP7_75t_L g272 ( .A(n_189), .B(n_273), .Y(n_272) );
INVx1_ASAP7_75t_SL g284 ( .A(n_189), .Y(n_284) );
INVx2_ASAP7_75t_L g295 ( .A(n_189), .Y(n_295) );
BUFx2_ASAP7_75t_L g319 ( .A(n_189), .Y(n_319) );
AND2x2_ASAP7_75t_SL g376 ( .A(n_189), .B(n_377), .Y(n_376) );
AOI21xp5_ASAP7_75t_L g527 ( .A1(n_194), .A2(n_528), .B(n_529), .Y(n_527) );
O2A1O1Ixp5_ASAP7_75t_L g571 ( .A1(n_194), .A2(n_513), .B(n_572), .C(n_573), .Y(n_571) );
INVx2_ASAP7_75t_L g194 ( .A(n_195), .Y(n_194) );
INVx4_ASAP7_75t_L g241 ( .A(n_195), .Y(n_241) );
OAI22xp5_ASAP7_75t_L g488 ( .A1(n_195), .A2(n_489), .B1(n_490), .B2(n_491), .Y(n_488) );
OAI22xp5_ASAP7_75t_L g539 ( .A1(n_195), .A2(n_490), .B1(n_540), .B2(n_541), .Y(n_539) );
INVx1_ASAP7_75t_L g216 ( .A(n_199), .Y(n_216) );
INVx2_ASAP7_75t_L g235 ( .A(n_199), .Y(n_235) );
OA21x2_ASAP7_75t_L g247 ( .A1(n_199), .A2(n_248), .B(n_257), .Y(n_247) );
OA21x2_ASAP7_75t_L g521 ( .A1(n_199), .A2(n_522), .B(n_531), .Y(n_521) );
OA21x2_ASAP7_75t_L g545 ( .A1(n_199), .A2(n_546), .B(n_553), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g200 ( .A(n_201), .B(n_202), .Y(n_200) );
AOI332xp33_ASAP7_75t_L g297 ( .A1(n_201), .A2(n_298), .A3(n_302), .B1(n_303), .B2(n_307), .B3(n_310), .C1(n_311), .C2(n_313), .Y(n_297) );
NAND2x1_ASAP7_75t_L g382 ( .A(n_201), .B(n_273), .Y(n_382) );
NAND2xp5_ASAP7_75t_L g433 ( .A(n_201), .B(n_287), .Y(n_433) );
A2O1A1Ixp33_ASAP7_75t_SL g315 ( .A1(n_202), .A2(n_316), .B(n_319), .C(n_320), .Y(n_315) );
AND2x2_ASAP7_75t_L g454 ( .A(n_202), .B(n_295), .Y(n_454) );
INVx3_ASAP7_75t_SL g202 ( .A(n_203), .Y(n_202) );
OR2x2_ASAP7_75t_L g351 ( .A(n_203), .B(n_352), .Y(n_351) );
OR2x2_ASAP7_75t_L g356 ( .A(n_203), .B(n_353), .Y(n_356) );
INVx1_ASAP7_75t_L g287 ( .A(n_204), .Y(n_287) );
AND2x2_ASAP7_75t_L g390 ( .A(n_204), .B(n_349), .Y(n_390) );
AND2x2_ASAP7_75t_L g391 ( .A(n_204), .B(n_330), .Y(n_391) );
NAND2xp5_ASAP7_75t_L g400 ( .A(n_204), .B(n_401), .Y(n_400) );
NAND2xp5_ASAP7_75t_L g416 ( .A(n_204), .B(n_308), .Y(n_416) );
INVx3_ASAP7_75t_L g204 ( .A(n_205), .Y(n_204) );
INVx3_ASAP7_75t_L g273 ( .A(n_205), .Y(n_273) );
O2A1O1Ixp33_ASAP7_75t_L g209 ( .A1(n_210), .A2(n_211), .B(n_212), .C(n_213), .Y(n_209) );
INVx2_ASAP7_75t_L g490 ( .A(n_211), .Y(n_490) );
AOI21xp5_ASAP7_75t_L g498 ( .A1(n_211), .A2(n_499), .B(n_500), .Y(n_498) );
AOI21xp5_ASAP7_75t_L g568 ( .A1(n_211), .A2(n_569), .B(n_570), .Y(n_568) );
O2A1O1Ixp33_ASAP7_75t_L g508 ( .A1(n_213), .A2(n_509), .B(n_510), .C(n_511), .Y(n_508) );
NOR2xp33_ASAP7_75t_L g214 ( .A(n_215), .B(n_216), .Y(n_214) );
NOR2xp33_ASAP7_75t_L g244 ( .A(n_216), .B(n_245), .Y(n_244) );
NOR2xp33_ASAP7_75t_L g268 ( .A(n_216), .B(n_269), .Y(n_268) );
OAI31xp33_ASAP7_75t_L g455 ( .A1(n_217), .A2(n_376), .A3(n_383), .B(n_456), .Y(n_455) );
AND2x2_ASAP7_75t_L g217 ( .A(n_218), .B(n_232), .Y(n_217) );
AND2x2_ASAP7_75t_L g258 ( .A(n_218), .B(n_259), .Y(n_258) );
NAND2x1_ASAP7_75t_SL g278 ( .A(n_218), .B(n_279), .Y(n_278) );
HB1xp67_ASAP7_75t_L g365 ( .A(n_218), .Y(n_365) );
AND2x2_ASAP7_75t_L g370 ( .A(n_218), .B(n_281), .Y(n_370) );
INVx3_ASAP7_75t_L g218 ( .A(n_219), .Y(n_218) );
A2O1A1Ixp33_ASAP7_75t_L g282 ( .A1(n_219), .A2(n_283), .B(n_285), .C(n_288), .Y(n_282) );
OR2x2_ASAP7_75t_L g299 ( .A(n_219), .B(n_300), .Y(n_299) );
INVx1_ASAP7_75t_L g312 ( .A(n_219), .Y(n_312) );
AND2x2_ASAP7_75t_L g318 ( .A(n_219), .B(n_260), .Y(n_318) );
INVx2_ASAP7_75t_L g336 ( .A(n_219), .Y(n_336) );
AND2x2_ASAP7_75t_L g347 ( .A(n_219), .B(n_301), .Y(n_347) );
AND2x2_ASAP7_75t_L g379 ( .A(n_219), .B(n_337), .Y(n_379) );
AND2x2_ASAP7_75t_L g383 ( .A(n_219), .B(n_306), .Y(n_383) );
NAND2xp5_ASAP7_75t_L g388 ( .A(n_219), .B(n_232), .Y(n_388) );
AND2x2_ASAP7_75t_L g422 ( .A(n_219), .B(n_423), .Y(n_422) );
NOR2xp33_ASAP7_75t_L g456 ( .A(n_219), .B(n_325), .Y(n_456) );
OR2x6_ASAP7_75t_L g219 ( .A(n_220), .B(n_230), .Y(n_219) );
AOI21xp5_ASAP7_75t_SL g220 ( .A1(n_221), .A2(n_222), .B(n_229), .Y(n_220) );
AOI21xp5_ASAP7_75t_L g223 ( .A1(n_224), .A2(n_225), .B(n_226), .Y(n_223) );
AOI21xp5_ASAP7_75t_L g264 ( .A1(n_226), .A2(n_265), .B(n_266), .Y(n_264) );
INVx2_ASAP7_75t_L g226 ( .A(n_227), .Y(n_226) );
INVx2_ASAP7_75t_L g227 ( .A(n_228), .Y(n_227) );
INVx1_ASAP7_75t_L g256 ( .A(n_228), .Y(n_256) );
INVx1_ASAP7_75t_L g267 ( .A(n_229), .Y(n_267) );
OA21x2_ASAP7_75t_L g506 ( .A1(n_229), .A2(n_507), .B(n_516), .Y(n_506) );
OA21x2_ASAP7_75t_L g566 ( .A1(n_229), .A2(n_567), .B(n_574), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g286 ( .A(n_232), .B(n_287), .Y(n_286) );
INVx1_ASAP7_75t_L g364 ( .A(n_232), .Y(n_364) );
AND2x2_ASAP7_75t_L g426 ( .A(n_232), .B(n_347), .Y(n_426) );
AND2x2_ASAP7_75t_L g232 ( .A(n_233), .B(n_246), .Y(n_232) );
OR2x2_ASAP7_75t_L g280 ( .A(n_233), .B(n_281), .Y(n_280) );
AND2x2_ASAP7_75t_L g290 ( .A(n_233), .B(n_291), .Y(n_290) );
NAND2xp5_ASAP7_75t_L g300 ( .A(n_233), .B(n_301), .Y(n_300) );
INVx1_ASAP7_75t_L g398 ( .A(n_233), .Y(n_398) );
AND2x2_ASAP7_75t_L g415 ( .A(n_233), .B(n_260), .Y(n_415) );
INVx2_ASAP7_75t_L g233 ( .A(n_234), .Y(n_233) );
AND2x2_ASAP7_75t_L g306 ( .A(n_234), .B(n_246), .Y(n_306) );
AND2x2_ASAP7_75t_L g335 ( .A(n_234), .B(n_336), .Y(n_335) );
INVx1_ASAP7_75t_L g346 ( .A(n_234), .Y(n_346) );
NAND2xp5_ASAP7_75t_L g437 ( .A(n_234), .B(n_301), .Y(n_437) );
AO21x2_ASAP7_75t_L g234 ( .A1(n_235), .A2(n_236), .B(n_244), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g236 ( .A(n_237), .B(n_243), .Y(n_236) );
AOI21xp5_ASAP7_75t_L g238 ( .A1(n_239), .A2(n_240), .B(n_242), .Y(n_238) );
INVx1_ASAP7_75t_L g246 ( .A(n_247), .Y(n_246) );
AND2x2_ASAP7_75t_L g259 ( .A(n_247), .B(n_260), .Y(n_259) );
INVx2_ASAP7_75t_L g281 ( .A(n_247), .Y(n_281) );
AND2x2_ASAP7_75t_L g337 ( .A(n_247), .B(n_301), .Y(n_337) );
NOR2xp33_ASAP7_75t_L g254 ( .A(n_253), .B(n_255), .Y(n_254) );
INVx1_ASAP7_75t_L g511 ( .A(n_253), .Y(n_511) );
AOI21xp5_ASAP7_75t_L g550 ( .A1(n_253), .A2(n_551), .B(n_552), .Y(n_550) );
INVx1_ASAP7_75t_L g439 ( .A(n_258), .Y(n_439) );
INVx1_ASAP7_75t_L g443 ( .A(n_259), .Y(n_443) );
INVx2_ASAP7_75t_L g301 ( .A(n_260), .Y(n_301) );
AO21x2_ASAP7_75t_L g260 ( .A1(n_261), .A2(n_267), .B(n_268), .Y(n_260) );
NOR2xp33_ASAP7_75t_L g270 ( .A(n_271), .B(n_274), .Y(n_270) );
INVx1_ASAP7_75t_SL g271 ( .A(n_272), .Y(n_271) );
NAND2xp5_ASAP7_75t_L g417 ( .A(n_272), .B(n_418), .Y(n_417) );
NAND2xp5_ASAP7_75t_L g435 ( .A(n_272), .B(n_377), .Y(n_435) );
OR2x2_ASAP7_75t_L g276 ( .A(n_273), .B(n_274), .Y(n_276) );
INVx1_ASAP7_75t_SL g328 ( .A(n_273), .Y(n_328) );
INVx1_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
INVx1_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
AOI221xp5_ASAP7_75t_L g331 ( .A1(n_279), .A2(n_332), .B1(n_334), .B2(n_338), .C(n_339), .Y(n_331) );
INVx2_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
OR2x2_ASAP7_75t_L g359 ( .A(n_280), .B(n_323), .Y(n_359) );
INVx2_ASAP7_75t_L g291 ( .A(n_281), .Y(n_291) );
INVx1_ASAP7_75t_L g317 ( .A(n_281), .Y(n_317) );
NAND2xp5_ASAP7_75t_L g325 ( .A(n_281), .B(n_301), .Y(n_325) );
NAND2xp5_ASAP7_75t_L g411 ( .A(n_281), .B(n_304), .Y(n_411) );
INVx1_ASAP7_75t_L g419 ( .A(n_281), .Y(n_419) );
NAND2xp5_ASAP7_75t_L g333 ( .A(n_283), .B(n_287), .Y(n_333) );
AND2x4_ASAP7_75t_L g308 ( .A(n_284), .B(n_309), .Y(n_308) );
INVx1_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
AND2x2_ASAP7_75t_L g421 ( .A(n_287), .B(n_377), .Y(n_421) );
NOR2xp33_ASAP7_75t_L g288 ( .A(n_289), .B(n_292), .Y(n_288) );
INVx1_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
NAND2xp5_ASAP7_75t_L g321 ( .A(n_290), .B(n_322), .Y(n_321) );
INVxp67_ASAP7_75t_L g429 ( .A(n_291), .Y(n_429) );
INVxp67_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
AND2x2_ASAP7_75t_L g293 ( .A(n_294), .B(n_296), .Y(n_293) );
INVx1_ASAP7_75t_SL g294 ( .A(n_295), .Y(n_294) );
AND2x2_ASAP7_75t_L g329 ( .A(n_295), .B(n_330), .Y(n_329) );
AND2x2_ASAP7_75t_L g401 ( .A(n_295), .B(n_377), .Y(n_401) );
NAND2xp5_ASAP7_75t_L g407 ( .A(n_295), .B(n_314), .Y(n_407) );
AOI322xp5_ASAP7_75t_L g361 ( .A1(n_296), .A2(n_330), .A3(n_337), .B1(n_362), .B2(n_365), .C1(n_366), .C2(n_368), .Y(n_361) );
NAND2xp5_ASAP7_75t_L g404 ( .A(n_296), .B(n_405), .Y(n_404) );
INVx1_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
OR2x2_ASAP7_75t_L g427 ( .A(n_299), .B(n_428), .Y(n_427) );
INVx1_ASAP7_75t_L g373 ( .A(n_300), .Y(n_373) );
INVx2_ASAP7_75t_L g304 ( .A(n_301), .Y(n_304) );
INVx1_ASAP7_75t_L g363 ( .A(n_301), .Y(n_363) );
CKINVDCx16_ASAP7_75t_R g310 ( .A(n_302), .Y(n_310) );
NOR2xp33_ASAP7_75t_L g303 ( .A(n_304), .B(n_305), .Y(n_303) );
AND2x2_ASAP7_75t_L g399 ( .A(n_304), .B(n_312), .Y(n_399) );
INVx1_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
AND2x2_ASAP7_75t_L g311 ( .A(n_306), .B(n_312), .Y(n_311) );
AND2x2_ASAP7_75t_L g354 ( .A(n_306), .B(n_347), .Y(n_354) );
AND2x2_ASAP7_75t_L g358 ( .A(n_306), .B(n_318), .Y(n_358) );
OAI21xp33_ASAP7_75t_SL g368 ( .A1(n_307), .A2(n_369), .B(n_371), .Y(n_368) );
OAI22xp33_ASAP7_75t_L g438 ( .A1(n_307), .A2(n_439), .B1(n_440), .B2(n_442), .Y(n_438) );
INVx3_ASAP7_75t_SL g307 ( .A(n_308), .Y(n_307) );
AND2x2_ASAP7_75t_L g313 ( .A(n_308), .B(n_314), .Y(n_313) );
NAND2xp5_ASAP7_75t_L g340 ( .A(n_308), .B(n_328), .Y(n_340) );
NAND2xp5_ASAP7_75t_L g447 ( .A(n_310), .B(n_448), .Y(n_447) );
AND2x2_ASAP7_75t_L g316 ( .A(n_317), .B(n_318), .Y(n_316) );
INVx1_ASAP7_75t_L g450 ( .A(n_317), .Y(n_450) );
INVx4_ASAP7_75t_L g323 ( .A(n_318), .Y(n_323) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_318), .B(n_345), .Y(n_393) );
INVx1_ASAP7_75t_SL g405 ( .A(n_319), .Y(n_405) );
INVx1_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
INVx1_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
NOR2xp67_ASAP7_75t_L g418 ( .A(n_323), .B(n_419), .Y(n_418) );
OAI211xp5_ASAP7_75t_SL g324 ( .A1(n_325), .A2(n_326), .B(n_331), .C(n_348), .Y(n_324) );
OAI221xp5_ASAP7_75t_SL g444 ( .A1(n_326), .A2(n_364), .B1(n_443), .B2(n_445), .C(n_447), .Y(n_444) );
INVx1_ASAP7_75t_SL g326 ( .A(n_327), .Y(n_326) );
AND2x2_ASAP7_75t_L g327 ( .A(n_328), .B(n_329), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g440 ( .A(n_328), .B(n_441), .Y(n_440) );
OAI31xp33_ASAP7_75t_L g420 ( .A1(n_329), .A2(n_406), .A3(n_421), .B(n_422), .Y(n_420) );
INVx1_ASAP7_75t_L g360 ( .A(n_330), .Y(n_360) );
INVx1_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
AND2x2_ASAP7_75t_L g334 ( .A(n_335), .B(n_337), .Y(n_334) );
INVx1_ASAP7_75t_L g410 ( .A(n_335), .Y(n_410) );
AND2x2_ASAP7_75t_L g423 ( .A(n_337), .B(n_346), .Y(n_423) );
AOI21xp33_ASAP7_75t_L g339 ( .A1(n_340), .A2(n_341), .B(n_343), .Y(n_339) );
INVx1_ASAP7_75t_SL g341 ( .A(n_342), .Y(n_341) );
INVxp67_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
AND2x2_ASAP7_75t_L g344 ( .A(n_345), .B(n_347), .Y(n_344) );
INVx1_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
NAND2xp5_ASAP7_75t_L g449 ( .A(n_347), .B(n_450), .Y(n_449) );
OAI21xp33_ASAP7_75t_L g348 ( .A1(n_349), .A2(n_350), .B(n_354), .Y(n_348) );
INVx1_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
INVx1_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
OAI221xp5_ASAP7_75t_SL g355 ( .A1(n_356), .A2(n_357), .B1(n_359), .B2(n_360), .C(n_361), .Y(n_355) );
A2O1A1Ixp33_ASAP7_75t_L g424 ( .A1(n_356), .A2(n_425), .B(n_427), .C(n_430), .Y(n_424) );
CKINVDCx16_ASAP7_75t_R g357 ( .A(n_358), .Y(n_357) );
NAND2xp5_ASAP7_75t_SL g408 ( .A(n_359), .B(n_409), .Y(n_408) );
NOR2xp33_ASAP7_75t_L g362 ( .A(n_363), .B(n_364), .Y(n_362) );
INVx1_ASAP7_75t_L g386 ( .A(n_367), .Y(n_386) );
INVx1_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
AND2x2_ASAP7_75t_L g372 ( .A(n_370), .B(n_373), .Y(n_372) );
AND2x2_ASAP7_75t_L g414 ( .A(n_370), .B(n_415), .Y(n_414) );
INVx2_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
OAI211xp5_ASAP7_75t_L g374 ( .A1(n_375), .A2(n_378), .B(n_380), .C(n_389), .Y(n_374) );
INVx1_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
OAI221xp5_ASAP7_75t_L g451 ( .A1(n_378), .A2(n_388), .B1(n_452), .B2(n_453), .C(n_455), .Y(n_451) );
INVx1_ASAP7_75t_SL g378 ( .A(n_379), .Y(n_378) );
AOI22xp5_ASAP7_75t_L g380 ( .A1(n_381), .A2(n_383), .B1(n_384), .B2(n_387), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
AND2x2_ASAP7_75t_L g384 ( .A(n_385), .B(n_386), .Y(n_384) );
INVx1_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
OAI21xp5_ASAP7_75t_SL g389 ( .A1(n_390), .A2(n_391), .B(n_392), .Y(n_389) );
INVx1_ASAP7_75t_SL g452 ( .A(n_391), .Y(n_452) );
INVxp67_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
NOR4xp25_ASAP7_75t_L g394 ( .A(n_395), .B(n_424), .C(n_444), .D(n_451), .Y(n_394) );
OAI211xp5_ASAP7_75t_L g395 ( .A1(n_396), .A2(n_400), .B(n_402), .C(n_420), .Y(n_395) );
NAND2xp5_ASAP7_75t_L g396 ( .A(n_397), .B(n_399), .Y(n_396) );
INVxp67_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
O2A1O1Ixp33_ASAP7_75t_L g402 ( .A1(n_403), .A2(n_406), .B(n_408), .C(n_412), .Y(n_402) );
INVx1_ASAP7_75t_SL g403 ( .A(n_404), .Y(n_403) );
INVx1_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
INVx1_ASAP7_75t_SL g431 ( .A(n_409), .Y(n_431) );
OR2x2_ASAP7_75t_L g409 ( .A(n_410), .B(n_411), .Y(n_409) );
OR2x2_ASAP7_75t_L g442 ( .A(n_410), .B(n_443), .Y(n_442) );
OAI21xp33_ASAP7_75t_L g412 ( .A1(n_413), .A2(n_416), .B(n_417), .Y(n_412) );
INVx1_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
INVx1_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
HB1xp67_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
AOI221xp5_ASAP7_75t_L g430 ( .A1(n_431), .A2(n_432), .B1(n_434), .B2(n_436), .C(n_438), .Y(n_430) );
INVx1_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
INVx1_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
INVxp67_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
NAND2xp5_ASAP7_75t_L g445 ( .A(n_441), .B(n_446), .Y(n_445) );
INVx1_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
INVx1_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
INVx1_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
INVx1_ASAP7_75t_SL g458 ( .A(n_459), .Y(n_458) );
INVx1_ASAP7_75t_SL g459 ( .A(n_460), .Y(n_459) );
BUFx2_ASAP7_75t_L g467 ( .A(n_460), .Y(n_467) );
NOR2x2_ASAP7_75t_L g770 ( .A(n_461), .B(n_477), .Y(n_770) );
INVx2_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
OR2x2_ASAP7_75t_L g476 ( .A(n_462), .B(n_477), .Y(n_476) );
AND2x2_ASAP7_75t_L g462 ( .A(n_463), .B(n_464), .Y(n_462) );
INVx1_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
INVx2_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
INVx2_ASAP7_75t_L g767 ( .A(n_472), .Y(n_767) );
INVx1_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
INVx2_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
INVx1_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
INVx1_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
INVx2_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
AND2x2_ASAP7_75t_SL g480 ( .A(n_481), .B(n_690), .Y(n_480) );
NOR5xp2_ASAP7_75t_L g481 ( .A(n_482), .B(n_603), .C(n_649), .D(n_662), .E(n_674), .Y(n_481) );
OAI211xp5_ASAP7_75t_L g482 ( .A1(n_483), .A2(n_517), .B(n_557), .C(n_584), .Y(n_482) );
INVx1_ASAP7_75t_SL g685 ( .A(n_483), .Y(n_685) );
OR2x2_ASAP7_75t_L g483 ( .A(n_484), .B(n_493), .Y(n_483) );
AND2x2_ASAP7_75t_L g609 ( .A(n_484), .B(n_494), .Y(n_609) );
AND2x2_ASAP7_75t_L g637 ( .A(n_484), .B(n_583), .Y(n_637) );
AND2x2_ASAP7_75t_L g645 ( .A(n_484), .B(n_588), .Y(n_645) );
INVx3_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
AND2x2_ASAP7_75t_L g575 ( .A(n_485), .B(n_495), .Y(n_575) );
INVx2_ASAP7_75t_L g587 ( .A(n_485), .Y(n_587) );
AND2x2_ASAP7_75t_L g712 ( .A(n_485), .B(n_654), .Y(n_712) );
OR2x2_ASAP7_75t_L g714 ( .A(n_485), .B(n_715), .Y(n_714) );
AND2x4_ASAP7_75t_L g485 ( .A(n_486), .B(n_487), .Y(n_485) );
INVx1_ASAP7_75t_L g581 ( .A(n_486), .Y(n_581) );
AOI21xp5_ASAP7_75t_L g501 ( .A1(n_490), .A2(n_502), .B(n_503), .Y(n_501) );
O2A1O1Ixp33_ASAP7_75t_L g512 ( .A1(n_490), .A2(n_513), .B(n_514), .C(n_515), .Y(n_512) );
OAI21xp5_ASAP7_75t_L g567 ( .A1(n_492), .A2(n_568), .B(n_571), .Y(n_567) );
INVx2_ASAP7_75t_SL g493 ( .A(n_494), .Y(n_493) );
AND2x2_ASAP7_75t_L g625 ( .A(n_494), .B(n_597), .Y(n_625) );
NOR2xp33_ASAP7_75t_L g653 ( .A(n_494), .B(n_654), .Y(n_653) );
AND2x2_ASAP7_75t_L g739 ( .A(n_494), .B(n_579), .Y(n_739) );
AND2x2_ASAP7_75t_L g494 ( .A(n_495), .B(n_506), .Y(n_494) );
AND2x2_ASAP7_75t_L g582 ( .A(n_495), .B(n_583), .Y(n_582) );
INVx2_ASAP7_75t_L g629 ( .A(n_495), .Y(n_629) );
AND2x2_ASAP7_75t_L g654 ( .A(n_495), .B(n_566), .Y(n_654) );
NAND2xp5_ASAP7_75t_L g724 ( .A(n_495), .B(n_687), .Y(n_724) );
INVx3_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
AND2x2_ASAP7_75t_L g588 ( .A(n_496), .B(n_566), .Y(n_588) );
AND2x2_ASAP7_75t_L g602 ( .A(n_496), .B(n_565), .Y(n_602) );
AND2x2_ASAP7_75t_L g619 ( .A(n_496), .B(n_506), .Y(n_619) );
AND2x2_ASAP7_75t_L g676 ( .A(n_496), .B(n_677), .Y(n_676) );
NAND2xp5_ASAP7_75t_L g689 ( .A(n_496), .B(n_583), .Y(n_689) );
AND2x2_ASAP7_75t_L g741 ( .A(n_496), .B(n_666), .Y(n_741) );
INVx2_ASAP7_75t_L g513 ( .A(n_504), .Y(n_513) );
AND2x2_ASAP7_75t_L g564 ( .A(n_506), .B(n_565), .Y(n_564) );
INVx2_ASAP7_75t_L g583 ( .A(n_506), .Y(n_583) );
NAND2xp5_ASAP7_75t_L g660 ( .A(n_506), .B(n_566), .Y(n_660) );
AOI21xp5_ASAP7_75t_L g517 ( .A1(n_518), .A2(n_542), .B(n_554), .Y(n_517) );
INVx1_ASAP7_75t_SL g673 ( .A(n_518), .Y(n_673) );
AND2x4_ASAP7_75t_L g518 ( .A(n_519), .B(n_532), .Y(n_518) );
BUFx3_ASAP7_75t_L g519 ( .A(n_520), .Y(n_519) );
AND2x2_ASAP7_75t_SL g561 ( .A(n_520), .B(n_562), .Y(n_561) );
INVx1_ASAP7_75t_L g520 ( .A(n_521), .Y(n_520) );
INVx2_ASAP7_75t_L g556 ( .A(n_521), .Y(n_556) );
INVx1_ASAP7_75t_L g593 ( .A(n_521), .Y(n_593) );
AND2x2_ASAP7_75t_L g614 ( .A(n_521), .B(n_537), .Y(n_614) );
AND2x2_ASAP7_75t_L g648 ( .A(n_521), .B(n_538), .Y(n_648) );
OR2x2_ASAP7_75t_L g667 ( .A(n_521), .B(n_544), .Y(n_667) );
HB1xp67_ASAP7_75t_L g681 ( .A(n_521), .Y(n_681) );
AND2x2_ASAP7_75t_L g694 ( .A(n_521), .B(n_695), .Y(n_694) );
AOI21xp5_ASAP7_75t_L g523 ( .A1(n_524), .A2(n_525), .B(n_526), .Y(n_523) );
AOI22xp5_ASAP7_75t_L g615 ( .A1(n_532), .A2(n_616), .B1(n_617), .B2(n_626), .Y(n_615) );
AND2x2_ASAP7_75t_L g699 ( .A(n_532), .B(n_700), .Y(n_699) );
AND2x2_ASAP7_75t_L g532 ( .A(n_533), .B(n_537), .Y(n_532) );
INVx1_ASAP7_75t_L g560 ( .A(n_533), .Y(n_560) );
BUFx6f_ASAP7_75t_L g597 ( .A(n_533), .Y(n_597) );
INVx1_ASAP7_75t_L g608 ( .A(n_533), .Y(n_608) );
AND2x2_ASAP7_75t_L g623 ( .A(n_533), .B(n_538), .Y(n_623) );
OR2x2_ASAP7_75t_L g577 ( .A(n_537), .B(n_562), .Y(n_577) );
AND2x2_ASAP7_75t_L g607 ( .A(n_537), .B(n_608), .Y(n_607) );
NOR2xp67_ASAP7_75t_L g695 ( .A(n_537), .B(n_696), .Y(n_695) );
INVx2_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
AND2x2_ASAP7_75t_L g555 ( .A(n_538), .B(n_556), .Y(n_555) );
BUFx2_ASAP7_75t_L g664 ( .A(n_538), .Y(n_664) );
NAND2xp5_ASAP7_75t_L g679 ( .A(n_542), .B(n_680), .Y(n_679) );
BUFx2_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
AND2x2_ASAP7_75t_L g642 ( .A(n_543), .B(n_608), .Y(n_642) );
INVx2_ASAP7_75t_L g543 ( .A(n_544), .Y(n_543) );
AND2x2_ASAP7_75t_L g554 ( .A(n_544), .B(n_555), .Y(n_554) );
INVx1_ASAP7_75t_L g613 ( .A(n_544), .Y(n_613) );
INVx2_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
INVx2_ASAP7_75t_L g562 ( .A(n_545), .Y(n_562) );
OR2x2_ASAP7_75t_L g592 ( .A(n_545), .B(n_593), .Y(n_592) );
HB1xp67_ASAP7_75t_L g647 ( .A(n_545), .Y(n_647) );
AOI32xp33_ASAP7_75t_L g684 ( .A1(n_554), .A2(n_614), .A3(n_685), .B1(n_686), .B2(n_688), .Y(n_684) );
AND2x2_ASAP7_75t_L g610 ( .A(n_555), .B(n_611), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g708 ( .A(n_555), .B(n_709), .Y(n_708) );
NAND2xp5_ASAP7_75t_L g728 ( .A(n_555), .B(n_642), .Y(n_728) );
INVx1_ASAP7_75t_L g733 ( .A(n_555), .Y(n_733) );
AOI22xp5_ASAP7_75t_L g557 ( .A1(n_558), .A2(n_563), .B1(n_576), .B2(n_578), .Y(n_557) );
AND2x2_ASAP7_75t_L g558 ( .A(n_559), .B(n_561), .Y(n_558) );
AND2x2_ASAP7_75t_L g663 ( .A(n_559), .B(n_664), .Y(n_663) );
HB1xp67_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g707 ( .A(n_560), .B(n_562), .Y(n_707) );
AOI22xp5_ASAP7_75t_L g584 ( .A1(n_561), .A2(n_585), .B1(n_589), .B2(n_599), .Y(n_584) );
AND2x2_ASAP7_75t_L g606 ( .A(n_561), .B(n_607), .Y(n_606) );
A2O1A1Ixp33_ASAP7_75t_L g657 ( .A1(n_561), .A2(n_575), .B(n_623), .C(n_658), .Y(n_657) );
OAI332xp33_ASAP7_75t_L g662 ( .A1(n_561), .A2(n_663), .A3(n_665), .B1(n_667), .B2(n_668), .B3(n_670), .C1(n_671), .C2(n_673), .Y(n_662) );
INVx2_ASAP7_75t_L g703 ( .A(n_561), .Y(n_703) );
HB1xp67_ASAP7_75t_L g621 ( .A(n_562), .Y(n_621) );
INVx1_ASAP7_75t_L g696 ( .A(n_562), .Y(n_696) );
AND2x2_ASAP7_75t_L g750 ( .A(n_562), .B(n_614), .Y(n_750) );
AND2x2_ASAP7_75t_L g563 ( .A(n_564), .B(n_575), .Y(n_563) );
AND2x2_ASAP7_75t_L g630 ( .A(n_565), .B(n_580), .Y(n_630) );
INVx2_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
AND2x2_ASAP7_75t_L g579 ( .A(n_566), .B(n_580), .Y(n_579) );
OR2x2_ASAP7_75t_L g678 ( .A(n_566), .B(n_580), .Y(n_678) );
INVx1_ASAP7_75t_L g687 ( .A(n_566), .Y(n_687) );
INVx1_ASAP7_75t_L g661 ( .A(n_575), .Y(n_661) );
INVxp67_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
OR2x2_ASAP7_75t_L g745 ( .A(n_577), .B(n_597), .Y(n_745) );
INVx1_ASAP7_75t_SL g656 ( .A(n_578), .Y(n_656) );
AND2x2_ASAP7_75t_L g578 ( .A(n_579), .B(n_582), .Y(n_578) );
AND2x2_ASAP7_75t_L g683 ( .A(n_579), .B(n_641), .Y(n_683) );
INVx1_ASAP7_75t_L g702 ( .A(n_579), .Y(n_702) );
NAND2xp5_ASAP7_75t_SL g704 ( .A(n_579), .B(n_669), .Y(n_704) );
INVx1_ASAP7_75t_L g601 ( .A(n_580), .Y(n_601) );
AND2x2_ASAP7_75t_L g605 ( .A(n_582), .B(n_586), .Y(n_605) );
AND2x2_ASAP7_75t_L g672 ( .A(n_582), .B(n_630), .Y(n_672) );
INVx2_ASAP7_75t_L g715 ( .A(n_582), .Y(n_715) );
INVx2_ASAP7_75t_L g598 ( .A(n_583), .Y(n_598) );
AND2x2_ASAP7_75t_L g600 ( .A(n_583), .B(n_601), .Y(n_600) );
AND2x2_ASAP7_75t_L g585 ( .A(n_586), .B(n_588), .Y(n_585) );
INVx1_ASAP7_75t_L g616 ( .A(n_586), .Y(n_616) );
INVx2_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
NOR2xp33_ASAP7_75t_L g666 ( .A(n_587), .B(n_660), .Y(n_666) );
OR2x2_ASAP7_75t_L g730 ( .A(n_587), .B(n_689), .Y(n_730) );
INVx1_ASAP7_75t_L g754 ( .A(n_587), .Y(n_754) );
INVx1_ASAP7_75t_L g710 ( .A(n_588), .Y(n_710) );
AND2x2_ASAP7_75t_L g755 ( .A(n_588), .B(n_598), .Y(n_755) );
INVx1_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
NAND2xp5_ASAP7_75t_L g590 ( .A(n_591), .B(n_594), .Y(n_590) );
INVx2_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
OAI22xp5_ASAP7_75t_L g617 ( .A1(n_592), .A2(n_618), .B1(n_620), .B2(n_624), .Y(n_617) );
INVx1_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
OAI322xp33_ASAP7_75t_SL g701 ( .A1(n_595), .A2(n_702), .A3(n_703), .B1(n_704), .B2(n_705), .C1(n_708), .C2(n_710), .Y(n_701) );
OR2x2_ASAP7_75t_L g595 ( .A(n_596), .B(n_598), .Y(n_595) );
AND2x2_ASAP7_75t_L g698 ( .A(n_596), .B(n_614), .Y(n_698) );
OR2x2_ASAP7_75t_L g732 ( .A(n_596), .B(n_733), .Y(n_732) );
OR2x2_ASAP7_75t_L g735 ( .A(n_596), .B(n_667), .Y(n_735) );
INVx2_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
AND2x2_ASAP7_75t_L g680 ( .A(n_597), .B(n_681), .Y(n_680) );
OR2x2_ASAP7_75t_L g736 ( .A(n_597), .B(n_667), .Y(n_736) );
INVx3_ASAP7_75t_L g669 ( .A(n_598), .Y(n_669) );
AND2x2_ASAP7_75t_L g599 ( .A(n_600), .B(n_602), .Y(n_599) );
INVx1_ASAP7_75t_L g725 ( .A(n_600), .Y(n_725) );
AOI222xp33_ASAP7_75t_L g604 ( .A1(n_602), .A2(n_605), .B1(n_606), .B2(n_609), .C1(n_610), .C2(n_612), .Y(n_604) );
INVx1_ASAP7_75t_L g635 ( .A(n_602), .Y(n_635) );
NAND3xp33_ASAP7_75t_SL g603 ( .A(n_604), .B(n_615), .C(n_632), .Y(n_603) );
AND2x2_ASAP7_75t_L g720 ( .A(n_607), .B(n_621), .Y(n_720) );
BUFx2_ASAP7_75t_L g611 ( .A(n_608), .Y(n_611) );
INVx1_ASAP7_75t_L g652 ( .A(n_608), .Y(n_652) );
AOI221xp5_ASAP7_75t_L g697 ( .A1(n_609), .A2(n_645), .B1(n_698), .B2(n_699), .C(n_701), .Y(n_697) );
NAND2xp5_ASAP7_75t_L g693 ( .A(n_611), .B(n_694), .Y(n_693) );
AND2x2_ASAP7_75t_L g612 ( .A(n_613), .B(n_614), .Y(n_612) );
HB1xp67_ASAP7_75t_L g638 ( .A(n_614), .Y(n_638) );
AND2x2_ASAP7_75t_L g651 ( .A(n_614), .B(n_652), .Y(n_651) );
INVx1_ASAP7_75t_SL g618 ( .A(n_619), .Y(n_618) );
NAND2xp5_ASAP7_75t_L g631 ( .A(n_619), .B(n_630), .Y(n_631) );
OR2x2_ASAP7_75t_L g620 ( .A(n_621), .B(n_622), .Y(n_620) );
OAI21xp33_ASAP7_75t_L g626 ( .A1(n_621), .A2(n_627), .B(n_631), .Y(n_626) );
NAND2xp5_ASAP7_75t_L g650 ( .A(n_621), .B(n_651), .Y(n_650) );
INVx1_ASAP7_75t_SL g622 ( .A(n_623), .Y(n_622) );
AND2x2_ASAP7_75t_L g718 ( .A(n_623), .B(n_700), .Y(n_718) );
INVx1_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
INVx1_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
AND2x2_ASAP7_75t_L g628 ( .A(n_629), .B(n_630), .Y(n_628) );
INVx1_ASAP7_75t_L g641 ( .A(n_629), .Y(n_641) );
NAND2xp5_ASAP7_75t_L g640 ( .A(n_630), .B(n_641), .Y(n_640) );
INVx2_ASAP7_75t_L g747 ( .A(n_630), .Y(n_747) );
AOI221xp5_ASAP7_75t_L g632 ( .A1(n_633), .A2(n_638), .B1(n_639), .B2(n_642), .C(n_643), .Y(n_632) );
INVx2_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
NAND2xp5_ASAP7_75t_SL g722 ( .A(n_634), .B(n_723), .Y(n_722) );
OR2x2_ASAP7_75t_L g634 ( .A(n_635), .B(n_636), .Y(n_634) );
INVx1_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
INVx1_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
AND2x2_ASAP7_75t_L g743 ( .A(n_642), .B(n_648), .Y(n_743) );
INVxp67_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g644 ( .A(n_645), .B(n_646), .Y(n_644) );
OAI31xp33_ASAP7_75t_SL g711 ( .A1(n_646), .A2(n_685), .A3(n_712), .B(n_713), .Y(n_711) );
AND2x2_ASAP7_75t_L g646 ( .A(n_647), .B(n_648), .Y(n_646) );
INVx1_ASAP7_75t_L g700 ( .A(n_647), .Y(n_700) );
NAND2xp5_ASAP7_75t_SL g751 ( .A(n_648), .B(n_652), .Y(n_751) );
OAI221xp5_ASAP7_75t_SL g649 ( .A1(n_650), .A2(n_653), .B1(n_655), .B2(n_656), .C(n_657), .Y(n_649) );
INVx1_ASAP7_75t_L g655 ( .A(n_651), .Y(n_655) );
NAND2xp5_ASAP7_75t_L g668 ( .A(n_654), .B(n_669), .Y(n_668) );
INVx1_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
OR2x2_ASAP7_75t_L g659 ( .A(n_660), .B(n_661), .Y(n_659) );
INVx1_ASAP7_75t_L g670 ( .A(n_663), .Y(n_670) );
INVx2_ASAP7_75t_L g706 ( .A(n_664), .Y(n_706) );
INVx1_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
OR2x2_ASAP7_75t_L g692 ( .A(n_669), .B(n_678), .Y(n_692) );
A2O1A1Ixp33_ASAP7_75t_L g742 ( .A1(n_669), .A2(n_686), .B(n_743), .C(n_744), .Y(n_742) );
OAI221xp5_ASAP7_75t_SL g674 ( .A1(n_670), .A2(n_675), .B1(n_679), .B2(n_682), .C(n_684), .Y(n_674) );
INVx1_ASAP7_75t_SL g671 ( .A(n_672), .Y(n_671) );
A2O1A1Ixp33_ASAP7_75t_L g737 ( .A1(n_673), .A2(n_738), .B(n_740), .C(n_742), .Y(n_737) );
INVx1_ASAP7_75t_L g675 ( .A(n_676), .Y(n_675) );
AOI221xp5_ASAP7_75t_L g726 ( .A1(n_676), .A2(n_727), .B1(n_729), .B2(n_731), .C(n_734), .Y(n_726) );
INVx1_ASAP7_75t_SL g677 ( .A(n_678), .Y(n_677) );
INVx1_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
INVx1_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
INVx1_ASAP7_75t_SL g688 ( .A(n_689), .Y(n_688) );
NOR4xp25_ASAP7_75t_L g690 ( .A(n_691), .B(n_716), .C(n_737), .D(n_748), .Y(n_690) );
OAI211xp5_ASAP7_75t_SL g691 ( .A1(n_692), .A2(n_693), .B(n_697), .C(n_711), .Y(n_691) );
INVx1_ASAP7_75t_SL g746 ( .A(n_698), .Y(n_746) );
OR2x2_ASAP7_75t_L g705 ( .A(n_706), .B(n_707), .Y(n_705) );
INVx1_ASAP7_75t_SL g709 ( .A(n_707), .Y(n_709) );
INVx1_ASAP7_75t_L g713 ( .A(n_714), .Y(n_713) );
OAI22xp5_ASAP7_75t_L g734 ( .A1(n_714), .A2(n_723), .B1(n_735), .B2(n_736), .Y(n_734) );
A2O1A1Ixp33_ASAP7_75t_L g716 ( .A1(n_717), .A2(n_719), .B(n_721), .C(n_726), .Y(n_716) );
INVx1_ASAP7_75t_L g717 ( .A(n_718), .Y(n_717) );
AOI31xp33_ASAP7_75t_L g748 ( .A1(n_719), .A2(n_749), .A3(n_751), .B(n_752), .Y(n_748) );
INVx1_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
INVxp67_ASAP7_75t_L g721 ( .A(n_722), .Y(n_721) );
OR2x2_ASAP7_75t_L g723 ( .A(n_724), .B(n_725), .Y(n_723) );
INVx1_ASAP7_75t_L g727 ( .A(n_728), .Y(n_727) );
INVx1_ASAP7_75t_SL g729 ( .A(n_730), .Y(n_729) );
INVx1_ASAP7_75t_L g731 ( .A(n_732), .Y(n_731) );
INVx1_ASAP7_75t_L g738 ( .A(n_739), .Y(n_738) );
INVx1_ASAP7_75t_SL g740 ( .A(n_741), .Y(n_740) );
AOI21xp5_ASAP7_75t_L g744 ( .A1(n_745), .A2(n_746), .B(n_747), .Y(n_744) );
INVx1_ASAP7_75t_L g749 ( .A(n_750), .Y(n_749) );
NAND2xp5_ASAP7_75t_L g752 ( .A(n_753), .B(n_755), .Y(n_752) );
INVx1_ASAP7_75t_L g753 ( .A(n_754), .Y(n_753) );
CKINVDCx20_ASAP7_75t_R g756 ( .A(n_757), .Y(n_756) );
CKINVDCx14_ASAP7_75t_R g759 ( .A(n_760), .Y(n_759) );
INVx1_ASAP7_75t_L g764 ( .A(n_761), .Y(n_764) );
INVx1_ASAP7_75t_SL g768 ( .A(n_769), .Y(n_768) );
INVx3_ASAP7_75t_SL g769 ( .A(n_770), .Y(n_769) );
CKINVDCx20_ASAP7_75t_R g771 ( .A(n_772), .Y(n_771) );
endmodule