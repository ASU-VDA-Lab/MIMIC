module fake_jpeg_25218_n_41 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_41);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_41;

wire n_13;
wire n_21;
wire n_33;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_14;
wire n_40;
wire n_19;
wire n_20;
wire n_18;
wire n_35;
wire n_34;
wire n_30;
wire n_39;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

BUFx6f_ASAP7_75t_L g7 ( 
.A(n_6),
.Y(n_7)
);

INVx3_ASAP7_75t_L g8 ( 
.A(n_6),
.Y(n_8)
);

NOR2xp33_ASAP7_75t_SL g9 ( 
.A(n_2),
.B(n_0),
.Y(n_9)
);

NOR2xp33_ASAP7_75t_L g10 ( 
.A(n_2),
.B(n_4),
.Y(n_10)
);

INVx2_ASAP7_75t_L g11 ( 
.A(n_2),
.Y(n_11)
);

INVx2_ASAP7_75t_L g12 ( 
.A(n_3),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_5),
.Y(n_13)
);

INVx4_ASAP7_75t_L g14 ( 
.A(n_7),
.Y(n_14)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_9),
.B(n_0),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_SL g21 ( 
.A(n_15),
.B(n_16),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_9),
.B(n_0),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_10),
.B(n_1),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_17),
.B(n_20),
.Y(n_23)
);

AOI22xp33_ASAP7_75t_SL g18 ( 
.A1(n_8),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_18)
);

OAI21xp5_ASAP7_75t_L g22 ( 
.A1(n_18),
.A2(n_19),
.B(n_10),
.Y(n_22)
);

AOI22xp33_ASAP7_75t_SL g19 ( 
.A1(n_8),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_19)
);

AND2x6_ASAP7_75t_L g20 ( 
.A(n_11),
.B(n_5),
.Y(n_20)
);

OAI22xp5_ASAP7_75t_L g27 ( 
.A1(n_22),
.A2(n_12),
.B1(n_8),
.B2(n_14),
.Y(n_27)
);

OAI21xp5_ASAP7_75t_SL g25 ( 
.A1(n_20),
.A2(n_11),
.B(n_12),
.Y(n_25)
);

MAJIxp5_ASAP7_75t_L g29 ( 
.A(n_25),
.B(n_7),
.C(n_13),
.Y(n_29)
);

OAI322xp33_ASAP7_75t_L g26 ( 
.A1(n_23),
.A2(n_20),
.A3(n_15),
.B1(n_16),
.B2(n_19),
.C1(n_18),
.C2(n_17),
.Y(n_26)
);

MAJIxp5_ASAP7_75t_L g32 ( 
.A(n_26),
.B(n_30),
.C(n_21),
.Y(n_32)
);

AND2x2_ASAP7_75t_L g34 ( 
.A(n_27),
.B(n_28),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_25),
.B(n_14),
.Y(n_28)
);

MAJIxp5_ASAP7_75t_L g33 ( 
.A(n_29),
.B(n_24),
.C(n_30),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_SL g30 ( 
.A1(n_22),
.A2(n_24),
.B1(n_13),
.B2(n_7),
.Y(n_30)
);

XNOR2xp5_ASAP7_75t_L g31 ( 
.A(n_29),
.B(n_21),
.Y(n_31)
);

XNOR2xp5_ASAP7_75t_L g37 ( 
.A(n_31),
.B(n_32),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_L g35 ( 
.A1(n_33),
.A2(n_27),
.B1(n_26),
.B2(n_28),
.Y(n_35)
);

OAI21xp5_ASAP7_75t_SL g39 ( 
.A1(n_35),
.A2(n_36),
.B(n_34),
.Y(n_39)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_34),
.Y(n_36)
);

INVxp67_ASAP7_75t_L g38 ( 
.A(n_37),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_38),
.B(n_39),
.Y(n_40)
);

XOR2xp5_ASAP7_75t_L g41 ( 
.A(n_40),
.B(n_37),
.Y(n_41)
);


endmodule