module fake_jpeg_20569_n_105 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_105);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_105;

wire n_10;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

BUFx6f_ASAP7_75t_L g10 ( 
.A(n_1),
.Y(n_10)
);

BUFx12f_ASAP7_75t_L g11 ( 
.A(n_4),
.Y(n_11)
);

INVx2_ASAP7_75t_L g12 ( 
.A(n_7),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_3),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_2),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_4),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

INVx3_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

INVx3_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

BUFx10_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_2),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_21),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_22),
.Y(n_32)
);

OR2x2_ASAP7_75t_L g23 ( 
.A(n_20),
.B(n_0),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_23),
.B(n_25),
.Y(n_36)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_24),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_26),
.B(n_27),
.Y(n_29)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

AO22x1_ASAP7_75t_SL g31 ( 
.A1(n_24),
.A2(n_19),
.B1(n_10),
.B2(n_15),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_31),
.B(n_34),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_23),
.B(n_20),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_33),
.B(n_14),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_23),
.B(n_19),
.Y(n_34)
);

MAJIxp5_ASAP7_75t_L g35 ( 
.A(n_26),
.B(n_19),
.C(n_18),
.Y(n_35)
);

AOI22xp5_ASAP7_75t_SL g37 ( 
.A1(n_35),
.A2(n_24),
.B1(n_27),
.B2(n_12),
.Y(n_37)
);

OAI21xp5_ASAP7_75t_SL g51 ( 
.A1(n_37),
.A2(n_47),
.B(n_31),
.Y(n_51)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_39),
.B(n_40),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_28),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_36),
.B(n_12),
.Y(n_41)
);

CKINVDCx16_ASAP7_75t_R g52 ( 
.A(n_41),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_34),
.B(n_14),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_42),
.B(n_44),
.Y(n_56)
);

A2O1A1Ixp33_ASAP7_75t_L g43 ( 
.A1(n_36),
.A2(n_13),
.B(n_16),
.C(n_19),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_43),
.B(n_48),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_28),
.B(n_17),
.Y(n_44)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_30),
.Y(n_45)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_45),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_SL g47 ( 
.A1(n_35),
.A2(n_17),
.B1(n_18),
.B2(n_13),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_30),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_51),
.A2(n_54),
.B1(n_59),
.B2(n_21),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_46),
.A2(n_32),
.B1(n_31),
.B2(n_22),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_38),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_55),
.B(n_26),
.Y(n_63)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_48),
.Y(n_57)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_57),
.Y(n_65)
);

AOI21xp5_ASAP7_75t_L g58 ( 
.A1(n_46),
.A2(n_32),
.B(n_26),
.Y(n_58)
);

INVxp67_ASAP7_75t_L g71 ( 
.A(n_58),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_L g59 ( 
.A1(n_47),
.A2(n_22),
.B1(n_21),
.B2(n_16),
.Y(n_59)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_45),
.Y(n_61)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_61),
.Y(n_68)
);

XNOR2xp5_ASAP7_75t_L g62 ( 
.A(n_60),
.B(n_37),
.Y(n_62)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_62),
.B(n_67),
.C(n_72),
.Y(n_76)
);

CKINVDCx16_ASAP7_75t_R g74 ( 
.A(n_63),
.Y(n_74)
);

HB1xp67_ASAP7_75t_L g64 ( 
.A(n_58),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_64),
.Y(n_75)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_57),
.Y(n_66)
);

INVxp67_ASAP7_75t_L g80 ( 
.A(n_66),
.Y(n_80)
);

XNOR2xp5_ASAP7_75t_L g67 ( 
.A(n_60),
.B(n_43),
.Y(n_67)
);

FAx1_ASAP7_75t_SL g69 ( 
.A(n_56),
.B(n_26),
.CI(n_25),
.CON(n_69),
.SN(n_69)
);

NOR2xp33_ASAP7_75t_SL g79 ( 
.A(n_69),
.B(n_49),
.Y(n_79)
);

OAI21xp5_ASAP7_75t_SL g78 ( 
.A1(n_70),
.A2(n_50),
.B(n_53),
.Y(n_78)
);

XNOR2xp5_ASAP7_75t_L g72 ( 
.A(n_51),
.B(n_25),
.Y(n_72)
);

AOI21xp5_ASAP7_75t_L g73 ( 
.A1(n_71),
.A2(n_55),
.B(n_52),
.Y(n_73)
);

CKINVDCx14_ASAP7_75t_R g87 ( 
.A(n_73),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_65),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_77),
.B(n_78),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_79),
.B(n_76),
.Y(n_86)
);

A2O1A1O1Ixp25_ASAP7_75t_L g81 ( 
.A1(n_71),
.A2(n_67),
.B(n_72),
.C(n_69),
.D(n_50),
.Y(n_81)
);

NAND3xp33_ASAP7_75t_L g82 ( 
.A(n_81),
.B(n_68),
.C(n_61),
.Y(n_82)
);

AO22x1_ASAP7_75t_L g89 ( 
.A1(n_82),
.A2(n_81),
.B1(n_88),
.B2(n_87),
.Y(n_89)
);

AOI21xp5_ASAP7_75t_L g83 ( 
.A1(n_75),
.A2(n_53),
.B(n_1),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_83),
.B(n_86),
.Y(n_93)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_80),
.Y(n_84)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_84),
.Y(n_90)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_80),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_85),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_89),
.B(n_92),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_85),
.B(n_76),
.C(n_74),
.Y(n_92)
);

AOI322xp5_ASAP7_75t_L g95 ( 
.A1(n_93),
.A2(n_83),
.A3(n_15),
.B1(n_7),
.B2(n_9),
.C1(n_6),
.C2(n_8),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_95),
.B(n_25),
.C(n_9),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g96 ( 
.A(n_92),
.B(n_8),
.Y(n_96)
);

AOI31xp33_ASAP7_75t_L g101 ( 
.A1(n_96),
.A2(n_97),
.A3(n_0),
.B(n_2),
.Y(n_101)
);

OR2x2_ASAP7_75t_L g97 ( 
.A(n_91),
.B(n_89),
.Y(n_97)
);

NOR2xp67_ASAP7_75t_SL g98 ( 
.A(n_94),
.B(n_90),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_L g102 ( 
.A1(n_98),
.A2(n_99),
.B(n_100),
.Y(n_102)
);

XNOR2x2_ASAP7_75t_SL g100 ( 
.A(n_95),
.B(n_0),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_L g103 ( 
.A1(n_101),
.A2(n_4),
.B(n_5),
.Y(n_103)
);

AOI21xp5_ASAP7_75t_L g104 ( 
.A1(n_103),
.A2(n_5),
.B(n_102),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_104),
.B(n_5),
.Y(n_105)
);


endmodule