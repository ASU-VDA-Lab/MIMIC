module fake_jpeg_1282_n_188 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_188);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_188;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g48 ( 
.A(n_31),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_4),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_17),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_8),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_47),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_1),
.Y(n_53)
);

BUFx12_ASAP7_75t_L g54 ( 
.A(n_30),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_1),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_16),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_42),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_21),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_18),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_25),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_0),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_6),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_12),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_39),
.Y(n_64)
);

INVx2_ASAP7_75t_SL g65 ( 
.A(n_44),
.Y(n_65)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_13),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_12),
.Y(n_67)
);

BUFx5_ASAP7_75t_L g68 ( 
.A(n_37),
.Y(n_68)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_49),
.Y(n_69)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_69),
.Y(n_84)
);

INVx2_ASAP7_75t_SL g70 ( 
.A(n_68),
.Y(n_70)
);

OR2x2_ASAP7_75t_L g86 ( 
.A(n_70),
.B(n_65),
.Y(n_86)
);

CKINVDCx16_ASAP7_75t_R g71 ( 
.A(n_62),
.Y(n_71)
);

CKINVDCx16_ASAP7_75t_R g83 ( 
.A(n_71),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_62),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_72),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_55),
.B(n_0),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_73),
.B(n_76),
.Y(n_82)
);

BUFx12f_ASAP7_75t_L g74 ( 
.A(n_54),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_74),
.Y(n_79)
);

INVx11_ASAP7_75t_L g75 ( 
.A(n_49),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_75),
.Y(n_85)
);

INVx5_ASAP7_75t_L g76 ( 
.A(n_49),
.Y(n_76)
);

AND2x2_ASAP7_75t_SL g77 ( 
.A(n_69),
.B(n_66),
.Y(n_77)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_77),
.B(n_80),
.Y(n_93)
);

AOI21xp5_ASAP7_75t_L g80 ( 
.A1(n_70),
.A2(n_65),
.B(n_66),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_70),
.B(n_63),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_81),
.B(n_74),
.Y(n_96)
);

INVx2_ASAP7_75t_SL g107 ( 
.A(n_86),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_72),
.A2(n_67),
.B1(n_56),
.B2(n_51),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_87),
.A2(n_72),
.B1(n_76),
.B2(n_52),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_75),
.A2(n_51),
.B1(n_66),
.B2(n_67),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_88),
.A2(n_74),
.B1(n_52),
.B2(n_68),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_71),
.B(n_53),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_89),
.B(n_50),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_81),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_90),
.B(n_106),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_91),
.B(n_96),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_92),
.A2(n_79),
.B1(n_54),
.B2(n_27),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_94),
.A2(n_100),
.B1(n_105),
.B2(n_93),
.Y(n_112)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_84),
.Y(n_95)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_95),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_82),
.B(n_56),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_97),
.B(n_98),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_86),
.B(n_48),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_77),
.B(n_61),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_99),
.B(n_103),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_87),
.A2(n_64),
.B1(n_58),
.B2(n_57),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_78),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_101),
.Y(n_113)
);

HB1xp67_ASAP7_75t_L g102 ( 
.A(n_84),
.Y(n_102)
);

CKINVDCx16_ASAP7_75t_R g109 ( 
.A(n_102),
.Y(n_109)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_78),
.Y(n_103)
);

FAx1_ASAP7_75t_SL g104 ( 
.A(n_77),
.B(n_80),
.CI(n_85),
.CON(n_104),
.SN(n_104)
);

OR2x2_ASAP7_75t_L g120 ( 
.A(n_104),
.B(n_24),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_L g105 ( 
.A1(n_83),
.A2(n_60),
.B1(n_59),
.B2(n_74),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_85),
.B(n_2),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_93),
.A2(n_79),
.B1(n_54),
.B2(n_4),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_108),
.A2(n_116),
.B1(n_121),
.B2(n_7),
.Y(n_129)
);

OR2x2_ASAP7_75t_L g142 ( 
.A(n_112),
.B(n_34),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_105),
.B(n_2),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_114),
.B(n_115),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_107),
.B(n_3),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_101),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_117),
.B(n_118),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_107),
.B(n_100),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_L g133 ( 
.A1(n_120),
.A2(n_126),
.B(n_9),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_L g121 ( 
.A1(n_104),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_121)
);

BUFx24_ASAP7_75t_L g122 ( 
.A(n_104),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_122),
.Y(n_146)
);

INVx5_ASAP7_75t_L g123 ( 
.A(n_94),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_123),
.B(n_124),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_90),
.B(n_5),
.Y(n_124)
);

AOI21xp5_ASAP7_75t_L g126 ( 
.A1(n_93),
.A2(n_7),
.B(n_8),
.Y(n_126)
);

AND2x2_ASAP7_75t_SL g128 ( 
.A(n_122),
.B(n_29),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g149 ( 
.A(n_128),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_129),
.A2(n_142),
.B1(n_144),
.B2(n_14),
.Y(n_155)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_125),
.Y(n_132)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_132),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_L g150 ( 
.A1(n_133),
.A2(n_148),
.B(n_116),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_L g134 ( 
.A(n_111),
.B(n_32),
.Y(n_134)
);

XOR2xp5_ASAP7_75t_L g161 ( 
.A(n_134),
.B(n_140),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_119),
.B(n_9),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_136),
.B(n_138),
.Y(n_160)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_109),
.Y(n_137)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_137),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_120),
.B(n_33),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_127),
.B(n_110),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g163 ( 
.A(n_139),
.B(n_141),
.Y(n_163)
);

XOR2xp5_ASAP7_75t_L g140 ( 
.A(n_122),
.B(n_28),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_126),
.B(n_10),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_121),
.B(n_10),
.Y(n_143)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_143),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_123),
.A2(n_35),
.B1(n_46),
.B2(n_45),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_113),
.Y(n_145)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_145),
.Y(n_162)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_113),
.Y(n_147)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_147),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_108),
.B(n_11),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_150),
.B(n_155),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_SL g151 ( 
.A(n_128),
.B(n_11),
.C(n_13),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_151),
.B(n_152),
.Y(n_164)
);

OAI21xp33_ASAP7_75t_L g152 ( 
.A1(n_146),
.A2(n_26),
.B(n_43),
.Y(n_152)
);

INVxp67_ASAP7_75t_L g169 ( 
.A(n_152),
.Y(n_169)
);

BUFx3_ASAP7_75t_L g158 ( 
.A(n_144),
.Y(n_158)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_158),
.Y(n_168)
);

INVxp33_ASAP7_75t_SL g159 ( 
.A(n_130),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_159),
.A2(n_135),
.B1(n_133),
.B2(n_142),
.Y(n_165)
);

OR2x2_ASAP7_75t_L g177 ( 
.A(n_164),
.B(n_166),
.Y(n_177)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_165),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_159),
.A2(n_131),
.B1(n_129),
.B2(n_140),
.Y(n_166)
);

NAND4xp25_ASAP7_75t_L g167 ( 
.A(n_149),
.B(n_138),
.C(n_128),
.D(n_134),
.Y(n_167)
);

AOI321xp33_ASAP7_75t_L g175 ( 
.A1(n_167),
.A2(n_163),
.A3(n_154),
.B1(n_160),
.B2(n_157),
.C(n_14),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_161),
.B(n_23),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g176 ( 
.A(n_171),
.B(n_15),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_SL g173 ( 
.A(n_171),
.B(n_149),
.Y(n_173)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_173),
.B(n_169),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_168),
.A2(n_156),
.B1(n_153),
.B2(n_162),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_174),
.A2(n_170),
.B1(n_169),
.B2(n_15),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_175),
.B(n_176),
.Y(n_179)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_174),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_178),
.A2(n_180),
.B1(n_172),
.B2(n_177),
.Y(n_182)
);

AOI21xp5_ASAP7_75t_L g183 ( 
.A1(n_181),
.A2(n_19),
.B(n_20),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_182),
.B(n_183),
.C(n_179),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_184),
.B(n_181),
.Y(n_185)
);

FAx1_ASAP7_75t_SL g186 ( 
.A(n_185),
.B(n_22),
.CI(n_36),
.CON(n_186),
.SN(n_186)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_186),
.B(n_38),
.C(n_40),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_187),
.B(n_41),
.Y(n_188)
);


endmodule