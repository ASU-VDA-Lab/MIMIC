module real_aes_647_n_105 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_104, n_21, n_31, n_8, n_834, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_833, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_105);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_104;
input n_21;
input n_31;
input n_8;
input n_834;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_833;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_105;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_485;
wire n_822;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_364;
wire n_319;
wire n_421;
wire n_555;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_666;
wire n_551;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_786;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_732;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_781;
wire n_748;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_812;
wire n_782;
wire n_443;
wire n_565;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_505;
wire n_434;
wire n_769;
wire n_502;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_402;
wire n_552;
wire n_602;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_807;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_810;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_765;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_831;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_789;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_717;
wire n_456;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_479;
wire n_338;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_719;
wire n_473;
wire n_465;
wire n_566;
wire n_474;
wire n_829;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_729;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_804;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_802;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
NAND2xp5_ASAP7_75t_L g222 ( .A(n_0), .B(n_144), .Y(n_222) );
NAND2xp5_ASAP7_75t_L g827 ( .A(n_1), .B(n_828), .Y(n_827) );
NAND2xp5_ASAP7_75t_L g163 ( .A(n_2), .B(n_150), .Y(n_163) );
INVx1_ASAP7_75t_L g137 ( .A(n_3), .Y(n_137) );
NAND2xp33_ASAP7_75t_SL g214 ( .A(n_4), .B(n_148), .Y(n_214) );
INVx1_ASAP7_75t_L g195 ( .A(n_5), .Y(n_195) );
NAND2xp5_ASAP7_75t_SL g541 ( .A(n_6), .B(n_168), .Y(n_541) );
OAI22xp5_ASAP7_75t_SL g110 ( .A1(n_7), .A2(n_111), .B1(n_112), .B2(n_114), .Y(n_110) );
CKINVDCx20_ASAP7_75t_R g111 ( .A(n_7), .Y(n_111) );
INVx1_ASAP7_75t_L g521 ( .A(n_8), .Y(n_521) );
CKINVDCx16_ASAP7_75t_R g828 ( .A(n_9), .Y(n_828) );
AND2x2_ASAP7_75t_L g161 ( .A(n_10), .B(n_154), .Y(n_161) );
CKINVDCx5p33_ASAP7_75t_R g488 ( .A(n_11), .Y(n_488) );
INVx2_ASAP7_75t_L g155 ( .A(n_12), .Y(n_155) );
CKINVDCx20_ASAP7_75t_R g113 ( .A(n_13), .Y(n_113) );
CKINVDCx16_ASAP7_75t_R g120 ( .A(n_14), .Y(n_120) );
NOR2xp33_ASAP7_75t_L g717 ( .A(n_14), .B(n_27), .Y(n_717) );
AND3x1_ASAP7_75t_L g825 ( .A(n_14), .B(n_37), .C(n_826), .Y(n_825) );
INVx1_ASAP7_75t_L g549 ( .A(n_15), .Y(n_549) );
OAI22xp5_ASAP7_75t_SL g808 ( .A1(n_16), .A2(n_27), .B1(n_771), .B2(n_809), .Y(n_808) );
CKINVDCx20_ASAP7_75t_R g809 ( .A(n_16), .Y(n_809) );
AOI221x1_ASAP7_75t_L g208 ( .A1(n_17), .A2(n_132), .B1(n_209), .B2(n_211), .C(n_213), .Y(n_208) );
NAND2xp5_ASAP7_75t_SL g183 ( .A(n_18), .B(n_150), .Y(n_183) );
INVx1_ASAP7_75t_L g783 ( .A(n_19), .Y(n_783) );
INVx1_ASAP7_75t_L g547 ( .A(n_20), .Y(n_547) );
INVx1_ASAP7_75t_SL g470 ( .A(n_21), .Y(n_470) );
NAND2xp5_ASAP7_75t_SL g537 ( .A(n_22), .B(n_151), .Y(n_537) );
AOI21xp5_ASAP7_75t_L g164 ( .A1(n_23), .A2(n_132), .B(n_165), .Y(n_164) );
AOI221xp5_ASAP7_75t_SL g175 ( .A1(n_24), .A2(n_40), .B1(n_132), .B2(n_150), .C(n_176), .Y(n_175) );
NAND2xp5_ASAP7_75t_L g166 ( .A(n_25), .B(n_144), .Y(n_166) );
AOI33xp33_ASAP7_75t_L g507 ( .A1(n_26), .A2(n_53), .A3(n_198), .B1(n_204), .B2(n_508), .B3(n_509), .Y(n_507) );
INVx1_ASAP7_75t_L g771 ( .A(n_27), .Y(n_771) );
INVx1_ASAP7_75t_L g481 ( .A(n_28), .Y(n_481) );
OR2x2_ASAP7_75t_L g156 ( .A(n_29), .B(n_94), .Y(n_156) );
OA21x2_ASAP7_75t_L g189 ( .A1(n_29), .A2(n_94), .B(n_155), .Y(n_189) );
NAND2xp5_ASAP7_75t_L g187 ( .A(n_30), .B(n_140), .Y(n_187) );
INVxp67_ASAP7_75t_L g207 ( .A(n_31), .Y(n_207) );
AND2x2_ASAP7_75t_L g238 ( .A(n_32), .B(n_153), .Y(n_238) );
NAND2xp5_ASAP7_75t_L g467 ( .A(n_33), .B(n_196), .Y(n_467) );
AOI21xp5_ASAP7_75t_L g220 ( .A1(n_34), .A2(n_132), .B(n_221), .Y(n_220) );
NAND2xp5_ASAP7_75t_L g177 ( .A(n_35), .B(n_140), .Y(n_177) );
AND2x2_ASAP7_75t_L g133 ( .A(n_36), .B(n_134), .Y(n_133) );
AND2x2_ASAP7_75t_L g148 ( .A(n_36), .B(n_137), .Y(n_148) );
INVx1_ASAP7_75t_L g203 ( .A(n_36), .Y(n_203) );
OR2x6_ASAP7_75t_L g781 ( .A(n_37), .B(n_782), .Y(n_781) );
CKINVDCx20_ASAP7_75t_R g483 ( .A(n_38), .Y(n_483) );
NAND2xp5_ASAP7_75t_L g495 ( .A(n_39), .B(n_196), .Y(n_495) );
AOI22xp5_ASAP7_75t_L g530 ( .A1(n_41), .A2(n_168), .B1(n_212), .B2(n_531), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_42), .B(n_539), .Y(n_538) );
AOI22xp5_ASAP7_75t_L g274 ( .A1(n_43), .A2(n_84), .B1(n_132), .B2(n_201), .Y(n_274) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_44), .B(n_151), .Y(n_471) );
NAND2xp5_ASAP7_75t_L g236 ( .A(n_45), .B(n_144), .Y(n_236) );
INVx1_ASAP7_75t_L g779 ( .A(n_46), .Y(n_779) );
XNOR2xp5_ASAP7_75t_L g811 ( .A(n_47), .B(n_88), .Y(n_811) );
NAND2xp5_ASAP7_75t_SL g523 ( .A(n_48), .B(n_188), .Y(n_523) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_49), .B(n_151), .Y(n_522) );
CKINVDCx5p33_ASAP7_75t_R g534 ( .A(n_50), .Y(n_534) );
AND2x2_ASAP7_75t_L g225 ( .A(n_51), .B(n_153), .Y(n_225) );
NAND2xp5_ASAP7_75t_L g179 ( .A(n_52), .B(n_153), .Y(n_179) );
XOR2xp5_ASAP7_75t_L g803 ( .A(n_52), .B(n_804), .Y(n_803) );
NAND2xp5_ASAP7_75t_L g499 ( .A(n_54), .B(n_151), .Y(n_499) );
INVx1_ASAP7_75t_L g136 ( .A(n_55), .Y(n_136) );
INVx1_ASAP7_75t_L g146 ( .A(n_55), .Y(n_146) );
AND2x2_ASAP7_75t_L g500 ( .A(n_56), .B(n_153), .Y(n_500) );
AOI221xp5_ASAP7_75t_L g519 ( .A1(n_57), .A2(n_77), .B1(n_196), .B2(n_201), .C(n_520), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g464 ( .A(n_58), .B(n_196), .Y(n_464) );
NAND2xp5_ASAP7_75t_SL g237 ( .A(n_59), .B(n_150), .Y(n_237) );
OAI22xp5_ASAP7_75t_SL g109 ( .A1(n_60), .A2(n_110), .B1(n_115), .B2(n_116), .Y(n_109) );
CKINVDCx20_ASAP7_75t_R g115 ( .A(n_60), .Y(n_115) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_61), .B(n_212), .Y(n_490) );
AOI21xp5_ASAP7_75t_SL g459 ( .A1(n_62), .A2(n_201), .B(n_460), .Y(n_459) );
AND2x2_ASAP7_75t_L g157 ( .A(n_63), .B(n_153), .Y(n_157) );
AOI22xp5_ASAP7_75t_L g105 ( .A1(n_64), .A2(n_106), .B1(n_820), .B2(n_829), .Y(n_105) );
NAND2xp5_ASAP7_75t_L g223 ( .A(n_65), .B(n_140), .Y(n_223) );
NAND2xp5_ASAP7_75t_L g143 ( .A(n_66), .B(n_144), .Y(n_143) );
AND2x2_ASAP7_75t_SL g190 ( .A(n_67), .B(n_154), .Y(n_190) );
INVx1_ASAP7_75t_L g544 ( .A(n_68), .Y(n_544) );
XNOR2xp5_ASAP7_75t_L g112 ( .A(n_69), .B(n_113), .Y(n_112) );
AOI21xp5_ASAP7_75t_L g233 ( .A1(n_70), .A2(n_132), .B(n_234), .Y(n_233) );
INVx1_ASAP7_75t_L g498 ( .A(n_71), .Y(n_498) );
NAND2xp5_ASAP7_75t_L g167 ( .A(n_72), .B(n_140), .Y(n_167) );
AND2x2_ASAP7_75t_SL g275 ( .A(n_73), .B(n_188), .Y(n_275) );
AOI21xp5_ASAP7_75t_L g496 ( .A1(n_74), .A2(n_201), .B(n_497), .Y(n_496) );
INVx1_ASAP7_75t_L g134 ( .A(n_75), .Y(n_134) );
INVx1_ASAP7_75t_L g142 ( .A(n_75), .Y(n_142) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_76), .B(n_196), .Y(n_510) );
AND2x2_ASAP7_75t_L g472 ( .A(n_78), .B(n_211), .Y(n_472) );
INVx1_ASAP7_75t_L g545 ( .A(n_79), .Y(n_545) );
AOI21xp5_ASAP7_75t_L g468 ( .A1(n_80), .A2(n_201), .B(n_469), .Y(n_468) );
A2O1A1Ixp33_ASAP7_75t_L g535 ( .A1(n_81), .A2(n_201), .B(n_271), .C(n_536), .Y(n_535) );
NAND2xp5_ASAP7_75t_SL g149 ( .A(n_82), .B(n_150), .Y(n_149) );
AOI22xp5_ASAP7_75t_L g273 ( .A1(n_83), .A2(n_87), .B1(n_150), .B2(n_196), .Y(n_273) );
INVx1_ASAP7_75t_L g784 ( .A(n_85), .Y(n_784) );
AND2x2_ASAP7_75t_SL g457 ( .A(n_86), .B(n_211), .Y(n_457) );
AOI22xp5_ASAP7_75t_L g504 ( .A1(n_89), .A2(n_201), .B1(n_505), .B2(n_506), .Y(n_504) );
NAND2xp5_ASAP7_75t_L g186 ( .A(n_90), .B(n_144), .Y(n_186) );
NAND2xp5_ASAP7_75t_L g178 ( .A(n_91), .B(n_144), .Y(n_178) );
NAND2xp5_ASAP7_75t_SL g785 ( .A(n_92), .B(n_786), .Y(n_785) );
AOI21xp5_ASAP7_75t_L g131 ( .A1(n_93), .A2(n_132), .B(n_138), .Y(n_131) );
INVx1_ASAP7_75t_L g461 ( .A(n_95), .Y(n_461) );
NAND2xp5_ASAP7_75t_L g139 ( .A(n_96), .B(n_140), .Y(n_139) );
AND2x2_ASAP7_75t_L g511 ( .A(n_97), .B(n_211), .Y(n_511) );
A2O1A1Ixp33_ASAP7_75t_L g478 ( .A1(n_98), .A2(n_479), .B(n_480), .C(n_482), .Y(n_478) );
INVxp67_ASAP7_75t_L g210 ( .A(n_99), .Y(n_210) );
NAND2xp5_ASAP7_75t_L g224 ( .A(n_100), .B(n_150), .Y(n_224) );
NAND2xp5_ASAP7_75t_L g235 ( .A(n_101), .B(n_140), .Y(n_235) );
AOI21xp5_ASAP7_75t_L g184 ( .A1(n_102), .A2(n_132), .B(n_185), .Y(n_184) );
BUFx2_ASAP7_75t_SL g777 ( .A(n_103), .Y(n_777) );
BUFx2_ASAP7_75t_L g795 ( .A(n_103), .Y(n_795) );
NAND2xp5_ASAP7_75t_L g463 ( .A(n_104), .B(n_151), .Y(n_463) );
AND2x4_ASAP7_75t_L g106 ( .A(n_107), .B(n_796), .Y(n_106) );
AOI21xp5_ASAP7_75t_L g107 ( .A1(n_108), .A2(n_773), .B(n_790), .Y(n_107) );
NOR2xp33_ASAP7_75t_L g108 ( .A(n_109), .B(n_117), .Y(n_108) );
CKINVDCx16_ASAP7_75t_R g819 ( .A(n_109), .Y(n_819) );
INVxp33_ASAP7_75t_L g116 ( .A(n_110), .Y(n_116) );
INVx1_ASAP7_75t_L g114 ( .A(n_112), .Y(n_114) );
INVx1_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
HB1xp67_ASAP7_75t_L g818 ( .A(n_118), .Y(n_818) );
OAI21x1_ASAP7_75t_L g118 ( .A1(n_119), .A2(n_121), .B(n_447), .Y(n_118) );
HB1xp67_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
CKINVDCx16_ASAP7_75t_R g772 ( .A(n_120), .Y(n_772) );
OR2x2_ASAP7_75t_L g780 ( .A(n_120), .B(n_781), .Y(n_780) );
NAND2xp5_ASAP7_75t_L g788 ( .A(n_120), .B(n_789), .Y(n_788) );
AND2x4_ASAP7_75t_L g121 ( .A(n_122), .B(n_386), .Y(n_121) );
NOR3xp33_ASAP7_75t_L g122 ( .A(n_123), .B(n_279), .C(n_330), .Y(n_122) );
OAI211xp5_ASAP7_75t_SL g123 ( .A1(n_124), .A2(n_169), .B(n_226), .C(n_257), .Y(n_123) );
INVxp67_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
NOR2xp33_ASAP7_75t_L g125 ( .A(n_126), .B(n_158), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
HB1xp67_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
NAND2xp5_ASAP7_75t_L g394 ( .A(n_128), .B(n_231), .Y(n_394) );
INVx1_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
AND2x2_ASAP7_75t_L g239 ( .A(n_129), .B(n_160), .Y(n_239) );
NAND2xp5_ASAP7_75t_L g245 ( .A(n_129), .B(n_246), .Y(n_245) );
OR2x2_ASAP7_75t_L g256 ( .A(n_129), .B(n_246), .Y(n_256) );
NAND2xp5_ASAP7_75t_L g277 ( .A(n_129), .B(n_278), .Y(n_277) );
AND2x2_ASAP7_75t_L g293 ( .A(n_129), .B(n_269), .Y(n_293) );
INVx2_ASAP7_75t_L g319 ( .A(n_129), .Y(n_319) );
AND2x4_ASAP7_75t_L g328 ( .A(n_129), .B(n_329), .Y(n_328) );
AND2x2_ASAP7_75t_L g433 ( .A(n_129), .B(n_300), .Y(n_433) );
AO21x2_ASAP7_75t_L g129 ( .A1(n_130), .A2(n_152), .B(n_157), .Y(n_129) );
NAND2xp5_ASAP7_75t_L g130 ( .A(n_131), .B(n_149), .Y(n_130) );
AND2x6_ASAP7_75t_L g132 ( .A(n_133), .B(n_135), .Y(n_132) );
BUFx3_ASAP7_75t_L g200 ( .A(n_133), .Y(n_200) );
AND2x6_ASAP7_75t_L g144 ( .A(n_134), .B(n_145), .Y(n_144) );
INVx2_ASAP7_75t_L g205 ( .A(n_134), .Y(n_205) );
AND2x4_ASAP7_75t_L g201 ( .A(n_135), .B(n_202), .Y(n_201) );
AND2x2_ASAP7_75t_L g135 ( .A(n_136), .B(n_137), .Y(n_135) );
AND2x4_ASAP7_75t_L g140 ( .A(n_136), .B(n_141), .Y(n_140) );
INVx2_ASAP7_75t_L g198 ( .A(n_136), .Y(n_198) );
HB1xp67_ASAP7_75t_L g199 ( .A(n_137), .Y(n_199) );
AOI21xp5_ASAP7_75t_L g138 ( .A1(n_139), .A2(n_143), .B(n_147), .Y(n_138) );
INVxp67_ASAP7_75t_L g550 ( .A(n_140), .Y(n_550) );
AND2x4_ASAP7_75t_L g151 ( .A(n_141), .B(n_145), .Y(n_151) );
INVx2_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
INVxp67_ASAP7_75t_L g548 ( .A(n_144), .Y(n_548) );
INVx2_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
AOI21xp5_ASAP7_75t_L g165 ( .A1(n_147), .A2(n_166), .B(n_167), .Y(n_165) );
AOI21xp5_ASAP7_75t_L g176 ( .A1(n_147), .A2(n_177), .B(n_178), .Y(n_176) );
AOI21xp5_ASAP7_75t_L g185 ( .A1(n_147), .A2(n_186), .B(n_187), .Y(n_185) );
AOI21xp5_ASAP7_75t_L g221 ( .A1(n_147), .A2(n_222), .B(n_223), .Y(n_221) );
AOI21xp5_ASAP7_75t_L g234 ( .A1(n_147), .A2(n_235), .B(n_236), .Y(n_234) );
O2A1O1Ixp33_ASAP7_75t_L g460 ( .A1(n_147), .A2(n_461), .B(n_462), .C(n_463), .Y(n_460) );
O2A1O1Ixp33_ASAP7_75t_SL g469 ( .A1(n_147), .A2(n_462), .B(n_470), .C(n_471), .Y(n_469) );
O2A1O1Ixp33_ASAP7_75t_L g497 ( .A1(n_147), .A2(n_462), .B(n_498), .C(n_499), .Y(n_497) );
INVx1_ASAP7_75t_L g505 ( .A(n_147), .Y(n_505) );
O2A1O1Ixp33_ASAP7_75t_SL g520 ( .A1(n_147), .A2(n_462), .B(n_521), .C(n_522), .Y(n_520) );
AOI21xp5_ASAP7_75t_L g536 ( .A1(n_147), .A2(n_537), .B(n_538), .Y(n_536) );
NOR2xp33_ASAP7_75t_L g551 ( .A(n_147), .B(n_168), .Y(n_551) );
INVx5_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
AND2x4_ASAP7_75t_L g150 ( .A(n_148), .B(n_151), .Y(n_150) );
HB1xp67_ASAP7_75t_L g482 ( .A(n_148), .Y(n_482) );
INVx1_ASAP7_75t_L g215 ( .A(n_151), .Y(n_215) );
AO21x2_ASAP7_75t_L g231 ( .A1(n_152), .A2(n_232), .B(n_238), .Y(n_231) );
AO21x2_ASAP7_75t_L g246 ( .A1(n_152), .A2(n_232), .B(n_238), .Y(n_246) );
AO21x2_ASAP7_75t_L g465 ( .A1(n_152), .A2(n_466), .B(n_472), .Y(n_465) );
CKINVDCx5p33_ASAP7_75t_R g152 ( .A(n_153), .Y(n_152) );
OA21x2_ASAP7_75t_L g174 ( .A1(n_153), .A2(n_175), .B(n_179), .Y(n_174) );
BUFx6f_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
AND2x2_ASAP7_75t_SL g154 ( .A(n_155), .B(n_156), .Y(n_154) );
AND2x4_ASAP7_75t_L g168 ( .A(n_155), .B(n_156), .Y(n_168) );
AND2x2_ASAP7_75t_L g317 ( .A(n_158), .B(n_318), .Y(n_317) );
OAI32xp33_ASAP7_75t_L g400 ( .A1(n_158), .A2(n_322), .A3(n_326), .B1(n_333), .B2(n_401), .Y(n_400) );
NAND2xp5_ASAP7_75t_L g432 ( .A(n_158), .B(n_433), .Y(n_432) );
INVx2_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
AND2x2_ASAP7_75t_L g254 ( .A(n_159), .B(n_255), .Y(n_254) );
NAND3xp33_ASAP7_75t_L g327 ( .A(n_159), .B(n_249), .C(n_328), .Y(n_327) );
OR2x2_ASAP7_75t_L g353 ( .A(n_159), .B(n_256), .Y(n_353) );
INVx2_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
HB1xp67_ASAP7_75t_L g243 ( .A(n_160), .Y(n_243) );
INVx5_ASAP7_75t_L g278 ( .A(n_160), .Y(n_278) );
AND2x4_ASAP7_75t_L g334 ( .A(n_160), .B(n_246), .Y(n_334) );
OR2x2_ASAP7_75t_L g349 ( .A(n_160), .B(n_269), .Y(n_349) );
OR2x2_ASAP7_75t_L g375 ( .A(n_160), .B(n_231), .Y(n_375) );
AND2x2_ASAP7_75t_L g383 ( .A(n_160), .B(n_329), .Y(n_383) );
AND2x4_ASAP7_75t_SL g408 ( .A(n_160), .B(n_328), .Y(n_408) );
OR2x6_ASAP7_75t_L g160 ( .A(n_161), .B(n_162), .Y(n_160) );
AOI21xp5_ASAP7_75t_L g162 ( .A1(n_163), .A2(n_164), .B(n_168), .Y(n_162) );
NOR2xp33_ASAP7_75t_L g194 ( .A(n_168), .B(n_195), .Y(n_194) );
NOR2xp33_ASAP7_75t_L g206 ( .A(n_168), .B(n_207), .Y(n_206) );
NOR2xp33_ASAP7_75t_L g209 ( .A(n_168), .B(n_210), .Y(n_209) );
NOR3xp33_ASAP7_75t_L g213 ( .A(n_168), .B(n_214), .C(n_215), .Y(n_213) );
AOI21xp5_ASAP7_75t_L g458 ( .A1(n_168), .A2(n_459), .B(n_464), .Y(n_458) );
INVx1_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
NAND2xp5_ASAP7_75t_L g404 ( .A(n_170), .B(n_328), .Y(n_404) );
AND2x2_ASAP7_75t_L g170 ( .A(n_171), .B(n_180), .Y(n_170) );
NAND2xp5_ASAP7_75t_L g302 ( .A(n_171), .B(n_303), .Y(n_302) );
INVx1_ASAP7_75t_L g171 ( .A(n_172), .Y(n_171) );
OR2x6_ASAP7_75t_SL g228 ( .A(n_172), .B(n_229), .Y(n_228) );
INVxp67_ASAP7_75t_SL g172 ( .A(n_173), .Y(n_172) );
INVx1_ASAP7_75t_L g253 ( .A(n_173), .Y(n_253) );
NAND2xp5_ASAP7_75t_L g306 ( .A(n_173), .B(n_288), .Y(n_306) );
HB1xp67_ASAP7_75t_L g444 ( .A(n_173), .Y(n_444) );
INVx1_ASAP7_75t_L g173 ( .A(n_174), .Y(n_173) );
INVx2_ASAP7_75t_L g261 ( .A(n_174), .Y(n_261) );
AND2x2_ASAP7_75t_L g286 ( .A(n_174), .B(n_217), .Y(n_286) );
INVx2_ASAP7_75t_L g314 ( .A(n_174), .Y(n_314) );
NAND2xp5_ASAP7_75t_L g355 ( .A(n_174), .B(n_181), .Y(n_355) );
BUFx3_ASAP7_75t_L g379 ( .A(n_174), .Y(n_379) );
OR2x2_ASAP7_75t_L g391 ( .A(n_174), .B(n_181), .Y(n_391) );
HB1xp67_ASAP7_75t_L g399 ( .A(n_174), .Y(n_399) );
AOI22xp5_ASAP7_75t_L g421 ( .A1(n_180), .A2(n_422), .B1(n_425), .B2(n_426), .Y(n_421) );
AND2x2_ASAP7_75t_L g180 ( .A(n_181), .B(n_191), .Y(n_180) );
INVx1_ASAP7_75t_L g249 ( .A(n_181), .Y(n_249) );
OR2x2_ASAP7_75t_L g260 ( .A(n_181), .B(n_261), .Y(n_260) );
INVx2_ASAP7_75t_L g267 ( .A(n_181), .Y(n_267) );
AND2x4_ASAP7_75t_SL g284 ( .A(n_181), .B(n_192), .Y(n_284) );
AND2x4_ASAP7_75t_L g289 ( .A(n_181), .B(n_290), .Y(n_289) );
INVx2_ASAP7_75t_L g298 ( .A(n_181), .Y(n_298) );
OR2x2_ASAP7_75t_L g304 ( .A(n_181), .B(n_192), .Y(n_304) );
OR2x2_ASAP7_75t_L g305 ( .A(n_181), .B(n_306), .Y(n_305) );
HB1xp67_ASAP7_75t_L g416 ( .A(n_181), .Y(n_416) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_181), .B(n_286), .Y(n_420) );
OR2x2_ASAP7_75t_L g436 ( .A(n_181), .B(n_339), .Y(n_436) );
OR2x6_ASAP7_75t_L g181 ( .A(n_182), .B(n_190), .Y(n_181) );
AOI21xp5_ASAP7_75t_L g182 ( .A1(n_183), .A2(n_184), .B(n_188), .Y(n_182) );
INVx2_ASAP7_75t_SL g271 ( .A(n_188), .Y(n_271) );
OA21x2_ASAP7_75t_L g518 ( .A1(n_188), .A2(n_519), .B(n_523), .Y(n_518) );
BUFx4f_ASAP7_75t_L g188 ( .A(n_189), .Y(n_188) );
INVx3_ASAP7_75t_L g212 ( .A(n_189), .Y(n_212) );
NAND2xp5_ASAP7_75t_L g248 ( .A(n_191), .B(n_249), .Y(n_248) );
INVx1_ASAP7_75t_L g262 ( .A(n_191), .Y(n_262) );
AND2x2_ASAP7_75t_SL g369 ( .A(n_191), .B(n_253), .Y(n_369) );
AND2x4_ASAP7_75t_L g191 ( .A(n_192), .B(n_216), .Y(n_191) );
NAND2xp5_ASAP7_75t_L g229 ( .A(n_192), .B(n_217), .Y(n_229) );
NOR2xp33_ASAP7_75t_L g250 ( .A(n_192), .B(n_251), .Y(n_250) );
NAND2xp5_ASAP7_75t_L g265 ( .A(n_192), .B(n_261), .Y(n_265) );
INVx3_ASAP7_75t_L g290 ( .A(n_192), .Y(n_290) );
INVx1_ASAP7_75t_L g323 ( .A(n_192), .Y(n_323) );
AND2x2_ASAP7_75t_L g403 ( .A(n_192), .B(n_267), .Y(n_403) );
AND2x4_ASAP7_75t_L g192 ( .A(n_193), .B(n_208), .Y(n_192) );
AOI22xp5_ASAP7_75t_L g193 ( .A1(n_194), .A2(n_196), .B1(n_201), .B2(n_206), .Y(n_193) );
INVx1_ASAP7_75t_L g491 ( .A(n_196), .Y(n_491) );
AND2x4_ASAP7_75t_L g196 ( .A(n_197), .B(n_200), .Y(n_196) );
INVx1_ASAP7_75t_L g532 ( .A(n_197), .Y(n_532) );
AND2x2_ASAP7_75t_L g197 ( .A(n_198), .B(n_199), .Y(n_197) );
OR2x6_ASAP7_75t_L g462 ( .A(n_198), .B(n_205), .Y(n_462) );
INVxp33_ASAP7_75t_L g508 ( .A(n_198), .Y(n_508) );
INVx1_ASAP7_75t_L g533 ( .A(n_200), .Y(n_533) );
INVxp67_ASAP7_75t_L g489 ( .A(n_201), .Y(n_489) );
NOR2x1p5_ASAP7_75t_L g202 ( .A(n_203), .B(n_204), .Y(n_202) );
INVx1_ASAP7_75t_L g509 ( .A(n_204), .Y(n_509) );
INVx3_ASAP7_75t_L g204 ( .A(n_205), .Y(n_204) );
OAI22xp5_ASAP7_75t_L g477 ( .A1(n_211), .A2(n_478), .B1(n_483), .B2(n_484), .Y(n_477) );
INVx3_ASAP7_75t_L g484 ( .A(n_211), .Y(n_484) );
INVx4_ASAP7_75t_L g211 ( .A(n_212), .Y(n_211) );
AOI21x1_ASAP7_75t_L g218 ( .A1(n_212), .A2(n_219), .B(n_225), .Y(n_218) );
NAND2xp5_ASAP7_75t_L g486 ( .A(n_212), .B(n_487), .Y(n_486) );
NOR2xp33_ASAP7_75t_L g480 ( .A(n_215), .B(n_481), .Y(n_480) );
OAI22xp5_ASAP7_75t_L g543 ( .A1(n_215), .A2(n_462), .B1(n_544), .B2(n_545), .Y(n_543) );
INVx2_ASAP7_75t_L g216 ( .A(n_217), .Y(n_216) );
NAND2xp5_ASAP7_75t_L g266 ( .A(n_217), .B(n_267), .Y(n_266) );
INVx1_ASAP7_75t_L g288 ( .A(n_217), .Y(n_288) );
AND2x2_ASAP7_75t_L g313 ( .A(n_217), .B(n_314), .Y(n_313) );
OR2x2_ASAP7_75t_L g339 ( .A(n_217), .B(n_261), .Y(n_339) );
NAND2xp5_ASAP7_75t_L g356 ( .A(n_217), .B(n_290), .Y(n_356) );
INVx1_ASAP7_75t_L g362 ( .A(n_217), .Y(n_362) );
INVx3_ASAP7_75t_L g217 ( .A(n_218), .Y(n_217) );
NAND2xp5_ASAP7_75t_L g219 ( .A(n_220), .B(n_224), .Y(n_219) );
AOI222xp33_ASAP7_75t_SL g226 ( .A1(n_227), .A2(n_230), .B1(n_240), .B2(n_247), .C1(n_250), .C2(n_254), .Y(n_226) );
CKINVDCx16_ASAP7_75t_R g227 ( .A(n_228), .Y(n_227) );
AND2x2_ASAP7_75t_L g230 ( .A(n_231), .B(n_239), .Y(n_230) );
NOR2xp33_ASAP7_75t_L g351 ( .A(n_231), .B(n_300), .Y(n_351) );
AND2x4_ASAP7_75t_L g367 ( .A(n_231), .B(n_278), .Y(n_367) );
NAND2xp5_ASAP7_75t_L g232 ( .A(n_233), .B(n_237), .Y(n_232) );
INVx2_ASAP7_75t_L g240 ( .A(n_241), .Y(n_240) );
NAND2xp5_ASAP7_75t_SL g241 ( .A(n_242), .B(n_244), .Y(n_241) );
INVx1_ASAP7_75t_L g242 ( .A(n_243), .Y(n_242) );
AND2x2_ASAP7_75t_L g292 ( .A(n_243), .B(n_293), .Y(n_292) );
AOI222xp33_ASAP7_75t_L g257 ( .A1(n_244), .A2(n_258), .B1(n_263), .B2(n_268), .C1(n_276), .C2(n_833), .Y(n_257) );
INVx1_ASAP7_75t_L g244 ( .A(n_245), .Y(n_244) );
OR2x2_ASAP7_75t_L g396 ( .A(n_245), .B(n_300), .Y(n_396) );
OR2x2_ASAP7_75t_L g439 ( .A(n_245), .B(n_345), .Y(n_439) );
AND2x2_ASAP7_75t_L g268 ( .A(n_246), .B(n_269), .Y(n_268) );
INVx2_ASAP7_75t_L g329 ( .A(n_246), .Y(n_329) );
HB1xp67_ASAP7_75t_L g344 ( .A(n_246), .Y(n_344) );
O2A1O1Ixp33_ASAP7_75t_L g357 ( .A1(n_247), .A2(n_358), .B(n_363), .C(n_364), .Y(n_357) );
INVx1_ASAP7_75t_SL g247 ( .A(n_248), .Y(n_247) );
INVx1_ASAP7_75t_L g385 ( .A(n_249), .Y(n_385) );
INVx1_ASAP7_75t_L g251 ( .A(n_252), .Y(n_251) );
HB1xp67_ASAP7_75t_L g252 ( .A(n_253), .Y(n_252) );
INVx2_ASAP7_75t_L g315 ( .A(n_254), .Y(n_315) );
AND2x2_ASAP7_75t_L g299 ( .A(n_255), .B(n_300), .Y(n_299) );
AND2x2_ASAP7_75t_L g308 ( .A(n_255), .B(n_309), .Y(n_308) );
INVx2_ASAP7_75t_L g255 ( .A(n_256), .Y(n_255) );
OAI31xp33_ASAP7_75t_L g350 ( .A1(n_258), .A2(n_276), .A3(n_351), .B(n_352), .Y(n_350) );
INVx1_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
A2O1A1Ixp33_ASAP7_75t_L g352 ( .A1(n_259), .A2(n_309), .B(n_353), .C(n_354), .Y(n_352) );
OR2x2_ASAP7_75t_L g259 ( .A(n_260), .B(n_262), .Y(n_259) );
OR2x2_ASAP7_75t_L g341 ( .A(n_260), .B(n_290), .Y(n_341) );
INVx2_ASAP7_75t_SL g263 ( .A(n_264), .Y(n_263) );
OR2x2_ASAP7_75t_L g264 ( .A(n_265), .B(n_266), .Y(n_264) );
BUFx2_ASAP7_75t_L g309 ( .A(n_269), .Y(n_309) );
AND2x2_ASAP7_75t_L g318 ( .A(n_269), .B(n_319), .Y(n_318) );
INVx2_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
BUFx6f_ASAP7_75t_L g300 ( .A(n_270), .Y(n_300) );
AOI21x1_ASAP7_75t_L g270 ( .A1(n_271), .A2(n_272), .B(n_275), .Y(n_270) );
AO21x2_ASAP7_75t_L g502 ( .A1(n_271), .A2(n_503), .B(n_511), .Y(n_502) );
AO21x2_ASAP7_75t_L g562 ( .A1(n_271), .A2(n_503), .B(n_511), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g272 ( .A(n_273), .B(n_274), .Y(n_272) );
INVx1_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
NAND2xp5_ASAP7_75t_L g427 ( .A(n_278), .B(n_335), .Y(n_427) );
OAI211xp5_ASAP7_75t_L g279 ( .A1(n_280), .A2(n_291), .B(n_294), .C(n_316), .Y(n_279) );
INVxp33_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
NAND2xp5_ASAP7_75t_SL g281 ( .A(n_282), .B(n_287), .Y(n_281) );
OR2x2_ASAP7_75t_L g282 ( .A(n_283), .B(n_285), .Y(n_282) );
INVx1_ASAP7_75t_SL g283 ( .A(n_284), .Y(n_283) );
AND2x2_ASAP7_75t_L g320 ( .A(n_284), .B(n_313), .Y(n_320) );
OR2x2_ASAP7_75t_L g296 ( .A(n_285), .B(n_297), .Y(n_296) );
OR2x2_ASAP7_75t_L g326 ( .A(n_285), .B(n_300), .Y(n_326) );
INVx2_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
AND2x2_ASAP7_75t_L g402 ( .A(n_286), .B(n_403), .Y(n_402) );
INVx1_ASAP7_75t_L g425 ( .A(n_287), .Y(n_425) );
NAND2xp5_ASAP7_75t_L g287 ( .A(n_288), .B(n_289), .Y(n_287) );
NAND2xp5_ASAP7_75t_L g337 ( .A(n_289), .B(n_338), .Y(n_337) );
NAND2xp5_ASAP7_75t_L g359 ( .A(n_289), .B(n_360), .Y(n_359) );
AND2x2_ASAP7_75t_L g437 ( .A(n_289), .B(n_313), .Y(n_437) );
NAND2xp5_ASAP7_75t_L g442 ( .A(n_289), .B(n_443), .Y(n_442) );
AND2x2_ASAP7_75t_L g380 ( .A(n_290), .B(n_362), .Y(n_380) );
INVx1_ASAP7_75t_SL g291 ( .A(n_292), .Y(n_291) );
AOI322xp5_ASAP7_75t_L g434 ( .A1(n_293), .A2(n_313), .A3(n_367), .B1(n_392), .B2(n_435), .C1(n_437), .C2(n_438), .Y(n_434) );
AOI211xp5_ASAP7_75t_SL g294 ( .A1(n_295), .A2(n_299), .B(n_301), .C(n_310), .Y(n_294) );
INVx1_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
NAND2xp5_ASAP7_75t_L g347 ( .A(n_297), .B(n_325), .Y(n_347) );
INVx1_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
AND2x2_ASAP7_75t_L g312 ( .A(n_298), .B(n_313), .Y(n_312) );
NOR2x1p5_ASAP7_75t_L g378 ( .A(n_298), .B(n_379), .Y(n_378) );
HB1xp67_ASAP7_75t_L g411 ( .A(n_298), .Y(n_411) );
O2A1O1Ixp33_ASAP7_75t_L g316 ( .A1(n_299), .A2(n_317), .B(n_320), .C(n_321), .Y(n_316) );
AND2x4_ASAP7_75t_L g335 ( .A(n_300), .B(n_319), .Y(n_335) );
INVx2_ASAP7_75t_L g345 ( .A(n_300), .Y(n_345) );
NAND2xp5_ASAP7_75t_SL g365 ( .A(n_300), .B(n_334), .Y(n_365) );
AND2x2_ASAP7_75t_L g407 ( .A(n_300), .B(n_408), .Y(n_407) );
NOR2xp33_ASAP7_75t_L g445 ( .A(n_300), .B(n_424), .Y(n_445) );
AND2x2_ASAP7_75t_L g446 ( .A(n_300), .B(n_328), .Y(n_446) );
AOI21xp33_ASAP7_75t_L g301 ( .A1(n_302), .A2(n_305), .B(n_307), .Y(n_301) );
AND2x2_ASAP7_75t_L g397 ( .A(n_303), .B(n_398), .Y(n_397) );
INVx1_ASAP7_75t_SL g303 ( .A(n_304), .Y(n_303) );
INVx1_ASAP7_75t_L g325 ( .A(n_306), .Y(n_325) );
INVx2_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
NOR2xp33_ASAP7_75t_L g310 ( .A(n_311), .B(n_315), .Y(n_310) );
INVx1_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
NAND2xp5_ASAP7_75t_L g373 ( .A(n_318), .B(n_374), .Y(n_373) );
INVx1_ASAP7_75t_L g412 ( .A(n_318), .Y(n_412) );
O2A1O1Ixp33_ASAP7_75t_SL g321 ( .A1(n_322), .A2(n_324), .B(n_326), .C(n_327), .Y(n_321) );
INVx1_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
INVx1_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
HB1xp67_ASAP7_75t_L g409 ( .A(n_325), .Y(n_409) );
INVx3_ASAP7_75t_SL g424 ( .A(n_328), .Y(n_424) );
NAND5xp2_ASAP7_75t_L g330 ( .A(n_331), .B(n_350), .C(n_357), .D(n_370), .E(n_381), .Y(n_330) );
AOI222xp33_ASAP7_75t_L g331 ( .A1(n_332), .A2(n_336), .B1(n_340), .B2(n_342), .C1(n_346), .C2(n_348), .Y(n_331) );
NOR2xp33_ASAP7_75t_L g332 ( .A(n_333), .B(n_335), .Y(n_332) );
AOI22xp5_ASAP7_75t_L g413 ( .A1(n_333), .A2(n_414), .B1(n_418), .B2(n_419), .Y(n_413) );
INVx2_ASAP7_75t_SL g333 ( .A(n_334), .Y(n_333) );
AND2x2_ASAP7_75t_L g363 ( .A(n_334), .B(n_335), .Y(n_363) );
INVx1_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
INVx1_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
INVx1_ASAP7_75t_SL g340 ( .A(n_341), .Y(n_340) );
NOR2xp33_ASAP7_75t_L g342 ( .A(n_343), .B(n_345), .Y(n_342) );
INVx1_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
NAND2xp5_ASAP7_75t_SL g430 ( .A(n_344), .B(n_431), .Y(n_430) );
NAND2xp5_ASAP7_75t_L g366 ( .A(n_345), .B(n_367), .Y(n_366) );
AND2x2_ASAP7_75t_L g382 ( .A(n_345), .B(n_383), .Y(n_382) );
OR2x2_ASAP7_75t_L g393 ( .A(n_345), .B(n_394), .Y(n_393) );
INVx1_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
INVx1_ASAP7_75t_SL g348 ( .A(n_349), .Y(n_348) );
OR2x2_ASAP7_75t_L g423 ( .A(n_349), .B(n_424), .Y(n_423) );
OR2x2_ASAP7_75t_L g354 ( .A(n_355), .B(n_356), .Y(n_354) );
INVx1_ASAP7_75t_L g371 ( .A(n_356), .Y(n_371) );
INVxp67_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
INVxp67_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
HB1xp67_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
AOI21xp33_ASAP7_75t_L g364 ( .A1(n_365), .A2(n_366), .B(n_368), .Y(n_364) );
AOI22xp33_ASAP7_75t_L g370 ( .A1(n_367), .A2(n_371), .B1(n_372), .B2(n_376), .Y(n_370) );
HB1xp67_ASAP7_75t_L g418 ( .A(n_367), .Y(n_418) );
INVx2_ASAP7_75t_SL g368 ( .A(n_369), .Y(n_368) );
AND2x2_ASAP7_75t_L g384 ( .A(n_369), .B(n_385), .Y(n_384) );
AND2x2_ASAP7_75t_L g389 ( .A(n_371), .B(n_390), .Y(n_389) );
INVx1_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
INVx1_ASAP7_75t_SL g374 ( .A(n_375), .Y(n_374) );
INVx1_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
NAND2xp5_ASAP7_75t_L g377 ( .A(n_378), .B(n_380), .Y(n_377) );
INVx1_ASAP7_75t_SL g417 ( .A(n_380), .Y(n_417) );
NAND2xp5_ASAP7_75t_L g381 ( .A(n_382), .B(n_384), .Y(n_381) );
NOR3xp33_ASAP7_75t_L g386 ( .A(n_387), .B(n_405), .C(n_428), .Y(n_386) );
NAND2xp5_ASAP7_75t_SL g387 ( .A(n_388), .B(n_404), .Y(n_387) );
AOI221xp5_ASAP7_75t_L g388 ( .A1(n_389), .A2(n_392), .B1(n_395), .B2(n_397), .C(n_400), .Y(n_388) );
INVx1_ASAP7_75t_SL g390 ( .A(n_391), .Y(n_390) );
OR2x2_ASAP7_75t_L g429 ( .A(n_391), .B(n_417), .Y(n_429) );
INVx1_ASAP7_75t_SL g392 ( .A(n_393), .Y(n_392) );
INVx1_ASAP7_75t_SL g395 ( .A(n_396), .Y(n_395) );
HB1xp67_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
INVx1_ASAP7_75t_SL g401 ( .A(n_402), .Y(n_401) );
OAI321xp33_ASAP7_75t_L g405 ( .A1(n_406), .A2(n_409), .A3(n_410), .B1(n_412), .B2(n_413), .C(n_421), .Y(n_405) );
INVx1_ASAP7_75t_SL g406 ( .A(n_407), .Y(n_406) );
INVx1_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
INVx1_ASAP7_75t_SL g414 ( .A(n_415), .Y(n_414) );
OR2x2_ASAP7_75t_L g415 ( .A(n_416), .B(n_417), .Y(n_415) );
AOI22xp33_ASAP7_75t_L g440 ( .A1(n_419), .A2(n_441), .B1(n_445), .B2(n_446), .Y(n_440) );
INVx1_ASAP7_75t_SL g419 ( .A(n_420), .Y(n_419) );
INVx1_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
INVx1_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
OAI211xp5_ASAP7_75t_SL g428 ( .A1(n_429), .A2(n_430), .B(n_434), .C(n_440), .Y(n_428) );
INVx1_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
INVx1_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
INVx1_ASAP7_75t_SL g438 ( .A(n_439), .Y(n_438) );
INVx1_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
INVxp67_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
NOR2x1_ASAP7_75t_L g447 ( .A(n_448), .B(n_768), .Y(n_447) );
NAND2xp5_ASAP7_75t_L g448 ( .A(n_449), .B(n_718), .Y(n_448) );
OAI21xp5_ASAP7_75t_L g449 ( .A1(n_450), .A2(n_658), .B(n_717), .Y(n_449) );
NOR3xp33_ASAP7_75t_L g768 ( .A(n_450), .B(n_719), .C(n_769), .Y(n_768) );
INVx1_ASAP7_75t_L g814 ( .A(n_450), .Y(n_814) );
NAND2xp5_ASAP7_75t_L g450 ( .A(n_451), .B(n_622), .Y(n_450) );
NOR3xp33_ASAP7_75t_L g451 ( .A(n_452), .B(n_563), .C(n_592), .Y(n_451) );
NAND2xp5_ASAP7_75t_SL g452 ( .A(n_453), .B(n_552), .Y(n_452) );
AOI22xp5_ASAP7_75t_L g453 ( .A1(n_454), .A2(n_473), .B1(n_512), .B2(n_524), .Y(n_453) );
NAND2x1_ASAP7_75t_L g754 ( .A(n_454), .B(n_553), .Y(n_754) );
INVx2_ASAP7_75t_SL g454 ( .A(n_455), .Y(n_454) );
OR2x2_ASAP7_75t_L g455 ( .A(n_456), .B(n_465), .Y(n_455) );
INVx2_ASAP7_75t_L g526 ( .A(n_456), .Y(n_526) );
INVx4_ASAP7_75t_L g568 ( .A(n_456), .Y(n_568) );
BUFx6f_ASAP7_75t_L g588 ( .A(n_456), .Y(n_588) );
AND2x4_ASAP7_75t_L g599 ( .A(n_456), .B(n_567), .Y(n_599) );
AND2x2_ASAP7_75t_L g605 ( .A(n_456), .B(n_529), .Y(n_605) );
NOR2x1_ASAP7_75t_SL g678 ( .A(n_456), .B(n_540), .Y(n_678) );
OR2x6_ASAP7_75t_L g456 ( .A(n_457), .B(n_458), .Y(n_456) );
INVxp67_ASAP7_75t_L g479 ( .A(n_462), .Y(n_479) );
INVx2_ASAP7_75t_L g539 ( .A(n_462), .Y(n_539) );
INVx2_ASAP7_75t_L g571 ( .A(n_465), .Y(n_571) );
HB1xp67_ASAP7_75t_L g585 ( .A(n_465), .Y(n_585) );
INVx1_ASAP7_75t_L g596 ( .A(n_465), .Y(n_596) );
HB1xp67_ASAP7_75t_L g608 ( .A(n_465), .Y(n_608) );
AND2x2_ASAP7_75t_L g640 ( .A(n_465), .B(n_540), .Y(n_640) );
INVx1_ASAP7_75t_L g666 ( .A(n_465), .Y(n_666) );
AND2x2_ASAP7_75t_L g728 ( .A(n_465), .B(n_556), .Y(n_728) );
NAND2xp5_ASAP7_75t_L g466 ( .A(n_467), .B(n_468), .Y(n_466) );
AND2x2_ASAP7_75t_L g473 ( .A(n_474), .B(n_492), .Y(n_473) );
INVx1_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
AND2x2_ASAP7_75t_L g621 ( .A(n_475), .B(n_560), .Y(n_621) );
INVx2_ASAP7_75t_L g663 ( .A(n_475), .Y(n_663) );
AND2x2_ASAP7_75t_L g765 ( .A(n_475), .B(n_492), .Y(n_765) );
INVx1_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
NAND2xp5_ASAP7_75t_L g559 ( .A(n_476), .B(n_515), .Y(n_559) );
INVx2_ASAP7_75t_L g580 ( .A(n_476), .Y(n_580) );
AND2x4_ASAP7_75t_L g602 ( .A(n_476), .B(n_603), .Y(n_602) );
INVx1_ASAP7_75t_L g637 ( .A(n_476), .Y(n_637) );
AND2x2_ASAP7_75t_L g761 ( .A(n_476), .B(n_518), .Y(n_761) );
OR2x2_ASAP7_75t_L g476 ( .A(n_477), .B(n_485), .Y(n_476) );
AO21x2_ASAP7_75t_L g493 ( .A1(n_484), .A2(n_494), .B(n_500), .Y(n_493) );
AO21x2_ASAP7_75t_L g515 ( .A1(n_484), .A2(n_494), .B(n_500), .Y(n_515) );
OAI22xp5_ASAP7_75t_L g485 ( .A1(n_486), .A2(n_489), .B1(n_490), .B2(n_491), .Y(n_485) );
INVx1_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
INVx1_ASAP7_75t_L g735 ( .A(n_492), .Y(n_735) );
AND2x2_ASAP7_75t_L g492 ( .A(n_493), .B(n_501), .Y(n_492) );
NOR2xp67_ASAP7_75t_L g610 ( .A(n_493), .B(n_580), .Y(n_610) );
AND2x2_ASAP7_75t_L g615 ( .A(n_493), .B(n_580), .Y(n_615) );
INVx2_ASAP7_75t_L g628 ( .A(n_493), .Y(n_628) );
NOR2x1_ASAP7_75t_L g693 ( .A(n_493), .B(n_694), .Y(n_693) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_495), .B(n_496), .Y(n_494) );
AND2x4_ASAP7_75t_L g601 ( .A(n_501), .B(n_514), .Y(n_601) );
AND2x2_ASAP7_75t_L g616 ( .A(n_501), .B(n_617), .Y(n_616) );
INVx1_ASAP7_75t_L g671 ( .A(n_501), .Y(n_671) );
INVx2_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
NAND2xp5_ASAP7_75t_L g591 ( .A(n_502), .B(n_518), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g669 ( .A(n_502), .B(n_515), .Y(n_669) );
NAND2xp5_ASAP7_75t_SL g503 ( .A(n_504), .B(n_510), .Y(n_503) );
INVx1_ASAP7_75t_L g506 ( .A(n_507), .Y(n_506) );
INVxp33_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
NAND2x1p5_ASAP7_75t_L g513 ( .A(n_514), .B(n_516), .Y(n_513) );
INVx3_ASAP7_75t_L g577 ( .A(n_514), .Y(n_577) );
INVx3_ASAP7_75t_L g514 ( .A(n_515), .Y(n_514) );
HB1xp67_ASAP7_75t_L g575 ( .A(n_515), .Y(n_575) );
AND2x2_ASAP7_75t_L g689 ( .A(n_515), .B(n_690), .Y(n_689) );
INVx3_ASAP7_75t_L g632 ( .A(n_516), .Y(n_632) );
NAND2xp5_ASAP7_75t_L g712 ( .A(n_516), .B(n_671), .Y(n_712) );
BUFx3_ASAP7_75t_L g516 ( .A(n_517), .Y(n_516) );
AND2x2_ASAP7_75t_L g579 ( .A(n_517), .B(n_580), .Y(n_579) );
INVx1_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
AND2x4_ASAP7_75t_L g560 ( .A(n_518), .B(n_561), .Y(n_560) );
INVx2_ASAP7_75t_L g603 ( .A(n_518), .Y(n_603) );
INVxp67_ASAP7_75t_L g617 ( .A(n_518), .Y(n_617) );
HB1xp67_ASAP7_75t_L g690 ( .A(n_518), .Y(n_690) );
INVx1_ASAP7_75t_L g694 ( .A(n_518), .Y(n_694) );
INVx1_ASAP7_75t_L g672 ( .A(n_524), .Y(n_672) );
NOR2x1_ASAP7_75t_L g524 ( .A(n_525), .B(n_527), .Y(n_524) );
NOR2x1_ASAP7_75t_L g649 ( .A(n_525), .B(n_650), .Y(n_649) );
INVx1_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
AND2x2_ASAP7_75t_L g714 ( .A(n_526), .B(n_555), .Y(n_714) );
OR2x2_ASAP7_75t_L g766 ( .A(n_527), .B(n_767), .Y(n_766) );
INVx2_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
AND2x2_ASAP7_75t_L g665 ( .A(n_528), .B(n_666), .Y(n_665) );
AND2x2_ASAP7_75t_L g701 ( .A(n_528), .B(n_588), .Y(n_701) );
AND2x2_ASAP7_75t_L g528 ( .A(n_529), .B(n_540), .Y(n_528) );
AND2x4_ASAP7_75t_L g555 ( .A(n_529), .B(n_556), .Y(n_555) );
INVx1_ASAP7_75t_L g567 ( .A(n_529), .Y(n_567) );
INVx2_ASAP7_75t_L g584 ( .A(n_529), .Y(n_584) );
HB1xp67_ASAP7_75t_L g710 ( .A(n_529), .Y(n_710) );
AND2x2_ASAP7_75t_L g529 ( .A(n_530), .B(n_535), .Y(n_529) );
NOR3xp33_ASAP7_75t_L g531 ( .A(n_532), .B(n_533), .C(n_534), .Y(n_531) );
INVx3_ASAP7_75t_L g556 ( .A(n_540), .Y(n_556) );
INVx2_ASAP7_75t_L g650 ( .A(n_540), .Y(n_650) );
AND2x4_ASAP7_75t_L g540 ( .A(n_541), .B(n_542), .Y(n_540) );
OAI21xp5_ASAP7_75t_L g542 ( .A1(n_543), .A2(n_546), .B(n_551), .Y(n_542) );
OAI22xp5_ASAP7_75t_L g546 ( .A1(n_547), .A2(n_548), .B1(n_549), .B2(n_550), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g552 ( .A(n_553), .B(n_557), .Y(n_552) );
INVx2_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
NOR2xp33_ASAP7_75t_L g647 ( .A(n_554), .B(n_630), .Y(n_647) );
NOR2x1_ASAP7_75t_L g739 ( .A(n_554), .B(n_568), .Y(n_739) );
INVx4_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
NAND2xp5_ASAP7_75t_L g716 ( .A(n_555), .B(n_630), .Y(n_716) );
AND2x2_ASAP7_75t_L g583 ( .A(n_556), .B(n_584), .Y(n_583) );
INVx1_ASAP7_75t_L g597 ( .A(n_556), .Y(n_597) );
AOI22xp5_ASAP7_75t_SL g645 ( .A1(n_557), .A2(n_646), .B1(n_647), .B2(n_648), .Y(n_645) );
AND2x2_ASAP7_75t_L g557 ( .A(n_558), .B(n_560), .Y(n_557) );
NAND2x1p5_ASAP7_75t_L g642 ( .A(n_558), .B(n_616), .Y(n_642) );
INVx2_ASAP7_75t_SL g558 ( .A(n_559), .Y(n_558) );
OR2x2_ASAP7_75t_L g750 ( .A(n_559), .B(n_591), .Y(n_750) );
AND2x2_ASAP7_75t_L g573 ( .A(n_560), .B(n_574), .Y(n_573) );
AND2x4_ASAP7_75t_L g609 ( .A(n_560), .B(n_610), .Y(n_609) );
AND2x2_ASAP7_75t_L g752 ( .A(n_560), .B(n_663), .Y(n_752) );
INVx2_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
AND2x4_ASAP7_75t_L g627 ( .A(n_562), .B(n_628), .Y(n_627) );
INVx1_ASAP7_75t_L g653 ( .A(n_562), .Y(n_653) );
AND2x2_ASAP7_75t_L g688 ( .A(n_562), .B(n_580), .Y(n_688) );
OAI221xp5_ASAP7_75t_L g563 ( .A1(n_564), .A2(n_572), .B1(n_576), .B2(n_581), .C(n_586), .Y(n_563) );
INVx1_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
AND2x2_ASAP7_75t_L g565 ( .A(n_566), .B(n_569), .Y(n_565) );
INVx1_ASAP7_75t_L g644 ( .A(n_566), .Y(n_644) );
NAND2xp5_ASAP7_75t_L g707 ( .A(n_566), .B(n_640), .Y(n_707) );
NAND2xp5_ASAP7_75t_L g727 ( .A(n_566), .B(n_728), .Y(n_727) );
AND2x4_ASAP7_75t_L g566 ( .A(n_567), .B(n_568), .Y(n_566) );
NOR2xp67_ASAP7_75t_SL g612 ( .A(n_568), .B(n_613), .Y(n_612) );
HB1xp67_ASAP7_75t_L g625 ( .A(n_568), .Y(n_625) );
AND2x4_ASAP7_75t_SL g709 ( .A(n_568), .B(n_710), .Y(n_709) );
OR2x2_ASAP7_75t_L g756 ( .A(n_568), .B(n_757), .Y(n_756) );
HB1xp67_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
INVx3_ASAP7_75t_L g630 ( .A(n_570), .Y(n_630) );
INVx2_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
HB1xp67_ASAP7_75t_L g767 ( .A(n_571), .Y(n_767) );
INVx1_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
AOI221x1_ASAP7_75t_L g720 ( .A1(n_573), .A2(n_721), .B1(n_723), .B2(n_724), .C(n_726), .Y(n_720) );
AND2x2_ASAP7_75t_L g646 ( .A(n_574), .B(n_602), .Y(n_646) );
INVx1_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
OR2x2_ASAP7_75t_L g576 ( .A(n_577), .B(n_578), .Y(n_576) );
AND2x2_ASAP7_75t_L g589 ( .A(n_577), .B(n_590), .Y(n_589) );
NAND2xp5_ASAP7_75t_L g763 ( .A(n_577), .B(n_579), .Y(n_763) );
INVx2_ASAP7_75t_L g578 ( .A(n_579), .Y(n_578) );
INVx2_ASAP7_75t_L g581 ( .A(n_582), .Y(n_581) );
AND2x2_ASAP7_75t_L g582 ( .A(n_583), .B(n_585), .Y(n_582) );
AND2x2_ASAP7_75t_SL g587 ( .A(n_583), .B(n_588), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g613 ( .A(n_583), .B(n_596), .Y(n_613) );
INVx2_ASAP7_75t_L g620 ( .A(n_583), .Y(n_620) );
INVx1_ASAP7_75t_L g682 ( .A(n_584), .Y(n_682) );
BUFx2_ASAP7_75t_L g702 ( .A(n_585), .Y(n_702) );
NAND2xp33_ASAP7_75t_SL g586 ( .A(n_587), .B(n_589), .Y(n_586) );
OR2x6_ASAP7_75t_L g619 ( .A(n_588), .B(n_620), .Y(n_619) );
AND2x2_ASAP7_75t_L g748 ( .A(n_588), .B(n_640), .Y(n_748) );
INVx2_ASAP7_75t_L g590 ( .A(n_591), .Y(n_590) );
NAND2xp5_ASAP7_75t_L g592 ( .A(n_593), .B(n_611), .Y(n_592) );
AOI22xp5_ASAP7_75t_L g593 ( .A1(n_594), .A2(n_600), .B1(n_604), .B2(n_609), .Y(n_593) );
NOR2xp33_ASAP7_75t_L g594 ( .A(n_595), .B(n_598), .Y(n_594) );
AND2x2_ASAP7_75t_SL g657 ( .A(n_595), .B(n_599), .Y(n_657) );
AND2x4_ASAP7_75t_L g723 ( .A(n_595), .B(n_681), .Y(n_723) );
AND2x4_ASAP7_75t_SL g595 ( .A(n_596), .B(n_597), .Y(n_595) );
HB1xp67_ASAP7_75t_L g738 ( .A(n_596), .Y(n_738) );
INVx2_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
NOR2xp33_ASAP7_75t_L g638 ( .A(n_599), .B(n_639), .Y(n_638) );
HB1xp67_ASAP7_75t_L g691 ( .A(n_599), .Y(n_691) );
NAND2xp5_ASAP7_75t_L g722 ( .A(n_599), .B(n_630), .Y(n_722) );
AND2x2_ASAP7_75t_L g600 ( .A(n_601), .B(n_602), .Y(n_600) );
AND2x2_ASAP7_75t_L g743 ( .A(n_601), .B(n_662), .Y(n_743) );
INVx3_ASAP7_75t_L g654 ( .A(n_602), .Y(n_654) );
AND2x2_ASAP7_75t_L g675 ( .A(n_602), .B(n_627), .Y(n_675) );
NAND2x1_ASAP7_75t_SL g746 ( .A(n_602), .B(n_653), .Y(n_746) );
AND2x2_ASAP7_75t_L g604 ( .A(n_605), .B(n_606), .Y(n_604) );
INVx1_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
INVx1_ASAP7_75t_L g607 ( .A(n_608), .Y(n_607) );
AOI22xp5_ASAP7_75t_L g611 ( .A1(n_612), .A2(n_614), .B1(n_618), .B2(n_621), .Y(n_611) );
BUFx2_ASAP7_75t_L g667 ( .A(n_613), .Y(n_667) );
AOI22xp33_ASAP7_75t_L g713 ( .A1(n_614), .A2(n_705), .B1(n_714), .B2(n_715), .Y(n_713) );
AND2x2_ASAP7_75t_L g614 ( .A(n_615), .B(n_616), .Y(n_614) );
NAND2x1p5_ASAP7_75t_L g670 ( .A(n_615), .B(n_671), .Y(n_670) );
AND2x2_ASAP7_75t_L g635 ( .A(n_616), .B(n_636), .Y(n_635) );
INVx2_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
NAND3xp33_ASAP7_75t_L g699 ( .A(n_620), .B(n_700), .C(n_702), .Y(n_699) );
INVx1_ASAP7_75t_L g655 ( .A(n_621), .Y(n_655) );
AOI211x1_ASAP7_75t_L g622 ( .A1(n_623), .A2(n_631), .B(n_633), .C(n_651), .Y(n_622) );
INVx1_ASAP7_75t_L g623 ( .A(n_624), .Y(n_623) );
NAND2xp5_ASAP7_75t_L g624 ( .A(n_625), .B(n_626), .Y(n_624) );
NAND2xp5_ASAP7_75t_SL g733 ( .A(n_626), .B(n_714), .Y(n_733) );
AND2x2_ASAP7_75t_L g626 ( .A(n_627), .B(n_629), .Y(n_626) );
NAND2xp5_ASAP7_75t_L g661 ( .A(n_627), .B(n_662), .Y(n_661) );
AND2x2_ASAP7_75t_L g705 ( .A(n_627), .B(n_663), .Y(n_705) );
AND2x2_ASAP7_75t_L g760 ( .A(n_627), .B(n_761), .Y(n_760) );
INVx1_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
INVx1_ASAP7_75t_L g683 ( .A(n_630), .Y(n_683) );
INVx1_ASAP7_75t_L g631 ( .A(n_632), .Y(n_631) );
OR2x2_ASAP7_75t_L g725 ( .A(n_632), .B(n_670), .Y(n_725) );
NAND2xp5_ASAP7_75t_L g633 ( .A(n_634), .B(n_645), .Y(n_633) );
AOI22xp5_ASAP7_75t_SL g634 ( .A1(n_635), .A2(n_638), .B1(n_641), .B2(n_643), .Y(n_634) );
BUFx2_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
AND2x2_ASAP7_75t_L g698 ( .A(n_637), .B(n_693), .Y(n_698) );
INVx1_ASAP7_75t_SL g740 ( .A(n_637), .Y(n_740) );
INVx1_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
AND2x2_ASAP7_75t_SL g708 ( .A(n_640), .B(n_709), .Y(n_708) );
INVx3_ASAP7_75t_L g641 ( .A(n_642), .Y(n_641) );
INVxp67_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
HB1xp67_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
AND2x2_ASAP7_75t_L g744 ( .A(n_649), .B(n_666), .Y(n_744) );
AOI21xp5_ASAP7_75t_L g651 ( .A1(n_652), .A2(n_655), .B(n_656), .Y(n_651) );
OR2x2_ASAP7_75t_L g652 ( .A(n_653), .B(n_654), .Y(n_652) );
NAND2xp5_ASAP7_75t_L g697 ( .A(n_653), .B(n_698), .Y(n_697) );
OR2x2_ASAP7_75t_L g668 ( .A(n_654), .B(n_669), .Y(n_668) );
INVx1_ASAP7_75t_SL g656 ( .A(n_657), .Y(n_656) );
INVxp67_ASAP7_75t_SL g816 ( .A(n_658), .Y(n_816) );
NAND3x1_ASAP7_75t_L g658 ( .A(n_659), .B(n_695), .C(n_703), .Y(n_658) );
NAND4xp25_ASAP7_75t_L g769 ( .A(n_659), .B(n_695), .C(n_703), .D(n_770), .Y(n_769) );
NOR2x1_ASAP7_75t_L g659 ( .A(n_660), .B(n_673), .Y(n_659) );
OAI222xp33_ASAP7_75t_L g660 ( .A1(n_661), .A2(n_664), .B1(n_667), .B2(n_668), .C1(n_670), .C2(n_672), .Y(n_660) );
INVx1_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
INVx1_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
OAI21xp5_ASAP7_75t_SL g747 ( .A1(n_665), .A2(n_748), .B(n_749), .Y(n_747) );
NAND2xp5_ASAP7_75t_SL g730 ( .A(n_666), .B(n_681), .Y(n_730) );
OAI22xp5_ASAP7_75t_L g726 ( .A1(n_669), .A2(n_727), .B1(n_729), .B2(n_730), .Y(n_726) );
NAND2xp5_ASAP7_75t_L g673 ( .A(n_674), .B(n_684), .Y(n_673) );
NAND2xp5_ASAP7_75t_SL g674 ( .A(n_675), .B(n_676), .Y(n_674) );
NAND2xp5_ASAP7_75t_L g676 ( .A(n_677), .B(n_679), .Y(n_676) );
NAND2xp5_ASAP7_75t_L g685 ( .A(n_677), .B(n_686), .Y(n_685) );
INVx1_ASAP7_75t_L g677 ( .A(n_678), .Y(n_677) );
NAND2xp5_ASAP7_75t_L g679 ( .A(n_680), .B(n_683), .Y(n_679) );
INVx2_ASAP7_75t_SL g680 ( .A(n_681), .Y(n_680) );
NAND2xp5_ASAP7_75t_L g686 ( .A(n_681), .B(n_683), .Y(n_686) );
INVx2_ASAP7_75t_L g681 ( .A(n_682), .Y(n_681) );
AOI22xp5_ASAP7_75t_L g684 ( .A1(n_685), .A2(n_687), .B1(n_691), .B2(n_692), .Y(n_684) );
AND2x4_ASAP7_75t_L g687 ( .A(n_688), .B(n_689), .Y(n_687) );
AND2x2_ASAP7_75t_L g692 ( .A(n_688), .B(n_693), .Y(n_692) );
NAND2xp5_ASAP7_75t_SL g695 ( .A(n_696), .B(n_699), .Y(n_695) );
INVx1_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
INVx1_ASAP7_75t_L g729 ( .A(n_698), .Y(n_729) );
INVx1_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
AND2x2_ASAP7_75t_L g703 ( .A(n_704), .B(n_713), .Y(n_703) );
AOI22xp5_ASAP7_75t_SL g704 ( .A1(n_705), .A2(n_706), .B1(n_708), .B2(n_711), .Y(n_704) );
INVx1_ASAP7_75t_L g706 ( .A(n_707), .Y(n_706) );
INVxp67_ASAP7_75t_L g711 ( .A(n_712), .Y(n_711) );
INVx1_ASAP7_75t_L g715 ( .A(n_716), .Y(n_715) );
NAND2xp33_ASAP7_75t_L g718 ( .A(n_717), .B(n_719), .Y(n_718) );
INVx1_ASAP7_75t_L g815 ( .A(n_719), .Y(n_815) );
NAND3x1_ASAP7_75t_L g719 ( .A(n_720), .B(n_731), .C(n_751), .Y(n_719) );
INVx1_ASAP7_75t_L g721 ( .A(n_722), .Y(n_721) );
AOI22xp5_ASAP7_75t_L g742 ( .A1(n_723), .A2(n_743), .B1(n_744), .B2(n_745), .Y(n_742) );
INVx1_ASAP7_75t_L g724 ( .A(n_725), .Y(n_724) );
INVx1_ASAP7_75t_SL g757 ( .A(n_728), .Y(n_757) );
NOR2x1_ASAP7_75t_L g731 ( .A(n_732), .B(n_741), .Y(n_731) );
AOI21xp5_ASAP7_75t_SL g732 ( .A1(n_733), .A2(n_734), .B(n_740), .Y(n_732) );
NAND2xp5_ASAP7_75t_L g734 ( .A(n_735), .B(n_736), .Y(n_734) );
INVx1_ASAP7_75t_L g736 ( .A(n_737), .Y(n_736) );
NAND2xp5_ASAP7_75t_L g737 ( .A(n_738), .B(n_739), .Y(n_737) );
NAND2xp5_ASAP7_75t_L g741 ( .A(n_742), .B(n_747), .Y(n_741) );
INVx2_ASAP7_75t_SL g745 ( .A(n_746), .Y(n_745) );
NAND2xp5_ASAP7_75t_L g758 ( .A(n_746), .B(n_759), .Y(n_758) );
INVx1_ASAP7_75t_SL g749 ( .A(n_750), .Y(n_749) );
AOI221xp5_ASAP7_75t_L g751 ( .A1(n_752), .A2(n_753), .B1(n_755), .B2(n_758), .C(n_762), .Y(n_751) );
INVx1_ASAP7_75t_L g753 ( .A(n_754), .Y(n_753) );
INVxp67_ASAP7_75t_L g755 ( .A(n_756), .Y(n_755) );
INVx2_ASAP7_75t_L g759 ( .A(n_760), .Y(n_759) );
AOI21xp5_ASAP7_75t_L g762 ( .A1(n_763), .A2(n_764), .B(n_766), .Y(n_762) );
INVx1_ASAP7_75t_L g764 ( .A(n_765), .Y(n_764) );
NOR2xp33_ASAP7_75t_L g770 ( .A(n_771), .B(n_772), .Y(n_770) );
INVxp67_ASAP7_75t_L g773 ( .A(n_774), .Y(n_773) );
NOR3xp33_ASAP7_75t_L g817 ( .A(n_774), .B(n_818), .C(n_819), .Y(n_817) );
NAND2xp5_ASAP7_75t_L g774 ( .A(n_775), .B(n_785), .Y(n_774) );
INVxp33_ASAP7_75t_L g792 ( .A(n_775), .Y(n_792) );
NOR2xp33_ASAP7_75t_L g775 ( .A(n_776), .B(n_778), .Y(n_775) );
CKINVDCx8_ASAP7_75t_R g776 ( .A(n_777), .Y(n_776) );
NOR2xp33_ASAP7_75t_L g778 ( .A(n_779), .B(n_780), .Y(n_778) );
CKINVDCx5p33_ASAP7_75t_R g789 ( .A(n_781), .Y(n_789) );
OAI32xp33_ASAP7_75t_L g790 ( .A1(n_781), .A2(n_791), .A3(n_792), .B1(n_793), .B2(n_834), .Y(n_790) );
INVx1_ASAP7_75t_L g824 ( .A(n_782), .Y(n_824) );
NAND2xp5_ASAP7_75t_L g782 ( .A(n_783), .B(n_784), .Y(n_782) );
CKINVDCx20_ASAP7_75t_R g791 ( .A(n_785), .Y(n_791) );
INVx1_ASAP7_75t_SL g786 ( .A(n_787), .Y(n_786) );
BUFx2_ASAP7_75t_L g787 ( .A(n_788), .Y(n_787) );
NOR2x1_ASAP7_75t_R g794 ( .A(n_788), .B(n_795), .Y(n_794) );
NOR2xp33_ASAP7_75t_L g797 ( .A(n_791), .B(n_798), .Y(n_797) );
INVx1_ASAP7_75t_L g793 ( .A(n_794), .Y(n_793) );
HB1xp67_ASAP7_75t_L g802 ( .A(n_795), .Y(n_802) );
AOI21xp5_ASAP7_75t_L g796 ( .A1(n_797), .A2(n_803), .B(n_817), .Y(n_796) );
HB1xp67_ASAP7_75t_L g798 ( .A(n_799), .Y(n_798) );
CKINVDCx5p33_ASAP7_75t_R g799 ( .A(n_800), .Y(n_799) );
BUFx3_ASAP7_75t_L g800 ( .A(n_801), .Y(n_800) );
CKINVDCx20_ASAP7_75t_R g801 ( .A(n_802), .Y(n_801) );
AOI22xp33_ASAP7_75t_SL g804 ( .A1(n_805), .A2(n_806), .B1(n_812), .B2(n_813), .Y(n_804) );
INVx1_ASAP7_75t_L g805 ( .A(n_806), .Y(n_805) );
OAI22xp5_ASAP7_75t_L g806 ( .A1(n_807), .A2(n_808), .B1(n_810), .B2(n_811), .Y(n_806) );
INVx1_ASAP7_75t_L g807 ( .A(n_808), .Y(n_807) );
CKINVDCx5p33_ASAP7_75t_R g810 ( .A(n_811), .Y(n_810) );
INVx1_ASAP7_75t_L g812 ( .A(n_813), .Y(n_812) );
AND3x2_ASAP7_75t_L g813 ( .A(n_814), .B(n_815), .C(n_816), .Y(n_813) );
BUFx4f_ASAP7_75t_SL g820 ( .A(n_821), .Y(n_820) );
INVx1_ASAP7_75t_L g821 ( .A(n_822), .Y(n_821) );
INVx1_ASAP7_75t_SL g831 ( .A(n_822), .Y(n_831) );
CKINVDCx5p33_ASAP7_75t_R g822 ( .A(n_823), .Y(n_822) );
AND2x2_ASAP7_75t_SL g823 ( .A(n_824), .B(n_825), .Y(n_823) );
INVx2_ASAP7_75t_L g826 ( .A(n_827), .Y(n_826) );
INVx4_ASAP7_75t_SL g829 ( .A(n_830), .Y(n_829) );
BUFx4f_ASAP7_75t_SL g830 ( .A(n_831), .Y(n_830) );
endmodule