module fake_ariane_332_n_259 (n_8, n_56, n_60, n_64, n_38, n_47, n_18, n_75, n_67, n_34, n_69, n_74, n_33, n_19, n_40, n_12, n_53, n_21, n_66, n_71, n_24, n_7, n_49, n_20, n_17, n_50, n_62, n_51, n_76, n_79, n_26, n_3, n_46, n_0, n_36, n_72, n_44, n_30, n_31, n_42, n_57, n_70, n_10, n_6, n_48, n_4, n_2, n_32, n_37, n_58, n_65, n_9, n_45, n_11, n_52, n_73, n_77, n_15, n_23, n_61, n_22, n_43, n_1, n_13, n_27, n_29, n_41, n_55, n_28, n_80, n_14, n_68, n_78, n_39, n_59, n_63, n_16, n_5, n_35, n_54, n_25, n_259);

input n_8;
input n_56;
input n_60;
input n_64;
input n_38;
input n_47;
input n_18;
input n_75;
input n_67;
input n_34;
input n_69;
input n_74;
input n_33;
input n_19;
input n_40;
input n_12;
input n_53;
input n_21;
input n_66;
input n_71;
input n_24;
input n_7;
input n_49;
input n_20;
input n_17;
input n_50;
input n_62;
input n_51;
input n_76;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_36;
input n_72;
input n_44;
input n_30;
input n_31;
input n_42;
input n_57;
input n_70;
input n_10;
input n_6;
input n_48;
input n_4;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_9;
input n_45;
input n_11;
input n_52;
input n_73;
input n_77;
input n_15;
input n_23;
input n_61;
input n_22;
input n_43;
input n_1;
input n_13;
input n_27;
input n_29;
input n_41;
input n_55;
input n_28;
input n_80;
input n_14;
input n_68;
input n_78;
input n_39;
input n_59;
input n_63;
input n_16;
input n_5;
input n_35;
input n_54;
input n_25;

output n_259;

wire n_83;
wire n_233;
wire n_170;
wire n_190;
wire n_160;
wire n_179;
wire n_180;
wire n_119;
wire n_124;
wire n_167;
wire n_90;
wire n_195;
wire n_213;
wire n_110;
wire n_153;
wire n_197;
wire n_221;
wire n_86;
wire n_89;
wire n_176;
wire n_149;
wire n_158;
wire n_237;
wire n_172;
wire n_95;
wire n_175;
wire n_92;
wire n_143;
wire n_183;
wire n_203;
wire n_150;
wire n_98;
wire n_113;
wire n_114;
wire n_181;
wire n_152;
wire n_120;
wire n_169;
wire n_106;
wire n_173;
wire n_111;
wire n_242;
wire n_115;
wire n_133;
wire n_205;
wire n_236;
wire n_109;
wire n_208;
wire n_245;
wire n_96;
wire n_156;
wire n_209;
wire n_174;
wire n_100;
wire n_187;
wire n_132;
wire n_225;
wire n_210;
wire n_147;
wire n_204;
wire n_235;
wire n_200;
wire n_166;
wire n_253;
wire n_218;
wire n_103;
wire n_244;
wire n_226;
wire n_246;
wire n_220;
wire n_84;
wire n_247;
wire n_199;
wire n_91;
wire n_159;
wire n_107;
wire n_189;
wire n_128;
wire n_105;
wire n_217;
wire n_240;
wire n_82;
wire n_178;
wire n_224;
wire n_131;
wire n_201;
wire n_229;
wire n_250;
wire n_222;
wire n_117;
wire n_139;
wire n_165;
wire n_85;
wire n_130;
wire n_144;
wire n_256;
wire n_214;
wire n_227;
wire n_94;
wire n_101;
wire n_243;
wire n_134;
wire n_188;
wire n_185;
wire n_249;
wire n_212;
wire n_123;
wire n_138;
wire n_112;
wire n_162;
wire n_129;
wire n_126;
wire n_137;
wire n_255;
wire n_122;
wire n_257;
wire n_198;
wire n_148;
wire n_232;
wire n_164;
wire n_157;
wire n_248;
wire n_184;
wire n_177;
wire n_135;
wire n_258;
wire n_171;
wire n_228;
wire n_118;
wire n_121;
wire n_93;
wire n_108;
wire n_102;
wire n_182;
wire n_196;
wire n_125;
wire n_168;
wire n_81;
wire n_87;
wire n_206;
wire n_207;
wire n_241;
wire n_254;
wire n_238;
wire n_219;
wire n_140;
wire n_191;
wire n_151;
wire n_136;
wire n_231;
wire n_192;
wire n_146;
wire n_234;
wire n_230;
wire n_211;
wire n_194;
wire n_97;
wire n_154;
wire n_215;
wire n_252;
wire n_142;
wire n_251;
wire n_161;
wire n_163;
wire n_88;
wire n_186;
wire n_141;
wire n_116;
wire n_104;
wire n_202;
wire n_145;
wire n_193;
wire n_99;
wire n_216;
wire n_155;
wire n_127;
wire n_239;
wire n_223;

INVx1_ASAP7_75t_L g81 ( 
.A(n_38),
.Y(n_81)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_42),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_66),
.Y(n_83)
);

CKINVDCx5p33_ASAP7_75t_R g84 ( 
.A(n_80),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_61),
.Y(n_85)
);

HB1xp67_ASAP7_75t_L g86 ( 
.A(n_12),
.Y(n_86)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_74),
.Y(n_87)
);

INVxp67_ASAP7_75t_SL g88 ( 
.A(n_59),
.Y(n_88)
);

CKINVDCx5p33_ASAP7_75t_R g89 ( 
.A(n_64),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_6),
.Y(n_90)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_28),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_16),
.Y(n_92)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_70),
.Y(n_93)
);

CKINVDCx5p33_ASAP7_75t_R g94 ( 
.A(n_18),
.Y(n_94)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_35),
.Y(n_95)
);

BUFx3_ASAP7_75t_L g96 ( 
.A(n_27),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_45),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_32),
.Y(n_98)
);

INVxp33_ASAP7_75t_L g99 ( 
.A(n_17),
.Y(n_99)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_77),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_72),
.B(n_55),
.Y(n_101)
);

INVx1_ASAP7_75t_SL g102 ( 
.A(n_1),
.Y(n_102)
);

BUFx3_ASAP7_75t_L g103 ( 
.A(n_13),
.Y(n_103)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_33),
.Y(n_104)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_73),
.Y(n_105)
);

CKINVDCx5p33_ASAP7_75t_R g106 ( 
.A(n_56),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_4),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_3),
.Y(n_108)
);

INVxp67_ASAP7_75t_SL g109 ( 
.A(n_34),
.Y(n_109)
);

INVx2_ASAP7_75t_SL g110 ( 
.A(n_3),
.Y(n_110)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_37),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_31),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_14),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_50),
.Y(n_114)
);

INVxp67_ASAP7_75t_SL g115 ( 
.A(n_46),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_0),
.Y(n_116)
);

CKINVDCx5p33_ASAP7_75t_R g117 ( 
.A(n_58),
.Y(n_117)
);

CKINVDCx16_ASAP7_75t_R g118 ( 
.A(n_78),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_49),
.Y(n_119)
);

CKINVDCx5p33_ASAP7_75t_R g120 ( 
.A(n_63),
.Y(n_120)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_107),
.Y(n_121)
);

AND2x4_ASAP7_75t_L g122 ( 
.A(n_110),
.B(n_0),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_108),
.Y(n_123)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_116),
.Y(n_124)
);

BUFx2_ASAP7_75t_L g125 ( 
.A(n_102),
.Y(n_125)
);

HB1xp67_ASAP7_75t_L g126 ( 
.A(n_86),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_96),
.Y(n_127)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_103),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_81),
.Y(n_129)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_82),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_83),
.B(n_1),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_85),
.Y(n_132)
);

NOR2x1_ASAP7_75t_L g133 ( 
.A(n_90),
.B(n_44),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_91),
.B(n_2),
.Y(n_134)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_118),
.Y(n_135)
);

BUFx2_ASAP7_75t_L g136 ( 
.A(n_112),
.Y(n_136)
);

HB1xp67_ASAP7_75t_L g137 ( 
.A(n_125),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_126),
.A2(n_113),
.B1(n_119),
.B2(n_115),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_124),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_135),
.B(n_99),
.Y(n_140)
);

AND2x4_ASAP7_75t_L g141 ( 
.A(n_128),
.B(n_88),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_127),
.B(n_97),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_127),
.Y(n_143)
);

BUFx3_ASAP7_75t_L g144 ( 
.A(n_132),
.Y(n_144)
);

BUFx10_ASAP7_75t_L g145 ( 
.A(n_122),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_124),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_131),
.B(n_134),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_129),
.B(n_92),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_121),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_123),
.Y(n_150)
);

BUFx3_ASAP7_75t_L g151 ( 
.A(n_132),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_130),
.B(n_98),
.Y(n_152)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_123),
.Y(n_153)
);

AND2x6_ASAP7_75t_L g154 ( 
.A(n_133),
.B(n_100),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_136),
.Y(n_155)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_153),
.Y(n_156)
);

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_137),
.Y(n_157)
);

NAND2x1p5_ASAP7_75t_L g158 ( 
.A(n_144),
.B(n_136),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_139),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g160 ( 
.A(n_150),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_145),
.B(n_114),
.Y(n_161)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_149),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_146),
.Y(n_163)
);

AND3x1_ASAP7_75t_SL g164 ( 
.A(n_155),
.B(n_2),
.C(n_4),
.Y(n_164)
);

INVx1_ASAP7_75t_SL g165 ( 
.A(n_151),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_152),
.Y(n_166)
);

INVx5_ASAP7_75t_L g167 ( 
.A(n_143),
.Y(n_167)
);

O2A1O1Ixp33_ASAP7_75t_L g168 ( 
.A1(n_147),
.A2(n_109),
.B(n_105),
.C(n_111),
.Y(n_168)
);

HB1xp67_ASAP7_75t_L g169 ( 
.A(n_141),
.Y(n_169)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_150),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_138),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_141),
.B(n_84),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_142),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_150),
.Y(n_174)
);

NAND2x1p5_ASAP7_75t_L g175 ( 
.A(n_143),
.B(n_104),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_148),
.B(n_89),
.Y(n_176)
);

NOR2x1p5_ASAP7_75t_L g177 ( 
.A(n_140),
.B(n_94),
.Y(n_177)
);

INVx4_ASAP7_75t_L g178 ( 
.A(n_154),
.Y(n_178)
);

AND2x4_ASAP7_75t_L g179 ( 
.A(n_178),
.B(n_154),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g180 ( 
.A(n_160),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_157),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_166),
.B(n_106),
.Y(n_182)
);

INVx4_ASAP7_75t_L g183 ( 
.A(n_160),
.Y(n_183)
);

INVx3_ASAP7_75t_L g184 ( 
.A(n_160),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_L g185 ( 
.A1(n_163),
.A2(n_101),
.B(n_95),
.Y(n_185)
);

HB1xp67_ASAP7_75t_L g186 ( 
.A(n_169),
.Y(n_186)
);

BUFx2_ASAP7_75t_L g187 ( 
.A(n_158),
.Y(n_187)
);

INVx4_ASAP7_75t_L g188 ( 
.A(n_167),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_161),
.B(n_120),
.Y(n_189)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_162),
.Y(n_190)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_156),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_171),
.A2(n_117),
.B1(n_93),
.B2(n_87),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_173),
.B(n_79),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_159),
.Y(n_194)
);

A2O1A1Ixp33_ASAP7_75t_L g195 ( 
.A1(n_168),
.A2(n_5),
.B(n_7),
.C(n_8),
.Y(n_195)
);

AOI21xp5_ASAP7_75t_L g196 ( 
.A1(n_172),
.A2(n_9),
.B(n_10),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_174),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_176),
.B(n_76),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_170),
.Y(n_199)
);

OAI21x1_ASAP7_75t_L g200 ( 
.A1(n_193),
.A2(n_175),
.B(n_177),
.Y(n_200)
);

BUFx2_ASAP7_75t_L g201 ( 
.A(n_181),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_194),
.Y(n_202)
);

AO21x2_ASAP7_75t_L g203 ( 
.A1(n_185),
.A2(n_198),
.B(n_196),
.Y(n_203)
);

NOR2xp67_ASAP7_75t_L g204 ( 
.A(n_183),
.B(n_188),
.Y(n_204)
);

OAI21x1_ASAP7_75t_L g205 ( 
.A1(n_184),
.A2(n_167),
.B(n_164),
.Y(n_205)
);

A2O1A1Ixp33_ASAP7_75t_L g206 ( 
.A1(n_189),
.A2(n_165),
.B(n_167),
.C(n_19),
.Y(n_206)
);

INVx8_ASAP7_75t_L g207 ( 
.A(n_179),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_182),
.A2(n_11),
.B1(n_15),
.B2(n_20),
.Y(n_208)
);

BUFx4_ASAP7_75t_SL g209 ( 
.A(n_187),
.Y(n_209)
);

OAI21x1_ASAP7_75t_L g210 ( 
.A1(n_184),
.A2(n_21),
.B(n_22),
.Y(n_210)
);

OA21x2_ASAP7_75t_L g211 ( 
.A1(n_199),
.A2(n_23),
.B(n_24),
.Y(n_211)
);

OAI21x1_ASAP7_75t_L g212 ( 
.A1(n_199),
.A2(n_25),
.B(n_26),
.Y(n_212)
);

OAI21x1_ASAP7_75t_L g213 ( 
.A1(n_197),
.A2(n_29),
.B(n_30),
.Y(n_213)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_190),
.Y(n_214)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_191),
.Y(n_215)
);

AOI22xp33_ASAP7_75t_L g216 ( 
.A1(n_214),
.A2(n_192),
.B1(n_186),
.B2(n_179),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_202),
.Y(n_217)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_215),
.Y(n_218)
);

AOI22xp33_ASAP7_75t_SL g219 ( 
.A1(n_201),
.A2(n_207),
.B1(n_208),
.B2(n_205),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_200),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_206),
.A2(n_195),
.B1(n_180),
.B2(n_188),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_207),
.B(n_180),
.Y(n_222)
);

AOI21xp5_ASAP7_75t_L g223 ( 
.A1(n_203),
.A2(n_36),
.B(n_39),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_204),
.B(n_40),
.Y(n_224)
);

BUFx6f_ASAP7_75t_L g225 ( 
.A(n_222),
.Y(n_225)
);

OR2x2_ASAP7_75t_L g226 ( 
.A(n_217),
.B(n_209),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_218),
.Y(n_227)
);

AND2x2_ASAP7_75t_L g228 ( 
.A(n_216),
.B(n_209),
.Y(n_228)
);

INVxp67_ASAP7_75t_SL g229 ( 
.A(n_220),
.Y(n_229)
);

AND2x2_ASAP7_75t_L g230 ( 
.A(n_219),
.B(n_208),
.Y(n_230)
);

AND2x2_ASAP7_75t_L g231 ( 
.A(n_228),
.B(n_211),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_227),
.Y(n_232)
);

AND2x2_ASAP7_75t_L g233 ( 
.A(n_226),
.B(n_211),
.Y(n_233)
);

AND2x2_ASAP7_75t_L g234 ( 
.A(n_230),
.B(n_203),
.Y(n_234)
);

OR2x2_ASAP7_75t_L g235 ( 
.A(n_225),
.B(n_221),
.Y(n_235)
);

OAI21xp5_ASAP7_75t_L g236 ( 
.A1(n_229),
.A2(n_221),
.B(n_223),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_225),
.Y(n_237)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_232),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_234),
.Y(n_239)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_237),
.Y(n_240)
);

AND2x4_ASAP7_75t_SL g241 ( 
.A(n_233),
.B(n_231),
.Y(n_241)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_235),
.Y(n_242)
);

AND2x2_ASAP7_75t_L g243 ( 
.A(n_236),
.B(n_213),
.Y(n_243)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_238),
.Y(n_244)
);

AND2x4_ASAP7_75t_L g245 ( 
.A(n_242),
.B(n_236),
.Y(n_245)
);

AND2x2_ASAP7_75t_L g246 ( 
.A(n_241),
.B(n_210),
.Y(n_246)
);

AND2x2_ASAP7_75t_L g247 ( 
.A(n_239),
.B(n_212),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_244),
.Y(n_248)
);

AOI322xp5_ASAP7_75t_L g249 ( 
.A1(n_248),
.A2(n_245),
.A3(n_243),
.B1(n_247),
.B2(n_240),
.C1(n_246),
.C2(n_224),
.Y(n_249)
);

OAI21xp33_ASAP7_75t_L g250 ( 
.A1(n_249),
.A2(n_41),
.B(n_43),
.Y(n_250)
);

AOI211xp5_ASAP7_75t_L g251 ( 
.A1(n_250),
.A2(n_75),
.B(n_47),
.C(n_48),
.Y(n_251)
);

NAND2xp33_ASAP7_75t_SL g252 ( 
.A(n_251),
.B(n_51),
.Y(n_252)
);

AOI211xp5_ASAP7_75t_L g253 ( 
.A1(n_252),
.A2(n_52),
.B(n_53),
.C(n_54),
.Y(n_253)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_253),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_254),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_255),
.Y(n_256)
);

AOI21xp5_ASAP7_75t_L g257 ( 
.A1(n_256),
.A2(n_57),
.B(n_60),
.Y(n_257)
);

AOI21xp5_ASAP7_75t_L g258 ( 
.A1(n_257),
.A2(n_62),
.B(n_65),
.Y(n_258)
);

AOI221xp5_ASAP7_75t_L g259 ( 
.A1(n_258),
.A2(n_67),
.B1(n_68),
.B2(n_69),
.C(n_71),
.Y(n_259)
);


endmodule