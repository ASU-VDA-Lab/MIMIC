module fake_jpeg_28572_n_117 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_117);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_117;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_93;
wire n_91;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_43;
wire n_100;
wire n_82;
wire n_96;

INVx13_ASAP7_75t_L g38 ( 
.A(n_27),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_35),
.Y(n_39)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_9),
.Y(n_40)
);

BUFx4f_ASAP7_75t_L g41 ( 
.A(n_8),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_21),
.B(n_6),
.Y(n_42)
);

BUFx12_ASAP7_75t_L g43 ( 
.A(n_20),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_13),
.B(n_23),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_37),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_2),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_16),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_10),
.B(n_18),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_6),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_42),
.B(n_0),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_50),
.B(n_42),
.Y(n_58)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_41),
.Y(n_51)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_51),
.Y(n_65)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_52),
.Y(n_67)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_41),
.Y(n_53)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_53),
.Y(n_68)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

CKINVDCx6p67_ASAP7_75t_R g59 ( 
.A(n_54),
.Y(n_59)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_49),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_55),
.B(n_46),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_L g56 ( 
.A1(n_41),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_56),
.A2(n_39),
.B1(n_3),
.B2(n_4),
.Y(n_66)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_57),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_58),
.B(n_63),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_60),
.B(n_61),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_50),
.B(n_44),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_55),
.B(n_48),
.Y(n_63)
);

OAI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_51),
.A2(n_47),
.B1(n_45),
.B2(n_39),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_64),
.A2(n_53),
.B1(n_52),
.B2(n_39),
.Y(n_71)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_66),
.B(n_69),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_57),
.B(n_43),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_54),
.B(n_43),
.Y(n_70)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_70),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_71),
.A2(n_62),
.B1(n_9),
.B2(n_8),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_SL g73 ( 
.A1(n_64),
.A2(n_38),
.B(n_43),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_73),
.B(n_80),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_65),
.A2(n_19),
.B1(n_34),
.B2(n_33),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_76),
.A2(n_77),
.B1(n_36),
.B2(n_14),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_68),
.A2(n_17),
.B1(n_32),
.B2(n_31),
.Y(n_77)
);

INVxp67_ASAP7_75t_L g78 ( 
.A(n_59),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_78),
.B(n_83),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_L g79 ( 
.A1(n_59),
.A2(n_1),
.B(n_3),
.Y(n_79)
);

OR2x2_ASAP7_75t_L g87 ( 
.A(n_79),
.B(n_5),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_59),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_68),
.Y(n_81)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_81),
.Y(n_95)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_67),
.Y(n_82)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_82),
.Y(n_96)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_67),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_72),
.A2(n_62),
.B1(n_5),
.B2(n_7),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_85),
.A2(n_92),
.B1(n_94),
.B2(n_15),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_84),
.B(n_4),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_86),
.B(n_89),
.Y(n_99)
);

AOI21xp5_ASAP7_75t_L g100 ( 
.A1(n_87),
.A2(n_93),
.B(n_78),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_75),
.B(n_7),
.Y(n_89)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_79),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_91),
.B(n_97),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_72),
.B(n_11),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_74),
.B(n_12),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_100),
.B(n_101),
.Y(n_108)
);

HB1xp67_ASAP7_75t_L g101 ( 
.A(n_96),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_93),
.B(n_83),
.C(n_22),
.Y(n_102)
);

XNOR2xp5_ASAP7_75t_L g107 ( 
.A(n_102),
.B(n_92),
.Y(n_107)
);

BUFx4f_ASAP7_75t_SL g103 ( 
.A(n_88),
.Y(n_103)
);

BUFx2_ASAP7_75t_L g106 ( 
.A(n_103),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_91),
.B(n_90),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_L g109 ( 
.A1(n_104),
.A2(n_105),
.B(n_87),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_L g111 ( 
.A(n_107),
.B(n_109),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_108),
.B(n_98),
.C(n_99),
.Y(n_110)
);

XOR2xp5_ASAP7_75t_L g113 ( 
.A(n_110),
.B(n_112),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_106),
.B(n_98),
.C(n_103),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_113),
.A2(n_111),
.B1(n_95),
.B2(n_26),
.Y(n_114)
);

BUFx24_ASAP7_75t_SL g115 ( 
.A(n_114),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_115),
.A2(n_24),
.B1(n_25),
.B2(n_28),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_L g117 ( 
.A1(n_116),
.A2(n_29),
.B(n_30),
.Y(n_117)
);


endmodule