module fake_jpeg_11150_n_536 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_536);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_536;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_511;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

INVx3_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

INVx5_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_13),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_17),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_14),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_17),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_13),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_14),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_4),
.Y(n_37)
);

BUFx12_ASAP7_75t_L g38 ( 
.A(n_6),
.Y(n_38)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_8),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_13),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_14),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_1),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_16),
.Y(n_43)
);

BUFx16f_ASAP7_75t_L g44 ( 
.A(n_11),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_18),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_2),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_10),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_17),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_10),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_15),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_16),
.Y(n_51)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_9),
.Y(n_52)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_48),
.Y(n_53)
);

HB1xp67_ASAP7_75t_L g124 ( 
.A(n_53),
.Y(n_124)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_24),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g122 ( 
.A(n_54),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_19),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_55),
.Y(n_134)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_24),
.Y(n_56)
);

INVx5_ASAP7_75t_L g110 ( 
.A(n_56),
.Y(n_110)
);

INVx11_ASAP7_75t_L g57 ( 
.A(n_44),
.Y(n_57)
);

INVx5_ASAP7_75t_SL g117 ( 
.A(n_57),
.Y(n_117)
);

INVx1_ASAP7_75t_SL g58 ( 
.A(n_31),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g112 ( 
.A(n_58),
.B(n_90),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_19),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_59),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_19),
.Y(n_60)
);

INVx6_ASAP7_75t_L g115 ( 
.A(n_60),
.Y(n_115)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_24),
.Y(n_61)
);

INVx5_ASAP7_75t_L g151 ( 
.A(n_61),
.Y(n_151)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_37),
.Y(n_62)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_62),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_45),
.B(n_18),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_63),
.B(n_67),
.Y(n_147)
);

BUFx5_ASAP7_75t_L g64 ( 
.A(n_19),
.Y(n_64)
);

INVx4_ASAP7_75t_L g120 ( 
.A(n_64),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_22),
.Y(n_65)
);

INVx6_ASAP7_75t_L g125 ( 
.A(n_65),
.Y(n_125)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_48),
.Y(n_66)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_66),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_45),
.B(n_18),
.Y(n_67)
);

CKINVDCx6p67_ASAP7_75t_R g68 ( 
.A(n_48),
.Y(n_68)
);

INVx4_ASAP7_75t_SL g114 ( 
.A(n_68),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_31),
.B(n_28),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_69),
.B(n_77),
.Y(n_106)
);

INVx11_ASAP7_75t_L g70 ( 
.A(n_44),
.Y(n_70)
);

INVx8_ASAP7_75t_L g155 ( 
.A(n_70),
.Y(n_155)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_22),
.Y(n_71)
);

INVx6_ASAP7_75t_L g140 ( 
.A(n_71),
.Y(n_140)
);

CKINVDCx16_ASAP7_75t_R g72 ( 
.A(n_44),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_72),
.B(n_83),
.Y(n_118)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_48),
.Y(n_73)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_73),
.Y(n_111)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_37),
.Y(n_74)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_74),
.Y(n_105)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_32),
.Y(n_75)
);

INVx4_ASAP7_75t_L g128 ( 
.A(n_75),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_22),
.Y(n_76)
);

INVx6_ASAP7_75t_L g142 ( 
.A(n_76),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_25),
.B(n_0),
.Y(n_77)
);

BUFx10_ASAP7_75t_L g78 ( 
.A(n_44),
.Y(n_78)
);

INVx4_ASAP7_75t_L g143 ( 
.A(n_78),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_22),
.Y(n_79)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_79),
.Y(n_121)
);

INVx8_ASAP7_75t_L g80 ( 
.A(n_27),
.Y(n_80)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_80),
.Y(n_133)
);

INVx5_ASAP7_75t_L g81 ( 
.A(n_28),
.Y(n_81)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_81),
.Y(n_141)
);

BUFx12f_ASAP7_75t_L g82 ( 
.A(n_32),
.Y(n_82)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_82),
.Y(n_146)
);

OR2x2_ASAP7_75t_L g83 ( 
.A(n_31),
.B(n_20),
.Y(n_83)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_37),
.Y(n_84)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_84),
.Y(n_126)
);

INVx2_ASAP7_75t_SL g85 ( 
.A(n_21),
.Y(n_85)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_85),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_27),
.Y(n_86)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_86),
.Y(n_130)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_20),
.Y(n_87)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_87),
.Y(n_123)
);

BUFx12f_ASAP7_75t_L g88 ( 
.A(n_32),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_88),
.B(n_44),
.Y(n_119)
);

BUFx3_ASAP7_75t_L g89 ( 
.A(n_49),
.Y(n_89)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_89),
.Y(n_136)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_48),
.B(n_0),
.Y(n_90)
);

INVx2_ASAP7_75t_SL g91 ( 
.A(n_21),
.Y(n_91)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_91),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_27),
.Y(n_92)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_92),
.Y(n_145)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_48),
.Y(n_93)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_93),
.Y(n_149)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_21),
.Y(n_94)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_94),
.Y(n_152)
);

INVx8_ASAP7_75t_L g95 ( 
.A(n_27),
.Y(n_95)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_95),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_29),
.Y(n_96)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_96),
.Y(n_159)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_23),
.Y(n_97)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_97),
.Y(n_161)
);

BUFx3_ASAP7_75t_L g98 ( 
.A(n_49),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g150 ( 
.A(n_98),
.B(n_99),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_29),
.Y(n_99)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_23),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_100),
.B(n_49),
.Y(n_160)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_47),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_101),
.B(n_51),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_28),
.B(n_0),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_102),
.B(n_46),
.Y(n_148)
);

INVx8_ASAP7_75t_L g103 ( 
.A(n_29),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_103),
.A2(n_70),
.B1(n_57),
.B2(n_78),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g208 ( 
.A(n_109),
.Y(n_208)
);

AOI21xp33_ASAP7_75t_L g207 ( 
.A1(n_113),
.A2(n_148),
.B(n_154),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_83),
.B(n_30),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g185 ( 
.A(n_116),
.B(n_129),
.Y(n_185)
);

INVxp67_ASAP7_75t_L g216 ( 
.A(n_119),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_68),
.A2(n_52),
.B1(n_29),
.B2(n_50),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_127),
.A2(n_158),
.B1(n_39),
.B2(n_33),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_68),
.B(n_25),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_90),
.A2(n_52),
.B1(n_40),
.B2(n_50),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_131),
.A2(n_43),
.B1(n_35),
.B2(n_41),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_54),
.B(n_30),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_132),
.B(n_135),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_78),
.Y(n_135)
);

AND2x4_ASAP7_75t_SL g137 ( 
.A(n_53),
.B(n_23),
.Y(n_137)
);

AND2x4_ASAP7_75t_SL g217 ( 
.A(n_137),
.B(n_42),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_54),
.B(n_34),
.Y(n_138)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_138),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_82),
.B(n_34),
.Y(n_144)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_144),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_85),
.B(n_33),
.C(n_50),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_153),
.B(n_150),
.C(n_40),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_SL g154 ( 
.A(n_82),
.B(n_46),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_55),
.A2(n_52),
.B1(n_33),
.B2(n_50),
.Y(n_158)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_160),
.Y(n_204)
);

INVx1_ASAP7_75t_SL g162 ( 
.A(n_117),
.Y(n_162)
);

AND2x2_ASAP7_75t_L g221 ( 
.A(n_162),
.B(n_212),
.Y(n_221)
);

INVx4_ASAP7_75t_L g163 ( 
.A(n_114),
.Y(n_163)
);

INVx3_ASAP7_75t_L g223 ( 
.A(n_163),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_106),
.A2(n_79),
.B1(n_99),
.B2(n_59),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_164),
.A2(n_167),
.B1(n_168),
.B2(n_179),
.Y(n_233)
);

AOI32xp33_ASAP7_75t_L g165 ( 
.A1(n_147),
.A2(n_91),
.A3(n_88),
.B1(n_94),
.B2(n_97),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_165),
.B(n_110),
.Y(n_224)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_117),
.Y(n_166)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_166),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_131),
.A2(n_60),
.B1(n_65),
.B2(n_96),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_112),
.A2(n_56),
.B1(n_98),
.B2(n_75),
.Y(n_170)
);

CKINVDCx16_ASAP7_75t_R g220 ( 
.A(n_170),
.Y(n_220)
);

BUFx2_ASAP7_75t_L g172 ( 
.A(n_110),
.Y(n_172)
);

BUFx3_ASAP7_75t_L g226 ( 
.A(n_172),
.Y(n_226)
);

INVx4_ASAP7_75t_L g173 ( 
.A(n_114),
.Y(n_173)
);

INVx3_ASAP7_75t_L g259 ( 
.A(n_173),
.Y(n_259)
);

INVx5_ASAP7_75t_L g174 ( 
.A(n_143),
.Y(n_174)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_174),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_112),
.B(n_51),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_175),
.B(n_189),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_L g218 ( 
.A1(n_176),
.A2(n_182),
.B1(n_188),
.B2(n_195),
.Y(n_218)
);

O2A1O1Ixp33_ASAP7_75t_SL g177 ( 
.A1(n_137),
.A2(n_103),
.B(n_95),
.C(n_71),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_177),
.B(n_203),
.Y(n_241)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_123),
.Y(n_178)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_178),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_153),
.A2(n_92),
.B1(n_86),
.B2(n_76),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g180 ( 
.A(n_134),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g266 ( 
.A(n_180),
.Y(n_266)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_124),
.Y(n_181)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_181),
.Y(n_228)
);

AOI22xp33_ASAP7_75t_L g182 ( 
.A1(n_127),
.A2(n_80),
.B1(n_36),
.B2(n_47),
.Y(n_182)
);

HB1xp67_ASAP7_75t_L g183 ( 
.A(n_161),
.Y(n_183)
);

CKINVDCx16_ASAP7_75t_R g229 ( 
.A(n_183),
.Y(n_229)
);

BUFx3_ASAP7_75t_L g184 ( 
.A(n_122),
.Y(n_184)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_184),
.Y(n_245)
);

AOI22xp33_ASAP7_75t_SL g186 ( 
.A1(n_108),
.A2(n_39),
.B1(n_26),
.B2(n_35),
.Y(n_186)
);

CKINVDCx16_ASAP7_75t_R g258 ( 
.A(n_186),
.Y(n_258)
);

INVx3_ASAP7_75t_L g187 ( 
.A(n_155),
.Y(n_187)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_187),
.Y(n_253)
);

AOI22xp33_ASAP7_75t_SL g188 ( 
.A1(n_157),
.A2(n_39),
.B1(n_26),
.B2(n_35),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_118),
.B(n_36),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_107),
.Y(n_190)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_190),
.Y(n_231)
);

BUFx12f_ASAP7_75t_L g191 ( 
.A(n_122),
.Y(n_191)
);

INVx6_ASAP7_75t_L g239 ( 
.A(n_191),
.Y(n_239)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_130),
.Y(n_192)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_192),
.Y(n_260)
);

BUFx3_ASAP7_75t_L g193 ( 
.A(n_146),
.Y(n_193)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_193),
.Y(n_235)
);

AOI22xp33_ASAP7_75t_SL g195 ( 
.A1(n_141),
.A2(n_39),
.B1(n_26),
.B2(n_41),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_104),
.B(n_43),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_196),
.B(n_200),
.Y(n_248)
);

INVx4_ASAP7_75t_L g197 ( 
.A(n_155),
.Y(n_197)
);

INVx6_ASAP7_75t_L g251 ( 
.A(n_197),
.Y(n_251)
);

AOI22xp33_ASAP7_75t_SL g198 ( 
.A1(n_141),
.A2(n_43),
.B1(n_41),
.B2(n_89),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g243 ( 
.A1(n_198),
.A2(n_202),
.B1(n_120),
.B2(n_151),
.Y(n_243)
);

INVx5_ASAP7_75t_L g199 ( 
.A(n_143),
.Y(n_199)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_199),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_105),
.B(n_73),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_109),
.A2(n_42),
.B1(n_40),
.B2(n_33),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_201),
.A2(n_139),
.B1(n_140),
.B2(n_133),
.Y(n_244)
);

AOI22xp33_ASAP7_75t_SL g202 ( 
.A1(n_128),
.A2(n_61),
.B1(n_42),
.B2(n_40),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_150),
.Y(n_203)
);

INVx8_ASAP7_75t_L g205 ( 
.A(n_140),
.Y(n_205)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_205),
.Y(n_247)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_145),
.Y(n_206)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_206),
.Y(n_249)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_136),
.Y(n_209)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_209),
.Y(n_255)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_126),
.Y(n_210)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_210),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_137),
.B(n_66),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_211),
.B(n_1),
.Y(n_263)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_159),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_213),
.B(n_215),
.C(n_146),
.Y(n_234)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_107),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_214),
.B(n_111),
.Y(n_254)
);

AND2x2_ASAP7_75t_SL g215 ( 
.A(n_149),
.B(n_88),
.Y(n_215)
);

OAI21x1_ASAP7_75t_SL g265 ( 
.A1(n_217),
.A2(n_38),
.B(n_3),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_176),
.A2(n_121),
.B1(n_115),
.B2(n_142),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_219),
.A2(n_237),
.B1(n_242),
.B2(n_256),
.Y(n_267)
);

AND2x2_ASAP7_75t_L g309 ( 
.A(n_224),
.B(n_263),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_185),
.B(n_189),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_SL g300 ( 
.A(n_225),
.B(n_238),
.Y(n_300)
);

XOR2xp5_ASAP7_75t_L g304 ( 
.A(n_234),
.B(n_174),
.Y(n_304)
);

NOR3xp33_ASAP7_75t_L g236 ( 
.A(n_175),
.B(n_42),
.C(n_134),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g268 ( 
.A(n_236),
.B(n_252),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_213),
.A2(n_121),
.B1(n_125),
.B2(n_115),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_SL g238 ( 
.A(n_207),
.B(n_128),
.Y(n_238)
);

MAJx2_ASAP7_75t_L g240 ( 
.A(n_204),
.B(n_152),
.C(n_156),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_240),
.B(n_181),
.C(n_210),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_208),
.A2(n_142),
.B1(n_125),
.B2(n_139),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_243),
.A2(n_264),
.B1(n_172),
.B2(n_184),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_244),
.A2(n_170),
.B1(n_173),
.B2(n_163),
.Y(n_275)
);

AOI22x1_ASAP7_75t_SL g250 ( 
.A1(n_177),
.A2(n_120),
.B1(n_151),
.B2(n_133),
.Y(n_250)
);

INVxp67_ASAP7_75t_L g311 ( 
.A(n_250),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_194),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_254),
.B(n_257),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_L g256 ( 
.A1(n_208),
.A2(n_111),
.B1(n_38),
.B2(n_2),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_169),
.B(n_0),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_211),
.A2(n_38),
.B1(n_2),
.B2(n_3),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_261),
.A2(n_162),
.B1(n_166),
.B2(n_168),
.Y(n_272)
);

OAI22xp33_ASAP7_75t_SL g264 ( 
.A1(n_216),
.A2(n_38),
.B1(n_3),
.B2(n_4),
.Y(n_264)
);

A2O1A1O1Ixp25_ASAP7_75t_L g287 ( 
.A1(n_265),
.A2(n_190),
.B(n_3),
.C(n_4),
.D(n_5),
.Y(n_287)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_227),
.Y(n_269)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_269),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_221),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_270),
.B(n_289),
.Y(n_317)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_231),
.Y(n_271)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_271),
.Y(n_337)
);

OAI22xp33_ASAP7_75t_SL g344 ( 
.A1(n_272),
.A2(n_284),
.B1(n_226),
.B2(n_245),
.Y(n_344)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_224),
.A2(n_218),
.B1(n_219),
.B2(n_237),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_L g318 ( 
.A1(n_273),
.A2(n_274),
.B1(n_277),
.B2(n_250),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_220),
.A2(n_217),
.B1(n_196),
.B2(n_216),
.Y(n_274)
);

AOI22xp33_ASAP7_75t_L g313 ( 
.A1(n_275),
.A2(n_285),
.B1(n_290),
.B2(n_305),
.Y(n_313)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_227),
.Y(n_276)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_276),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_248),
.A2(n_217),
.B1(n_215),
.B2(n_200),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_248),
.B(n_178),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_278),
.B(n_292),
.Y(n_316)
);

OAI21xp5_ASAP7_75t_L g279 ( 
.A1(n_241),
.A2(n_215),
.B(n_171),
.Y(n_279)
);

INVxp67_ASAP7_75t_L g312 ( 
.A(n_279),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_221),
.Y(n_280)
);

INVxp67_ASAP7_75t_SL g336 ( 
.A(n_280),
.Y(n_336)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_222),
.Y(n_281)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_281),
.Y(n_330)
);

XNOR2xp5_ASAP7_75t_SL g346 ( 
.A(n_283),
.B(n_307),
.Y(n_346)
);

OAI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_233),
.A2(n_205),
.B1(n_192),
.B2(n_206),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_221),
.Y(n_286)
);

INVxp67_ASAP7_75t_SL g351 ( 
.A(n_286),
.Y(n_351)
);

OAI21xp5_ASAP7_75t_SL g325 ( 
.A1(n_287),
.A2(n_245),
.B(n_235),
.Y(n_325)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_222),
.Y(n_288)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_288),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_231),
.Y(n_289)
);

AOI22xp33_ASAP7_75t_L g290 ( 
.A1(n_242),
.A2(n_212),
.B1(n_187),
.B2(n_209),
.Y(n_290)
);

CKINVDCx16_ASAP7_75t_R g291 ( 
.A(n_229),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_291),
.B(n_297),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_263),
.B(n_234),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_261),
.B(n_197),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_293),
.B(n_294),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_232),
.B(n_193),
.Y(n_294)
);

INVx4_ASAP7_75t_L g295 ( 
.A(n_251),
.Y(n_295)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_295),
.Y(n_340)
);

INVx4_ASAP7_75t_L g296 ( 
.A(n_251),
.Y(n_296)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_296),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_262),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_228),
.Y(n_298)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_298),
.Y(n_345)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_228),
.Y(n_299)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_299),
.Y(n_352)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_262),
.Y(n_301)
);

INVx1_ASAP7_75t_SL g314 ( 
.A(n_301),
.Y(n_314)
);

HB1xp67_ASAP7_75t_L g302 ( 
.A(n_253),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_302),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_232),
.B(n_199),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g341 ( 
.A(n_303),
.B(n_259),
.Y(n_341)
);

MAJIxp5_ASAP7_75t_L g349 ( 
.A(n_304),
.B(n_266),
.C(n_239),
.Y(n_349)
);

OAI22xp5_ASAP7_75t_SL g305 ( 
.A1(n_233),
.A2(n_180),
.B1(n_191),
.B2(n_38),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_249),
.Y(n_306)
);

INVxp67_ASAP7_75t_L g347 ( 
.A(n_306),
.Y(n_347)
);

XNOR2xp5_ASAP7_75t_SL g307 ( 
.A(n_240),
.B(n_191),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_255),
.B(n_1),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_SL g323 ( 
.A(n_308),
.B(n_223),
.Y(n_323)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_249),
.Y(n_310)
);

BUFx3_ASAP7_75t_L g320 ( 
.A(n_310),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_L g356 ( 
.A1(n_318),
.A2(n_344),
.B1(n_348),
.B2(n_350),
.Y(n_356)
);

OAI32xp33_ASAP7_75t_L g321 ( 
.A1(n_278),
.A2(n_265),
.A3(n_258),
.B1(n_247),
.B2(n_253),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_321),
.B(n_324),
.Y(n_358)
);

XOR2xp5_ASAP7_75t_L g322 ( 
.A(n_304),
.B(n_255),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g380 ( 
.A(n_322),
.B(n_349),
.C(n_287),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_SL g377 ( 
.A(n_323),
.B(n_333),
.Y(n_377)
);

OAI32xp33_ASAP7_75t_L g324 ( 
.A1(n_293),
.A2(n_247),
.A3(n_246),
.B1(n_260),
.B2(n_230),
.Y(n_324)
);

INVxp67_ASAP7_75t_L g365 ( 
.A(n_325),
.Y(n_365)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_289),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_326),
.B(n_327),
.Y(n_357)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_282),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g332 ( 
.A(n_294),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_332),
.B(n_334),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_SL g333 ( 
.A(n_300),
.B(n_223),
.Y(n_333)
);

CKINVDCx16_ASAP7_75t_R g334 ( 
.A(n_279),
.Y(n_334)
);

CKINVDCx14_ASAP7_75t_R g335 ( 
.A(n_268),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g376 ( 
.A(n_335),
.B(n_334),
.Y(n_376)
);

OAI32xp33_ASAP7_75t_L g339 ( 
.A1(n_303),
.A2(n_246),
.A3(n_260),
.B1(n_230),
.B2(n_235),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_339),
.B(n_275),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_SL g363 ( 
.A(n_341),
.B(n_283),
.Y(n_363)
);

AOI21xp5_ASAP7_75t_L g342 ( 
.A1(n_311),
.A2(n_259),
.B(n_244),
.Y(n_342)
);

AOI21xp5_ASAP7_75t_L g354 ( 
.A1(n_342),
.A2(n_284),
.B(n_267),
.Y(n_354)
);

OAI22xp5_ASAP7_75t_SL g348 ( 
.A1(n_273),
.A2(n_266),
.B1(n_226),
.B2(n_239),
.Y(n_348)
);

OAI22xp5_ASAP7_75t_SL g350 ( 
.A1(n_311),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_350)
);

CKINVDCx14_ASAP7_75t_R g353 ( 
.A(n_317),
.Y(n_353)
);

CKINVDCx16_ASAP7_75t_R g405 ( 
.A(n_353),
.Y(n_405)
);

AOI21xp5_ASAP7_75t_L g389 ( 
.A1(n_354),
.A2(n_359),
.B(n_364),
.Y(n_389)
);

XOR2xp5_ASAP7_75t_SL g355 ( 
.A(n_316),
.B(n_309),
.Y(n_355)
);

XNOR2xp5_ASAP7_75t_L g388 ( 
.A(n_355),
.B(n_346),
.Y(n_388)
);

AOI21xp5_ASAP7_75t_L g359 ( 
.A1(n_342),
.A2(n_309),
.B(n_274),
.Y(n_359)
);

OAI22xp5_ASAP7_75t_L g360 ( 
.A1(n_332),
.A2(n_267),
.B1(n_277),
.B2(n_272),
.Y(n_360)
);

AOI22xp5_ASAP7_75t_L g395 ( 
.A1(n_360),
.A2(n_370),
.B1(n_387),
.B2(n_352),
.Y(n_395)
);

INVx2_ASAP7_75t_L g361 ( 
.A(n_337),
.Y(n_361)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_361),
.Y(n_394)
);

AOI22xp5_ASAP7_75t_L g362 ( 
.A1(n_318),
.A2(n_285),
.B1(n_309),
.B2(n_305),
.Y(n_362)
);

OAI22xp5_ASAP7_75t_L g413 ( 
.A1(n_362),
.A2(n_367),
.B1(n_374),
.B2(n_379),
.Y(n_413)
);

XNOR2xp5_ASAP7_75t_SL g418 ( 
.A(n_363),
.B(n_343),
.Y(n_418)
);

AO21x1_ASAP7_75t_L g364 ( 
.A1(n_336),
.A2(n_307),
.B(n_292),
.Y(n_364)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_366),
.Y(n_402)
);

AOI22xp5_ASAP7_75t_L g367 ( 
.A1(n_348),
.A2(n_286),
.B1(n_280),
.B2(n_281),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_319),
.Y(n_368)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_368),
.Y(n_397)
);

CKINVDCx16_ASAP7_75t_R g369 ( 
.A(n_329),
.Y(n_369)
);

AOI22xp33_ASAP7_75t_L g396 ( 
.A1(n_369),
.A2(n_375),
.B1(n_384),
.B2(n_314),
.Y(n_396)
);

OAI22xp5_ASAP7_75t_SL g370 ( 
.A1(n_331),
.A2(n_288),
.B1(n_276),
.B2(n_269),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_319),
.Y(n_371)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_371),
.Y(n_399)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_328),
.Y(n_373)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_373),
.Y(n_417)
);

AOI22xp5_ASAP7_75t_L g374 ( 
.A1(n_331),
.A2(n_298),
.B1(n_299),
.B2(n_271),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_328),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_SL g390 ( 
.A(n_376),
.B(n_385),
.Y(n_390)
);

XOR2xp5_ASAP7_75t_L g378 ( 
.A(n_346),
.B(n_322),
.Y(n_378)
);

MAJIxp5_ASAP7_75t_L g391 ( 
.A(n_378),
.B(n_380),
.C(n_312),
.Y(n_391)
);

AOI22xp5_ASAP7_75t_L g379 ( 
.A1(n_312),
.A2(n_310),
.B1(n_306),
.B2(n_301),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_326),
.B(n_296),
.Y(n_381)
);

CKINVDCx20_ASAP7_75t_R g392 ( 
.A(n_381),
.Y(n_392)
);

OAI21xp5_ASAP7_75t_L g382 ( 
.A1(n_351),
.A2(n_295),
.B(n_7),
.Y(n_382)
);

OAI21xp5_ASAP7_75t_L g393 ( 
.A1(n_382),
.A2(n_350),
.B(n_323),
.Y(n_393)
);

CKINVDCx20_ASAP7_75t_R g383 ( 
.A(n_315),
.Y(n_383)
);

CKINVDCx20_ASAP7_75t_R g398 ( 
.A(n_383),
.Y(n_398)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_330),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_L g385 ( 
.A(n_327),
.B(n_5),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_316),
.B(n_7),
.Y(n_386)
);

CKINVDCx16_ASAP7_75t_R g411 ( 
.A(n_386),
.Y(n_411)
);

OAI22xp5_ASAP7_75t_L g387 ( 
.A1(n_313),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_387)
);

MAJx2_ASAP7_75t_L g446 ( 
.A(n_388),
.B(n_391),
.C(n_377),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_393),
.B(n_382),
.Y(n_421)
);

OAI22xp5_ASAP7_75t_L g434 ( 
.A1(n_395),
.A2(n_414),
.B1(n_419),
.B2(n_356),
.Y(n_434)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_396),
.Y(n_426)
);

MAJIxp5_ASAP7_75t_L g400 ( 
.A(n_378),
.B(n_349),
.C(n_341),
.Y(n_400)
);

MAJIxp5_ASAP7_75t_L g435 ( 
.A(n_400),
.B(n_406),
.C(n_407),
.Y(n_435)
);

AOI22xp5_ASAP7_75t_L g401 ( 
.A1(n_360),
.A2(n_333),
.B1(n_347),
.B2(n_314),
.Y(n_401)
);

OAI22xp5_ASAP7_75t_SL g441 ( 
.A1(n_401),
.A2(n_409),
.B1(n_362),
.B2(n_379),
.Y(n_441)
);

XOR2xp5_ASAP7_75t_L g403 ( 
.A(n_364),
.B(n_363),
.Y(n_403)
);

XOR2xp5_ASAP7_75t_L g433 ( 
.A(n_403),
.B(n_404),
.Y(n_433)
);

XNOR2xp5_ASAP7_75t_L g404 ( 
.A(n_364),
.B(n_325),
.Y(n_404)
);

MAJIxp5_ASAP7_75t_L g406 ( 
.A(n_380),
.B(n_347),
.C(n_352),
.Y(n_406)
);

MAJIxp5_ASAP7_75t_L g407 ( 
.A(n_355),
.B(n_345),
.C(n_338),
.Y(n_407)
);

XNOR2xp5_ASAP7_75t_L g408 ( 
.A(n_372),
.B(n_345),
.Y(n_408)
);

MAJIxp5_ASAP7_75t_L g436 ( 
.A(n_408),
.B(n_410),
.C(n_412),
.Y(n_436)
);

AOI22xp5_ASAP7_75t_L g409 ( 
.A1(n_366),
.A2(n_338),
.B1(n_330),
.B2(n_321),
.Y(n_409)
);

XOR2xp5_ASAP7_75t_L g410 ( 
.A(n_372),
.B(n_339),
.Y(n_410)
);

XOR2xp5_ASAP7_75t_L g412 ( 
.A(n_376),
.B(n_324),
.Y(n_412)
);

AOI22xp33_ASAP7_75t_L g414 ( 
.A1(n_357),
.A2(n_369),
.B1(n_370),
.B2(n_383),
.Y(n_414)
);

OAI21xp5_ASAP7_75t_L g415 ( 
.A1(n_359),
.A2(n_315),
.B(n_320),
.Y(n_415)
);

OAI21xp5_ASAP7_75t_L g428 ( 
.A1(n_415),
.A2(n_354),
.B(n_358),
.Y(n_428)
);

OAI22x1_ASAP7_75t_SL g416 ( 
.A1(n_356),
.A2(n_320),
.B1(n_340),
.B2(n_343),
.Y(n_416)
);

AOI22xp5_ASAP7_75t_L g439 ( 
.A1(n_416),
.A2(n_358),
.B1(n_384),
.B2(n_371),
.Y(n_439)
);

XNOR2xp5_ASAP7_75t_L g440 ( 
.A(n_418),
.B(n_388),
.Y(n_440)
);

OAI22xp5_ASAP7_75t_L g419 ( 
.A1(n_353),
.A2(n_337),
.B1(n_340),
.B2(n_11),
.Y(n_419)
);

NOR2xp33_ASAP7_75t_L g420 ( 
.A(n_390),
.B(n_357),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_420),
.B(n_421),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_398),
.B(n_381),
.Y(n_422)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_422),
.Y(n_447)
);

CKINVDCx20_ASAP7_75t_R g423 ( 
.A(n_392),
.Y(n_423)
);

BUFx12f_ASAP7_75t_L g463 ( 
.A(n_423),
.Y(n_463)
);

CKINVDCx20_ASAP7_75t_R g424 ( 
.A(n_401),
.Y(n_424)
);

OAI21xp5_ASAP7_75t_SL g468 ( 
.A1(n_424),
.A2(n_439),
.B(n_8),
.Y(n_468)
);

NOR2xp33_ASAP7_75t_SL g425 ( 
.A(n_405),
.B(n_385),
.Y(n_425)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_425),
.Y(n_448)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_417),
.Y(n_427)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_427),
.Y(n_449)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_428),
.Y(n_456)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_417),
.Y(n_429)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_429),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_408),
.B(n_374),
.Y(n_430)
);

XNOR2xp5_ASAP7_75t_L g455 ( 
.A(n_430),
.B(n_432),
.Y(n_455)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_397),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_SL g465 ( 
.A(n_431),
.B(n_445),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_395),
.B(n_386),
.Y(n_432)
);

AOI22xp5_ASAP7_75t_L g450 ( 
.A1(n_434),
.A2(n_441),
.B1(n_402),
.B2(n_415),
.Y(n_450)
);

MAJIxp5_ASAP7_75t_L g437 ( 
.A(n_400),
.B(n_406),
.C(n_391),
.Y(n_437)
);

MAJIxp5_ASAP7_75t_L g451 ( 
.A(n_437),
.B(n_438),
.C(n_444),
.Y(n_451)
);

MAJIxp5_ASAP7_75t_L g438 ( 
.A(n_403),
.B(n_365),
.C(n_367),
.Y(n_438)
);

XNOR2xp5_ASAP7_75t_L g462 ( 
.A(n_440),
.B(n_442),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_413),
.B(n_375),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_411),
.B(n_373),
.Y(n_443)
);

XOR2xp5_ASAP7_75t_L g452 ( 
.A(n_443),
.B(n_409),
.Y(n_452)
);

MAJIxp5_ASAP7_75t_L g444 ( 
.A(n_418),
.B(n_368),
.C(n_361),
.Y(n_444)
);

AOI22xp5_ASAP7_75t_L g445 ( 
.A1(n_402),
.A2(n_416),
.B1(n_410),
.B2(n_412),
.Y(n_445)
);

MAJIxp5_ASAP7_75t_L g453 ( 
.A(n_446),
.B(n_407),
.C(n_404),
.Y(n_453)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_450),
.Y(n_470)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_452),
.Y(n_477)
);

MAJx2_ASAP7_75t_L g472 ( 
.A(n_453),
.B(n_446),
.C(n_440),
.Y(n_472)
);

AOI22xp5_ASAP7_75t_L g457 ( 
.A1(n_441),
.A2(n_424),
.B1(n_426),
.B2(n_442),
.Y(n_457)
);

HB1xp67_ASAP7_75t_L g469 ( 
.A(n_457),
.Y(n_469)
);

XOR2xp5_ASAP7_75t_L g458 ( 
.A(n_436),
.B(n_389),
.Y(n_458)
);

XNOR2xp5_ASAP7_75t_SL g481 ( 
.A(n_458),
.B(n_461),
.Y(n_481)
);

MAJIxp5_ASAP7_75t_L g459 ( 
.A(n_435),
.B(n_389),
.C(n_394),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_459),
.B(n_467),
.Y(n_475)
);

XOR2xp5_ASAP7_75t_L g461 ( 
.A(n_436),
.B(n_393),
.Y(n_461)
);

FAx1_ASAP7_75t_SL g464 ( 
.A(n_438),
.B(n_377),
.CI(n_387),
.CON(n_464),
.SN(n_464)
);

NOR2xp33_ASAP7_75t_L g483 ( 
.A(n_464),
.B(n_421),
.Y(n_483)
);

OAI21xp5_ASAP7_75t_SL g466 ( 
.A1(n_435),
.A2(n_423),
.B(n_422),
.Y(n_466)
);

AOI21xp5_ASAP7_75t_L g478 ( 
.A1(n_466),
.A2(n_445),
.B(n_443),
.Y(n_478)
);

MAJIxp5_ASAP7_75t_L g467 ( 
.A(n_437),
.B(n_394),
.C(n_399),
.Y(n_467)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_468),
.Y(n_480)
);

XNOR2x1_ASAP7_75t_L g471 ( 
.A(n_458),
.B(n_433),
.Y(n_471)
);

XOR2xp5_ASAP7_75t_L g486 ( 
.A(n_471),
.B(n_485),
.Y(n_486)
);

MAJIxp5_ASAP7_75t_L g495 ( 
.A(n_472),
.B(n_473),
.C(n_451),
.Y(n_495)
);

MAJIxp5_ASAP7_75t_L g473 ( 
.A(n_467),
.B(n_444),
.C(n_433),
.Y(n_473)
);

AOI22xp5_ASAP7_75t_L g474 ( 
.A1(n_452),
.A2(n_426),
.B1(n_428),
.B2(n_432),
.Y(n_474)
);

OAI22xp33_ASAP7_75t_SL g490 ( 
.A1(n_474),
.A2(n_476),
.B1(n_447),
.B2(n_469),
.Y(n_490)
);

AOI22xp5_ASAP7_75t_L g476 ( 
.A1(n_448),
.A2(n_429),
.B1(n_427),
.B2(n_425),
.Y(n_476)
);

OAI21xp5_ASAP7_75t_SL g489 ( 
.A1(n_478),
.A2(n_483),
.B(n_453),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_454),
.B(n_431),
.Y(n_479)
);

NOR2xp33_ASAP7_75t_L g492 ( 
.A(n_479),
.B(n_482),
.Y(n_492)
);

BUFx24_ASAP7_75t_SL g482 ( 
.A(n_464),
.Y(n_482)
);

NOR2xp33_ASAP7_75t_L g484 ( 
.A(n_464),
.B(n_439),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_484),
.B(n_459),
.Y(n_487)
);

XNOR2xp5_ASAP7_75t_L g485 ( 
.A(n_451),
.B(n_430),
.Y(n_485)
);

INVxp67_ASAP7_75t_L g510 ( 
.A(n_487),
.Y(n_510)
);

AOI21xp5_ASAP7_75t_L g488 ( 
.A1(n_470),
.A2(n_456),
.B(n_465),
.Y(n_488)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_488),
.Y(n_502)
);

MAJx2_ASAP7_75t_L g511 ( 
.A(n_489),
.B(n_495),
.C(n_12),
.Y(n_511)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_490),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_480),
.B(n_463),
.Y(n_491)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_491),
.Y(n_514)
);

AOI21xp5_ASAP7_75t_L g493 ( 
.A1(n_474),
.A2(n_457),
.B(n_450),
.Y(n_493)
);

XNOR2xp5_ASAP7_75t_L g509 ( 
.A(n_493),
.B(n_497),
.Y(n_509)
);

AOI22xp5_ASAP7_75t_L g494 ( 
.A1(n_477),
.A2(n_461),
.B1(n_449),
.B2(n_460),
.Y(n_494)
);

OAI22xp5_ASAP7_75t_SL g513 ( 
.A1(n_494),
.A2(n_15),
.B1(n_16),
.B2(n_501),
.Y(n_513)
);

INVx11_ASAP7_75t_L g496 ( 
.A(n_475),
.Y(n_496)
);

AOI22xp5_ASAP7_75t_L g503 ( 
.A1(n_496),
.A2(n_501),
.B1(n_472),
.B2(n_462),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_485),
.B(n_463),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_473),
.B(n_463),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_SL g504 ( 
.A(n_498),
.B(n_499),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_481),
.B(n_455),
.Y(n_499)
);

MAJIxp5_ASAP7_75t_L g500 ( 
.A(n_481),
.B(n_462),
.C(n_455),
.Y(n_500)
);

NOR2xp33_ASAP7_75t_L g506 ( 
.A(n_500),
.B(n_8),
.Y(n_506)
);

INVx1_ASAP7_75t_SL g501 ( 
.A(n_471),
.Y(n_501)
);

OAI21x1_ASAP7_75t_SL g519 ( 
.A1(n_503),
.A2(n_508),
.B(n_488),
.Y(n_519)
);

AOI22xp5_ASAP7_75t_L g505 ( 
.A1(n_496),
.A2(n_468),
.B1(n_10),
.B2(n_11),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_505),
.B(n_506),
.Y(n_522)
);

AOI22xp5_ASAP7_75t_L g508 ( 
.A1(n_491),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_508)
);

XNOR2xp5_ASAP7_75t_L g521 ( 
.A(n_511),
.B(n_499),
.Y(n_521)
);

NOR2xp33_ASAP7_75t_SL g512 ( 
.A(n_492),
.B(n_13),
.Y(n_512)
);

NOR2xp33_ASAP7_75t_L g518 ( 
.A(n_512),
.B(n_15),
.Y(n_518)
);

INVx1_ASAP7_75t_SL g517 ( 
.A(n_513),
.Y(n_517)
);

AOI21x1_ASAP7_75t_SL g515 ( 
.A1(n_504),
.A2(n_489),
.B(n_498),
.Y(n_515)
);

OAI21xp5_ASAP7_75t_L g527 ( 
.A1(n_515),
.A2(n_520),
.B(n_507),
.Y(n_527)
);

MAJIxp5_ASAP7_75t_L g516 ( 
.A(n_510),
.B(n_495),
.C(n_487),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_SL g526 ( 
.A(n_516),
.B(n_521),
.Y(n_526)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_518),
.Y(n_524)
);

A2O1A1Ixp33_ASAP7_75t_SL g525 ( 
.A1(n_519),
.A2(n_493),
.B(n_514),
.C(n_502),
.Y(n_525)
);

OAI21xp5_ASAP7_75t_SL g520 ( 
.A1(n_510),
.A2(n_497),
.B(n_494),
.Y(n_520)
);

INVxp67_ASAP7_75t_L g523 ( 
.A(n_522),
.Y(n_523)
);

AOI221xp5_ASAP7_75t_SL g529 ( 
.A1(n_523),
.A2(n_525),
.B1(n_511),
.B2(n_509),
.C(n_486),
.Y(n_529)
);

AOI21xp5_ASAP7_75t_L g528 ( 
.A1(n_527),
.A2(n_509),
.B(n_486),
.Y(n_528)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_528),
.Y(n_531)
);

AO21x2_ASAP7_75t_L g532 ( 
.A1(n_529),
.A2(n_530),
.B(n_524),
.Y(n_532)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_526),
.Y(n_530)
);

O2A1O1Ixp33_ASAP7_75t_L g533 ( 
.A1(n_532),
.A2(n_517),
.B(n_518),
.C(n_500),
.Y(n_533)
);

AOI21xp5_ASAP7_75t_SL g534 ( 
.A1(n_533),
.A2(n_531),
.B(n_517),
.Y(n_534)
);

NOR2xp33_ASAP7_75t_L g535 ( 
.A(n_534),
.B(n_508),
.Y(n_535)
);

NOR2xp33_ASAP7_75t_L g536 ( 
.A(n_535),
.B(n_16),
.Y(n_536)
);


endmodule