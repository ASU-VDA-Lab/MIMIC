module fake_ariane_2738_n_1842 (n_83, n_8, n_56, n_60, n_160, n_64, n_119, n_124, n_167, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_149, n_34, n_158, n_69, n_95, n_92, n_143, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_152, n_120, n_106, n_12, n_53, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_166, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_159, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_148, n_164, n_52, n_157, n_135, n_73, n_77, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_151, n_136, n_28, n_80, n_146, n_97, n_154, n_142, n_161, n_14, n_163, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_1842);

input n_83;
input n_8;
input n_56;
input n_60;
input n_160;
input n_64;
input n_119;
input n_124;
input n_167;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_149;
input n_34;
input n_158;
input n_69;
input n_95;
input n_92;
input n_143;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_152;
input n_120;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_166;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_159;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_164;
input n_52;
input n_157;
input n_135;
input n_73;
input n_77;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_151;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1842;

wire n_913;
wire n_1681;
wire n_1486;
wire n_1507;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_610;
wire n_245;
wire n_1713;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_187;
wire n_1463;
wire n_1238;
wire n_1515;
wire n_817;
wire n_1837;
wire n_924;
wire n_781;
wire n_1566;
wire n_189;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_524;
wire n_634;
wire n_1214;
wire n_1839;
wire n_1246;
wire n_1138;
wire n_214;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_232;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1835;
wire n_1457;
wire n_377;
wire n_1682;
wire n_1836;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_958;
wire n_945;
wire n_813;
wire n_419;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1184;
wire n_202;
wire n_1535;
wire n_500;
wire n_754;
wire n_665;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1277;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_672;
wire n_740;
wire n_1283;
wire n_1736;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_242;
wire n_645;
wire n_331;
wire n_559;
wire n_267;
wire n_495;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_200;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_587;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_352;
wire n_206;
wire n_899;
wire n_1703;
wire n_611;
wire n_1295;
wire n_238;
wire n_365;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_192;
wire n_661;
wire n_1751;
wire n_300;
wire n_533;
wire n_438;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_1811;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_1840;
wire n_376;
wire n_512;
wire n_1597;
wire n_1771;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_237;
wire n_780;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_209;
wire n_490;
wire n_1461;
wire n_1391;
wire n_225;
wire n_1599;
wire n_1006;
wire n_1830;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_1838;
wire n_1594;
wire n_680;
wire n_287;
wire n_1716;
wire n_302;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_212;
wire n_851;
wire n_444;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_1819;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_182;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_1833;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_460;
wire n_1555;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_179;
wire n_1292;
wire n_1178;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_306;
wire n_203;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1787;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_1717;
wire n_1812;
wire n_824;
wire n_428;
wire n_892;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_990;
wire n_1623;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_1780;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1825;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1832;
wire n_1841;
wire n_1680;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_1731;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_698;
wire n_1674;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_172;
wire n_1058;
wire n_347;
wire n_1042;
wire n_183;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_205;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_1728;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_1817;
wire n_348;
wire n_552;
wire n_670;
wire n_1826;
wire n_379;
wire n_264;
wire n_441;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_1743;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_194;
wire n_1802;
wire n_1163;
wire n_186;
wire n_1795;
wire n_1384;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1648;
wire n_1413;
wire n_855;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_647;
wire n_1423;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_529;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1828;
wire n_1798;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_1105;
wire n_547;
wire n_439;
wire n_677;
wire n_604;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_727;
wire n_699;
wire n_301;
wire n_1726;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_325;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1693;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1823;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_221;
wire n_321;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_888;
wire n_845;
wire n_1649;
wire n_1677;
wire n_1297;
wire n_178;
wire n_551;
wire n_417;
wire n_1708;
wire n_343;
wire n_1222;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_534;
wire n_1791;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_451;
wire n_745;
wire n_1741;
wire n_1572;
wire n_1793;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_769;
wire n_1797;
wire n_1753;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_982;
wire n_1800;
wire n_915;
wire n_215;
wire n_1075;
wire n_454;
wire n_298;
wire n_1331;
wire n_1529;
wire n_1227;
wire n_655;
wire n_1734;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_509;
wire n_666;
wire n_1747;
wire n_430;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_456;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_873;
wire n_1301;
wire n_1748;
wire n_1243;
wire n_1400;
wire n_342;
wire n_1466;
wire n_1513;
wire n_1527;
wire n_358;
wire n_1783;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1668;
wire n_1605;
wire n_1078;
wire n_266;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_1786;
wire n_480;
wire n_1327;
wire n_1475;
wire n_211;
wire n_642;
wire n_1804;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_1757;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_1632;
wire n_1769;
wire n_474;
wire n_805;
wire n_295;
wire n_1658;
wire n_190;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_180;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1258;
wire n_197;
wire n_640;
wire n_463;
wire n_1476;
wire n_1524;
wire n_1733;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_1807;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_1784;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_283;
wire n_806;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_1824;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_1822;
wire n_682;
wire n_1616;
wire n_819;
wire n_586;
wire n_1324;
wire n_1429;
wire n_1778;
wire n_1776;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1759;
wire n_1829;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_1815;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_198;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_169;
wire n_1288;
wire n_1201;
wire n_173;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_1367;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1023;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_467;
wire n_1511;
wire n_1422;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_538;
wire n_1517;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1773;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_810;
wire n_1290;
wire n_181;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_414;
wire n_571;
wire n_1521;
wire n_1694;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_409;
wire n_171;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1444;
wire n_1803;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_1739;
wire n_1814;
wire n_532;
wire n_1789;
wire n_763;
wire n_540;
wire n_216;
wire n_692;
wire n_984;
wire n_1687;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_1816;
wire n_1756;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_1772;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_493;
wire n_1311;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1335;
wire n_1715;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_1785;
wire n_792;
wire n_1262;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1183;
wire n_1326;
wire n_1805;
wire n_981;
wire n_1110;
wire n_1758;
wire n_243;
wire n_1407;
wire n_185;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_184;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_1054;
wire n_508;
wire n_1679;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_191;
wire n_1834;
wire n_978;
wire n_1011;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_170;
wire n_1536;
wire n_1471;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_176;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_541;
wire n_499;
wire n_1775;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_1663;
wire n_1625;
wire n_318;
wire n_1458;
wire n_244;
wire n_679;
wire n_1630;
wire n_220;
wire n_663;
wire n_1720;
wire n_443;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_1735;
wire n_1788;
wire n_391;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_765;
wire n_1809;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_857;
wire n_898;
wire n_363;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_1755;
wire n_1285;
wire n_193;
wire n_733;
wire n_761;
wire n_731;
wire n_336;
wire n_1813;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1106;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_1770;
wire n_701;
wire n_1003;
wire n_1125;
wire n_1710;
wire n_309;
wire n_1344;
wire n_1390;
wire n_401;
wire n_485;
wire n_1792;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_567;
wire n_369;
wire n_240;
wire n_1727;
wire n_1575;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_188;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1806;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_1696;
wire n_498;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1831;
wire n_1497;
wire n_459;
wire n_1136;
wire n_1782;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1316;
wire n_175;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_1781;
wire n_709;
wire n_809;
wire n_1686;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_199;
wire n_217;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_308;
wire n_1223;
wire n_201;
wire n_1768;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_948;
wire n_922;
wire n_1004;
wire n_1810;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_1764;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_196;
wire n_1337;
wire n_774;
wire n_933;
wire n_1779;
wire n_596;
wire n_954;
wire n_1168;
wire n_1821;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_252;
wire n_664;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1732;
wire n_415;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1799;
wire n_1126;
wire n_195;
wire n_938;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_946;
wire n_757;
wire n_375;
wire n_1655;
wire n_1818;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_265;
wire n_1583;
wire n_1604;
wire n_208;
wire n_1631;
wire n_1702;
wire n_174;
wire n_275;
wire n_1794;
wire n_1375;
wire n_204;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_1827;
wire n_866;
wire n_246;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_1569;
wire n_289;
wire n_548;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_177;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1228;
wire n_1244;
wire n_1796;
wire n_484;
wire n_411;
wire n_849;
wire n_1820;
wire n_357;
wire n_412;
wire n_1251;
wire n_447;
wire n_1421;
wire n_1762;
wire n_1233;
wire n_1808;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_56),
.Y(n_169)
);

HB1xp67_ASAP7_75t_L g170 ( 
.A(n_121),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_71),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_115),
.Y(n_172)
);

INVxp33_ASAP7_75t_SL g173 ( 
.A(n_112),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_21),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_79),
.Y(n_175)
);

BUFx10_ASAP7_75t_L g176 ( 
.A(n_161),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_55),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_95),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_130),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_141),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_80),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_143),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g183 ( 
.A(n_54),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_140),
.Y(n_184)
);

INVx2_ASAP7_75t_SL g185 ( 
.A(n_109),
.Y(n_185)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_47),
.Y(n_186)
);

BUFx3_ASAP7_75t_L g187 ( 
.A(n_55),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_84),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_167),
.Y(n_189)
);

BUFx3_ASAP7_75t_L g190 ( 
.A(n_59),
.Y(n_190)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_113),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_86),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_123),
.Y(n_193)
);

INVx2_ASAP7_75t_SL g194 ( 
.A(n_107),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_62),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_99),
.Y(n_196)
);

CKINVDCx16_ASAP7_75t_R g197 ( 
.A(n_26),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_96),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_83),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_152),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_11),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_110),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_129),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_153),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_159),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_59),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_100),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_147),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_50),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_50),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_97),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_63),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_11),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_19),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_135),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_144),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_114),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_88),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_10),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_23),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_43),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_68),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_42),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_146),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_49),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_8),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_74),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_150),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_128),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_165),
.Y(n_230)
);

BUFx3_ASAP7_75t_L g231 ( 
.A(n_26),
.Y(n_231)
);

CKINVDCx16_ASAP7_75t_R g232 ( 
.A(n_30),
.Y(n_232)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_117),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_73),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_91),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_31),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_3),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_116),
.Y(n_238)
);

INVxp67_ASAP7_75t_L g239 ( 
.A(n_1),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_82),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_77),
.Y(n_241)
);

BUFx5_ASAP7_75t_L g242 ( 
.A(n_15),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_2),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_3),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_33),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_162),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_40),
.Y(n_247)
);

HB1xp67_ASAP7_75t_L g248 ( 
.A(n_28),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_36),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_131),
.Y(n_250)
);

INVxp67_ASAP7_75t_L g251 ( 
.A(n_53),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_22),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_106),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_132),
.Y(n_254)
);

INVx1_ASAP7_75t_SL g255 ( 
.A(n_31),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_104),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_76),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_23),
.Y(n_258)
);

INVxp67_ASAP7_75t_L g259 ( 
.A(n_52),
.Y(n_259)
);

INVx1_ASAP7_75t_SL g260 ( 
.A(n_102),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_25),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_63),
.Y(n_262)
);

BUFx6f_ASAP7_75t_L g263 ( 
.A(n_119),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_148),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_22),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_4),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_101),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_154),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_92),
.Y(n_269)
);

BUFx10_ASAP7_75t_L g270 ( 
.A(n_75),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_52),
.Y(n_271)
);

CKINVDCx16_ASAP7_75t_R g272 ( 
.A(n_6),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_137),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_13),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_29),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_160),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_58),
.Y(n_277)
);

INVxp67_ASAP7_75t_SL g278 ( 
.A(n_66),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_36),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_13),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_142),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_40),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_8),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_2),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_45),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_45),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_168),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_27),
.Y(n_288)
);

INVx2_ASAP7_75t_SL g289 ( 
.A(n_25),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_149),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_1),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_134),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_78),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_49),
.Y(n_294)
);

INVx1_ASAP7_75t_SL g295 ( 
.A(n_5),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_118),
.Y(n_296)
);

INVx2_ASAP7_75t_SL g297 ( 
.A(n_18),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_14),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_28),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_67),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_38),
.Y(n_301)
);

BUFx2_ASAP7_75t_L g302 ( 
.A(n_72),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_124),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_6),
.Y(n_304)
);

BUFx3_ASAP7_75t_L g305 ( 
.A(n_16),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_32),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_145),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_120),
.Y(n_308)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_53),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_93),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_17),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_66),
.Y(n_312)
);

INVx1_ASAP7_75t_SL g313 ( 
.A(n_122),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_166),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_38),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_51),
.Y(n_316)
);

BUFx6f_ASAP7_75t_L g317 ( 
.A(n_164),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_7),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_90),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_139),
.Y(n_320)
);

INVx1_ASAP7_75t_SL g321 ( 
.A(n_87),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_155),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_9),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_58),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_111),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_44),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_81),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_157),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_136),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_133),
.Y(n_330)
);

INVx2_ASAP7_75t_L g331 ( 
.A(n_46),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_151),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_51),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_103),
.Y(n_334)
);

HB1xp67_ASAP7_75t_L g335 ( 
.A(n_15),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_19),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_175),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_216),
.Y(n_338)
);

INVx2_ASAP7_75t_L g339 ( 
.A(n_242),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_222),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_242),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_242),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_224),
.Y(n_343)
);

BUFx3_ASAP7_75t_L g344 ( 
.A(n_302),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_242),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_267),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_242),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_273),
.Y(n_348)
);

CKINVDCx16_ASAP7_75t_R g349 ( 
.A(n_197),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_242),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_307),
.Y(n_351)
);

INVx2_ASAP7_75t_L g352 ( 
.A(n_242),
.Y(n_352)
);

CKINVDCx20_ASAP7_75t_R g353 ( 
.A(n_322),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_329),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_197),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_242),
.Y(n_356)
);

INVx2_ASAP7_75t_L g357 ( 
.A(n_242),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_171),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_171),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_180),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_180),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_181),
.Y(n_362)
);

CKINVDCx20_ASAP7_75t_R g363 ( 
.A(n_169),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_181),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_182),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_182),
.Y(n_366)
);

INVxp33_ASAP7_75t_L g367 ( 
.A(n_248),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_188),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_188),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_200),
.Y(n_370)
);

CKINVDCx20_ASAP7_75t_R g371 ( 
.A(n_213),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_232),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_200),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_232),
.Y(n_374)
);

BUFx3_ASAP7_75t_L g375 ( 
.A(n_302),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_272),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_272),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_205),
.Y(n_378)
);

CKINVDCx20_ASAP7_75t_R g379 ( 
.A(n_277),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_205),
.Y(n_380)
);

HB1xp67_ASAP7_75t_L g381 ( 
.A(n_335),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_174),
.Y(n_382)
);

BUFx6f_ASAP7_75t_L g383 ( 
.A(n_263),
.Y(n_383)
);

BUFx2_ASAP7_75t_L g384 ( 
.A(n_190),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_211),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_211),
.Y(n_386)
);

INVxp67_ASAP7_75t_L g387 ( 
.A(n_195),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_177),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_201),
.Y(n_389)
);

CKINVDCx20_ASAP7_75t_R g390 ( 
.A(n_286),
.Y(n_390)
);

CKINVDCx20_ASAP7_75t_R g391 ( 
.A(n_176),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_217),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_217),
.Y(n_393)
);

CKINVDCx20_ASAP7_75t_R g394 ( 
.A(n_176),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_230),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_230),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_209),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_235),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_212),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_235),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_214),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_238),
.Y(n_402)
);

BUFx2_ASAP7_75t_L g403 ( 
.A(n_190),
.Y(n_403)
);

BUFx2_ASAP7_75t_L g404 ( 
.A(n_231),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_238),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_220),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_225),
.Y(n_407)
);

CKINVDCx16_ASAP7_75t_R g408 ( 
.A(n_176),
.Y(n_408)
);

OR2x2_ASAP7_75t_L g409 ( 
.A(n_186),
.B(n_0),
.Y(n_409)
);

INVxp33_ASAP7_75t_L g410 ( 
.A(n_195),
.Y(n_410)
);

CKINVDCx20_ASAP7_75t_R g411 ( 
.A(n_176),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_170),
.B(n_0),
.Y(n_412)
);

CKINVDCx20_ASAP7_75t_R g413 ( 
.A(n_270),
.Y(n_413)
);

CKINVDCx20_ASAP7_75t_R g414 ( 
.A(n_270),
.Y(n_414)
);

CKINVDCx20_ASAP7_75t_R g415 ( 
.A(n_270),
.Y(n_415)
);

CKINVDCx20_ASAP7_75t_R g416 ( 
.A(n_270),
.Y(n_416)
);

CKINVDCx20_ASAP7_75t_R g417 ( 
.A(n_236),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_240),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_341),
.Y(n_419)
);

INVx3_ASAP7_75t_L g420 ( 
.A(n_339),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_341),
.Y(n_421)
);

NAND2x1p5_ASAP7_75t_L g422 ( 
.A(n_409),
.B(n_240),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_358),
.B(n_250),
.Y(n_423)
);

BUFx6f_ASAP7_75t_L g424 ( 
.A(n_383),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_342),
.Y(n_425)
);

INVx6_ASAP7_75t_L g426 ( 
.A(n_383),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_342),
.Y(n_427)
);

INVx2_ASAP7_75t_L g428 ( 
.A(n_383),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_345),
.Y(n_429)
);

HB1xp67_ASAP7_75t_L g430 ( 
.A(n_349),
.Y(n_430)
);

NAND2xp33_ASAP7_75t_L g431 ( 
.A(n_358),
.B(n_183),
.Y(n_431)
);

INVx2_ASAP7_75t_L g432 ( 
.A(n_383),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_345),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_347),
.Y(n_434)
);

NAND2xp33_ASAP7_75t_L g435 ( 
.A(n_359),
.B(n_183),
.Y(n_435)
);

AND2x4_ASAP7_75t_L g436 ( 
.A(n_359),
.B(n_187),
.Y(n_436)
);

INVx2_ASAP7_75t_L g437 ( 
.A(n_383),
.Y(n_437)
);

BUFx6f_ASAP7_75t_L g438 ( 
.A(n_339),
.Y(n_438)
);

AND2x2_ASAP7_75t_L g439 ( 
.A(n_360),
.B(n_187),
.Y(n_439)
);

BUFx6f_ASAP7_75t_L g440 ( 
.A(n_352),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_347),
.Y(n_441)
);

BUFx6f_ASAP7_75t_L g442 ( 
.A(n_352),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_350),
.Y(n_443)
);

BUFx6f_ASAP7_75t_L g444 ( 
.A(n_357),
.Y(n_444)
);

HB1xp67_ASAP7_75t_L g445 ( 
.A(n_349),
.Y(n_445)
);

AND2x2_ASAP7_75t_L g446 ( 
.A(n_360),
.B(n_187),
.Y(n_446)
);

INVxp67_ASAP7_75t_L g447 ( 
.A(n_384),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_SL g448 ( 
.A(n_412),
.B(n_183),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_350),
.Y(n_449)
);

HB1xp67_ASAP7_75t_L g450 ( 
.A(n_355),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_356),
.Y(n_451)
);

OA21x2_ASAP7_75t_L g452 ( 
.A1(n_361),
.A2(n_257),
.B(n_250),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_361),
.B(n_362),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_362),
.B(n_257),
.Y(n_454)
);

BUFx6f_ASAP7_75t_L g455 ( 
.A(n_357),
.Y(n_455)
);

INVx5_ASAP7_75t_L g456 ( 
.A(n_384),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_364),
.B(n_268),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_364),
.B(n_268),
.Y(n_458)
);

INVx3_ASAP7_75t_L g459 ( 
.A(n_356),
.Y(n_459)
);

AND2x2_ASAP7_75t_L g460 ( 
.A(n_365),
.B(n_231),
.Y(n_460)
);

BUFx6f_ASAP7_75t_L g461 ( 
.A(n_365),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_SL g462 ( 
.A(n_408),
.B(n_183),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_366),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_366),
.B(n_308),
.Y(n_464)
);

BUFx6f_ASAP7_75t_L g465 ( 
.A(n_368),
.Y(n_465)
);

CKINVDCx8_ASAP7_75t_R g466 ( 
.A(n_340),
.Y(n_466)
);

BUFx6f_ASAP7_75t_L g467 ( 
.A(n_368),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_369),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_369),
.Y(n_469)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_370),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_370),
.Y(n_471)
);

NOR2xp33_ASAP7_75t_L g472 ( 
.A(n_344),
.B(n_173),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_373),
.Y(n_473)
);

AND2x2_ASAP7_75t_L g474 ( 
.A(n_373),
.B(n_305),
.Y(n_474)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_378),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_378),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_380),
.Y(n_477)
);

NOR2xp33_ASAP7_75t_SL g478 ( 
.A(n_391),
.B(n_255),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_380),
.Y(n_479)
);

INVx2_ASAP7_75t_L g480 ( 
.A(n_385),
.Y(n_480)
);

AND2x2_ASAP7_75t_L g481 ( 
.A(n_385),
.B(n_305),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_386),
.Y(n_482)
);

AND2x2_ASAP7_75t_L g483 ( 
.A(n_386),
.B(n_186),
.Y(n_483)
);

NOR2xp33_ASAP7_75t_L g484 ( 
.A(n_344),
.B(n_308),
.Y(n_484)
);

INVx2_ASAP7_75t_L g485 ( 
.A(n_392),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_392),
.Y(n_486)
);

HB1xp67_ASAP7_75t_L g487 ( 
.A(n_372),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_393),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_393),
.B(n_310),
.Y(n_489)
);

BUFx6f_ASAP7_75t_L g490 ( 
.A(n_395),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_395),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_396),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_461),
.Y(n_493)
);

INVx2_ASAP7_75t_SL g494 ( 
.A(n_456),
.Y(n_494)
);

INVx3_ASAP7_75t_L g495 ( 
.A(n_461),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_SL g496 ( 
.A(n_456),
.B(n_382),
.Y(n_496)
);

BUFx4f_ASAP7_75t_L g497 ( 
.A(n_452),
.Y(n_497)
);

INVxp67_ASAP7_75t_SL g498 ( 
.A(n_453),
.Y(n_498)
);

OR2x2_ASAP7_75t_L g499 ( 
.A(n_447),
.B(n_381),
.Y(n_499)
);

INVx4_ASAP7_75t_L g500 ( 
.A(n_461),
.Y(n_500)
);

INVx2_ASAP7_75t_L g501 ( 
.A(n_420),
.Y(n_501)
);

INVx3_ASAP7_75t_L g502 ( 
.A(n_461),
.Y(n_502)
);

AND2x2_ASAP7_75t_L g503 ( 
.A(n_483),
.B(n_410),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_461),
.Y(n_504)
);

INVx3_ASAP7_75t_L g505 ( 
.A(n_461),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_SL g506 ( 
.A(n_456),
.B(n_388),
.Y(n_506)
);

AND2x2_ASAP7_75t_SL g507 ( 
.A(n_452),
.B(n_409),
.Y(n_507)
);

AND2x2_ASAP7_75t_L g508 ( 
.A(n_483),
.B(n_403),
.Y(n_508)
);

BUFx3_ASAP7_75t_L g509 ( 
.A(n_419),
.Y(n_509)
);

NOR2xp33_ASAP7_75t_L g510 ( 
.A(n_462),
.B(n_389),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g511 ( 
.A(n_422),
.B(n_375),
.Y(n_511)
);

BUFx2_ASAP7_75t_L g512 ( 
.A(n_430),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_SL g513 ( 
.A(n_456),
.B(n_397),
.Y(n_513)
);

CKINVDCx6p67_ASAP7_75t_R g514 ( 
.A(n_430),
.Y(n_514)
);

BUFx3_ASAP7_75t_L g515 ( 
.A(n_419),
.Y(n_515)
);

BUFx3_ASAP7_75t_L g516 ( 
.A(n_421),
.Y(n_516)
);

INVx2_ASAP7_75t_SL g517 ( 
.A(n_456),
.Y(n_517)
);

BUFx6f_ASAP7_75t_L g518 ( 
.A(n_438),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_461),
.Y(n_519)
);

AOI22xp33_ASAP7_75t_L g520 ( 
.A1(n_422),
.A2(n_375),
.B1(n_367),
.B2(n_396),
.Y(n_520)
);

AND2x2_ASAP7_75t_L g521 ( 
.A(n_483),
.B(n_403),
.Y(n_521)
);

INVx4_ASAP7_75t_L g522 ( 
.A(n_461),
.Y(n_522)
);

INVx4_ASAP7_75t_L g523 ( 
.A(n_465),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_SL g524 ( 
.A(n_456),
.B(n_399),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_465),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_422),
.B(n_398),
.Y(n_526)
);

INVx5_ASAP7_75t_L g527 ( 
.A(n_424),
.Y(n_527)
);

INVx5_ASAP7_75t_L g528 ( 
.A(n_424),
.Y(n_528)
);

AND2x6_ASAP7_75t_L g529 ( 
.A(n_475),
.B(n_310),
.Y(n_529)
);

INVx2_ASAP7_75t_L g530 ( 
.A(n_420),
.Y(n_530)
);

INVx2_ASAP7_75t_L g531 ( 
.A(n_420),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_465),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_422),
.B(n_398),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_L g534 ( 
.A(n_456),
.B(n_463),
.Y(n_534)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_420),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_465),
.Y(n_536)
);

BUFx6f_ASAP7_75t_L g537 ( 
.A(n_438),
.Y(n_537)
);

AOI22xp5_ASAP7_75t_L g538 ( 
.A1(n_484),
.A2(n_295),
.B1(n_278),
.B2(n_289),
.Y(n_538)
);

BUFx6f_ASAP7_75t_L g539 ( 
.A(n_438),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_SL g540 ( 
.A(n_456),
.B(n_401),
.Y(n_540)
);

BUFx8_ASAP7_75t_SL g541 ( 
.A(n_466),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_SL g542 ( 
.A(n_472),
.B(n_406),
.Y(n_542)
);

INVx2_ASAP7_75t_L g543 ( 
.A(n_420),
.Y(n_543)
);

AOI22xp5_ASAP7_75t_L g544 ( 
.A1(n_484),
.A2(n_289),
.B1(n_297),
.B2(n_259),
.Y(n_544)
);

BUFx3_ASAP7_75t_L g545 ( 
.A(n_421),
.Y(n_545)
);

INVx2_ASAP7_75t_SL g546 ( 
.A(n_462),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_465),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_SL g548 ( 
.A(n_472),
.B(n_407),
.Y(n_548)
);

NAND2xp33_ASAP7_75t_L g549 ( 
.A(n_465),
.B(n_183),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_465),
.Y(n_550)
);

OAI22xp33_ASAP7_75t_L g551 ( 
.A1(n_478),
.A2(n_377),
.B1(n_376),
.B2(n_374),
.Y(n_551)
);

AND2x6_ASAP7_75t_L g552 ( 
.A(n_475),
.B(n_314),
.Y(n_552)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_459),
.Y(n_553)
);

NOR2xp33_ASAP7_75t_L g554 ( 
.A(n_447),
.B(n_463),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_465),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_467),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_SL g557 ( 
.A(n_450),
.B(n_417),
.Y(n_557)
);

INVx4_ASAP7_75t_L g558 ( 
.A(n_467),
.Y(n_558)
);

BUFx4f_ASAP7_75t_L g559 ( 
.A(n_452),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_467),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_467),
.Y(n_561)
);

BUFx10_ASAP7_75t_L g562 ( 
.A(n_450),
.Y(n_562)
);

OR2x6_ASAP7_75t_L g563 ( 
.A(n_445),
.B(n_297),
.Y(n_563)
);

NOR2xp33_ASAP7_75t_L g564 ( 
.A(n_468),
.B(n_394),
.Y(n_564)
);

NAND2xp33_ASAP7_75t_L g565 ( 
.A(n_467),
.B(n_183),
.Y(n_565)
);

BUFx3_ASAP7_75t_L g566 ( 
.A(n_425),
.Y(n_566)
);

AND2x6_ASAP7_75t_L g567 ( 
.A(n_475),
.B(n_314),
.Y(n_567)
);

INVx2_ASAP7_75t_L g568 ( 
.A(n_459),
.Y(n_568)
);

BUFx4f_ASAP7_75t_L g569 ( 
.A(n_452),
.Y(n_569)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_459),
.Y(n_570)
);

AND2x6_ASAP7_75t_L g571 ( 
.A(n_475),
.B(n_325),
.Y(n_571)
);

OR2x6_ASAP7_75t_L g572 ( 
.A(n_445),
.B(n_400),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_467),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_L g574 ( 
.A(n_468),
.B(n_400),
.Y(n_574)
);

BUFx6f_ASAP7_75t_L g575 ( 
.A(n_438),
.Y(n_575)
);

INVx2_ASAP7_75t_L g576 ( 
.A(n_459),
.Y(n_576)
);

AND2x6_ASAP7_75t_L g577 ( 
.A(n_470),
.B(n_325),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_L g578 ( 
.A(n_469),
.B(n_402),
.Y(n_578)
);

BUFx6f_ASAP7_75t_L g579 ( 
.A(n_438),
.Y(n_579)
);

AND3x2_ASAP7_75t_L g580 ( 
.A(n_478),
.B(n_404),
.C(n_251),
.Y(n_580)
);

BUFx3_ASAP7_75t_L g581 ( 
.A(n_425),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_467),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_L g583 ( 
.A(n_469),
.B(n_402),
.Y(n_583)
);

INVx2_ASAP7_75t_SL g584 ( 
.A(n_439),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_L g585 ( 
.A(n_471),
.B(n_405),
.Y(n_585)
);

AOI22xp33_ASAP7_75t_L g586 ( 
.A1(n_452),
.A2(n_418),
.B1(n_405),
.B2(n_415),
.Y(n_586)
);

AND2x2_ASAP7_75t_L g587 ( 
.A(n_460),
.B(n_474),
.Y(n_587)
);

INVx2_ASAP7_75t_L g588 ( 
.A(n_459),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_467),
.Y(n_589)
);

NOR3xp33_ASAP7_75t_L g590 ( 
.A(n_487),
.B(n_239),
.C(n_387),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_490),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_490),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_490),
.Y(n_593)
);

INVx3_ASAP7_75t_L g594 ( 
.A(n_490),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_427),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_SL g596 ( 
.A(n_487),
.B(n_343),
.Y(n_596)
);

AOI21x1_ASAP7_75t_L g597 ( 
.A1(n_427),
.A2(n_418),
.B(n_233),
.Y(n_597)
);

INVx2_ASAP7_75t_L g598 ( 
.A(n_429),
.Y(n_598)
);

XOR2x2_ASAP7_75t_L g599 ( 
.A(n_466),
.B(n_363),
.Y(n_599)
);

AND3x2_ASAP7_75t_L g600 ( 
.A(n_460),
.B(n_404),
.C(n_210),
.Y(n_600)
);

INVx3_ASAP7_75t_L g601 ( 
.A(n_490),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_471),
.B(n_473),
.Y(n_602)
);

XNOR2xp5_ASAP7_75t_L g603 ( 
.A(n_466),
.B(n_371),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_490),
.Y(n_604)
);

INVx4_ASAP7_75t_L g605 ( 
.A(n_490),
.Y(n_605)
);

AND2x2_ASAP7_75t_L g606 ( 
.A(n_460),
.B(n_206),
.Y(n_606)
);

AND2x2_ASAP7_75t_L g607 ( 
.A(n_474),
.B(n_206),
.Y(n_607)
);

AOI22xp33_ASAP7_75t_L g608 ( 
.A1(n_452),
.A2(n_416),
.B1(n_414),
.B2(n_413),
.Y(n_608)
);

INVx2_ASAP7_75t_L g609 ( 
.A(n_429),
.Y(n_609)
);

INVx2_ASAP7_75t_SL g610 ( 
.A(n_439),
.Y(n_610)
);

INVx1_ASAP7_75t_SL g611 ( 
.A(n_474),
.Y(n_611)
);

INVx1_ASAP7_75t_SL g612 ( 
.A(n_481),
.Y(n_612)
);

BUFx6f_ASAP7_75t_L g613 ( 
.A(n_438),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_490),
.Y(n_614)
);

INVx2_ASAP7_75t_L g615 ( 
.A(n_433),
.Y(n_615)
);

OR2x2_ASAP7_75t_L g616 ( 
.A(n_453),
.B(n_346),
.Y(n_616)
);

INVx8_ASAP7_75t_L g617 ( 
.A(n_436),
.Y(n_617)
);

INVx4_ASAP7_75t_L g618 ( 
.A(n_438),
.Y(n_618)
);

OR2x6_ASAP7_75t_L g619 ( 
.A(n_436),
.B(n_309),
.Y(n_619)
);

INVx8_ASAP7_75t_L g620 ( 
.A(n_436),
.Y(n_620)
);

AND2x6_ASAP7_75t_L g621 ( 
.A(n_470),
.B(n_191),
.Y(n_621)
);

INVx2_ASAP7_75t_L g622 ( 
.A(n_433),
.Y(n_622)
);

INVx2_ASAP7_75t_L g623 ( 
.A(n_434),
.Y(n_623)
);

INVx2_ASAP7_75t_L g624 ( 
.A(n_434),
.Y(n_624)
);

AOI22xp33_ASAP7_75t_L g625 ( 
.A1(n_436),
.A2(n_411),
.B1(n_309),
.B2(n_331),
.Y(n_625)
);

INVxp67_ASAP7_75t_SL g626 ( 
.A(n_438),
.Y(n_626)
);

INVx2_ASAP7_75t_L g627 ( 
.A(n_441),
.Y(n_627)
);

BUFx3_ASAP7_75t_L g628 ( 
.A(n_441),
.Y(n_628)
);

AND2x2_ASAP7_75t_L g629 ( 
.A(n_481),
.B(n_210),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_470),
.Y(n_630)
);

INVx2_ASAP7_75t_L g631 ( 
.A(n_443),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g632 ( 
.A(n_473),
.B(n_260),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_480),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_SL g634 ( 
.A(n_436),
.B(n_348),
.Y(n_634)
);

INVx2_ASAP7_75t_L g635 ( 
.A(n_443),
.Y(n_635)
);

NOR2x1p5_ASAP7_75t_L g636 ( 
.A(n_423),
.B(n_351),
.Y(n_636)
);

INVx2_ASAP7_75t_L g637 ( 
.A(n_449),
.Y(n_637)
);

AND2x2_ASAP7_75t_L g638 ( 
.A(n_481),
.B(n_219),
.Y(n_638)
);

AND3x2_ASAP7_75t_L g639 ( 
.A(n_439),
.B(n_221),
.C(n_219),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_480),
.Y(n_640)
);

AND2x2_ASAP7_75t_L g641 ( 
.A(n_446),
.B(n_221),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_480),
.Y(n_642)
);

NAND3xp33_ASAP7_75t_L g643 ( 
.A(n_476),
.B(n_226),
.C(n_223),
.Y(n_643)
);

INVx2_ASAP7_75t_L g644 ( 
.A(n_595),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_SL g645 ( 
.A(n_497),
.B(n_449),
.Y(n_645)
);

NOR2xp33_ASAP7_75t_SL g646 ( 
.A(n_541),
.B(n_354),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_SL g647 ( 
.A(n_497),
.B(n_451),
.Y(n_647)
);

INVx2_ASAP7_75t_SL g648 ( 
.A(n_572),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_498),
.B(n_476),
.Y(n_649)
);

AOI22xp5_ASAP7_75t_L g650 ( 
.A1(n_510),
.A2(n_448),
.B1(n_491),
.B2(n_482),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_SL g651 ( 
.A(n_497),
.B(n_451),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_554),
.B(n_477),
.Y(n_652)
);

INVx2_ASAP7_75t_SL g653 ( 
.A(n_572),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_L g654 ( 
.A(n_526),
.B(n_477),
.Y(n_654)
);

OR2x6_ASAP7_75t_L g655 ( 
.A(n_572),
.B(n_446),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_509),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_L g657 ( 
.A(n_533),
.B(n_479),
.Y(n_657)
);

AND2x4_ASAP7_75t_L g658 ( 
.A(n_619),
.B(n_446),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_SL g659 ( 
.A(n_559),
.B(n_479),
.Y(n_659)
);

NAND2xp33_ASAP7_75t_L g660 ( 
.A(n_617),
.B(n_482),
.Y(n_660)
);

INVxp67_ASAP7_75t_SL g661 ( 
.A(n_559),
.Y(n_661)
);

INVx2_ASAP7_75t_L g662 ( 
.A(n_595),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_509),
.Y(n_663)
);

INVx2_ASAP7_75t_L g664 ( 
.A(n_598),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_515),
.Y(n_665)
);

BUFx6f_ASAP7_75t_SL g666 ( 
.A(n_562),
.Y(n_666)
);

NOR2xp33_ASAP7_75t_L g667 ( 
.A(n_546),
.B(n_448),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_515),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_546),
.B(n_486),
.Y(n_669)
);

NAND2xp33_ASAP7_75t_L g670 ( 
.A(n_617),
.B(n_486),
.Y(n_670)
);

AOI22xp33_ASAP7_75t_L g671 ( 
.A1(n_507),
.A2(n_491),
.B1(n_488),
.B2(n_492),
.Y(n_671)
);

NOR2xp33_ASAP7_75t_L g672 ( 
.A(n_616),
.B(n_488),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_SL g673 ( 
.A(n_559),
.B(n_492),
.Y(n_673)
);

INVx8_ASAP7_75t_L g674 ( 
.A(n_617),
.Y(n_674)
);

O2A1O1Ixp33_ASAP7_75t_L g675 ( 
.A1(n_584),
.A2(n_489),
.B(n_464),
.C(n_458),
.Y(n_675)
);

NOR2xp33_ASAP7_75t_L g676 ( 
.A(n_616),
.B(n_485),
.Y(n_676)
);

AND2x2_ASAP7_75t_L g677 ( 
.A(n_503),
.B(n_337),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_L g678 ( 
.A(n_611),
.B(n_485),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_SL g679 ( 
.A(n_569),
.B(n_440),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_SL g680 ( 
.A(n_569),
.B(n_440),
.Y(n_680)
);

INVx4_ASAP7_75t_L g681 ( 
.A(n_617),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_L g682 ( 
.A(n_611),
.B(n_485),
.Y(n_682)
);

INVx2_ASAP7_75t_L g683 ( 
.A(n_598),
.Y(n_683)
);

INVxp67_ASAP7_75t_SL g684 ( 
.A(n_569),
.Y(n_684)
);

INVx2_ASAP7_75t_L g685 ( 
.A(n_609),
.Y(n_685)
);

BUFx3_ASAP7_75t_L g686 ( 
.A(n_617),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_516),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_L g688 ( 
.A(n_584),
.B(n_423),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_L g689 ( 
.A(n_610),
.B(n_454),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_SL g690 ( 
.A(n_507),
.B(n_440),
.Y(n_690)
);

INVx2_ASAP7_75t_L g691 ( 
.A(n_609),
.Y(n_691)
);

AOI22xp5_ASAP7_75t_L g692 ( 
.A1(n_507),
.A2(n_489),
.B1(n_464),
.B2(n_458),
.Y(n_692)
);

OAI22xp5_ASAP7_75t_L g693 ( 
.A1(n_516),
.A2(n_457),
.B1(n_454),
.B2(n_243),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_L g694 ( 
.A(n_610),
.B(n_457),
.Y(n_694)
);

OR2x6_ASAP7_75t_L g695 ( 
.A(n_572),
.B(n_338),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_L g696 ( 
.A(n_586),
.B(n_440),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_612),
.B(n_440),
.Y(n_697)
);

OR2x2_ASAP7_75t_L g698 ( 
.A(n_499),
.B(n_353),
.Y(n_698)
);

INVx2_ASAP7_75t_L g699 ( 
.A(n_615),
.Y(n_699)
);

AOI21xp5_ASAP7_75t_L g700 ( 
.A1(n_626),
.A2(n_442),
.B(n_440),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_SL g701 ( 
.A(n_553),
.B(n_440),
.Y(n_701)
);

INVx3_ASAP7_75t_L g702 ( 
.A(n_620),
.Y(n_702)
);

INVx3_ASAP7_75t_L g703 ( 
.A(n_620),
.Y(n_703)
);

AOI22xp33_ASAP7_75t_L g704 ( 
.A1(n_538),
.A2(n_619),
.B1(n_625),
.B2(n_566),
.Y(n_704)
);

NOR2xp33_ASAP7_75t_L g705 ( 
.A(n_511),
.B(n_440),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_L g706 ( 
.A(n_632),
.B(n_442),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_503),
.B(n_442),
.Y(n_707)
);

BUFx3_ASAP7_75t_L g708 ( 
.A(n_620),
.Y(n_708)
);

INVx2_ASAP7_75t_L g709 ( 
.A(n_615),
.Y(n_709)
);

INVx3_ASAP7_75t_L g710 ( 
.A(n_620),
.Y(n_710)
);

INVx3_ASAP7_75t_L g711 ( 
.A(n_620),
.Y(n_711)
);

AND2x2_ASAP7_75t_L g712 ( 
.A(n_572),
.B(n_564),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_L g713 ( 
.A(n_587),
.B(n_442),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_SL g714 ( 
.A(n_553),
.B(n_442),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_L g715 ( 
.A(n_587),
.B(n_442),
.Y(n_715)
);

AND2x2_ASAP7_75t_L g716 ( 
.A(n_499),
.B(n_379),
.Y(n_716)
);

INVx2_ASAP7_75t_L g717 ( 
.A(n_622),
.Y(n_717)
);

AND2x2_ASAP7_75t_L g718 ( 
.A(n_512),
.B(n_390),
.Y(n_718)
);

NAND3xp33_ASAP7_75t_L g719 ( 
.A(n_520),
.B(n_244),
.C(n_237),
.Y(n_719)
);

AOI22xp33_ASAP7_75t_L g720 ( 
.A1(n_538),
.A2(n_331),
.B1(n_444),
.B2(n_442),
.Y(n_720)
);

INVxp67_ASAP7_75t_L g721 ( 
.A(n_512),
.Y(n_721)
);

NOR2xp33_ASAP7_75t_L g722 ( 
.A(n_542),
.B(n_442),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_L g723 ( 
.A(n_545),
.B(n_444),
.Y(n_723)
);

INVx2_ASAP7_75t_L g724 ( 
.A(n_622),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_L g725 ( 
.A(n_545),
.B(n_444),
.Y(n_725)
);

INVx2_ASAP7_75t_L g726 ( 
.A(n_623),
.Y(n_726)
);

HB1xp67_ASAP7_75t_L g727 ( 
.A(n_563),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_L g728 ( 
.A(n_566),
.B(n_444),
.Y(n_728)
);

INVx8_ASAP7_75t_L g729 ( 
.A(n_563),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_SL g730 ( 
.A(n_568),
.B(n_444),
.Y(n_730)
);

BUFx6f_ASAP7_75t_SL g731 ( 
.A(n_562),
.Y(n_731)
);

AND2x2_ASAP7_75t_L g732 ( 
.A(n_508),
.B(n_223),
.Y(n_732)
);

NOR2xp33_ASAP7_75t_L g733 ( 
.A(n_548),
.B(n_444),
.Y(n_733)
);

NOR3xp33_ASAP7_75t_L g734 ( 
.A(n_557),
.B(n_590),
.C(n_596),
.Y(n_734)
);

INVxp33_ASAP7_75t_L g735 ( 
.A(n_603),
.Y(n_735)
);

OAI22xp5_ASAP7_75t_L g736 ( 
.A1(n_581),
.A2(n_271),
.B1(n_336),
.B2(n_252),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_581),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_628),
.Y(n_738)
);

AND2x2_ASAP7_75t_L g739 ( 
.A(n_508),
.B(n_226),
.Y(n_739)
);

INVx2_ASAP7_75t_L g740 ( 
.A(n_623),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_SL g741 ( 
.A(n_568),
.B(n_444),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_628),
.Y(n_742)
);

INVxp67_ASAP7_75t_L g743 ( 
.A(n_603),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_L g744 ( 
.A(n_641),
.B(n_444),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_L g745 ( 
.A(n_641),
.B(n_455),
.Y(n_745)
);

NOR2xp33_ASAP7_75t_L g746 ( 
.A(n_634),
.B(n_455),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_606),
.B(n_455),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_SL g748 ( 
.A(n_570),
.B(n_455),
.Y(n_748)
);

NOR2xp33_ASAP7_75t_L g749 ( 
.A(n_619),
.B(n_455),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_602),
.Y(n_750)
);

INVx8_ASAP7_75t_L g751 ( 
.A(n_563),
.Y(n_751)
);

NOR2xp33_ASAP7_75t_SL g752 ( 
.A(n_514),
.B(n_313),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_630),
.Y(n_753)
);

AND2x2_ASAP7_75t_L g754 ( 
.A(n_521),
.B(n_247),
.Y(n_754)
);

INVx2_ASAP7_75t_L g755 ( 
.A(n_624),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_SL g756 ( 
.A(n_570),
.B(n_455),
.Y(n_756)
);

NAND2x1p5_ASAP7_75t_L g757 ( 
.A(n_494),
.B(n_321),
.Y(n_757)
);

BUFx3_ASAP7_75t_L g758 ( 
.A(n_562),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_606),
.B(n_455),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_630),
.Y(n_760)
);

INVx2_ASAP7_75t_SL g761 ( 
.A(n_562),
.Y(n_761)
);

NAND3xp33_ASAP7_75t_L g762 ( 
.A(n_544),
.B(n_258),
.C(n_245),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_607),
.B(n_629),
.Y(n_763)
);

AND2x4_ASAP7_75t_L g764 ( 
.A(n_619),
.B(n_247),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_SL g765 ( 
.A(n_576),
.B(n_588),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_607),
.B(n_455),
.Y(n_766)
);

AOI22xp33_ASAP7_75t_L g767 ( 
.A1(n_619),
.A2(n_185),
.B1(n_194),
.B2(n_431),
.Y(n_767)
);

INVxp67_ASAP7_75t_L g768 ( 
.A(n_521),
.Y(n_768)
);

INVx2_ASAP7_75t_L g769 ( 
.A(n_624),
.Y(n_769)
);

AND2x6_ASAP7_75t_L g770 ( 
.A(n_576),
.B(n_191),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_629),
.B(n_249),
.Y(n_771)
);

BUFx4f_ASAP7_75t_L g772 ( 
.A(n_514),
.Y(n_772)
);

NOR3xp33_ASAP7_75t_L g773 ( 
.A(n_551),
.B(n_265),
.C(n_249),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_L g774 ( 
.A(n_638),
.B(n_265),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_638),
.B(n_266),
.Y(n_775)
);

INVx3_ASAP7_75t_L g776 ( 
.A(n_627),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_L g777 ( 
.A(n_574),
.B(n_266),
.Y(n_777)
);

INVx2_ASAP7_75t_L g778 ( 
.A(n_627),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_633),
.Y(n_779)
);

NOR2xp33_ASAP7_75t_R g780 ( 
.A(n_580),
.B(n_431),
.Y(n_780)
);

NAND2xp33_ASAP7_75t_SL g781 ( 
.A(n_636),
.B(n_274),
.Y(n_781)
);

INVx8_ASAP7_75t_L g782 ( 
.A(n_563),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_L g783 ( 
.A(n_578),
.B(n_274),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_583),
.B(n_275),
.Y(n_784)
);

INVx2_ASAP7_75t_L g785 ( 
.A(n_631),
.Y(n_785)
);

NOR2xp33_ASAP7_75t_L g786 ( 
.A(n_588),
.B(n_261),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_L g787 ( 
.A(n_585),
.B(n_631),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_640),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_635),
.B(n_275),
.Y(n_789)
);

AND2x4_ASAP7_75t_L g790 ( 
.A(n_563),
.B(n_279),
.Y(n_790)
);

INVx2_ASAP7_75t_L g791 ( 
.A(n_635),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_640),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_642),
.Y(n_793)
);

AOI22xp5_ASAP7_75t_L g794 ( 
.A1(n_636),
.A2(n_194),
.B1(n_185),
.B2(n_229),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_L g795 ( 
.A(n_637),
.B(n_279),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_L g796 ( 
.A(n_637),
.B(n_285),
.Y(n_796)
);

AOI22xp5_ASAP7_75t_L g797 ( 
.A1(n_544),
.A2(n_203),
.B1(n_218),
.B2(n_215),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_SL g798 ( 
.A(n_518),
.B(n_233),
.Y(n_798)
);

O2A1O1Ixp33_ASAP7_75t_L g799 ( 
.A1(n_642),
.A2(n_304),
.B(n_285),
.C(n_288),
.Y(n_799)
);

CKINVDCx5p33_ASAP7_75t_R g800 ( 
.A(n_599),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_501),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_L g802 ( 
.A(n_501),
.B(n_288),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_SL g803 ( 
.A(n_518),
.B(n_263),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_SL g804 ( 
.A(n_518),
.B(n_263),
.Y(n_804)
);

AOI22xp5_ASAP7_75t_L g805 ( 
.A1(n_496),
.A2(n_198),
.B1(n_204),
.B2(n_202),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_SL g806 ( 
.A(n_518),
.B(n_263),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_L g807 ( 
.A(n_530),
.B(n_300),
.Y(n_807)
);

BUFx8_ASAP7_75t_L g808 ( 
.A(n_577),
.Y(n_808)
);

INVx2_ASAP7_75t_L g809 ( 
.A(n_530),
.Y(n_809)
);

INVx8_ASAP7_75t_L g810 ( 
.A(n_529),
.Y(n_810)
);

CKINVDCx20_ASAP7_75t_R g811 ( 
.A(n_599),
.Y(n_811)
);

NOR2xp33_ASAP7_75t_L g812 ( 
.A(n_500),
.B(n_262),
.Y(n_812)
);

NAND2x1_ASAP7_75t_L g813 ( 
.A(n_500),
.B(n_426),
.Y(n_813)
);

NOR3xp33_ASAP7_75t_L g814 ( 
.A(n_643),
.B(n_300),
.C(n_304),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_SL g815 ( 
.A(n_518),
.B(n_263),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_672),
.B(n_608),
.Y(n_816)
);

OR2x2_ASAP7_75t_L g817 ( 
.A(n_698),
.B(n_716),
.Y(n_817)
);

INVx2_ASAP7_75t_L g818 ( 
.A(n_776),
.Y(n_818)
);

AOI21xp5_ASAP7_75t_L g819 ( 
.A1(n_645),
.A2(n_534),
.B(n_618),
.Y(n_819)
);

OAI21xp5_ASAP7_75t_L g820 ( 
.A1(n_690),
.A2(n_673),
.B(n_659),
.Y(n_820)
);

A2O1A1Ixp33_ASAP7_75t_L g821 ( 
.A1(n_672),
.A2(n_643),
.B(n_311),
.C(n_306),
.Y(n_821)
);

AO21x1_ASAP7_75t_L g822 ( 
.A1(n_645),
.A2(n_597),
.B(n_522),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_753),
.Y(n_823)
);

AOI21xp5_ASAP7_75t_L g824 ( 
.A1(n_647),
.A2(n_618),
.B(n_513),
.Y(n_824)
);

INVx4_ASAP7_75t_L g825 ( 
.A(n_674),
.Y(n_825)
);

OAI21xp33_ASAP7_75t_L g826 ( 
.A1(n_652),
.A2(n_282),
.B(n_280),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_L g827 ( 
.A(n_676),
.B(n_531),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_L g828 ( 
.A(n_676),
.B(n_531),
.Y(n_828)
);

CKINVDCx16_ASAP7_75t_R g829 ( 
.A(n_646),
.Y(n_829)
);

INVx2_ASAP7_75t_L g830 ( 
.A(n_776),
.Y(n_830)
);

AOI21xp5_ASAP7_75t_L g831 ( 
.A1(n_647),
.A2(n_618),
.B(n_524),
.Y(n_831)
);

BUFx2_ASAP7_75t_L g832 ( 
.A(n_718),
.Y(n_832)
);

INVxp67_ASAP7_75t_L g833 ( 
.A(n_677),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_750),
.B(n_535),
.Y(n_834)
);

BUFx6f_ASAP7_75t_L g835 ( 
.A(n_674),
.Y(n_835)
);

OAI21xp33_ASAP7_75t_L g836 ( 
.A1(n_763),
.A2(n_284),
.B(n_283),
.Y(n_836)
);

INVx2_ASAP7_75t_L g837 ( 
.A(n_644),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_SL g838 ( 
.A(n_681),
.B(n_537),
.Y(n_838)
);

A2O1A1Ixp33_ASAP7_75t_L g839 ( 
.A1(n_692),
.A2(n_306),
.B(n_311),
.C(n_535),
.Y(n_839)
);

INVx3_ASAP7_75t_L g840 ( 
.A(n_681),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_L g841 ( 
.A(n_688),
.B(n_689),
.Y(n_841)
);

HB1xp67_ASAP7_75t_L g842 ( 
.A(n_655),
.Y(n_842)
);

OR2x2_ASAP7_75t_L g843 ( 
.A(n_721),
.B(n_543),
.Y(n_843)
);

OAI21x1_ASAP7_75t_L g844 ( 
.A1(n_679),
.A2(n_597),
.B(n_504),
.Y(n_844)
);

AOI21xp5_ASAP7_75t_L g845 ( 
.A1(n_651),
.A2(n_618),
.B(n_540),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_SL g846 ( 
.A(n_681),
.B(n_537),
.Y(n_846)
);

AOI21xp5_ASAP7_75t_L g847 ( 
.A1(n_651),
.A2(n_680),
.B(n_679),
.Y(n_847)
);

INVx3_ASAP7_75t_L g848 ( 
.A(n_674),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_694),
.B(n_543),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_760),
.Y(n_850)
);

INVx2_ASAP7_75t_L g851 ( 
.A(n_644),
.Y(n_851)
);

OAI21xp5_ASAP7_75t_L g852 ( 
.A1(n_690),
.A2(n_504),
.B(n_493),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_L g853 ( 
.A(n_678),
.B(n_600),
.Y(n_853)
);

OAI21xp33_ASAP7_75t_L g854 ( 
.A1(n_786),
.A2(n_294),
.B(n_291),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_L g855 ( 
.A(n_682),
.B(n_639),
.Y(n_855)
);

INVx3_ASAP7_75t_L g856 ( 
.A(n_686),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_648),
.B(n_494),
.Y(n_857)
);

INVx2_ASAP7_75t_L g858 ( 
.A(n_662),
.Y(n_858)
);

BUFx6f_ASAP7_75t_L g859 ( 
.A(n_686),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_L g860 ( 
.A(n_653),
.B(n_517),
.Y(n_860)
);

OR2x2_ASAP7_75t_L g861 ( 
.A(n_695),
.B(n_298),
.Y(n_861)
);

NOR2xp33_ASAP7_75t_L g862 ( 
.A(n_712),
.B(n_500),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_L g863 ( 
.A(n_704),
.B(n_517),
.Y(n_863)
);

NOR2xp33_ASAP7_75t_L g864 ( 
.A(n_768),
.B(n_500),
.Y(n_864)
);

AOI21xp5_ASAP7_75t_L g865 ( 
.A1(n_680),
.A2(n_506),
.B(n_493),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_L g866 ( 
.A(n_649),
.B(n_522),
.Y(n_866)
);

AOI21xp5_ASAP7_75t_L g867 ( 
.A1(n_659),
.A2(n_673),
.B(n_765),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_SL g868 ( 
.A(n_702),
.B(n_537),
.Y(n_868)
);

BUFx3_ASAP7_75t_L g869 ( 
.A(n_708),
.Y(n_869)
);

AOI21xp5_ASAP7_75t_L g870 ( 
.A1(n_765),
.A2(n_700),
.B(n_787),
.Y(n_870)
);

OAI22xp5_ASAP7_75t_L g871 ( 
.A1(n_671),
.A2(n_523),
.B1(n_522),
.B2(n_558),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_SL g872 ( 
.A(n_702),
.B(n_537),
.Y(n_872)
);

INVxp67_ASAP7_75t_L g873 ( 
.A(n_752),
.Y(n_873)
);

AOI21xp5_ASAP7_75t_L g874 ( 
.A1(n_654),
.A2(n_525),
.B(n_519),
.Y(n_874)
);

AOI21xp5_ASAP7_75t_L g875 ( 
.A1(n_657),
.A2(n_525),
.B(n_519),
.Y(n_875)
);

NOR2xp33_ASAP7_75t_SL g876 ( 
.A(n_772),
.B(n_529),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_L g877 ( 
.A(n_707),
.B(n_522),
.Y(n_877)
);

OAI21xp5_ASAP7_75t_L g878 ( 
.A1(n_713),
.A2(n_536),
.B(n_532),
.Y(n_878)
);

AOI22xp5_ASAP7_75t_L g879 ( 
.A1(n_655),
.A2(n_523),
.B1(n_558),
.B2(n_605),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_SL g880 ( 
.A(n_703),
.B(n_537),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_779),
.Y(n_881)
);

A2O1A1Ixp33_ASAP7_75t_L g882 ( 
.A1(n_675),
.A2(n_556),
.B(n_614),
.C(n_550),
.Y(n_882)
);

AOI21xp5_ASAP7_75t_L g883 ( 
.A1(n_701),
.A2(n_536),
.B(n_532),
.Y(n_883)
);

AND2x2_ASAP7_75t_L g884 ( 
.A(n_732),
.B(n_299),
.Y(n_884)
);

OAI21xp5_ASAP7_75t_L g885 ( 
.A1(n_715),
.A2(n_745),
.B(n_744),
.Y(n_885)
);

AOI21xp5_ASAP7_75t_L g886 ( 
.A1(n_701),
.A2(n_550),
.B(n_547),
.Y(n_886)
);

AOI21xp5_ASAP7_75t_L g887 ( 
.A1(n_714),
.A2(n_741),
.B(n_730),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_658),
.B(n_523),
.Y(n_888)
);

CKINVDCx5p33_ASAP7_75t_R g889 ( 
.A(n_772),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_L g890 ( 
.A(n_658),
.B(n_523),
.Y(n_890)
);

AOI21xp5_ASAP7_75t_L g891 ( 
.A1(n_714),
.A2(n_555),
.B(n_547),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_788),
.Y(n_892)
);

AOI21xp5_ASAP7_75t_L g893 ( 
.A1(n_730),
.A2(n_556),
.B(n_555),
.Y(n_893)
);

NAND2x1p5_ASAP7_75t_L g894 ( 
.A(n_708),
.B(n_558),
.Y(n_894)
);

NOR2xp33_ASAP7_75t_L g895 ( 
.A(n_655),
.B(n_558),
.Y(n_895)
);

A2O1A1Ixp33_ASAP7_75t_L g896 ( 
.A1(n_773),
.A2(n_591),
.B(n_614),
.C(n_573),
.Y(n_896)
);

AOI21xp5_ASAP7_75t_L g897 ( 
.A1(n_741),
.A2(n_561),
.B(n_560),
.Y(n_897)
);

NOR2xp33_ASAP7_75t_L g898 ( 
.A(n_656),
.B(n_605),
.Y(n_898)
);

AOI21x1_ASAP7_75t_L g899 ( 
.A1(n_748),
.A2(n_561),
.B(n_560),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_L g900 ( 
.A(n_658),
.B(n_605),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_669),
.B(n_605),
.Y(n_901)
);

INVx11_ASAP7_75t_L g902 ( 
.A(n_808),
.Y(n_902)
);

BUFx6f_ASAP7_75t_L g903 ( 
.A(n_703),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_792),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_793),
.Y(n_905)
);

NOR3xp33_ASAP7_75t_L g906 ( 
.A(n_762),
.B(n_312),
.C(n_301),
.Y(n_906)
);

AOI21xp5_ASAP7_75t_L g907 ( 
.A1(n_748),
.A2(n_582),
.B(n_573),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_662),
.Y(n_908)
);

AND2x4_ASAP7_75t_L g909 ( 
.A(n_758),
.B(n_495),
.Y(n_909)
);

AOI21xp5_ASAP7_75t_L g910 ( 
.A1(n_756),
.A2(n_589),
.B(n_582),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_L g911 ( 
.A(n_739),
.B(n_495),
.Y(n_911)
);

OAI21xp5_ASAP7_75t_L g912 ( 
.A1(n_747),
.A2(n_591),
.B(n_589),
.Y(n_912)
);

INVx2_ASAP7_75t_L g913 ( 
.A(n_664),
.Y(n_913)
);

AOI21xp5_ASAP7_75t_L g914 ( 
.A1(n_756),
.A2(n_592),
.B(n_593),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_L g915 ( 
.A(n_754),
.B(n_764),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_L g916 ( 
.A(n_764),
.B(n_495),
.Y(n_916)
);

OAI22xp5_ASAP7_75t_L g917 ( 
.A1(n_710),
.A2(n_502),
.B1(n_505),
.B2(n_594),
.Y(n_917)
);

AOI21x1_ASAP7_75t_L g918 ( 
.A1(n_798),
.A2(n_604),
.B(n_592),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_L g919 ( 
.A(n_764),
.B(n_502),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_L g920 ( 
.A(n_667),
.B(n_502),
.Y(n_920)
);

OAI21xp5_ASAP7_75t_L g921 ( 
.A1(n_759),
.A2(n_604),
.B(n_593),
.Y(n_921)
);

INVx1_ASAP7_75t_SL g922 ( 
.A(n_695),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_L g923 ( 
.A(n_667),
.B(n_505),
.Y(n_923)
);

O2A1O1Ixp33_ASAP7_75t_L g924 ( 
.A1(n_766),
.A2(n_601),
.B(n_594),
.C(n_505),
.Y(n_924)
);

BUFx6f_ASAP7_75t_L g925 ( 
.A(n_710),
.Y(n_925)
);

BUFx6f_ASAP7_75t_L g926 ( 
.A(n_711),
.Y(n_926)
);

NOR2xp33_ASAP7_75t_L g927 ( 
.A(n_663),
.B(n_594),
.Y(n_927)
);

AOI21xp5_ASAP7_75t_L g928 ( 
.A1(n_723),
.A2(n_601),
.B(n_613),
.Y(n_928)
);

AOI21xp5_ASAP7_75t_L g929 ( 
.A1(n_725),
.A2(n_601),
.B(n_613),
.Y(n_929)
);

AOI21xp5_ASAP7_75t_L g930 ( 
.A1(n_728),
.A2(n_575),
.B(n_613),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_L g931 ( 
.A(n_771),
.B(n_539),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_L g932 ( 
.A(n_774),
.B(n_539),
.Y(n_932)
);

INVx1_ASAP7_75t_L g933 ( 
.A(n_683),
.Y(n_933)
);

AOI21xp5_ASAP7_75t_L g934 ( 
.A1(n_661),
.A2(n_575),
.B(n_613),
.Y(n_934)
);

NOR2xp33_ASAP7_75t_L g935 ( 
.A(n_665),
.B(n_539),
.Y(n_935)
);

AO21x1_ASAP7_75t_L g936 ( 
.A1(n_705),
.A2(n_549),
.B(n_565),
.Y(n_936)
);

INVx3_ASAP7_75t_L g937 ( 
.A(n_711),
.Y(n_937)
);

BUFx6f_ASAP7_75t_L g938 ( 
.A(n_810),
.Y(n_938)
);

A2O1A1Ixp33_ASAP7_75t_L g939 ( 
.A1(n_814),
.A2(n_435),
.B(n_316),
.C(n_326),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_L g940 ( 
.A(n_775),
.B(n_539),
.Y(n_940)
);

AOI21xp5_ASAP7_75t_L g941 ( 
.A1(n_684),
.A2(n_706),
.B(n_670),
.Y(n_941)
);

AND2x2_ASAP7_75t_L g942 ( 
.A(n_695),
.B(n_315),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_L g943 ( 
.A(n_668),
.B(n_539),
.Y(n_943)
);

AOI21xp5_ASAP7_75t_L g944 ( 
.A1(n_660),
.A2(n_575),
.B(n_613),
.Y(n_944)
);

O2A1O1Ixp33_ASAP7_75t_L g945 ( 
.A1(n_693),
.A2(n_435),
.B(n_437),
.C(n_432),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_SL g946 ( 
.A(n_722),
.B(n_575),
.Y(n_946)
);

O2A1O1Ixp5_ASAP7_75t_L g947 ( 
.A1(n_812),
.A2(n_437),
.B(n_432),
.C(n_428),
.Y(n_947)
);

AOI21xp5_ASAP7_75t_L g948 ( 
.A1(n_705),
.A2(n_579),
.B(n_575),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_SL g949 ( 
.A(n_722),
.B(n_733),
.Y(n_949)
);

AOI21xp5_ASAP7_75t_L g950 ( 
.A1(n_813),
.A2(n_579),
.B(n_527),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_683),
.Y(n_951)
);

AOI33xp33_ASAP7_75t_L g952 ( 
.A1(n_799),
.A2(n_318),
.A3(n_323),
.B1(n_324),
.B2(n_333),
.B3(n_10),
.Y(n_952)
);

A2O1A1Ixp33_ASAP7_75t_L g953 ( 
.A1(n_650),
.A2(n_709),
.B(n_724),
.C(n_726),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_L g954 ( 
.A(n_687),
.B(n_579),
.Y(n_954)
);

AOI21xp5_ASAP7_75t_L g955 ( 
.A1(n_809),
.A2(n_579),
.B(n_527),
.Y(n_955)
);

O2A1O1Ixp5_ASAP7_75t_L g956 ( 
.A1(n_812),
.A2(n_437),
.B(n_432),
.C(n_428),
.Y(n_956)
);

OAI21xp5_ASAP7_75t_L g957 ( 
.A1(n_685),
.A2(n_552),
.B(n_571),
.Y(n_957)
);

BUFx3_ASAP7_75t_L g958 ( 
.A(n_729),
.Y(n_958)
);

OAI21xp5_ASAP7_75t_L g959 ( 
.A1(n_685),
.A2(n_552),
.B(n_571),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_L g960 ( 
.A(n_737),
.B(n_579),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_L g961 ( 
.A(n_738),
.B(n_577),
.Y(n_961)
);

OAI22xp5_ASAP7_75t_L g962 ( 
.A1(n_742),
.A2(n_528),
.B1(n_527),
.B2(n_320),
.Y(n_962)
);

NOR3xp33_ASAP7_75t_L g963 ( 
.A(n_781),
.B(n_290),
.C(n_287),
.Y(n_963)
);

INVx2_ASAP7_75t_L g964 ( 
.A(n_691),
.Y(n_964)
);

AOI21xp5_ASAP7_75t_L g965 ( 
.A1(n_809),
.A2(n_527),
.B(n_528),
.Y(n_965)
);

AOI21x1_ASAP7_75t_L g966 ( 
.A1(n_798),
.A2(n_428),
.B(n_528),
.Y(n_966)
);

NOR2xp33_ASAP7_75t_L g967 ( 
.A(n_727),
.B(n_4),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_L g968 ( 
.A(n_790),
.B(n_761),
.Y(n_968)
);

AOI33xp33_ASAP7_75t_L g969 ( 
.A1(n_790),
.A2(n_5),
.A3(n_7),
.B1(n_9),
.B2(n_12),
.B3(n_14),
.Y(n_969)
);

AOI21xp5_ASAP7_75t_L g970 ( 
.A1(n_801),
.A2(n_527),
.B(n_528),
.Y(n_970)
);

AOI21xp5_ASAP7_75t_L g971 ( 
.A1(n_699),
.A2(n_527),
.B(n_528),
.Y(n_971)
);

INVx2_ASAP7_75t_L g972 ( 
.A(n_699),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_L g973 ( 
.A(n_790),
.B(n_577),
.Y(n_973)
);

AOI21xp5_ASAP7_75t_L g974 ( 
.A1(n_709),
.A2(n_724),
.B(n_717),
.Y(n_974)
);

AOI21xp5_ASAP7_75t_L g975 ( 
.A1(n_717),
.A2(n_528),
.B(n_172),
.Y(n_975)
);

AOI21xp5_ASAP7_75t_L g976 ( 
.A1(n_726),
.A2(n_269),
.B(n_179),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_L g977 ( 
.A(n_786),
.B(n_577),
.Y(n_977)
);

AOI21xp5_ASAP7_75t_L g978 ( 
.A1(n_740),
.A2(n_276),
.B(n_184),
.Y(n_978)
);

NOR3xp33_ASAP7_75t_L g979 ( 
.A(n_781),
.B(n_264),
.C(n_281),
.Y(n_979)
);

AOI21x1_ASAP7_75t_L g980 ( 
.A1(n_803),
.A2(n_621),
.B(n_529),
.Y(n_980)
);

OAI21xp5_ASAP7_75t_L g981 ( 
.A1(n_740),
.A2(n_571),
.B(n_567),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_SL g982 ( 
.A(n_733),
.B(n_424),
.Y(n_982)
);

HB1xp67_ASAP7_75t_L g983 ( 
.A(n_729),
.Y(n_983)
);

AOI21xp5_ASAP7_75t_L g984 ( 
.A1(n_755),
.A2(n_791),
.B(n_785),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_L g985 ( 
.A(n_777),
.B(n_577),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_L g986 ( 
.A(n_783),
.B(n_784),
.Y(n_986)
);

CKINVDCx5p33_ASAP7_75t_R g987 ( 
.A(n_800),
.Y(n_987)
);

AOI22xp33_ASAP7_75t_L g988 ( 
.A1(n_755),
.A2(n_577),
.B1(n_552),
.B2(n_571),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_L g989 ( 
.A(n_697),
.B(n_577),
.Y(n_989)
);

OAI21xp33_ASAP7_75t_L g990 ( 
.A1(n_797),
.A2(n_292),
.B(n_334),
.Y(n_990)
);

AOI21xp5_ASAP7_75t_L g991 ( 
.A1(n_769),
.A2(n_785),
.B(n_791),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_L g992 ( 
.A(n_758),
.B(n_757),
.Y(n_992)
);

AOI21xp5_ASAP7_75t_L g993 ( 
.A1(n_769),
.A2(n_178),
.B(n_189),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_L g994 ( 
.A(n_757),
.B(n_529),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_778),
.Y(n_995)
);

A2O1A1Ixp33_ASAP7_75t_L g996 ( 
.A1(n_778),
.A2(n_749),
.B(n_746),
.C(n_734),
.Y(n_996)
);

AOI21xp5_ASAP7_75t_L g997 ( 
.A1(n_749),
.A2(n_293),
.B(n_193),
.Y(n_997)
);

INVx1_ASAP7_75t_L g998 ( 
.A(n_802),
.Y(n_998)
);

BUFx3_ASAP7_75t_L g999 ( 
.A(n_729),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_L g1000 ( 
.A(n_720),
.B(n_529),
.Y(n_1000)
);

AOI21xp5_ASAP7_75t_L g1001 ( 
.A1(n_746),
.A2(n_296),
.B(n_196),
.Y(n_1001)
);

OAI22xp5_ASAP7_75t_L g1002 ( 
.A1(n_751),
.A2(n_254),
.B1(n_253),
.B2(n_246),
.Y(n_1002)
);

AOI21xp5_ASAP7_75t_L g1003 ( 
.A1(n_807),
.A2(n_192),
.B(n_199),
.Y(n_1003)
);

AOI21xp5_ASAP7_75t_L g1004 ( 
.A1(n_803),
.A2(n_319),
.B(n_208),
.Y(n_1004)
);

O2A1O1Ixp33_ASAP7_75t_L g1005 ( 
.A1(n_736),
.A2(n_529),
.B(n_552),
.C(n_567),
.Y(n_1005)
);

O2A1O1Ixp33_ASAP7_75t_L g1006 ( 
.A1(n_854),
.A2(n_789),
.B(n_795),
.C(n_796),
.Y(n_1006)
);

CKINVDCx5p33_ASAP7_75t_R g1007 ( 
.A(n_829),
.Y(n_1007)
);

BUFx4f_ASAP7_75t_SL g1008 ( 
.A(n_832),
.Y(n_1008)
);

AND2x2_ASAP7_75t_L g1009 ( 
.A(n_884),
.B(n_743),
.Y(n_1009)
);

INVx3_ASAP7_75t_L g1010 ( 
.A(n_825),
.Y(n_1010)
);

A2O1A1Ixp33_ASAP7_75t_L g1011 ( 
.A1(n_996),
.A2(n_794),
.B(n_719),
.C(n_782),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_SL g1012 ( 
.A(n_835),
.B(n_751),
.Y(n_1012)
);

AOI22xp5_ASAP7_75t_L g1013 ( 
.A1(n_987),
.A2(n_666),
.B1(n_731),
.B2(n_811),
.Y(n_1013)
);

OAI21xp5_ASAP7_75t_L g1014 ( 
.A1(n_882),
.A2(n_696),
.B(n_805),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_823),
.Y(n_1015)
);

INVx1_ASAP7_75t_L g1016 ( 
.A(n_850),
.Y(n_1016)
);

AOI21xp5_ASAP7_75t_L g1017 ( 
.A1(n_870),
.A2(n_810),
.B(n_815),
.Y(n_1017)
);

CKINVDCx5p33_ASAP7_75t_R g1018 ( 
.A(n_889),
.Y(n_1018)
);

INVx3_ASAP7_75t_L g1019 ( 
.A(n_825),
.Y(n_1019)
);

INVx1_ASAP7_75t_L g1020 ( 
.A(n_881),
.Y(n_1020)
);

INVx1_ASAP7_75t_L g1021 ( 
.A(n_892),
.Y(n_1021)
);

A2O1A1Ixp33_ASAP7_75t_L g1022 ( 
.A1(n_996),
.A2(n_782),
.B(n_751),
.C(n_810),
.Y(n_1022)
);

OAI211xp5_ASAP7_75t_SL g1023 ( 
.A1(n_952),
.A2(n_767),
.B(n_806),
.C(n_804),
.Y(n_1023)
);

AOI21xp5_ASAP7_75t_L g1024 ( 
.A1(n_885),
.A2(n_815),
.B(n_806),
.Y(n_1024)
);

NAND2xp5_ASAP7_75t_SL g1025 ( 
.A(n_835),
.B(n_782),
.Y(n_1025)
);

INVx3_ASAP7_75t_L g1026 ( 
.A(n_835),
.Y(n_1026)
);

O2A1O1Ixp33_ASAP7_75t_L g1027 ( 
.A1(n_841),
.A2(n_804),
.B(n_735),
.C(n_811),
.Y(n_1027)
);

OAI21xp33_ASAP7_75t_SL g1028 ( 
.A1(n_862),
.A2(n_969),
.B(n_986),
.Y(n_1028)
);

AND2x4_ASAP7_75t_L g1029 ( 
.A(n_958),
.B(n_770),
.Y(n_1029)
);

NOR2xp33_ASAP7_75t_L g1030 ( 
.A(n_817),
.B(n_735),
.Y(n_1030)
);

AOI21xp5_ASAP7_75t_L g1031 ( 
.A1(n_948),
.A2(n_424),
.B(n_263),
.Y(n_1031)
);

AOI21xp5_ASAP7_75t_L g1032 ( 
.A1(n_847),
.A2(n_424),
.B(n_317),
.Y(n_1032)
);

BUFx3_ASAP7_75t_L g1033 ( 
.A(n_958),
.Y(n_1033)
);

INVx1_ASAP7_75t_SL g1034 ( 
.A(n_922),
.Y(n_1034)
);

HB1xp67_ASAP7_75t_L g1035 ( 
.A(n_833),
.Y(n_1035)
);

HB1xp67_ASAP7_75t_L g1036 ( 
.A(n_915),
.Y(n_1036)
);

AOI21xp5_ASAP7_75t_L g1037 ( 
.A1(n_941),
.A2(n_424),
.B(n_317),
.Y(n_1037)
);

INVx3_ASAP7_75t_L g1038 ( 
.A(n_835),
.Y(n_1038)
);

NOR2xp33_ASAP7_75t_L g1039 ( 
.A(n_816),
.B(n_666),
.Y(n_1039)
);

INVx1_ASAP7_75t_L g1040 ( 
.A(n_904),
.Y(n_1040)
);

NAND3xp33_ASAP7_75t_L g1041 ( 
.A(n_821),
.B(n_808),
.C(n_330),
.Y(n_1041)
);

INVxp67_ASAP7_75t_L g1042 ( 
.A(n_967),
.Y(n_1042)
);

INVx1_ASAP7_75t_L g1043 ( 
.A(n_905),
.Y(n_1043)
);

AO32x2_ASAP7_75t_L g1044 ( 
.A1(n_871),
.A2(n_917),
.A3(n_962),
.B1(n_839),
.B2(n_936),
.Y(n_1044)
);

BUFx6f_ASAP7_75t_L g1045 ( 
.A(n_999),
.Y(n_1045)
);

INVx2_ASAP7_75t_SL g1046 ( 
.A(n_902),
.Y(n_1046)
);

NAND2x1p5_ASAP7_75t_L g1047 ( 
.A(n_999),
.B(n_808),
.Y(n_1047)
);

OA22x2_ASAP7_75t_L g1048 ( 
.A1(n_942),
.A2(n_731),
.B1(n_780),
.B2(n_529),
.Y(n_1048)
);

INVxp67_ASAP7_75t_L g1049 ( 
.A(n_967),
.Y(n_1049)
);

INVx2_ASAP7_75t_L g1050 ( 
.A(n_837),
.Y(n_1050)
);

INVx2_ASAP7_75t_L g1051 ( 
.A(n_851),
.Y(n_1051)
);

NAND2xp5_ASAP7_75t_L g1052 ( 
.A(n_998),
.B(n_780),
.Y(n_1052)
);

NAND2xp5_ASAP7_75t_L g1053 ( 
.A(n_968),
.B(n_770),
.Y(n_1053)
);

NAND2xp5_ASAP7_75t_L g1054 ( 
.A(n_862),
.B(n_864),
.Y(n_1054)
);

CKINVDCx5p33_ASAP7_75t_R g1055 ( 
.A(n_873),
.Y(n_1055)
);

NAND2xp5_ASAP7_75t_SL g1056 ( 
.A(n_859),
.B(n_869),
.Y(n_1056)
);

CKINVDCx11_ASAP7_75t_R g1057 ( 
.A(n_859),
.Y(n_1057)
);

OA22x2_ASAP7_75t_L g1058 ( 
.A1(n_853),
.A2(n_842),
.B1(n_855),
.B2(n_836),
.Y(n_1058)
);

OAI22x1_ASAP7_75t_SL g1059 ( 
.A1(n_969),
.A2(n_227),
.B1(n_228),
.B2(n_207),
.Y(n_1059)
);

INVx2_ASAP7_75t_L g1060 ( 
.A(n_858),
.Y(n_1060)
);

OAI21x1_ASAP7_75t_L g1061 ( 
.A1(n_844),
.A2(n_770),
.B(n_552),
.Y(n_1061)
);

NOR2xp33_ASAP7_75t_R g1062 ( 
.A(n_876),
.B(n_869),
.Y(n_1062)
);

AOI21xp5_ASAP7_75t_L g1063 ( 
.A1(n_949),
.A2(n_424),
.B(n_317),
.Y(n_1063)
);

NAND2xp5_ASAP7_75t_SL g1064 ( 
.A(n_859),
.B(n_328),
.Y(n_1064)
);

BUFx6f_ASAP7_75t_L g1065 ( 
.A(n_859),
.Y(n_1065)
);

INVx1_ASAP7_75t_L g1066 ( 
.A(n_908),
.Y(n_1066)
);

OAI21x1_ASAP7_75t_L g1067 ( 
.A1(n_867),
.A2(n_966),
.B(n_899),
.Y(n_1067)
);

NAND2xp5_ASAP7_75t_L g1068 ( 
.A(n_864),
.B(n_843),
.Y(n_1068)
);

OAI21xp33_ASAP7_75t_SL g1069 ( 
.A1(n_977),
.A2(n_12),
.B(n_16),
.Y(n_1069)
);

AOI22xp5_ASAP7_75t_L g1070 ( 
.A1(n_895),
.A2(n_770),
.B1(n_571),
.B2(n_567),
.Y(n_1070)
);

NAND2xp5_ASAP7_75t_L g1071 ( 
.A(n_842),
.B(n_770),
.Y(n_1071)
);

NOR2xp67_ASAP7_75t_SL g1072 ( 
.A(n_848),
.B(n_856),
.Y(n_1072)
);

NAND2xp5_ASAP7_75t_SL g1073 ( 
.A(n_856),
.B(n_327),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_L g1074 ( 
.A(n_911),
.B(n_571),
.Y(n_1074)
);

NAND2xp5_ASAP7_75t_SL g1075 ( 
.A(n_848),
.B(n_332),
.Y(n_1075)
);

INVx3_ASAP7_75t_L g1076 ( 
.A(n_938),
.Y(n_1076)
);

NAND2xp5_ASAP7_75t_L g1077 ( 
.A(n_821),
.B(n_571),
.Y(n_1077)
);

AOI21xp5_ASAP7_75t_L g1078 ( 
.A1(n_949),
.A2(n_424),
.B(n_317),
.Y(n_1078)
);

INVx2_ASAP7_75t_L g1079 ( 
.A(n_913),
.Y(n_1079)
);

OAI22xp5_ASAP7_75t_L g1080 ( 
.A1(n_888),
.A2(n_303),
.B1(n_256),
.B2(n_241),
.Y(n_1080)
);

INVx1_ASAP7_75t_L g1081 ( 
.A(n_933),
.Y(n_1081)
);

NOR2xp33_ASAP7_75t_L g1082 ( 
.A(n_861),
.B(n_234),
.Y(n_1082)
);

AOI21xp5_ASAP7_75t_L g1083 ( 
.A1(n_827),
.A2(n_828),
.B(n_931),
.Y(n_1083)
);

NOR2xp33_ASAP7_75t_L g1084 ( 
.A(n_826),
.B(n_17),
.Y(n_1084)
);

AOI21xp5_ASAP7_75t_L g1085 ( 
.A1(n_866),
.A2(n_317),
.B(n_567),
.Y(n_1085)
);

HB1xp67_ASAP7_75t_L g1086 ( 
.A(n_973),
.Y(n_1086)
);

AOI21xp5_ASAP7_75t_L g1087 ( 
.A1(n_932),
.A2(n_317),
.B(n_567),
.Y(n_1087)
);

BUFx6f_ASAP7_75t_L g1088 ( 
.A(n_938),
.Y(n_1088)
);

INVx1_ASAP7_75t_L g1089 ( 
.A(n_951),
.Y(n_1089)
);

CKINVDCx5p33_ASAP7_75t_R g1090 ( 
.A(n_983),
.Y(n_1090)
);

INVx1_ASAP7_75t_L g1091 ( 
.A(n_995),
.Y(n_1091)
);

INVx1_ASAP7_75t_L g1092 ( 
.A(n_834),
.Y(n_1092)
);

INVxp67_ASAP7_75t_L g1093 ( 
.A(n_818),
.Y(n_1093)
);

A2O1A1Ixp33_ASAP7_75t_L g1094 ( 
.A1(n_839),
.A2(n_567),
.B(n_552),
.C(n_621),
.Y(n_1094)
);

INVx2_ASAP7_75t_L g1095 ( 
.A(n_964),
.Y(n_1095)
);

AOI21xp5_ASAP7_75t_L g1096 ( 
.A1(n_940),
.A2(n_567),
.B(n_552),
.Y(n_1096)
);

NOR2xp33_ASAP7_75t_R g1097 ( 
.A(n_938),
.B(n_621),
.Y(n_1097)
);

O2A1O1Ixp33_ASAP7_75t_SL g1098 ( 
.A1(n_838),
.A2(n_18),
.B(n_20),
.C(n_21),
.Y(n_1098)
);

AOI33xp33_ASAP7_75t_L g1099 ( 
.A1(n_952),
.A2(n_20),
.A3(n_24),
.B1(n_27),
.B2(n_29),
.B3(n_30),
.Y(n_1099)
);

BUFx3_ASAP7_75t_L g1100 ( 
.A(n_983),
.Y(n_1100)
);

NOR2xp33_ASAP7_75t_L g1101 ( 
.A(n_992),
.B(n_24),
.Y(n_1101)
);

AOI21xp5_ASAP7_75t_L g1102 ( 
.A1(n_819),
.A2(n_621),
.B(n_426),
.Y(n_1102)
);

INVx2_ASAP7_75t_L g1103 ( 
.A(n_972),
.Y(n_1103)
);

O2A1O1Ixp33_ASAP7_75t_L g1104 ( 
.A1(n_882),
.A2(n_32),
.B(n_33),
.C(n_34),
.Y(n_1104)
);

O2A1O1Ixp33_ASAP7_75t_L g1105 ( 
.A1(n_896),
.A2(n_34),
.B(n_35),
.C(n_37),
.Y(n_1105)
);

AOI21xp5_ASAP7_75t_L g1106 ( 
.A1(n_930),
.A2(n_621),
.B(n_125),
.Y(n_1106)
);

NAND2xp5_ASAP7_75t_SL g1107 ( 
.A(n_903),
.B(n_621),
.Y(n_1107)
);

NAND2xp5_ASAP7_75t_L g1108 ( 
.A(n_849),
.B(n_621),
.Y(n_1108)
);

AOI22xp5_ASAP7_75t_L g1109 ( 
.A1(n_895),
.A2(n_426),
.B1(n_37),
.B2(n_39),
.Y(n_1109)
);

INVxp67_ASAP7_75t_SL g1110 ( 
.A(n_890),
.Y(n_1110)
);

INVx6_ASAP7_75t_L g1111 ( 
.A(n_909),
.Y(n_1111)
);

AOI21xp5_ASAP7_75t_L g1112 ( 
.A1(n_877),
.A2(n_108),
.B(n_163),
.Y(n_1112)
);

INVx2_ASAP7_75t_L g1113 ( 
.A(n_830),
.Y(n_1113)
);

OAI21xp5_ASAP7_75t_L g1114 ( 
.A1(n_852),
.A2(n_426),
.B(n_39),
.Y(n_1114)
);

AOI22xp5_ASAP7_75t_L g1115 ( 
.A1(n_963),
.A2(n_979),
.B1(n_990),
.B2(n_906),
.Y(n_1115)
);

NOR2xp33_ASAP7_75t_L g1116 ( 
.A(n_900),
.B(n_35),
.Y(n_1116)
);

INVx1_ASAP7_75t_L g1117 ( 
.A(n_927),
.Y(n_1117)
);

NOR2xp33_ASAP7_75t_R g1118 ( 
.A(n_938),
.B(n_158),
.Y(n_1118)
);

AOI21xp5_ASAP7_75t_L g1119 ( 
.A1(n_865),
.A2(n_426),
.B(n_42),
.Y(n_1119)
);

O2A1O1Ixp33_ASAP7_75t_L g1120 ( 
.A1(n_896),
.A2(n_41),
.B(n_43),
.C(n_44),
.Y(n_1120)
);

AOI21xp5_ASAP7_75t_L g1121 ( 
.A1(n_887),
.A2(n_426),
.B(n_46),
.Y(n_1121)
);

NAND2xp5_ASAP7_75t_L g1122 ( 
.A(n_863),
.B(n_41),
.Y(n_1122)
);

AOI21xp5_ASAP7_75t_L g1123 ( 
.A1(n_912),
.A2(n_47),
.B(n_48),
.Y(n_1123)
);

OR2x4_ASAP7_75t_L g1124 ( 
.A(n_903),
.B(n_48),
.Y(n_1124)
);

INVx1_ASAP7_75t_L g1125 ( 
.A(n_927),
.Y(n_1125)
);

OR2x2_ASAP7_75t_L g1126 ( 
.A(n_1002),
.B(n_54),
.Y(n_1126)
);

AOI21xp5_ASAP7_75t_L g1127 ( 
.A1(n_921),
.A2(n_56),
.B(n_57),
.Y(n_1127)
);

OAI22xp5_ASAP7_75t_L g1128 ( 
.A1(n_840),
.A2(n_57),
.B1(n_60),
.B2(n_61),
.Y(n_1128)
);

O2A1O1Ixp33_ASAP7_75t_L g1129 ( 
.A1(n_820),
.A2(n_939),
.B(n_985),
.C(n_920),
.Y(n_1129)
);

NAND2xp5_ASAP7_75t_L g1130 ( 
.A(n_909),
.B(n_60),
.Y(n_1130)
);

INVx1_ASAP7_75t_L g1131 ( 
.A(n_916),
.Y(n_1131)
);

NAND2xp5_ASAP7_75t_L g1132 ( 
.A(n_919),
.B(n_61),
.Y(n_1132)
);

AO31x2_ASAP7_75t_L g1133 ( 
.A1(n_953),
.A2(n_89),
.A3(n_138),
.B(n_127),
.Y(n_1133)
);

INVx1_ASAP7_75t_L g1134 ( 
.A(n_961),
.Y(n_1134)
);

INVx1_ASAP7_75t_L g1135 ( 
.A(n_943),
.Y(n_1135)
);

AOI21xp5_ASAP7_75t_L g1136 ( 
.A1(n_928),
.A2(n_62),
.B(n_64),
.Y(n_1136)
);

NOR2xp67_ASAP7_75t_L g1137 ( 
.A(n_857),
.B(n_85),
.Y(n_1137)
);

INVx1_ASAP7_75t_SL g1138 ( 
.A(n_994),
.Y(n_1138)
);

AOI21xp5_ASAP7_75t_L g1139 ( 
.A1(n_929),
.A2(n_64),
.B(n_65),
.Y(n_1139)
);

BUFx4f_ASAP7_75t_SL g1140 ( 
.A(n_903),
.Y(n_1140)
);

NOR3xp33_ASAP7_75t_SL g1141 ( 
.A(n_939),
.B(n_65),
.C(n_67),
.Y(n_1141)
);

AOI21xp5_ASAP7_75t_L g1142 ( 
.A1(n_878),
.A2(n_69),
.B(n_70),
.Y(n_1142)
);

CKINVDCx20_ASAP7_75t_R g1143 ( 
.A(n_903),
.Y(n_1143)
);

AOI21xp5_ASAP7_75t_L g1144 ( 
.A1(n_923),
.A2(n_94),
.B(n_98),
.Y(n_1144)
);

OAI22x1_ASAP7_75t_L g1145 ( 
.A1(n_879),
.A2(n_105),
.B1(n_126),
.B2(n_156),
.Y(n_1145)
);

OAI22xp5_ASAP7_75t_L g1146 ( 
.A1(n_840),
.A2(n_901),
.B1(n_898),
.B2(n_937),
.Y(n_1146)
);

OAI22xp5_ASAP7_75t_L g1147 ( 
.A1(n_898),
.A2(n_937),
.B1(n_894),
.B2(n_925),
.Y(n_1147)
);

NOR2xp33_ASAP7_75t_L g1148 ( 
.A(n_860),
.B(n_954),
.Y(n_1148)
);

INVx1_ASAP7_75t_L g1149 ( 
.A(n_960),
.Y(n_1149)
);

AND2x2_ASAP7_75t_L g1150 ( 
.A(n_997),
.B(n_988),
.Y(n_1150)
);

NAND2xp5_ASAP7_75t_SL g1151 ( 
.A(n_925),
.B(n_926),
.Y(n_1151)
);

INVx2_ASAP7_75t_SL g1152 ( 
.A(n_925),
.Y(n_1152)
);

INVx3_ASAP7_75t_L g1153 ( 
.A(n_925),
.Y(n_1153)
);

AOI21xp5_ASAP7_75t_L g1154 ( 
.A1(n_924),
.A2(n_875),
.B(n_874),
.Y(n_1154)
);

AOI21xp5_ASAP7_75t_L g1155 ( 
.A1(n_824),
.A2(n_845),
.B(n_831),
.Y(n_1155)
);

NOR2xp67_ASAP7_75t_L g1156 ( 
.A(n_935),
.B(n_1001),
.Y(n_1156)
);

O2A1O1Ixp33_ASAP7_75t_L g1157 ( 
.A1(n_868),
.A2(n_872),
.B(n_880),
.C(n_1005),
.Y(n_1157)
);

AND2x4_ASAP7_75t_L g1158 ( 
.A(n_926),
.B(n_838),
.Y(n_1158)
);

NAND2xp5_ASAP7_75t_SL g1159 ( 
.A(n_926),
.B(n_894),
.Y(n_1159)
);

NAND3xp33_ASAP7_75t_L g1160 ( 
.A(n_1003),
.B(n_953),
.C(n_993),
.Y(n_1160)
);

OAI22xp5_ASAP7_75t_L g1161 ( 
.A1(n_1054),
.A2(n_926),
.B1(n_935),
.B2(n_988),
.Y(n_1161)
);

INVx1_ASAP7_75t_L g1162 ( 
.A(n_1015),
.Y(n_1162)
);

OAI21x1_ASAP7_75t_L g1163 ( 
.A1(n_1067),
.A2(n_918),
.B(n_956),
.Y(n_1163)
);

AOI21xp5_ASAP7_75t_L g1164 ( 
.A1(n_1083),
.A2(n_944),
.B(n_934),
.Y(n_1164)
);

BUFx2_ASAP7_75t_L g1165 ( 
.A(n_1008),
.Y(n_1165)
);

AND2x2_ASAP7_75t_L g1166 ( 
.A(n_1009),
.B(n_957),
.Y(n_1166)
);

INVx3_ASAP7_75t_L g1167 ( 
.A(n_1088),
.Y(n_1167)
);

AO31x2_ASAP7_75t_L g1168 ( 
.A1(n_1083),
.A2(n_1096),
.A3(n_1154),
.B(n_1031),
.Y(n_1168)
);

NAND2xp5_ASAP7_75t_L g1169 ( 
.A(n_1036),
.B(n_974),
.Y(n_1169)
);

INVx1_ASAP7_75t_L g1170 ( 
.A(n_1016),
.Y(n_1170)
);

AOI21xp5_ASAP7_75t_L g1171 ( 
.A1(n_1154),
.A2(n_846),
.B(n_946),
.Y(n_1171)
);

OAI21x1_ASAP7_75t_L g1172 ( 
.A1(n_1155),
.A2(n_947),
.B(n_991),
.Y(n_1172)
);

INVx3_ASAP7_75t_L g1173 ( 
.A(n_1088),
.Y(n_1173)
);

INVx1_ASAP7_75t_L g1174 ( 
.A(n_1020),
.Y(n_1174)
);

OR2x2_ASAP7_75t_L g1175 ( 
.A(n_1030),
.B(n_1035),
.Y(n_1175)
);

OR2x2_ASAP7_75t_L g1176 ( 
.A(n_1042),
.B(n_1000),
.Y(n_1176)
);

AO31x2_ASAP7_75t_L g1177 ( 
.A1(n_1096),
.A2(n_822),
.A3(n_984),
.B(n_989),
.Y(n_1177)
);

AOI21xp5_ASAP7_75t_L g1178 ( 
.A1(n_1155),
.A2(n_846),
.B(n_946),
.Y(n_1178)
);

AND2x4_ASAP7_75t_L g1179 ( 
.A(n_1143),
.B(n_981),
.Y(n_1179)
);

CKINVDCx5p33_ASAP7_75t_R g1180 ( 
.A(n_1018),
.Y(n_1180)
);

OAI22xp5_ASAP7_75t_L g1181 ( 
.A1(n_1049),
.A2(n_868),
.B1(n_872),
.B2(n_880),
.Y(n_1181)
);

AOI221xp5_ASAP7_75t_SL g1182 ( 
.A1(n_1123),
.A2(n_976),
.B1(n_978),
.B2(n_891),
.C(n_893),
.Y(n_1182)
);

AOI21xp5_ASAP7_75t_L g1183 ( 
.A1(n_1037),
.A2(n_982),
.B(n_965),
.Y(n_1183)
);

OR2x2_ASAP7_75t_L g1184 ( 
.A(n_1034),
.B(n_959),
.Y(n_1184)
);

A2O1A1Ixp33_ASAP7_75t_L g1185 ( 
.A1(n_1084),
.A2(n_975),
.B(n_982),
.C(n_955),
.Y(n_1185)
);

OAI21x1_ASAP7_75t_L g1186 ( 
.A1(n_1032),
.A2(n_1037),
.B(n_1031),
.Y(n_1186)
);

AO31x2_ASAP7_75t_L g1187 ( 
.A1(n_1063),
.A2(n_971),
.A3(n_886),
.B(n_897),
.Y(n_1187)
);

AOI21xp5_ASAP7_75t_L g1188 ( 
.A1(n_1017),
.A2(n_950),
.B(n_907),
.Y(n_1188)
);

AOI21xp5_ASAP7_75t_L g1189 ( 
.A1(n_1017),
.A2(n_1146),
.B(n_1114),
.Y(n_1189)
);

AOI21xp5_ASAP7_75t_L g1190 ( 
.A1(n_1129),
.A2(n_883),
.B(n_910),
.Y(n_1190)
);

CKINVDCx20_ASAP7_75t_R g1191 ( 
.A(n_1007),
.Y(n_1191)
);

BUFx2_ASAP7_75t_L g1192 ( 
.A(n_1090),
.Y(n_1192)
);

AO31x2_ASAP7_75t_L g1193 ( 
.A1(n_1063),
.A2(n_914),
.A3(n_970),
.B(n_1004),
.Y(n_1193)
);

NAND2xp5_ASAP7_75t_L g1194 ( 
.A(n_1052),
.B(n_945),
.Y(n_1194)
);

INVx1_ASAP7_75t_SL g1195 ( 
.A(n_1055),
.Y(n_1195)
);

NAND2xp5_ASAP7_75t_L g1196 ( 
.A(n_1039),
.B(n_980),
.Y(n_1196)
);

O2A1O1Ixp33_ASAP7_75t_L g1197 ( 
.A1(n_1126),
.A2(n_1028),
.B(n_1120),
.C(n_1105),
.Y(n_1197)
);

AOI222xp33_ASAP7_75t_L g1198 ( 
.A1(n_1059),
.A2(n_1082),
.B1(n_1040),
.B2(n_1021),
.C1(n_1043),
.C2(n_1092),
.Y(n_1198)
);

O2A1O1Ixp5_ASAP7_75t_L g1199 ( 
.A1(n_1123),
.A2(n_1127),
.B(n_1121),
.C(n_1119),
.Y(n_1199)
);

INVx2_ASAP7_75t_SL g1200 ( 
.A(n_1033),
.Y(n_1200)
);

AOI21xp5_ASAP7_75t_L g1201 ( 
.A1(n_1024),
.A2(n_1142),
.B(n_1068),
.Y(n_1201)
);

NOR2xp33_ASAP7_75t_L g1202 ( 
.A(n_1111),
.B(n_1124),
.Y(n_1202)
);

AOI21xp5_ASAP7_75t_L g1203 ( 
.A1(n_1024),
.A2(n_1142),
.B(n_1157),
.Y(n_1203)
);

AOI22xp5_ASAP7_75t_L g1204 ( 
.A1(n_1116),
.A2(n_1101),
.B1(n_1109),
.B2(n_1141),
.Y(n_1204)
);

AOI21xp5_ASAP7_75t_L g1205 ( 
.A1(n_1160),
.A2(n_1022),
.B(n_1032),
.Y(n_1205)
);

AO31x2_ASAP7_75t_L g1206 ( 
.A1(n_1078),
.A2(n_1087),
.A3(n_1121),
.B(n_1085),
.Y(n_1206)
);

AOI21xp5_ASAP7_75t_SL g1207 ( 
.A1(n_1110),
.A2(n_1145),
.B(n_1094),
.Y(n_1207)
);

AOI22xp5_ASAP7_75t_L g1208 ( 
.A1(n_1117),
.A2(n_1125),
.B1(n_1023),
.B2(n_1127),
.Y(n_1208)
);

INVx3_ASAP7_75t_L g1209 ( 
.A(n_1088),
.Y(n_1209)
);

AOI221xp5_ASAP7_75t_SL g1210 ( 
.A1(n_1104),
.A2(n_1128),
.B1(n_1136),
.B2(n_1139),
.C(n_1069),
.Y(n_1210)
);

OAI21xp5_ASAP7_75t_L g1211 ( 
.A1(n_1122),
.A2(n_1014),
.B(n_1119),
.Y(n_1211)
);

AOI21xp5_ASAP7_75t_L g1212 ( 
.A1(n_1147),
.A2(n_1156),
.B(n_1112),
.Y(n_1212)
);

A2O1A1Ixp33_ASAP7_75t_L g1213 ( 
.A1(n_1115),
.A2(n_1011),
.B(n_1006),
.C(n_1027),
.Y(n_1213)
);

AO32x2_ASAP7_75t_L g1214 ( 
.A1(n_1058),
.A2(n_1152),
.A3(n_1044),
.B1(n_1080),
.B2(n_1099),
.Y(n_1214)
);

A2O1A1Ixp33_ASAP7_75t_L g1215 ( 
.A1(n_1148),
.A2(n_1041),
.B(n_1150),
.C(n_1131),
.Y(n_1215)
);

INVx5_ASAP7_75t_L g1216 ( 
.A(n_1045),
.Y(n_1216)
);

AOI21xp5_ASAP7_75t_L g1217 ( 
.A1(n_1102),
.A2(n_1078),
.B(n_1144),
.Y(n_1217)
);

OAI21x1_ASAP7_75t_L g1218 ( 
.A1(n_1061),
.A2(n_1102),
.B(n_1087),
.Y(n_1218)
);

OAI21x1_ASAP7_75t_L g1219 ( 
.A1(n_1106),
.A2(n_1144),
.B(n_1139),
.Y(n_1219)
);

INVx3_ASAP7_75t_L g1220 ( 
.A(n_1065),
.Y(n_1220)
);

OAI22x1_ASAP7_75t_L g1221 ( 
.A1(n_1013),
.A2(n_1124),
.B1(n_1047),
.B2(n_1070),
.Y(n_1221)
);

OA21x2_ASAP7_75t_L g1222 ( 
.A1(n_1136),
.A2(n_1108),
.B(n_1074),
.Y(n_1222)
);

NAND2xp5_ASAP7_75t_L g1223 ( 
.A(n_1100),
.B(n_1111),
.Y(n_1223)
);

AOI22xp5_ASAP7_75t_L g1224 ( 
.A1(n_1048),
.A2(n_1077),
.B1(n_1086),
.B2(n_1132),
.Y(n_1224)
);

AOI21xp33_ASAP7_75t_L g1225 ( 
.A1(n_1058),
.A2(n_1048),
.B(n_1053),
.Y(n_1225)
);

INVx1_ASAP7_75t_L g1226 ( 
.A(n_1066),
.Y(n_1226)
);

OAI21x1_ASAP7_75t_L g1227 ( 
.A1(n_1134),
.A2(n_1107),
.B(n_1159),
.Y(n_1227)
);

O2A1O1Ixp33_ASAP7_75t_L g1228 ( 
.A1(n_1098),
.A2(n_1130),
.B(n_1073),
.C(n_1075),
.Y(n_1228)
);

OAI21xp5_ASAP7_75t_L g1229 ( 
.A1(n_1135),
.A2(n_1149),
.B(n_1064),
.Y(n_1229)
);

OAI22x1_ASAP7_75t_L g1230 ( 
.A1(n_1047),
.A2(n_1093),
.B1(n_1113),
.B2(n_1091),
.Y(n_1230)
);

AOI21xp5_ASAP7_75t_L g1231 ( 
.A1(n_1151),
.A2(n_1158),
.B(n_1056),
.Y(n_1231)
);

NOR2xp33_ASAP7_75t_L g1232 ( 
.A(n_1111),
.B(n_1046),
.Y(n_1232)
);

BUFx10_ASAP7_75t_L g1233 ( 
.A(n_1045),
.Y(n_1233)
);

O2A1O1Ixp33_ASAP7_75t_L g1234 ( 
.A1(n_1071),
.A2(n_1010),
.B(n_1019),
.C(n_1012),
.Y(n_1234)
);

AOI21xp5_ASAP7_75t_L g1235 ( 
.A1(n_1158),
.A2(n_1137),
.B(n_1153),
.Y(n_1235)
);

AOI21xp5_ASAP7_75t_L g1236 ( 
.A1(n_1153),
.A2(n_1138),
.B(n_1010),
.Y(n_1236)
);

AOI21xp5_ASAP7_75t_L g1237 ( 
.A1(n_1019),
.A2(n_1025),
.B(n_1089),
.Y(n_1237)
);

AOI22xp5_ASAP7_75t_L g1238 ( 
.A1(n_1029),
.A2(n_1057),
.B1(n_1081),
.B2(n_1140),
.Y(n_1238)
);

OR2x6_ASAP7_75t_L g1239 ( 
.A(n_1045),
.B(n_1029),
.Y(n_1239)
);

OAI21x1_ASAP7_75t_L g1240 ( 
.A1(n_1076),
.A2(n_1026),
.B(n_1038),
.Y(n_1240)
);

AOI21xp5_ASAP7_75t_L g1241 ( 
.A1(n_1076),
.A2(n_1065),
.B(n_1044),
.Y(n_1241)
);

INVx2_ASAP7_75t_L g1242 ( 
.A(n_1050),
.Y(n_1242)
);

NAND2xp5_ASAP7_75t_SL g1243 ( 
.A(n_1062),
.B(n_1065),
.Y(n_1243)
);

OAI21xp5_ASAP7_75t_L g1244 ( 
.A1(n_1072),
.A2(n_1026),
.B(n_1038),
.Y(n_1244)
);

OAI22xp5_ASAP7_75t_L g1245 ( 
.A1(n_1051),
.A2(n_1060),
.B1(n_1079),
.B2(n_1095),
.Y(n_1245)
);

OA21x2_ASAP7_75t_L g1246 ( 
.A1(n_1103),
.A2(n_1044),
.B(n_1133),
.Y(n_1246)
);

INVx2_ASAP7_75t_SL g1247 ( 
.A(n_1118),
.Y(n_1247)
);

INVx1_ASAP7_75t_L g1248 ( 
.A(n_1133),
.Y(n_1248)
);

AO32x2_ASAP7_75t_L g1249 ( 
.A1(n_1133),
.A2(n_1128),
.A3(n_1146),
.B1(n_1147),
.B2(n_693),
.Y(n_1249)
);

OAI21xp5_ASAP7_75t_L g1250 ( 
.A1(n_1097),
.A2(n_1054),
.B(n_1049),
.Y(n_1250)
);

AOI21xp5_ASAP7_75t_SL g1251 ( 
.A1(n_1054),
.A2(n_1022),
.B(n_1110),
.Y(n_1251)
);

AND2x4_ASAP7_75t_L g1252 ( 
.A(n_1143),
.B(n_958),
.Y(n_1252)
);

AOI22xp33_ASAP7_75t_L g1253 ( 
.A1(n_1009),
.A2(n_811),
.B1(n_608),
.B2(n_599),
.Y(n_1253)
);

NAND2xp5_ASAP7_75t_L g1254 ( 
.A(n_1036),
.B(n_768),
.Y(n_1254)
);

NAND3xp33_ASAP7_75t_L g1255 ( 
.A(n_1084),
.B(n_564),
.C(n_1141),
.Y(n_1255)
);

INVx2_ASAP7_75t_SL g1256 ( 
.A(n_1008),
.Y(n_1256)
);

AOI21xp5_ASAP7_75t_L g1257 ( 
.A1(n_1054),
.A2(n_1083),
.B(n_1154),
.Y(n_1257)
);

NAND2xp5_ASAP7_75t_L g1258 ( 
.A(n_1036),
.B(n_768),
.Y(n_1258)
);

AOI221x1_ASAP7_75t_L g1259 ( 
.A1(n_1123),
.A2(n_1127),
.B1(n_1121),
.B2(n_1142),
.C(n_1084),
.Y(n_1259)
);

AOI21xp5_ASAP7_75t_L g1260 ( 
.A1(n_1054),
.A2(n_1083),
.B(n_1154),
.Y(n_1260)
);

O2A1O1Ixp33_ASAP7_75t_SL g1261 ( 
.A1(n_1054),
.A2(n_1125),
.B(n_1117),
.C(n_846),
.Y(n_1261)
);

OAI22xp5_ASAP7_75t_L g1262 ( 
.A1(n_1054),
.A2(n_1042),
.B1(n_1049),
.B2(n_1068),
.Y(n_1262)
);

AOI221xp5_ASAP7_75t_SL g1263 ( 
.A1(n_1123),
.A2(n_1127),
.B1(n_1049),
.B2(n_1042),
.C(n_1120),
.Y(n_1263)
);

AND2x2_ASAP7_75t_L g1264 ( 
.A(n_1009),
.B(n_677),
.Y(n_1264)
);

O2A1O1Ixp33_ASAP7_75t_SL g1265 ( 
.A1(n_1054),
.A2(n_1125),
.B(n_1117),
.C(n_846),
.Y(n_1265)
);

AOI21xp5_ASAP7_75t_L g1266 ( 
.A1(n_1054),
.A2(n_1083),
.B(n_1154),
.Y(n_1266)
);

A2O1A1Ixp33_ASAP7_75t_L g1267 ( 
.A1(n_1084),
.A2(n_510),
.B(n_1028),
.C(n_672),
.Y(n_1267)
);

A2O1A1Ixp33_ASAP7_75t_L g1268 ( 
.A1(n_1084),
.A2(n_510),
.B(n_1028),
.C(n_672),
.Y(n_1268)
);

A2O1A1Ixp33_ASAP7_75t_L g1269 ( 
.A1(n_1084),
.A2(n_510),
.B(n_1028),
.C(n_672),
.Y(n_1269)
);

BUFx10_ASAP7_75t_L g1270 ( 
.A(n_1018),
.Y(n_1270)
);

INVx2_ASAP7_75t_SL g1271 ( 
.A(n_1008),
.Y(n_1271)
);

NAND2xp5_ASAP7_75t_SL g1272 ( 
.A(n_1054),
.B(n_712),
.Y(n_1272)
);

AND2x4_ASAP7_75t_L g1273 ( 
.A(n_1143),
.B(n_958),
.Y(n_1273)
);

AOI21xp5_ASAP7_75t_L g1274 ( 
.A1(n_1054),
.A2(n_1083),
.B(n_1154),
.Y(n_1274)
);

OAI21x1_ASAP7_75t_L g1275 ( 
.A1(n_1067),
.A2(n_1155),
.B(n_1032),
.Y(n_1275)
);

AOI22xp5_ASAP7_75t_L g1276 ( 
.A1(n_1084),
.A2(n_712),
.B1(n_816),
.B2(n_773),
.Y(n_1276)
);

OAI22xp5_ASAP7_75t_L g1277 ( 
.A1(n_1054),
.A2(n_1042),
.B1(n_1049),
.B2(n_1068),
.Y(n_1277)
);

NAND2xp5_ASAP7_75t_L g1278 ( 
.A(n_1036),
.B(n_768),
.Y(n_1278)
);

AOI21xp5_ASAP7_75t_L g1279 ( 
.A1(n_1054),
.A2(n_1083),
.B(n_1154),
.Y(n_1279)
);

OAI21x1_ASAP7_75t_L g1280 ( 
.A1(n_1067),
.A2(n_1155),
.B(n_1032),
.Y(n_1280)
);

OAI21x1_ASAP7_75t_L g1281 ( 
.A1(n_1067),
.A2(n_1155),
.B(n_1032),
.Y(n_1281)
);

INVx2_ASAP7_75t_SL g1282 ( 
.A(n_1008),
.Y(n_1282)
);

AOI222xp33_ASAP7_75t_L g1283 ( 
.A1(n_1059),
.A2(n_599),
.B1(n_478),
.B2(n_811),
.C1(n_816),
.C2(n_716),
.Y(n_1283)
);

INVx1_ASAP7_75t_L g1284 ( 
.A(n_1015),
.Y(n_1284)
);

INVx1_ASAP7_75t_L g1285 ( 
.A(n_1015),
.Y(n_1285)
);

O2A1O1Ixp33_ASAP7_75t_SL g1286 ( 
.A1(n_1054),
.A2(n_1125),
.B(n_1117),
.C(n_846),
.Y(n_1286)
);

AOI21xp5_ASAP7_75t_L g1287 ( 
.A1(n_1054),
.A2(n_1083),
.B(n_1154),
.Y(n_1287)
);

NAND2xp5_ASAP7_75t_L g1288 ( 
.A(n_1036),
.B(n_768),
.Y(n_1288)
);

CKINVDCx11_ASAP7_75t_R g1289 ( 
.A(n_1057),
.Y(n_1289)
);

OA21x2_ASAP7_75t_L g1290 ( 
.A1(n_1155),
.A2(n_1037),
.B(n_1154),
.Y(n_1290)
);

NAND2xp5_ASAP7_75t_L g1291 ( 
.A(n_1036),
.B(n_768),
.Y(n_1291)
);

AOI21xp5_ASAP7_75t_L g1292 ( 
.A1(n_1054),
.A2(n_1083),
.B(n_1154),
.Y(n_1292)
);

INVx1_ASAP7_75t_L g1293 ( 
.A(n_1015),
.Y(n_1293)
);

INVxp67_ASAP7_75t_SL g1294 ( 
.A(n_1068),
.Y(n_1294)
);

NAND2xp5_ASAP7_75t_L g1295 ( 
.A(n_1036),
.B(n_768),
.Y(n_1295)
);

AO31x2_ASAP7_75t_L g1296 ( 
.A1(n_1083),
.A2(n_1096),
.A3(n_1154),
.B(n_953),
.Y(n_1296)
);

INVx1_ASAP7_75t_L g1297 ( 
.A(n_1015),
.Y(n_1297)
);

BUFx10_ASAP7_75t_L g1298 ( 
.A(n_1018),
.Y(n_1298)
);

INVx1_ASAP7_75t_L g1299 ( 
.A(n_1015),
.Y(n_1299)
);

INVx1_ASAP7_75t_L g1300 ( 
.A(n_1015),
.Y(n_1300)
);

AOI21x1_ASAP7_75t_L g1301 ( 
.A1(n_1037),
.A2(n_1032),
.B(n_1031),
.Y(n_1301)
);

NAND2x1_ASAP7_75t_L g1302 ( 
.A(n_1072),
.B(n_1153),
.Y(n_1302)
);

AOI21xp5_ASAP7_75t_L g1303 ( 
.A1(n_1054),
.A2(n_1083),
.B(n_1154),
.Y(n_1303)
);

INVx2_ASAP7_75t_L g1304 ( 
.A(n_1050),
.Y(n_1304)
);

NAND2xp5_ASAP7_75t_L g1305 ( 
.A(n_1036),
.B(n_768),
.Y(n_1305)
);

AND2x4_ASAP7_75t_L g1306 ( 
.A(n_1143),
.B(n_958),
.Y(n_1306)
);

AOI21xp5_ASAP7_75t_L g1307 ( 
.A1(n_1054),
.A2(n_1083),
.B(n_1154),
.Y(n_1307)
);

NAND3xp33_ASAP7_75t_L g1308 ( 
.A(n_1084),
.B(n_1141),
.C(n_1127),
.Y(n_1308)
);

AOI21xp5_ASAP7_75t_L g1309 ( 
.A1(n_1054),
.A2(n_1083),
.B(n_1154),
.Y(n_1309)
);

AO31x2_ASAP7_75t_L g1310 ( 
.A1(n_1083),
.A2(n_1096),
.A3(n_1154),
.B(n_953),
.Y(n_1310)
);

AOI21xp5_ASAP7_75t_L g1311 ( 
.A1(n_1054),
.A2(n_1083),
.B(n_1154),
.Y(n_1311)
);

NAND2xp5_ASAP7_75t_L g1312 ( 
.A(n_1036),
.B(n_768),
.Y(n_1312)
);

CKINVDCx16_ASAP7_75t_R g1313 ( 
.A(n_1143),
.Y(n_1313)
);

A2O1A1Ixp33_ASAP7_75t_L g1314 ( 
.A1(n_1084),
.A2(n_510),
.B(n_1028),
.C(n_672),
.Y(n_1314)
);

A2O1A1Ixp33_ASAP7_75t_L g1315 ( 
.A1(n_1084),
.A2(n_510),
.B(n_1028),
.C(n_672),
.Y(n_1315)
);

OAI21xp5_ASAP7_75t_L g1316 ( 
.A1(n_1054),
.A2(n_1049),
.B(n_1042),
.Y(n_1316)
);

AOI21xp5_ASAP7_75t_SL g1317 ( 
.A1(n_1054),
.A2(n_1022),
.B(n_1110),
.Y(n_1317)
);

BUFx4f_ASAP7_75t_SL g1318 ( 
.A(n_1046),
.Y(n_1318)
);

AOI21xp5_ASAP7_75t_L g1319 ( 
.A1(n_1054),
.A2(n_1083),
.B(n_1154),
.Y(n_1319)
);

INVx1_ASAP7_75t_L g1320 ( 
.A(n_1015),
.Y(n_1320)
);

AND2x2_ASAP7_75t_L g1321 ( 
.A(n_1166),
.B(n_1226),
.Y(n_1321)
);

NAND2x1p5_ASAP7_75t_L g1322 ( 
.A(n_1216),
.B(n_1243),
.Y(n_1322)
);

BUFx8_ASAP7_75t_SL g1323 ( 
.A(n_1191),
.Y(n_1323)
);

INVxp67_ASAP7_75t_SL g1324 ( 
.A(n_1294),
.Y(n_1324)
);

CKINVDCx20_ASAP7_75t_R g1325 ( 
.A(n_1289),
.Y(n_1325)
);

OAI22xp33_ASAP7_75t_L g1326 ( 
.A1(n_1204),
.A2(n_1255),
.B1(n_1308),
.B2(n_1276),
.Y(n_1326)
);

CKINVDCx6p67_ASAP7_75t_R g1327 ( 
.A(n_1313),
.Y(n_1327)
);

AOI22xp33_ASAP7_75t_L g1328 ( 
.A1(n_1253),
.A2(n_1283),
.B1(n_1198),
.B2(n_1308),
.Y(n_1328)
);

AOI22xp33_ASAP7_75t_L g1329 ( 
.A1(n_1204),
.A2(n_1276),
.B1(n_1264),
.B2(n_1272),
.Y(n_1329)
);

INVx2_ASAP7_75t_L g1330 ( 
.A(n_1246),
.Y(n_1330)
);

INVx3_ASAP7_75t_L g1331 ( 
.A(n_1227),
.Y(n_1331)
);

AND2x2_ASAP7_75t_L g1332 ( 
.A(n_1162),
.B(n_1170),
.Y(n_1332)
);

CKINVDCx20_ASAP7_75t_R g1333 ( 
.A(n_1318),
.Y(n_1333)
);

CKINVDCx11_ASAP7_75t_R g1334 ( 
.A(n_1270),
.Y(n_1334)
);

INVx2_ASAP7_75t_L g1335 ( 
.A(n_1168),
.Y(n_1335)
);

INVx2_ASAP7_75t_L g1336 ( 
.A(n_1168),
.Y(n_1336)
);

INVx2_ASAP7_75t_L g1337 ( 
.A(n_1168),
.Y(n_1337)
);

INVx2_ASAP7_75t_L g1338 ( 
.A(n_1301),
.Y(n_1338)
);

INVx1_ASAP7_75t_L g1339 ( 
.A(n_1174),
.Y(n_1339)
);

INVx1_ASAP7_75t_SL g1340 ( 
.A(n_1192),
.Y(n_1340)
);

AOI22xp33_ASAP7_75t_SL g1341 ( 
.A1(n_1179),
.A2(n_1211),
.B1(n_1262),
.B2(n_1277),
.Y(n_1341)
);

AOI22xp33_ASAP7_75t_L g1342 ( 
.A1(n_1225),
.A2(n_1179),
.B1(n_1221),
.B2(n_1242),
.Y(n_1342)
);

OAI22xp5_ASAP7_75t_L g1343 ( 
.A1(n_1267),
.A2(n_1269),
.B1(n_1268),
.B2(n_1315),
.Y(n_1343)
);

AOI22xp33_ASAP7_75t_L g1344 ( 
.A1(n_1304),
.A2(n_1224),
.B1(n_1247),
.B2(n_1184),
.Y(n_1344)
);

NAND2xp5_ASAP7_75t_L g1345 ( 
.A(n_1316),
.B(n_1254),
.Y(n_1345)
);

INVx4_ASAP7_75t_SL g1346 ( 
.A(n_1296),
.Y(n_1346)
);

AOI22xp33_ASAP7_75t_L g1347 ( 
.A1(n_1224),
.A2(n_1230),
.B1(n_1250),
.B2(n_1245),
.Y(n_1347)
);

BUFx3_ASAP7_75t_L g1348 ( 
.A(n_1165),
.Y(n_1348)
);

INVx2_ASAP7_75t_SL g1349 ( 
.A(n_1216),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_1284),
.Y(n_1350)
);

OAI22x1_ASAP7_75t_L g1351 ( 
.A1(n_1208),
.A2(n_1238),
.B1(n_1248),
.B2(n_1320),
.Y(n_1351)
);

OAI21xp5_ASAP7_75t_SL g1352 ( 
.A1(n_1197),
.A2(n_1314),
.B(n_1259),
.Y(n_1352)
);

OAI22xp5_ASAP7_75t_L g1353 ( 
.A1(n_1208),
.A2(n_1213),
.B1(n_1175),
.B2(n_1312),
.Y(n_1353)
);

OAI22xp5_ASAP7_75t_L g1354 ( 
.A1(n_1258),
.A2(n_1288),
.B1(n_1278),
.B2(n_1305),
.Y(n_1354)
);

INVxp67_ASAP7_75t_SL g1355 ( 
.A(n_1169),
.Y(n_1355)
);

AOI22xp5_ASAP7_75t_SL g1356 ( 
.A1(n_1202),
.A2(n_1252),
.B1(n_1306),
.B2(n_1273),
.Y(n_1356)
);

AOI22xp33_ASAP7_75t_SL g1357 ( 
.A1(n_1161),
.A2(n_1229),
.B1(n_1196),
.B2(n_1194),
.Y(n_1357)
);

NAND2x1p5_ASAP7_75t_L g1358 ( 
.A(n_1216),
.B(n_1238),
.Y(n_1358)
);

NAND2xp5_ASAP7_75t_L g1359 ( 
.A(n_1291),
.B(n_1295),
.Y(n_1359)
);

AOI22xp33_ASAP7_75t_L g1360 ( 
.A1(n_1176),
.A2(n_1297),
.B1(n_1293),
.B2(n_1299),
.Y(n_1360)
);

CKINVDCx6p67_ASAP7_75t_R g1361 ( 
.A(n_1270),
.Y(n_1361)
);

BUFx3_ASAP7_75t_L g1362 ( 
.A(n_1252),
.Y(n_1362)
);

AOI22xp33_ASAP7_75t_SL g1363 ( 
.A1(n_1273),
.A2(n_1306),
.B1(n_1189),
.B2(n_1285),
.Y(n_1363)
);

BUFx3_ASAP7_75t_L g1364 ( 
.A(n_1256),
.Y(n_1364)
);

CKINVDCx6p67_ASAP7_75t_R g1365 ( 
.A(n_1298),
.Y(n_1365)
);

AOI22xp33_ASAP7_75t_L g1366 ( 
.A1(n_1300),
.A2(n_1222),
.B1(n_1239),
.B2(n_1181),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_1214),
.Y(n_1367)
);

CKINVDCx5p33_ASAP7_75t_R g1368 ( 
.A(n_1180),
.Y(n_1368)
);

OAI22xp33_ASAP7_75t_SL g1369 ( 
.A1(n_1223),
.A2(n_1239),
.B1(n_1195),
.B2(n_1200),
.Y(n_1369)
);

AOI22xp33_ASAP7_75t_L g1370 ( 
.A1(n_1222),
.A2(n_1239),
.B1(n_1203),
.B2(n_1231),
.Y(n_1370)
);

AND2x2_ASAP7_75t_L g1371 ( 
.A(n_1214),
.B(n_1241),
.Y(n_1371)
);

INVx1_ASAP7_75t_L g1372 ( 
.A(n_1214),
.Y(n_1372)
);

CKINVDCx20_ASAP7_75t_R g1373 ( 
.A(n_1298),
.Y(n_1373)
);

BUFx2_ASAP7_75t_L g1374 ( 
.A(n_1167),
.Y(n_1374)
);

NAND2xp5_ASAP7_75t_L g1375 ( 
.A(n_1215),
.B(n_1232),
.Y(n_1375)
);

CKINVDCx20_ASAP7_75t_R g1376 ( 
.A(n_1271),
.Y(n_1376)
);

BUFx6f_ASAP7_75t_L g1377 ( 
.A(n_1233),
.Y(n_1377)
);

INVx1_ASAP7_75t_L g1378 ( 
.A(n_1220),
.Y(n_1378)
);

AND2x2_ASAP7_75t_L g1379 ( 
.A(n_1249),
.B(n_1263),
.Y(n_1379)
);

BUFx3_ASAP7_75t_L g1380 ( 
.A(n_1282),
.Y(n_1380)
);

CKINVDCx5p33_ASAP7_75t_R g1381 ( 
.A(n_1233),
.Y(n_1381)
);

AND2x2_ASAP7_75t_L g1382 ( 
.A(n_1249),
.B(n_1310),
.Y(n_1382)
);

BUFx12f_ASAP7_75t_L g1383 ( 
.A(n_1167),
.Y(n_1383)
);

INVx2_ASAP7_75t_SL g1384 ( 
.A(n_1173),
.Y(n_1384)
);

INVx3_ASAP7_75t_L g1385 ( 
.A(n_1310),
.Y(n_1385)
);

AOI22xp33_ASAP7_75t_L g1386 ( 
.A1(n_1201),
.A2(n_1235),
.B1(n_1237),
.B2(n_1236),
.Y(n_1386)
);

BUFx6f_ASAP7_75t_L g1387 ( 
.A(n_1302),
.Y(n_1387)
);

AOI22xp33_ASAP7_75t_L g1388 ( 
.A1(n_1205),
.A2(n_1209),
.B1(n_1244),
.B2(n_1217),
.Y(n_1388)
);

AOI22xp33_ASAP7_75t_L g1389 ( 
.A1(n_1257),
.A2(n_1287),
.B1(n_1311),
.B2(n_1260),
.Y(n_1389)
);

NAND2xp5_ASAP7_75t_L g1390 ( 
.A(n_1251),
.B(n_1317),
.Y(n_1390)
);

OAI22xp33_ASAP7_75t_L g1391 ( 
.A1(n_1212),
.A2(n_1303),
.B1(n_1279),
.B2(n_1266),
.Y(n_1391)
);

INVx1_ASAP7_75t_L g1392 ( 
.A(n_1240),
.Y(n_1392)
);

INVx2_ASAP7_75t_L g1393 ( 
.A(n_1186),
.Y(n_1393)
);

OAI22xp33_ASAP7_75t_L g1394 ( 
.A1(n_1274),
.A2(n_1319),
.B1(n_1307),
.B2(n_1292),
.Y(n_1394)
);

INVx1_ASAP7_75t_SL g1395 ( 
.A(n_1178),
.Y(n_1395)
);

INVxp67_ASAP7_75t_SL g1396 ( 
.A(n_1309),
.Y(n_1396)
);

INVx1_ASAP7_75t_L g1397 ( 
.A(n_1234),
.Y(n_1397)
);

BUFx8_ASAP7_75t_L g1398 ( 
.A(n_1249),
.Y(n_1398)
);

NAND2xp5_ASAP7_75t_L g1399 ( 
.A(n_1228),
.B(n_1207),
.Y(n_1399)
);

AOI22xp5_ASAP7_75t_L g1400 ( 
.A1(n_1210),
.A2(n_1182),
.B1(n_1261),
.B2(n_1286),
.Y(n_1400)
);

HB1xp67_ASAP7_75t_L g1401 ( 
.A(n_1177),
.Y(n_1401)
);

INVx6_ASAP7_75t_L g1402 ( 
.A(n_1265),
.Y(n_1402)
);

INVx6_ASAP7_75t_L g1403 ( 
.A(n_1199),
.Y(n_1403)
);

BUFx4f_ASAP7_75t_SL g1404 ( 
.A(n_1185),
.Y(n_1404)
);

INVx6_ASAP7_75t_L g1405 ( 
.A(n_1171),
.Y(n_1405)
);

AOI22xp5_ASAP7_75t_L g1406 ( 
.A1(n_1219),
.A2(n_1183),
.B1(n_1190),
.B2(n_1218),
.Y(n_1406)
);

INVx1_ASAP7_75t_L g1407 ( 
.A(n_1177),
.Y(n_1407)
);

BUFx3_ASAP7_75t_L g1408 ( 
.A(n_1275),
.Y(n_1408)
);

BUFx2_ASAP7_75t_SL g1409 ( 
.A(n_1290),
.Y(n_1409)
);

NAND2xp5_ASAP7_75t_L g1410 ( 
.A(n_1290),
.B(n_1177),
.Y(n_1410)
);

BUFx3_ASAP7_75t_L g1411 ( 
.A(n_1280),
.Y(n_1411)
);

AOI22xp33_ASAP7_75t_L g1412 ( 
.A1(n_1164),
.A2(n_1188),
.B1(n_1163),
.B2(n_1281),
.Y(n_1412)
);

AOI22xp33_ASAP7_75t_L g1413 ( 
.A1(n_1172),
.A2(n_1206),
.B1(n_1193),
.B2(n_1187),
.Y(n_1413)
);

OAI21xp33_ASAP7_75t_L g1414 ( 
.A1(n_1206),
.A2(n_1187),
.B(n_1193),
.Y(n_1414)
);

CKINVDCx6p67_ASAP7_75t_R g1415 ( 
.A(n_1206),
.Y(n_1415)
);

AOI22xp33_ASAP7_75t_SL g1416 ( 
.A1(n_1193),
.A2(n_478),
.B1(n_811),
.B2(n_338),
.Y(n_1416)
);

CKINVDCx6p67_ASAP7_75t_R g1417 ( 
.A(n_1187),
.Y(n_1417)
);

BUFx12f_ASAP7_75t_L g1418 ( 
.A(n_1289),
.Y(n_1418)
);

OAI22xp5_ASAP7_75t_L g1419 ( 
.A1(n_1204),
.A2(n_1042),
.B1(n_1049),
.B2(n_1255),
.Y(n_1419)
);

CKINVDCx6p67_ASAP7_75t_R g1420 ( 
.A(n_1289),
.Y(n_1420)
);

BUFx10_ASAP7_75t_L g1421 ( 
.A(n_1180),
.Y(n_1421)
);

AOI22xp33_ASAP7_75t_L g1422 ( 
.A1(n_1253),
.A2(n_811),
.B1(n_1283),
.B2(n_608),
.Y(n_1422)
);

OAI22xp5_ASAP7_75t_L g1423 ( 
.A1(n_1204),
.A2(n_1042),
.B1(n_1049),
.B2(n_1255),
.Y(n_1423)
);

INVxp67_ASAP7_75t_SL g1424 ( 
.A(n_1294),
.Y(n_1424)
);

BUFx10_ASAP7_75t_L g1425 ( 
.A(n_1180),
.Y(n_1425)
);

INVx6_ASAP7_75t_L g1426 ( 
.A(n_1216),
.Y(n_1426)
);

BUFx3_ASAP7_75t_L g1427 ( 
.A(n_1165),
.Y(n_1427)
);

INVx1_ASAP7_75t_SL g1428 ( 
.A(n_1192),
.Y(n_1428)
);

INVx6_ASAP7_75t_L g1429 ( 
.A(n_1216),
.Y(n_1429)
);

INVx1_ASAP7_75t_SL g1430 ( 
.A(n_1192),
.Y(n_1430)
);

AOI22xp5_ASAP7_75t_L g1431 ( 
.A1(n_1204),
.A2(n_712),
.B1(n_1198),
.B2(n_1255),
.Y(n_1431)
);

AND2x2_ASAP7_75t_L g1432 ( 
.A(n_1166),
.B(n_1226),
.Y(n_1432)
);

OAI22xp33_ASAP7_75t_L g1433 ( 
.A1(n_1204),
.A2(n_1255),
.B1(n_1124),
.B2(n_478),
.Y(n_1433)
);

OAI221xp5_ASAP7_75t_L g1434 ( 
.A1(n_1204),
.A2(n_1255),
.B1(n_1268),
.B2(n_1269),
.C(n_1267),
.Y(n_1434)
);

AOI22xp5_ASAP7_75t_L g1435 ( 
.A1(n_1204),
.A2(n_712),
.B1(n_1198),
.B2(n_1255),
.Y(n_1435)
);

BUFx6f_ASAP7_75t_L g1436 ( 
.A(n_1239),
.Y(n_1436)
);

INVx2_ASAP7_75t_SL g1437 ( 
.A(n_1216),
.Y(n_1437)
);

AOI22xp33_ASAP7_75t_L g1438 ( 
.A1(n_1253),
.A2(n_811),
.B1(n_1283),
.B2(n_608),
.Y(n_1438)
);

CKINVDCx20_ASAP7_75t_R g1439 ( 
.A(n_1289),
.Y(n_1439)
);

INVx2_ASAP7_75t_SL g1440 ( 
.A(n_1216),
.Y(n_1440)
);

BUFx6f_ASAP7_75t_L g1441 ( 
.A(n_1239),
.Y(n_1441)
);

CKINVDCx11_ASAP7_75t_R g1442 ( 
.A(n_1289),
.Y(n_1442)
);

OAI22xp5_ASAP7_75t_L g1443 ( 
.A1(n_1204),
.A2(n_1042),
.B1(n_1049),
.B2(n_1255),
.Y(n_1443)
);

INVx2_ASAP7_75t_SL g1444 ( 
.A(n_1216),
.Y(n_1444)
);

INVx2_ASAP7_75t_SL g1445 ( 
.A(n_1216),
.Y(n_1445)
);

OAI22xp33_ASAP7_75t_L g1446 ( 
.A1(n_1204),
.A2(n_1255),
.B1(n_1124),
.B2(n_478),
.Y(n_1446)
);

INVx1_ASAP7_75t_L g1447 ( 
.A(n_1162),
.Y(n_1447)
);

BUFx4_ASAP7_75t_SL g1448 ( 
.A(n_1191),
.Y(n_1448)
);

AOI21x1_ASAP7_75t_L g1449 ( 
.A1(n_1390),
.A2(n_1343),
.B(n_1338),
.Y(n_1449)
);

NAND2xp5_ASAP7_75t_L g1450 ( 
.A(n_1321),
.B(n_1432),
.Y(n_1450)
);

AO32x2_ASAP7_75t_L g1451 ( 
.A1(n_1353),
.A2(n_1354),
.A3(n_1443),
.B1(n_1419),
.B2(n_1423),
.Y(n_1451)
);

AOI21x1_ASAP7_75t_L g1452 ( 
.A1(n_1338),
.A2(n_1399),
.B(n_1410),
.Y(n_1452)
);

INVx1_ASAP7_75t_L g1453 ( 
.A(n_1330),
.Y(n_1453)
);

OAI21x1_ASAP7_75t_L g1454 ( 
.A1(n_1412),
.A2(n_1389),
.B(n_1413),
.Y(n_1454)
);

INVx1_ASAP7_75t_L g1455 ( 
.A(n_1330),
.Y(n_1455)
);

INVx1_ASAP7_75t_L g1456 ( 
.A(n_1355),
.Y(n_1456)
);

INVx1_ASAP7_75t_L g1457 ( 
.A(n_1379),
.Y(n_1457)
);

AND2x4_ASAP7_75t_L g1458 ( 
.A(n_1346),
.B(n_1392),
.Y(n_1458)
);

INVx1_ASAP7_75t_L g1459 ( 
.A(n_1379),
.Y(n_1459)
);

CKINVDCx6p67_ASAP7_75t_R g1460 ( 
.A(n_1333),
.Y(n_1460)
);

A2O1A1Ixp33_ASAP7_75t_L g1461 ( 
.A1(n_1328),
.A2(n_1431),
.B(n_1435),
.C(n_1352),
.Y(n_1461)
);

INVx1_ASAP7_75t_L g1462 ( 
.A(n_1371),
.Y(n_1462)
);

INVx3_ASAP7_75t_L g1463 ( 
.A(n_1403),
.Y(n_1463)
);

INVx4_ASAP7_75t_SL g1464 ( 
.A(n_1404),
.Y(n_1464)
);

INVx1_ASAP7_75t_L g1465 ( 
.A(n_1371),
.Y(n_1465)
);

BUFx3_ASAP7_75t_L g1466 ( 
.A(n_1358),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_1407),
.Y(n_1467)
);

AND2x2_ASAP7_75t_L g1468 ( 
.A(n_1321),
.B(n_1432),
.Y(n_1468)
);

AO21x2_ASAP7_75t_L g1469 ( 
.A1(n_1414),
.A2(n_1391),
.B(n_1337),
.Y(n_1469)
);

AND2x2_ASAP7_75t_L g1470 ( 
.A(n_1382),
.B(n_1332),
.Y(n_1470)
);

OR2x2_ASAP7_75t_L g1471 ( 
.A(n_1324),
.B(n_1424),
.Y(n_1471)
);

NOR2xp33_ASAP7_75t_L g1472 ( 
.A(n_1368),
.B(n_1340),
.Y(n_1472)
);

BUFx2_ASAP7_75t_L g1473 ( 
.A(n_1403),
.Y(n_1473)
);

NAND2xp5_ASAP7_75t_L g1474 ( 
.A(n_1357),
.B(n_1341),
.Y(n_1474)
);

OR2x2_ASAP7_75t_L g1475 ( 
.A(n_1367),
.B(n_1372),
.Y(n_1475)
);

OAI21x1_ASAP7_75t_L g1476 ( 
.A1(n_1393),
.A2(n_1406),
.B(n_1386),
.Y(n_1476)
);

AOI22xp33_ASAP7_75t_L g1477 ( 
.A1(n_1422),
.A2(n_1438),
.B1(n_1416),
.B2(n_1398),
.Y(n_1477)
);

HB1xp67_ASAP7_75t_L g1478 ( 
.A(n_1332),
.Y(n_1478)
);

INVx1_ASAP7_75t_L g1479 ( 
.A(n_1401),
.Y(n_1479)
);

OAI21xp33_ASAP7_75t_L g1480 ( 
.A1(n_1434),
.A2(n_1326),
.B(n_1329),
.Y(n_1480)
);

INVx1_ASAP7_75t_SL g1481 ( 
.A(n_1374),
.Y(n_1481)
);

INVx3_ASAP7_75t_L g1482 ( 
.A(n_1403),
.Y(n_1482)
);

HB1xp67_ASAP7_75t_L g1483 ( 
.A(n_1339),
.Y(n_1483)
);

OAI21x1_ASAP7_75t_L g1484 ( 
.A1(n_1393),
.A2(n_1331),
.B(n_1336),
.Y(n_1484)
);

NAND2xp5_ASAP7_75t_L g1485 ( 
.A(n_1359),
.B(n_1345),
.Y(n_1485)
);

AOI22xp33_ASAP7_75t_L g1486 ( 
.A1(n_1398),
.A2(n_1433),
.B1(n_1446),
.B2(n_1342),
.Y(n_1486)
);

BUFx2_ASAP7_75t_SL g1487 ( 
.A(n_1349),
.Y(n_1487)
);

INVx1_ASAP7_75t_L g1488 ( 
.A(n_1350),
.Y(n_1488)
);

INVx1_ASAP7_75t_SL g1489 ( 
.A(n_1362),
.Y(n_1489)
);

AOI22xp33_ASAP7_75t_SL g1490 ( 
.A1(n_1398),
.A2(n_1356),
.B1(n_1375),
.B2(n_1402),
.Y(n_1490)
);

INVx4_ASAP7_75t_L g1491 ( 
.A(n_1402),
.Y(n_1491)
);

INVx1_ASAP7_75t_L g1492 ( 
.A(n_1447),
.Y(n_1492)
);

AOI221xp5_ASAP7_75t_L g1493 ( 
.A1(n_1351),
.A2(n_1360),
.B1(n_1347),
.B2(n_1397),
.C(n_1363),
.Y(n_1493)
);

BUFx6f_ASAP7_75t_L g1494 ( 
.A(n_1405),
.Y(n_1494)
);

AOI21xp5_ASAP7_75t_L g1495 ( 
.A1(n_1394),
.A2(n_1396),
.B(n_1395),
.Y(n_1495)
);

BUFx8_ASAP7_75t_SL g1496 ( 
.A(n_1323),
.Y(n_1496)
);

AND2x4_ASAP7_75t_L g1497 ( 
.A(n_1346),
.B(n_1331),
.Y(n_1497)
);

HB1xp67_ASAP7_75t_L g1498 ( 
.A(n_1378),
.Y(n_1498)
);

AOI21xp33_ASAP7_75t_L g1499 ( 
.A1(n_1400),
.A2(n_1366),
.B(n_1335),
.Y(n_1499)
);

HB1xp67_ASAP7_75t_L g1500 ( 
.A(n_1384),
.Y(n_1500)
);

INVx1_ASAP7_75t_L g1501 ( 
.A(n_1385),
.Y(n_1501)
);

BUFx6f_ASAP7_75t_L g1502 ( 
.A(n_1405),
.Y(n_1502)
);

INVx1_ASAP7_75t_L g1503 ( 
.A(n_1385),
.Y(n_1503)
);

INVx1_ASAP7_75t_L g1504 ( 
.A(n_1331),
.Y(n_1504)
);

OR2x2_ASAP7_75t_L g1505 ( 
.A(n_1417),
.B(n_1415),
.Y(n_1505)
);

OR2x2_ASAP7_75t_L g1506 ( 
.A(n_1417),
.B(n_1415),
.Y(n_1506)
);

AND2x2_ASAP7_75t_L g1507 ( 
.A(n_1346),
.B(n_1370),
.Y(n_1507)
);

NAND2xp5_ASAP7_75t_L g1508 ( 
.A(n_1344),
.B(n_1388),
.Y(n_1508)
);

CKINVDCx20_ASAP7_75t_R g1509 ( 
.A(n_1323),
.Y(n_1509)
);

INVx1_ASAP7_75t_L g1510 ( 
.A(n_1409),
.Y(n_1510)
);

INVx2_ASAP7_75t_L g1511 ( 
.A(n_1408),
.Y(n_1511)
);

NAND2xp5_ASAP7_75t_L g1512 ( 
.A(n_1428),
.B(n_1430),
.Y(n_1512)
);

OAI21x1_ASAP7_75t_L g1513 ( 
.A1(n_1322),
.A2(n_1411),
.B(n_1402),
.Y(n_1513)
);

INVx1_ASAP7_75t_L g1514 ( 
.A(n_1411),
.Y(n_1514)
);

AO21x2_ASAP7_75t_L g1515 ( 
.A1(n_1402),
.A2(n_1369),
.B(n_1387),
.Y(n_1515)
);

INVx1_ASAP7_75t_L g1516 ( 
.A(n_1387),
.Y(n_1516)
);

HB1xp67_ASAP7_75t_L g1517 ( 
.A(n_1348),
.Y(n_1517)
);

BUFx2_ASAP7_75t_L g1518 ( 
.A(n_1383),
.Y(n_1518)
);

INVxp67_ASAP7_75t_SL g1519 ( 
.A(n_1437),
.Y(n_1519)
);

INVx1_ASAP7_75t_L g1520 ( 
.A(n_1437),
.Y(n_1520)
);

INVx2_ASAP7_75t_SL g1521 ( 
.A(n_1426),
.Y(n_1521)
);

BUFx2_ASAP7_75t_SL g1522 ( 
.A(n_1440),
.Y(n_1522)
);

AND2x2_ASAP7_75t_L g1523 ( 
.A(n_1468),
.B(n_1327),
.Y(n_1523)
);

AND2x2_ASAP7_75t_L g1524 ( 
.A(n_1468),
.B(n_1470),
.Y(n_1524)
);

AND2x2_ASAP7_75t_L g1525 ( 
.A(n_1470),
.B(n_1327),
.Y(n_1525)
);

INVx4_ASAP7_75t_L g1526 ( 
.A(n_1464),
.Y(n_1526)
);

NOR2xp33_ASAP7_75t_L g1527 ( 
.A(n_1474),
.B(n_1427),
.Y(n_1527)
);

NOR2xp33_ASAP7_75t_L g1528 ( 
.A(n_1474),
.B(n_1427),
.Y(n_1528)
);

AND2x2_ASAP7_75t_L g1529 ( 
.A(n_1478),
.B(n_1348),
.Y(n_1529)
);

NOR2xp33_ASAP7_75t_L g1530 ( 
.A(n_1480),
.B(n_1365),
.Y(n_1530)
);

NAND2xp5_ASAP7_75t_L g1531 ( 
.A(n_1485),
.B(n_1364),
.Y(n_1531)
);

BUFx4f_ASAP7_75t_SL g1532 ( 
.A(n_1509),
.Y(n_1532)
);

AND2x2_ASAP7_75t_L g1533 ( 
.A(n_1450),
.B(n_1364),
.Y(n_1533)
);

INVx1_ASAP7_75t_L g1534 ( 
.A(n_1483),
.Y(n_1534)
);

A2O1A1Ixp33_ASAP7_75t_L g1535 ( 
.A1(n_1461),
.A2(n_1445),
.B(n_1444),
.C(n_1440),
.Y(n_1535)
);

AOI22xp5_ASAP7_75t_L g1536 ( 
.A1(n_1480),
.A2(n_1373),
.B1(n_1376),
.B2(n_1436),
.Y(n_1536)
);

AND2x2_ASAP7_75t_L g1537 ( 
.A(n_1517),
.B(n_1380),
.Y(n_1537)
);

NOR2xp33_ASAP7_75t_L g1538 ( 
.A(n_1481),
.B(n_1361),
.Y(n_1538)
);

OA21x2_ASAP7_75t_L g1539 ( 
.A1(n_1476),
.A2(n_1381),
.B(n_1429),
.Y(n_1539)
);

BUFx8_ASAP7_75t_SL g1540 ( 
.A(n_1496),
.Y(n_1540)
);

HB1xp67_ASAP7_75t_L g1541 ( 
.A(n_1471),
.Y(n_1541)
);

OAI21xp5_ASAP7_75t_L g1542 ( 
.A1(n_1495),
.A2(n_1373),
.B(n_1376),
.Y(n_1542)
);

OA21x2_ASAP7_75t_L g1543 ( 
.A1(n_1454),
.A2(n_1381),
.B(n_1429),
.Y(n_1543)
);

OAI21xp5_ASAP7_75t_L g1544 ( 
.A1(n_1508),
.A2(n_1368),
.B(n_1439),
.Y(n_1544)
);

NAND2xp5_ASAP7_75t_L g1545 ( 
.A(n_1481),
.B(n_1365),
.Y(n_1545)
);

OAI22xp5_ASAP7_75t_L g1546 ( 
.A1(n_1486),
.A2(n_1361),
.B1(n_1420),
.B2(n_1439),
.Y(n_1546)
);

O2A1O1Ixp33_ASAP7_75t_L g1547 ( 
.A1(n_1508),
.A2(n_1333),
.B(n_1325),
.C(n_1448),
.Y(n_1547)
);

INVxp67_ASAP7_75t_L g1548 ( 
.A(n_1500),
.Y(n_1548)
);

OAI211xp5_ASAP7_75t_SL g1549 ( 
.A1(n_1512),
.A2(n_1334),
.B(n_1442),
.C(n_1421),
.Y(n_1549)
);

INVx1_ASAP7_75t_L g1550 ( 
.A(n_1488),
.Y(n_1550)
);

OAI21xp5_ASAP7_75t_L g1551 ( 
.A1(n_1493),
.A2(n_1325),
.B(n_1334),
.Y(n_1551)
);

OAI21xp5_ASAP7_75t_L g1552 ( 
.A1(n_1449),
.A2(n_1451),
.B(n_1499),
.Y(n_1552)
);

AO21x1_ASAP7_75t_SL g1553 ( 
.A1(n_1457),
.A2(n_1442),
.B(n_1418),
.Y(n_1553)
);

A2O1A1Ixp33_ASAP7_75t_L g1554 ( 
.A1(n_1451),
.A2(n_1441),
.B(n_1377),
.C(n_1418),
.Y(n_1554)
);

INVxp67_ASAP7_75t_SL g1555 ( 
.A(n_1471),
.Y(n_1555)
);

OAI21xp5_ASAP7_75t_L g1556 ( 
.A1(n_1449),
.A2(n_1425),
.B(n_1377),
.Y(n_1556)
);

AND2x2_ASAP7_75t_L g1557 ( 
.A(n_1462),
.B(n_1377),
.Y(n_1557)
);

AOI21xp5_ASAP7_75t_L g1558 ( 
.A1(n_1491),
.A2(n_1441),
.B(n_1469),
.Y(n_1558)
);

BUFx3_ASAP7_75t_L g1559 ( 
.A(n_1518),
.Y(n_1559)
);

NOR2xp33_ASAP7_75t_L g1560 ( 
.A(n_1491),
.B(n_1473),
.Y(n_1560)
);

AO32x2_ASAP7_75t_L g1561 ( 
.A1(n_1521),
.A2(n_1491),
.A3(n_1459),
.B1(n_1462),
.B2(n_1465),
.Y(n_1561)
);

OAI22xp5_ASAP7_75t_L g1562 ( 
.A1(n_1477),
.A2(n_1490),
.B1(n_1451),
.B2(n_1482),
.Y(n_1562)
);

OAI22xp5_ASAP7_75t_L g1563 ( 
.A1(n_1451),
.A2(n_1463),
.B1(n_1482),
.B2(n_1518),
.Y(n_1563)
);

OA21x2_ASAP7_75t_L g1564 ( 
.A1(n_1454),
.A2(n_1484),
.B(n_1499),
.Y(n_1564)
);

AND2x4_ASAP7_75t_L g1565 ( 
.A(n_1497),
.B(n_1473),
.Y(n_1565)
);

HB1xp67_ASAP7_75t_L g1566 ( 
.A(n_1452),
.Y(n_1566)
);

OR2x2_ASAP7_75t_L g1567 ( 
.A(n_1475),
.B(n_1492),
.Y(n_1567)
);

AND2x4_ASAP7_75t_L g1568 ( 
.A(n_1497),
.B(n_1458),
.Y(n_1568)
);

AOI221xp5_ASAP7_75t_L g1569 ( 
.A1(n_1456),
.A2(n_1492),
.B1(n_1479),
.B2(n_1467),
.C(n_1514),
.Y(n_1569)
);

AND2x4_ASAP7_75t_L g1570 ( 
.A(n_1458),
.B(n_1507),
.Y(n_1570)
);

OR2x2_ASAP7_75t_L g1571 ( 
.A(n_1475),
.B(n_1456),
.Y(n_1571)
);

AND2x4_ASAP7_75t_L g1572 ( 
.A(n_1458),
.B(n_1507),
.Y(n_1572)
);

A2O1A1Ixp33_ASAP7_75t_L g1573 ( 
.A1(n_1464),
.A2(n_1513),
.B(n_1505),
.C(n_1506),
.Y(n_1573)
);

NOR2xp33_ASAP7_75t_L g1574 ( 
.A(n_1530),
.B(n_1472),
.Y(n_1574)
);

OR2x2_ASAP7_75t_L g1575 ( 
.A(n_1541),
.B(n_1469),
.Y(n_1575)
);

AOI22xp33_ASAP7_75t_L g1576 ( 
.A1(n_1551),
.A2(n_1464),
.B1(n_1515),
.B2(n_1469),
.Y(n_1576)
);

OAI222xp33_ASAP7_75t_L g1577 ( 
.A1(n_1562),
.A2(n_1506),
.B1(n_1489),
.B2(n_1466),
.C1(n_1453),
.C2(n_1455),
.Y(n_1577)
);

AOI22xp33_ASAP7_75t_L g1578 ( 
.A1(n_1552),
.A2(n_1464),
.B1(n_1515),
.B2(n_1469),
.Y(n_1578)
);

NAND2xp5_ASAP7_75t_L g1579 ( 
.A(n_1555),
.B(n_1479),
.Y(n_1579)
);

BUFx2_ASAP7_75t_L g1580 ( 
.A(n_1561),
.Y(n_1580)
);

AND2x2_ASAP7_75t_L g1581 ( 
.A(n_1561),
.B(n_1504),
.Y(n_1581)
);

OR2x2_ASAP7_75t_L g1582 ( 
.A(n_1541),
.B(n_1510),
.Y(n_1582)
);

OR2x2_ASAP7_75t_L g1583 ( 
.A(n_1571),
.B(n_1567),
.Y(n_1583)
);

AND2x2_ASAP7_75t_L g1584 ( 
.A(n_1561),
.B(n_1504),
.Y(n_1584)
);

NAND2xp5_ASAP7_75t_SL g1585 ( 
.A(n_1554),
.B(n_1464),
.Y(n_1585)
);

INVx2_ASAP7_75t_L g1586 ( 
.A(n_1561),
.Y(n_1586)
);

INVx2_ASAP7_75t_L g1587 ( 
.A(n_1550),
.Y(n_1587)
);

AOI22xp33_ASAP7_75t_L g1588 ( 
.A1(n_1527),
.A2(n_1515),
.B1(n_1467),
.B2(n_1498),
.Y(n_1588)
);

AND2x2_ASAP7_75t_L g1589 ( 
.A(n_1524),
.B(n_1511),
.Y(n_1589)
);

AOI22xp33_ASAP7_75t_L g1590 ( 
.A1(n_1527),
.A2(n_1515),
.B1(n_1494),
.B2(n_1502),
.Y(n_1590)
);

HB1xp67_ASAP7_75t_L g1591 ( 
.A(n_1548),
.Y(n_1591)
);

AND2x4_ASAP7_75t_L g1592 ( 
.A(n_1568),
.B(n_1458),
.Y(n_1592)
);

NAND2xp5_ASAP7_75t_SL g1593 ( 
.A(n_1554),
.B(n_1563),
.Y(n_1593)
);

BUFx2_ASAP7_75t_L g1594 ( 
.A(n_1565),
.Y(n_1594)
);

OAI221xp5_ASAP7_75t_L g1595 ( 
.A1(n_1535),
.A2(n_1510),
.B1(n_1514),
.B2(n_1516),
.C(n_1519),
.Y(n_1595)
);

OAI22xp5_ASAP7_75t_L g1596 ( 
.A1(n_1536),
.A2(n_1522),
.B1(n_1487),
.B2(n_1460),
.Y(n_1596)
);

INVx1_ASAP7_75t_L g1597 ( 
.A(n_1534),
.Y(n_1597)
);

HB1xp67_ASAP7_75t_L g1598 ( 
.A(n_1548),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1566),
.Y(n_1599)
);

NAND2xp5_ASAP7_75t_L g1600 ( 
.A(n_1569),
.B(n_1452),
.Y(n_1600)
);

INVx1_ASAP7_75t_L g1601 ( 
.A(n_1566),
.Y(n_1601)
);

AND2x2_ASAP7_75t_L g1602 ( 
.A(n_1594),
.B(n_1529),
.Y(n_1602)
);

INVx1_ASAP7_75t_L g1603 ( 
.A(n_1587),
.Y(n_1603)
);

INVx1_ASAP7_75t_L g1604 ( 
.A(n_1587),
.Y(n_1604)
);

INVx1_ASAP7_75t_L g1605 ( 
.A(n_1587),
.Y(n_1605)
);

INVx2_ASAP7_75t_L g1606 ( 
.A(n_1581),
.Y(n_1606)
);

NOR2xp67_ASAP7_75t_L g1607 ( 
.A(n_1575),
.B(n_1526),
.Y(n_1607)
);

INVx2_ASAP7_75t_L g1608 ( 
.A(n_1581),
.Y(n_1608)
);

AOI221x1_ASAP7_75t_L g1609 ( 
.A1(n_1600),
.A2(n_1535),
.B1(n_1546),
.B2(n_1549),
.C(n_1556),
.Y(n_1609)
);

OAI31xp33_ASAP7_75t_L g1610 ( 
.A1(n_1593),
.A2(n_1528),
.A3(n_1573),
.B(n_1525),
.Y(n_1610)
);

INVx2_ASAP7_75t_L g1611 ( 
.A(n_1581),
.Y(n_1611)
);

HB1xp67_ASAP7_75t_L g1612 ( 
.A(n_1591),
.Y(n_1612)
);

INVx2_ASAP7_75t_SL g1613 ( 
.A(n_1592),
.Y(n_1613)
);

AOI22xp5_ASAP7_75t_L g1614 ( 
.A1(n_1593),
.A2(n_1528),
.B1(n_1542),
.B2(n_1531),
.Y(n_1614)
);

AOI21xp5_ASAP7_75t_L g1615 ( 
.A1(n_1600),
.A2(n_1543),
.B(n_1558),
.Y(n_1615)
);

HB1xp67_ASAP7_75t_L g1616 ( 
.A(n_1591),
.Y(n_1616)
);

HB1xp67_ASAP7_75t_L g1617 ( 
.A(n_1598),
.Y(n_1617)
);

INVxp67_ASAP7_75t_L g1618 ( 
.A(n_1598),
.Y(n_1618)
);

INVx2_ASAP7_75t_L g1619 ( 
.A(n_1584),
.Y(n_1619)
);

INVxp67_ASAP7_75t_L g1620 ( 
.A(n_1574),
.Y(n_1620)
);

OAI33xp33_ASAP7_75t_L g1621 ( 
.A1(n_1575),
.A2(n_1545),
.A3(n_1547),
.B1(n_1520),
.B2(n_1501),
.B3(n_1503),
.Y(n_1621)
);

NAND4xp75_ASAP7_75t_L g1622 ( 
.A(n_1585),
.B(n_1544),
.C(n_1543),
.D(n_1539),
.Y(n_1622)
);

NAND2xp5_ASAP7_75t_L g1623 ( 
.A(n_1579),
.B(n_1533),
.Y(n_1623)
);

INVx2_ASAP7_75t_L g1624 ( 
.A(n_1584),
.Y(n_1624)
);

AND2x2_ASAP7_75t_L g1625 ( 
.A(n_1594),
.B(n_1537),
.Y(n_1625)
);

INVx1_ASAP7_75t_SL g1626 ( 
.A(n_1582),
.Y(n_1626)
);

OAI22xp5_ASAP7_75t_L g1627 ( 
.A1(n_1580),
.A2(n_1523),
.B1(n_1526),
.B2(n_1560),
.Y(n_1627)
);

BUFx3_ASAP7_75t_L g1628 ( 
.A(n_1592),
.Y(n_1628)
);

INVx1_ASAP7_75t_L g1629 ( 
.A(n_1599),
.Y(n_1629)
);

INVx1_ASAP7_75t_L g1630 ( 
.A(n_1599),
.Y(n_1630)
);

NAND2xp5_ASAP7_75t_L g1631 ( 
.A(n_1579),
.B(n_1557),
.Y(n_1631)
);

AOI22xp33_ASAP7_75t_L g1632 ( 
.A1(n_1576),
.A2(n_1572),
.B1(n_1570),
.B2(n_1543),
.Y(n_1632)
);

OAI221xp5_ASAP7_75t_L g1633 ( 
.A1(n_1576),
.A2(n_1573),
.B1(n_1564),
.B2(n_1539),
.C(n_1538),
.Y(n_1633)
);

AND2x2_ASAP7_75t_L g1634 ( 
.A(n_1606),
.B(n_1580),
.Y(n_1634)
);

INVxp67_ASAP7_75t_SL g1635 ( 
.A(n_1612),
.Y(n_1635)
);

INVx2_ASAP7_75t_L g1636 ( 
.A(n_1606),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_1629),
.Y(n_1637)
);

AND2x2_ASAP7_75t_L g1638 ( 
.A(n_1606),
.B(n_1580),
.Y(n_1638)
);

INVx1_ASAP7_75t_SL g1639 ( 
.A(n_1616),
.Y(n_1639)
);

AND2x4_ASAP7_75t_L g1640 ( 
.A(n_1628),
.B(n_1586),
.Y(n_1640)
);

OR2x2_ASAP7_75t_L g1641 ( 
.A(n_1626),
.B(n_1583),
.Y(n_1641)
);

BUFx3_ASAP7_75t_L g1642 ( 
.A(n_1629),
.Y(n_1642)
);

OR2x2_ASAP7_75t_L g1643 ( 
.A(n_1626),
.B(n_1583),
.Y(n_1643)
);

NAND3xp33_ASAP7_75t_SL g1644 ( 
.A(n_1610),
.B(n_1574),
.C(n_1586),
.Y(n_1644)
);

INVx1_ASAP7_75t_L g1645 ( 
.A(n_1630),
.Y(n_1645)
);

NAND2xp5_ASAP7_75t_L g1646 ( 
.A(n_1630),
.B(n_1586),
.Y(n_1646)
);

NAND2xp5_ASAP7_75t_L g1647 ( 
.A(n_1617),
.B(n_1586),
.Y(n_1647)
);

NAND2xp5_ASAP7_75t_L g1648 ( 
.A(n_1618),
.B(n_1601),
.Y(n_1648)
);

OR2x2_ASAP7_75t_L g1649 ( 
.A(n_1608),
.B(n_1601),
.Y(n_1649)
);

NAND2xp5_ASAP7_75t_L g1650 ( 
.A(n_1620),
.B(n_1597),
.Y(n_1650)
);

OR2x2_ASAP7_75t_L g1651 ( 
.A(n_1608),
.B(n_1583),
.Y(n_1651)
);

OR2x2_ASAP7_75t_L g1652 ( 
.A(n_1611),
.B(n_1582),
.Y(n_1652)
);

INVx1_ASAP7_75t_L g1653 ( 
.A(n_1603),
.Y(n_1653)
);

INVx1_ASAP7_75t_L g1654 ( 
.A(n_1604),
.Y(n_1654)
);

OR2x2_ASAP7_75t_L g1655 ( 
.A(n_1611),
.B(n_1582),
.Y(n_1655)
);

INVx1_ASAP7_75t_L g1656 ( 
.A(n_1605),
.Y(n_1656)
);

AND2x4_ASAP7_75t_SL g1657 ( 
.A(n_1625),
.B(n_1592),
.Y(n_1657)
);

BUFx2_ASAP7_75t_L g1658 ( 
.A(n_1628),
.Y(n_1658)
);

INVx4_ASAP7_75t_L g1659 ( 
.A(n_1628),
.Y(n_1659)
);

AND2x4_ASAP7_75t_L g1660 ( 
.A(n_1613),
.B(n_1592),
.Y(n_1660)
);

AND2x2_ASAP7_75t_L g1661 ( 
.A(n_1619),
.B(n_1624),
.Y(n_1661)
);

AND2x2_ASAP7_75t_L g1662 ( 
.A(n_1624),
.B(n_1589),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_1637),
.Y(n_1663)
);

INVx2_ASAP7_75t_L g1664 ( 
.A(n_1661),
.Y(n_1664)
);

NAND2xp5_ASAP7_75t_L g1665 ( 
.A(n_1639),
.B(n_1614),
.Y(n_1665)
);

OR2x2_ASAP7_75t_L g1666 ( 
.A(n_1641),
.B(n_1624),
.Y(n_1666)
);

NAND2xp5_ASAP7_75t_L g1667 ( 
.A(n_1639),
.B(n_1614),
.Y(n_1667)
);

AND2x4_ASAP7_75t_L g1668 ( 
.A(n_1657),
.B(n_1613),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_1650),
.Y(n_1669)
);

NAND2xp5_ASAP7_75t_L g1670 ( 
.A(n_1650),
.B(n_1610),
.Y(n_1670)
);

AOI322xp5_ASAP7_75t_L g1671 ( 
.A1(n_1644),
.A2(n_1632),
.A3(n_1578),
.B1(n_1588),
.B2(n_1585),
.C1(n_1609),
.C2(n_1590),
.Y(n_1671)
);

NAND2xp5_ASAP7_75t_L g1672 ( 
.A(n_1635),
.B(n_1609),
.Y(n_1672)
);

INVx1_ASAP7_75t_L g1673 ( 
.A(n_1637),
.Y(n_1673)
);

INVxp67_ASAP7_75t_SL g1674 ( 
.A(n_1642),
.Y(n_1674)
);

INVx1_ASAP7_75t_L g1675 ( 
.A(n_1645),
.Y(n_1675)
);

OR2x2_ASAP7_75t_L g1676 ( 
.A(n_1641),
.B(n_1623),
.Y(n_1676)
);

INVx2_ASAP7_75t_L g1677 ( 
.A(n_1661),
.Y(n_1677)
);

NAND2x1p5_ASAP7_75t_L g1678 ( 
.A(n_1659),
.B(n_1539),
.Y(n_1678)
);

OR2x2_ASAP7_75t_L g1679 ( 
.A(n_1643),
.B(n_1623),
.Y(n_1679)
);

INVx1_ASAP7_75t_L g1680 ( 
.A(n_1645),
.Y(n_1680)
);

INVx2_ASAP7_75t_SL g1681 ( 
.A(n_1657),
.Y(n_1681)
);

INVx1_ASAP7_75t_L g1682 ( 
.A(n_1643),
.Y(n_1682)
);

INVx1_ASAP7_75t_L g1683 ( 
.A(n_1646),
.Y(n_1683)
);

AND2x2_ASAP7_75t_L g1684 ( 
.A(n_1657),
.B(n_1613),
.Y(n_1684)
);

HB1xp67_ASAP7_75t_L g1685 ( 
.A(n_1642),
.Y(n_1685)
);

INVx1_ASAP7_75t_L g1686 ( 
.A(n_1642),
.Y(n_1686)
);

NOR2xp67_ASAP7_75t_L g1687 ( 
.A(n_1644),
.B(n_1633),
.Y(n_1687)
);

OR2x2_ASAP7_75t_L g1688 ( 
.A(n_1651),
.B(n_1631),
.Y(n_1688)
);

HB1xp67_ASAP7_75t_L g1689 ( 
.A(n_1648),
.Y(n_1689)
);

O2A1O1Ixp33_ASAP7_75t_L g1690 ( 
.A1(n_1635),
.A2(n_1633),
.B(n_1615),
.C(n_1621),
.Y(n_1690)
);

AND2x2_ASAP7_75t_L g1691 ( 
.A(n_1660),
.B(n_1625),
.Y(n_1691)
);

INVx2_ASAP7_75t_L g1692 ( 
.A(n_1661),
.Y(n_1692)
);

INVx2_ASAP7_75t_L g1693 ( 
.A(n_1636),
.Y(n_1693)
);

OR2x2_ASAP7_75t_L g1694 ( 
.A(n_1651),
.B(n_1631),
.Y(n_1694)
);

INVx1_ASAP7_75t_L g1695 ( 
.A(n_1646),
.Y(n_1695)
);

AND2x2_ASAP7_75t_L g1696 ( 
.A(n_1660),
.B(n_1602),
.Y(n_1696)
);

INVx1_ASAP7_75t_L g1697 ( 
.A(n_1653),
.Y(n_1697)
);

NOR4xp25_ASAP7_75t_L g1698 ( 
.A(n_1647),
.B(n_1597),
.C(n_1595),
.D(n_1627),
.Y(n_1698)
);

INVx1_ASAP7_75t_L g1699 ( 
.A(n_1648),
.Y(n_1699)
);

INVxp67_ASAP7_75t_SL g1700 ( 
.A(n_1647),
.Y(n_1700)
);

INVx1_ASAP7_75t_L g1701 ( 
.A(n_1653),
.Y(n_1701)
);

INVx1_ASAP7_75t_L g1702 ( 
.A(n_1654),
.Y(n_1702)
);

AND2x2_ASAP7_75t_L g1703 ( 
.A(n_1660),
.B(n_1602),
.Y(n_1703)
);

INVx1_ASAP7_75t_L g1704 ( 
.A(n_1654),
.Y(n_1704)
);

INVx1_ASAP7_75t_L g1705 ( 
.A(n_1656),
.Y(n_1705)
);

OR2x2_ASAP7_75t_L g1706 ( 
.A(n_1676),
.B(n_1652),
.Y(n_1706)
);

NAND2xp5_ASAP7_75t_L g1707 ( 
.A(n_1670),
.B(n_1662),
.Y(n_1707)
);

NAND2xp5_ASAP7_75t_L g1708 ( 
.A(n_1665),
.B(n_1667),
.Y(n_1708)
);

OR2x2_ASAP7_75t_L g1709 ( 
.A(n_1676),
.B(n_1652),
.Y(n_1709)
);

INVx1_ASAP7_75t_L g1710 ( 
.A(n_1663),
.Y(n_1710)
);

NAND2xp5_ASAP7_75t_L g1711 ( 
.A(n_1672),
.B(n_1662),
.Y(n_1711)
);

NAND2xp5_ASAP7_75t_L g1712 ( 
.A(n_1669),
.B(n_1662),
.Y(n_1712)
);

INVx2_ASAP7_75t_L g1713 ( 
.A(n_1664),
.Y(n_1713)
);

AND2x2_ASAP7_75t_L g1714 ( 
.A(n_1691),
.B(n_1660),
.Y(n_1714)
);

NAND2xp5_ASAP7_75t_L g1715 ( 
.A(n_1698),
.B(n_1634),
.Y(n_1715)
);

NAND2x1_ASAP7_75t_L g1716 ( 
.A(n_1668),
.B(n_1681),
.Y(n_1716)
);

BUFx2_ASAP7_75t_L g1717 ( 
.A(n_1674),
.Y(n_1717)
);

OAI22xp33_ASAP7_75t_L g1718 ( 
.A1(n_1687),
.A2(n_1615),
.B1(n_1595),
.B2(n_1575),
.Y(n_1718)
);

NAND2x2_ASAP7_75t_L g1719 ( 
.A(n_1681),
.B(n_1540),
.Y(n_1719)
);

AND2x2_ASAP7_75t_L g1720 ( 
.A(n_1691),
.B(n_1660),
.Y(n_1720)
);

INVx1_ASAP7_75t_SL g1721 ( 
.A(n_1685),
.Y(n_1721)
);

AOI22xp33_ASAP7_75t_L g1722 ( 
.A1(n_1682),
.A2(n_1578),
.B1(n_1621),
.B2(n_1640),
.Y(n_1722)
);

AND2x2_ASAP7_75t_L g1723 ( 
.A(n_1696),
.B(n_1658),
.Y(n_1723)
);

OR2x2_ASAP7_75t_L g1724 ( 
.A(n_1679),
.B(n_1652),
.Y(n_1724)
);

AND2x2_ASAP7_75t_L g1725 ( 
.A(n_1696),
.B(n_1658),
.Y(n_1725)
);

INVx2_ASAP7_75t_L g1726 ( 
.A(n_1664),
.Y(n_1726)
);

OAI211xp5_ASAP7_75t_L g1727 ( 
.A1(n_1690),
.A2(n_1659),
.B(n_1538),
.C(n_1559),
.Y(n_1727)
);

NAND2xp5_ASAP7_75t_L g1728 ( 
.A(n_1689),
.B(n_1634),
.Y(n_1728)
);

NOR2x1p5_ASAP7_75t_L g1729 ( 
.A(n_1682),
.B(n_1659),
.Y(n_1729)
);

OR2x2_ASAP7_75t_L g1730 ( 
.A(n_1679),
.B(n_1655),
.Y(n_1730)
);

INVx1_ASAP7_75t_L g1731 ( 
.A(n_1663),
.Y(n_1731)
);

OR2x2_ASAP7_75t_L g1732 ( 
.A(n_1688),
.B(n_1655),
.Y(n_1732)
);

NAND2xp5_ASAP7_75t_L g1733 ( 
.A(n_1699),
.B(n_1634),
.Y(n_1733)
);

INVx2_ASAP7_75t_L g1734 ( 
.A(n_1677),
.Y(n_1734)
);

INVx2_ASAP7_75t_L g1735 ( 
.A(n_1677),
.Y(n_1735)
);

NAND2xp5_ASAP7_75t_L g1736 ( 
.A(n_1686),
.B(n_1638),
.Y(n_1736)
);

AND2x2_ASAP7_75t_L g1737 ( 
.A(n_1703),
.B(n_1659),
.Y(n_1737)
);

OR2x2_ASAP7_75t_L g1738 ( 
.A(n_1688),
.B(n_1655),
.Y(n_1738)
);

AND2x2_ASAP7_75t_L g1739 ( 
.A(n_1703),
.B(n_1640),
.Y(n_1739)
);

OR2x2_ASAP7_75t_L g1740 ( 
.A(n_1694),
.B(n_1649),
.Y(n_1740)
);

INVx1_ASAP7_75t_L g1741 ( 
.A(n_1673),
.Y(n_1741)
);

NOR2xp67_ASAP7_75t_SL g1742 ( 
.A(n_1727),
.B(n_1622),
.Y(n_1742)
);

NAND2xp5_ASAP7_75t_L g1743 ( 
.A(n_1721),
.B(n_1700),
.Y(n_1743)
);

HB1xp67_ASAP7_75t_L g1744 ( 
.A(n_1717),
.Y(n_1744)
);

NAND2xp5_ASAP7_75t_L g1745 ( 
.A(n_1721),
.B(n_1692),
.Y(n_1745)
);

AND2x2_ASAP7_75t_L g1746 ( 
.A(n_1723),
.B(n_1668),
.Y(n_1746)
);

NAND2xp5_ASAP7_75t_L g1747 ( 
.A(n_1717),
.B(n_1692),
.Y(n_1747)
);

AOI221xp5_ASAP7_75t_L g1748 ( 
.A1(n_1715),
.A2(n_1683),
.B1(n_1695),
.B2(n_1638),
.C(n_1705),
.Y(n_1748)
);

OAI21xp5_ASAP7_75t_L g1749 ( 
.A1(n_1718),
.A2(n_1671),
.B(n_1622),
.Y(n_1749)
);

INVx1_ASAP7_75t_SL g1750 ( 
.A(n_1708),
.Y(n_1750)
);

AOI22xp33_ASAP7_75t_L g1751 ( 
.A1(n_1722),
.A2(n_1678),
.B1(n_1693),
.B2(n_1640),
.Y(n_1751)
);

NAND2xp5_ASAP7_75t_L g1752 ( 
.A(n_1707),
.B(n_1694),
.Y(n_1752)
);

INVx2_ASAP7_75t_L g1753 ( 
.A(n_1713),
.Y(n_1753)
);

INVxp67_ASAP7_75t_L g1754 ( 
.A(n_1716),
.Y(n_1754)
);

OAI31xp33_ASAP7_75t_L g1755 ( 
.A1(n_1711),
.A2(n_1678),
.A3(n_1729),
.B(n_1577),
.Y(n_1755)
);

AOI211xp5_ASAP7_75t_SL g1756 ( 
.A1(n_1723),
.A2(n_1532),
.B(n_1596),
.C(n_1540),
.Y(n_1756)
);

AND2x2_ASAP7_75t_L g1757 ( 
.A(n_1725),
.B(n_1668),
.Y(n_1757)
);

NOR2xp33_ASAP7_75t_L g1758 ( 
.A(n_1716),
.B(n_1532),
.Y(n_1758)
);

INVx1_ASAP7_75t_L g1759 ( 
.A(n_1710),
.Y(n_1759)
);

NOR2xp33_ASAP7_75t_L g1760 ( 
.A(n_1706),
.B(n_1709),
.Y(n_1760)
);

INVx1_ASAP7_75t_L g1761 ( 
.A(n_1710),
.Y(n_1761)
);

BUFx2_ASAP7_75t_L g1762 ( 
.A(n_1729),
.Y(n_1762)
);

OAI31xp33_ASAP7_75t_SL g1763 ( 
.A1(n_1725),
.A2(n_1596),
.A3(n_1640),
.B(n_1684),
.Y(n_1763)
);

INVx1_ASAP7_75t_L g1764 ( 
.A(n_1731),
.Y(n_1764)
);

AOI22xp33_ASAP7_75t_L g1765 ( 
.A1(n_1713),
.A2(n_1734),
.B1(n_1735),
.B2(n_1726),
.Y(n_1765)
);

OAI22xp33_ASAP7_75t_L g1766 ( 
.A1(n_1706),
.A2(n_1678),
.B1(n_1666),
.B2(n_1607),
.Y(n_1766)
);

INVx1_ASAP7_75t_L g1767 ( 
.A(n_1731),
.Y(n_1767)
);

NAND2xp5_ASAP7_75t_L g1768 ( 
.A(n_1760),
.B(n_1726),
.Y(n_1768)
);

AOI22xp33_ASAP7_75t_SL g1769 ( 
.A1(n_1749),
.A2(n_1728),
.B1(n_1739),
.B2(n_1733),
.Y(n_1769)
);

INVx1_ASAP7_75t_L g1770 ( 
.A(n_1744),
.Y(n_1770)
);

OAI221xp5_ASAP7_75t_SL g1771 ( 
.A1(n_1755),
.A2(n_1724),
.B1(n_1709),
.B2(n_1730),
.C(n_1738),
.Y(n_1771)
);

NAND2xp5_ASAP7_75t_SL g1772 ( 
.A(n_1763),
.B(n_1737),
.Y(n_1772)
);

INVx2_ASAP7_75t_L g1773 ( 
.A(n_1753),
.Y(n_1773)
);

OAI221xp5_ASAP7_75t_L g1774 ( 
.A1(n_1755),
.A2(n_1719),
.B1(n_1736),
.B2(n_1724),
.C(n_1730),
.Y(n_1774)
);

INVxp67_ASAP7_75t_L g1775 ( 
.A(n_1758),
.Y(n_1775)
);

AND2x2_ASAP7_75t_L g1776 ( 
.A(n_1746),
.B(n_1739),
.Y(n_1776)
);

NAND2xp5_ASAP7_75t_L g1777 ( 
.A(n_1750),
.B(n_1734),
.Y(n_1777)
);

NAND2xp5_ASAP7_75t_L g1778 ( 
.A(n_1748),
.B(n_1735),
.Y(n_1778)
);

INVx1_ASAP7_75t_L g1779 ( 
.A(n_1753),
.Y(n_1779)
);

INVx1_ASAP7_75t_L g1780 ( 
.A(n_1753),
.Y(n_1780)
);

INVx1_ASAP7_75t_L g1781 ( 
.A(n_1759),
.Y(n_1781)
);

INVx3_ASAP7_75t_L g1782 ( 
.A(n_1746),
.Y(n_1782)
);

AOI21xp33_ASAP7_75t_L g1783 ( 
.A1(n_1750),
.A2(n_1743),
.B(n_1742),
.Y(n_1783)
);

HB1xp67_ASAP7_75t_L g1784 ( 
.A(n_1754),
.Y(n_1784)
);

INVx3_ASAP7_75t_L g1785 ( 
.A(n_1757),
.Y(n_1785)
);

NAND2xp5_ASAP7_75t_L g1786 ( 
.A(n_1752),
.B(n_1765),
.Y(n_1786)
);

HB1xp67_ASAP7_75t_L g1787 ( 
.A(n_1745),
.Y(n_1787)
);

INVx1_ASAP7_75t_L g1788 ( 
.A(n_1779),
.Y(n_1788)
);

OAI22xp5_ASAP7_75t_L g1789 ( 
.A1(n_1771),
.A2(n_1719),
.B1(n_1751),
.B2(n_1732),
.Y(n_1789)
);

AO22x2_ASAP7_75t_L g1790 ( 
.A1(n_1770),
.A2(n_1767),
.B1(n_1764),
.B2(n_1759),
.Y(n_1790)
);

AOI22xp5_ASAP7_75t_L g1791 ( 
.A1(n_1774),
.A2(n_1742),
.B1(n_1757),
.B2(n_1747),
.Y(n_1791)
);

INVx1_ASAP7_75t_L g1792 ( 
.A(n_1779),
.Y(n_1792)
);

INVx1_ASAP7_75t_L g1793 ( 
.A(n_1780),
.Y(n_1793)
);

AOI22xp5_ASAP7_75t_L g1794 ( 
.A1(n_1783),
.A2(n_1766),
.B1(n_1719),
.B2(n_1762),
.Y(n_1794)
);

NAND2xp5_ASAP7_75t_L g1795 ( 
.A(n_1782),
.B(n_1762),
.Y(n_1795)
);

INVxp67_ASAP7_75t_SL g1796 ( 
.A(n_1782),
.Y(n_1796)
);

A2O1A1Ixp33_ASAP7_75t_L g1797 ( 
.A1(n_1783),
.A2(n_1763),
.B(n_1756),
.C(n_1767),
.Y(n_1797)
);

INVx1_ASAP7_75t_L g1798 ( 
.A(n_1780),
.Y(n_1798)
);

XOR2xp5_ASAP7_75t_L g1799 ( 
.A(n_1769),
.B(n_1732),
.Y(n_1799)
);

INVx2_ASAP7_75t_SL g1800 ( 
.A(n_1795),
.Y(n_1800)
);

NAND4xp25_ASAP7_75t_L g1801 ( 
.A(n_1791),
.B(n_1785),
.C(n_1782),
.D(n_1775),
.Y(n_1801)
);

INVx1_ASAP7_75t_L g1802 ( 
.A(n_1790),
.Y(n_1802)
);

AOI211x1_ASAP7_75t_L g1803 ( 
.A1(n_1789),
.A2(n_1778),
.B(n_1772),
.C(n_1786),
.Y(n_1803)
);

OR2x2_ASAP7_75t_L g1804 ( 
.A(n_1796),
.B(n_1768),
.Y(n_1804)
);

NAND2xp5_ASAP7_75t_L g1805 ( 
.A(n_1799),
.B(n_1785),
.Y(n_1805)
);

NAND2xp5_ASAP7_75t_L g1806 ( 
.A(n_1797),
.B(n_1785),
.Y(n_1806)
);

NOR2xp33_ASAP7_75t_L g1807 ( 
.A(n_1794),
.B(n_1776),
.Y(n_1807)
);

AOI21xp5_ASAP7_75t_L g1808 ( 
.A1(n_1790),
.A2(n_1778),
.B(n_1777),
.Y(n_1808)
);

AND2x2_ASAP7_75t_L g1809 ( 
.A(n_1788),
.B(n_1776),
.Y(n_1809)
);

OAI211xp5_ASAP7_75t_L g1810 ( 
.A1(n_1792),
.A2(n_1787),
.B(n_1784),
.C(n_1770),
.Y(n_1810)
);

NAND4xp25_ASAP7_75t_L g1811 ( 
.A(n_1803),
.B(n_1756),
.C(n_1781),
.D(n_1793),
.Y(n_1811)
);

INVx1_ASAP7_75t_L g1812 ( 
.A(n_1809),
.Y(n_1812)
);

AOI22xp5_ASAP7_75t_L g1813 ( 
.A1(n_1802),
.A2(n_1773),
.B1(n_1798),
.B2(n_1781),
.Y(n_1813)
);

NOR2x1_ASAP7_75t_L g1814 ( 
.A(n_1801),
.B(n_1773),
.Y(n_1814)
);

AND4x1_ASAP7_75t_L g1815 ( 
.A(n_1807),
.B(n_1764),
.C(n_1761),
.D(n_1737),
.Y(n_1815)
);

AOI22xp5_ASAP7_75t_L g1816 ( 
.A1(n_1814),
.A2(n_1808),
.B1(n_1805),
.B2(n_1806),
.Y(n_1816)
);

AOI22xp5_ASAP7_75t_L g1817 ( 
.A1(n_1813),
.A2(n_1800),
.B1(n_1804),
.B2(n_1810),
.Y(n_1817)
);

AOI311xp33_ASAP7_75t_L g1818 ( 
.A1(n_1812),
.A2(n_1761),
.A3(n_1741),
.B(n_1733),
.C(n_1675),
.Y(n_1818)
);

OAI22xp5_ASAP7_75t_L g1819 ( 
.A1(n_1815),
.A2(n_1738),
.B1(n_1740),
.B2(n_1712),
.Y(n_1819)
);

OAI211xp5_ASAP7_75t_SL g1820 ( 
.A1(n_1811),
.A2(n_1741),
.B(n_1740),
.C(n_1683),
.Y(n_1820)
);

NAND2xp5_ASAP7_75t_SL g1821 ( 
.A(n_1815),
.B(n_1714),
.Y(n_1821)
);

INVx2_ASAP7_75t_L g1822 ( 
.A(n_1821),
.Y(n_1822)
);

NOR2x1_ASAP7_75t_L g1823 ( 
.A(n_1820),
.B(n_1673),
.Y(n_1823)
);

INVx1_ASAP7_75t_L g1824 ( 
.A(n_1819),
.Y(n_1824)
);

INVx1_ASAP7_75t_L g1825 ( 
.A(n_1817),
.Y(n_1825)
);

XNOR2x1_ASAP7_75t_L g1826 ( 
.A(n_1816),
.B(n_1666),
.Y(n_1826)
);

BUFx3_ASAP7_75t_L g1827 ( 
.A(n_1825),
.Y(n_1827)
);

NAND2xp5_ASAP7_75t_L g1828 ( 
.A(n_1822),
.B(n_1675),
.Y(n_1828)
);

AOI322xp5_ASAP7_75t_L g1829 ( 
.A1(n_1823),
.A2(n_1818),
.A3(n_1638),
.B1(n_1695),
.B2(n_1693),
.C1(n_1640),
.C2(n_1702),
.Y(n_1829)
);

INVx2_ASAP7_75t_L g1830 ( 
.A(n_1827),
.Y(n_1830)
);

HB1xp67_ASAP7_75t_L g1831 ( 
.A(n_1830),
.Y(n_1831)
);

INVx1_ASAP7_75t_L g1832 ( 
.A(n_1831),
.Y(n_1832)
);

AOI22xp5_ASAP7_75t_L g1833 ( 
.A1(n_1831),
.A2(n_1826),
.B1(n_1824),
.B2(n_1828),
.Y(n_1833)
);

CKINVDCx20_ASAP7_75t_R g1834 ( 
.A(n_1833),
.Y(n_1834)
);

INVx1_ASAP7_75t_L g1835 ( 
.A(n_1832),
.Y(n_1835)
);

OAI22xp5_ASAP7_75t_L g1836 ( 
.A1(n_1835),
.A2(n_1829),
.B1(n_1720),
.B2(n_1714),
.Y(n_1836)
);

AOI22xp33_ASAP7_75t_L g1837 ( 
.A1(n_1834),
.A2(n_1705),
.B1(n_1704),
.B2(n_1702),
.Y(n_1837)
);

AOI22xp5_ASAP7_75t_L g1838 ( 
.A1(n_1836),
.A2(n_1720),
.B1(n_1704),
.B2(n_1701),
.Y(n_1838)
);

OAI21xp5_ASAP7_75t_L g1839 ( 
.A1(n_1838),
.A2(n_1837),
.B(n_1701),
.Y(n_1839)
);

INVx1_ASAP7_75t_L g1840 ( 
.A(n_1839),
.Y(n_1840)
);

OAI221xp5_ASAP7_75t_R g1841 ( 
.A1(n_1840),
.A2(n_1553),
.B1(n_1680),
.B2(n_1697),
.C(n_1684),
.Y(n_1841)
);

AOI211xp5_ASAP7_75t_L g1842 ( 
.A1(n_1841),
.A2(n_1680),
.B(n_1697),
.C(n_1559),
.Y(n_1842)
);


endmodule