module fake_netlist_1_7392_n_39 (n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_39);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_39;
wire n_20;
wire n_38;
wire n_36;
wire n_37;
wire n_34;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_11;
wire n_25;
wire n_30;
wire n_26;
wire n_13;
wire n_16;
wire n_33;
wire n_18;
wire n_32;
wire n_35;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_27;
CKINVDCx5p33_ASAP7_75t_R g11 ( .A(n_6), .Y(n_11) );
CKINVDCx5p33_ASAP7_75t_R g12 ( .A(n_8), .Y(n_12) );
CKINVDCx5p33_ASAP7_75t_R g13 ( .A(n_6), .Y(n_13) );
CKINVDCx5p33_ASAP7_75t_R g14 ( .A(n_1), .Y(n_14) );
CKINVDCx5p33_ASAP7_75t_R g15 ( .A(n_1), .Y(n_15) );
CKINVDCx20_ASAP7_75t_R g16 ( .A(n_8), .Y(n_16) );
CKINVDCx20_ASAP7_75t_R g17 ( .A(n_2), .Y(n_17) );
OAI22xp5_ASAP7_75t_L g18 ( .A1(n_14), .A2(n_0), .B1(n_1), .B2(n_2), .Y(n_18) );
AOI21xp5_ASAP7_75t_L g19 ( .A1(n_15), .A2(n_0), .B(n_2), .Y(n_19) );
BUFx2_ASAP7_75t_L g20 ( .A(n_17), .Y(n_20) );
O2A1O1Ixp5_ASAP7_75t_L g21 ( .A1(n_13), .A2(n_0), .B(n_3), .C(n_4), .Y(n_21) );
NAND2xp5_ASAP7_75t_SL g22 ( .A(n_11), .B(n_3), .Y(n_22) );
OAI21xp5_ASAP7_75t_L g23 ( .A1(n_19), .A2(n_13), .B(n_12), .Y(n_23) );
NOR2xp33_ASAP7_75t_R g24 ( .A(n_20), .B(n_17), .Y(n_24) );
NAND2xp33_ASAP7_75t_R g25 ( .A(n_21), .B(n_4), .Y(n_25) );
NAND2xp5_ASAP7_75t_L g26 ( .A(n_23), .B(n_22), .Y(n_26) );
INVx1_ASAP7_75t_L g27 ( .A(n_23), .Y(n_27) );
HB1xp67_ASAP7_75t_L g28 ( .A(n_24), .Y(n_28) );
A2O1A1Ixp33_ASAP7_75t_L g29 ( .A1(n_27), .A2(n_18), .B(n_22), .C(n_25), .Y(n_29) );
INVx1_ASAP7_75t_L g30 ( .A(n_27), .Y(n_30) );
INVx2_ASAP7_75t_L g31 ( .A(n_30), .Y(n_31) );
OAI221xp5_ASAP7_75t_L g32 ( .A1(n_29), .A2(n_28), .B1(n_26), .B2(n_16), .C(n_10), .Y(n_32) );
INVx1_ASAP7_75t_SL g33 ( .A(n_31), .Y(n_33) );
CKINVDCx16_ASAP7_75t_R g34 ( .A(n_32), .Y(n_34) );
NAND2x1p5_ASAP7_75t_L g35 ( .A(n_31), .B(n_30), .Y(n_35) );
AO22x2_ASAP7_75t_L g36 ( .A1(n_33), .A2(n_26), .B1(n_16), .B2(n_9), .Y(n_36) );
OR3x2_ASAP7_75t_L g37 ( .A(n_34), .B(n_5), .C(n_7), .Y(n_37) );
INVx2_ASAP7_75t_L g38 ( .A(n_35), .Y(n_38) );
AOI222xp33_ASAP7_75t_L g39 ( .A1(n_36), .A2(n_5), .B1(n_10), .B2(n_35), .C1(n_37), .C2(n_38), .Y(n_39) );
endmodule