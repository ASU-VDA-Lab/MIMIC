module fake_netlist_5_896_n_1988 (n_137, n_294, n_431, n_318, n_380, n_419, n_444, n_469, n_82, n_194, n_316, n_389, n_418, n_248, n_124, n_86, n_136, n_146, n_315, n_268, n_451, n_408, n_61, n_376, n_127, n_75, n_235, n_226, n_74, n_57, n_353, n_351, n_367, n_452, n_397, n_111, n_483, n_155, n_43, n_116, n_22, n_467, n_423, n_284, n_46, n_245, n_21, n_139, n_38, n_105, n_280, n_4, n_378, n_17, n_382, n_254, n_33, n_23, n_302, n_265, n_293, n_372, n_443, n_244, n_47, n_173, n_198, n_447, n_247, n_314, n_368, n_433, n_8, n_321, n_292, n_100, n_455, n_417, n_212, n_385, n_119, n_275, n_252, n_26, n_295, n_133, n_330, n_2, n_6, n_39, n_147, n_373, n_67, n_307, n_439, n_87, n_150, n_106, n_209, n_259, n_448, n_375, n_301, n_68, n_93, n_186, n_134, n_191, n_51, n_63, n_171, n_153, n_399, n_341, n_204, n_394, n_250, n_260, n_298, n_320, n_286, n_122, n_282, n_331, n_10, n_24, n_406, n_470, n_325, n_449, n_132, n_90, n_101, n_281, n_240, n_381, n_189, n_220, n_291, n_231, n_257, n_390, n_31, n_456, n_13, n_371, n_481, n_152, n_317, n_9, n_323, n_195, n_42, n_356, n_227, n_45, n_271, n_94, n_335, n_123, n_370, n_167, n_234, n_343, n_308, n_379, n_428, n_267, n_457, n_297, n_156, n_5, n_225, n_377, n_484, n_219, n_442, n_157, n_131, n_192, n_223, n_392, n_158, n_138, n_264, n_109, n_472, n_454, n_387, n_374, n_163, n_276, n_339, n_95, n_183, n_185, n_243, n_398, n_396, n_347, n_169, n_59, n_255, n_215, n_350, n_196, n_459, n_211, n_218, n_400, n_181, n_436, n_3, n_290, n_221, n_178, n_386, n_287, n_344, n_473, n_422, n_475, n_72, n_104, n_41, n_415, n_56, n_141, n_485, n_355, n_486, n_15, n_336, n_145, n_48, n_50, n_337, n_430, n_313, n_88, n_479, n_216, n_168, n_395, n_164, n_432, n_311, n_208, n_142, n_214, n_328, n_140, n_299, n_303, n_369, n_296, n_241, n_357, n_184, n_446, n_445, n_65, n_78, n_144, n_114, n_96, n_165, n_468, n_213, n_129, n_342, n_482, n_98, n_361, n_464, n_363, n_402, n_413, n_197, n_107, n_69, n_236, n_388, n_1, n_249, n_304, n_329, n_203, n_274, n_384, n_460, n_80, n_35, n_73, n_277, n_92, n_19, n_338, n_149, n_477, n_461, n_333, n_309, n_30, n_14, n_84, n_462, n_130, n_322, n_258, n_29, n_79, n_151, n_25, n_306, n_458, n_288, n_188, n_190, n_201, n_263, n_471, n_44, n_224, n_40, n_34, n_228, n_283, n_383, n_474, n_112, n_85, n_463, n_488, n_239, n_466, n_420, n_55, n_49, n_310, n_54, n_12, n_465, n_76, n_358, n_362, n_170, n_332, n_27, n_77, n_102, n_161, n_273, n_349, n_270, n_230, n_81, n_118, n_279, n_70, n_253, n_261, n_174, n_289, n_172, n_206, n_217, n_440, n_478, n_441, n_450, n_312, n_476, n_429, n_345, n_210, n_365, n_91, n_176, n_182, n_143, n_83, n_354, n_480, n_237, n_425, n_407, n_180, n_340, n_207, n_37, n_346, n_393, n_229, n_108, n_487, n_437, n_66, n_177, n_60, n_403, n_453, n_421, n_16, n_0, n_58, n_405, n_18, n_359, n_117, n_326, n_233, n_404, n_205, n_366, n_113, n_246, n_179, n_125, n_410, n_269, n_128, n_285, n_412, n_120, n_232, n_327, n_135, n_126, n_202, n_266, n_272, n_427, n_193, n_251, n_352, n_53, n_160, n_426, n_409, n_154, n_62, n_148, n_71, n_300, n_435, n_159, n_334, n_391, n_434, n_175, n_262, n_238, n_99, n_411, n_414, n_319, n_364, n_20, n_121, n_242, n_360, n_36, n_200, n_162, n_64, n_222, n_28, n_89, n_438, n_115, n_324, n_416, n_199, n_187, n_32, n_401, n_103, n_348, n_97, n_166, n_11, n_424, n_7, n_256, n_305, n_52, n_278, n_110, n_1988);

input n_137;
input n_294;
input n_431;
input n_318;
input n_380;
input n_419;
input n_444;
input n_469;
input n_82;
input n_194;
input n_316;
input n_389;
input n_418;
input n_248;
input n_124;
input n_86;
input n_136;
input n_146;
input n_315;
input n_268;
input n_451;
input n_408;
input n_61;
input n_376;
input n_127;
input n_75;
input n_235;
input n_226;
input n_74;
input n_57;
input n_353;
input n_351;
input n_367;
input n_452;
input n_397;
input n_111;
input n_483;
input n_155;
input n_43;
input n_116;
input n_22;
input n_467;
input n_423;
input n_284;
input n_46;
input n_245;
input n_21;
input n_139;
input n_38;
input n_105;
input n_280;
input n_4;
input n_378;
input n_17;
input n_382;
input n_254;
input n_33;
input n_23;
input n_302;
input n_265;
input n_293;
input n_372;
input n_443;
input n_244;
input n_47;
input n_173;
input n_198;
input n_447;
input n_247;
input n_314;
input n_368;
input n_433;
input n_8;
input n_321;
input n_292;
input n_100;
input n_455;
input n_417;
input n_212;
input n_385;
input n_119;
input n_275;
input n_252;
input n_26;
input n_295;
input n_133;
input n_330;
input n_2;
input n_6;
input n_39;
input n_147;
input n_373;
input n_67;
input n_307;
input n_439;
input n_87;
input n_150;
input n_106;
input n_209;
input n_259;
input n_448;
input n_375;
input n_301;
input n_68;
input n_93;
input n_186;
input n_134;
input n_191;
input n_51;
input n_63;
input n_171;
input n_153;
input n_399;
input n_341;
input n_204;
input n_394;
input n_250;
input n_260;
input n_298;
input n_320;
input n_286;
input n_122;
input n_282;
input n_331;
input n_10;
input n_24;
input n_406;
input n_470;
input n_325;
input n_449;
input n_132;
input n_90;
input n_101;
input n_281;
input n_240;
input n_381;
input n_189;
input n_220;
input n_291;
input n_231;
input n_257;
input n_390;
input n_31;
input n_456;
input n_13;
input n_371;
input n_481;
input n_152;
input n_317;
input n_9;
input n_323;
input n_195;
input n_42;
input n_356;
input n_227;
input n_45;
input n_271;
input n_94;
input n_335;
input n_123;
input n_370;
input n_167;
input n_234;
input n_343;
input n_308;
input n_379;
input n_428;
input n_267;
input n_457;
input n_297;
input n_156;
input n_5;
input n_225;
input n_377;
input n_484;
input n_219;
input n_442;
input n_157;
input n_131;
input n_192;
input n_223;
input n_392;
input n_158;
input n_138;
input n_264;
input n_109;
input n_472;
input n_454;
input n_387;
input n_374;
input n_163;
input n_276;
input n_339;
input n_95;
input n_183;
input n_185;
input n_243;
input n_398;
input n_396;
input n_347;
input n_169;
input n_59;
input n_255;
input n_215;
input n_350;
input n_196;
input n_459;
input n_211;
input n_218;
input n_400;
input n_181;
input n_436;
input n_3;
input n_290;
input n_221;
input n_178;
input n_386;
input n_287;
input n_344;
input n_473;
input n_422;
input n_475;
input n_72;
input n_104;
input n_41;
input n_415;
input n_56;
input n_141;
input n_485;
input n_355;
input n_486;
input n_15;
input n_336;
input n_145;
input n_48;
input n_50;
input n_337;
input n_430;
input n_313;
input n_88;
input n_479;
input n_216;
input n_168;
input n_395;
input n_164;
input n_432;
input n_311;
input n_208;
input n_142;
input n_214;
input n_328;
input n_140;
input n_299;
input n_303;
input n_369;
input n_296;
input n_241;
input n_357;
input n_184;
input n_446;
input n_445;
input n_65;
input n_78;
input n_144;
input n_114;
input n_96;
input n_165;
input n_468;
input n_213;
input n_129;
input n_342;
input n_482;
input n_98;
input n_361;
input n_464;
input n_363;
input n_402;
input n_413;
input n_197;
input n_107;
input n_69;
input n_236;
input n_388;
input n_1;
input n_249;
input n_304;
input n_329;
input n_203;
input n_274;
input n_384;
input n_460;
input n_80;
input n_35;
input n_73;
input n_277;
input n_92;
input n_19;
input n_338;
input n_149;
input n_477;
input n_461;
input n_333;
input n_309;
input n_30;
input n_14;
input n_84;
input n_462;
input n_130;
input n_322;
input n_258;
input n_29;
input n_79;
input n_151;
input n_25;
input n_306;
input n_458;
input n_288;
input n_188;
input n_190;
input n_201;
input n_263;
input n_471;
input n_44;
input n_224;
input n_40;
input n_34;
input n_228;
input n_283;
input n_383;
input n_474;
input n_112;
input n_85;
input n_463;
input n_488;
input n_239;
input n_466;
input n_420;
input n_55;
input n_49;
input n_310;
input n_54;
input n_12;
input n_465;
input n_76;
input n_358;
input n_362;
input n_170;
input n_332;
input n_27;
input n_77;
input n_102;
input n_161;
input n_273;
input n_349;
input n_270;
input n_230;
input n_81;
input n_118;
input n_279;
input n_70;
input n_253;
input n_261;
input n_174;
input n_289;
input n_172;
input n_206;
input n_217;
input n_440;
input n_478;
input n_441;
input n_450;
input n_312;
input n_476;
input n_429;
input n_345;
input n_210;
input n_365;
input n_91;
input n_176;
input n_182;
input n_143;
input n_83;
input n_354;
input n_480;
input n_237;
input n_425;
input n_407;
input n_180;
input n_340;
input n_207;
input n_37;
input n_346;
input n_393;
input n_229;
input n_108;
input n_487;
input n_437;
input n_66;
input n_177;
input n_60;
input n_403;
input n_453;
input n_421;
input n_16;
input n_0;
input n_58;
input n_405;
input n_18;
input n_359;
input n_117;
input n_326;
input n_233;
input n_404;
input n_205;
input n_366;
input n_113;
input n_246;
input n_179;
input n_125;
input n_410;
input n_269;
input n_128;
input n_285;
input n_412;
input n_120;
input n_232;
input n_327;
input n_135;
input n_126;
input n_202;
input n_266;
input n_272;
input n_427;
input n_193;
input n_251;
input n_352;
input n_53;
input n_160;
input n_426;
input n_409;
input n_154;
input n_62;
input n_148;
input n_71;
input n_300;
input n_435;
input n_159;
input n_334;
input n_391;
input n_434;
input n_175;
input n_262;
input n_238;
input n_99;
input n_411;
input n_414;
input n_319;
input n_364;
input n_20;
input n_121;
input n_242;
input n_360;
input n_36;
input n_200;
input n_162;
input n_64;
input n_222;
input n_28;
input n_89;
input n_438;
input n_115;
input n_324;
input n_416;
input n_199;
input n_187;
input n_32;
input n_401;
input n_103;
input n_348;
input n_97;
input n_166;
input n_11;
input n_424;
input n_7;
input n_256;
input n_305;
input n_52;
input n_278;
input n_110;

output n_1988;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1729;
wire n_1166;
wire n_1751;
wire n_1508;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1859;
wire n_1677;
wire n_1150;
wire n_1780;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_1738;
wire n_1021;
wire n_1960;
wire n_551;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1695;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_1789;
wire n_1666;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_1545;
wire n_864;
wire n_859;
wire n_951;
wire n_1947;
wire n_1264;
wire n_1494;
wire n_625;
wire n_854;
wire n_1462;
wire n_1799;
wire n_1580;
wire n_674;
wire n_1939;
wire n_1806;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_1869;
wire n_1607;
wire n_1563;
wire n_606;
wire n_877;
wire n_1696;
wire n_755;
wire n_1118;
wire n_1686;
wire n_947;
wire n_1285;
wire n_1860;
wire n_1359;
wire n_530;
wire n_1107;
wire n_1728;
wire n_556;
wire n_1230;
wire n_668;
wire n_1896;
wire n_929;
wire n_1124;
wire n_1818;
wire n_902;
wire n_1576;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1705;
wire n_1257;
wire n_1182;
wire n_579;
wire n_1698;
wire n_1261;
wire n_938;
wire n_1098;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_519;
wire n_1016;
wire n_1243;
wire n_546;
wire n_1280;
wire n_1845;
wire n_731;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_1236;
wire n_1633;
wire n_569;
wire n_1778;
wire n_920;
wire n_1289;
wire n_1517;
wire n_1669;
wire n_976;
wire n_1949;
wire n_1449;
wire n_1946;
wire n_1566;
wire n_1078;
wire n_1670;
wire n_775;
wire n_600;
wire n_1484;
wire n_1374;
wire n_1328;
wire n_1948;
wire n_1984;
wire n_1877;
wire n_1831;
wire n_1598;
wire n_1723;
wire n_955;
wire n_1850;
wire n_1146;
wire n_882;
wire n_1097;
wire n_1036;
wire n_1749;
wire n_550;
wire n_696;
wire n_897;
wire n_798;
wire n_646;
wire n_1428;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_580;
wire n_1040;
wire n_1872;
wire n_1852;
wire n_578;
wire n_926;
wire n_1218;
wire n_1931;
wire n_1070;
wire n_777;
wire n_1547;
wire n_1030;
wire n_1755;
wire n_1071;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1801;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_663;
wire n_845;
wire n_1862;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_1796;
wire n_680;
wire n_1473;
wire n_1587;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_1748;
wire n_1672;
wire n_675;
wire n_888;
wire n_1880;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1384;
wire n_1556;
wire n_1863;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_1706;
wire n_1582;
wire n_1069;
wire n_1784;
wire n_1075;
wire n_1836;
wire n_1450;
wire n_1322;
wire n_1471;
wire n_1986;
wire n_1750;
wire n_1459;
wire n_889;
wire n_973;
wire n_1700;
wire n_571;
wire n_1585;
wire n_1971;
wire n_1599;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_1950;
wire n_907;
wire n_1447;
wire n_1377;
wire n_989;
wire n_1039;
wire n_1403;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_1667;
wire n_838;
wire n_1053;
wire n_1224;
wire n_1926;
wire n_1248;
wire n_1331;
wire n_953;
wire n_1014;
wire n_1241;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_793;
wire n_1819;
wire n_1527;
wire n_534;
wire n_1882;
wire n_884;
wire n_944;
wire n_1754;
wire n_1623;
wire n_1854;
wire n_1565;
wire n_1809;
wire n_1856;
wire n_647;
wire n_1072;
wire n_832;
wire n_857;
wire n_561;
wire n_1319;
wire n_1825;
wire n_1951;
wire n_1883;
wire n_1906;
wire n_1712;
wire n_1387;
wire n_1532;
wire n_1027;
wire n_971;
wire n_1156;
wire n_794;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1775;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_1709;
wire n_728;
wire n_1162;
wire n_1538;
wire n_1838;
wire n_1199;
wire n_1847;
wire n_1779;
wire n_1884;
wire n_1038;
wire n_520;
wire n_1369;
wire n_1841;
wire n_1660;
wire n_887;
wire n_1905;
wire n_809;
wire n_870;
wire n_931;
wire n_599;
wire n_1711;
wire n_1662;
wire n_1891;
wire n_1481;
wire n_1942;
wire n_1978;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_1629;
wire n_1293;
wire n_965;
wire n_1876;
wire n_1743;
wire n_935;
wire n_1175;
wire n_817;
wire n_1479;
wire n_1810;
wire n_1888;
wire n_759;
wire n_1892;
wire n_806;
wire n_1766;
wire n_1477;
wire n_1635;
wire n_1963;
wire n_1571;
wire n_1189;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_784;
wire n_1733;
wire n_1244;
wire n_1194;
wire n_1925;
wire n_1815;
wire n_851;
wire n_615;
wire n_1759;
wire n_843;
wire n_1788;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_1679;
wire n_776;
wire n_1798;
wire n_1790;
wire n_1415;
wire n_525;
wire n_1260;
wire n_1746;
wire n_1647;
wire n_1829;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_1674;
wire n_1833;
wire n_1830;
wire n_1710;
wire n_1128;
wire n_1734;
wire n_744;
wire n_590;
wire n_629;
wire n_1308;
wire n_1767;
wire n_1680;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_526;
wire n_1916;
wire n_677;
wire n_1333;
wire n_1121;
wire n_604;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_498;
wire n_1468;
wire n_1559;
wire n_1765;
wire n_1866;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_624;
wire n_1380;
wire n_1744;
wire n_1617;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_1839;
wire n_1837;
wire n_610;
wire n_1760;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_1832;
wire n_1851;
wire n_758;
wire n_999;
wire n_1933;
wire n_1656;
wire n_1158;
wire n_1509;
wire n_1874;
wire n_563;
wire n_1987;
wire n_1145;
wire n_878;
wire n_524;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_1871;
wire n_1964;
wire n_1163;
wire n_906;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_1781;
wire n_658;
wire n_1740;
wire n_1362;
wire n_1586;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_1923;
wire n_1773;
wire n_592;
wire n_1169;
wire n_1596;
wire n_1692;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_1095;
wire n_1828;
wire n_1614;
wire n_514;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_1431;
wire n_1593;
wire n_1033;
wire n_636;
wire n_660;
wire n_1640;
wire n_1732;
wire n_1009;
wire n_1148;
wire n_750;
wire n_742;
wire n_995;
wire n_1609;
wire n_1887;
wire n_1383;
wire n_1073;
wire n_662;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1920;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1721;
wire n_1959;
wire n_1758;
wire n_1574;
wire n_1921;
wire n_1309;
wire n_1878;
wire n_1426;
wire n_1043;
wire n_1800;
wire n_1548;
wire n_614;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_743;
wire n_613;
wire n_1119;
wire n_1240;
wire n_1820;
wire n_829;
wire n_1612;
wire n_1416;
wire n_1724;
wire n_700;
wire n_1237;
wire n_573;
wire n_1420;
wire n_1132;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1785;
wire n_1568;
wire n_1006;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_1870;
wire n_512;
wire n_1591;
wire n_1682;
wire n_1980;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1927;
wire n_1349;
wire n_1093;
wire n_1031;
wire n_609;
wire n_1041;
wire n_1265;
wire n_1909;
wire n_1562;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_1965;
wire n_630;
wire n_1902;
wire n_1941;
wire n_1913;
wire n_504;
wire n_1823;
wire n_511;
wire n_874;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_1875;
wire n_1982;
wire n_1304;
wire n_1324;
wire n_987;
wire n_1846;
wire n_1885;
wire n_1455;
wire n_767;
wire n_993;
wire n_1903;
wire n_1407;
wire n_1551;
wire n_545;
wire n_860;
wire n_1805;
wire n_1816;
wire n_948;
wire n_1217;
wire n_628;
wire n_1849;
wire n_729;
wire n_1131;
wire n_1084;
wire n_1961;
wire n_970;
wire n_1935;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_824;
wire n_1645;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_1684;
wire n_1717;
wire n_572;
wire n_815;
wire n_1795;
wire n_1821;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_1708;
wire n_1438;
wire n_1082;
wire n_1840;
wire n_589;
wire n_716;
wire n_1630;
wire n_562;
wire n_1436;
wire n_1691;
wire n_952;
wire n_1229;
wire n_701;
wire n_1437;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_1776;
wire n_531;
wire n_1757;
wire n_890;
wire n_1897;
wire n_764;
wire n_1919;
wire n_1056;
wire n_1424;
wire n_960;
wire n_1893;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_634;
wire n_1958;
wire n_1252;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_1311;
wire n_1519;
wire n_950;
wire n_1553;
wire n_1811;
wire n_1346;
wire n_1299;
wire n_1808;
wire n_1060;
wire n_1141;
wire n_912;
wire n_968;
wire n_619;
wire n_1386;
wire n_1699;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_885;
wire n_1432;
wire n_1357;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_1954;
wire n_1608;
wire n_983;
wire n_1844;
wire n_1305;
wire n_873;
wire n_1826;
wire n_1112;
wire n_762;
wire n_1283;
wire n_1644;
wire n_690;
wire n_1974;
wire n_583;
wire n_1343;
wire n_1203;
wire n_1631;
wire n_821;
wire n_1763;
wire n_1966;
wire n_1768;
wire n_1179;
wire n_753;
wire n_621;
wire n_1048;
wire n_1719;
wire n_1288;
wire n_507;
wire n_1560;
wire n_1605;
wire n_1228;
wire n_972;
wire n_692;
wire n_1953;
wire n_1938;
wire n_820;
wire n_1200;
wire n_1911;
wire n_1301;
wire n_1363;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_1967;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_1688;
wire n_945;
wire n_492;
wire n_1504;
wire n_943;
wire n_992;
wire n_1932;
wire n_543;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_1643;
wire n_883;
wire n_1983;
wire n_1594;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_856;
wire n_1793;
wire n_1976;
wire n_918;
wire n_942;
wire n_1804;
wire n_1147;
wire n_1557;
wire n_1977;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_894;
wire n_1636;
wire n_1730;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1865;
wire n_1470;
wire n_1096;
wire n_1575;
wire n_1735;
wire n_1697;
wire n_833;
wire n_1646;
wire n_1307;
wire n_1881;
wire n_988;
wire n_1940;
wire n_814;
wire n_1549;
wire n_1934;
wire n_1201;
wire n_1114;
wire n_655;
wire n_1616;
wire n_1446;
wire n_669;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_1807;
wire n_1149;
wire n_1671;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_1824;
wire n_1917;
wire n_1219;
wire n_1204;
wire n_1814;
wire n_1035;
wire n_555;
wire n_783;
wire n_1848;
wire n_1928;
wire n_1188;
wire n_1722;
wire n_661;
wire n_1802;
wire n_849;
wire n_681;
wire n_584;
wire n_1638;
wire n_1786;
wire n_510;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_875;
wire n_1110;
wire n_1655;
wire n_749;
wire n_1895;
wire n_1134;
wire n_1358;
wire n_717;
wire n_939;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_1338;
wire n_577;
wire n_1522;
wire n_1687;
wire n_1637;
wire n_1419;
wire n_1653;
wire n_693;
wire n_1506;
wire n_836;
wire n_990;
wire n_1886;
wire n_1389;
wire n_1894;
wire n_975;
wire n_1908;
wire n_1256;
wire n_1702;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_770;
wire n_1375;
wire n_1102;
wire n_1843;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1929;
wire n_1164;
wire n_1659;
wire n_1834;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_1572;
wire n_1968;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1736;
wire n_1685;
wire n_601;
wire n_917;
wire n_1714;
wire n_966;
wire n_1116;
wire n_1661;
wire n_1212;
wire n_1541;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_1731;
wire n_818;
wire n_1970;
wire n_861;
wire n_1713;
wire n_1183;
wire n_1658;
wire n_899;
wire n_1253;
wire n_1737;
wire n_1904;
wire n_774;
wire n_1628;
wire n_1335;
wire n_1514;
wire n_1777;
wire n_1957;
wire n_1059;
wire n_1345;
wire n_1133;
wire n_1771;
wire n_1912;
wire n_1899;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_1168;
wire n_707;
wire n_937;
wire n_1427;
wire n_1726;
wire n_665;
wire n_1835;
wire n_1584;
wire n_1440;
wire n_1853;
wire n_1356;
wire n_1787;
wire n_910;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1774;
wire n_1725;
wire n_1313;
wire n_1136;
wire n_1491;
wire n_754;
wire n_1496;
wire n_1125;
wire n_708;
wire n_529;
wire n_1812;
wire n_735;
wire n_1915;
wire n_1109;
wire n_895;
wire n_1310;
wire n_1803;
wire n_1399;
wire n_1543;
wire n_1979;
wire n_791;
wire n_732;
wire n_1533;
wire n_808;
wire n_797;
wire n_1025;
wire n_1930;
wire n_1955;
wire n_500;
wire n_1067;
wire n_1720;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1742;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_594;
wire n_1291;
wire n_1297;
wire n_1753;
wire n_1782;
wire n_1155;
wire n_1418;
wire n_1972;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_985;
wire n_1855;
wire n_869;
wire n_810;
wire n_827;
wire n_1703;
wire n_1352;
wire n_626;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_676;
wire n_653;
wire n_642;
wire n_1602;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_664;
wire n_503;
wire n_1372;
wire n_605;
wire n_1273;
wire n_1822;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_1783;
wire n_780;
wire n_998;
wire n_1454;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_1907;
wire n_501;
wire n_823;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_1985;
wire n_1898;
wire n_581;
wire n_554;
wire n_1625;
wire n_898;
wire n_1762;
wire n_1013;
wire n_1452;
wire n_718;
wire n_1120;
wire n_719;
wire n_1791;
wire n_1890;
wire n_1747;
wire n_714;
wire n_1817;
wire n_1683;
wire n_909;
wire n_1944;
wire n_1530;
wire n_1497;
wire n_997;
wire n_932;
wire n_612;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_1981;
wire n_508;
wire n_506;
wire n_1320;
wire n_1663;
wire n_737;
wire n_1718;
wire n_986;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1715;
wire n_1281;
wire n_1952;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_1889;
wire n_1792;
wire n_1564;
wire n_1868;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1922;
wire n_1376;
wire n_941;
wire n_981;
wire n_1569;
wire n_867;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_1238;
wire n_548;
wire n_812;
wire n_518;
wire n_505;
wire n_1772;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1861;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1901;
wire n_1900;
wire n_1620;
wire n_1330;
wire n_1867;
wire n_1945;
wire n_1675;
wire n_1924;
wire n_1727;
wire n_1554;
wire n_1745;
wire n_769;
wire n_1046;
wire n_934;
wire n_1618;
wire n_826;
wire n_1813;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_1341;
wire n_570;
wire n_1641;
wire n_1361;
wire n_1707;
wire n_853;
wire n_751;
wire n_1973;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_704;
wire n_787;
wire n_1770;
wire n_961;
wire n_1756;
wire n_771;
wire n_1716;
wire n_1225;
wire n_1520;
wire n_522;
wire n_1287;
wire n_1262;
wire n_930;
wire n_1873;
wire n_1411;
wire n_622;
wire n_1962;
wire n_1577;
wire n_1087;
wire n_994;
wire n_1701;
wire n_848;
wire n_1550;
wire n_1498;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1857;
wire n_1344;
wire n_631;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_1797;
wire n_1769;
wire n_839;
wire n_1210;
wire n_1364;
wire n_1250;
wire n_1842;
wire n_871;
wire n_685;
wire n_598;
wire n_928;
wire n_608;
wire n_1367;
wire n_1943;
wire n_1460;
wire n_772;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_1086;
wire n_796;
wire n_1858;
wire n_1619;
wire n_1502;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_903;
wire n_1525;
wire n_1752;
wire n_740;
wire n_1404;
wire n_1794;
wire n_1315;
wire n_1061;
wire n_1910;
wire n_1298;
wire n_1652;
wire n_1193;
wire n_1676;
wire n_1255;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_844;
wire n_852;
wire n_1487;
wire n_1864;
wire n_1028;
wire n_1601;
wire n_781;
wire n_542;
wire n_1546;
wire n_595;
wire n_502;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_1673;
wire n_1321;
wire n_1975;
wire n_1937;
wire n_585;
wire n_1739;
wire n_616;
wire n_1914;
wire n_745;
wire n_1654;
wire n_1103;
wire n_648;
wire n_1379;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_1761;
wire n_641;
wire n_730;
wire n_1325;
wire n_1595;
wire n_575;
wire n_795;
wire n_695;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_1936;
wire n_1956;
wire n_1642;
wire n_1130;
wire n_720;
wire n_1918;
wire n_1526;
wire n_863;
wire n_805;
wire n_1604;
wire n_1275;
wire n_1764;
wire n_712;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_1493;
wire n_657;
wire n_644;
wire n_1741;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_1621;
wire n_566;
wire n_565;
wire n_1448;
wire n_1507;
wire n_1398;
wire n_1879;
wire n_597;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_651;
wire n_1340;
wire n_811;
wire n_1558;
wire n_807;
wire n_835;
wire n_666;
wire n_1433;
wire n_1704;
wire n_1254;
wire n_1026;
wire n_1969;
wire n_1234;
wire n_1138;
wire n_927;
wire n_1089;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_1681;
wire n_1018;
wire n_1693;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_1180;
wire n_1827;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;

INVxp67_ASAP7_75t_L g489 ( 
.A(n_315),
.Y(n_489)
);

CKINVDCx5p33_ASAP7_75t_R g490 ( 
.A(n_375),
.Y(n_490)
);

BUFx3_ASAP7_75t_L g491 ( 
.A(n_426),
.Y(n_491)
);

CKINVDCx5p33_ASAP7_75t_R g492 ( 
.A(n_281),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_399),
.Y(n_493)
);

CKINVDCx20_ASAP7_75t_R g494 ( 
.A(n_220),
.Y(n_494)
);

CKINVDCx5p33_ASAP7_75t_R g495 ( 
.A(n_449),
.Y(n_495)
);

CKINVDCx5p33_ASAP7_75t_R g496 ( 
.A(n_471),
.Y(n_496)
);

CKINVDCx5p33_ASAP7_75t_R g497 ( 
.A(n_484),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_164),
.Y(n_498)
);

BUFx5_ASAP7_75t_L g499 ( 
.A(n_66),
.Y(n_499)
);

INVx2_ASAP7_75t_L g500 ( 
.A(n_354),
.Y(n_500)
);

BUFx6f_ASAP7_75t_L g501 ( 
.A(n_162),
.Y(n_501)
);

CKINVDCx5p33_ASAP7_75t_R g502 ( 
.A(n_339),
.Y(n_502)
);

INVx1_ASAP7_75t_SL g503 ( 
.A(n_226),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_17),
.Y(n_504)
);

CKINVDCx5p33_ASAP7_75t_R g505 ( 
.A(n_79),
.Y(n_505)
);

CKINVDCx5p33_ASAP7_75t_R g506 ( 
.A(n_61),
.Y(n_506)
);

INVx2_ASAP7_75t_L g507 ( 
.A(n_430),
.Y(n_507)
);

CKINVDCx20_ASAP7_75t_R g508 ( 
.A(n_347),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_178),
.Y(n_509)
);

INVx1_ASAP7_75t_SL g510 ( 
.A(n_166),
.Y(n_510)
);

CKINVDCx5p33_ASAP7_75t_R g511 ( 
.A(n_228),
.Y(n_511)
);

CKINVDCx5p33_ASAP7_75t_R g512 ( 
.A(n_480),
.Y(n_512)
);

CKINVDCx5p33_ASAP7_75t_R g513 ( 
.A(n_180),
.Y(n_513)
);

CKINVDCx5p33_ASAP7_75t_R g514 ( 
.A(n_483),
.Y(n_514)
);

CKINVDCx5p33_ASAP7_75t_R g515 ( 
.A(n_183),
.Y(n_515)
);

CKINVDCx5p33_ASAP7_75t_R g516 ( 
.A(n_235),
.Y(n_516)
);

CKINVDCx5p33_ASAP7_75t_R g517 ( 
.A(n_451),
.Y(n_517)
);

CKINVDCx5p33_ASAP7_75t_R g518 ( 
.A(n_169),
.Y(n_518)
);

CKINVDCx5p33_ASAP7_75t_R g519 ( 
.A(n_173),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_159),
.Y(n_520)
);

INVx1_ASAP7_75t_SL g521 ( 
.A(n_470),
.Y(n_521)
);

CKINVDCx5p33_ASAP7_75t_R g522 ( 
.A(n_42),
.Y(n_522)
);

CKINVDCx5p33_ASAP7_75t_R g523 ( 
.A(n_239),
.Y(n_523)
);

HB1xp67_ASAP7_75t_L g524 ( 
.A(n_422),
.Y(n_524)
);

CKINVDCx5p33_ASAP7_75t_R g525 ( 
.A(n_398),
.Y(n_525)
);

CKINVDCx5p33_ASAP7_75t_R g526 ( 
.A(n_302),
.Y(n_526)
);

CKINVDCx5p33_ASAP7_75t_R g527 ( 
.A(n_176),
.Y(n_527)
);

CKINVDCx5p33_ASAP7_75t_R g528 ( 
.A(n_444),
.Y(n_528)
);

CKINVDCx5p33_ASAP7_75t_R g529 ( 
.A(n_435),
.Y(n_529)
);

CKINVDCx5p33_ASAP7_75t_R g530 ( 
.A(n_3),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_487),
.Y(n_531)
);

CKINVDCx20_ASAP7_75t_R g532 ( 
.A(n_350),
.Y(n_532)
);

CKINVDCx5p33_ASAP7_75t_R g533 ( 
.A(n_79),
.Y(n_533)
);

CKINVDCx5p33_ASAP7_75t_R g534 ( 
.A(n_181),
.Y(n_534)
);

INVx2_ASAP7_75t_SL g535 ( 
.A(n_38),
.Y(n_535)
);

CKINVDCx5p33_ASAP7_75t_R g536 ( 
.A(n_200),
.Y(n_536)
);

CKINVDCx5p33_ASAP7_75t_R g537 ( 
.A(n_20),
.Y(n_537)
);

INVx2_ASAP7_75t_SL g538 ( 
.A(n_394),
.Y(n_538)
);

CKINVDCx5p33_ASAP7_75t_R g539 ( 
.A(n_39),
.Y(n_539)
);

BUFx6f_ASAP7_75t_L g540 ( 
.A(n_14),
.Y(n_540)
);

INVx2_ASAP7_75t_L g541 ( 
.A(n_482),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_336),
.Y(n_542)
);

CKINVDCx5p33_ASAP7_75t_R g543 ( 
.A(n_253),
.Y(n_543)
);

CKINVDCx5p33_ASAP7_75t_R g544 ( 
.A(n_2),
.Y(n_544)
);

BUFx2_ASAP7_75t_L g545 ( 
.A(n_230),
.Y(n_545)
);

CKINVDCx5p33_ASAP7_75t_R g546 ( 
.A(n_3),
.Y(n_546)
);

BUFx6f_ASAP7_75t_L g547 ( 
.A(n_456),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_176),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_254),
.Y(n_549)
);

CKINVDCx5p33_ASAP7_75t_R g550 ( 
.A(n_277),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_72),
.Y(n_551)
);

CKINVDCx5p33_ASAP7_75t_R g552 ( 
.A(n_244),
.Y(n_552)
);

CKINVDCx5p33_ASAP7_75t_R g553 ( 
.A(n_89),
.Y(n_553)
);

CKINVDCx5p33_ASAP7_75t_R g554 ( 
.A(n_464),
.Y(n_554)
);

CKINVDCx5p33_ASAP7_75t_R g555 ( 
.A(n_88),
.Y(n_555)
);

CKINVDCx20_ASAP7_75t_R g556 ( 
.A(n_227),
.Y(n_556)
);

CKINVDCx20_ASAP7_75t_R g557 ( 
.A(n_18),
.Y(n_557)
);

INVx2_ASAP7_75t_SL g558 ( 
.A(n_76),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_57),
.Y(n_559)
);

INVx2_ASAP7_75t_L g560 ( 
.A(n_294),
.Y(n_560)
);

BUFx5_ASAP7_75t_L g561 ( 
.A(n_81),
.Y(n_561)
);

CKINVDCx5p33_ASAP7_75t_R g562 ( 
.A(n_121),
.Y(n_562)
);

CKINVDCx5p33_ASAP7_75t_R g563 ( 
.A(n_46),
.Y(n_563)
);

CKINVDCx5p33_ASAP7_75t_R g564 ( 
.A(n_128),
.Y(n_564)
);

CKINVDCx5p33_ASAP7_75t_R g565 ( 
.A(n_340),
.Y(n_565)
);

CKINVDCx20_ASAP7_75t_R g566 ( 
.A(n_57),
.Y(n_566)
);

CKINVDCx5p33_ASAP7_75t_R g567 ( 
.A(n_186),
.Y(n_567)
);

CKINVDCx5p33_ASAP7_75t_R g568 ( 
.A(n_47),
.Y(n_568)
);

CKINVDCx5p33_ASAP7_75t_R g569 ( 
.A(n_369),
.Y(n_569)
);

CKINVDCx20_ASAP7_75t_R g570 ( 
.A(n_417),
.Y(n_570)
);

CKINVDCx5p33_ASAP7_75t_R g571 ( 
.A(n_131),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_154),
.Y(n_572)
);

INVx1_ASAP7_75t_SL g573 ( 
.A(n_365),
.Y(n_573)
);

CKINVDCx5p33_ASAP7_75t_R g574 ( 
.A(n_189),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_370),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_55),
.Y(n_576)
);

CKINVDCx5p33_ASAP7_75t_R g577 ( 
.A(n_382),
.Y(n_577)
);

INVx2_ASAP7_75t_SL g578 ( 
.A(n_306),
.Y(n_578)
);

CKINVDCx16_ASAP7_75t_R g579 ( 
.A(n_296),
.Y(n_579)
);

CKINVDCx5p33_ASAP7_75t_R g580 ( 
.A(n_330),
.Y(n_580)
);

CKINVDCx16_ASAP7_75t_R g581 ( 
.A(n_210),
.Y(n_581)
);

CKINVDCx5p33_ASAP7_75t_R g582 ( 
.A(n_224),
.Y(n_582)
);

CKINVDCx20_ASAP7_75t_R g583 ( 
.A(n_147),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_266),
.Y(n_584)
);

CKINVDCx20_ASAP7_75t_R g585 ( 
.A(n_320),
.Y(n_585)
);

INVx1_ASAP7_75t_SL g586 ( 
.A(n_65),
.Y(n_586)
);

BUFx10_ASAP7_75t_L g587 ( 
.A(n_160),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_74),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_469),
.Y(n_589)
);

INVx3_ASAP7_75t_L g590 ( 
.A(n_49),
.Y(n_590)
);

CKINVDCx5p33_ASAP7_75t_R g591 ( 
.A(n_127),
.Y(n_591)
);

CKINVDCx5p33_ASAP7_75t_R g592 ( 
.A(n_40),
.Y(n_592)
);

CKINVDCx20_ASAP7_75t_R g593 ( 
.A(n_290),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_357),
.Y(n_594)
);

CKINVDCx20_ASAP7_75t_R g595 ( 
.A(n_288),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_436),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_206),
.Y(n_597)
);

CKINVDCx5p33_ASAP7_75t_R g598 ( 
.A(n_207),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_181),
.Y(n_599)
);

CKINVDCx20_ASAP7_75t_R g600 ( 
.A(n_54),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_22),
.Y(n_601)
);

BUFx10_ASAP7_75t_L g602 ( 
.A(n_160),
.Y(n_602)
);

INVx2_ASAP7_75t_L g603 ( 
.A(n_207),
.Y(n_603)
);

INVx2_ASAP7_75t_L g604 ( 
.A(n_462),
.Y(n_604)
);

CKINVDCx5p33_ASAP7_75t_R g605 ( 
.A(n_393),
.Y(n_605)
);

CKINVDCx5p33_ASAP7_75t_R g606 ( 
.A(n_392),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_96),
.Y(n_607)
);

CKINVDCx5p33_ASAP7_75t_R g608 ( 
.A(n_26),
.Y(n_608)
);

CKINVDCx5p33_ASAP7_75t_R g609 ( 
.A(n_303),
.Y(n_609)
);

CKINVDCx5p33_ASAP7_75t_R g610 ( 
.A(n_317),
.Y(n_610)
);

CKINVDCx5p33_ASAP7_75t_R g611 ( 
.A(n_415),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_29),
.Y(n_612)
);

CKINVDCx5p33_ASAP7_75t_R g613 ( 
.A(n_318),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_103),
.Y(n_614)
);

CKINVDCx5p33_ASAP7_75t_R g615 ( 
.A(n_283),
.Y(n_615)
);

CKINVDCx20_ASAP7_75t_R g616 ( 
.A(n_150),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_1),
.Y(n_617)
);

BUFx2_ASAP7_75t_L g618 ( 
.A(n_366),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_250),
.Y(n_619)
);

INVx2_ASAP7_75t_L g620 ( 
.A(n_319),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_485),
.Y(n_621)
);

CKINVDCx20_ASAP7_75t_R g622 ( 
.A(n_292),
.Y(n_622)
);

INVx2_ASAP7_75t_SL g623 ( 
.A(n_84),
.Y(n_623)
);

INVx2_ASAP7_75t_L g624 ( 
.A(n_63),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_385),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_278),
.Y(n_626)
);

CKINVDCx5p33_ASAP7_75t_R g627 ( 
.A(n_169),
.Y(n_627)
);

CKINVDCx5p33_ASAP7_75t_R g628 ( 
.A(n_130),
.Y(n_628)
);

CKINVDCx5p33_ASAP7_75t_R g629 ( 
.A(n_178),
.Y(n_629)
);

BUFx10_ASAP7_75t_L g630 ( 
.A(n_44),
.Y(n_630)
);

CKINVDCx5p33_ASAP7_75t_R g631 ( 
.A(n_113),
.Y(n_631)
);

BUFx6f_ASAP7_75t_L g632 ( 
.A(n_177),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_437),
.Y(n_633)
);

CKINVDCx5p33_ASAP7_75t_R g634 ( 
.A(n_159),
.Y(n_634)
);

CKINVDCx20_ASAP7_75t_R g635 ( 
.A(n_384),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_387),
.Y(n_636)
);

CKINVDCx20_ASAP7_75t_R g637 ( 
.A(n_275),
.Y(n_637)
);

BUFx10_ASAP7_75t_L g638 ( 
.A(n_110),
.Y(n_638)
);

BUFx3_ASAP7_75t_L g639 ( 
.A(n_270),
.Y(n_639)
);

CKINVDCx5p33_ASAP7_75t_R g640 ( 
.A(n_106),
.Y(n_640)
);

CKINVDCx5p33_ASAP7_75t_R g641 ( 
.A(n_222),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_55),
.Y(n_642)
);

CKINVDCx20_ASAP7_75t_R g643 ( 
.A(n_133),
.Y(n_643)
);

CKINVDCx5p33_ASAP7_75t_R g644 ( 
.A(n_33),
.Y(n_644)
);

CKINVDCx5p33_ASAP7_75t_R g645 ( 
.A(n_237),
.Y(n_645)
);

CKINVDCx5p33_ASAP7_75t_R g646 ( 
.A(n_148),
.Y(n_646)
);

BUFx5_ASAP7_75t_L g647 ( 
.A(n_453),
.Y(n_647)
);

INVx1_ASAP7_75t_SL g648 ( 
.A(n_472),
.Y(n_648)
);

CKINVDCx5p33_ASAP7_75t_R g649 ( 
.A(n_179),
.Y(n_649)
);

CKINVDCx5p33_ASAP7_75t_R g650 ( 
.A(n_423),
.Y(n_650)
);

CKINVDCx5p33_ASAP7_75t_R g651 ( 
.A(n_165),
.Y(n_651)
);

CKINVDCx5p33_ASAP7_75t_R g652 ( 
.A(n_272),
.Y(n_652)
);

INVx2_ASAP7_75t_L g653 ( 
.A(n_133),
.Y(n_653)
);

CKINVDCx5p33_ASAP7_75t_R g654 ( 
.A(n_327),
.Y(n_654)
);

CKINVDCx5p33_ASAP7_75t_R g655 ( 
.A(n_211),
.Y(n_655)
);

CKINVDCx5p33_ASAP7_75t_R g656 ( 
.A(n_223),
.Y(n_656)
);

CKINVDCx5p33_ASAP7_75t_R g657 ( 
.A(n_220),
.Y(n_657)
);

CKINVDCx20_ASAP7_75t_R g658 ( 
.A(n_246),
.Y(n_658)
);

BUFx3_ASAP7_75t_L g659 ( 
.A(n_234),
.Y(n_659)
);

CKINVDCx5p33_ASAP7_75t_R g660 ( 
.A(n_221),
.Y(n_660)
);

CKINVDCx5p33_ASAP7_75t_R g661 ( 
.A(n_117),
.Y(n_661)
);

CKINVDCx5p33_ASAP7_75t_R g662 ( 
.A(n_460),
.Y(n_662)
);

HB1xp67_ASAP7_75t_L g663 ( 
.A(n_258),
.Y(n_663)
);

BUFx3_ASAP7_75t_L g664 ( 
.A(n_53),
.Y(n_664)
);

INVxp67_ASAP7_75t_L g665 ( 
.A(n_323),
.Y(n_665)
);

INVx2_ASAP7_75t_SL g666 ( 
.A(n_477),
.Y(n_666)
);

CKINVDCx5p33_ASAP7_75t_R g667 ( 
.A(n_468),
.Y(n_667)
);

CKINVDCx16_ASAP7_75t_R g668 ( 
.A(n_242),
.Y(n_668)
);

CKINVDCx5p33_ASAP7_75t_R g669 ( 
.A(n_88),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_499),
.Y(n_670)
);

CKINVDCx20_ASAP7_75t_R g671 ( 
.A(n_494),
.Y(n_671)
);

CKINVDCx16_ASAP7_75t_R g672 ( 
.A(n_581),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_499),
.Y(n_673)
);

CKINVDCx5p33_ASAP7_75t_R g674 ( 
.A(n_490),
.Y(n_674)
);

INVx2_ASAP7_75t_L g675 ( 
.A(n_499),
.Y(n_675)
);

HB1xp67_ASAP7_75t_L g676 ( 
.A(n_505),
.Y(n_676)
);

INVx2_ASAP7_75t_L g677 ( 
.A(n_499),
.Y(n_677)
);

CKINVDCx5p33_ASAP7_75t_R g678 ( 
.A(n_492),
.Y(n_678)
);

HB1xp67_ASAP7_75t_L g679 ( 
.A(n_506),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_499),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_499),
.Y(n_681)
);

CKINVDCx14_ASAP7_75t_R g682 ( 
.A(n_545),
.Y(n_682)
);

BUFx2_ASAP7_75t_L g683 ( 
.A(n_664),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_561),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_561),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_561),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_561),
.Y(n_687)
);

INVx2_ASAP7_75t_L g688 ( 
.A(n_561),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_561),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_664),
.Y(n_690)
);

CKINVDCx5p33_ASAP7_75t_R g691 ( 
.A(n_495),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_590),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_590),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_501),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_501),
.Y(n_695)
);

CKINVDCx20_ASAP7_75t_R g696 ( 
.A(n_557),
.Y(n_696)
);

INVxp67_ASAP7_75t_SL g697 ( 
.A(n_524),
.Y(n_697)
);

CKINVDCx5p33_ASAP7_75t_R g698 ( 
.A(n_496),
.Y(n_698)
);

INVxp67_ASAP7_75t_SL g699 ( 
.A(n_663),
.Y(n_699)
);

CKINVDCx14_ASAP7_75t_R g700 ( 
.A(n_618),
.Y(n_700)
);

CKINVDCx5p33_ASAP7_75t_R g701 ( 
.A(n_497),
.Y(n_701)
);

CKINVDCx16_ASAP7_75t_R g702 ( 
.A(n_579),
.Y(n_702)
);

CKINVDCx20_ASAP7_75t_R g703 ( 
.A(n_566),
.Y(n_703)
);

BUFx2_ASAP7_75t_L g704 ( 
.A(n_513),
.Y(n_704)
);

CKINVDCx5p33_ASAP7_75t_R g705 ( 
.A(n_502),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_540),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_540),
.Y(n_707)
);

BUFx6f_ASAP7_75t_L g708 ( 
.A(n_547),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_540),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_632),
.Y(n_710)
);

CKINVDCx20_ASAP7_75t_R g711 ( 
.A(n_583),
.Y(n_711)
);

INVxp33_ASAP7_75t_SL g712 ( 
.A(n_515),
.Y(n_712)
);

CKINVDCx5p33_ASAP7_75t_R g713 ( 
.A(n_511),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_632),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_632),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_632),
.Y(n_716)
);

INVx2_ASAP7_75t_L g717 ( 
.A(n_647),
.Y(n_717)
);

CKINVDCx16_ASAP7_75t_R g718 ( 
.A(n_668),
.Y(n_718)
);

CKINVDCx5p33_ASAP7_75t_R g719 ( 
.A(n_512),
.Y(n_719)
);

INVxp67_ASAP7_75t_L g720 ( 
.A(n_587),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_498),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_504),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_509),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_520),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_548),
.Y(n_725)
);

INVxp33_ASAP7_75t_SL g726 ( 
.A(n_518),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_551),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_559),
.Y(n_728)
);

CKINVDCx20_ASAP7_75t_R g729 ( 
.A(n_600),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_572),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_576),
.Y(n_731)
);

CKINVDCx20_ASAP7_75t_R g732 ( 
.A(n_616),
.Y(n_732)
);

CKINVDCx5p33_ASAP7_75t_R g733 ( 
.A(n_519),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_588),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_597),
.Y(n_735)
);

CKINVDCx5p33_ASAP7_75t_R g736 ( 
.A(n_514),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_599),
.Y(n_737)
);

CKINVDCx5p33_ASAP7_75t_R g738 ( 
.A(n_516),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_601),
.Y(n_739)
);

CKINVDCx5p33_ASAP7_75t_R g740 ( 
.A(n_517),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_607),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_612),
.Y(n_742)
);

BUFx6f_ASAP7_75t_L g743 ( 
.A(n_547),
.Y(n_743)
);

CKINVDCx5p33_ASAP7_75t_R g744 ( 
.A(n_523),
.Y(n_744)
);

CKINVDCx5p33_ASAP7_75t_R g745 ( 
.A(n_525),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_614),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_617),
.Y(n_747)
);

CKINVDCx5p33_ASAP7_75t_R g748 ( 
.A(n_526),
.Y(n_748)
);

HB1xp67_ASAP7_75t_L g749 ( 
.A(n_522),
.Y(n_749)
);

INVx2_ASAP7_75t_L g750 ( 
.A(n_647),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_642),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_491),
.Y(n_752)
);

INVx2_ASAP7_75t_L g753 ( 
.A(n_647),
.Y(n_753)
);

CKINVDCx5p33_ASAP7_75t_R g754 ( 
.A(n_528),
.Y(n_754)
);

CKINVDCx20_ASAP7_75t_R g755 ( 
.A(n_643),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_491),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_639),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_639),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_659),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_659),
.Y(n_760)
);

BUFx6f_ASAP7_75t_L g761 ( 
.A(n_708),
.Y(n_761)
);

INVx3_ASAP7_75t_L g762 ( 
.A(n_708),
.Y(n_762)
);

AND2x4_ASAP7_75t_L g763 ( 
.A(n_692),
.B(n_538),
.Y(n_763)
);

INVx2_ASAP7_75t_L g764 ( 
.A(n_708),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_694),
.Y(n_765)
);

HB1xp67_ASAP7_75t_L g766 ( 
.A(n_683),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_695),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_706),
.Y(n_768)
);

BUFx6f_ASAP7_75t_L g769 ( 
.A(n_708),
.Y(n_769)
);

BUFx6f_ASAP7_75t_L g770 ( 
.A(n_743),
.Y(n_770)
);

INVx5_ASAP7_75t_L g771 ( 
.A(n_743),
.Y(n_771)
);

OAI22xp5_ASAP7_75t_SL g772 ( 
.A1(n_682),
.A2(n_510),
.B1(n_586),
.B2(n_530),
.Y(n_772)
);

CKINVDCx5p33_ASAP7_75t_R g773 ( 
.A(n_674),
.Y(n_773)
);

OAI22xp5_ASAP7_75t_SL g774 ( 
.A1(n_682),
.A2(n_527),
.B1(n_534),
.B2(n_533),
.Y(n_774)
);

BUFx6f_ASAP7_75t_L g775 ( 
.A(n_743),
.Y(n_775)
);

INVx2_ASAP7_75t_L g776 ( 
.A(n_743),
.Y(n_776)
);

AND2x6_ASAP7_75t_L g777 ( 
.A(n_675),
.B(n_547),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_707),
.Y(n_778)
);

AND2x2_ASAP7_75t_L g779 ( 
.A(n_676),
.B(n_503),
.Y(n_779)
);

XOR2xp5_ASAP7_75t_L g780 ( 
.A(n_671),
.B(n_508),
.Y(n_780)
);

NOR2x1_ASAP7_75t_L g781 ( 
.A(n_709),
.B(n_493),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_L g782 ( 
.A(n_678),
.B(n_666),
.Y(n_782)
);

INVx6_ASAP7_75t_L g783 ( 
.A(n_702),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_691),
.B(n_578),
.Y(n_784)
);

AND2x4_ASAP7_75t_L g785 ( 
.A(n_693),
.B(n_500),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_SL g786 ( 
.A(n_718),
.B(n_535),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_710),
.Y(n_787)
);

INVx2_ASAP7_75t_L g788 ( 
.A(n_675),
.Y(n_788)
);

OAI22xp5_ASAP7_75t_SL g789 ( 
.A1(n_700),
.A2(n_536),
.B1(n_539),
.B2(n_537),
.Y(n_789)
);

CKINVDCx20_ASAP7_75t_R g790 ( 
.A(n_671),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_L g791 ( 
.A(n_698),
.B(n_507),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_714),
.Y(n_792)
);

INVx2_ASAP7_75t_L g793 ( 
.A(n_677),
.Y(n_793)
);

AND2x2_ASAP7_75t_L g794 ( 
.A(n_679),
.B(n_521),
.Y(n_794)
);

BUFx2_ASAP7_75t_L g795 ( 
.A(n_733),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_715),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_701),
.B(n_507),
.Y(n_797)
);

AND2x4_ASAP7_75t_L g798 ( 
.A(n_697),
.B(n_489),
.Y(n_798)
);

BUFx8_ASAP7_75t_SL g799 ( 
.A(n_696),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_L g800 ( 
.A(n_705),
.B(n_541),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_716),
.Y(n_801)
);

INVx2_ASAP7_75t_L g802 ( 
.A(n_677),
.Y(n_802)
);

INVx4_ASAP7_75t_L g803 ( 
.A(n_713),
.Y(n_803)
);

HB1xp67_ASAP7_75t_L g804 ( 
.A(n_749),
.Y(n_804)
);

AND2x4_ASAP7_75t_L g805 ( 
.A(n_752),
.B(n_541),
.Y(n_805)
);

INVx2_ASAP7_75t_L g806 ( 
.A(n_688),
.Y(n_806)
);

NOR2xp33_ASAP7_75t_L g807 ( 
.A(n_699),
.B(n_712),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_L g808 ( 
.A(n_719),
.B(n_560),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_670),
.Y(n_809)
);

OA21x2_ASAP7_75t_L g810 ( 
.A1(n_673),
.A2(n_604),
.B(n_560),
.Y(n_810)
);

OAI22xp5_ASAP7_75t_L g811 ( 
.A1(n_700),
.A2(n_544),
.B1(n_553),
.B2(n_546),
.Y(n_811)
);

AND2x2_ASAP7_75t_SL g812 ( 
.A(n_672),
.B(n_604),
.Y(n_812)
);

HB1xp67_ASAP7_75t_L g813 ( 
.A(n_733),
.Y(n_813)
);

OAI22xp5_ASAP7_75t_SL g814 ( 
.A1(n_696),
.A2(n_562),
.B1(n_563),
.B2(n_555),
.Y(n_814)
);

INVx3_ASAP7_75t_L g815 ( 
.A(n_688),
.Y(n_815)
);

AND2x4_ASAP7_75t_L g816 ( 
.A(n_756),
.B(n_620),
.Y(n_816)
);

INVx2_ASAP7_75t_L g817 ( 
.A(n_680),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_788),
.Y(n_818)
);

AOI21x1_ASAP7_75t_L g819 ( 
.A1(n_809),
.A2(n_684),
.B(n_681),
.Y(n_819)
);

NOR2xp33_ASAP7_75t_L g820 ( 
.A(n_791),
.B(n_736),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_788),
.Y(n_821)
);

INVx2_ASAP7_75t_L g822 ( 
.A(n_793),
.Y(n_822)
);

INVx2_ASAP7_75t_L g823 ( 
.A(n_793),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_L g824 ( 
.A(n_797),
.B(n_738),
.Y(n_824)
);

INVx2_ASAP7_75t_L g825 ( 
.A(n_802),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_802),
.Y(n_826)
);

INVx2_ASAP7_75t_L g827 ( 
.A(n_806),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_SL g828 ( 
.A(n_779),
.B(n_740),
.Y(n_828)
);

AOI21x1_ASAP7_75t_L g829 ( 
.A1(n_810),
.A2(n_817),
.B(n_806),
.Y(n_829)
);

BUFx10_ASAP7_75t_L g830 ( 
.A(n_807),
.Y(n_830)
);

INVx2_ASAP7_75t_L g831 ( 
.A(n_815),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_817),
.Y(n_832)
);

INVx2_ASAP7_75t_L g833 ( 
.A(n_764),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_765),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_SL g835 ( 
.A(n_794),
.B(n_744),
.Y(n_835)
);

NOR2x1p5_ASAP7_75t_L g836 ( 
.A(n_803),
.B(n_603),
.Y(n_836)
);

NOR2xp33_ASAP7_75t_L g837 ( 
.A(n_800),
.B(n_745),
.Y(n_837)
);

NOR2xp33_ASAP7_75t_L g838 ( 
.A(n_808),
.B(n_748),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_L g839 ( 
.A(n_782),
.B(n_784),
.Y(n_839)
);

INVx2_ASAP7_75t_L g840 ( 
.A(n_764),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_767),
.Y(n_841)
);

INVx2_ASAP7_75t_L g842 ( 
.A(n_776),
.Y(n_842)
);

INVx2_ASAP7_75t_L g843 ( 
.A(n_776),
.Y(n_843)
);

INVx2_ASAP7_75t_L g844 ( 
.A(n_761),
.Y(n_844)
);

NOR2xp33_ASAP7_75t_L g845 ( 
.A(n_807),
.B(n_754),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_L g846 ( 
.A(n_798),
.B(n_685),
.Y(n_846)
);

INVx2_ASAP7_75t_L g847 ( 
.A(n_761),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_768),
.Y(n_848)
);

INVx2_ASAP7_75t_L g849 ( 
.A(n_761),
.Y(n_849)
);

AND2x2_ASAP7_75t_L g850 ( 
.A(n_805),
.B(n_757),
.Y(n_850)
);

INVx2_ASAP7_75t_L g851 ( 
.A(n_761),
.Y(n_851)
);

INVx2_ASAP7_75t_L g852 ( 
.A(n_769),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_SL g853 ( 
.A(n_812),
.B(n_712),
.Y(n_853)
);

INVx2_ASAP7_75t_L g854 ( 
.A(n_769),
.Y(n_854)
);

INVx2_ASAP7_75t_L g855 ( 
.A(n_769),
.Y(n_855)
);

INVx3_ASAP7_75t_L g856 ( 
.A(n_769),
.Y(n_856)
);

INVx8_ASAP7_75t_L g857 ( 
.A(n_777),
.Y(n_857)
);

NOR2xp33_ASAP7_75t_L g858 ( 
.A(n_803),
.B(n_726),
.Y(n_858)
);

OR2x2_ASAP7_75t_L g859 ( 
.A(n_766),
.B(n_704),
.Y(n_859)
);

INVx2_ASAP7_75t_L g860 ( 
.A(n_770),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_778),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_798),
.B(n_686),
.Y(n_862)
);

BUFx3_ASAP7_75t_L g863 ( 
.A(n_762),
.Y(n_863)
);

INVx2_ASAP7_75t_SL g864 ( 
.A(n_766),
.Y(n_864)
);

INVx2_ASAP7_75t_L g865 ( 
.A(n_770),
.Y(n_865)
);

INVx2_ASAP7_75t_L g866 ( 
.A(n_770),
.Y(n_866)
);

NAND2xp33_ASAP7_75t_L g867 ( 
.A(n_777),
.B(n_647),
.Y(n_867)
);

INVxp67_ASAP7_75t_SL g868 ( 
.A(n_762),
.Y(n_868)
);

INVx2_ASAP7_75t_L g869 ( 
.A(n_770),
.Y(n_869)
);

INVxp33_ASAP7_75t_L g870 ( 
.A(n_780),
.Y(n_870)
);

INVx2_ASAP7_75t_L g871 ( 
.A(n_775),
.Y(n_871)
);

INVx4_ASAP7_75t_L g872 ( 
.A(n_771),
.Y(n_872)
);

NAND3xp33_ASAP7_75t_L g873 ( 
.A(n_816),
.B(n_689),
.C(n_687),
.Y(n_873)
);

BUFx6f_ASAP7_75t_SL g874 ( 
.A(n_812),
.Y(n_874)
);

INVx2_ASAP7_75t_SL g875 ( 
.A(n_804),
.Y(n_875)
);

NOR2xp33_ASAP7_75t_L g876 ( 
.A(n_786),
.B(n_726),
.Y(n_876)
);

BUFx10_ASAP7_75t_L g877 ( 
.A(n_773),
.Y(n_877)
);

INVx2_ASAP7_75t_L g878 ( 
.A(n_775),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_787),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_792),
.Y(n_880)
);

INVx2_ASAP7_75t_L g881 ( 
.A(n_775),
.Y(n_881)
);

INVx3_ASAP7_75t_L g882 ( 
.A(n_771),
.Y(n_882)
);

OR2x2_ASAP7_75t_L g883 ( 
.A(n_811),
.B(n_720),
.Y(n_883)
);

INVx2_ASAP7_75t_L g884 ( 
.A(n_810),
.Y(n_884)
);

INVx3_ASAP7_75t_L g885 ( 
.A(n_771),
.Y(n_885)
);

AND2x2_ASAP7_75t_L g886 ( 
.A(n_805),
.B(n_758),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_796),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_801),
.Y(n_888)
);

INVx2_ASAP7_75t_L g889 ( 
.A(n_810),
.Y(n_889)
);

INVx2_ASAP7_75t_L g890 ( 
.A(n_771),
.Y(n_890)
);

BUFx10_ASAP7_75t_L g891 ( 
.A(n_783),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_816),
.Y(n_892)
);

INVx2_ASAP7_75t_L g893 ( 
.A(n_816),
.Y(n_893)
);

INVx2_ASAP7_75t_L g894 ( 
.A(n_805),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_785),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_SL g896 ( 
.A(n_772),
.B(n_532),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_893),
.Y(n_897)
);

NOR2xp33_ASAP7_75t_L g898 ( 
.A(n_839),
.B(n_813),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_L g899 ( 
.A(n_884),
.B(n_763),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_894),
.Y(n_900)
);

NAND2x1p5_ASAP7_75t_L g901 ( 
.A(n_892),
.B(n_895),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_892),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_L g903 ( 
.A(n_884),
.B(n_763),
.Y(n_903)
);

AND2x2_ASAP7_75t_L g904 ( 
.A(n_875),
.B(n_813),
.Y(n_904)
);

INVx2_ASAP7_75t_SL g905 ( 
.A(n_836),
.Y(n_905)
);

XNOR2xp5_ASAP7_75t_L g906 ( 
.A(n_870),
.B(n_790),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_834),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_841),
.Y(n_908)
);

NAND2xp33_ASAP7_75t_SL g909 ( 
.A(n_874),
.B(n_774),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_841),
.Y(n_910)
);

XOR2xp5_ASAP7_75t_L g911 ( 
.A(n_896),
.B(n_790),
.Y(n_911)
);

CKINVDCx20_ASAP7_75t_R g912 ( 
.A(n_877),
.Y(n_912)
);

INVxp67_ASAP7_75t_L g913 ( 
.A(n_875),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_L g914 ( 
.A(n_889),
.B(n_763),
.Y(n_914)
);

OAI21xp5_ASAP7_75t_L g915 ( 
.A1(n_889),
.A2(n_786),
.B(n_804),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_848),
.Y(n_916)
);

NOR2xp33_ASAP7_75t_L g917 ( 
.A(n_845),
.B(n_795),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_848),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_861),
.Y(n_919)
);

CKINVDCx20_ASAP7_75t_R g920 ( 
.A(n_877),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_879),
.Y(n_921)
);

NOR2xp33_ASAP7_75t_L g922 ( 
.A(n_820),
.B(n_783),
.Y(n_922)
);

INVx2_ASAP7_75t_L g923 ( 
.A(n_831),
.Y(n_923)
);

AND2x2_ASAP7_75t_L g924 ( 
.A(n_864),
.B(n_783),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_879),
.Y(n_925)
);

INVx2_ASAP7_75t_SL g926 ( 
.A(n_836),
.Y(n_926)
);

AND2x4_ASAP7_75t_L g927 ( 
.A(n_895),
.B(n_721),
.Y(n_927)
);

INVx2_ASAP7_75t_SL g928 ( 
.A(n_864),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_880),
.Y(n_929)
);

XOR2xp5_ASAP7_75t_L g930 ( 
.A(n_859),
.B(n_703),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_880),
.Y(n_931)
);

OAI21xp5_ASAP7_75t_L g932 ( 
.A1(n_829),
.A2(n_665),
.B(n_785),
.Y(n_932)
);

AND2x2_ASAP7_75t_L g933 ( 
.A(n_830),
.B(n_759),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_887),
.Y(n_934)
);

NOR2xp33_ASAP7_75t_R g935 ( 
.A(n_891),
.B(n_703),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_888),
.Y(n_936)
);

NOR2xp33_ASAP7_75t_L g937 ( 
.A(n_837),
.B(n_789),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_L g938 ( 
.A(n_832),
.B(n_717),
.Y(n_938)
);

OAI21xp5_ASAP7_75t_L g939 ( 
.A1(n_829),
.A2(n_781),
.B(n_542),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_850),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_886),
.Y(n_941)
);

XNOR2xp5_ASAP7_75t_L g942 ( 
.A(n_853),
.B(n_711),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_886),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_L g944 ( 
.A(n_846),
.B(n_862),
.Y(n_944)
);

INVx1_ASAP7_75t_L g945 ( 
.A(n_833),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_833),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_L g947 ( 
.A(n_838),
.B(n_717),
.Y(n_947)
);

NOR2xp33_ASAP7_75t_L g948 ( 
.A(n_824),
.B(n_828),
.Y(n_948)
);

AND2x2_ASAP7_75t_L g949 ( 
.A(n_830),
.B(n_760),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_840),
.Y(n_950)
);

INVx2_ASAP7_75t_L g951 ( 
.A(n_822),
.Y(n_951)
);

NAND2xp33_ASAP7_75t_SL g952 ( 
.A(n_874),
.B(n_556),
.Y(n_952)
);

AND2x2_ASAP7_75t_L g953 ( 
.A(n_830),
.B(n_690),
.Y(n_953)
);

AND2x2_ASAP7_75t_L g954 ( 
.A(n_876),
.B(n_722),
.Y(n_954)
);

INVx1_ASAP7_75t_L g955 ( 
.A(n_842),
.Y(n_955)
);

INVx1_ASAP7_75t_SL g956 ( 
.A(n_859),
.Y(n_956)
);

AND2x2_ASAP7_75t_L g957 ( 
.A(n_891),
.B(n_723),
.Y(n_957)
);

INVx1_ASAP7_75t_L g958 ( 
.A(n_843),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_843),
.Y(n_959)
);

OR2x6_ASAP7_75t_L g960 ( 
.A(n_883),
.B(n_814),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_L g961 ( 
.A(n_818),
.B(n_750),
.Y(n_961)
);

XNOR2xp5_ASAP7_75t_L g962 ( 
.A(n_835),
.B(n_711),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_868),
.Y(n_963)
);

INVx2_ASAP7_75t_L g964 ( 
.A(n_823),
.Y(n_964)
);

INVx1_ASAP7_75t_L g965 ( 
.A(n_818),
.Y(n_965)
);

INVx2_ASAP7_75t_L g966 ( 
.A(n_823),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_821),
.Y(n_967)
);

NOR2xp67_ASAP7_75t_L g968 ( 
.A(n_858),
.B(n_742),
.Y(n_968)
);

AND2x2_ASAP7_75t_L g969 ( 
.A(n_891),
.B(n_724),
.Y(n_969)
);

BUFx2_ASAP7_75t_L g970 ( 
.A(n_883),
.Y(n_970)
);

AND2x2_ASAP7_75t_L g971 ( 
.A(n_877),
.B(n_725),
.Y(n_971)
);

NAND2xp33_ASAP7_75t_R g972 ( 
.A(n_874),
.B(n_529),
.Y(n_972)
);

INVx1_ASAP7_75t_L g973 ( 
.A(n_821),
.Y(n_973)
);

INVx2_ASAP7_75t_L g974 ( 
.A(n_825),
.Y(n_974)
);

OR2x2_ASAP7_75t_L g975 ( 
.A(n_873),
.B(n_751),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_L g976 ( 
.A(n_826),
.B(n_750),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_826),
.Y(n_977)
);

AND2x6_ASAP7_75t_L g978 ( 
.A(n_825),
.B(n_620),
.Y(n_978)
);

CKINVDCx5p33_ASAP7_75t_R g979 ( 
.A(n_877),
.Y(n_979)
);

CKINVDCx5p33_ASAP7_75t_R g980 ( 
.A(n_863),
.Y(n_980)
);

XOR2xp5_ASAP7_75t_L g981 ( 
.A(n_873),
.B(n_729),
.Y(n_981)
);

AOI21x1_ASAP7_75t_L g982 ( 
.A1(n_819),
.A2(n_753),
.B(n_549),
.Y(n_982)
);

INVx1_ASAP7_75t_L g983 ( 
.A(n_863),
.Y(n_983)
);

AND2x4_ASAP7_75t_L g984 ( 
.A(n_844),
.B(n_727),
.Y(n_984)
);

NOR2xp67_ASAP7_75t_L g985 ( 
.A(n_827),
.B(n_728),
.Y(n_985)
);

AND2x2_ASAP7_75t_L g986 ( 
.A(n_819),
.B(n_730),
.Y(n_986)
);

NOR2xp33_ASAP7_75t_L g987 ( 
.A(n_856),
.B(n_729),
.Y(n_987)
);

OR2x2_ASAP7_75t_L g988 ( 
.A(n_844),
.B(n_734),
.Y(n_988)
);

INVx1_ASAP7_75t_L g989 ( 
.A(n_847),
.Y(n_989)
);

INVx3_ASAP7_75t_L g990 ( 
.A(n_849),
.Y(n_990)
);

OR2x2_ASAP7_75t_L g991 ( 
.A(n_849),
.B(n_735),
.Y(n_991)
);

INVx1_ASAP7_75t_L g992 ( 
.A(n_851),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_851),
.Y(n_993)
);

XOR2xp5_ASAP7_75t_L g994 ( 
.A(n_852),
.B(n_732),
.Y(n_994)
);

NAND2x1p5_ASAP7_75t_L g995 ( 
.A(n_856),
.B(n_531),
.Y(n_995)
);

INVx1_ASAP7_75t_L g996 ( 
.A(n_852),
.Y(n_996)
);

INVxp33_ASAP7_75t_L g997 ( 
.A(n_854),
.Y(n_997)
);

INVx1_ASAP7_75t_L g998 ( 
.A(n_854),
.Y(n_998)
);

INVx1_ASAP7_75t_SL g999 ( 
.A(n_867),
.Y(n_999)
);

INVxp33_ASAP7_75t_L g1000 ( 
.A(n_855),
.Y(n_1000)
);

INVx1_ASAP7_75t_L g1001 ( 
.A(n_855),
.Y(n_1001)
);

XOR2xp5_ASAP7_75t_L g1002 ( 
.A(n_860),
.B(n_755),
.Y(n_1002)
);

AND2x2_ASAP7_75t_L g1003 ( 
.A(n_860),
.B(n_731),
.Y(n_1003)
);

INVx2_ASAP7_75t_L g1004 ( 
.A(n_865),
.Y(n_1004)
);

INVx2_ASAP7_75t_SL g1005 ( 
.A(n_928),
.Y(n_1005)
);

INVx2_ASAP7_75t_SL g1006 ( 
.A(n_924),
.Y(n_1006)
);

INVx2_ASAP7_75t_SL g1007 ( 
.A(n_904),
.Y(n_1007)
);

AND2x6_ASAP7_75t_SL g1008 ( 
.A(n_937),
.B(n_799),
.Y(n_1008)
);

OR2x6_ASAP7_75t_L g1009 ( 
.A(n_913),
.B(n_857),
.Y(n_1009)
);

AOI22xp5_ASAP7_75t_L g1010 ( 
.A1(n_948),
.A2(n_570),
.B1(n_593),
.B2(n_585),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_L g1011 ( 
.A(n_944),
.B(n_866),
.Y(n_1011)
);

INVx8_ASAP7_75t_L g1012 ( 
.A(n_980),
.Y(n_1012)
);

AOI22xp5_ASAP7_75t_L g1013 ( 
.A1(n_898),
.A2(n_595),
.B1(n_635),
.B2(n_622),
.Y(n_1013)
);

NOR2xp67_ASAP7_75t_L g1014 ( 
.A(n_979),
.B(n_737),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_L g1015 ( 
.A(n_947),
.B(n_954),
.Y(n_1015)
);

OAI22xp5_ASAP7_75t_SL g1016 ( 
.A1(n_911),
.A2(n_755),
.B1(n_658),
.B2(n_637),
.Y(n_1016)
);

AOI22xp33_ASAP7_75t_L g1017 ( 
.A1(n_986),
.A2(n_902),
.B1(n_903),
.B2(n_899),
.Y(n_1017)
);

INVx3_ASAP7_75t_L g1018 ( 
.A(n_990),
.Y(n_1018)
);

AOI22xp33_ASAP7_75t_L g1019 ( 
.A1(n_899),
.A2(n_584),
.B1(n_589),
.B2(n_575),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_SL g1020 ( 
.A(n_913),
.B(n_573),
.Y(n_1020)
);

AOI22xp5_ASAP7_75t_L g1021 ( 
.A1(n_999),
.A2(n_866),
.B1(n_871),
.B2(n_869),
.Y(n_1021)
);

OAI22xp5_ASAP7_75t_L g1022 ( 
.A1(n_999),
.A2(n_648),
.B1(n_594),
.B2(n_596),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_L g1023 ( 
.A(n_947),
.B(n_869),
.Y(n_1023)
);

INVx2_ASAP7_75t_SL g1024 ( 
.A(n_971),
.Y(n_1024)
);

NOR2xp33_ASAP7_75t_L g1025 ( 
.A(n_917),
.B(n_799),
.Y(n_1025)
);

NAND2xp33_ASAP7_75t_L g1026 ( 
.A(n_903),
.B(n_914),
.Y(n_1026)
);

NOR2xp33_ASAP7_75t_L g1027 ( 
.A(n_922),
.B(n_564),
.Y(n_1027)
);

HB1xp67_ASAP7_75t_L g1028 ( 
.A(n_956),
.Y(n_1028)
);

AND2x2_ASAP7_75t_L g1029 ( 
.A(n_953),
.B(n_587),
.Y(n_1029)
);

INVx3_ASAP7_75t_L g1030 ( 
.A(n_990),
.Y(n_1030)
);

NOR2xp33_ASAP7_75t_L g1031 ( 
.A(n_956),
.B(n_567),
.Y(n_1031)
);

NOR2xp33_ASAP7_75t_L g1032 ( 
.A(n_970),
.B(n_933),
.Y(n_1032)
);

NAND2xp5_ASAP7_75t_L g1033 ( 
.A(n_907),
.B(n_908),
.Y(n_1033)
);

AND2x6_ASAP7_75t_SL g1034 ( 
.A(n_960),
.B(n_739),
.Y(n_1034)
);

NAND2xp5_ASAP7_75t_L g1035 ( 
.A(n_910),
.B(n_878),
.Y(n_1035)
);

AOI22xp5_ASAP7_75t_L g1036 ( 
.A1(n_968),
.A2(n_881),
.B1(n_878),
.B2(n_619),
.Y(n_1036)
);

INVx1_ASAP7_75t_L g1037 ( 
.A(n_900),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_SL g1038 ( 
.A(n_915),
.B(n_543),
.Y(n_1038)
);

NAND2xp5_ASAP7_75t_SL g1039 ( 
.A(n_957),
.B(n_550),
.Y(n_1039)
);

INVx2_ASAP7_75t_L g1040 ( 
.A(n_951),
.Y(n_1040)
);

BUFx6f_ASAP7_75t_L g1041 ( 
.A(n_901),
.Y(n_1041)
);

AOI22xp33_ASAP7_75t_L g1042 ( 
.A1(n_914),
.A2(n_625),
.B1(n_626),
.B2(n_621),
.Y(n_1042)
);

NAND2xp5_ASAP7_75t_L g1043 ( 
.A(n_916),
.B(n_633),
.Y(n_1043)
);

OR2x6_ASAP7_75t_L g1044 ( 
.A(n_905),
.B(n_857),
.Y(n_1044)
);

NOR2xp33_ASAP7_75t_L g1045 ( 
.A(n_949),
.B(n_568),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_L g1046 ( 
.A(n_918),
.B(n_636),
.Y(n_1046)
);

NAND3xp33_ASAP7_75t_L g1047 ( 
.A(n_987),
.B(n_574),
.C(n_571),
.Y(n_1047)
);

INVx1_ASAP7_75t_L g1048 ( 
.A(n_965),
.Y(n_1048)
);

AND2x2_ASAP7_75t_L g1049 ( 
.A(n_969),
.B(n_602),
.Y(n_1049)
);

NAND2xp5_ASAP7_75t_SL g1050 ( 
.A(n_926),
.B(n_552),
.Y(n_1050)
);

NAND3xp33_ASAP7_75t_L g1051 ( 
.A(n_942),
.B(n_592),
.C(n_591),
.Y(n_1051)
);

BUFx3_ASAP7_75t_L g1052 ( 
.A(n_912),
.Y(n_1052)
);

NAND2xp5_ASAP7_75t_SL g1053 ( 
.A(n_919),
.B(n_554),
.Y(n_1053)
);

AOI22xp33_ASAP7_75t_L g1054 ( 
.A1(n_940),
.A2(n_943),
.B1(n_941),
.B2(n_921),
.Y(n_1054)
);

AND2x2_ASAP7_75t_L g1055 ( 
.A(n_927),
.B(n_602),
.Y(n_1055)
);

CKINVDCx5p33_ASAP7_75t_R g1056 ( 
.A(n_935),
.Y(n_1056)
);

AOI22xp33_ASAP7_75t_L g1057 ( 
.A1(n_925),
.A2(n_647),
.B1(n_547),
.B2(n_857),
.Y(n_1057)
);

OAI221xp5_ASAP7_75t_L g1058 ( 
.A1(n_929),
.A2(n_623),
.B1(n_558),
.B2(n_598),
.C(n_608),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_967),
.Y(n_1059)
);

O2A1O1Ixp33_ASAP7_75t_L g1060 ( 
.A1(n_975),
.A2(n_603),
.B(n_653),
.C(n_624),
.Y(n_1060)
);

NAND2xp5_ASAP7_75t_L g1061 ( 
.A(n_931),
.B(n_565),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_L g1062 ( 
.A(n_934),
.B(n_569),
.Y(n_1062)
);

INVx2_ASAP7_75t_SL g1063 ( 
.A(n_988),
.Y(n_1063)
);

AND2x2_ASAP7_75t_L g1064 ( 
.A(n_927),
.B(n_630),
.Y(n_1064)
);

INVx1_ASAP7_75t_L g1065 ( 
.A(n_973),
.Y(n_1065)
);

NAND2xp5_ASAP7_75t_L g1066 ( 
.A(n_936),
.B(n_577),
.Y(n_1066)
);

AOI21xp5_ASAP7_75t_L g1067 ( 
.A1(n_932),
.A2(n_857),
.B(n_882),
.Y(n_1067)
);

INVx1_ASAP7_75t_L g1068 ( 
.A(n_977),
.Y(n_1068)
);

BUFx6f_ASAP7_75t_SL g1069 ( 
.A(n_960),
.Y(n_1069)
);

NAND2xp5_ASAP7_75t_L g1070 ( 
.A(n_963),
.B(n_580),
.Y(n_1070)
);

NOR2xp67_ASAP7_75t_SL g1071 ( 
.A(n_983),
.B(n_653),
.Y(n_1071)
);

OAI22xp5_ASAP7_75t_L g1072 ( 
.A1(n_901),
.A2(n_857),
.B1(n_582),
.B2(n_605),
.Y(n_1072)
);

BUFx4_ASAP7_75t_L g1073 ( 
.A(n_920),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_SL g1074 ( 
.A(n_984),
.B(n_606),
.Y(n_1074)
);

NOR2xp67_ASAP7_75t_L g1075 ( 
.A(n_923),
.B(n_225),
.Y(n_1075)
);

NAND2xp5_ASAP7_75t_SL g1076 ( 
.A(n_984),
.B(n_609),
.Y(n_1076)
);

BUFx6f_ASAP7_75t_L g1077 ( 
.A(n_991),
.Y(n_1077)
);

AOI22xp5_ASAP7_75t_L g1078 ( 
.A1(n_909),
.A2(n_610),
.B1(n_613),
.B2(n_611),
.Y(n_1078)
);

AND2x4_ASAP7_75t_L g1079 ( 
.A(n_1003),
.B(n_741),
.Y(n_1079)
);

NAND2xp5_ASAP7_75t_SL g1080 ( 
.A(n_952),
.B(n_615),
.Y(n_1080)
);

INVxp67_ASAP7_75t_L g1081 ( 
.A(n_994),
.Y(n_1081)
);

NOR2xp33_ASAP7_75t_L g1082 ( 
.A(n_981),
.B(n_627),
.Y(n_1082)
);

INVxp67_ASAP7_75t_L g1083 ( 
.A(n_1002),
.Y(n_1083)
);

OR2x6_ASAP7_75t_L g1084 ( 
.A(n_960),
.B(n_746),
.Y(n_1084)
);

NAND2xp33_ASAP7_75t_L g1085 ( 
.A(n_932),
.B(n_995),
.Y(n_1085)
);

INVx2_ASAP7_75t_L g1086 ( 
.A(n_964),
.Y(n_1086)
);

O2A1O1Ixp33_ASAP7_75t_L g1087 ( 
.A1(n_938),
.A2(n_747),
.B(n_890),
.C(n_885),
.Y(n_1087)
);

NOR2xp33_ASAP7_75t_L g1088 ( 
.A(n_930),
.B(n_628),
.Y(n_1088)
);

NOR2xp33_ASAP7_75t_L g1089 ( 
.A(n_962),
.B(n_629),
.Y(n_1089)
);

INVx2_ASAP7_75t_L g1090 ( 
.A(n_966),
.Y(n_1090)
);

INVx2_ASAP7_75t_L g1091 ( 
.A(n_974),
.Y(n_1091)
);

NOR2xp33_ASAP7_75t_SL g1092 ( 
.A(n_985),
.B(n_630),
.Y(n_1092)
);

NAND2xp5_ASAP7_75t_L g1093 ( 
.A(n_997),
.B(n_641),
.Y(n_1093)
);

AND2x4_ASAP7_75t_L g1094 ( 
.A(n_989),
.B(n_229),
.Y(n_1094)
);

INVx2_ASAP7_75t_SL g1095 ( 
.A(n_906),
.Y(n_1095)
);

NOR2xp33_ASAP7_75t_L g1096 ( 
.A(n_1000),
.B(n_631),
.Y(n_1096)
);

INVx1_ASAP7_75t_L g1097 ( 
.A(n_945),
.Y(n_1097)
);

AND2x2_ASAP7_75t_L g1098 ( 
.A(n_995),
.B(n_638),
.Y(n_1098)
);

NAND2xp5_ASAP7_75t_L g1099 ( 
.A(n_946),
.B(n_645),
.Y(n_1099)
);

INVx2_ASAP7_75t_SL g1100 ( 
.A(n_1004),
.Y(n_1100)
);

OAI22xp33_ASAP7_75t_L g1101 ( 
.A1(n_972),
.A2(n_640),
.B1(n_644),
.B2(n_634),
.Y(n_1101)
);

NAND2xp5_ASAP7_75t_L g1102 ( 
.A(n_950),
.B(n_650),
.Y(n_1102)
);

NAND2xp5_ASAP7_75t_L g1103 ( 
.A(n_955),
.B(n_652),
.Y(n_1103)
);

AOI22xp33_ASAP7_75t_L g1104 ( 
.A1(n_958),
.A2(n_647),
.B1(n_777),
.B2(n_656),
.Y(n_1104)
);

NAND2xp5_ASAP7_75t_L g1105 ( 
.A(n_959),
.B(n_992),
.Y(n_1105)
);

NAND2xp5_ASAP7_75t_L g1106 ( 
.A(n_993),
.B(n_996),
.Y(n_1106)
);

INVx1_ASAP7_75t_L g1107 ( 
.A(n_1001),
.Y(n_1107)
);

INVx2_ASAP7_75t_L g1108 ( 
.A(n_998),
.Y(n_1108)
);

HB1xp67_ASAP7_75t_L g1109 ( 
.A(n_961),
.Y(n_1109)
);

INVx1_ASAP7_75t_L g1110 ( 
.A(n_961),
.Y(n_1110)
);

INVx2_ASAP7_75t_L g1111 ( 
.A(n_976),
.Y(n_1111)
);

NOR2x1p5_ASAP7_75t_L g1112 ( 
.A(n_976),
.B(n_646),
.Y(n_1112)
);

INVx1_ASAP7_75t_L g1113 ( 
.A(n_978),
.Y(n_1113)
);

NAND2xp5_ASAP7_75t_SL g1114 ( 
.A(n_939),
.B(n_654),
.Y(n_1114)
);

INVx2_ASAP7_75t_L g1115 ( 
.A(n_982),
.Y(n_1115)
);

NOR2xp33_ASAP7_75t_L g1116 ( 
.A(n_939),
.B(n_649),
.Y(n_1116)
);

INVxp67_ASAP7_75t_L g1117 ( 
.A(n_978),
.Y(n_1117)
);

AND2x2_ASAP7_75t_L g1118 ( 
.A(n_978),
.B(n_638),
.Y(n_1118)
);

AO22x1_ASAP7_75t_L g1119 ( 
.A1(n_978),
.A2(n_655),
.B1(n_657),
.B2(n_651),
.Y(n_1119)
);

AOI21xp5_ASAP7_75t_L g1120 ( 
.A1(n_899),
.A2(n_885),
.B(n_882),
.Y(n_1120)
);

BUFx8_ASAP7_75t_L g1121 ( 
.A(n_904),
.Y(n_1121)
);

INVx5_ASAP7_75t_L g1122 ( 
.A(n_924),
.Y(n_1122)
);

BUFx3_ASAP7_75t_L g1123 ( 
.A(n_924),
.Y(n_1123)
);

AND2x6_ASAP7_75t_SL g1124 ( 
.A(n_937),
.B(n_661),
.Y(n_1124)
);

AOI21xp5_ASAP7_75t_L g1125 ( 
.A1(n_899),
.A2(n_885),
.B(n_882),
.Y(n_1125)
);

INVxp67_ASAP7_75t_L g1126 ( 
.A(n_904),
.Y(n_1126)
);

NAND2xp33_ASAP7_75t_L g1127 ( 
.A(n_999),
.B(n_660),
.Y(n_1127)
);

OAI22xp5_ASAP7_75t_L g1128 ( 
.A1(n_999),
.A2(n_667),
.B1(n_662),
.B2(n_669),
.Y(n_1128)
);

INVx2_ASAP7_75t_L g1129 ( 
.A(n_897),
.Y(n_1129)
);

NAND2xp5_ASAP7_75t_L g1130 ( 
.A(n_944),
.B(n_777),
.Y(n_1130)
);

INVx1_ASAP7_75t_L g1131 ( 
.A(n_897),
.Y(n_1131)
);

NAND2xp5_ASAP7_75t_L g1132 ( 
.A(n_944),
.B(n_872),
.Y(n_1132)
);

NAND2xp5_ASAP7_75t_L g1133 ( 
.A(n_944),
.B(n_0),
.Y(n_1133)
);

NAND2xp5_ASAP7_75t_L g1134 ( 
.A(n_944),
.B(n_0),
.Y(n_1134)
);

NAND2xp5_ASAP7_75t_L g1135 ( 
.A(n_944),
.B(n_1),
.Y(n_1135)
);

NAND2xp5_ASAP7_75t_L g1136 ( 
.A(n_944),
.B(n_2),
.Y(n_1136)
);

A2O1A1Ixp33_ASAP7_75t_L g1137 ( 
.A1(n_937),
.A2(n_6),
.B(n_4),
.C(n_5),
.Y(n_1137)
);

AND2x6_ASAP7_75t_SL g1138 ( 
.A(n_937),
.B(n_4),
.Y(n_1138)
);

NAND2xp5_ASAP7_75t_L g1139 ( 
.A(n_944),
.B(n_5),
.Y(n_1139)
);

NOR2xp33_ASAP7_75t_L g1140 ( 
.A(n_917),
.B(n_6),
.Y(n_1140)
);

NAND2xp5_ASAP7_75t_SL g1141 ( 
.A(n_948),
.B(n_231),
.Y(n_1141)
);

INVx2_ASAP7_75t_L g1142 ( 
.A(n_897),
.Y(n_1142)
);

NAND2xp5_ASAP7_75t_SL g1143 ( 
.A(n_948),
.B(n_232),
.Y(n_1143)
);

NAND2xp5_ASAP7_75t_SL g1144 ( 
.A(n_948),
.B(n_233),
.Y(n_1144)
);

NAND2xp5_ASAP7_75t_L g1145 ( 
.A(n_944),
.B(n_7),
.Y(n_1145)
);

AO221x1_ASAP7_75t_L g1146 ( 
.A1(n_970),
.A2(n_9),
.B1(n_7),
.B2(n_8),
.C(n_10),
.Y(n_1146)
);

AND2x2_ASAP7_75t_L g1147 ( 
.A(n_898),
.B(n_8),
.Y(n_1147)
);

INVx1_ASAP7_75t_L g1148 ( 
.A(n_897),
.Y(n_1148)
);

OAI221xp5_ASAP7_75t_L g1149 ( 
.A1(n_937),
.A2(n_11),
.B1(n_9),
.B2(n_10),
.C(n_12),
.Y(n_1149)
);

INVx2_ASAP7_75t_L g1150 ( 
.A(n_897),
.Y(n_1150)
);

INVx1_ASAP7_75t_L g1151 ( 
.A(n_897),
.Y(n_1151)
);

NOR2xp67_ASAP7_75t_L g1152 ( 
.A(n_947),
.B(n_236),
.Y(n_1152)
);

INVx1_ASAP7_75t_L g1153 ( 
.A(n_897),
.Y(n_1153)
);

NOR2xp33_ASAP7_75t_R g1154 ( 
.A(n_979),
.B(n_238),
.Y(n_1154)
);

AOI22xp33_ASAP7_75t_L g1155 ( 
.A1(n_937),
.A2(n_13),
.B1(n_11),
.B2(n_12),
.Y(n_1155)
);

NAND2xp5_ASAP7_75t_L g1156 ( 
.A(n_944),
.B(n_13),
.Y(n_1156)
);

INVx2_ASAP7_75t_L g1157 ( 
.A(n_897),
.Y(n_1157)
);

INVx4_ASAP7_75t_L g1158 ( 
.A(n_980),
.Y(n_1158)
);

NAND2xp5_ASAP7_75t_L g1159 ( 
.A(n_944),
.B(n_14),
.Y(n_1159)
);

NAND2xp5_ASAP7_75t_L g1160 ( 
.A(n_944),
.B(n_15),
.Y(n_1160)
);

BUFx4f_ASAP7_75t_L g1161 ( 
.A(n_924),
.Y(n_1161)
);

NAND2xp5_ASAP7_75t_SL g1162 ( 
.A(n_948),
.B(n_240),
.Y(n_1162)
);

INVx2_ASAP7_75t_L g1163 ( 
.A(n_897),
.Y(n_1163)
);

NAND2xp5_ASAP7_75t_L g1164 ( 
.A(n_944),
.B(n_15),
.Y(n_1164)
);

NAND2xp5_ASAP7_75t_L g1165 ( 
.A(n_944),
.B(n_16),
.Y(n_1165)
);

NOR2xp33_ASAP7_75t_R g1166 ( 
.A(n_1056),
.B(n_241),
.Y(n_1166)
);

BUFx6f_ASAP7_75t_L g1167 ( 
.A(n_1041),
.Y(n_1167)
);

NAND2xp5_ASAP7_75t_L g1168 ( 
.A(n_1015),
.B(n_16),
.Y(n_1168)
);

BUFx6f_ASAP7_75t_L g1169 ( 
.A(n_1041),
.Y(n_1169)
);

NAND2xp5_ASAP7_75t_L g1170 ( 
.A(n_1109),
.B(n_18),
.Y(n_1170)
);

INVx2_ASAP7_75t_SL g1171 ( 
.A(n_1028),
.Y(n_1171)
);

BUFx6f_ASAP7_75t_L g1172 ( 
.A(n_1041),
.Y(n_1172)
);

INVx1_ASAP7_75t_L g1173 ( 
.A(n_1048),
.Y(n_1173)
);

NOR2xp33_ASAP7_75t_L g1174 ( 
.A(n_1013),
.B(n_19),
.Y(n_1174)
);

INVx2_ASAP7_75t_SL g1175 ( 
.A(n_1005),
.Y(n_1175)
);

INVx2_ASAP7_75t_L g1176 ( 
.A(n_1129),
.Y(n_1176)
);

BUFx2_ASAP7_75t_L g1177 ( 
.A(n_1121),
.Y(n_1177)
);

AND2x4_ASAP7_75t_L g1178 ( 
.A(n_1122),
.B(n_1123),
.Y(n_1178)
);

HB1xp67_ASAP7_75t_L g1179 ( 
.A(n_1007),
.Y(n_1179)
);

INVx1_ASAP7_75t_SL g1180 ( 
.A(n_1012),
.Y(n_1180)
);

AND2x4_ASAP7_75t_L g1181 ( 
.A(n_1122),
.B(n_243),
.Y(n_1181)
);

BUFx3_ASAP7_75t_L g1182 ( 
.A(n_1012),
.Y(n_1182)
);

INVx1_ASAP7_75t_L g1183 ( 
.A(n_1059),
.Y(n_1183)
);

INVx1_ASAP7_75t_L g1184 ( 
.A(n_1065),
.Y(n_1184)
);

CKINVDCx5p33_ASAP7_75t_R g1185 ( 
.A(n_1012),
.Y(n_1185)
);

BUFx3_ASAP7_75t_L g1186 ( 
.A(n_1121),
.Y(n_1186)
);

NAND2xp5_ASAP7_75t_L g1187 ( 
.A(n_1027),
.B(n_19),
.Y(n_1187)
);

BUFx2_ASAP7_75t_L g1188 ( 
.A(n_1126),
.Y(n_1188)
);

NAND2xp5_ASAP7_75t_L g1189 ( 
.A(n_1147),
.B(n_20),
.Y(n_1189)
);

BUFx2_ASAP7_75t_L g1190 ( 
.A(n_1084),
.Y(n_1190)
);

INVx1_ASAP7_75t_L g1191 ( 
.A(n_1068),
.Y(n_1191)
);

AND2x4_ASAP7_75t_L g1192 ( 
.A(n_1122),
.B(n_245),
.Y(n_1192)
);

NAND2xp33_ASAP7_75t_R g1193 ( 
.A(n_1154),
.B(n_1025),
.Y(n_1193)
);

BUFx3_ASAP7_75t_L g1194 ( 
.A(n_1052),
.Y(n_1194)
);

NAND2xp5_ASAP7_75t_L g1195 ( 
.A(n_1010),
.B(n_21),
.Y(n_1195)
);

BUFx3_ASAP7_75t_L g1196 ( 
.A(n_1158),
.Y(n_1196)
);

NAND2xp5_ASAP7_75t_L g1197 ( 
.A(n_1133),
.B(n_21),
.Y(n_1197)
);

NAND2xp5_ASAP7_75t_L g1198 ( 
.A(n_1134),
.B(n_22),
.Y(n_1198)
);

BUFx10_ASAP7_75t_L g1199 ( 
.A(n_1031),
.Y(n_1199)
);

INVxp67_ASAP7_75t_L g1200 ( 
.A(n_1032),
.Y(n_1200)
);

INVx2_ASAP7_75t_L g1201 ( 
.A(n_1142),
.Y(n_1201)
);

A2O1A1Ixp33_ASAP7_75t_L g1202 ( 
.A1(n_1140),
.A2(n_25),
.B(n_23),
.C(n_24),
.Y(n_1202)
);

A2O1A1Ixp33_ASAP7_75t_L g1203 ( 
.A1(n_1116),
.A2(n_25),
.B(n_23),
.C(n_24),
.Y(n_1203)
);

NAND2xp5_ASAP7_75t_L g1204 ( 
.A(n_1135),
.B(n_26),
.Y(n_1204)
);

BUFx4f_ASAP7_75t_L g1205 ( 
.A(n_1084),
.Y(n_1205)
);

AOI22xp5_ASAP7_75t_L g1206 ( 
.A1(n_1024),
.A2(n_248),
.B1(n_249),
.B2(n_247),
.Y(n_1206)
);

INVx4_ASAP7_75t_L g1207 ( 
.A(n_1161),
.Y(n_1207)
);

NOR3xp33_ASAP7_75t_SL g1208 ( 
.A(n_1016),
.B(n_27),
.C(n_28),
.Y(n_1208)
);

INVx2_ASAP7_75t_L g1209 ( 
.A(n_1150),
.Y(n_1209)
);

NAND2xp5_ASAP7_75t_L g1210 ( 
.A(n_1136),
.B(n_27),
.Y(n_1210)
);

NOR3xp33_ASAP7_75t_SL g1211 ( 
.A(n_1088),
.B(n_28),
.C(n_29),
.Y(n_1211)
);

INVx2_ASAP7_75t_L g1212 ( 
.A(n_1157),
.Y(n_1212)
);

NAND2xp33_ASAP7_75t_SL g1213 ( 
.A(n_1069),
.B(n_30),
.Y(n_1213)
);

INVx1_ASAP7_75t_L g1214 ( 
.A(n_1037),
.Y(n_1214)
);

NOR3xp33_ASAP7_75t_SL g1215 ( 
.A(n_1051),
.B(n_31),
.C(n_32),
.Y(n_1215)
);

CKINVDCx20_ASAP7_75t_R g1216 ( 
.A(n_1095),
.Y(n_1216)
);

AND2x4_ASAP7_75t_L g1217 ( 
.A(n_1006),
.B(n_251),
.Y(n_1217)
);

OR2x6_ASAP7_75t_L g1218 ( 
.A(n_1158),
.B(n_34),
.Y(n_1218)
);

AOI21xp5_ASAP7_75t_L g1219 ( 
.A1(n_1085),
.A2(n_1026),
.B(n_1067),
.Y(n_1219)
);

OR2x2_ASAP7_75t_L g1220 ( 
.A(n_1063),
.B(n_34),
.Y(n_1220)
);

AND2x4_ASAP7_75t_L g1221 ( 
.A(n_1077),
.B(n_252),
.Y(n_1221)
);

INVx2_ASAP7_75t_L g1222 ( 
.A(n_1163),
.Y(n_1222)
);

NAND2xp5_ASAP7_75t_L g1223 ( 
.A(n_1139),
.B(n_35),
.Y(n_1223)
);

NAND2xp5_ASAP7_75t_SL g1224 ( 
.A(n_1077),
.B(n_255),
.Y(n_1224)
);

CKINVDCx5p33_ASAP7_75t_R g1225 ( 
.A(n_1008),
.Y(n_1225)
);

INVx1_ASAP7_75t_L g1226 ( 
.A(n_1131),
.Y(n_1226)
);

NAND2xp5_ASAP7_75t_L g1227 ( 
.A(n_1145),
.B(n_35),
.Y(n_1227)
);

NOR2xp33_ASAP7_75t_L g1228 ( 
.A(n_1089),
.B(n_36),
.Y(n_1228)
);

OAI21xp5_ASAP7_75t_L g1229 ( 
.A1(n_1017),
.A2(n_257),
.B(n_256),
.Y(n_1229)
);

AND2x4_ASAP7_75t_L g1230 ( 
.A(n_1079),
.B(n_259),
.Y(n_1230)
);

OR2x6_ASAP7_75t_L g1231 ( 
.A(n_1084),
.B(n_36),
.Y(n_1231)
);

NOR3xp33_ASAP7_75t_SL g1232 ( 
.A(n_1082),
.B(n_37),
.C(n_38),
.Y(n_1232)
);

AND2x2_ASAP7_75t_L g1233 ( 
.A(n_1029),
.B(n_37),
.Y(n_1233)
);

INVx2_ASAP7_75t_L g1234 ( 
.A(n_1148),
.Y(n_1234)
);

INVx1_ASAP7_75t_L g1235 ( 
.A(n_1151),
.Y(n_1235)
);

CKINVDCx5p33_ASAP7_75t_R g1236 ( 
.A(n_1034),
.Y(n_1236)
);

NOR2xp33_ASAP7_75t_L g1237 ( 
.A(n_1045),
.B(n_39),
.Y(n_1237)
);

CKINVDCx5p33_ASAP7_75t_R g1238 ( 
.A(n_1069),
.Y(n_1238)
);

AND2x4_ASAP7_75t_L g1239 ( 
.A(n_1079),
.B(n_260),
.Y(n_1239)
);

INVx1_ASAP7_75t_L g1240 ( 
.A(n_1153),
.Y(n_1240)
);

BUFx6f_ASAP7_75t_L g1241 ( 
.A(n_1161),
.Y(n_1241)
);

NOR3xp33_ASAP7_75t_SL g1242 ( 
.A(n_1149),
.B(n_40),
.C(n_41),
.Y(n_1242)
);

INVx5_ASAP7_75t_L g1243 ( 
.A(n_1009),
.Y(n_1243)
);

HB1xp67_ASAP7_75t_L g1244 ( 
.A(n_1049),
.Y(n_1244)
);

NAND2xp5_ASAP7_75t_L g1245 ( 
.A(n_1156),
.B(n_41),
.Y(n_1245)
);

INVx2_ASAP7_75t_L g1246 ( 
.A(n_1040),
.Y(n_1246)
);

AND2x4_ASAP7_75t_L g1247 ( 
.A(n_1112),
.B(n_261),
.Y(n_1247)
);

NAND2xp5_ASAP7_75t_L g1248 ( 
.A(n_1159),
.B(n_42),
.Y(n_1248)
);

INVx4_ASAP7_75t_L g1249 ( 
.A(n_1044),
.Y(n_1249)
);

INVx1_ASAP7_75t_L g1250 ( 
.A(n_1097),
.Y(n_1250)
);

BUFx2_ASAP7_75t_L g1251 ( 
.A(n_1081),
.Y(n_1251)
);

INVxp67_ASAP7_75t_SL g1252 ( 
.A(n_1018),
.Y(n_1252)
);

INVx3_ASAP7_75t_L g1253 ( 
.A(n_1094),
.Y(n_1253)
);

INVx1_ASAP7_75t_L g1254 ( 
.A(n_1033),
.Y(n_1254)
);

INVx1_ASAP7_75t_L g1255 ( 
.A(n_1105),
.Y(n_1255)
);

INVx1_ASAP7_75t_SL g1256 ( 
.A(n_1073),
.Y(n_1256)
);

NAND2xp5_ASAP7_75t_SL g1257 ( 
.A(n_1160),
.B(n_262),
.Y(n_1257)
);

INVx2_ASAP7_75t_L g1258 ( 
.A(n_1086),
.Y(n_1258)
);

BUFx6f_ASAP7_75t_L g1259 ( 
.A(n_1009),
.Y(n_1259)
);

BUFx12f_ASAP7_75t_L g1260 ( 
.A(n_1124),
.Y(n_1260)
);

INVx2_ASAP7_75t_L g1261 ( 
.A(n_1090),
.Y(n_1261)
);

AND2x4_ASAP7_75t_L g1262 ( 
.A(n_1054),
.B(n_263),
.Y(n_1262)
);

NAND2xp5_ASAP7_75t_L g1263 ( 
.A(n_1164),
.B(n_43),
.Y(n_1263)
);

NAND2xp5_ASAP7_75t_L g1264 ( 
.A(n_1165),
.B(n_43),
.Y(n_1264)
);

INVx2_ASAP7_75t_L g1265 ( 
.A(n_1091),
.Y(n_1265)
);

BUFx2_ASAP7_75t_L g1266 ( 
.A(n_1083),
.Y(n_1266)
);

BUFx2_ASAP7_75t_L g1267 ( 
.A(n_1055),
.Y(n_1267)
);

NOR2x1_ASAP7_75t_L g1268 ( 
.A(n_1047),
.B(n_1044),
.Y(n_1268)
);

BUFx6f_ASAP7_75t_L g1269 ( 
.A(n_1009),
.Y(n_1269)
);

INVx1_ASAP7_75t_L g1270 ( 
.A(n_1035),
.Y(n_1270)
);

INVx2_ASAP7_75t_L g1271 ( 
.A(n_1108),
.Y(n_1271)
);

NAND2xp5_ASAP7_75t_L g1272 ( 
.A(n_1110),
.B(n_44),
.Y(n_1272)
);

INVx2_ASAP7_75t_L g1273 ( 
.A(n_1107),
.Y(n_1273)
);

NAND2xp5_ASAP7_75t_L g1274 ( 
.A(n_1111),
.B(n_45),
.Y(n_1274)
);

AOI22xp5_ASAP7_75t_L g1275 ( 
.A1(n_1096),
.A2(n_265),
.B1(n_267),
.B2(n_264),
.Y(n_1275)
);

OAI31xp33_ASAP7_75t_SL g1276 ( 
.A1(n_1058),
.A2(n_48),
.A3(n_45),
.B(n_47),
.Y(n_1276)
);

BUFx6f_ASAP7_75t_L g1277 ( 
.A(n_1094),
.Y(n_1277)
);

INVxp67_ASAP7_75t_SL g1278 ( 
.A(n_1018),
.Y(n_1278)
);

CKINVDCx5p33_ASAP7_75t_R g1279 ( 
.A(n_1138),
.Y(n_1279)
);

INVx3_ASAP7_75t_L g1280 ( 
.A(n_1100),
.Y(n_1280)
);

NAND2xp5_ASAP7_75t_L g1281 ( 
.A(n_1011),
.B(n_49),
.Y(n_1281)
);

INVx2_ASAP7_75t_L g1282 ( 
.A(n_1030),
.Y(n_1282)
);

NAND2xp5_ASAP7_75t_L g1283 ( 
.A(n_1132),
.B(n_50),
.Y(n_1283)
);

AND2x4_ASAP7_75t_L g1284 ( 
.A(n_1044),
.B(n_268),
.Y(n_1284)
);

BUFx4f_ASAP7_75t_L g1285 ( 
.A(n_1064),
.Y(n_1285)
);

INVx1_ASAP7_75t_L g1286 ( 
.A(n_1106),
.Y(n_1286)
);

BUFx2_ASAP7_75t_L g1287 ( 
.A(n_1118),
.Y(n_1287)
);

BUFx3_ASAP7_75t_L g1288 ( 
.A(n_1098),
.Y(n_1288)
);

BUFx2_ASAP7_75t_L g1289 ( 
.A(n_1093),
.Y(n_1289)
);

AND2x4_ASAP7_75t_L g1290 ( 
.A(n_1050),
.B(n_269),
.Y(n_1290)
);

INVx2_ASAP7_75t_L g1291 ( 
.A(n_1115),
.Y(n_1291)
);

AND2x4_ASAP7_75t_L g1292 ( 
.A(n_1014),
.B(n_271),
.Y(n_1292)
);

AND2x6_ASAP7_75t_L g1293 ( 
.A(n_1113),
.B(n_273),
.Y(n_1293)
);

NAND2xp5_ASAP7_75t_SL g1294 ( 
.A(n_1092),
.B(n_274),
.Y(n_1294)
);

OR2x6_ASAP7_75t_L g1295 ( 
.A(n_1060),
.B(n_51),
.Y(n_1295)
);

XOR2xp5_ASAP7_75t_L g1296 ( 
.A(n_1078),
.B(n_52),
.Y(n_1296)
);

AOI22xp5_ASAP7_75t_L g1297 ( 
.A1(n_1039),
.A2(n_1127),
.B1(n_1053),
.B2(n_1038),
.Y(n_1297)
);

NAND2xp5_ASAP7_75t_SL g1298 ( 
.A(n_1070),
.B(n_276),
.Y(n_1298)
);

BUFx4f_ASAP7_75t_L g1299 ( 
.A(n_1146),
.Y(n_1299)
);

AOI22xp33_ASAP7_75t_L g1300 ( 
.A1(n_1155),
.A2(n_54),
.B1(n_52),
.B2(n_53),
.Y(n_1300)
);

INVx4_ASAP7_75t_L g1301 ( 
.A(n_1071),
.Y(n_1301)
);

AOI22xp33_ASAP7_75t_L g1302 ( 
.A1(n_1141),
.A2(n_59),
.B1(n_56),
.B2(n_58),
.Y(n_1302)
);

INVx6_ASAP7_75t_L g1303 ( 
.A(n_1101),
.Y(n_1303)
);

INVx2_ASAP7_75t_L g1304 ( 
.A(n_1021),
.Y(n_1304)
);

CKINVDCx5p33_ASAP7_75t_R g1305 ( 
.A(n_1128),
.Y(n_1305)
);

NAND2xp5_ASAP7_75t_L g1306 ( 
.A(n_1023),
.B(n_56),
.Y(n_1306)
);

NOR2xp33_ASAP7_75t_R g1307 ( 
.A(n_1061),
.B(n_279),
.Y(n_1307)
);

BUFx6f_ASAP7_75t_L g1308 ( 
.A(n_1143),
.Y(n_1308)
);

INVx1_ASAP7_75t_L g1309 ( 
.A(n_1043),
.Y(n_1309)
);

NAND3xp33_ASAP7_75t_SL g1310 ( 
.A(n_1137),
.B(n_59),
.C(n_60),
.Y(n_1310)
);

NOR2xp33_ASAP7_75t_R g1311 ( 
.A(n_1062),
.B(n_280),
.Y(n_1311)
);

BUFx6f_ASAP7_75t_L g1312 ( 
.A(n_1144),
.Y(n_1312)
);

BUFx3_ASAP7_75t_L g1313 ( 
.A(n_1046),
.Y(n_1313)
);

OAI22xp5_ASAP7_75t_L g1314 ( 
.A1(n_1130),
.A2(n_284),
.B1(n_285),
.B2(n_282),
.Y(n_1314)
);

NOR2xp33_ASAP7_75t_L g1315 ( 
.A(n_1020),
.B(n_60),
.Y(n_1315)
);

INVx1_ASAP7_75t_L g1316 ( 
.A(n_1099),
.Y(n_1316)
);

INVx8_ASAP7_75t_L g1317 ( 
.A(n_1074),
.Y(n_1317)
);

AND2x4_ASAP7_75t_L g1318 ( 
.A(n_1117),
.B(n_286),
.Y(n_1318)
);

HB1xp67_ASAP7_75t_L g1319 ( 
.A(n_1066),
.Y(n_1319)
);

BUFx6f_ASAP7_75t_L g1320 ( 
.A(n_1162),
.Y(n_1320)
);

BUFx3_ASAP7_75t_L g1321 ( 
.A(n_1102),
.Y(n_1321)
);

INVx2_ASAP7_75t_L g1322 ( 
.A(n_1103),
.Y(n_1322)
);

BUFx6f_ASAP7_75t_L g1323 ( 
.A(n_1080),
.Y(n_1323)
);

BUFx6f_ASAP7_75t_L g1324 ( 
.A(n_1076),
.Y(n_1324)
);

INVx2_ASAP7_75t_L g1325 ( 
.A(n_1114),
.Y(n_1325)
);

INVx2_ASAP7_75t_L g1326 ( 
.A(n_1036),
.Y(n_1326)
);

AND2x4_ASAP7_75t_L g1327 ( 
.A(n_1152),
.B(n_287),
.Y(n_1327)
);

NAND2xp5_ASAP7_75t_L g1328 ( 
.A(n_1022),
.B(n_62),
.Y(n_1328)
);

INVx1_ASAP7_75t_SL g1329 ( 
.A(n_1119),
.Y(n_1329)
);

AND2x4_ASAP7_75t_L g1330 ( 
.A(n_1152),
.B(n_289),
.Y(n_1330)
);

HB1xp67_ASAP7_75t_L g1331 ( 
.A(n_1075),
.Y(n_1331)
);

AND2x4_ASAP7_75t_L g1332 ( 
.A(n_1120),
.B(n_291),
.Y(n_1332)
);

CKINVDCx5p33_ASAP7_75t_R g1333 ( 
.A(n_1072),
.Y(n_1333)
);

NAND2xp5_ASAP7_75t_L g1334 ( 
.A(n_1254),
.B(n_1019),
.Y(n_1334)
);

AOI21xp5_ASAP7_75t_L g1335 ( 
.A1(n_1219),
.A2(n_1125),
.B(n_1087),
.Y(n_1335)
);

NAND2xp5_ASAP7_75t_L g1336 ( 
.A(n_1255),
.B(n_1042),
.Y(n_1336)
);

NAND2xp5_ASAP7_75t_SL g1337 ( 
.A(n_1199),
.B(n_1057),
.Y(n_1337)
);

AOI21x1_ASAP7_75t_L g1338 ( 
.A1(n_1283),
.A2(n_1104),
.B(n_293),
.Y(n_1338)
);

AND2x4_ASAP7_75t_L g1339 ( 
.A(n_1207),
.B(n_488),
.Y(n_1339)
);

AND2x2_ASAP7_75t_L g1340 ( 
.A(n_1200),
.B(n_64),
.Y(n_1340)
);

OAI22xp5_ASAP7_75t_L g1341 ( 
.A1(n_1253),
.A2(n_68),
.B1(n_66),
.B2(n_67),
.Y(n_1341)
);

INVx3_ASAP7_75t_L g1342 ( 
.A(n_1196),
.Y(n_1342)
);

OAI21x1_ASAP7_75t_L g1343 ( 
.A1(n_1229),
.A2(n_297),
.B(n_295),
.Y(n_1343)
);

NAND2xp5_ASAP7_75t_L g1344 ( 
.A(n_1286),
.B(n_67),
.Y(n_1344)
);

OAI21x1_ASAP7_75t_SL g1345 ( 
.A1(n_1272),
.A2(n_1325),
.B(n_1249),
.Y(n_1345)
);

NAND2xp5_ASAP7_75t_L g1346 ( 
.A(n_1309),
.B(n_68),
.Y(n_1346)
);

NAND2xp5_ASAP7_75t_L g1347 ( 
.A(n_1316),
.B(n_69),
.Y(n_1347)
);

BUFx6f_ASAP7_75t_L g1348 ( 
.A(n_1241),
.Y(n_1348)
);

NAND2xp5_ASAP7_75t_L g1349 ( 
.A(n_1262),
.B(n_69),
.Y(n_1349)
);

OAI21xp5_ASAP7_75t_L g1350 ( 
.A1(n_1187),
.A2(n_299),
.B(n_298),
.Y(n_1350)
);

INVx1_ASAP7_75t_L g1351 ( 
.A(n_1173),
.Y(n_1351)
);

AOI21xp5_ASAP7_75t_L g1352 ( 
.A1(n_1322),
.A2(n_301),
.B(n_300),
.Y(n_1352)
);

OAI21x1_ASAP7_75t_L g1353 ( 
.A1(n_1268),
.A2(n_305),
.B(n_304),
.Y(n_1353)
);

BUFx3_ASAP7_75t_L g1354 ( 
.A(n_1182),
.Y(n_1354)
);

NOR2xp33_ASAP7_75t_L g1355 ( 
.A(n_1319),
.B(n_70),
.Y(n_1355)
);

INVx4_ASAP7_75t_L g1356 ( 
.A(n_1241),
.Y(n_1356)
);

INVx1_ASAP7_75t_L g1357 ( 
.A(n_1183),
.Y(n_1357)
);

NAND2xp5_ASAP7_75t_SL g1358 ( 
.A(n_1199),
.B(n_70),
.Y(n_1358)
);

OR2x6_ASAP7_75t_L g1359 ( 
.A(n_1241),
.B(n_307),
.Y(n_1359)
);

OAI21x1_ASAP7_75t_L g1360 ( 
.A1(n_1291),
.A2(n_309),
.B(n_308),
.Y(n_1360)
);

BUFx3_ASAP7_75t_L g1361 ( 
.A(n_1194),
.Y(n_1361)
);

OAI21x1_ASAP7_75t_L g1362 ( 
.A1(n_1304),
.A2(n_311),
.B(n_310),
.Y(n_1362)
);

AND2x4_ASAP7_75t_L g1363 ( 
.A(n_1178),
.B(n_486),
.Y(n_1363)
);

AOI21x1_ASAP7_75t_L g1364 ( 
.A1(n_1306),
.A2(n_313),
.B(n_312),
.Y(n_1364)
);

AOI21xp5_ASAP7_75t_L g1365 ( 
.A1(n_1332),
.A2(n_316),
.B(n_314),
.Y(n_1365)
);

AOI22xp5_ASAP7_75t_SL g1366 ( 
.A1(n_1296),
.A2(n_73),
.B1(n_71),
.B2(n_72),
.Y(n_1366)
);

NAND2xp5_ASAP7_75t_L g1367 ( 
.A(n_1262),
.B(n_71),
.Y(n_1367)
);

BUFx6f_ASAP7_75t_L g1368 ( 
.A(n_1167),
.Y(n_1368)
);

OR2x6_ASAP7_75t_L g1369 ( 
.A(n_1186),
.B(n_321),
.Y(n_1369)
);

NOR2x1_ASAP7_75t_L g1370 ( 
.A(n_1216),
.B(n_322),
.Y(n_1370)
);

AOI21xp5_ASAP7_75t_L g1371 ( 
.A1(n_1270),
.A2(n_325),
.B(n_324),
.Y(n_1371)
);

AO31x2_ASAP7_75t_L g1372 ( 
.A1(n_1237),
.A2(n_75),
.A3(n_73),
.B(n_74),
.Y(n_1372)
);

NAND2x1p5_ASAP7_75t_L g1373 ( 
.A(n_1243),
.B(n_326),
.Y(n_1373)
);

INVx3_ASAP7_75t_L g1374 ( 
.A(n_1178),
.Y(n_1374)
);

OAI21x1_ASAP7_75t_L g1375 ( 
.A1(n_1257),
.A2(n_329),
.B(n_328),
.Y(n_1375)
);

INVx1_ASAP7_75t_L g1376 ( 
.A(n_1184),
.Y(n_1376)
);

AOI21xp5_ASAP7_75t_L g1377 ( 
.A1(n_1331),
.A2(n_1297),
.B(n_1298),
.Y(n_1377)
);

OAI21x1_ASAP7_75t_L g1378 ( 
.A1(n_1281),
.A2(n_1314),
.B(n_1274),
.Y(n_1378)
);

OAI21x1_ASAP7_75t_L g1379 ( 
.A1(n_1197),
.A2(n_332),
.B(n_331),
.Y(n_1379)
);

A2O1A1Ixp33_ASAP7_75t_L g1380 ( 
.A1(n_1228),
.A2(n_78),
.B(n_76),
.C(n_77),
.Y(n_1380)
);

NAND2xp5_ASAP7_75t_L g1381 ( 
.A(n_1313),
.B(n_1289),
.Y(n_1381)
);

OAI21x1_ASAP7_75t_L g1382 ( 
.A1(n_1198),
.A2(n_334),
.B(n_333),
.Y(n_1382)
);

AOI21x1_ASAP7_75t_L g1383 ( 
.A1(n_1204),
.A2(n_481),
.B(n_337),
.Y(n_1383)
);

AOI21xp5_ASAP7_75t_L g1384 ( 
.A1(n_1327),
.A2(n_1330),
.B(n_1326),
.Y(n_1384)
);

INVx1_ASAP7_75t_L g1385 ( 
.A(n_1191),
.Y(n_1385)
);

NAND2x1p5_ASAP7_75t_L g1386 ( 
.A(n_1243),
.B(n_335),
.Y(n_1386)
);

OAI21x1_ASAP7_75t_L g1387 ( 
.A1(n_1210),
.A2(n_341),
.B(n_338),
.Y(n_1387)
);

NAND2xp5_ASAP7_75t_L g1388 ( 
.A(n_1321),
.B(n_77),
.Y(n_1388)
);

OAI21xp5_ASAP7_75t_L g1389 ( 
.A1(n_1168),
.A2(n_343),
.B(n_342),
.Y(n_1389)
);

AOI21xp33_ASAP7_75t_L g1390 ( 
.A1(n_1174),
.A2(n_78),
.B(n_80),
.Y(n_1390)
);

OAI21x1_ASAP7_75t_L g1391 ( 
.A1(n_1223),
.A2(n_345),
.B(n_344),
.Y(n_1391)
);

AOI21xp5_ASAP7_75t_L g1392 ( 
.A1(n_1327),
.A2(n_348),
.B(n_346),
.Y(n_1392)
);

BUFx6f_ASAP7_75t_L g1393 ( 
.A(n_1167),
.Y(n_1393)
);

NAND2xp5_ASAP7_75t_L g1394 ( 
.A(n_1305),
.B(n_80),
.Y(n_1394)
);

OAI22xp5_ASAP7_75t_L g1395 ( 
.A1(n_1277),
.A2(n_84),
.B1(n_82),
.B2(n_83),
.Y(n_1395)
);

AOI21x1_ASAP7_75t_L g1396 ( 
.A1(n_1227),
.A2(n_351),
.B(n_349),
.Y(n_1396)
);

OR2x6_ASAP7_75t_L g1397 ( 
.A(n_1177),
.B(n_352),
.Y(n_1397)
);

A2O1A1Ixp33_ASAP7_75t_L g1398 ( 
.A1(n_1315),
.A2(n_86),
.B(n_83),
.C(n_85),
.Y(n_1398)
);

OAI21x1_ASAP7_75t_L g1399 ( 
.A1(n_1245),
.A2(n_355),
.B(n_353),
.Y(n_1399)
);

AOI21x1_ASAP7_75t_L g1400 ( 
.A1(n_1248),
.A2(n_479),
.B(n_358),
.Y(n_1400)
);

OAI21x1_ASAP7_75t_L g1401 ( 
.A1(n_1263),
.A2(n_359),
.B(n_356),
.Y(n_1401)
);

AND2x2_ASAP7_75t_SL g1402 ( 
.A(n_1276),
.B(n_85),
.Y(n_1402)
);

OAI21xp5_ASAP7_75t_L g1403 ( 
.A1(n_1264),
.A2(n_361),
.B(n_360),
.Y(n_1403)
);

OR2x6_ASAP7_75t_L g1404 ( 
.A(n_1284),
.B(n_362),
.Y(n_1404)
);

INVx1_ASAP7_75t_SL g1405 ( 
.A(n_1171),
.Y(n_1405)
);

NAND2xp5_ASAP7_75t_SL g1406 ( 
.A(n_1285),
.B(n_1244),
.Y(n_1406)
);

NAND2xp5_ASAP7_75t_L g1407 ( 
.A(n_1170),
.B(n_86),
.Y(n_1407)
);

OAI21x1_ASAP7_75t_L g1408 ( 
.A1(n_1282),
.A2(n_364),
.B(n_363),
.Y(n_1408)
);

NOR2xp33_ASAP7_75t_L g1409 ( 
.A(n_1303),
.B(n_87),
.Y(n_1409)
);

OAI21x1_ASAP7_75t_L g1410 ( 
.A1(n_1176),
.A2(n_368),
.B(n_367),
.Y(n_1410)
);

NAND2xp5_ASAP7_75t_L g1411 ( 
.A(n_1195),
.B(n_87),
.Y(n_1411)
);

INVx1_ASAP7_75t_SL g1412 ( 
.A(n_1188),
.Y(n_1412)
);

AO31x2_ASAP7_75t_L g1413 ( 
.A1(n_1203),
.A2(n_91),
.A3(n_89),
.B(n_90),
.Y(n_1413)
);

A2O1A1Ixp33_ASAP7_75t_L g1414 ( 
.A1(n_1189),
.A2(n_92),
.B(n_90),
.C(n_91),
.Y(n_1414)
);

NAND2xp5_ASAP7_75t_L g1415 ( 
.A(n_1277),
.B(n_92),
.Y(n_1415)
);

INVx3_ASAP7_75t_SL g1416 ( 
.A(n_1185),
.Y(n_1416)
);

INVx2_ASAP7_75t_SL g1417 ( 
.A(n_1288),
.Y(n_1417)
);

AOI22xp5_ASAP7_75t_L g1418 ( 
.A1(n_1303),
.A2(n_1193),
.B1(n_1267),
.B2(n_1290),
.Y(n_1418)
);

AND2x2_ASAP7_75t_L g1419 ( 
.A(n_1233),
.B(n_1287),
.Y(n_1419)
);

BUFx2_ASAP7_75t_SL g1420 ( 
.A(n_1175),
.Y(n_1420)
);

AOI21xp5_ASAP7_75t_L g1421 ( 
.A1(n_1308),
.A2(n_372),
.B(n_371),
.Y(n_1421)
);

OAI21x1_ASAP7_75t_L g1422 ( 
.A1(n_1201),
.A2(n_374),
.B(n_373),
.Y(n_1422)
);

OAI21xp5_ASAP7_75t_L g1423 ( 
.A1(n_1299),
.A2(n_377),
.B(n_376),
.Y(n_1423)
);

A2O1A1Ixp33_ASAP7_75t_L g1424 ( 
.A1(n_1328),
.A2(n_95),
.B(n_93),
.C(n_94),
.Y(n_1424)
);

OAI21x1_ASAP7_75t_L g1425 ( 
.A1(n_1209),
.A2(n_379),
.B(n_378),
.Y(n_1425)
);

AOI21xp5_ASAP7_75t_L g1426 ( 
.A1(n_1308),
.A2(n_381),
.B(n_380),
.Y(n_1426)
);

OAI22xp5_ASAP7_75t_L g1427 ( 
.A1(n_1277),
.A2(n_95),
.B1(n_93),
.B2(n_94),
.Y(n_1427)
);

NOR3xp33_ASAP7_75t_L g1428 ( 
.A(n_1310),
.B(n_97),
.C(n_98),
.Y(n_1428)
);

NOR2xp33_ASAP7_75t_L g1429 ( 
.A(n_1251),
.B(n_99),
.Y(n_1429)
);

NAND2xp5_ASAP7_75t_L g1430 ( 
.A(n_1234),
.B(n_99),
.Y(n_1430)
);

OAI21x1_ASAP7_75t_L g1431 ( 
.A1(n_1212),
.A2(n_386),
.B(n_383),
.Y(n_1431)
);

OAI22xp5_ASAP7_75t_L g1432 ( 
.A1(n_1333),
.A2(n_102),
.B1(n_100),
.B2(n_101),
.Y(n_1432)
);

NAND2xp5_ASAP7_75t_L g1433 ( 
.A(n_1273),
.B(n_100),
.Y(n_1433)
);

BUFx6f_ASAP7_75t_L g1434 ( 
.A(n_1167),
.Y(n_1434)
);

OAI21x1_ASAP7_75t_L g1435 ( 
.A1(n_1222),
.A2(n_389),
.B(n_388),
.Y(n_1435)
);

AOI21xp33_ASAP7_75t_L g1436 ( 
.A1(n_1300),
.A2(n_101),
.B(n_102),
.Y(n_1436)
);

BUFx5_ASAP7_75t_L g1437 ( 
.A(n_1293),
.Y(n_1437)
);

AOI22xp33_ASAP7_75t_L g1438 ( 
.A1(n_1296),
.A2(n_103),
.B1(n_104),
.B2(n_105),
.Y(n_1438)
);

INVx1_ASAP7_75t_L g1439 ( 
.A(n_1214),
.Y(n_1439)
);

AOI21xp5_ASAP7_75t_L g1440 ( 
.A1(n_1308),
.A2(n_391),
.B(n_390),
.Y(n_1440)
);

NOR2xp33_ASAP7_75t_L g1441 ( 
.A(n_1266),
.B(n_104),
.Y(n_1441)
);

INVx1_ASAP7_75t_SL g1442 ( 
.A(n_1179),
.Y(n_1442)
);

OAI21xp5_ASAP7_75t_L g1443 ( 
.A1(n_1271),
.A2(n_396),
.B(n_395),
.Y(n_1443)
);

OAI21x1_ASAP7_75t_L g1444 ( 
.A1(n_1224),
.A2(n_1235),
.B(n_1226),
.Y(n_1444)
);

OAI21x1_ASAP7_75t_L g1445 ( 
.A1(n_1240),
.A2(n_400),
.B(n_397),
.Y(n_1445)
);

INVx1_ASAP7_75t_L g1446 ( 
.A(n_1250),
.Y(n_1446)
);

NAND2xp5_ASAP7_75t_L g1447 ( 
.A(n_1329),
.B(n_105),
.Y(n_1447)
);

NOR2xp33_ASAP7_75t_L g1448 ( 
.A(n_1280),
.B(n_106),
.Y(n_1448)
);

OAI21xp5_ASAP7_75t_L g1449 ( 
.A1(n_1246),
.A2(n_402),
.B(n_401),
.Y(n_1449)
);

INVx1_ASAP7_75t_L g1450 ( 
.A(n_1258),
.Y(n_1450)
);

NAND2xp5_ASAP7_75t_L g1451 ( 
.A(n_1221),
.B(n_107),
.Y(n_1451)
);

NAND2xp5_ASAP7_75t_L g1452 ( 
.A(n_1221),
.B(n_107),
.Y(n_1452)
);

OAI22xp5_ASAP7_75t_L g1453 ( 
.A1(n_1252),
.A2(n_108),
.B1(n_109),
.B2(n_110),
.Y(n_1453)
);

OAI21x1_ASAP7_75t_L g1454 ( 
.A1(n_1261),
.A2(n_1265),
.B(n_1278),
.Y(n_1454)
);

INVx1_ASAP7_75t_L g1455 ( 
.A(n_1217),
.Y(n_1455)
);

OAI21xp5_ASAP7_75t_L g1456 ( 
.A1(n_1302),
.A2(n_404),
.B(n_403),
.Y(n_1456)
);

AO31x2_ASAP7_75t_L g1457 ( 
.A1(n_1202),
.A2(n_108),
.A3(n_109),
.B(n_111),
.Y(n_1457)
);

BUFx6f_ASAP7_75t_L g1458 ( 
.A(n_1169),
.Y(n_1458)
);

NAND2xp5_ASAP7_75t_SL g1459 ( 
.A(n_1324),
.B(n_111),
.Y(n_1459)
);

OAI21x1_ASAP7_75t_SL g1460 ( 
.A1(n_1206),
.A2(n_406),
.B(n_405),
.Y(n_1460)
);

A2O1A1Ixp33_ASAP7_75t_L g1461 ( 
.A1(n_1242),
.A2(n_112),
.B(n_113),
.C(n_114),
.Y(n_1461)
);

BUFx2_ASAP7_75t_L g1462 ( 
.A(n_1190),
.Y(n_1462)
);

NOR2x1_ASAP7_75t_L g1463 ( 
.A(n_1294),
.B(n_407),
.Y(n_1463)
);

OAI22xp5_ASAP7_75t_L g1464 ( 
.A1(n_1312),
.A2(n_112),
.B1(n_114),
.B2(n_115),
.Y(n_1464)
);

INVx2_ASAP7_75t_L g1465 ( 
.A(n_1169),
.Y(n_1465)
);

INVx2_ASAP7_75t_L g1466 ( 
.A(n_1169),
.Y(n_1466)
);

BUFx6f_ASAP7_75t_L g1467 ( 
.A(n_1172),
.Y(n_1467)
);

BUFx6f_ASAP7_75t_L g1468 ( 
.A(n_1172),
.Y(n_1468)
);

BUFx10_ASAP7_75t_L g1469 ( 
.A(n_1238),
.Y(n_1469)
);

INVx3_ASAP7_75t_L g1470 ( 
.A(n_1172),
.Y(n_1470)
);

AOI21xp5_ASAP7_75t_L g1471 ( 
.A1(n_1312),
.A2(n_1320),
.B(n_1192),
.Y(n_1471)
);

HB1xp67_ASAP7_75t_L g1472 ( 
.A(n_1220),
.Y(n_1472)
);

NAND2xp5_ASAP7_75t_L g1473 ( 
.A(n_1230),
.B(n_116),
.Y(n_1473)
);

NAND2xp5_ASAP7_75t_L g1474 ( 
.A(n_1230),
.B(n_118),
.Y(n_1474)
);

OAI21x1_ASAP7_75t_L g1475 ( 
.A1(n_1275),
.A2(n_409),
.B(n_408),
.Y(n_1475)
);

INVx2_ASAP7_75t_L g1476 ( 
.A(n_1217),
.Y(n_1476)
);

INVx2_ASAP7_75t_L g1477 ( 
.A(n_1318),
.Y(n_1477)
);

AO31x2_ASAP7_75t_L g1478 ( 
.A1(n_1301),
.A2(n_118),
.A3(n_119),
.B(n_120),
.Y(n_1478)
);

AOI21xp5_ASAP7_75t_L g1479 ( 
.A1(n_1312),
.A2(n_411),
.B(n_410),
.Y(n_1479)
);

INVx1_ASAP7_75t_L g1480 ( 
.A(n_1318),
.Y(n_1480)
);

NAND2xp5_ASAP7_75t_L g1481 ( 
.A(n_1239),
.B(n_119),
.Y(n_1481)
);

OAI21x1_ASAP7_75t_L g1482 ( 
.A1(n_1259),
.A2(n_1269),
.B(n_1320),
.Y(n_1482)
);

OAI21x1_ASAP7_75t_L g1483 ( 
.A1(n_1259),
.A2(n_413),
.B(n_412),
.Y(n_1483)
);

AND2x2_ASAP7_75t_L g1484 ( 
.A(n_1215),
.B(n_120),
.Y(n_1484)
);

NAND2xp5_ASAP7_75t_L g1485 ( 
.A(n_1239),
.B(n_1324),
.Y(n_1485)
);

BUFx10_ASAP7_75t_L g1486 ( 
.A(n_1247),
.Y(n_1486)
);

AO31x2_ASAP7_75t_L g1487 ( 
.A1(n_1295),
.A2(n_121),
.A3(n_122),
.B(n_123),
.Y(n_1487)
);

XNOR2xp5_ASAP7_75t_L g1488 ( 
.A(n_1256),
.B(n_414),
.Y(n_1488)
);

AND2x2_ASAP7_75t_L g1489 ( 
.A(n_1211),
.B(n_122),
.Y(n_1489)
);

AOI31xp33_ASAP7_75t_L g1490 ( 
.A1(n_1423),
.A2(n_1225),
.A3(n_1213),
.B(n_1236),
.Y(n_1490)
);

INVx4_ASAP7_75t_L g1491 ( 
.A(n_1348),
.Y(n_1491)
);

INVx1_ASAP7_75t_L g1492 ( 
.A(n_1351),
.Y(n_1492)
);

NAND3xp33_ASAP7_75t_SL g1493 ( 
.A(n_1438),
.B(n_1208),
.C(n_1232),
.Y(n_1493)
);

BUFx6f_ASAP7_75t_L g1494 ( 
.A(n_1361),
.Y(n_1494)
);

O2A1O1Ixp33_ASAP7_75t_L g1495 ( 
.A1(n_1380),
.A2(n_1231),
.B(n_1218),
.C(n_1295),
.Y(n_1495)
);

INVx1_ASAP7_75t_L g1496 ( 
.A(n_1357),
.Y(n_1496)
);

INVx2_ASAP7_75t_R g1497 ( 
.A(n_1416),
.Y(n_1497)
);

BUFx2_ASAP7_75t_L g1498 ( 
.A(n_1462),
.Y(n_1498)
);

AOI21xp5_ASAP7_75t_L g1499 ( 
.A1(n_1335),
.A2(n_1284),
.B(n_1192),
.Y(n_1499)
);

AOI21xp5_ASAP7_75t_L g1500 ( 
.A1(n_1384),
.A2(n_1181),
.B(n_1290),
.Y(n_1500)
);

OAI21x1_ASAP7_75t_L g1501 ( 
.A1(n_1454),
.A2(n_1269),
.B(n_1259),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_1376),
.Y(n_1502)
);

INVx1_ASAP7_75t_L g1503 ( 
.A(n_1385),
.Y(n_1503)
);

A2O1A1Ixp33_ASAP7_75t_L g1504 ( 
.A1(n_1456),
.A2(n_1205),
.B(n_1317),
.C(n_1292),
.Y(n_1504)
);

OAI22xp5_ASAP7_75t_L g1505 ( 
.A1(n_1418),
.A2(n_1180),
.B1(n_1324),
.B2(n_1317),
.Y(n_1505)
);

A2O1A1Ixp33_ASAP7_75t_L g1506 ( 
.A1(n_1377),
.A2(n_1292),
.B(n_1247),
.C(n_1323),
.Y(n_1506)
);

BUFx3_ASAP7_75t_L g1507 ( 
.A(n_1354),
.Y(n_1507)
);

BUFx12f_ASAP7_75t_L g1508 ( 
.A(n_1469),
.Y(n_1508)
);

A2O1A1Ixp33_ASAP7_75t_L g1509 ( 
.A1(n_1409),
.A2(n_1323),
.B(n_1181),
.C(n_1269),
.Y(n_1509)
);

OAI21x1_ASAP7_75t_L g1510 ( 
.A1(n_1360),
.A2(n_1323),
.B(n_1293),
.Y(n_1510)
);

OAI21xp5_ASAP7_75t_L g1511 ( 
.A1(n_1378),
.A2(n_1231),
.B(n_1218),
.Y(n_1511)
);

INVx2_ASAP7_75t_SL g1512 ( 
.A(n_1342),
.Y(n_1512)
);

AO31x2_ASAP7_75t_L g1513 ( 
.A1(n_1365),
.A2(n_1311),
.A3(n_1307),
.B(n_478),
.Y(n_1513)
);

NOR2xp67_ASAP7_75t_L g1514 ( 
.A(n_1374),
.B(n_1381),
.Y(n_1514)
);

AO21x1_ASAP7_75t_L g1515 ( 
.A1(n_1350),
.A2(n_123),
.B(n_124),
.Y(n_1515)
);

AOI21x1_ASAP7_75t_L g1516 ( 
.A1(n_1338),
.A2(n_1166),
.B(n_418),
.Y(n_1516)
);

NOR2xp33_ASAP7_75t_L g1517 ( 
.A(n_1412),
.B(n_1279),
.Y(n_1517)
);

CKINVDCx11_ASAP7_75t_R g1518 ( 
.A(n_1486),
.Y(n_1518)
);

AOI22xp5_ASAP7_75t_L g1519 ( 
.A1(n_1402),
.A2(n_1260),
.B1(n_125),
.B2(n_126),
.Y(n_1519)
);

AO32x2_ASAP7_75t_L g1520 ( 
.A1(n_1453),
.A2(n_124),
.A3(n_125),
.B1(n_126),
.B2(n_127),
.Y(n_1520)
);

AOI22xp5_ASAP7_75t_L g1521 ( 
.A1(n_1349),
.A2(n_128),
.B1(n_129),
.B2(n_130),
.Y(n_1521)
);

INVx2_ASAP7_75t_SL g1522 ( 
.A(n_1417),
.Y(n_1522)
);

OAI22xp5_ASAP7_75t_L g1523 ( 
.A1(n_1480),
.A2(n_131),
.B1(n_132),
.B2(n_134),
.Y(n_1523)
);

CKINVDCx20_ASAP7_75t_R g1524 ( 
.A(n_1488),
.Y(n_1524)
);

AOI221xp5_ASAP7_75t_L g1525 ( 
.A1(n_1390),
.A2(n_132),
.B1(n_134),
.B2(n_135),
.C(n_136),
.Y(n_1525)
);

AOI221x1_ASAP7_75t_L g1526 ( 
.A1(n_1428),
.A2(n_135),
.B1(n_136),
.B2(n_137),
.C(n_138),
.Y(n_1526)
);

BUFx6f_ASAP7_75t_L g1527 ( 
.A(n_1348),
.Y(n_1527)
);

NOR2xp33_ASAP7_75t_L g1528 ( 
.A(n_1394),
.B(n_416),
.Y(n_1528)
);

AND2x2_ASAP7_75t_L g1529 ( 
.A(n_1419),
.B(n_137),
.Y(n_1529)
);

INVx1_ASAP7_75t_L g1530 ( 
.A(n_1439),
.Y(n_1530)
);

A2O1A1Ixp33_ASAP7_75t_L g1531 ( 
.A1(n_1436),
.A2(n_138),
.B(n_139),
.C(n_140),
.Y(n_1531)
);

INVxp67_ASAP7_75t_L g1532 ( 
.A(n_1442),
.Y(n_1532)
);

OAI21xp5_ASAP7_75t_L g1533 ( 
.A1(n_1334),
.A2(n_139),
.B(n_140),
.Y(n_1533)
);

OAI21x1_ASAP7_75t_L g1534 ( 
.A1(n_1410),
.A2(n_476),
.B(n_475),
.Y(n_1534)
);

BUFx10_ASAP7_75t_L g1535 ( 
.A(n_1355),
.Y(n_1535)
);

AOI21x1_ASAP7_75t_SL g1536 ( 
.A1(n_1367),
.A2(n_1411),
.B(n_1489),
.Y(n_1536)
);

O2A1O1Ixp33_ASAP7_75t_L g1537 ( 
.A1(n_1461),
.A2(n_1398),
.B(n_1358),
.C(n_1424),
.Y(n_1537)
);

AOI21xp33_ASAP7_75t_L g1538 ( 
.A1(n_1336),
.A2(n_141),
.B(n_142),
.Y(n_1538)
);

AOI21xp5_ASAP7_75t_L g1539 ( 
.A1(n_1389),
.A2(n_474),
.B(n_473),
.Y(n_1539)
);

NOR2xp33_ASAP7_75t_L g1540 ( 
.A(n_1405),
.B(n_419),
.Y(n_1540)
);

INVx2_ASAP7_75t_L g1541 ( 
.A(n_1446),
.Y(n_1541)
);

O2A1O1Ixp33_ASAP7_75t_SL g1542 ( 
.A1(n_1414),
.A2(n_141),
.B(n_142),
.C(n_143),
.Y(n_1542)
);

OAI21x1_ASAP7_75t_L g1543 ( 
.A1(n_1422),
.A2(n_467),
.B(n_466),
.Y(n_1543)
);

AOI21x1_ASAP7_75t_L g1544 ( 
.A1(n_1345),
.A2(n_465),
.B(n_463),
.Y(n_1544)
);

NAND2xp5_ASAP7_75t_L g1545 ( 
.A(n_1472),
.B(n_144),
.Y(n_1545)
);

AOI22xp5_ASAP7_75t_L g1546 ( 
.A1(n_1485),
.A2(n_144),
.B1(n_145),
.B2(n_146),
.Y(n_1546)
);

AOI21xp5_ASAP7_75t_L g1547 ( 
.A1(n_1471),
.A2(n_461),
.B(n_459),
.Y(n_1547)
);

AOI21x1_ASAP7_75t_L g1548 ( 
.A1(n_1364),
.A2(n_439),
.B(n_457),
.Y(n_1548)
);

A2O1A1Ixp33_ASAP7_75t_L g1549 ( 
.A1(n_1403),
.A2(n_145),
.B(n_146),
.C(n_147),
.Y(n_1549)
);

BUFx4_ASAP7_75t_SL g1550 ( 
.A(n_1369),
.Y(n_1550)
);

INVx2_ASAP7_75t_L g1551 ( 
.A(n_1450),
.Y(n_1551)
);

AOI21xp5_ASAP7_75t_L g1552 ( 
.A1(n_1443),
.A2(n_458),
.B(n_455),
.Y(n_1552)
);

AND2x2_ASAP7_75t_L g1553 ( 
.A(n_1340),
.B(n_148),
.Y(n_1553)
);

NAND2xp5_ASAP7_75t_L g1554 ( 
.A(n_1344),
.B(n_149),
.Y(n_1554)
);

OAI21x1_ASAP7_75t_L g1555 ( 
.A1(n_1425),
.A2(n_454),
.B(n_452),
.Y(n_1555)
);

AO32x2_ASAP7_75t_L g1556 ( 
.A1(n_1432),
.A2(n_149),
.A3(n_150),
.B1(n_151),
.B2(n_152),
.Y(n_1556)
);

BUFx2_ASAP7_75t_L g1557 ( 
.A(n_1444),
.Y(n_1557)
);

AND2x4_ASAP7_75t_L g1558 ( 
.A(n_1356),
.B(n_420),
.Y(n_1558)
);

OAI22xp5_ASAP7_75t_L g1559 ( 
.A1(n_1477),
.A2(n_1455),
.B1(n_1476),
.B2(n_1406),
.Y(n_1559)
);

AO21x2_ASAP7_75t_L g1560 ( 
.A1(n_1343),
.A2(n_450),
.B(n_448),
.Y(n_1560)
);

AOI21xp5_ASAP7_75t_L g1561 ( 
.A1(n_1449),
.A2(n_447),
.B(n_446),
.Y(n_1561)
);

AOI21xp5_ASAP7_75t_L g1562 ( 
.A1(n_1337),
.A2(n_445),
.B(n_443),
.Y(n_1562)
);

A2O1A1Ixp33_ASAP7_75t_L g1563 ( 
.A1(n_1407),
.A2(n_151),
.B(n_152),
.C(n_153),
.Y(n_1563)
);

INVx1_ASAP7_75t_L g1564 ( 
.A(n_1430),
.Y(n_1564)
);

AOI21xp5_ASAP7_75t_L g1565 ( 
.A1(n_1352),
.A2(n_442),
.B(n_441),
.Y(n_1565)
);

BUFx6f_ASAP7_75t_L g1566 ( 
.A(n_1348),
.Y(n_1566)
);

OR2x2_ASAP7_75t_L g1567 ( 
.A(n_1347),
.B(n_153),
.Y(n_1567)
);

CKINVDCx20_ASAP7_75t_R g1568 ( 
.A(n_1486),
.Y(n_1568)
);

OAI21x1_ASAP7_75t_L g1569 ( 
.A1(n_1431),
.A2(n_440),
.B(n_438),
.Y(n_1569)
);

OAI21x1_ASAP7_75t_L g1570 ( 
.A1(n_1435),
.A2(n_434),
.B(n_433),
.Y(n_1570)
);

INVx1_ASAP7_75t_L g1571 ( 
.A(n_1433),
.Y(n_1571)
);

BUFx4f_ASAP7_75t_L g1572 ( 
.A(n_1359),
.Y(n_1572)
);

AND2x2_ASAP7_75t_L g1573 ( 
.A(n_1484),
.B(n_155),
.Y(n_1573)
);

NOR2xp67_ASAP7_75t_SL g1574 ( 
.A(n_1420),
.B(n_156),
.Y(n_1574)
);

INVx5_ASAP7_75t_L g1575 ( 
.A(n_1368),
.Y(n_1575)
);

NAND2xp5_ASAP7_75t_L g1576 ( 
.A(n_1346),
.B(n_157),
.Y(n_1576)
);

NAND2xp5_ASAP7_75t_L g1577 ( 
.A(n_1451),
.B(n_157),
.Y(n_1577)
);

AOI21xp5_ASAP7_75t_L g1578 ( 
.A1(n_1371),
.A2(n_432),
.B(n_431),
.Y(n_1578)
);

NOR2x1_ASAP7_75t_SL g1579 ( 
.A(n_1359),
.B(n_429),
.Y(n_1579)
);

INVx1_ASAP7_75t_SL g1580 ( 
.A(n_1388),
.Y(n_1580)
);

AOI21xp5_ASAP7_75t_L g1581 ( 
.A1(n_1392),
.A2(n_428),
.B(n_427),
.Y(n_1581)
);

BUFx3_ASAP7_75t_L g1582 ( 
.A(n_1368),
.Y(n_1582)
);

BUFx3_ASAP7_75t_L g1583 ( 
.A(n_1368),
.Y(n_1583)
);

OAI21x1_ASAP7_75t_L g1584 ( 
.A1(n_1408),
.A2(n_425),
.B(n_424),
.Y(n_1584)
);

AND2x4_ASAP7_75t_L g1585 ( 
.A(n_1363),
.B(n_421),
.Y(n_1585)
);

NAND2xp5_ASAP7_75t_L g1586 ( 
.A(n_1452),
.B(n_158),
.Y(n_1586)
);

OAI21xp5_ASAP7_75t_L g1587 ( 
.A1(n_1475),
.A2(n_161),
.B(n_163),
.Y(n_1587)
);

NAND3xp33_ASAP7_75t_L g1588 ( 
.A(n_1429),
.B(n_164),
.C(n_165),
.Y(n_1588)
);

NAND2xp5_ASAP7_75t_L g1589 ( 
.A(n_1473),
.B(n_167),
.Y(n_1589)
);

OA21x2_ASAP7_75t_L g1590 ( 
.A1(n_1379),
.A2(n_168),
.B(n_170),
.Y(n_1590)
);

AOI21x1_ASAP7_75t_L g1591 ( 
.A1(n_1383),
.A2(n_168),
.B(n_170),
.Y(n_1591)
);

INVxp67_ASAP7_75t_SL g1592 ( 
.A(n_1465),
.Y(n_1592)
);

NAND2xp5_ASAP7_75t_L g1593 ( 
.A(n_1474),
.B(n_171),
.Y(n_1593)
);

INVxp67_ASAP7_75t_SL g1594 ( 
.A(n_1466),
.Y(n_1594)
);

AOI21xp5_ASAP7_75t_L g1595 ( 
.A1(n_1421),
.A2(n_171),
.B(n_172),
.Y(n_1595)
);

NAND2xp5_ASAP7_75t_L g1596 ( 
.A(n_1481),
.B(n_172),
.Y(n_1596)
);

INVx6_ASAP7_75t_L g1597 ( 
.A(n_1393),
.Y(n_1597)
);

BUFx6f_ASAP7_75t_L g1598 ( 
.A(n_1393),
.Y(n_1598)
);

OR2x2_ASAP7_75t_L g1599 ( 
.A(n_1415),
.B(n_1404),
.Y(n_1599)
);

INVx4_ASAP7_75t_L g1600 ( 
.A(n_1393),
.Y(n_1600)
);

AOI21xp5_ASAP7_75t_L g1601 ( 
.A1(n_1426),
.A2(n_173),
.B(n_174),
.Y(n_1601)
);

A2O1A1Ixp33_ASAP7_75t_L g1602 ( 
.A1(n_1463),
.A2(n_174),
.B(n_175),
.C(n_177),
.Y(n_1602)
);

BUFx4f_ASAP7_75t_L g1603 ( 
.A(n_1404),
.Y(n_1603)
);

AND2x6_ASAP7_75t_L g1604 ( 
.A(n_1339),
.B(n_175),
.Y(n_1604)
);

BUFx3_ASAP7_75t_L g1605 ( 
.A(n_1434),
.Y(n_1605)
);

OAI22xp5_ASAP7_75t_L g1606 ( 
.A1(n_1366),
.A2(n_179),
.B1(n_180),
.B2(n_182),
.Y(n_1606)
);

OAI22x1_ASAP7_75t_L g1607 ( 
.A1(n_1459),
.A2(n_182),
.B1(n_183),
.B2(n_184),
.Y(n_1607)
);

BUFx2_ASAP7_75t_L g1608 ( 
.A(n_1470),
.Y(n_1608)
);

AND2x4_ASAP7_75t_L g1609 ( 
.A(n_1363),
.B(n_184),
.Y(n_1609)
);

AND2x2_ASAP7_75t_L g1610 ( 
.A(n_1448),
.B(n_185),
.Y(n_1610)
);

BUFx2_ASAP7_75t_L g1611 ( 
.A(n_1482),
.Y(n_1611)
);

OAI21xp33_ASAP7_75t_SL g1612 ( 
.A1(n_1445),
.A2(n_185),
.B(n_186),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1457),
.Y(n_1613)
);

AND2x2_ASAP7_75t_L g1614 ( 
.A(n_1441),
.B(n_187),
.Y(n_1614)
);

CKINVDCx5p33_ASAP7_75t_R g1615 ( 
.A(n_1369),
.Y(n_1615)
);

OAI21x1_ASAP7_75t_L g1616 ( 
.A1(n_1362),
.A2(n_187),
.B(n_188),
.Y(n_1616)
);

NAND2xp5_ASAP7_75t_SL g1617 ( 
.A(n_1339),
.B(n_188),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_1457),
.Y(n_1618)
);

AOI21xp5_ASAP7_75t_L g1619 ( 
.A1(n_1440),
.A2(n_219),
.B(n_190),
.Y(n_1619)
);

NOR2xp33_ASAP7_75t_L g1620 ( 
.A(n_1447),
.B(n_189),
.Y(n_1620)
);

NOR2xp33_ASAP7_75t_SL g1621 ( 
.A(n_1370),
.B(n_190),
.Y(n_1621)
);

AOI21xp5_ASAP7_75t_L g1622 ( 
.A1(n_1479),
.A2(n_219),
.B(n_192),
.Y(n_1622)
);

INVx5_ASAP7_75t_L g1623 ( 
.A(n_1434),
.Y(n_1623)
);

OAI21x1_ASAP7_75t_L g1624 ( 
.A1(n_1382),
.A2(n_191),
.B(n_193),
.Y(n_1624)
);

AOI21xp5_ASAP7_75t_L g1625 ( 
.A1(n_1460),
.A2(n_218),
.B(n_195),
.Y(n_1625)
);

AOI22xp33_ASAP7_75t_L g1626 ( 
.A1(n_1493),
.A2(n_1464),
.B1(n_1427),
.B2(n_1395),
.Y(n_1626)
);

AOI22xp33_ASAP7_75t_L g1627 ( 
.A1(n_1533),
.A2(n_1341),
.B1(n_1397),
.B2(n_1437),
.Y(n_1627)
);

CKINVDCx6p67_ASAP7_75t_R g1628 ( 
.A(n_1508),
.Y(n_1628)
);

OAI22xp5_ASAP7_75t_L g1629 ( 
.A1(n_1572),
.A2(n_1397),
.B1(n_1386),
.B2(n_1373),
.Y(n_1629)
);

INVx2_ASAP7_75t_SL g1630 ( 
.A(n_1494),
.Y(n_1630)
);

AOI22xp33_ASAP7_75t_SL g1631 ( 
.A1(n_1621),
.A2(n_1437),
.B1(n_1353),
.B2(n_1483),
.Y(n_1631)
);

BUFx2_ASAP7_75t_SL g1632 ( 
.A(n_1568),
.Y(n_1632)
);

CKINVDCx20_ASAP7_75t_R g1633 ( 
.A(n_1518),
.Y(n_1633)
);

AOI22xp33_ASAP7_75t_L g1634 ( 
.A1(n_1519),
.A2(n_1437),
.B1(n_1375),
.B2(n_1399),
.Y(n_1634)
);

NAND2xp5_ASAP7_75t_L g1635 ( 
.A(n_1580),
.B(n_1487),
.Y(n_1635)
);

NAND2xp5_ASAP7_75t_L g1636 ( 
.A(n_1564),
.B(n_1487),
.Y(n_1636)
);

BUFx2_ASAP7_75t_L g1637 ( 
.A(n_1498),
.Y(n_1637)
);

AOI22xp33_ASAP7_75t_L g1638 ( 
.A1(n_1525),
.A2(n_1437),
.B1(n_1391),
.B2(n_1401),
.Y(n_1638)
);

INVx2_ASAP7_75t_L g1639 ( 
.A(n_1541),
.Y(n_1639)
);

AOI22xp33_ASAP7_75t_SL g1640 ( 
.A1(n_1606),
.A2(n_1387),
.B1(n_1457),
.B2(n_1413),
.Y(n_1640)
);

CKINVDCx5p33_ASAP7_75t_R g1641 ( 
.A(n_1494),
.Y(n_1641)
);

INVx3_ASAP7_75t_L g1642 ( 
.A(n_1598),
.Y(n_1642)
);

CKINVDCx20_ASAP7_75t_R g1643 ( 
.A(n_1524),
.Y(n_1643)
);

BUFx3_ASAP7_75t_L g1644 ( 
.A(n_1507),
.Y(n_1644)
);

INVx1_ASAP7_75t_L g1645 ( 
.A(n_1613),
.Y(n_1645)
);

AOI22xp33_ASAP7_75t_L g1646 ( 
.A1(n_1588),
.A2(n_1434),
.B1(n_1468),
.B2(n_1467),
.Y(n_1646)
);

INVx6_ASAP7_75t_L g1647 ( 
.A(n_1575),
.Y(n_1647)
);

BUFx3_ASAP7_75t_L g1648 ( 
.A(n_1582),
.Y(n_1648)
);

INVx6_ASAP7_75t_L g1649 ( 
.A(n_1575),
.Y(n_1649)
);

INVx1_ASAP7_75t_L g1650 ( 
.A(n_1492),
.Y(n_1650)
);

NAND2x1p5_ASAP7_75t_L g1651 ( 
.A(n_1575),
.B(n_1468),
.Y(n_1651)
);

AOI22xp33_ASAP7_75t_SL g1652 ( 
.A1(n_1604),
.A2(n_1413),
.B1(n_1372),
.B2(n_1467),
.Y(n_1652)
);

BUFx12f_ASAP7_75t_L g1653 ( 
.A(n_1615),
.Y(n_1653)
);

NAND2xp5_ASAP7_75t_L g1654 ( 
.A(n_1571),
.B(n_1372),
.Y(n_1654)
);

INVx5_ASAP7_75t_L g1655 ( 
.A(n_1604),
.Y(n_1655)
);

BUFx6f_ASAP7_75t_L g1656 ( 
.A(n_1527),
.Y(n_1656)
);

CKINVDCx11_ASAP7_75t_R g1657 ( 
.A(n_1535),
.Y(n_1657)
);

INVx2_ASAP7_75t_SL g1658 ( 
.A(n_1597),
.Y(n_1658)
);

AND2x2_ASAP7_75t_L g1659 ( 
.A(n_1573),
.B(n_1529),
.Y(n_1659)
);

INVx1_ASAP7_75t_L g1660 ( 
.A(n_1496),
.Y(n_1660)
);

BUFx3_ASAP7_75t_L g1661 ( 
.A(n_1583),
.Y(n_1661)
);

AOI22xp33_ASAP7_75t_SL g1662 ( 
.A1(n_1604),
.A2(n_1413),
.B1(n_1372),
.B2(n_1467),
.Y(n_1662)
);

BUFx3_ASAP7_75t_L g1663 ( 
.A(n_1605),
.Y(n_1663)
);

INVx3_ASAP7_75t_L g1664 ( 
.A(n_1598),
.Y(n_1664)
);

AOI22xp33_ASAP7_75t_L g1665 ( 
.A1(n_1515),
.A2(n_1468),
.B1(n_1458),
.B2(n_1478),
.Y(n_1665)
);

INVx1_ASAP7_75t_L g1666 ( 
.A(n_1502),
.Y(n_1666)
);

CKINVDCx11_ASAP7_75t_R g1667 ( 
.A(n_1527),
.Y(n_1667)
);

INVx1_ASAP7_75t_L g1668 ( 
.A(n_1503),
.Y(n_1668)
);

BUFx8_ASAP7_75t_L g1669 ( 
.A(n_1608),
.Y(n_1669)
);

BUFx10_ASAP7_75t_L g1670 ( 
.A(n_1517),
.Y(n_1670)
);

INVx1_ASAP7_75t_L g1671 ( 
.A(n_1530),
.Y(n_1671)
);

INVx6_ASAP7_75t_L g1672 ( 
.A(n_1623),
.Y(n_1672)
);

INVx1_ASAP7_75t_L g1673 ( 
.A(n_1618),
.Y(n_1673)
);

CKINVDCx20_ASAP7_75t_R g1674 ( 
.A(n_1505),
.Y(n_1674)
);

INVx6_ASAP7_75t_L g1675 ( 
.A(n_1623),
.Y(n_1675)
);

BUFx2_ASAP7_75t_SL g1676 ( 
.A(n_1514),
.Y(n_1676)
);

INVx1_ASAP7_75t_SL g1677 ( 
.A(n_1522),
.Y(n_1677)
);

AOI22xp33_ASAP7_75t_L g1678 ( 
.A1(n_1528),
.A2(n_1458),
.B1(n_1478),
.B2(n_1400),
.Y(n_1678)
);

AOI22xp33_ASAP7_75t_SL g1679 ( 
.A1(n_1511),
.A2(n_1579),
.B1(n_1603),
.B2(n_1500),
.Y(n_1679)
);

CKINVDCx20_ASAP7_75t_R g1680 ( 
.A(n_1532),
.Y(n_1680)
);

INVx6_ASAP7_75t_L g1681 ( 
.A(n_1623),
.Y(n_1681)
);

BUFx6f_ASAP7_75t_L g1682 ( 
.A(n_1566),
.Y(n_1682)
);

AOI22xp33_ASAP7_75t_SL g1683 ( 
.A1(n_1539),
.A2(n_1458),
.B1(n_1396),
.B2(n_196),
.Y(n_1683)
);

BUFx2_ASAP7_75t_R g1684 ( 
.A(n_1617),
.Y(n_1684)
);

BUFx2_ASAP7_75t_SL g1685 ( 
.A(n_1512),
.Y(n_1685)
);

AOI22xp33_ASAP7_75t_L g1686 ( 
.A1(n_1538),
.A2(n_194),
.B1(n_195),
.B2(n_196),
.Y(n_1686)
);

AOI22xp33_ASAP7_75t_L g1687 ( 
.A1(n_1620),
.A2(n_194),
.B1(n_197),
.B2(n_198),
.Y(n_1687)
);

AOI22xp33_ASAP7_75t_L g1688 ( 
.A1(n_1521),
.A2(n_197),
.B1(n_198),
.B2(n_199),
.Y(n_1688)
);

OAI22xp33_ASAP7_75t_L g1689 ( 
.A1(n_1490),
.A2(n_199),
.B1(n_200),
.B2(n_201),
.Y(n_1689)
);

INVx2_ASAP7_75t_L g1690 ( 
.A(n_1551),
.Y(n_1690)
);

AOI22xp33_ASAP7_75t_SL g1691 ( 
.A1(n_1552),
.A2(n_201),
.B1(n_202),
.B2(n_203),
.Y(n_1691)
);

BUFx2_ASAP7_75t_SL g1692 ( 
.A(n_1491),
.Y(n_1692)
);

AOI22xp33_ASAP7_75t_L g1693 ( 
.A1(n_1607),
.A2(n_202),
.B1(n_203),
.B2(n_204),
.Y(n_1693)
);

INVx4_ASAP7_75t_L g1694 ( 
.A(n_1566),
.Y(n_1694)
);

OAI21xp5_ASAP7_75t_SL g1695 ( 
.A1(n_1495),
.A2(n_205),
.B(n_208),
.Y(n_1695)
);

INVx1_ASAP7_75t_SL g1696 ( 
.A(n_1599),
.Y(n_1696)
);

BUFx6f_ASAP7_75t_L g1697 ( 
.A(n_1597),
.Y(n_1697)
);

INVx5_ASAP7_75t_L g1698 ( 
.A(n_1600),
.Y(n_1698)
);

AOI22xp33_ASAP7_75t_L g1699 ( 
.A1(n_1574),
.A2(n_208),
.B1(n_209),
.B2(n_211),
.Y(n_1699)
);

CKINVDCx11_ASAP7_75t_R g1700 ( 
.A(n_1609),
.Y(n_1700)
);

AOI22xp33_ASAP7_75t_L g1701 ( 
.A1(n_1610),
.A2(n_209),
.B1(n_212),
.B2(n_213),
.Y(n_1701)
);

INVx6_ASAP7_75t_L g1702 ( 
.A(n_1585),
.Y(n_1702)
);

INVx11_ASAP7_75t_L g1703 ( 
.A(n_1550),
.Y(n_1703)
);

INVx2_ASAP7_75t_L g1704 ( 
.A(n_1611),
.Y(n_1704)
);

INVx1_ASAP7_75t_SL g1705 ( 
.A(n_1497),
.Y(n_1705)
);

CKINVDCx11_ASAP7_75t_R g1706 ( 
.A(n_1558),
.Y(n_1706)
);

BUFx3_ASAP7_75t_L g1707 ( 
.A(n_1545),
.Y(n_1707)
);

INVx1_ASAP7_75t_SL g1708 ( 
.A(n_1553),
.Y(n_1708)
);

AOI22xp33_ASAP7_75t_L g1709 ( 
.A1(n_1587),
.A2(n_212),
.B1(n_213),
.B2(n_214),
.Y(n_1709)
);

INVx1_ASAP7_75t_L g1710 ( 
.A(n_1611),
.Y(n_1710)
);

INVx1_ASAP7_75t_L g1711 ( 
.A(n_1592),
.Y(n_1711)
);

OAI22xp33_ASAP7_75t_L g1712 ( 
.A1(n_1526),
.A2(n_214),
.B1(n_215),
.B2(n_216),
.Y(n_1712)
);

INVx8_ASAP7_75t_L g1713 ( 
.A(n_1614),
.Y(n_1713)
);

INVx1_ASAP7_75t_L g1714 ( 
.A(n_1594),
.Y(n_1714)
);

AOI22x1_ASAP7_75t_SL g1715 ( 
.A1(n_1556),
.A2(n_215),
.B1(n_216),
.B2(n_217),
.Y(n_1715)
);

INVx1_ASAP7_75t_SL g1716 ( 
.A(n_1577),
.Y(n_1716)
);

BUFx10_ASAP7_75t_L g1717 ( 
.A(n_1540),
.Y(n_1717)
);

BUFx6f_ASAP7_75t_L g1718 ( 
.A(n_1501),
.Y(n_1718)
);

NAND2xp5_ASAP7_75t_L g1719 ( 
.A(n_1509),
.B(n_217),
.Y(n_1719)
);

INVx1_ASAP7_75t_L g1720 ( 
.A(n_1650),
.Y(n_1720)
);

AND2x2_ASAP7_75t_L g1721 ( 
.A(n_1704),
.B(n_1557),
.Y(n_1721)
);

INVx1_ASAP7_75t_L g1722 ( 
.A(n_1660),
.Y(n_1722)
);

HB1xp67_ASAP7_75t_L g1723 ( 
.A(n_1711),
.Y(n_1723)
);

INVx1_ASAP7_75t_L g1724 ( 
.A(n_1666),
.Y(n_1724)
);

OAI22xp5_ASAP7_75t_L g1725 ( 
.A1(n_1626),
.A2(n_1504),
.B1(n_1549),
.B2(n_1506),
.Y(n_1725)
);

INVx1_ASAP7_75t_L g1726 ( 
.A(n_1645),
.Y(n_1726)
);

HB1xp67_ASAP7_75t_L g1727 ( 
.A(n_1714),
.Y(n_1727)
);

AND2x2_ASAP7_75t_L g1728 ( 
.A(n_1668),
.B(n_1557),
.Y(n_1728)
);

HB1xp67_ASAP7_75t_L g1729 ( 
.A(n_1710),
.Y(n_1729)
);

HB1xp67_ASAP7_75t_L g1730 ( 
.A(n_1635),
.Y(n_1730)
);

NOR2xp33_ASAP7_75t_L g1731 ( 
.A(n_1680),
.B(n_1586),
.Y(n_1731)
);

INVx1_ASAP7_75t_L g1732 ( 
.A(n_1673),
.Y(n_1732)
);

AOI21x1_ASAP7_75t_L g1733 ( 
.A1(n_1636),
.A2(n_1591),
.B(n_1544),
.Y(n_1733)
);

AND2x2_ASAP7_75t_L g1734 ( 
.A(n_1671),
.B(n_1590),
.Y(n_1734)
);

AOI22xp33_ASAP7_75t_L g1735 ( 
.A1(n_1689),
.A2(n_1561),
.B1(n_1622),
.B2(n_1619),
.Y(n_1735)
);

INVx1_ASAP7_75t_L g1736 ( 
.A(n_1654),
.Y(n_1736)
);

INVx6_ASAP7_75t_L g1737 ( 
.A(n_1669),
.Y(n_1737)
);

NAND2xp5_ASAP7_75t_L g1738 ( 
.A(n_1696),
.B(n_1716),
.Y(n_1738)
);

NAND2xp5_ASAP7_75t_L g1739 ( 
.A(n_1639),
.B(n_1690),
.Y(n_1739)
);

INVx2_ASAP7_75t_L g1740 ( 
.A(n_1718),
.Y(n_1740)
);

INVx1_ASAP7_75t_L g1741 ( 
.A(n_1718),
.Y(n_1741)
);

OR2x6_ASAP7_75t_L g1742 ( 
.A(n_1718),
.B(n_1499),
.Y(n_1742)
);

INVx1_ASAP7_75t_L g1743 ( 
.A(n_1705),
.Y(n_1743)
);

INVx1_ASAP7_75t_L g1744 ( 
.A(n_1637),
.Y(n_1744)
);

OAI22xp5_ASAP7_75t_L g1745 ( 
.A1(n_1695),
.A2(n_1546),
.B1(n_1531),
.B2(n_1563),
.Y(n_1745)
);

INVx3_ASAP7_75t_L g1746 ( 
.A(n_1655),
.Y(n_1746)
);

BUFx3_ASAP7_75t_L g1747 ( 
.A(n_1669),
.Y(n_1747)
);

BUFx6f_ASAP7_75t_L g1748 ( 
.A(n_1655),
.Y(n_1748)
);

AND2x2_ASAP7_75t_L g1749 ( 
.A(n_1652),
.B(n_1662),
.Y(n_1749)
);

INVx1_ASAP7_75t_L g1750 ( 
.A(n_1715),
.Y(n_1750)
);

INVx1_ASAP7_75t_L g1751 ( 
.A(n_1640),
.Y(n_1751)
);

INVx1_ASAP7_75t_L g1752 ( 
.A(n_1678),
.Y(n_1752)
);

INVx2_ASAP7_75t_L g1753 ( 
.A(n_1647),
.Y(n_1753)
);

INVx1_ASAP7_75t_L g1754 ( 
.A(n_1715),
.Y(n_1754)
);

INVx2_ASAP7_75t_SL g1755 ( 
.A(n_1647),
.Y(n_1755)
);

AOI22xp33_ASAP7_75t_L g1756 ( 
.A1(n_1712),
.A2(n_1601),
.B1(n_1595),
.B2(n_1625),
.Y(n_1756)
);

INVx2_ASAP7_75t_L g1757 ( 
.A(n_1649),
.Y(n_1757)
);

INVx1_ASAP7_75t_L g1758 ( 
.A(n_1676),
.Y(n_1758)
);

INVx1_ASAP7_75t_L g1759 ( 
.A(n_1685),
.Y(n_1759)
);

INVx4_ASAP7_75t_L g1760 ( 
.A(n_1655),
.Y(n_1760)
);

INVx1_ASAP7_75t_L g1761 ( 
.A(n_1665),
.Y(n_1761)
);

INVx1_ASAP7_75t_L g1762 ( 
.A(n_1679),
.Y(n_1762)
);

INVx2_ASAP7_75t_L g1763 ( 
.A(n_1649),
.Y(n_1763)
);

INVx1_ASAP7_75t_L g1764 ( 
.A(n_1719),
.Y(n_1764)
);

HB1xp67_ASAP7_75t_L g1765 ( 
.A(n_1707),
.Y(n_1765)
);

INVx1_ASAP7_75t_L g1766 ( 
.A(n_1726),
.Y(n_1766)
);

INVx2_ASAP7_75t_L g1767 ( 
.A(n_1726),
.Y(n_1767)
);

HB1xp67_ASAP7_75t_L g1768 ( 
.A(n_1729),
.Y(n_1768)
);

INVx3_ASAP7_75t_L g1769 ( 
.A(n_1740),
.Y(n_1769)
);

BUFx3_ASAP7_75t_L g1770 ( 
.A(n_1748),
.Y(n_1770)
);

HB1xp67_ASAP7_75t_L g1771 ( 
.A(n_1734),
.Y(n_1771)
);

AOI22xp33_ASAP7_75t_L g1772 ( 
.A1(n_1745),
.A2(n_1687),
.B1(n_1688),
.B2(n_1709),
.Y(n_1772)
);

BUFx3_ASAP7_75t_L g1773 ( 
.A(n_1748),
.Y(n_1773)
);

BUFx2_ASAP7_75t_L g1774 ( 
.A(n_1740),
.Y(n_1774)
);

HB1xp67_ASAP7_75t_L g1775 ( 
.A(n_1734),
.Y(n_1775)
);

INVx2_ASAP7_75t_L g1776 ( 
.A(n_1732),
.Y(n_1776)
);

AND2x2_ASAP7_75t_L g1777 ( 
.A(n_1728),
.B(n_1659),
.Y(n_1777)
);

AND2x2_ASAP7_75t_L g1778 ( 
.A(n_1728),
.B(n_1736),
.Y(n_1778)
);

INVx1_ASAP7_75t_L g1779 ( 
.A(n_1720),
.Y(n_1779)
);

OAI21x1_ASAP7_75t_L g1780 ( 
.A1(n_1733),
.A2(n_1516),
.B(n_1548),
.Y(n_1780)
);

AO21x2_ASAP7_75t_L g1781 ( 
.A1(n_1751),
.A2(n_1542),
.B(n_1624),
.Y(n_1781)
);

AND2x2_ASAP7_75t_L g1782 ( 
.A(n_1721),
.B(n_1708),
.Y(n_1782)
);

AO21x2_ASAP7_75t_L g1783 ( 
.A1(n_1751),
.A2(n_1602),
.B(n_1616),
.Y(n_1783)
);

AOI22xp33_ASAP7_75t_L g1784 ( 
.A1(n_1750),
.A2(n_1691),
.B1(n_1693),
.B2(n_1701),
.Y(n_1784)
);

AND2x4_ASAP7_75t_L g1785 ( 
.A(n_1741),
.B(n_1510),
.Y(n_1785)
);

INVx1_ASAP7_75t_L g1786 ( 
.A(n_1722),
.Y(n_1786)
);

OR2x2_ASAP7_75t_L g1787 ( 
.A(n_1730),
.B(n_1723),
.Y(n_1787)
);

INVx1_ASAP7_75t_L g1788 ( 
.A(n_1724),
.Y(n_1788)
);

AND2x2_ASAP7_75t_L g1789 ( 
.A(n_1771),
.B(n_1749),
.Y(n_1789)
);

AND2x2_ASAP7_75t_L g1790 ( 
.A(n_1771),
.B(n_1749),
.Y(n_1790)
);

INVx2_ASAP7_75t_L g1791 ( 
.A(n_1776),
.Y(n_1791)
);

INVx1_ASAP7_75t_L g1792 ( 
.A(n_1766),
.Y(n_1792)
);

AND2x4_ASAP7_75t_L g1793 ( 
.A(n_1770),
.B(n_1773),
.Y(n_1793)
);

INVx2_ASAP7_75t_L g1794 ( 
.A(n_1776),
.Y(n_1794)
);

BUFx12f_ASAP7_75t_L g1795 ( 
.A(n_1782),
.Y(n_1795)
);

INVx1_ASAP7_75t_L g1796 ( 
.A(n_1776),
.Y(n_1796)
);

NAND2xp5_ASAP7_75t_L g1797 ( 
.A(n_1782),
.B(n_1743),
.Y(n_1797)
);

BUFx6f_ASAP7_75t_L g1798 ( 
.A(n_1770),
.Y(n_1798)
);

BUFx6f_ASAP7_75t_L g1799 ( 
.A(n_1770),
.Y(n_1799)
);

AND2x2_ASAP7_75t_L g1800 ( 
.A(n_1775),
.B(n_1744),
.Y(n_1800)
);

AND2x2_ASAP7_75t_L g1801 ( 
.A(n_1775),
.B(n_1765),
.Y(n_1801)
);

INVxp67_ASAP7_75t_L g1802 ( 
.A(n_1768),
.Y(n_1802)
);

INVx1_ASAP7_75t_L g1803 ( 
.A(n_1776),
.Y(n_1803)
);

AND2x2_ASAP7_75t_L g1804 ( 
.A(n_1778),
.B(n_1727),
.Y(n_1804)
);

INVx1_ASAP7_75t_L g1805 ( 
.A(n_1767),
.Y(n_1805)
);

AO31x2_ASAP7_75t_L g1806 ( 
.A1(n_1774),
.A2(n_1761),
.A3(n_1752),
.B(n_1760),
.Y(n_1806)
);

INVx2_ASAP7_75t_L g1807 ( 
.A(n_1767),
.Y(n_1807)
);

OR2x2_ASAP7_75t_L g1808 ( 
.A(n_1787),
.B(n_1752),
.Y(n_1808)
);

AND2x2_ASAP7_75t_L g1809 ( 
.A(n_1778),
.B(n_1742),
.Y(n_1809)
);

AND2x2_ASAP7_75t_L g1810 ( 
.A(n_1789),
.B(n_1777),
.Y(n_1810)
);

INVx4_ASAP7_75t_L g1811 ( 
.A(n_1798),
.Y(n_1811)
);

BUFx2_ASAP7_75t_L g1812 ( 
.A(n_1795),
.Y(n_1812)
);

INVx1_ASAP7_75t_L g1813 ( 
.A(n_1792),
.Y(n_1813)
);

AND2x4_ASAP7_75t_L g1814 ( 
.A(n_1793),
.B(n_1770),
.Y(n_1814)
);

INVx1_ASAP7_75t_L g1815 ( 
.A(n_1808),
.Y(n_1815)
);

NAND2xp5_ASAP7_75t_L g1816 ( 
.A(n_1797),
.B(n_1782),
.Y(n_1816)
);

INVx1_ASAP7_75t_L g1817 ( 
.A(n_1808),
.Y(n_1817)
);

AND2x2_ASAP7_75t_L g1818 ( 
.A(n_1789),
.B(n_1777),
.Y(n_1818)
);

OR2x2_ASAP7_75t_L g1819 ( 
.A(n_1790),
.B(n_1801),
.Y(n_1819)
);

INVx1_ASAP7_75t_L g1820 ( 
.A(n_1813),
.Y(n_1820)
);

INVx5_ASAP7_75t_SL g1821 ( 
.A(n_1814),
.Y(n_1821)
);

INVx1_ASAP7_75t_L g1822 ( 
.A(n_1810),
.Y(n_1822)
);

INVx2_ASAP7_75t_L g1823 ( 
.A(n_1810),
.Y(n_1823)
);

INVx1_ASAP7_75t_L g1824 ( 
.A(n_1818),
.Y(n_1824)
);

AND2x2_ASAP7_75t_L g1825 ( 
.A(n_1818),
.B(n_1790),
.Y(n_1825)
);

AND2x2_ASAP7_75t_L g1826 ( 
.A(n_1821),
.B(n_1814),
.Y(n_1826)
);

INVx1_ASAP7_75t_L g1827 ( 
.A(n_1820),
.Y(n_1827)
);

AND2x2_ASAP7_75t_L g1828 ( 
.A(n_1821),
.B(n_1814),
.Y(n_1828)
);

NAND2xp5_ASAP7_75t_L g1829 ( 
.A(n_1825),
.B(n_1819),
.Y(n_1829)
);

NAND2xp5_ASAP7_75t_L g1830 ( 
.A(n_1822),
.B(n_1815),
.Y(n_1830)
);

NAND2xp5_ASAP7_75t_L g1831 ( 
.A(n_1824),
.B(n_1823),
.Y(n_1831)
);

AND2x2_ASAP7_75t_L g1832 ( 
.A(n_1821),
.B(n_1812),
.Y(n_1832)
);

AND2x2_ASAP7_75t_L g1833 ( 
.A(n_1823),
.B(n_1811),
.Y(n_1833)
);

INVx2_ASAP7_75t_SL g1834 ( 
.A(n_1823),
.Y(n_1834)
);

NAND2xp5_ASAP7_75t_L g1835 ( 
.A(n_1832),
.B(n_1817),
.Y(n_1835)
);

NAND2xp33_ASAP7_75t_SL g1836 ( 
.A(n_1826),
.B(n_1633),
.Y(n_1836)
);

INVxp67_ASAP7_75t_L g1837 ( 
.A(n_1833),
.Y(n_1837)
);

NAND2xp33_ASAP7_75t_SL g1838 ( 
.A(n_1828),
.B(n_1754),
.Y(n_1838)
);

NAND2xp5_ASAP7_75t_L g1839 ( 
.A(n_1827),
.B(n_1811),
.Y(n_1839)
);

INVxp67_ASAP7_75t_L g1840 ( 
.A(n_1834),
.Y(n_1840)
);

NOR2x1_ASAP7_75t_L g1841 ( 
.A(n_1831),
.B(n_1811),
.Y(n_1841)
);

CKINVDCx5p33_ASAP7_75t_R g1842 ( 
.A(n_1831),
.Y(n_1842)
);

AO221x2_ASAP7_75t_L g1843 ( 
.A1(n_1830),
.A2(n_1725),
.B1(n_1629),
.B2(n_1762),
.C(n_1759),
.Y(n_1843)
);

OR2x2_ASAP7_75t_L g1844 ( 
.A(n_1829),
.B(n_1816),
.Y(n_1844)
);

NAND2xp5_ASAP7_75t_L g1845 ( 
.A(n_1830),
.B(n_1777),
.Y(n_1845)
);

INVx1_ASAP7_75t_L g1846 ( 
.A(n_1845),
.Y(n_1846)
);

INVx1_ASAP7_75t_L g1847 ( 
.A(n_1835),
.Y(n_1847)
);

HB1xp67_ASAP7_75t_L g1848 ( 
.A(n_1840),
.Y(n_1848)
);

INVx1_ASAP7_75t_L g1849 ( 
.A(n_1841),
.Y(n_1849)
);

INVx1_ASAP7_75t_L g1850 ( 
.A(n_1839),
.Y(n_1850)
);

NAND2x1p5_ASAP7_75t_L g1851 ( 
.A(n_1844),
.B(n_1747),
.Y(n_1851)
);

OR2x2_ASAP7_75t_L g1852 ( 
.A(n_1837),
.B(n_1842),
.Y(n_1852)
);

INVx1_ASAP7_75t_L g1853 ( 
.A(n_1843),
.Y(n_1853)
);

OAI32xp33_ASAP7_75t_L g1854 ( 
.A1(n_1853),
.A2(n_1838),
.A3(n_1836),
.B1(n_1843),
.B2(n_1762),
.Y(n_1854)
);

AOI221x1_ASAP7_75t_L g1855 ( 
.A1(n_1849),
.A2(n_1758),
.B1(n_1523),
.B2(n_1632),
.C(n_1798),
.Y(n_1855)
);

INVx1_ASAP7_75t_L g1856 ( 
.A(n_1848),
.Y(n_1856)
);

OAI221xp5_ASAP7_75t_L g1857 ( 
.A1(n_1852),
.A2(n_1772),
.B1(n_1784),
.B2(n_1737),
.C(n_1747),
.Y(n_1857)
);

INVx1_ASAP7_75t_L g1858 ( 
.A(n_1856),
.Y(n_1858)
);

INVx2_ASAP7_75t_L g1859 ( 
.A(n_1857),
.Y(n_1859)
);

INVx1_ASAP7_75t_L g1860 ( 
.A(n_1854),
.Y(n_1860)
);

INVxp67_ASAP7_75t_L g1861 ( 
.A(n_1855),
.Y(n_1861)
);

NAND2xp5_ASAP7_75t_L g1862 ( 
.A(n_1860),
.B(n_1847),
.Y(n_1862)
);

OAI21xp33_ASAP7_75t_L g1863 ( 
.A1(n_1859),
.A2(n_1851),
.B(n_1850),
.Y(n_1863)
);

NAND2xp5_ASAP7_75t_L g1864 ( 
.A(n_1861),
.B(n_1858),
.Y(n_1864)
);

AOI21xp33_ASAP7_75t_L g1865 ( 
.A1(n_1861),
.A2(n_1851),
.B(n_1846),
.Y(n_1865)
);

AOI21xp5_ASAP7_75t_L g1866 ( 
.A1(n_1861),
.A2(n_1731),
.B(n_1643),
.Y(n_1866)
);

INVx2_ASAP7_75t_L g1867 ( 
.A(n_1864),
.Y(n_1867)
);

INVx1_ASAP7_75t_L g1868 ( 
.A(n_1862),
.Y(n_1868)
);

AND2x2_ASAP7_75t_L g1869 ( 
.A(n_1866),
.B(n_1628),
.Y(n_1869)
);

HB1xp67_ASAP7_75t_L g1870 ( 
.A(n_1865),
.Y(n_1870)
);

INVx1_ASAP7_75t_L g1871 ( 
.A(n_1863),
.Y(n_1871)
);

INVx1_ASAP7_75t_L g1872 ( 
.A(n_1864),
.Y(n_1872)
);

INVx1_ASAP7_75t_L g1873 ( 
.A(n_1864),
.Y(n_1873)
);

INVx2_ASAP7_75t_L g1874 ( 
.A(n_1864),
.Y(n_1874)
);

NAND2xp5_ASAP7_75t_L g1875 ( 
.A(n_1866),
.B(n_1802),
.Y(n_1875)
);

INVx1_ASAP7_75t_L g1876 ( 
.A(n_1864),
.Y(n_1876)
);

NAND2xp5_ASAP7_75t_L g1877 ( 
.A(n_1870),
.B(n_1677),
.Y(n_1877)
);

NOR2x1_ASAP7_75t_L g1878 ( 
.A(n_1867),
.B(n_1874),
.Y(n_1878)
);

NAND3xp33_ASAP7_75t_SL g1879 ( 
.A(n_1872),
.B(n_1641),
.C(n_1699),
.Y(n_1879)
);

AOI211xp5_ASAP7_75t_L g1880 ( 
.A1(n_1871),
.A2(n_1630),
.B(n_1644),
.C(n_1703),
.Y(n_1880)
);

AND3x1_ASAP7_75t_L g1881 ( 
.A(n_1869),
.B(n_1657),
.C(n_1593),
.Y(n_1881)
);

NAND3xp33_ASAP7_75t_L g1882 ( 
.A(n_1873),
.B(n_1686),
.C(n_1576),
.Y(n_1882)
);

NOR2x1_ASAP7_75t_L g1883 ( 
.A(n_1876),
.B(n_1567),
.Y(n_1883)
);

AOI211x1_ASAP7_75t_L g1884 ( 
.A1(n_1875),
.A2(n_1738),
.B(n_1589),
.C(n_1596),
.Y(n_1884)
);

INVx2_ASAP7_75t_L g1885 ( 
.A(n_1875),
.Y(n_1885)
);

OAI322xp33_ASAP7_75t_L g1886 ( 
.A1(n_1868),
.A2(n_1554),
.A3(n_1799),
.B1(n_1798),
.B2(n_1537),
.C1(n_1562),
.C2(n_1658),
.Y(n_1886)
);

NAND2xp5_ASAP7_75t_L g1887 ( 
.A(n_1870),
.B(n_1801),
.Y(n_1887)
);

NOR3xp33_ASAP7_75t_L g1888 ( 
.A(n_1870),
.B(n_1700),
.C(n_1667),
.Y(n_1888)
);

NAND4xp25_ASAP7_75t_L g1889 ( 
.A(n_1888),
.B(n_1784),
.C(n_1772),
.D(n_1646),
.Y(n_1889)
);

OAI221xp5_ASAP7_75t_L g1890 ( 
.A1(n_1880),
.A2(n_1737),
.B1(n_1756),
.B2(n_1735),
.C(n_1760),
.Y(n_1890)
);

AOI211x1_ASAP7_75t_SL g1891 ( 
.A1(n_1887),
.A2(n_1799),
.B(n_1798),
.C(n_1670),
.Y(n_1891)
);

NAND2xp5_ASAP7_75t_L g1892 ( 
.A(n_1885),
.B(n_1713),
.Y(n_1892)
);

NOR3x1_ASAP7_75t_L g1893 ( 
.A(n_1877),
.B(n_1670),
.C(n_1755),
.Y(n_1893)
);

OAI211xp5_ASAP7_75t_SL g1894 ( 
.A1(n_1878),
.A2(n_1706),
.B(n_1627),
.C(n_1581),
.Y(n_1894)
);

AOI211xp5_ASAP7_75t_L g1895 ( 
.A1(n_1879),
.A2(n_1737),
.B(n_1798),
.C(n_1799),
.Y(n_1895)
);

AOI211xp5_ASAP7_75t_L g1896 ( 
.A1(n_1886),
.A2(n_1737),
.B(n_1799),
.C(n_1748),
.Y(n_1896)
);

NOR3xp33_ASAP7_75t_SL g1897 ( 
.A(n_1882),
.B(n_1547),
.C(n_1578),
.Y(n_1897)
);

NAND2xp5_ASAP7_75t_L g1898 ( 
.A(n_1884),
.B(n_1713),
.Y(n_1898)
);

NOR2xp67_ASAP7_75t_L g1899 ( 
.A(n_1881),
.B(n_1653),
.Y(n_1899)
);

NOR3xp33_ASAP7_75t_L g1900 ( 
.A(n_1883),
.B(n_1764),
.C(n_1760),
.Y(n_1900)
);

AOI211xp5_ASAP7_75t_SL g1901 ( 
.A1(n_1899),
.A2(n_1642),
.B(n_1664),
.C(n_1746),
.Y(n_1901)
);

AOI211xp5_ASAP7_75t_L g1902 ( 
.A1(n_1892),
.A2(n_1894),
.B(n_1895),
.C(n_1896),
.Y(n_1902)
);

NAND4xp25_ASAP7_75t_SL g1903 ( 
.A(n_1898),
.B(n_1674),
.C(n_1764),
.D(n_1634),
.Y(n_1903)
);

NAND2xp5_ASAP7_75t_L g1904 ( 
.A(n_1891),
.B(n_1799),
.Y(n_1904)
);

OAI211xp5_ASAP7_75t_L g1905 ( 
.A1(n_1900),
.A2(n_1698),
.B(n_1694),
.C(n_1663),
.Y(n_1905)
);

OAI211xp5_ASAP7_75t_L g1906 ( 
.A1(n_1897),
.A2(n_1698),
.B(n_1694),
.C(n_1661),
.Y(n_1906)
);

AOI221xp5_ASAP7_75t_L g1907 ( 
.A1(n_1889),
.A2(n_1890),
.B1(n_1893),
.B2(n_1793),
.C(n_1648),
.Y(n_1907)
);

INVx1_ASAP7_75t_L g1908 ( 
.A(n_1892),
.Y(n_1908)
);

NAND3xp33_ASAP7_75t_SL g1909 ( 
.A(n_1895),
.B(n_1651),
.C(n_1717),
.Y(n_1909)
);

O2A1O1Ixp5_ASAP7_75t_SL g1910 ( 
.A1(n_1892),
.A2(n_1642),
.B(n_1664),
.C(n_1768),
.Y(n_1910)
);

NOR3xp33_ASAP7_75t_L g1911 ( 
.A(n_1892),
.B(n_1565),
.C(n_1755),
.Y(n_1911)
);

AOI22xp5_ASAP7_75t_L g1912 ( 
.A1(n_1903),
.A2(n_1909),
.B1(n_1907),
.B2(n_1908),
.Y(n_1912)
);

NOR3xp33_ASAP7_75t_SL g1913 ( 
.A(n_1906),
.B(n_1612),
.C(n_1717),
.Y(n_1913)
);

NOR3xp33_ASAP7_75t_L g1914 ( 
.A(n_1902),
.B(n_1905),
.C(n_1904),
.Y(n_1914)
);

OA21x2_ASAP7_75t_L g1915 ( 
.A1(n_1901),
.A2(n_1793),
.B(n_1757),
.Y(n_1915)
);

AOI21xp5_ASAP7_75t_L g1916 ( 
.A1(n_1911),
.A2(n_1683),
.B(n_1753),
.Y(n_1916)
);

NAND2xp5_ASAP7_75t_L g1917 ( 
.A(n_1910),
.B(n_1806),
.Y(n_1917)
);

NAND4xp75_ASAP7_75t_L g1918 ( 
.A(n_1908),
.B(n_1800),
.C(n_1753),
.D(n_1763),
.Y(n_1918)
);

NAND4xp75_ASAP7_75t_L g1919 ( 
.A(n_1908),
.B(n_1800),
.C(n_1757),
.D(n_1763),
.Y(n_1919)
);

NAND2xp5_ASAP7_75t_L g1920 ( 
.A(n_1901),
.B(n_1806),
.Y(n_1920)
);

INVx1_ASAP7_75t_L g1921 ( 
.A(n_1904),
.Y(n_1921)
);

AOI211xp5_ASAP7_75t_L g1922 ( 
.A1(n_1909),
.A2(n_1748),
.B(n_1697),
.C(n_1656),
.Y(n_1922)
);

AND3x4_ASAP7_75t_L g1923 ( 
.A(n_1911),
.B(n_1773),
.C(n_1684),
.Y(n_1923)
);

OAI211xp5_ASAP7_75t_SL g1924 ( 
.A1(n_1902),
.A2(n_1746),
.B(n_1638),
.C(n_1631),
.Y(n_1924)
);

INVxp67_ASAP7_75t_L g1925 ( 
.A(n_1904),
.Y(n_1925)
);

HB1xp67_ASAP7_75t_L g1926 ( 
.A(n_1925),
.Y(n_1926)
);

NAND4xp75_ASAP7_75t_L g1927 ( 
.A(n_1921),
.B(n_1809),
.C(n_1761),
.D(n_1692),
.Y(n_1927)
);

NAND2xp5_ASAP7_75t_L g1928 ( 
.A(n_1914),
.B(n_1806),
.Y(n_1928)
);

NOR3xp33_ASAP7_75t_SL g1929 ( 
.A(n_1918),
.B(n_1559),
.C(n_1739),
.Y(n_1929)
);

NAND3xp33_ASAP7_75t_SL g1930 ( 
.A(n_1912),
.B(n_1787),
.C(n_1556),
.Y(n_1930)
);

NOR2x1_ASAP7_75t_L g1931 ( 
.A(n_1923),
.B(n_1697),
.Y(n_1931)
);

NAND2xp5_ASAP7_75t_L g1932 ( 
.A(n_1919),
.B(n_1806),
.Y(n_1932)
);

INVx1_ASAP7_75t_L g1933 ( 
.A(n_1917),
.Y(n_1933)
);

AND2x4_ASAP7_75t_L g1934 ( 
.A(n_1913),
.B(n_1773),
.Y(n_1934)
);

AND2x4_ASAP7_75t_L g1935 ( 
.A(n_1916),
.B(n_1773),
.Y(n_1935)
);

NAND2xp5_ASAP7_75t_L g1936 ( 
.A(n_1922),
.B(n_1806),
.Y(n_1936)
);

AND2x2_ASAP7_75t_SL g1937 ( 
.A(n_1915),
.B(n_1748),
.Y(n_1937)
);

INVx2_ASAP7_75t_L g1938 ( 
.A(n_1915),
.Y(n_1938)
);

NOR2xp67_ASAP7_75t_L g1939 ( 
.A(n_1920),
.B(n_1698),
.Y(n_1939)
);

OAI22xp5_ASAP7_75t_L g1940 ( 
.A1(n_1928),
.A2(n_1926),
.B1(n_1931),
.B2(n_1927),
.Y(n_1940)
);

INVx2_ASAP7_75t_L g1941 ( 
.A(n_1937),
.Y(n_1941)
);

INVx4_ASAP7_75t_L g1942 ( 
.A(n_1938),
.Y(n_1942)
);

INVx2_ASAP7_75t_L g1943 ( 
.A(n_1934),
.Y(n_1943)
);

NAND3xp33_ASAP7_75t_SL g1944 ( 
.A(n_1933),
.B(n_1924),
.C(n_1787),
.Y(n_1944)
);

AND2x2_ASAP7_75t_L g1945 ( 
.A(n_1935),
.B(n_1804),
.Y(n_1945)
);

AOI22xp5_ASAP7_75t_L g1946 ( 
.A1(n_1930),
.A2(n_1795),
.B1(n_1697),
.B2(n_1681),
.Y(n_1946)
);

NAND2xp5_ASAP7_75t_L g1947 ( 
.A(n_1939),
.B(n_1779),
.Y(n_1947)
);

OAI22xp5_ASAP7_75t_L g1948 ( 
.A1(n_1932),
.A2(n_1936),
.B1(n_1929),
.B2(n_1675),
.Y(n_1948)
);

NAND2xp5_ASAP7_75t_L g1949 ( 
.A(n_1934),
.B(n_1779),
.Y(n_1949)
);

AO22x2_ASAP7_75t_L g1950 ( 
.A1(n_1941),
.A2(n_1940),
.B1(n_1942),
.B2(n_1943),
.Y(n_1950)
);

INVx1_ASAP7_75t_L g1951 ( 
.A(n_1949),
.Y(n_1951)
);

OAI22xp5_ASAP7_75t_SL g1952 ( 
.A1(n_1948),
.A2(n_1681),
.B1(n_1675),
.B2(n_1672),
.Y(n_1952)
);

AO22x1_ASAP7_75t_L g1953 ( 
.A1(n_1945),
.A2(n_1682),
.B1(n_1656),
.B2(n_1746),
.Y(n_1953)
);

INVx1_ASAP7_75t_L g1954 ( 
.A(n_1947),
.Y(n_1954)
);

AOI22xp5_ASAP7_75t_L g1955 ( 
.A1(n_1944),
.A2(n_1672),
.B1(n_1682),
.B2(n_1656),
.Y(n_1955)
);

INVx1_ASAP7_75t_L g1956 ( 
.A(n_1946),
.Y(n_1956)
);

HB1xp67_ASAP7_75t_L g1957 ( 
.A(n_1941),
.Y(n_1957)
);

AOI22xp33_ASAP7_75t_L g1958 ( 
.A1(n_1943),
.A2(n_1682),
.B1(n_1774),
.B2(n_1769),
.Y(n_1958)
);

OAI22xp5_ASAP7_75t_SL g1959 ( 
.A1(n_1957),
.A2(n_1702),
.B1(n_1520),
.B2(n_1774),
.Y(n_1959)
);

INVx1_ASAP7_75t_L g1960 ( 
.A(n_1950),
.Y(n_1960)
);

INVxp33_ASAP7_75t_SL g1961 ( 
.A(n_1956),
.Y(n_1961)
);

INVx1_ASAP7_75t_L g1962 ( 
.A(n_1952),
.Y(n_1962)
);

OAI22x1_ASAP7_75t_L g1963 ( 
.A1(n_1954),
.A2(n_1769),
.B1(n_1791),
.B2(n_1794),
.Y(n_1963)
);

INVx1_ASAP7_75t_L g1964 ( 
.A(n_1951),
.Y(n_1964)
);

NAND2xp5_ASAP7_75t_L g1965 ( 
.A(n_1955),
.B(n_1513),
.Y(n_1965)
);

OAI21xp5_ASAP7_75t_L g1966 ( 
.A1(n_1958),
.A2(n_1584),
.B(n_1780),
.Y(n_1966)
);

OAI21xp5_ASAP7_75t_L g1967 ( 
.A1(n_1960),
.A2(n_1953),
.B(n_1780),
.Y(n_1967)
);

INVx1_ASAP7_75t_L g1968 ( 
.A(n_1964),
.Y(n_1968)
);

AO22x1_ASAP7_75t_L g1969 ( 
.A1(n_1961),
.A2(n_1809),
.B1(n_1520),
.B2(n_1769),
.Y(n_1969)
);

OA21x2_ASAP7_75t_L g1970 ( 
.A1(n_1962),
.A2(n_1780),
.B(n_1796),
.Y(n_1970)
);

OAI21xp5_ASAP7_75t_L g1971 ( 
.A1(n_1965),
.A2(n_1570),
.B(n_1569),
.Y(n_1971)
);

AOI22xp5_ASAP7_75t_L g1972 ( 
.A1(n_1959),
.A2(n_1702),
.B1(n_1804),
.B2(n_1769),
.Y(n_1972)
);

NAND2xp5_ASAP7_75t_SL g1973 ( 
.A(n_1963),
.B(n_1794),
.Y(n_1973)
);

CKINVDCx20_ASAP7_75t_R g1974 ( 
.A(n_1968),
.Y(n_1974)
);

INVx1_ASAP7_75t_SL g1975 ( 
.A(n_1967),
.Y(n_1975)
);

INVx1_ASAP7_75t_L g1976 ( 
.A(n_1972),
.Y(n_1976)
);

INVx1_ASAP7_75t_L g1977 ( 
.A(n_1973),
.Y(n_1977)
);

HB1xp67_ASAP7_75t_L g1978 ( 
.A(n_1970),
.Y(n_1978)
);

NAND4xp25_ASAP7_75t_SL g1979 ( 
.A(n_1969),
.B(n_1966),
.C(n_1796),
.D(n_1803),
.Y(n_1979)
);

AOI22xp5_ASAP7_75t_L g1980 ( 
.A1(n_1974),
.A2(n_1971),
.B1(n_1769),
.B2(n_1785),
.Y(n_1980)
);

INVx1_ASAP7_75t_L g1981 ( 
.A(n_1978),
.Y(n_1981)
);

AOI221xp5_ASAP7_75t_L g1982 ( 
.A1(n_1975),
.A2(n_1803),
.B1(n_1805),
.B2(n_1786),
.C(n_1788),
.Y(n_1982)
);

OAI22xp5_ASAP7_75t_L g1983 ( 
.A1(n_1981),
.A2(n_1976),
.B1(n_1977),
.B2(n_1979),
.Y(n_1983)
);

OAI22xp33_ASAP7_75t_L g1984 ( 
.A1(n_1980),
.A2(n_1791),
.B1(n_1807),
.B2(n_1805),
.Y(n_1984)
);

OAI21x1_ASAP7_75t_L g1985 ( 
.A1(n_1983),
.A2(n_1982),
.B(n_1536),
.Y(n_1985)
);

OAI21xp33_ASAP7_75t_L g1986 ( 
.A1(n_1985),
.A2(n_1984),
.B(n_1788),
.Y(n_1986)
);

AOI22xp5_ASAP7_75t_L g1987 ( 
.A1(n_1986),
.A2(n_1783),
.B1(n_1560),
.B2(n_1781),
.Y(n_1987)
);

AOI211xp5_ASAP7_75t_L g1988 ( 
.A1(n_1987),
.A2(n_1543),
.B(n_1534),
.C(n_1555),
.Y(n_1988)
);


endmodule