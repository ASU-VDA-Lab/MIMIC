module real_jpeg_14744_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

BUFx16f_ASAP7_75t_L g46 ( 
.A(n_1),
.Y(n_46)
);

BUFx12_ASAP7_75t_L g62 ( 
.A(n_2),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_3),
.A2(n_60),
.B1(n_61),
.B2(n_66),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_3),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_3),
.A2(n_55),
.B1(n_58),
.B2(n_66),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_3),
.A2(n_42),
.B1(n_43),
.B2(n_66),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_3),
.A2(n_30),
.B1(n_37),
.B2(n_66),
.Y(n_213)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_4),
.A2(n_55),
.B1(n_58),
.B2(n_74),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_4),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_4),
.A2(n_60),
.B1(n_61),
.B2(n_74),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_L g115 ( 
.A1(n_4),
.A2(n_42),
.B1(n_43),
.B2(n_74),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_4),
.A2(n_30),
.B1(n_37),
.B2(n_74),
.Y(n_171)
);

BUFx16f_ASAP7_75t_L g42 ( 
.A(n_5),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_6),
.A2(n_42),
.B1(n_43),
.B2(n_50),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_6),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_L g93 ( 
.A1(n_6),
.A2(n_50),
.B1(n_55),
.B2(n_58),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_L g111 ( 
.A1(n_6),
.A2(n_30),
.B1(n_37),
.B2(n_50),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g317 ( 
.A1(n_6),
.A2(n_50),
.B1(n_60),
.B2(n_61),
.Y(n_317)
);

AOI22xp33_ASAP7_75t_SL g155 ( 
.A1(n_7),
.A2(n_60),
.B1(n_61),
.B2(n_156),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_7),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_SL g199 ( 
.A1(n_7),
.A2(n_55),
.B1(n_58),
.B2(n_156),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g256 ( 
.A1(n_7),
.A2(n_42),
.B1(n_43),
.B2(n_156),
.Y(n_256)
);

OAI22xp33_ASAP7_75t_SL g263 ( 
.A1(n_7),
.A2(n_30),
.B1(n_37),
.B2(n_156),
.Y(n_263)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_8),
.Y(n_55)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_9),
.Y(n_175)
);

AOI21xp33_ASAP7_75t_L g195 ( 
.A1(n_9),
.A2(n_60),
.B(n_196),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_9),
.B(n_186),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_9),
.B(n_58),
.Y(n_234)
);

OAI22xp33_ASAP7_75t_L g248 ( 
.A1(n_9),
.A2(n_42),
.B1(n_43),
.B2(n_175),
.Y(n_248)
);

O2A1O1Ixp33_ASAP7_75t_L g250 ( 
.A1(n_9),
.A2(n_43),
.B(n_46),
.C(n_251),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_9),
.B(n_82),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_9),
.B(n_34),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_9),
.B(n_51),
.Y(n_275)
);

AOI21xp33_ASAP7_75t_L g284 ( 
.A1(n_9),
.A2(n_58),
.B(n_234),
.Y(n_284)
);

AOI22xp33_ASAP7_75t_L g182 ( 
.A1(n_10),
.A2(n_60),
.B1(n_61),
.B2(n_183),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_10),
.Y(n_183)
);

AOI22xp33_ASAP7_75t_SL g209 ( 
.A1(n_10),
.A2(n_55),
.B1(n_58),
.B2(n_183),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_L g249 ( 
.A1(n_10),
.A2(n_42),
.B1(n_43),
.B2(n_183),
.Y(n_249)
);

OAI22xp33_ASAP7_75t_SL g270 ( 
.A1(n_10),
.A2(n_30),
.B1(n_37),
.B2(n_183),
.Y(n_270)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_11),
.A2(n_60),
.B1(n_61),
.B2(n_64),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_11),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_11),
.A2(n_55),
.B1(n_58),
.B2(n_64),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_11),
.A2(n_42),
.B1(n_43),
.B2(n_64),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_11),
.A2(n_30),
.B1(n_37),
.B2(n_64),
.Y(n_237)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_12),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_13),
.A2(n_60),
.B1(n_61),
.B2(n_120),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_13),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g178 ( 
.A1(n_13),
.A2(n_55),
.B1(n_58),
.B2(n_120),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_SL g228 ( 
.A1(n_13),
.A2(n_42),
.B1(n_43),
.B2(n_120),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_13),
.A2(n_30),
.B1(n_37),
.B2(n_120),
.Y(n_258)
);

BUFx8_ASAP7_75t_L g57 ( 
.A(n_14),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g35 ( 
.A1(n_15),
.A2(n_30),
.B1(n_36),
.B2(n_37),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_15),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_15),
.A2(n_36),
.B1(n_42),
.B2(n_43),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_15),
.A2(n_36),
.B1(n_55),
.B2(n_58),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g326 ( 
.A1(n_15),
.A2(n_36),
.B1(n_60),
.B2(n_61),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_L g40 ( 
.A1(n_16),
.A2(n_41),
.B1(n_42),
.B2(n_43),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_16),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_16),
.A2(n_41),
.B1(n_55),
.B2(n_58),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_16),
.A2(n_41),
.B1(n_60),
.B2(n_61),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_16),
.A2(n_30),
.B1(n_37),
.B2(n_41),
.Y(n_147)
);

INVx11_ASAP7_75t_L g32 ( 
.A(n_17),
.Y(n_32)
);

XOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_322),
.Y(n_18)
);

AOI21xp5_ASAP7_75t_SL g19 ( 
.A1(n_20),
.A2(n_309),
.B(n_321),
.Y(n_19)
);

AO21x1_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_134),
.B(n_306),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_121),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_SL g22 ( 
.A(n_23),
.B(n_97),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_23),
.B(n_97),
.Y(n_307)
);

XOR2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_67),
.Y(n_23)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_24),
.B(n_83),
.C(n_95),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_28),
.B(n_52),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_25),
.A2(n_26),
.B1(n_100),
.B2(n_101),
.Y(n_99)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_38),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_27),
.A2(n_28),
.B1(n_52),
.B2(n_102),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_27),
.A2(n_28),
.B1(n_38),
.B2(n_39),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_28),
.Y(n_27)
);

OAI21xp5_ASAP7_75t_SL g28 ( 
.A1(n_29),
.A2(n_34),
.B(n_35),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_29),
.A2(n_34),
.B1(n_35),
.B2(n_110),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_29),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_29),
.A2(n_34),
.B1(n_147),
.B2(n_171),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_29),
.A2(n_34),
.B1(n_171),
.B2(n_213),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_29),
.A2(n_34),
.B1(n_213),
.B2(n_237),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_29),
.A2(n_34),
.B1(n_237),
.B2(n_258),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_29),
.A2(n_34),
.B1(n_175),
.B2(n_270),
.Y(n_269)
);

AOI22xp33_ASAP7_75t_L g274 ( 
.A1(n_29),
.A2(n_34),
.B1(n_263),
.B2(n_270),
.Y(n_274)
);

AND2x2_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_33),
.Y(n_29)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_30),
.Y(n_37)
);

OA22x2_ASAP7_75t_L g48 ( 
.A1(n_30),
.A2(n_37),
.B1(n_46),
.B2(n_47),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_30),
.B(n_272),
.Y(n_271)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_33),
.A2(n_111),
.B1(n_145),
.B2(n_146),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_33),
.A2(n_145),
.B1(n_262),
.B2(n_264),
.Y(n_261)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

OAI21xp33_ASAP7_75t_L g251 ( 
.A1(n_37),
.A2(n_47),
.B(n_175),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_39),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g39 ( 
.A1(n_40),
.A2(n_44),
.B1(n_49),
.B2(n_51),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_40),
.A2(n_44),
.B1(n_51),
.B2(n_114),
.Y(n_113)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_42),
.Y(n_43)
);

OAI22xp33_ASAP7_75t_L g45 ( 
.A1(n_42),
.A2(n_43),
.B1(n_46),
.B2(n_47),
.Y(n_45)
);

OA22x2_ASAP7_75t_L g77 ( 
.A1(n_42),
.A2(n_43),
.B1(n_78),
.B2(n_79),
.Y(n_77)
);

OAI32xp33_ASAP7_75t_L g232 ( 
.A1(n_42),
.A2(n_58),
.A3(n_79),
.B1(n_233),
.B2(n_235),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_43),
.B(n_78),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_44),
.A2(n_49),
.B1(n_51),
.B2(n_70),
.Y(n_69)
);

OAI21xp5_ASAP7_75t_L g89 ( 
.A1(n_44),
.A2(n_51),
.B(n_70),
.Y(n_89)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_44),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_44),
.A2(n_51),
.B1(n_150),
.B2(n_201),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_44),
.A2(n_51),
.B1(n_201),
.B2(n_227),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_44),
.A2(n_51),
.B1(n_248),
.B2(n_249),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_44),
.A2(n_51),
.B1(n_249),
.B2(n_256),
.Y(n_255)
);

AND2x2_ASAP7_75t_L g44 ( 
.A(n_45),
.B(n_48),
.Y(n_44)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_46),
.Y(n_47)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_48),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_48),
.A2(n_115),
.B1(n_149),
.B2(n_151),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_48),
.A2(n_151),
.B1(n_228),
.B2(n_286),
.Y(n_285)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_52),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_53),
.A2(n_54),
.B1(n_63),
.B2(n_65),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_53),
.A2(n_54),
.B1(n_65),
.B2(n_86),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_53),
.A2(n_54),
.B1(n_63),
.B2(n_119),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_53),
.A2(n_54),
.B1(n_86),
.B2(n_133),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_53),
.A2(n_54),
.B1(n_119),
.B2(n_155),
.Y(n_154)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_53),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_53),
.A2(n_54),
.B1(n_182),
.B2(n_195),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_54),
.B(n_59),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_54),
.Y(n_186)
);

OA22x2_ASAP7_75t_L g54 ( 
.A1(n_55),
.A2(n_56),
.B1(n_57),
.B2(n_58),
.Y(n_54)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_55),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_55),
.A2(n_58),
.B1(n_78),
.B2(n_79),
.Y(n_80)
);

OAI32xp33_ASAP7_75t_L g172 ( 
.A1(n_55),
.A2(n_57),
.A3(n_60),
.B1(n_173),
.B2(n_174),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_56),
.A2(n_57),
.B1(n_60),
.B2(n_61),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_56),
.B(n_58),
.Y(n_173)
);

INVx11_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_61),
.B(n_175),
.Y(n_174)
);

BUFx16f_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_68),
.A2(n_83),
.B1(n_95),
.B2(n_96),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_68),
.Y(n_95)
);

OAI21xp33_ASAP7_75t_L g104 ( 
.A1(n_68),
.A2(n_69),
.B(n_71),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_69),
.B(n_71),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_72),
.A2(n_75),
.B1(n_81),
.B2(n_82),
.Y(n_71)
);

INVxp67_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_73),
.A2(n_76),
.B1(n_77),
.B2(n_117),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_75),
.A2(n_81),
.B1(n_82),
.B2(n_92),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_75),
.A2(n_82),
.B1(n_177),
.B2(n_179),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_75),
.A2(n_82),
.B1(n_208),
.B2(n_210),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_SL g313 ( 
.A1(n_75),
.A2(n_82),
.B(n_314),
.Y(n_313)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_76),
.A2(n_77),
.B1(n_93),
.B2(n_131),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_76),
.A2(n_77),
.B1(n_117),
.B2(n_153),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_76),
.A2(n_77),
.B1(n_178),
.B2(n_199),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_76),
.A2(n_77),
.B1(n_209),
.B2(n_284),
.Y(n_283)
);

NAND2x1_ASAP7_75t_SL g76 ( 
.A(n_77),
.B(n_80),
.Y(n_76)
);

INVx1_ASAP7_75t_SL g82 ( 
.A(n_77),
.Y(n_82)
);

INVx8_ASAP7_75t_L g79 ( 
.A(n_78),
.Y(n_79)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_83),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_84),
.A2(n_85),
.B1(n_87),
.B2(n_88),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_84),
.A2(n_85),
.B1(n_126),
.B2(n_127),
.Y(n_125)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_85),
.B(n_89),
.C(n_91),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_85),
.B(n_124),
.C(n_127),
.Y(n_310)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_89),
.A2(n_90),
.B1(n_91),
.B2(n_94),
.Y(n_88)
);

CKINVDCx14_ASAP7_75t_R g94 ( 
.A(n_89),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_89),
.A2(n_94),
.B1(n_129),
.B2(n_130),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_89),
.B(n_130),
.C(n_132),
.Y(n_320)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

CKINVDCx14_ASAP7_75t_R g92 ( 
.A(n_93),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_103),
.C(n_105),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_98),
.A2(n_99),
.B1(n_103),
.B2(n_104),
.Y(n_158)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

XOR2xp5_ASAP7_75t_L g157 ( 
.A(n_105),
.B(n_158),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_106),
.B(n_116),
.C(n_118),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_106),
.A2(n_107),
.B1(n_138),
.B2(n_139),
.Y(n_137)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_112),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_108),
.A2(n_109),
.B1(n_112),
.B2(n_113),
.Y(n_166)
);

CKINVDCx14_ASAP7_75t_R g108 ( 
.A(n_109),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

CKINVDCx14_ASAP7_75t_R g112 ( 
.A(n_113),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

XOR2xp5_ASAP7_75t_L g139 ( 
.A(n_116),
.B(n_118),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_L g306 ( 
.A1(n_121),
.A2(n_307),
.B(n_308),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_123),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_122),
.B(n_123),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_125),
.Y(n_123)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_132),
.Y(n_127)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

CKINVDCx16_ASAP7_75t_R g314 ( 
.A(n_131),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_133),
.Y(n_316)
);

OAI21xp5_ASAP7_75t_L g134 ( 
.A1(n_135),
.A2(n_159),
.B(n_305),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_157),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_136),
.B(n_157),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_140),
.C(n_141),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_137),
.B(n_140),
.Y(n_188)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_141),
.B(n_188),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_152),
.C(n_154),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_142),
.A2(n_143),
.B1(n_164),
.B2(n_165),
.Y(n_163)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_148),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_144),
.B(n_148),
.Y(n_217)
);

CKINVDCx14_ASAP7_75t_R g146 ( 
.A(n_147),
.Y(n_146)
);

CKINVDCx16_ASAP7_75t_R g149 ( 
.A(n_150),
.Y(n_149)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_152),
.B(n_154),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g179 ( 
.A(n_153),
.Y(n_179)
);

INVxp67_ASAP7_75t_L g185 ( 
.A(n_155),
.Y(n_185)
);

AOI21xp5_ASAP7_75t_SL g159 ( 
.A1(n_160),
.A2(n_189),
.B(n_304),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_187),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_161),
.B(n_187),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_166),
.C(n_167),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_162),
.A2(n_163),
.B1(n_166),
.B2(n_302),
.Y(n_301)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_166),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_167),
.B(n_301),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_176),
.C(n_180),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_168),
.B(n_219),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_169),
.B(n_172),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_169),
.A2(n_170),
.B1(n_172),
.B2(n_205),
.Y(n_204)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_172),
.Y(n_205)
);

CKINVDCx16_ASAP7_75t_R g196 ( 
.A(n_174),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_176),
.B(n_180),
.Y(n_219)
);

INVxp67_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_181),
.A2(n_184),
.B1(n_185),
.B2(n_186),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_184),
.A2(n_186),
.B1(n_316),
.B2(n_317),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_SL g325 ( 
.A1(n_184),
.A2(n_186),
.B1(n_317),
.B2(n_326),
.Y(n_325)
);

A2O1A1Ixp33_ASAP7_75t_SL g189 ( 
.A1(n_190),
.A2(n_220),
.B(n_298),
.C(n_303),
.Y(n_189)
);

OR2x2_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_214),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_191),
.B(n_214),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_204),
.C(n_206),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_192),
.A2(n_193),
.B1(n_239),
.B2(n_240),
.Y(n_238)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_197),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_194),
.B(n_198),
.C(n_203),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_198),
.A2(n_200),
.B1(n_202),
.B2(n_203),
.Y(n_197)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_198),
.Y(n_202)
);

INVxp67_ASAP7_75t_L g210 ( 
.A(n_199),
.Y(n_210)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_200),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_SL g239 ( 
.A(n_204),
.B(n_206),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_211),
.C(n_212),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_SL g224 ( 
.A(n_207),
.B(n_225),
.Y(n_224)
);

INVxp67_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_211),
.B(n_212),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_218),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_217),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_216),
.B(n_217),
.C(n_218),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_221),
.B(n_297),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_L g221 ( 
.A1(n_222),
.A2(n_241),
.B(n_296),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_238),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g296 ( 
.A(n_223),
.B(n_238),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_226),
.C(n_229),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g292 ( 
.A(n_224),
.B(n_293),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_L g293 ( 
.A1(n_226),
.A2(n_229),
.B1(n_230),
.B2(n_294),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_226),
.Y(n_294)
);

INVxp67_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_236),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_231),
.A2(n_232),
.B1(n_236),
.B2(n_288),
.Y(n_287)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_236),
.Y(n_288)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_239),
.Y(n_240)
);

AOI21xp5_ASAP7_75t_L g241 ( 
.A1(n_242),
.A2(n_290),
.B(n_295),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_SL g242 ( 
.A1(n_243),
.A2(n_279),
.B(n_289),
.Y(n_242)
);

AOI21xp5_ASAP7_75t_L g243 ( 
.A1(n_244),
.A2(n_259),
.B(n_278),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_252),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_SL g278 ( 
.A(n_245),
.B(n_252),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_246),
.B(n_250),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_246),
.A2(n_247),
.B1(n_250),
.B2(n_266),
.Y(n_265)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_250),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_257),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_255),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_254),
.B(n_255),
.C(n_257),
.Y(n_280)
);

INVxp67_ASAP7_75t_L g286 ( 
.A(n_256),
.Y(n_286)
);

CKINVDCx14_ASAP7_75t_R g264 ( 
.A(n_258),
.Y(n_264)
);

OAI21xp5_ASAP7_75t_SL g259 ( 
.A1(n_260),
.A2(n_267),
.B(n_277),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_265),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_SL g277 ( 
.A(n_261),
.B(n_265),
.Y(n_277)
);

INVxp67_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

AOI21xp5_ASAP7_75t_L g267 ( 
.A1(n_268),
.A2(n_273),
.B(n_276),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_SL g268 ( 
.A(n_269),
.B(n_271),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_274),
.B(n_275),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_SL g276 ( 
.A(n_274),
.B(n_275),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_280),
.B(n_281),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_SL g289 ( 
.A(n_280),
.B(n_281),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_282),
.B(n_287),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_283),
.B(n_285),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_283),
.B(n_285),
.C(n_287),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_291),
.B(n_292),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_SL g295 ( 
.A(n_291),
.B(n_292),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_299),
.B(n_300),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_299),
.B(n_300),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_310),
.B(n_311),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_310),
.B(n_311),
.Y(n_321)
);

XNOR2xp5_ASAP7_75t_L g311 ( 
.A(n_312),
.B(n_320),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_313),
.A2(n_315),
.B1(n_318),
.B2(n_319),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_313),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_315),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_315),
.B(n_318),
.C(n_320),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_323),
.B(n_329),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_324),
.B(n_327),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_325),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_325),
.B(n_328),
.Y(n_329)
);

CKINVDCx14_ASAP7_75t_R g327 ( 
.A(n_328),
.Y(n_327)
);


endmodule