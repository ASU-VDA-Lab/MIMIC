module fake_jpeg_4116_n_202 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_202);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_202;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

BUFx12f_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_12),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_11),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

INVx11_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_9),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_5),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_14),
.B(n_13),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_31),
.Y(n_45)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_19),
.Y(n_32)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_32),
.A2(n_34),
.B1(n_25),
.B2(n_24),
.Y(n_54)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_20),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_33),
.B(n_40),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_SL g34 ( 
.A1(n_20),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_34)
);

INVx11_ASAP7_75t_L g35 ( 
.A(n_21),
.Y(n_35)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_35),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_24),
.B(n_25),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_36),
.B(n_38),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_19),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_37),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g38 ( 
.A(n_26),
.B(n_0),
.Y(n_38)
);

INVx5_ASAP7_75t_L g39 ( 
.A(n_20),
.Y(n_39)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_39),
.Y(n_50)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_19),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_41),
.B(n_27),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_39),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_42),
.B(n_43),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_39),
.Y(n_43)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_46),
.B(n_47),
.Y(n_76)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_40),
.Y(n_47)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_48),
.Y(n_74)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_31),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_49),
.Y(n_77)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_51),
.B(n_59),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

INVx5_ASAP7_75t_L g72 ( 
.A(n_52),
.Y(n_72)
);

CKINVDCx16_ASAP7_75t_R g71 ( 
.A(n_54),
.Y(n_71)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_33),
.Y(n_55)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_55),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_32),
.A2(n_40),
.B1(n_35),
.B2(n_33),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_L g66 ( 
.A1(n_58),
.A2(n_32),
.B1(n_35),
.B2(n_27),
.Y(n_66)
);

CKINVDCx16_ASAP7_75t_R g59 ( 
.A(n_31),
.Y(n_59)
);

INVx5_ASAP7_75t_L g60 ( 
.A(n_37),
.Y(n_60)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_60),
.Y(n_68)
);

AND2x2_ASAP7_75t_SL g61 ( 
.A(n_50),
.B(n_31),
.Y(n_61)
);

OAI21xp5_ASAP7_75t_SL g84 ( 
.A1(n_61),
.A2(n_50),
.B(n_31),
.Y(n_84)
);

AO22x1_ASAP7_75t_SL g62 ( 
.A1(n_54),
.A2(n_34),
.B1(n_32),
.B2(n_37),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_62),
.A2(n_69),
.B1(n_58),
.B2(n_28),
.Y(n_78)
);

A2O1A1Ixp33_ASAP7_75t_L g63 ( 
.A1(n_56),
.A2(n_38),
.B(n_29),
.C(n_18),
.Y(n_63)
);

AOI21xp5_ASAP7_75t_L g95 ( 
.A1(n_63),
.A2(n_45),
.B(n_15),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_66),
.A2(n_22),
.B1(n_21),
.B2(n_30),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_44),
.B(n_31),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_67),
.B(n_49),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_L g69 ( 
.A1(n_53),
.A2(n_17),
.B1(n_23),
.B2(n_18),
.Y(n_69)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_57),
.Y(n_70)
);

INVx11_ASAP7_75t_L g80 ( 
.A(n_70),
.Y(n_80)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_57),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_75),
.B(n_22),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_78),
.B(n_93),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_76),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_79),
.B(n_86),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_65),
.B(n_28),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_81),
.B(n_82),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_63),
.B(n_16),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_71),
.A2(n_53),
.B1(n_60),
.B2(n_55),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_83),
.A2(n_85),
.B1(n_87),
.B2(n_91),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_SL g101 ( 
.A1(n_84),
.A2(n_68),
.B(n_64),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_62),
.A2(n_43),
.B1(n_42),
.B2(n_23),
.Y(n_85)
);

CKINVDCx16_ASAP7_75t_R g86 ( 
.A(n_73),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_62),
.A2(n_17),
.B1(n_16),
.B2(n_52),
.Y(n_87)
);

CKINVDCx16_ASAP7_75t_R g88 ( 
.A(n_67),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_88),
.B(n_90),
.Y(n_103)
);

CKINVDCx14_ASAP7_75t_R g109 ( 
.A(n_89),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_77),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_61),
.A2(n_26),
.B1(n_22),
.B2(n_30),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_61),
.A2(n_41),
.B1(n_30),
.B2(n_21),
.Y(n_92)
);

CKINVDCx16_ASAP7_75t_R g114 ( 
.A(n_92),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_94),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_95),
.B(n_15),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_74),
.B(n_0),
.Y(n_96)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_96),
.Y(n_102)
);

BUFx4f_ASAP7_75t_SL g97 ( 
.A(n_80),
.Y(n_97)
);

HB1xp67_ASAP7_75t_L g118 ( 
.A(n_97),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_99),
.A2(n_95),
.B1(n_87),
.B2(n_86),
.Y(n_126)
);

INVx13_ASAP7_75t_L g100 ( 
.A(n_84),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_100),
.B(n_105),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_101),
.B(n_93),
.C(n_85),
.Y(n_119)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_80),
.Y(n_105)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_91),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_106),
.B(n_107),
.Y(n_120)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_83),
.Y(n_107)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_92),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_110),
.B(n_78),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_88),
.B(n_64),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_112),
.B(n_90),
.Y(n_129)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_97),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_116),
.B(n_121),
.Y(n_134)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_112),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_117),
.B(n_124),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_119),
.B(n_99),
.C(n_114),
.Y(n_136)
);

OR2x2_ASAP7_75t_L g121 ( 
.A(n_103),
.B(n_79),
.Y(n_121)
);

HB1xp67_ASAP7_75t_L g122 ( 
.A(n_97),
.Y(n_122)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_122),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_123),
.B(n_130),
.Y(n_138)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_111),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_108),
.B(n_81),
.Y(n_125)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_125),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g140 ( 
.A(n_126),
.B(n_98),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_108),
.B(n_82),
.Y(n_127)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_127),
.Y(n_133)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_97),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_128),
.Y(n_135)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_129),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_104),
.B(n_96),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_104),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_131),
.B(n_110),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_114),
.A2(n_68),
.B1(n_72),
.B2(n_75),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_132),
.A2(n_101),
.B1(n_107),
.B2(n_113),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_136),
.B(n_131),
.C(n_119),
.Y(n_153)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_139),
.Y(n_149)
);

XOR2xp5_ASAP7_75t_L g150 ( 
.A(n_140),
.B(n_136),
.Y(n_150)
);

INVx4_ASAP7_75t_L g141 ( 
.A(n_118),
.Y(n_141)
);

INVx13_ASAP7_75t_L g152 ( 
.A(n_141),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_SL g156 ( 
.A1(n_142),
.A2(n_124),
.B(n_121),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_117),
.B(n_104),
.Y(n_143)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_143),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_129),
.B(n_106),
.Y(n_144)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_144),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_130),
.B(n_98),
.Y(n_148)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_148),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_150),
.B(n_151),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_SL g151 ( 
.A(n_143),
.B(n_138),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_153),
.B(n_138),
.C(n_144),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_148),
.A2(n_115),
.B1(n_120),
.B2(n_113),
.Y(n_154)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_154),
.Y(n_167)
);

AOI21xp5_ASAP7_75t_L g166 ( 
.A1(n_156),
.A2(n_162),
.B(n_137),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_135),
.B(n_145),
.Y(n_157)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_157),
.Y(n_173)
);

BUFx2_ASAP7_75t_L g158 ( 
.A(n_141),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_158),
.B(n_159),
.Y(n_170)
);

NOR3xp33_ASAP7_75t_L g159 ( 
.A(n_134),
.B(n_100),
.C(n_102),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_SL g162 ( 
.A1(n_142),
.A2(n_116),
.B(n_132),
.Y(n_162)
);

NAND2xp33_ASAP7_75t_SL g163 ( 
.A(n_162),
.B(n_139),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_163),
.B(n_168),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_150),
.B(n_153),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_164),
.B(n_165),
.C(n_169),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_166),
.A2(n_160),
.B1(n_154),
.B2(n_102),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_149),
.A2(n_140),
.B1(n_137),
.B2(n_133),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_151),
.B(n_146),
.C(n_147),
.Y(n_169)
);

HB1xp67_ASAP7_75t_L g172 ( 
.A(n_158),
.Y(n_172)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_172),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_173),
.B(n_133),
.Y(n_176)
);

AOI21xp5_ASAP7_75t_L g185 ( 
.A1(n_176),
.A2(n_178),
.B(n_180),
.Y(n_185)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_170),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_171),
.B(n_155),
.C(n_161),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_179),
.B(n_175),
.C(n_174),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_169),
.B(n_156),
.Y(n_180)
);

AOI322xp5_ASAP7_75t_L g183 ( 
.A1(n_181),
.A2(n_165),
.A3(n_109),
.B1(n_171),
.B2(n_164),
.C1(n_152),
.C2(n_72),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_167),
.B(n_152),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_SL g188 ( 
.A1(n_182),
.A2(n_70),
.B(n_9),
.Y(n_188)
);

AOI21xp5_ASAP7_75t_L g190 ( 
.A1(n_183),
.A2(n_184),
.B(n_187),
.Y(n_190)
);

INVxp67_ASAP7_75t_L g184 ( 
.A(n_177),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_186),
.B(n_189),
.C(n_3),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_179),
.B(n_105),
.Y(n_187)
);

AOI21xp5_ASAP7_75t_L g194 ( 
.A1(n_188),
.A2(n_4),
.B(n_5),
.Y(n_194)
);

AOI322xp5_ASAP7_75t_L g189 ( 
.A1(n_175),
.A2(n_8),
.A3(n_12),
.B1(n_11),
.B2(n_45),
.C1(n_49),
.C2(n_7),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_184),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_191),
.B(n_193),
.C(n_194),
.Y(n_197)
);

INVxp67_ASAP7_75t_L g192 ( 
.A(n_185),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g196 ( 
.A(n_192),
.B(n_4),
.Y(n_196)
);

AND2x2_ASAP7_75t_L g195 ( 
.A(n_190),
.B(n_15),
.Y(n_195)
);

O2A1O1Ixp33_ASAP7_75t_L g198 ( 
.A1(n_195),
.A2(n_196),
.B(n_6),
.C(n_7),
.Y(n_198)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_198),
.Y(n_201)
);

INVxp67_ASAP7_75t_L g199 ( 
.A(n_197),
.Y(n_199)
);

MAJx2_ASAP7_75t_L g200 ( 
.A(n_199),
.B(n_6),
.C(n_7),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_200),
.B(n_201),
.Y(n_202)
);


endmodule