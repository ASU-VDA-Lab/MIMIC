module fake_jpeg_6139_n_29 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_29);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_29;

wire n_13;
wire n_21;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_14;
wire n_19;
wire n_20;
wire n_18;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_11;
wire n_17;
wire n_25;
wire n_12;
wire n_15;

AOI22xp33_ASAP7_75t_SL g10 ( 
.A1(n_3),
.A2(n_1),
.B1(n_5),
.B2(n_0),
.Y(n_10)
);

INVx2_ASAP7_75t_L g11 ( 
.A(n_6),
.Y(n_11)
);

INVx2_ASAP7_75t_L g12 ( 
.A(n_5),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_2),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_L g14 ( 
.A(n_6),
.B(n_7),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_8),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_4),
.B(n_3),
.Y(n_16)
);

AOI22xp33_ASAP7_75t_SL g17 ( 
.A1(n_4),
.A2(n_7),
.B1(n_9),
.B2(n_0),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_2),
.B(n_8),
.Y(n_18)
);

AO22x1_ASAP7_75t_SL g19 ( 
.A1(n_10),
.A2(n_0),
.B1(n_1),
.B2(n_9),
.Y(n_19)
);

XNOR2xp5_ASAP7_75t_L g25 ( 
.A(n_19),
.B(n_20),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_SL g20 ( 
.A1(n_17),
.A2(n_1),
.B1(n_11),
.B2(n_12),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_15),
.B(n_13),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_21),
.B(n_22),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_11),
.A2(n_12),
.B1(n_15),
.B2(n_13),
.Y(n_22)
);

XOR2xp5_ASAP7_75t_L g23 ( 
.A(n_14),
.B(n_18),
.Y(n_23)
);

AO221x1_ASAP7_75t_L g26 ( 
.A1(n_24),
.A2(n_19),
.B1(n_22),
.B2(n_20),
.C(n_14),
.Y(n_26)
);

OAI21x1_ASAP7_75t_L g28 ( 
.A1(n_26),
.A2(n_27),
.B(n_19),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_25),
.Y(n_27)
);

AOI322xp5_ASAP7_75t_L g29 ( 
.A1(n_28),
.A2(n_16),
.A3(n_18),
.B1(n_23),
.B2(n_25),
.C1(n_27),
.C2(n_26),
.Y(n_29)
);


endmodule