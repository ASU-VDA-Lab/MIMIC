module fake_netlist_5_639_n_2913 (n_137, n_294, n_431, n_318, n_380, n_419, n_444, n_469, n_82, n_194, n_316, n_389, n_549, n_418, n_248, n_124, n_86, n_136, n_146, n_315, n_268, n_523, n_451, n_532, n_408, n_61, n_376, n_503, n_127, n_75, n_235, n_226, n_74, n_515, n_57, n_353, n_351, n_367, n_452, n_397, n_493, n_111, n_525, n_483, n_544, n_155, n_552, n_547, n_43, n_116, n_22, n_467, n_423, n_284, n_46, n_245, n_21, n_501, n_139, n_38, n_105, n_280, n_4, n_378, n_551, n_17, n_382, n_554, n_254, n_33, n_23, n_302, n_265, n_526, n_293, n_372, n_443, n_244, n_47, n_173, n_198, n_447, n_247, n_314, n_368, n_433, n_8, n_321, n_292, n_100, n_455, n_417, n_212, n_385, n_498, n_516, n_507, n_119, n_497, n_275, n_252, n_26, n_295, n_133, n_330, n_508, n_506, n_2, n_6, n_509, n_39, n_147, n_373, n_67, n_307, n_439, n_87, n_150, n_530, n_106, n_209, n_259, n_448, n_375, n_301, n_68, n_93, n_186, n_537, n_134, n_191, n_51, n_63, n_492, n_171, n_153, n_524, n_399, n_341, n_204, n_394, n_250, n_548, n_543, n_260, n_298, n_320, n_518, n_505, n_286, n_122, n_282, n_331, n_10, n_24, n_406, n_519, n_470, n_325, n_449, n_132, n_90, n_546, n_101, n_281, n_240, n_381, n_189, n_220, n_291, n_231, n_257, n_390, n_31, n_456, n_13, n_371, n_481, n_535, n_152, n_540, n_317, n_9, n_323, n_195, n_42, n_356, n_227, n_45, n_271, n_94, n_335, n_123, n_370, n_167, n_234, n_343, n_308, n_379, n_428, n_267, n_514, n_457, n_297, n_156, n_5, n_225, n_377, n_484, n_219, n_442, n_157, n_131, n_192, n_223, n_392, n_158, n_138, n_264, n_109, n_472, n_454, n_387, n_374, n_163, n_276, n_339, n_95, n_183, n_185, n_243, n_398, n_396, n_347, n_169, n_59, n_522, n_550, n_255, n_215, n_350, n_196, n_459, n_211, n_218, n_400, n_181, n_436, n_3, n_290, n_221, n_178, n_386, n_287, n_344, n_473, n_422, n_475, n_72, n_104, n_41, n_415, n_56, n_141, n_485, n_496, n_355, n_486, n_15, n_336, n_145, n_48, n_521, n_50, n_337, n_430, n_313, n_88, n_479, n_528, n_510, n_216, n_168, n_395, n_164, n_432, n_553, n_311, n_208, n_142, n_214, n_328, n_140, n_299, n_303, n_369, n_296, n_241, n_357, n_184, n_446, n_445, n_65, n_78, n_144, n_114, n_96, n_165, n_468, n_499, n_213, n_129, n_342, n_482, n_517, n_98, n_361, n_464, n_363, n_402, n_413, n_197, n_107, n_69, n_236, n_388, n_1, n_249, n_304, n_329, n_203, n_274, n_384, n_460, n_80, n_35, n_73, n_277, n_92, n_19, n_338, n_149, n_477, n_461, n_333, n_309, n_30, n_512, n_14, n_84, n_462, n_130, n_322, n_258, n_29, n_79, n_151, n_25, n_306, n_458, n_288, n_188, n_190, n_201, n_263, n_471, n_44, n_224, n_40, n_34, n_228, n_283, n_383, n_474, n_112, n_542, n_85, n_463, n_488, n_502, n_239, n_466, n_420, n_489, n_55, n_49, n_310, n_54, n_504, n_511, n_12, n_465, n_76, n_358, n_362, n_170, n_332, n_27, n_77, n_102, n_161, n_273, n_349, n_270, n_230, n_81, n_118, n_279, n_70, n_253, n_261, n_174, n_289, n_172, n_206, n_217, n_440, n_478, n_545, n_441, n_450, n_312, n_476, n_429, n_534, n_345, n_210, n_494, n_365, n_91, n_176, n_182, n_143, n_83, n_354, n_480, n_237, n_425, n_513, n_407, n_527, n_180, n_340, n_207, n_37, n_346, n_393, n_229, n_108, n_487, n_495, n_437, n_66, n_177, n_60, n_403, n_453, n_421, n_16, n_0, n_58, n_405, n_18, n_359, n_490, n_117, n_326, n_233, n_404, n_205, n_366, n_113, n_246, n_179, n_125, n_410, n_269, n_529, n_128, n_285, n_412, n_120, n_232, n_327, n_135, n_126, n_202, n_266, n_272, n_491, n_427, n_193, n_251, n_352, n_53, n_160, n_426, n_520, n_409, n_500, n_154, n_62, n_148, n_71, n_300, n_435, n_159, n_334, n_541, n_391, n_434, n_539, n_175, n_538, n_262, n_238, n_99, n_411, n_414, n_319, n_364, n_20, n_536, n_531, n_121, n_242, n_360, n_36, n_200, n_162, n_64, n_222, n_28, n_89, n_438, n_115, n_324, n_416, n_199, n_187, n_32, n_401, n_103, n_348, n_97, n_166, n_11, n_424, n_7, n_256, n_305, n_533, n_52, n_278, n_110, n_2913);

input n_137;
input n_294;
input n_431;
input n_318;
input n_380;
input n_419;
input n_444;
input n_469;
input n_82;
input n_194;
input n_316;
input n_389;
input n_549;
input n_418;
input n_248;
input n_124;
input n_86;
input n_136;
input n_146;
input n_315;
input n_268;
input n_523;
input n_451;
input n_532;
input n_408;
input n_61;
input n_376;
input n_503;
input n_127;
input n_75;
input n_235;
input n_226;
input n_74;
input n_515;
input n_57;
input n_353;
input n_351;
input n_367;
input n_452;
input n_397;
input n_493;
input n_111;
input n_525;
input n_483;
input n_544;
input n_155;
input n_552;
input n_547;
input n_43;
input n_116;
input n_22;
input n_467;
input n_423;
input n_284;
input n_46;
input n_245;
input n_21;
input n_501;
input n_139;
input n_38;
input n_105;
input n_280;
input n_4;
input n_378;
input n_551;
input n_17;
input n_382;
input n_554;
input n_254;
input n_33;
input n_23;
input n_302;
input n_265;
input n_526;
input n_293;
input n_372;
input n_443;
input n_244;
input n_47;
input n_173;
input n_198;
input n_447;
input n_247;
input n_314;
input n_368;
input n_433;
input n_8;
input n_321;
input n_292;
input n_100;
input n_455;
input n_417;
input n_212;
input n_385;
input n_498;
input n_516;
input n_507;
input n_119;
input n_497;
input n_275;
input n_252;
input n_26;
input n_295;
input n_133;
input n_330;
input n_508;
input n_506;
input n_2;
input n_6;
input n_509;
input n_39;
input n_147;
input n_373;
input n_67;
input n_307;
input n_439;
input n_87;
input n_150;
input n_530;
input n_106;
input n_209;
input n_259;
input n_448;
input n_375;
input n_301;
input n_68;
input n_93;
input n_186;
input n_537;
input n_134;
input n_191;
input n_51;
input n_63;
input n_492;
input n_171;
input n_153;
input n_524;
input n_399;
input n_341;
input n_204;
input n_394;
input n_250;
input n_548;
input n_543;
input n_260;
input n_298;
input n_320;
input n_518;
input n_505;
input n_286;
input n_122;
input n_282;
input n_331;
input n_10;
input n_24;
input n_406;
input n_519;
input n_470;
input n_325;
input n_449;
input n_132;
input n_90;
input n_546;
input n_101;
input n_281;
input n_240;
input n_381;
input n_189;
input n_220;
input n_291;
input n_231;
input n_257;
input n_390;
input n_31;
input n_456;
input n_13;
input n_371;
input n_481;
input n_535;
input n_152;
input n_540;
input n_317;
input n_9;
input n_323;
input n_195;
input n_42;
input n_356;
input n_227;
input n_45;
input n_271;
input n_94;
input n_335;
input n_123;
input n_370;
input n_167;
input n_234;
input n_343;
input n_308;
input n_379;
input n_428;
input n_267;
input n_514;
input n_457;
input n_297;
input n_156;
input n_5;
input n_225;
input n_377;
input n_484;
input n_219;
input n_442;
input n_157;
input n_131;
input n_192;
input n_223;
input n_392;
input n_158;
input n_138;
input n_264;
input n_109;
input n_472;
input n_454;
input n_387;
input n_374;
input n_163;
input n_276;
input n_339;
input n_95;
input n_183;
input n_185;
input n_243;
input n_398;
input n_396;
input n_347;
input n_169;
input n_59;
input n_522;
input n_550;
input n_255;
input n_215;
input n_350;
input n_196;
input n_459;
input n_211;
input n_218;
input n_400;
input n_181;
input n_436;
input n_3;
input n_290;
input n_221;
input n_178;
input n_386;
input n_287;
input n_344;
input n_473;
input n_422;
input n_475;
input n_72;
input n_104;
input n_41;
input n_415;
input n_56;
input n_141;
input n_485;
input n_496;
input n_355;
input n_486;
input n_15;
input n_336;
input n_145;
input n_48;
input n_521;
input n_50;
input n_337;
input n_430;
input n_313;
input n_88;
input n_479;
input n_528;
input n_510;
input n_216;
input n_168;
input n_395;
input n_164;
input n_432;
input n_553;
input n_311;
input n_208;
input n_142;
input n_214;
input n_328;
input n_140;
input n_299;
input n_303;
input n_369;
input n_296;
input n_241;
input n_357;
input n_184;
input n_446;
input n_445;
input n_65;
input n_78;
input n_144;
input n_114;
input n_96;
input n_165;
input n_468;
input n_499;
input n_213;
input n_129;
input n_342;
input n_482;
input n_517;
input n_98;
input n_361;
input n_464;
input n_363;
input n_402;
input n_413;
input n_197;
input n_107;
input n_69;
input n_236;
input n_388;
input n_1;
input n_249;
input n_304;
input n_329;
input n_203;
input n_274;
input n_384;
input n_460;
input n_80;
input n_35;
input n_73;
input n_277;
input n_92;
input n_19;
input n_338;
input n_149;
input n_477;
input n_461;
input n_333;
input n_309;
input n_30;
input n_512;
input n_14;
input n_84;
input n_462;
input n_130;
input n_322;
input n_258;
input n_29;
input n_79;
input n_151;
input n_25;
input n_306;
input n_458;
input n_288;
input n_188;
input n_190;
input n_201;
input n_263;
input n_471;
input n_44;
input n_224;
input n_40;
input n_34;
input n_228;
input n_283;
input n_383;
input n_474;
input n_112;
input n_542;
input n_85;
input n_463;
input n_488;
input n_502;
input n_239;
input n_466;
input n_420;
input n_489;
input n_55;
input n_49;
input n_310;
input n_54;
input n_504;
input n_511;
input n_12;
input n_465;
input n_76;
input n_358;
input n_362;
input n_170;
input n_332;
input n_27;
input n_77;
input n_102;
input n_161;
input n_273;
input n_349;
input n_270;
input n_230;
input n_81;
input n_118;
input n_279;
input n_70;
input n_253;
input n_261;
input n_174;
input n_289;
input n_172;
input n_206;
input n_217;
input n_440;
input n_478;
input n_545;
input n_441;
input n_450;
input n_312;
input n_476;
input n_429;
input n_534;
input n_345;
input n_210;
input n_494;
input n_365;
input n_91;
input n_176;
input n_182;
input n_143;
input n_83;
input n_354;
input n_480;
input n_237;
input n_425;
input n_513;
input n_407;
input n_527;
input n_180;
input n_340;
input n_207;
input n_37;
input n_346;
input n_393;
input n_229;
input n_108;
input n_487;
input n_495;
input n_437;
input n_66;
input n_177;
input n_60;
input n_403;
input n_453;
input n_421;
input n_16;
input n_0;
input n_58;
input n_405;
input n_18;
input n_359;
input n_490;
input n_117;
input n_326;
input n_233;
input n_404;
input n_205;
input n_366;
input n_113;
input n_246;
input n_179;
input n_125;
input n_410;
input n_269;
input n_529;
input n_128;
input n_285;
input n_412;
input n_120;
input n_232;
input n_327;
input n_135;
input n_126;
input n_202;
input n_266;
input n_272;
input n_491;
input n_427;
input n_193;
input n_251;
input n_352;
input n_53;
input n_160;
input n_426;
input n_520;
input n_409;
input n_500;
input n_154;
input n_62;
input n_148;
input n_71;
input n_300;
input n_435;
input n_159;
input n_334;
input n_541;
input n_391;
input n_434;
input n_539;
input n_175;
input n_538;
input n_262;
input n_238;
input n_99;
input n_411;
input n_414;
input n_319;
input n_364;
input n_20;
input n_536;
input n_531;
input n_121;
input n_242;
input n_360;
input n_36;
input n_200;
input n_162;
input n_64;
input n_222;
input n_28;
input n_89;
input n_438;
input n_115;
input n_324;
input n_416;
input n_199;
input n_187;
input n_32;
input n_401;
input n_103;
input n_348;
input n_97;
input n_166;
input n_11;
input n_424;
input n_7;
input n_256;
input n_305;
input n_533;
input n_52;
input n_278;
input n_110;

output n_2913;

wire n_924;
wire n_1263;
wire n_1378;
wire n_977;
wire n_2253;
wire n_2417;
wire n_611;
wire n_2756;
wire n_1126;
wire n_1423;
wire n_1729;
wire n_2739;
wire n_1166;
wire n_2380;
wire n_1751;
wire n_1508;
wire n_2771;
wire n_785;
wire n_2617;
wire n_2200;
wire n_1161;
wire n_1859;
wire n_2746;
wire n_1677;
wire n_1150;
wire n_2327;
wire n_1780;
wire n_1488;
wire n_667;
wire n_2899;
wire n_790;
wire n_1055;
wire n_2386;
wire n_1501;
wire n_2395;
wire n_880;
wire n_1007;
wire n_2369;
wire n_1528;
wire n_2683;
wire n_1370;
wire n_1292;
wire n_2347;
wire n_2520;
wire n_2821;
wire n_1198;
wire n_1360;
wire n_2388;
wire n_1099;
wire n_2568;
wire n_956;
wire n_564;
wire n_1738;
wire n_2021;
wire n_2134;
wire n_2391;
wire n_1021;
wire n_1960;
wire n_2843;
wire n_2185;
wire n_2143;
wire n_2853;
wire n_2059;
wire n_1323;
wire n_1466;
wire n_1695;
wire n_688;
wire n_2487;
wire n_1353;
wire n_800;
wire n_1347;
wire n_2495;
wire n_2880;
wire n_1535;
wire n_1789;
wire n_1666;
wire n_2389;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_2302;
wire n_915;
wire n_1545;
wire n_2374;
wire n_864;
wire n_859;
wire n_951;
wire n_1947;
wire n_1264;
wire n_2114;
wire n_2001;
wire n_1494;
wire n_625;
wire n_1462;
wire n_854;
wire n_1799;
wire n_2069;
wire n_2396;
wire n_1580;
wire n_674;
wire n_1939;
wire n_2486;
wire n_1806;
wire n_933;
wire n_2244;
wire n_2257;
wire n_1152;
wire n_1869;
wire n_1607;
wire n_1563;
wire n_606;
wire n_2011;
wire n_2096;
wire n_877;
wire n_2105;
wire n_2538;
wire n_2024;
wire n_2530;
wire n_1696;
wire n_2483;
wire n_1118;
wire n_755;
wire n_1686;
wire n_947;
wire n_1285;
wire n_1860;
wire n_2543;
wire n_1359;
wire n_1107;
wire n_1728;
wire n_2031;
wire n_556;
wire n_2076;
wire n_2482;
wire n_2677;
wire n_1230;
wire n_668;
wire n_2165;
wire n_1896;
wire n_2147;
wire n_929;
wire n_2770;
wire n_1124;
wire n_1818;
wire n_2127;
wire n_1576;
wire n_902;
wire n_1104;
wire n_1294;
wire n_1705;
wire n_659;
wire n_2584;
wire n_1257;
wire n_2639;
wire n_1182;
wire n_579;
wire n_1698;
wire n_1261;
wire n_2329;
wire n_938;
wire n_1098;
wire n_2142;
wire n_1154;
wire n_2189;
wire n_1242;
wire n_1135;
wire n_2323;
wire n_2203;
wire n_2597;
wire n_1016;
wire n_1243;
wire n_2047;
wire n_1280;
wire n_1845;
wire n_2052;
wire n_2193;
wire n_2058;
wire n_2458;
wire n_2478;
wire n_2761;
wire n_731;
wire n_1483;
wire n_2888;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_1236;
wire n_1633;
wire n_2537;
wire n_569;
wire n_2669;
wire n_2144;
wire n_1778;
wire n_2306;
wire n_920;
wire n_2515;
wire n_1289;
wire n_1517;
wire n_2091;
wire n_2466;
wire n_2635;
wire n_2652;
wire n_2715;
wire n_2085;
wire n_1669;
wire n_2566;
wire n_976;
wire n_1949;
wire n_1449;
wire n_1946;
wire n_1566;
wire n_2032;
wire n_2587;
wire n_2149;
wire n_1078;
wire n_2782;
wire n_1670;
wire n_2672;
wire n_775;
wire n_2651;
wire n_600;
wire n_1484;
wire n_2071;
wire n_2561;
wire n_1374;
wire n_1328;
wire n_2643;
wire n_2141;
wire n_1948;
wire n_1984;
wire n_2099;
wire n_2408;
wire n_1877;
wire n_1831;
wire n_1598;
wire n_1723;
wire n_955;
wire n_1850;
wire n_1146;
wire n_882;
wire n_2384;
wire n_1036;
wire n_1097;
wire n_1749;
wire n_696;
wire n_897;
wire n_798;
wire n_646;
wire n_1428;
wire n_2663;
wire n_1394;
wire n_2659;
wire n_1414;
wire n_1216;
wire n_580;
wire n_2693;
wire n_1040;
wire n_2202;
wire n_2648;
wire n_1872;
wire n_1852;
wire n_2159;
wire n_578;
wire n_926;
wire n_2180;
wire n_2249;
wire n_2353;
wire n_1218;
wire n_1931;
wire n_2439;
wire n_2632;
wire n_2276;
wire n_1070;
wire n_1547;
wire n_777;
wire n_2089;
wire n_1030;
wire n_2470;
wire n_1755;
wire n_1071;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_1801;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_2908;
wire n_1600;
wire n_663;
wire n_845;
wire n_2235;
wire n_1862;
wire n_673;
wire n_837;
wire n_1239;
wire n_2300;
wire n_2791;
wire n_1796;
wire n_2551;
wire n_1473;
wire n_680;
wire n_1587;
wire n_2682;
wire n_901;
wire n_2432;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_2174;
wire n_2714;
wire n_1748;
wire n_1672;
wire n_2506;
wire n_675;
wire n_2699;
wire n_888;
wire n_1880;
wire n_2769;
wire n_2337;
wire n_1167;
wire n_1626;
wire n_637;
wire n_2615;
wire n_1384;
wire n_1556;
wire n_1863;
wire n_1064;
wire n_858;
wire n_2079;
wire n_2238;
wire n_923;
wire n_2118;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_2407;
wire n_1706;
wire n_2753;
wire n_1582;
wire n_1069;
wire n_1784;
wire n_2859;
wire n_2842;
wire n_1075;
wire n_1836;
wire n_2868;
wire n_1450;
wire n_1322;
wire n_2101;
wire n_1471;
wire n_1986;
wire n_2863;
wire n_2072;
wire n_2738;
wire n_1750;
wire n_1459;
wire n_889;
wire n_2358;
wire n_973;
wire n_1700;
wire n_2833;
wire n_571;
wire n_1585;
wire n_2684;
wire n_2712;
wire n_1971;
wire n_1599;
wire n_2275;
wire n_2855;
wire n_2713;
wire n_2644;
wire n_2700;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_2730;
wire n_1950;
wire n_1447;
wire n_907;
wire n_2251;
wire n_1377;
wire n_2370;
wire n_989;
wire n_2544;
wire n_1039;
wire n_2214;
wire n_2055;
wire n_1403;
wire n_2248;
wire n_2356;
wire n_736;
wire n_892;
wire n_2688;
wire n_1000;
wire n_1202;
wire n_2750;
wire n_2620;
wire n_1278;
wire n_2622;
wire n_2062;
wire n_2668;
wire n_1463;
wire n_1002;
wire n_1581;
wire n_2100;
wire n_593;
wire n_2258;
wire n_748;
wire n_1058;
wire n_586;
wire n_1667;
wire n_838;
wire n_2784;
wire n_1053;
wire n_1224;
wire n_2865;
wire n_2557;
wire n_1926;
wire n_2706;
wire n_1248;
wire n_1331;
wire n_953;
wire n_1014;
wire n_1241;
wire n_2150;
wire n_2241;
wire n_2757;
wire n_2152;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_793;
wire n_2590;
wire n_2776;
wire n_2140;
wire n_2385;
wire n_1819;
wire n_2330;
wire n_2139;
wire n_1527;
wire n_2042;
wire n_1882;
wire n_884;
wire n_944;
wire n_1754;
wire n_1623;
wire n_2862;
wire n_2175;
wire n_2720;
wire n_2324;
wire n_1854;
wire n_2606;
wire n_2674;
wire n_1565;
wire n_2828;
wire n_1809;
wire n_1856;
wire n_647;
wire n_1072;
wire n_2218;
wire n_2267;
wire n_832;
wire n_857;
wire n_2305;
wire n_2636;
wire n_2450;
wire n_561;
wire n_1319;
wire n_2379;
wire n_2616;
wire n_2911;
wire n_2154;
wire n_1825;
wire n_1951;
wire n_1906;
wire n_1883;
wire n_2759;
wire n_1712;
wire n_1387;
wire n_2262;
wire n_2462;
wire n_2514;
wire n_1532;
wire n_2322;
wire n_2271;
wire n_2625;
wire n_1027;
wire n_971;
wire n_1156;
wire n_794;
wire n_2798;
wire n_2331;
wire n_2293;
wire n_686;
wire n_2837;
wire n_847;
wire n_1393;
wire n_2319;
wire n_596;
wire n_1775;
wire n_2028;
wire n_1368;
wire n_2762;
wire n_558;
wire n_2808;
wire n_1276;
wire n_702;
wire n_2548;
wire n_822;
wire n_1412;
wire n_2679;
wire n_1709;
wire n_2676;
wire n_2108;
wire n_728;
wire n_1162;
wire n_1538;
wire n_1838;
wire n_1199;
wire n_1847;
wire n_1779;
wire n_2767;
wire n_2777;
wire n_2603;
wire n_1884;
wire n_2434;
wire n_2660;
wire n_1038;
wire n_1369;
wire n_2611;
wire n_1841;
wire n_1660;
wire n_887;
wire n_1905;
wire n_2553;
wire n_2581;
wire n_2195;
wire n_2529;
wire n_2698;
wire n_809;
wire n_1711;
wire n_870;
wire n_599;
wire n_1891;
wire n_1662;
wire n_931;
wire n_1481;
wire n_2626;
wire n_1942;
wire n_1978;
wire n_1544;
wire n_2510;
wire n_868;
wire n_2454;
wire n_639;
wire n_2804;
wire n_914;
wire n_2120;
wire n_2546;
wire n_1629;
wire n_1293;
wire n_2801;
wire n_965;
wire n_1876;
wire n_1743;
wire n_935;
wire n_1175;
wire n_817;
wire n_2763;
wire n_1479;
wire n_1810;
wire n_2350;
wire n_2813;
wire n_2825;
wire n_2009;
wire n_1888;
wire n_759;
wire n_2222;
wire n_1892;
wire n_806;
wire n_1997;
wire n_2667;
wire n_1766;
wire n_1477;
wire n_1635;
wire n_1963;
wire n_2226;
wire n_1571;
wire n_2891;
wire n_1189;
wire n_2690;
wire n_2215;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_2064;
wire n_784;
wire n_2449;
wire n_1733;
wire n_1244;
wire n_2413;
wire n_1194;
wire n_1925;
wire n_2297;
wire n_1815;
wire n_2621;
wire n_615;
wire n_851;
wire n_1759;
wire n_1788;
wire n_843;
wire n_2177;
wire n_2491;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_2227;
wire n_678;
wire n_2671;
wire n_697;
wire n_1222;
wire n_1679;
wire n_2190;
wire n_776;
wire n_2022;
wire n_1798;
wire n_1790;
wire n_2518;
wire n_2876;
wire n_1415;
wire n_2629;
wire n_2592;
wire n_1260;
wire n_1746;
wire n_1647;
wire n_2181;
wire n_2479;
wire n_2838;
wire n_1829;
wire n_1464;
wire n_649;
wire n_2563;
wire n_1444;
wire n_1191;
wire n_2387;
wire n_1674;
wire n_1833;
wire n_1830;
wire n_2517;
wire n_2073;
wire n_1710;
wire n_1128;
wire n_1734;
wire n_744;
wire n_590;
wire n_629;
wire n_2631;
wire n_1308;
wire n_2871;
wire n_2178;
wire n_1767;
wire n_2336;
wire n_1680;
wire n_1233;
wire n_2607;
wire n_1615;
wire n_1529;
wire n_2005;
wire n_1916;
wire n_677;
wire n_1333;
wire n_2469;
wire n_1121;
wire n_2723;
wire n_604;
wire n_2007;
wire n_949;
wire n_2539;
wire n_2582;
wire n_1443;
wire n_1008;
wire n_1539;
wire n_946;
wire n_2736;
wire n_1001;
wire n_1503;
wire n_2054;
wire n_1468;
wire n_1559;
wire n_1765;
wire n_1866;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_624;
wire n_1380;
wire n_1744;
wire n_2623;
wire n_1617;
wire n_1010;
wire n_1994;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_2718;
wire n_1195;
wire n_1837;
wire n_1839;
wire n_610;
wire n_2577;
wire n_1760;
wire n_2875;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_2796;
wire n_757;
wire n_2342;
wire n_633;
wire n_2856;
wire n_1832;
wire n_1851;
wire n_758;
wire n_999;
wire n_2046;
wire n_2848;
wire n_2741;
wire n_1933;
wire n_2290;
wire n_1656;
wire n_1158;
wire n_2045;
wire n_1509;
wire n_1874;
wire n_2040;
wire n_563;
wire n_2060;
wire n_2613;
wire n_1987;
wire n_2805;
wire n_1145;
wire n_878;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_2145;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_1871;
wire n_2580;
wire n_2545;
wire n_2787;
wire n_1964;
wire n_2869;
wire n_1163;
wire n_906;
wire n_2039;
wire n_1207;
wire n_919;
wire n_908;
wire n_2412;
wire n_2406;
wire n_2846;
wire n_724;
wire n_1781;
wire n_2084;
wire n_2035;
wire n_658;
wire n_2061;
wire n_2378;
wire n_2509;
wire n_1740;
wire n_2398;
wire n_1362;
wire n_2857;
wire n_1586;
wire n_959;
wire n_2459;
wire n_940;
wire n_1445;
wire n_1492;
wire n_2155;
wire n_2516;
wire n_1923;
wire n_1773;
wire n_592;
wire n_1169;
wire n_1596;
wire n_1692;
wire n_2666;
wire n_1017;
wire n_2481;
wire n_2171;
wire n_978;
wire n_2768;
wire n_2116;
wire n_2314;
wire n_1434;
wire n_1054;
wire n_2507;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_2420;
wire n_2900;
wire n_1095;
wire n_1828;
wire n_1614;
wire n_2886;
wire n_2093;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_2339;
wire n_2038;
wire n_2320;
wire n_2473;
wire n_2137;
wire n_603;
wire n_1431;
wire n_2583;
wire n_1593;
wire n_1033;
wire n_2299;
wire n_2540;
wire n_2873;
wire n_636;
wire n_660;
wire n_2087;
wire n_1640;
wire n_2162;
wire n_1732;
wire n_1009;
wire n_2847;
wire n_1148;
wire n_2051;
wire n_742;
wire n_2029;
wire n_750;
wire n_995;
wire n_2168;
wire n_2790;
wire n_1609;
wire n_1989;
wire n_2359;
wire n_1887;
wire n_2523;
wire n_1383;
wire n_1073;
wire n_2346;
wire n_2457;
wire n_662;
wire n_2312;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1920;
wire n_1065;
wire n_1592;
wire n_2536;
wire n_1336;
wire n_2882;
wire n_1721;
wire n_1959;
wire n_1758;
wire n_2338;
wire n_2737;
wire n_1574;
wire n_2399;
wire n_2812;
wire n_2048;
wire n_2355;
wire n_2133;
wire n_1921;
wire n_2721;
wire n_1309;
wire n_1878;
wire n_1426;
wire n_1043;
wire n_2585;
wire n_1800;
wire n_1548;
wire n_2725;
wire n_614;
wire n_1421;
wire n_2571;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_974;
wire n_2565;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_2124;
wire n_743;
wire n_2081;
wire n_613;
wire n_1119;
wire n_2156;
wire n_1240;
wire n_2261;
wire n_1820;
wire n_2729;
wire n_2418;
wire n_829;
wire n_2519;
wire n_2724;
wire n_1612;
wire n_2179;
wire n_1416;
wire n_2077;
wire n_2897;
wire n_2909;
wire n_1724;
wire n_2111;
wire n_2521;
wire n_1237;
wire n_700;
wire n_573;
wire n_1420;
wire n_1132;
wire n_1366;
wire n_1300;
wire n_2595;
wire n_1127;
wire n_2277;
wire n_761;
wire n_2477;
wire n_1785;
wire n_1568;
wire n_2829;
wire n_1006;
wire n_2110;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_2231;
wire n_1390;
wire n_2017;
wire n_2474;
wire n_2879;
wire n_2604;
wire n_2090;
wire n_1870;
wire n_2367;
wire n_1591;
wire n_2033;
wire n_1682;
wire n_1980;
wire n_2390;
wire n_2628;
wire n_1249;
wire n_2896;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1927;
wire n_2132;
wire n_1349;
wire n_1093;
wire n_2400;
wire n_1031;
wire n_609;
wire n_1041;
wire n_1265;
wire n_1909;
wire n_2681;
wire n_1562;
wire n_834;
wire n_765;
wire n_2255;
wire n_2424;
wire n_2272;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_1965;
wire n_630;
wire n_1902;
wire n_2151;
wire n_1941;
wire n_2106;
wire n_2775;
wire n_2716;
wire n_1913;
wire n_2878;
wire n_1823;
wire n_874;
wire n_2464;
wire n_1101;
wire n_2831;
wire n_1106;
wire n_1456;
wire n_2230;
wire n_2015;
wire n_2365;
wire n_1982;
wire n_1875;
wire n_1304;
wire n_2803;
wire n_1324;
wire n_2851;
wire n_987;
wire n_1846;
wire n_2066;
wire n_1885;
wire n_1455;
wire n_767;
wire n_993;
wire n_1903;
wire n_2490;
wire n_1407;
wire n_2452;
wire n_1551;
wire n_860;
wire n_2849;
wire n_1805;
wire n_2176;
wire n_2204;
wire n_2905;
wire n_1816;
wire n_948;
wire n_1217;
wire n_2220;
wire n_2455;
wire n_628;
wire n_1849;
wire n_2410;
wire n_1131;
wire n_729;
wire n_1084;
wire n_1961;
wire n_970;
wire n_1935;
wire n_911;
wire n_1430;
wire n_2645;
wire n_2467;
wire n_2727;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_2288;
wire n_1351;
wire n_2240;
wire n_2696;
wire n_1044;
wire n_1205;
wire n_2436;
wire n_1209;
wire n_1552;
wire n_2508;
wire n_602;
wire n_574;
wire n_2593;
wire n_1435;
wire n_879;
wire n_2416;
wire n_2405;
wire n_623;
wire n_2088;
wire n_824;
wire n_1645;
wire n_2461;
wire n_1327;
wire n_2858;
wire n_2243;
wire n_996;
wire n_921;
wire n_1684;
wire n_2658;
wire n_1717;
wire n_572;
wire n_2895;
wire n_815;
wire n_1795;
wire n_2128;
wire n_2578;
wire n_1821;
wire n_1381;
wire n_2555;
wire n_2662;
wire n_2740;
wire n_1611;
wire n_1037;
wire n_2368;
wire n_2656;
wire n_1080;
wire n_2301;
wire n_1274;
wire n_2890;
wire n_2554;
wire n_1316;
wire n_1708;
wire n_2419;
wire n_1438;
wire n_1082;
wire n_1840;
wire n_589;
wire n_1630;
wire n_2122;
wire n_716;
wire n_2512;
wire n_562;
wire n_1436;
wire n_1691;
wire n_952;
wire n_2786;
wire n_2534;
wire n_2092;
wire n_1229;
wire n_701;
wire n_1437;
wire n_1023;
wire n_2075;
wire n_645;
wire n_803;
wire n_1092;
wire n_2694;
wire n_1776;
wire n_2198;
wire n_2610;
wire n_2661;
wire n_2572;
wire n_2281;
wire n_2131;
wire n_2789;
wire n_2216;
wire n_1757;
wire n_890;
wire n_1897;
wire n_764;
wire n_1919;
wire n_1056;
wire n_1424;
wire n_960;
wire n_2308;
wire n_1893;
wire n_2910;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_2053;
wire n_2163;
wire n_634;
wire n_2328;
wire n_1958;
wire n_2254;
wire n_1252;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_2647;
wire n_1311;
wire n_2191;
wire n_2864;
wire n_1519;
wire n_950;
wire n_2428;
wire n_1553;
wire n_2664;
wire n_1811;
wire n_2443;
wire n_2624;
wire n_1346;
wire n_1299;
wire n_2158;
wire n_1808;
wire n_1060;
wire n_1141;
wire n_2266;
wire n_2465;
wire n_2824;
wire n_2650;
wire n_912;
wire n_968;
wire n_619;
wire n_2440;
wire n_1386;
wire n_1699;
wire n_967;
wire n_1442;
wire n_2541;
wire n_1139;
wire n_2731;
wire n_2333;
wire n_885;
wire n_1432;
wire n_1357;
wire n_2125;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_2402;
wire n_1157;
wire n_2403;
wire n_1050;
wire n_841;
wire n_802;
wire n_1954;
wire n_2265;
wire n_1608;
wire n_983;
wire n_1844;
wire n_2760;
wire n_2792;
wire n_2870;
wire n_1305;
wire n_873;
wire n_1826;
wire n_1112;
wire n_2304;
wire n_1283;
wire n_762;
wire n_1644;
wire n_2334;
wire n_2637;
wire n_690;
wire n_1974;
wire n_2463;
wire n_583;
wire n_2086;
wire n_2289;
wire n_1343;
wire n_2701;
wire n_2783;
wire n_2263;
wire n_2881;
wire n_1203;
wire n_1631;
wire n_2472;
wire n_821;
wire n_1763;
wire n_2341;
wire n_1966;
wire n_1768;
wire n_2294;
wire n_1179;
wire n_621;
wire n_753;
wire n_2475;
wire n_2733;
wire n_1048;
wire n_1719;
wire n_1288;
wire n_2785;
wire n_2556;
wire n_2269;
wire n_2732;
wire n_2309;
wire n_2415;
wire n_2646;
wire n_1560;
wire n_1605;
wire n_2236;
wire n_1228;
wire n_2816;
wire n_2123;
wire n_972;
wire n_692;
wire n_2037;
wire n_2685;
wire n_1953;
wire n_1938;
wire n_820;
wire n_1200;
wire n_2499;
wire n_1911;
wire n_2460;
wire n_2589;
wire n_1301;
wire n_1363;
wire n_1668;
wire n_1185;
wire n_991;
wire n_2903;
wire n_828;
wire n_1967;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_2233;
wire n_1329;
wire n_2743;
wire n_2675;
wire n_1312;
wire n_1439;
wire n_804;
wire n_2827;
wire n_1688;
wire n_945;
wire n_1504;
wire n_943;
wire n_992;
wire n_1932;
wire n_2755;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_2082;
wire n_1992;
wire n_2429;
wire n_1643;
wire n_1983;
wire n_883;
wire n_1594;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_2362;
wire n_856;
wire n_2609;
wire n_1793;
wire n_1976;
wire n_2223;
wire n_918;
wire n_942;
wire n_2169;
wire n_1804;
wire n_1147;
wire n_1557;
wire n_1977;
wire n_2153;
wire n_2468;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_2364;
wire n_2533;
wire n_618;
wire n_896;
wire n_2310;
wire n_2780;
wire n_2287;
wire n_2860;
wire n_2291;
wire n_2596;
wire n_1636;
wire n_894;
wire n_2056;
wire n_1730;
wire n_831;
wire n_2280;
wire n_2192;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1865;
wire n_1470;
wire n_1096;
wire n_2094;
wire n_2670;
wire n_1575;
wire n_1735;
wire n_1697;
wire n_2318;
wire n_833;
wire n_2393;
wire n_2020;
wire n_1646;
wire n_2502;
wire n_2504;
wire n_1307;
wire n_1881;
wire n_988;
wire n_2749;
wire n_2043;
wire n_2901;
wire n_1940;
wire n_814;
wire n_2707;
wire n_2751;
wire n_2793;
wire n_1549;
wire n_1934;
wire n_2311;
wire n_1201;
wire n_1114;
wire n_655;
wire n_2025;
wire n_1616;
wire n_1446;
wire n_2285;
wire n_2758;
wire n_1458;
wire n_669;
wire n_1176;
wire n_1472;
wire n_2298;
wire n_2471;
wire n_1807;
wire n_1149;
wire n_2618;
wire n_1671;
wire n_635;
wire n_2559;
wire n_763;
wire n_1020;
wire n_1062;
wire n_2303;
wire n_1824;
wire n_1917;
wire n_2295;
wire n_1219;
wire n_1204;
wire n_2840;
wire n_2810;
wire n_2325;
wire n_2747;
wire n_2446;
wire n_1814;
wire n_1035;
wire n_2822;
wire n_555;
wire n_783;
wire n_1848;
wire n_1928;
wire n_2126;
wire n_2893;
wire n_1188;
wire n_2588;
wire n_1722;
wire n_661;
wire n_2441;
wire n_1802;
wire n_2600;
wire n_849;
wire n_2795;
wire n_584;
wire n_681;
wire n_1638;
wire n_1786;
wire n_2002;
wire n_2282;
wire n_2800;
wire n_2371;
wire n_830;
wire n_2098;
wire n_1296;
wire n_2627;
wire n_2352;
wire n_1413;
wire n_801;
wire n_2207;
wire n_2080;
wire n_2377;
wire n_2619;
wire n_2340;
wire n_2444;
wire n_2068;
wire n_875;
wire n_1110;
wire n_1655;
wire n_2641;
wire n_749;
wire n_1895;
wire n_2574;
wire n_1134;
wire n_1358;
wire n_717;
wire n_939;
wire n_2361;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_2638;
wire n_866;
wire n_1401;
wire n_969;
wire n_2492;
wire n_1019;
wire n_1105;
wire n_1998;
wire n_1338;
wire n_577;
wire n_2016;
wire n_1522;
wire n_1687;
wire n_1637;
wire n_2034;
wire n_1419;
wire n_2711;
wire n_1653;
wire n_693;
wire n_2270;
wire n_1506;
wire n_2653;
wire n_836;
wire n_990;
wire n_2867;
wire n_2496;
wire n_1886;
wire n_1389;
wire n_1894;
wire n_975;
wire n_1908;
wire n_1256;
wire n_1702;
wire n_2259;
wire n_2794;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_2608;
wire n_2657;
wire n_770;
wire n_1375;
wire n_2494;
wire n_2649;
wire n_1102;
wire n_2852;
wire n_2392;
wire n_1843;
wire n_711;
wire n_1499;
wire n_1187;
wire n_2633;
wire n_1441;
wire n_2522;
wire n_2435;
wire n_1392;
wire n_1597;
wire n_1929;
wire n_2807;
wire n_1164;
wire n_1659;
wire n_2097;
wire n_1834;
wire n_2313;
wire n_2542;
wire n_1174;
wire n_2431;
wire n_2835;
wire n_2558;
wire n_1371;
wire n_617;
wire n_1303;
wire n_2206;
wire n_2063;
wire n_1572;
wire n_1968;
wire n_2564;
wire n_2252;
wire n_1516;
wire n_876;
wire n_1190;
wire n_1736;
wire n_1685;
wire n_2409;
wire n_601;
wire n_917;
wire n_1714;
wire n_966;
wire n_1116;
wire n_2000;
wire n_1661;
wire n_1212;
wire n_2074;
wire n_1541;
wire n_2576;
wire n_726;
wire n_982;
wire n_2575;
wire n_1573;
wire n_1453;
wire n_1731;
wire n_2217;
wire n_818;
wire n_2373;
wire n_1970;
wire n_861;
wire n_1713;
wire n_1183;
wire n_2307;
wire n_2766;
wire n_1658;
wire n_899;
wire n_1253;
wire n_1737;
wire n_2201;
wire n_2722;
wire n_2117;
wire n_2745;
wire n_1904;
wire n_2640;
wire n_1993;
wire n_774;
wire n_1628;
wire n_2493;
wire n_2205;
wire n_1335;
wire n_1514;
wire n_1777;
wire n_1957;
wire n_1059;
wire n_1345;
wire n_1133;
wire n_1912;
wire n_1771;
wire n_1899;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_2067;
wire n_1168;
wire n_707;
wire n_2219;
wire n_2437;
wire n_2885;
wire n_2877;
wire n_2148;
wire n_937;
wire n_2445;
wire n_1427;
wire n_2779;
wire n_1584;
wire n_665;
wire n_1835;
wire n_1726;
wire n_1440;
wire n_2164;
wire n_1988;
wire n_2115;
wire n_1853;
wire n_1356;
wire n_2845;
wire n_1787;
wire n_2634;
wire n_2232;
wire n_910;
wire n_2212;
wire n_2602;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1774;
wire n_1725;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_2811;
wire n_1496;
wire n_1125;
wire n_2547;
wire n_708;
wire n_1812;
wire n_735;
wire n_2501;
wire n_1915;
wire n_1109;
wire n_895;
wire n_2532;
wire n_1310;
wire n_2605;
wire n_2121;
wire n_1803;
wire n_2665;
wire n_1399;
wire n_1543;
wire n_1991;
wire n_1979;
wire n_791;
wire n_732;
wire n_1533;
wire n_2224;
wire n_808;
wire n_2484;
wire n_797;
wire n_1025;
wire n_1930;
wire n_1955;
wire n_2765;
wire n_1067;
wire n_1720;
wire n_2830;
wire n_2401;
wire n_2003;
wire n_1457;
wire n_766;
wire n_2692;
wire n_2354;
wire n_2246;
wire n_2008;
wire n_1117;
wire n_799;
wire n_2264;
wire n_2754;
wire n_687;
wire n_715;
wire n_1742;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_2489;
wire n_1266;
wire n_872;
wire n_2012;
wire n_594;
wire n_1291;
wire n_1297;
wire n_1753;
wire n_2283;
wire n_2866;
wire n_1782;
wire n_2245;
wire n_1155;
wire n_1418;
wire n_1972;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_2806;
wire n_1011;
wire n_1184;
wire n_2184;
wire n_985;
wire n_1855;
wire n_2425;
wire n_869;
wire n_810;
wire n_827;
wire n_1703;
wire n_1352;
wire n_626;
wire n_2197;
wire n_2199;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_2814;
wire n_1170;
wire n_2213;
wire n_2023;
wire n_2351;
wire n_2211;
wire n_2095;
wire n_676;
wire n_2103;
wire n_653;
wire n_2160;
wire n_642;
wire n_2228;
wire n_2527;
wire n_1602;
wire n_2498;
wire n_1178;
wire n_855;
wire n_1461;
wire n_2697;
wire n_850;
wire n_684;
wire n_2421;
wire n_2286;
wire n_2902;
wire n_664;
wire n_1999;
wire n_2372;
wire n_2065;
wire n_2136;
wire n_2480;
wire n_1372;
wire n_2861;
wire n_605;
wire n_2630;
wire n_1273;
wire n_1822;
wire n_620;
wire n_643;
wire n_2363;
wire n_2430;
wire n_916;
wire n_1081;
wire n_2549;
wire n_2705;
wire n_2332;
wire n_1235;
wire n_980;
wire n_1115;
wire n_698;
wire n_703;
wire n_2433;
wire n_1282;
wire n_1318;
wire n_1783;
wire n_780;
wire n_2601;
wire n_998;
wire n_2375;
wire n_2550;
wire n_1454;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_1907;
wire n_823;
wire n_2686;
wire n_2528;
wire n_725;
wire n_2344;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_2836;
wire n_2316;
wire n_672;
wire n_1985;
wire n_1898;
wire n_2107;
wire n_581;
wire n_2906;
wire n_1625;
wire n_2130;
wire n_2187;
wire n_2284;
wire n_898;
wire n_2817;
wire n_2773;
wire n_2598;
wire n_1762;
wire n_1013;
wire n_1452;
wire n_718;
wire n_2687;
wire n_1120;
wire n_719;
wire n_1791;
wire n_1890;
wire n_1747;
wire n_714;
wire n_2850;
wire n_1683;
wire n_1944;
wire n_909;
wire n_1817;
wire n_1497;
wire n_1530;
wire n_2654;
wire n_997;
wire n_932;
wire n_612;
wire n_2078;
wire n_1409;
wire n_788;
wire n_1326;
wire n_2884;
wire n_1268;
wire n_559;
wire n_825;
wire n_2819;
wire n_1981;
wire n_2186;
wire n_1320;
wire n_1663;
wire n_737;
wire n_1718;
wire n_986;
wire n_2315;
wire n_1317;
wire n_1518;
wire n_1715;
wire n_2102;
wire n_2562;
wire n_1281;
wire n_1952;
wire n_1192;
wire n_2221;
wire n_1024;
wire n_1063;
wire n_1889;
wire n_1792;
wire n_1564;
wire n_1868;
wire n_1613;
wire n_1489;
wire n_733;
wire n_1922;
wire n_1376;
wire n_941;
wire n_2326;
wire n_981;
wire n_2560;
wire n_1569;
wire n_2188;
wire n_867;
wire n_2348;
wire n_2422;
wire n_2239;
wire n_587;
wire n_792;
wire n_1429;
wire n_756;
wire n_1238;
wire n_2448;
wire n_812;
wire n_2104;
wire n_2748;
wire n_2057;
wire n_1772;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_2898;
wire n_782;
wire n_2717;
wire n_2818;
wire n_1100;
wire n_2129;
wire n_1861;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1901;
wire n_1900;
wire n_1620;
wire n_2889;
wire n_1330;
wire n_1867;
wire n_1945;
wire n_2772;
wire n_1675;
wire n_1924;
wire n_2573;
wire n_1727;
wire n_2710;
wire n_1554;
wire n_1745;
wire n_2735;
wire n_769;
wire n_2497;
wire n_2006;
wire n_2844;
wire n_1995;
wire n_2411;
wire n_2138;
wire n_1046;
wire n_934;
wire n_1618;
wire n_2260;
wire n_826;
wire n_2343;
wire n_1813;
wire n_2447;
wire n_886;
wire n_2014;
wire n_1221;
wire n_2345;
wire n_654;
wire n_1172;
wire n_2535;
wire n_1341;
wire n_2726;
wire n_570;
wire n_2774;
wire n_1641;
wire n_1361;
wire n_2382;
wire n_1707;
wire n_853;
wire n_2317;
wire n_751;
wire n_2799;
wire n_2172;
wire n_1973;
wire n_1083;
wire n_786;
wire n_1142;
wire n_2376;
wire n_2488;
wire n_1129;
wire n_2579;
wire n_2476;
wire n_704;
wire n_787;
wire n_1770;
wire n_2781;
wire n_2456;
wire n_961;
wire n_2250;
wire n_2678;
wire n_1756;
wire n_771;
wire n_2778;
wire n_1716;
wire n_2788;
wire n_2872;
wire n_1225;
wire n_1520;
wire n_2451;
wire n_2887;
wire n_1287;
wire n_1262;
wire n_2691;
wire n_930;
wire n_1873;
wire n_1411;
wire n_622;
wire n_1962;
wire n_1577;
wire n_2423;
wire n_1087;
wire n_2526;
wire n_2854;
wire n_994;
wire n_1701;
wire n_2194;
wire n_848;
wire n_1550;
wire n_2874;
wire n_2764;
wire n_2703;
wire n_1498;
wire n_2167;
wire n_1223;
wire n_1272;
wire n_2680;
wire n_1567;
wire n_682;
wire n_2567;
wire n_1247;
wire n_2709;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1857;
wire n_1344;
wire n_2041;
wire n_631;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_1797;
wire n_1769;
wire n_839;
wire n_1210;
wire n_1364;
wire n_2357;
wire n_2183;
wire n_2673;
wire n_2742;
wire n_2360;
wire n_2292;
wire n_1250;
wire n_2173;
wire n_1842;
wire n_871;
wire n_2442;
wire n_598;
wire n_685;
wire n_608;
wire n_1367;
wire n_928;
wire n_1943;
wire n_1460;
wire n_772;
wire n_2018;
wire n_1555;
wire n_2834;
wire n_2531;
wire n_1589;
wire n_1086;
wire n_2702;
wire n_2570;
wire n_796;
wire n_1858;
wire n_1619;
wire n_2815;
wire n_2119;
wire n_1502;
wire n_2157;
wire n_2552;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_2744;
wire n_1348;
wire n_2030;
wire n_903;
wire n_2453;
wire n_1525;
wire n_2397;
wire n_1752;
wire n_740;
wire n_2883;
wire n_2208;
wire n_1404;
wire n_2912;
wire n_1794;
wire n_2182;
wire n_1315;
wire n_2234;
wire n_1061;
wire n_1910;
wire n_1298;
wire n_1652;
wire n_2209;
wire n_2050;
wire n_2809;
wire n_1193;
wire n_2797;
wire n_1676;
wire n_1255;
wire n_1113;
wire n_2321;
wire n_1226;
wire n_1277;
wire n_722;
wire n_2591;
wire n_2146;
wire n_844;
wire n_852;
wire n_1487;
wire n_1864;
wire n_1028;
wire n_1601;
wire n_781;
wire n_1546;
wire n_595;
wire n_2612;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_2841;
wire n_1627;
wire n_1245;
wire n_846;
wire n_2427;
wire n_2438;
wire n_2505;
wire n_1673;
wire n_2832;
wire n_1321;
wire n_1975;
wire n_2296;
wire n_2070;
wire n_1937;
wire n_585;
wire n_2112;
wire n_1739;
wire n_616;
wire n_2278;
wire n_2594;
wire n_2394;
wire n_1914;
wire n_2135;
wire n_2335;
wire n_2904;
wire n_745;
wire n_2381;
wire n_1654;
wire n_2569;
wire n_2349;
wire n_1103;
wire n_648;
wire n_1379;
wire n_2734;
wire n_2196;
wire n_2170;
wire n_1076;
wire n_2823;
wire n_1091;
wire n_1408;
wire n_1761;
wire n_641;
wire n_730;
wire n_2036;
wire n_1325;
wire n_1595;
wire n_2161;
wire n_575;
wire n_795;
wire n_2404;
wire n_2083;
wire n_695;
wire n_656;
wire n_1606;
wire n_2503;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_2485;
wire n_1936;
wire n_1956;
wire n_1642;
wire n_2279;
wire n_2655;
wire n_2027;
wire n_2642;
wire n_1130;
wire n_720;
wire n_2500;
wire n_2366;
wire n_1918;
wire n_1526;
wire n_863;
wire n_2210;
wire n_805;
wire n_1604;
wire n_1275;
wire n_2513;
wire n_2525;
wire n_2695;
wire n_1764;
wire n_2892;
wire n_712;
wire n_2414;
wire n_2907;
wire n_1583;
wire n_2426;
wire n_2826;
wire n_1042;
wire n_1402;
wire n_2820;
wire n_2049;
wire n_2273;
wire n_2719;
wire n_1493;
wire n_657;
wire n_644;
wire n_1741;
wire n_2229;
wire n_1160;
wire n_1397;
wire n_1258;
wire n_1074;
wire n_2004;
wire n_1621;
wire n_2708;
wire n_2113;
wire n_566;
wire n_565;
wire n_2586;
wire n_1448;
wire n_2225;
wire n_1507;
wire n_1398;
wire n_2383;
wire n_1879;
wire n_597;
wire n_1996;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_2019;
wire n_651;
wire n_1340;
wire n_2274;
wire n_811;
wire n_1558;
wire n_807;
wire n_2166;
wire n_835;
wire n_666;
wire n_1433;
wire n_1704;
wire n_2256;
wire n_1254;
wire n_1026;
wire n_2026;
wire n_1969;
wire n_1234;
wire n_2109;
wire n_2044;
wire n_1138;
wire n_927;
wire n_1089;
wire n_2013;
wire n_1990;
wire n_2689;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_2614;
wire n_2511;
wire n_1681;
wire n_2010;
wire n_1018;
wire n_2242;
wire n_2247;
wire n_2752;
wire n_2894;
wire n_1693;
wire n_2599;
wire n_713;
wire n_2704;
wire n_904;
wire n_2839;
wire n_1588;
wire n_1622;
wire n_2237;
wire n_1180;
wire n_1827;
wire n_2524;
wire n_1271;
wire n_2802;
wire n_1542;
wire n_1251;
wire n_2728;
wire n_2268;

BUFx2_ASAP7_75t_L g555 ( 
.A(n_165),
.Y(n_555)
);

INVx2_ASAP7_75t_SL g556 ( 
.A(n_362),
.Y(n_556)
);

CKINVDCx5p33_ASAP7_75t_R g557 ( 
.A(n_139),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_35),
.Y(n_558)
);

CKINVDCx5p33_ASAP7_75t_R g559 ( 
.A(n_502),
.Y(n_559)
);

CKINVDCx5p33_ASAP7_75t_R g560 ( 
.A(n_457),
.Y(n_560)
);

CKINVDCx5p33_ASAP7_75t_R g561 ( 
.A(n_140),
.Y(n_561)
);

BUFx6f_ASAP7_75t_L g562 ( 
.A(n_499),
.Y(n_562)
);

CKINVDCx5p33_ASAP7_75t_R g563 ( 
.A(n_296),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_101),
.Y(n_564)
);

CKINVDCx20_ASAP7_75t_R g565 ( 
.A(n_416),
.Y(n_565)
);

CKINVDCx16_ASAP7_75t_R g566 ( 
.A(n_530),
.Y(n_566)
);

CKINVDCx14_ASAP7_75t_R g567 ( 
.A(n_473),
.Y(n_567)
);

CKINVDCx5p33_ASAP7_75t_R g568 ( 
.A(n_3),
.Y(n_568)
);

CKINVDCx20_ASAP7_75t_R g569 ( 
.A(n_94),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_15),
.Y(n_570)
);

CKINVDCx5p33_ASAP7_75t_R g571 ( 
.A(n_169),
.Y(n_571)
);

CKINVDCx14_ASAP7_75t_R g572 ( 
.A(n_167),
.Y(n_572)
);

CKINVDCx5p33_ASAP7_75t_R g573 ( 
.A(n_367),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_238),
.Y(n_574)
);

CKINVDCx5p33_ASAP7_75t_R g575 ( 
.A(n_507),
.Y(n_575)
);

INVxp67_ASAP7_75t_SL g576 ( 
.A(n_410),
.Y(n_576)
);

BUFx10_ASAP7_75t_L g577 ( 
.A(n_6),
.Y(n_577)
);

CKINVDCx5p33_ASAP7_75t_R g578 ( 
.A(n_488),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_348),
.Y(n_579)
);

INVx3_ASAP7_75t_L g580 ( 
.A(n_131),
.Y(n_580)
);

BUFx3_ASAP7_75t_L g581 ( 
.A(n_192),
.Y(n_581)
);

BUFx3_ASAP7_75t_L g582 ( 
.A(n_375),
.Y(n_582)
);

CKINVDCx5p33_ASAP7_75t_R g583 ( 
.A(n_532),
.Y(n_583)
);

INVx1_ASAP7_75t_SL g584 ( 
.A(n_521),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_86),
.Y(n_585)
);

INVx2_ASAP7_75t_SL g586 ( 
.A(n_445),
.Y(n_586)
);

BUFx6f_ASAP7_75t_L g587 ( 
.A(n_249),
.Y(n_587)
);

CKINVDCx20_ASAP7_75t_R g588 ( 
.A(n_366),
.Y(n_588)
);

CKINVDCx20_ASAP7_75t_R g589 ( 
.A(n_518),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_377),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_47),
.Y(n_591)
);

INVx1_ASAP7_75t_SL g592 ( 
.A(n_216),
.Y(n_592)
);

CKINVDCx5p33_ASAP7_75t_R g593 ( 
.A(n_420),
.Y(n_593)
);

INVx2_ASAP7_75t_SL g594 ( 
.A(n_520),
.Y(n_594)
);

CKINVDCx5p33_ASAP7_75t_R g595 ( 
.A(n_54),
.Y(n_595)
);

CKINVDCx5p33_ASAP7_75t_R g596 ( 
.A(n_461),
.Y(n_596)
);

CKINVDCx5p33_ASAP7_75t_R g597 ( 
.A(n_301),
.Y(n_597)
);

CKINVDCx5p33_ASAP7_75t_R g598 ( 
.A(n_6),
.Y(n_598)
);

BUFx10_ASAP7_75t_L g599 ( 
.A(n_97),
.Y(n_599)
);

CKINVDCx20_ASAP7_75t_R g600 ( 
.A(n_503),
.Y(n_600)
);

INVx2_ASAP7_75t_L g601 ( 
.A(n_220),
.Y(n_601)
);

INVx1_ASAP7_75t_SL g602 ( 
.A(n_242),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_536),
.Y(n_603)
);

CKINVDCx5p33_ASAP7_75t_R g604 ( 
.A(n_290),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_509),
.Y(n_605)
);

CKINVDCx5p33_ASAP7_75t_R g606 ( 
.A(n_270),
.Y(n_606)
);

CKINVDCx5p33_ASAP7_75t_R g607 ( 
.A(n_46),
.Y(n_607)
);

BUFx6f_ASAP7_75t_L g608 ( 
.A(n_41),
.Y(n_608)
);

CKINVDCx5p33_ASAP7_75t_R g609 ( 
.A(n_42),
.Y(n_609)
);

CKINVDCx5p33_ASAP7_75t_R g610 ( 
.A(n_204),
.Y(n_610)
);

INVx2_ASAP7_75t_L g611 ( 
.A(n_242),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_440),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_95),
.Y(n_613)
);

CKINVDCx5p33_ASAP7_75t_R g614 ( 
.A(n_205),
.Y(n_614)
);

CKINVDCx5p33_ASAP7_75t_R g615 ( 
.A(n_459),
.Y(n_615)
);

CKINVDCx5p33_ASAP7_75t_R g616 ( 
.A(n_98),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_446),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_495),
.Y(n_618)
);

INVx2_ASAP7_75t_L g619 ( 
.A(n_419),
.Y(n_619)
);

CKINVDCx5p33_ASAP7_75t_R g620 ( 
.A(n_251),
.Y(n_620)
);

BUFx2_ASAP7_75t_L g621 ( 
.A(n_513),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_396),
.Y(n_622)
);

CKINVDCx5p33_ASAP7_75t_R g623 ( 
.A(n_378),
.Y(n_623)
);

CKINVDCx20_ASAP7_75t_R g624 ( 
.A(n_87),
.Y(n_624)
);

CKINVDCx20_ASAP7_75t_R g625 ( 
.A(n_117),
.Y(n_625)
);

CKINVDCx5p33_ASAP7_75t_R g626 ( 
.A(n_281),
.Y(n_626)
);

CKINVDCx5p33_ASAP7_75t_R g627 ( 
.A(n_320),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_378),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_201),
.Y(n_629)
);

CKINVDCx5p33_ASAP7_75t_R g630 ( 
.A(n_535),
.Y(n_630)
);

INVx2_ASAP7_75t_SL g631 ( 
.A(n_67),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_122),
.Y(n_632)
);

CKINVDCx5p33_ASAP7_75t_R g633 ( 
.A(n_356),
.Y(n_633)
);

CKINVDCx5p33_ASAP7_75t_R g634 ( 
.A(n_280),
.Y(n_634)
);

CKINVDCx5p33_ASAP7_75t_R g635 ( 
.A(n_356),
.Y(n_635)
);

INVx2_ASAP7_75t_L g636 ( 
.A(n_374),
.Y(n_636)
);

CKINVDCx5p33_ASAP7_75t_R g637 ( 
.A(n_482),
.Y(n_637)
);

BUFx6f_ASAP7_75t_L g638 ( 
.A(n_471),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_205),
.Y(n_639)
);

BUFx6f_ASAP7_75t_L g640 ( 
.A(n_394),
.Y(n_640)
);

INVx2_ASAP7_75t_L g641 ( 
.A(n_62),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_292),
.Y(n_642)
);

CKINVDCx5p33_ASAP7_75t_R g643 ( 
.A(n_88),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_279),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_121),
.Y(n_645)
);

INVx2_ASAP7_75t_L g646 ( 
.A(n_316),
.Y(n_646)
);

INVx2_ASAP7_75t_L g647 ( 
.A(n_252),
.Y(n_647)
);

CKINVDCx5p33_ASAP7_75t_R g648 ( 
.A(n_59),
.Y(n_648)
);

INVx2_ASAP7_75t_L g649 ( 
.A(n_506),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_440),
.Y(n_650)
);

CKINVDCx5p33_ASAP7_75t_R g651 ( 
.A(n_78),
.Y(n_651)
);

CKINVDCx5p33_ASAP7_75t_R g652 ( 
.A(n_431),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_57),
.Y(n_653)
);

CKINVDCx5p33_ASAP7_75t_R g654 ( 
.A(n_436),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_435),
.Y(n_655)
);

CKINVDCx5p33_ASAP7_75t_R g656 ( 
.A(n_103),
.Y(n_656)
);

CKINVDCx5p33_ASAP7_75t_R g657 ( 
.A(n_539),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_179),
.Y(n_658)
);

BUFx6f_ASAP7_75t_L g659 ( 
.A(n_329),
.Y(n_659)
);

CKINVDCx5p33_ASAP7_75t_R g660 ( 
.A(n_443),
.Y(n_660)
);

CKINVDCx5p33_ASAP7_75t_R g661 ( 
.A(n_208),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_493),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_14),
.Y(n_663)
);

INVx1_ASAP7_75t_SL g664 ( 
.A(n_157),
.Y(n_664)
);

CKINVDCx16_ASAP7_75t_R g665 ( 
.A(n_463),
.Y(n_665)
);

INVx1_ASAP7_75t_SL g666 ( 
.A(n_491),
.Y(n_666)
);

BUFx2_ASAP7_75t_L g667 ( 
.A(n_288),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_28),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_24),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_268),
.Y(n_670)
);

CKINVDCx5p33_ASAP7_75t_R g671 ( 
.A(n_504),
.Y(n_671)
);

CKINVDCx5p33_ASAP7_75t_R g672 ( 
.A(n_2),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_544),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_34),
.Y(n_674)
);

CKINVDCx5p33_ASAP7_75t_R g675 ( 
.A(n_445),
.Y(n_675)
);

CKINVDCx5p33_ASAP7_75t_R g676 ( 
.A(n_540),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_227),
.Y(n_677)
);

CKINVDCx20_ASAP7_75t_R g678 ( 
.A(n_298),
.Y(n_678)
);

HB1xp67_ASAP7_75t_L g679 ( 
.A(n_232),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_220),
.Y(n_680)
);

CKINVDCx5p33_ASAP7_75t_R g681 ( 
.A(n_34),
.Y(n_681)
);

CKINVDCx5p33_ASAP7_75t_R g682 ( 
.A(n_457),
.Y(n_682)
);

CKINVDCx20_ASAP7_75t_R g683 ( 
.A(n_26),
.Y(n_683)
);

CKINVDCx5p33_ASAP7_75t_R g684 ( 
.A(n_12),
.Y(n_684)
);

CKINVDCx5p33_ASAP7_75t_R g685 ( 
.A(n_262),
.Y(n_685)
);

INVx1_ASAP7_75t_SL g686 ( 
.A(n_162),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_8),
.Y(n_687)
);

CKINVDCx5p33_ASAP7_75t_R g688 ( 
.A(n_204),
.Y(n_688)
);

CKINVDCx5p33_ASAP7_75t_R g689 ( 
.A(n_524),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_190),
.Y(n_690)
);

CKINVDCx5p33_ASAP7_75t_R g691 ( 
.A(n_144),
.Y(n_691)
);

CKINVDCx5p33_ASAP7_75t_R g692 ( 
.A(n_324),
.Y(n_692)
);

CKINVDCx5p33_ASAP7_75t_R g693 ( 
.A(n_60),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_324),
.Y(n_694)
);

BUFx2_ASAP7_75t_L g695 ( 
.A(n_545),
.Y(n_695)
);

CKINVDCx5p33_ASAP7_75t_R g696 ( 
.A(n_291),
.Y(n_696)
);

CKINVDCx5p33_ASAP7_75t_R g697 ( 
.A(n_143),
.Y(n_697)
);

CKINVDCx5p33_ASAP7_75t_R g698 ( 
.A(n_83),
.Y(n_698)
);

CKINVDCx5p33_ASAP7_75t_R g699 ( 
.A(n_30),
.Y(n_699)
);

CKINVDCx5p33_ASAP7_75t_R g700 ( 
.A(n_207),
.Y(n_700)
);

CKINVDCx20_ASAP7_75t_R g701 ( 
.A(n_58),
.Y(n_701)
);

CKINVDCx5p33_ASAP7_75t_R g702 ( 
.A(n_546),
.Y(n_702)
);

CKINVDCx5p33_ASAP7_75t_R g703 ( 
.A(n_398),
.Y(n_703)
);

CKINVDCx5p33_ASAP7_75t_R g704 ( 
.A(n_238),
.Y(n_704)
);

CKINVDCx5p33_ASAP7_75t_R g705 ( 
.A(n_52),
.Y(n_705)
);

BUFx2_ASAP7_75t_L g706 ( 
.A(n_483),
.Y(n_706)
);

CKINVDCx5p33_ASAP7_75t_R g707 ( 
.A(n_466),
.Y(n_707)
);

CKINVDCx5p33_ASAP7_75t_R g708 ( 
.A(n_253),
.Y(n_708)
);

CKINVDCx5p33_ASAP7_75t_R g709 ( 
.A(n_289),
.Y(n_709)
);

CKINVDCx5p33_ASAP7_75t_R g710 ( 
.A(n_349),
.Y(n_710)
);

CKINVDCx20_ASAP7_75t_R g711 ( 
.A(n_12),
.Y(n_711)
);

INVx2_ASAP7_75t_L g712 ( 
.A(n_343),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_33),
.Y(n_713)
);

CKINVDCx5p33_ASAP7_75t_R g714 ( 
.A(n_271),
.Y(n_714)
);

CKINVDCx5p33_ASAP7_75t_R g715 ( 
.A(n_494),
.Y(n_715)
);

CKINVDCx5p33_ASAP7_75t_R g716 ( 
.A(n_10),
.Y(n_716)
);

CKINVDCx5p33_ASAP7_75t_R g717 ( 
.A(n_487),
.Y(n_717)
);

CKINVDCx5p33_ASAP7_75t_R g718 ( 
.A(n_376),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_468),
.Y(n_719)
);

CKINVDCx5p33_ASAP7_75t_R g720 ( 
.A(n_538),
.Y(n_720)
);

INVx2_ASAP7_75t_L g721 ( 
.A(n_69),
.Y(n_721)
);

BUFx10_ASAP7_75t_L g722 ( 
.A(n_225),
.Y(n_722)
);

CKINVDCx5p33_ASAP7_75t_R g723 ( 
.A(n_441),
.Y(n_723)
);

BUFx3_ASAP7_75t_L g724 ( 
.A(n_376),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_179),
.Y(n_725)
);

CKINVDCx5p33_ASAP7_75t_R g726 ( 
.A(n_519),
.Y(n_726)
);

CKINVDCx5p33_ASAP7_75t_R g727 ( 
.A(n_379),
.Y(n_727)
);

CKINVDCx5p33_ASAP7_75t_R g728 ( 
.A(n_129),
.Y(n_728)
);

CKINVDCx5p33_ASAP7_75t_R g729 ( 
.A(n_515),
.Y(n_729)
);

CKINVDCx20_ASAP7_75t_R g730 ( 
.A(n_533),
.Y(n_730)
);

CKINVDCx5p33_ASAP7_75t_R g731 ( 
.A(n_268),
.Y(n_731)
);

INVx1_ASAP7_75t_SL g732 ( 
.A(n_458),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_123),
.Y(n_733)
);

CKINVDCx5p33_ASAP7_75t_R g734 ( 
.A(n_121),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_492),
.Y(n_735)
);

CKINVDCx5p33_ASAP7_75t_R g736 ( 
.A(n_322),
.Y(n_736)
);

CKINVDCx20_ASAP7_75t_R g737 ( 
.A(n_212),
.Y(n_737)
);

CKINVDCx5p33_ASAP7_75t_R g738 ( 
.A(n_460),
.Y(n_738)
);

CKINVDCx5p33_ASAP7_75t_R g739 ( 
.A(n_217),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_104),
.Y(n_740)
);

CKINVDCx5p33_ASAP7_75t_R g741 ( 
.A(n_403),
.Y(n_741)
);

INVx2_ASAP7_75t_L g742 ( 
.A(n_180),
.Y(n_742)
);

CKINVDCx5p33_ASAP7_75t_R g743 ( 
.A(n_103),
.Y(n_743)
);

CKINVDCx5p33_ASAP7_75t_R g744 ( 
.A(n_270),
.Y(n_744)
);

BUFx8_ASAP7_75t_SL g745 ( 
.A(n_194),
.Y(n_745)
);

INVx1_ASAP7_75t_SL g746 ( 
.A(n_278),
.Y(n_746)
);

CKINVDCx5p33_ASAP7_75t_R g747 ( 
.A(n_516),
.Y(n_747)
);

CKINVDCx20_ASAP7_75t_R g748 ( 
.A(n_534),
.Y(n_748)
);

INVx2_ASAP7_75t_SL g749 ( 
.A(n_415),
.Y(n_749)
);

CKINVDCx5p33_ASAP7_75t_R g750 ( 
.A(n_246),
.Y(n_750)
);

CKINVDCx5p33_ASAP7_75t_R g751 ( 
.A(n_165),
.Y(n_751)
);

BUFx6f_ASAP7_75t_L g752 ( 
.A(n_40),
.Y(n_752)
);

CKINVDCx5p33_ASAP7_75t_R g753 ( 
.A(n_214),
.Y(n_753)
);

INVx2_ASAP7_75t_L g754 ( 
.A(n_132),
.Y(n_754)
);

CKINVDCx5p33_ASAP7_75t_R g755 ( 
.A(n_226),
.Y(n_755)
);

CKINVDCx5p33_ASAP7_75t_R g756 ( 
.A(n_455),
.Y(n_756)
);

CKINVDCx5p33_ASAP7_75t_R g757 ( 
.A(n_74),
.Y(n_757)
);

CKINVDCx14_ASAP7_75t_R g758 ( 
.A(n_1),
.Y(n_758)
);

CKINVDCx5p33_ASAP7_75t_R g759 ( 
.A(n_329),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_552),
.Y(n_760)
);

INVx2_ASAP7_75t_L g761 ( 
.A(n_527),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_309),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_162),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_113),
.Y(n_764)
);

CKINVDCx5p33_ASAP7_75t_R g765 ( 
.A(n_429),
.Y(n_765)
);

CKINVDCx20_ASAP7_75t_R g766 ( 
.A(n_59),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_377),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_349),
.Y(n_768)
);

CKINVDCx5p33_ASAP7_75t_R g769 ( 
.A(n_517),
.Y(n_769)
);

CKINVDCx5p33_ASAP7_75t_R g770 ( 
.A(n_304),
.Y(n_770)
);

BUFx8_ASAP7_75t_SL g771 ( 
.A(n_202),
.Y(n_771)
);

CKINVDCx20_ASAP7_75t_R g772 ( 
.A(n_364),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_479),
.Y(n_773)
);

INVx2_ASAP7_75t_SL g774 ( 
.A(n_514),
.Y(n_774)
);

CKINVDCx5p33_ASAP7_75t_R g775 ( 
.A(n_62),
.Y(n_775)
);

CKINVDCx16_ASAP7_75t_R g776 ( 
.A(n_485),
.Y(n_776)
);

CKINVDCx5p33_ASAP7_75t_R g777 ( 
.A(n_448),
.Y(n_777)
);

BUFx2_ASAP7_75t_L g778 ( 
.A(n_525),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_476),
.Y(n_779)
);

INVx2_ASAP7_75t_L g780 ( 
.A(n_32),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_421),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_266),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_373),
.Y(n_783)
);

CKINVDCx14_ASAP7_75t_R g784 ( 
.A(n_455),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_323),
.Y(n_785)
);

CKINVDCx5p33_ASAP7_75t_R g786 ( 
.A(n_144),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_365),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_497),
.Y(n_788)
);

CKINVDCx5p33_ASAP7_75t_R g789 ( 
.A(n_232),
.Y(n_789)
);

CKINVDCx5p33_ASAP7_75t_R g790 ( 
.A(n_438),
.Y(n_790)
);

CKINVDCx5p33_ASAP7_75t_R g791 ( 
.A(n_194),
.Y(n_791)
);

CKINVDCx5p33_ASAP7_75t_R g792 ( 
.A(n_382),
.Y(n_792)
);

CKINVDCx5p33_ASAP7_75t_R g793 ( 
.A(n_541),
.Y(n_793)
);

CKINVDCx5p33_ASAP7_75t_R g794 ( 
.A(n_490),
.Y(n_794)
);

CKINVDCx5p33_ASAP7_75t_R g795 ( 
.A(n_306),
.Y(n_795)
);

CKINVDCx5p33_ASAP7_75t_R g796 ( 
.A(n_190),
.Y(n_796)
);

CKINVDCx5p33_ASAP7_75t_R g797 ( 
.A(n_78),
.Y(n_797)
);

CKINVDCx5p33_ASAP7_75t_R g798 ( 
.A(n_30),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_364),
.Y(n_799)
);

CKINVDCx5p33_ASAP7_75t_R g800 ( 
.A(n_392),
.Y(n_800)
);

CKINVDCx20_ASAP7_75t_R g801 ( 
.A(n_447),
.Y(n_801)
);

CKINVDCx5p33_ASAP7_75t_R g802 ( 
.A(n_542),
.Y(n_802)
);

CKINVDCx5p33_ASAP7_75t_R g803 ( 
.A(n_478),
.Y(n_803)
);

CKINVDCx5p33_ASAP7_75t_R g804 ( 
.A(n_522),
.Y(n_804)
);

CKINVDCx5p33_ASAP7_75t_R g805 ( 
.A(n_222),
.Y(n_805)
);

BUFx6f_ASAP7_75t_L g806 ( 
.A(n_66),
.Y(n_806)
);

CKINVDCx5p33_ASAP7_75t_R g807 ( 
.A(n_547),
.Y(n_807)
);

CKINVDCx5p33_ASAP7_75t_R g808 ( 
.A(n_452),
.Y(n_808)
);

CKINVDCx5p33_ASAP7_75t_R g809 ( 
.A(n_44),
.Y(n_809)
);

CKINVDCx5p33_ASAP7_75t_R g810 ( 
.A(n_336),
.Y(n_810)
);

CKINVDCx5p33_ASAP7_75t_R g811 ( 
.A(n_456),
.Y(n_811)
);

CKINVDCx5p33_ASAP7_75t_R g812 ( 
.A(n_300),
.Y(n_812)
);

CKINVDCx5p33_ASAP7_75t_R g813 ( 
.A(n_323),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_439),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_60),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_353),
.Y(n_816)
);

BUFx5_ASAP7_75t_L g817 ( 
.A(n_551),
.Y(n_817)
);

CKINVDCx5p33_ASAP7_75t_R g818 ( 
.A(n_374),
.Y(n_818)
);

CKINVDCx5p33_ASAP7_75t_R g819 ( 
.A(n_549),
.Y(n_819)
);

CKINVDCx5p33_ASAP7_75t_R g820 ( 
.A(n_212),
.Y(n_820)
);

CKINVDCx5p33_ASAP7_75t_R g821 ( 
.A(n_489),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_470),
.Y(n_822)
);

INVx2_ASAP7_75t_L g823 ( 
.A(n_371),
.Y(n_823)
);

CKINVDCx5p33_ASAP7_75t_R g824 ( 
.A(n_198),
.Y(n_824)
);

CKINVDCx20_ASAP7_75t_R g825 ( 
.A(n_390),
.Y(n_825)
);

BUFx3_ASAP7_75t_L g826 ( 
.A(n_273),
.Y(n_826)
);

CKINVDCx5p33_ASAP7_75t_R g827 ( 
.A(n_237),
.Y(n_827)
);

CKINVDCx5p33_ASAP7_75t_R g828 ( 
.A(n_481),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_79),
.Y(n_829)
);

CKINVDCx20_ASAP7_75t_R g830 ( 
.A(n_406),
.Y(n_830)
);

INVxp67_ASAP7_75t_L g831 ( 
.A(n_156),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_160),
.Y(n_832)
);

BUFx3_ASAP7_75t_L g833 ( 
.A(n_496),
.Y(n_833)
);

CKINVDCx5p33_ASAP7_75t_R g834 ( 
.A(n_304),
.Y(n_834)
);

CKINVDCx5p33_ASAP7_75t_R g835 ( 
.A(n_222),
.Y(n_835)
);

CKINVDCx5p33_ASAP7_75t_R g836 ( 
.A(n_55),
.Y(n_836)
);

BUFx10_ASAP7_75t_L g837 ( 
.A(n_66),
.Y(n_837)
);

CKINVDCx5p33_ASAP7_75t_R g838 ( 
.A(n_27),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_224),
.Y(n_839)
);

BUFx10_ASAP7_75t_L g840 ( 
.A(n_82),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_398),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_47),
.Y(n_842)
);

CKINVDCx5p33_ASAP7_75t_R g843 ( 
.A(n_432),
.Y(n_843)
);

CKINVDCx5p33_ASAP7_75t_R g844 ( 
.A(n_472),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_256),
.Y(n_845)
);

CKINVDCx5p33_ASAP7_75t_R g846 ( 
.A(n_500),
.Y(n_846)
);

INVx1_ASAP7_75t_SL g847 ( 
.A(n_435),
.Y(n_847)
);

CKINVDCx16_ASAP7_75t_R g848 ( 
.A(n_462),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_511),
.Y(n_849)
);

CKINVDCx5p33_ASAP7_75t_R g850 ( 
.A(n_273),
.Y(n_850)
);

CKINVDCx5p33_ASAP7_75t_R g851 ( 
.A(n_136),
.Y(n_851)
);

CKINVDCx5p33_ASAP7_75t_R g852 ( 
.A(n_118),
.Y(n_852)
);

BUFx2_ASAP7_75t_L g853 ( 
.A(n_166),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_404),
.Y(n_854)
);

CKINVDCx5p33_ASAP7_75t_R g855 ( 
.A(n_197),
.Y(n_855)
);

CKINVDCx16_ASAP7_75t_R g856 ( 
.A(n_459),
.Y(n_856)
);

CKINVDCx5p33_ASAP7_75t_R g857 ( 
.A(n_119),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_486),
.Y(n_858)
);

INVx2_ASAP7_75t_L g859 ( 
.A(n_177),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_152),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_208),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_429),
.Y(n_862)
);

CKINVDCx5p33_ASAP7_75t_R g863 ( 
.A(n_22),
.Y(n_863)
);

CKINVDCx5p33_ASAP7_75t_R g864 ( 
.A(n_24),
.Y(n_864)
);

CKINVDCx20_ASAP7_75t_R g865 ( 
.A(n_537),
.Y(n_865)
);

CKINVDCx5p33_ASAP7_75t_R g866 ( 
.A(n_4),
.Y(n_866)
);

CKINVDCx20_ASAP7_75t_R g867 ( 
.A(n_249),
.Y(n_867)
);

CKINVDCx5p33_ASAP7_75t_R g868 ( 
.A(n_174),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_86),
.Y(n_869)
);

CKINVDCx5p33_ASAP7_75t_R g870 ( 
.A(n_51),
.Y(n_870)
);

BUFx3_ASAP7_75t_L g871 ( 
.A(n_465),
.Y(n_871)
);

BUFx2_ASAP7_75t_L g872 ( 
.A(n_498),
.Y(n_872)
);

BUFx2_ASAP7_75t_L g873 ( 
.A(n_439),
.Y(n_873)
);

BUFx10_ASAP7_75t_L g874 ( 
.A(n_207),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_210),
.Y(n_875)
);

CKINVDCx5p33_ASAP7_75t_R g876 ( 
.A(n_18),
.Y(n_876)
);

CKINVDCx5p33_ASAP7_75t_R g877 ( 
.A(n_88),
.Y(n_877)
);

CKINVDCx5p33_ASAP7_75t_R g878 ( 
.A(n_299),
.Y(n_878)
);

CKINVDCx5p33_ASAP7_75t_R g879 ( 
.A(n_291),
.Y(n_879)
);

CKINVDCx20_ASAP7_75t_R g880 ( 
.A(n_173),
.Y(n_880)
);

CKINVDCx5p33_ASAP7_75t_R g881 ( 
.A(n_451),
.Y(n_881)
);

CKINVDCx5p33_ASAP7_75t_R g882 ( 
.A(n_76),
.Y(n_882)
);

CKINVDCx5p33_ASAP7_75t_R g883 ( 
.A(n_111),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_523),
.Y(n_884)
);

CKINVDCx20_ASAP7_75t_R g885 ( 
.A(n_108),
.Y(n_885)
);

CKINVDCx5p33_ASAP7_75t_R g886 ( 
.A(n_370),
.Y(n_886)
);

CKINVDCx5p33_ASAP7_75t_R g887 ( 
.A(n_252),
.Y(n_887)
);

INVx2_ASAP7_75t_SL g888 ( 
.A(n_444),
.Y(n_888)
);

CKINVDCx5p33_ASAP7_75t_R g889 ( 
.A(n_372),
.Y(n_889)
);

CKINVDCx20_ASAP7_75t_R g890 ( 
.A(n_285),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_186),
.Y(n_891)
);

CKINVDCx5p33_ASAP7_75t_R g892 ( 
.A(n_308),
.Y(n_892)
);

INVx2_ASAP7_75t_L g893 ( 
.A(n_428),
.Y(n_893)
);

BUFx6f_ASAP7_75t_L g894 ( 
.A(n_184),
.Y(n_894)
);

CKINVDCx5p33_ASAP7_75t_R g895 ( 
.A(n_147),
.Y(n_895)
);

INVx2_ASAP7_75t_L g896 ( 
.A(n_477),
.Y(n_896)
);

CKINVDCx5p33_ASAP7_75t_R g897 ( 
.A(n_255),
.Y(n_897)
);

CKINVDCx5p33_ASAP7_75t_R g898 ( 
.A(n_119),
.Y(n_898)
);

CKINVDCx5p33_ASAP7_75t_R g899 ( 
.A(n_350),
.Y(n_899)
);

CKINVDCx20_ASAP7_75t_R g900 ( 
.A(n_0),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_170),
.Y(n_901)
);

CKINVDCx5p33_ASAP7_75t_R g902 ( 
.A(n_221),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_122),
.Y(n_903)
);

INVx1_ASAP7_75t_SL g904 ( 
.A(n_288),
.Y(n_904)
);

INVx1_ASAP7_75t_SL g905 ( 
.A(n_275),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_508),
.Y(n_906)
);

CKINVDCx5p33_ASAP7_75t_R g907 ( 
.A(n_458),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_275),
.Y(n_908)
);

BUFx10_ASAP7_75t_L g909 ( 
.A(n_31),
.Y(n_909)
);

CKINVDCx5p33_ASAP7_75t_R g910 ( 
.A(n_345),
.Y(n_910)
);

CKINVDCx5p33_ASAP7_75t_R g911 ( 
.A(n_361),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_315),
.Y(n_912)
);

INVx1_ASAP7_75t_SL g913 ( 
.A(n_20),
.Y(n_913)
);

CKINVDCx5p33_ASAP7_75t_R g914 ( 
.A(n_187),
.Y(n_914)
);

INVx1_ASAP7_75t_SL g915 ( 
.A(n_131),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_480),
.Y(n_916)
);

CKINVDCx5p33_ASAP7_75t_R g917 ( 
.A(n_436),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_54),
.Y(n_918)
);

CKINVDCx5p33_ASAP7_75t_R g919 ( 
.A(n_449),
.Y(n_919)
);

BUFx10_ASAP7_75t_L g920 ( 
.A(n_105),
.Y(n_920)
);

INVx1_ASAP7_75t_SL g921 ( 
.A(n_444),
.Y(n_921)
);

CKINVDCx5p33_ASAP7_75t_R g922 ( 
.A(n_529),
.Y(n_922)
);

INVx2_ASAP7_75t_L g923 ( 
.A(n_199),
.Y(n_923)
);

CKINVDCx5p33_ASAP7_75t_R g924 ( 
.A(n_269),
.Y(n_924)
);

CKINVDCx5p33_ASAP7_75t_R g925 ( 
.A(n_510),
.Y(n_925)
);

CKINVDCx5p33_ASAP7_75t_R g926 ( 
.A(n_348),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_528),
.Y(n_927)
);

CKINVDCx5p33_ASAP7_75t_R g928 ( 
.A(n_161),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_453),
.Y(n_929)
);

CKINVDCx5p33_ASAP7_75t_R g930 ( 
.A(n_372),
.Y(n_930)
);

CKINVDCx5p33_ASAP7_75t_R g931 ( 
.A(n_139),
.Y(n_931)
);

INVx2_ASAP7_75t_L g932 ( 
.A(n_89),
.Y(n_932)
);

CKINVDCx5p33_ASAP7_75t_R g933 ( 
.A(n_434),
.Y(n_933)
);

CKINVDCx5p33_ASAP7_75t_R g934 ( 
.A(n_553),
.Y(n_934)
);

CKINVDCx5p33_ASAP7_75t_R g935 ( 
.A(n_321),
.Y(n_935)
);

CKINVDCx5p33_ASAP7_75t_R g936 ( 
.A(n_206),
.Y(n_936)
);

CKINVDCx5p33_ASAP7_75t_R g937 ( 
.A(n_413),
.Y(n_937)
);

CKINVDCx5p33_ASAP7_75t_R g938 ( 
.A(n_302),
.Y(n_938)
);

INVx2_ASAP7_75t_SL g939 ( 
.A(n_437),
.Y(n_939)
);

CKINVDCx5p33_ASAP7_75t_R g940 ( 
.A(n_200),
.Y(n_940)
);

CKINVDCx5p33_ASAP7_75t_R g941 ( 
.A(n_526),
.Y(n_941)
);

INVx1_ASAP7_75t_L g942 ( 
.A(n_290),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_11),
.Y(n_943)
);

CKINVDCx5p33_ASAP7_75t_R g944 ( 
.A(n_189),
.Y(n_944)
);

INVx1_ASAP7_75t_L g945 ( 
.A(n_450),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_343),
.Y(n_946)
);

CKINVDCx5p33_ASAP7_75t_R g947 ( 
.A(n_199),
.Y(n_947)
);

INVx1_ASAP7_75t_L g948 ( 
.A(n_237),
.Y(n_948)
);

CKINVDCx5p33_ASAP7_75t_R g949 ( 
.A(n_505),
.Y(n_949)
);

CKINVDCx5p33_ASAP7_75t_R g950 ( 
.A(n_27),
.Y(n_950)
);

CKINVDCx5p33_ASAP7_75t_R g951 ( 
.A(n_475),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_464),
.Y(n_952)
);

CKINVDCx5p33_ASAP7_75t_R g953 ( 
.A(n_39),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_369),
.Y(n_954)
);

CKINVDCx20_ASAP7_75t_R g955 ( 
.A(n_167),
.Y(n_955)
);

INVx1_ASAP7_75t_L g956 ( 
.A(n_168),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_286),
.Y(n_957)
);

CKINVDCx5p33_ASAP7_75t_R g958 ( 
.A(n_454),
.Y(n_958)
);

INVx2_ASAP7_75t_SL g959 ( 
.A(n_422),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_117),
.Y(n_960)
);

CKINVDCx5p33_ASAP7_75t_R g961 ( 
.A(n_172),
.Y(n_961)
);

BUFx10_ASAP7_75t_L g962 ( 
.A(n_550),
.Y(n_962)
);

CKINVDCx5p33_ASAP7_75t_R g963 ( 
.A(n_8),
.Y(n_963)
);

INVx1_ASAP7_75t_L g964 ( 
.A(n_548),
.Y(n_964)
);

CKINVDCx5p33_ASAP7_75t_R g965 ( 
.A(n_484),
.Y(n_965)
);

CKINVDCx20_ASAP7_75t_R g966 ( 
.A(n_428),
.Y(n_966)
);

HB1xp67_ASAP7_75t_L g967 ( 
.A(n_46),
.Y(n_967)
);

INVx2_ASAP7_75t_L g968 ( 
.A(n_61),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_276),
.Y(n_969)
);

CKINVDCx5p33_ASAP7_75t_R g970 ( 
.A(n_0),
.Y(n_970)
);

CKINVDCx5p33_ASAP7_75t_R g971 ( 
.A(n_241),
.Y(n_971)
);

CKINVDCx5p33_ASAP7_75t_R g972 ( 
.A(n_20),
.Y(n_972)
);

CKINVDCx5p33_ASAP7_75t_R g973 ( 
.A(n_330),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_501),
.Y(n_974)
);

CKINVDCx5p33_ASAP7_75t_R g975 ( 
.A(n_554),
.Y(n_975)
);

CKINVDCx5p33_ASAP7_75t_R g976 ( 
.A(n_474),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_410),
.Y(n_977)
);

CKINVDCx20_ASAP7_75t_R g978 ( 
.A(n_68),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_371),
.Y(n_979)
);

CKINVDCx5p33_ASAP7_75t_R g980 ( 
.A(n_512),
.Y(n_980)
);

CKINVDCx5p33_ASAP7_75t_R g981 ( 
.A(n_140),
.Y(n_981)
);

INVx1_ASAP7_75t_SL g982 ( 
.A(n_543),
.Y(n_982)
);

CKINVDCx5p33_ASAP7_75t_R g983 ( 
.A(n_442),
.Y(n_983)
);

INVx1_ASAP7_75t_L g984 ( 
.A(n_203),
.Y(n_984)
);

INVx2_ASAP7_75t_L g985 ( 
.A(n_281),
.Y(n_985)
);

BUFx2_ASAP7_75t_L g986 ( 
.A(n_299),
.Y(n_986)
);

CKINVDCx5p33_ASAP7_75t_R g987 ( 
.A(n_14),
.Y(n_987)
);

CKINVDCx20_ASAP7_75t_R g988 ( 
.A(n_104),
.Y(n_988)
);

BUFx10_ASAP7_75t_L g989 ( 
.A(n_265),
.Y(n_989)
);

CKINVDCx5p33_ASAP7_75t_R g990 ( 
.A(n_80),
.Y(n_990)
);

INVx1_ASAP7_75t_L g991 ( 
.A(n_201),
.Y(n_991)
);

INVx1_ASAP7_75t_L g992 ( 
.A(n_193),
.Y(n_992)
);

CKINVDCx5p33_ASAP7_75t_R g993 ( 
.A(n_256),
.Y(n_993)
);

INVx1_ASAP7_75t_L g994 ( 
.A(n_22),
.Y(n_994)
);

CKINVDCx20_ASAP7_75t_R g995 ( 
.A(n_389),
.Y(n_995)
);

INVx2_ASAP7_75t_L g996 ( 
.A(n_381),
.Y(n_996)
);

INVx2_ASAP7_75t_L g997 ( 
.A(n_109),
.Y(n_997)
);

BUFx3_ASAP7_75t_L g998 ( 
.A(n_531),
.Y(n_998)
);

CKINVDCx5p33_ASAP7_75t_R g999 ( 
.A(n_97),
.Y(n_999)
);

CKINVDCx5p33_ASAP7_75t_R g1000 ( 
.A(n_413),
.Y(n_1000)
);

CKINVDCx5p33_ASAP7_75t_R g1001 ( 
.A(n_219),
.Y(n_1001)
);

INVx2_ASAP7_75t_L g1002 ( 
.A(n_218),
.Y(n_1002)
);

BUFx3_ASAP7_75t_L g1003 ( 
.A(n_312),
.Y(n_1003)
);

CKINVDCx5p33_ASAP7_75t_R g1004 ( 
.A(n_278),
.Y(n_1004)
);

INVx2_ASAP7_75t_L g1005 ( 
.A(n_580),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_603),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_603),
.Y(n_1007)
);

BUFx6f_ASAP7_75t_L g1008 ( 
.A(n_562),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_605),
.Y(n_1009)
);

HB1xp67_ASAP7_75t_L g1010 ( 
.A(n_555),
.Y(n_1010)
);

INVx1_ASAP7_75t_L g1011 ( 
.A(n_605),
.Y(n_1011)
);

INVx1_ASAP7_75t_L g1012 ( 
.A(n_618),
.Y(n_1012)
);

INVx1_ASAP7_75t_L g1013 ( 
.A(n_618),
.Y(n_1013)
);

INVx1_ASAP7_75t_L g1014 ( 
.A(n_662),
.Y(n_1014)
);

BUFx2_ASAP7_75t_SL g1015 ( 
.A(n_589),
.Y(n_1015)
);

INVx1_ASAP7_75t_L g1016 ( 
.A(n_662),
.Y(n_1016)
);

INVx1_ASAP7_75t_L g1017 ( 
.A(n_673),
.Y(n_1017)
);

INVx1_ASAP7_75t_L g1018 ( 
.A(n_673),
.Y(n_1018)
);

INVx1_ASAP7_75t_L g1019 ( 
.A(n_719),
.Y(n_1019)
);

INVx1_ASAP7_75t_L g1020 ( 
.A(n_719),
.Y(n_1020)
);

INVx1_ASAP7_75t_L g1021 ( 
.A(n_735),
.Y(n_1021)
);

INVx1_ASAP7_75t_L g1022 ( 
.A(n_735),
.Y(n_1022)
);

HB1xp67_ASAP7_75t_L g1023 ( 
.A(n_555),
.Y(n_1023)
);

HB1xp67_ASAP7_75t_L g1024 ( 
.A(n_667),
.Y(n_1024)
);

INVxp33_ASAP7_75t_L g1025 ( 
.A(n_679),
.Y(n_1025)
);

CKINVDCx5p33_ASAP7_75t_R g1026 ( 
.A(n_745),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_760),
.Y(n_1027)
);

CKINVDCx5p33_ASAP7_75t_R g1028 ( 
.A(n_771),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_760),
.Y(n_1029)
);

CKINVDCx5p33_ASAP7_75t_R g1030 ( 
.A(n_572),
.Y(n_1030)
);

CKINVDCx5p33_ASAP7_75t_R g1031 ( 
.A(n_758),
.Y(n_1031)
);

INVx1_ASAP7_75t_L g1032 ( 
.A(n_773),
.Y(n_1032)
);

INVx1_ASAP7_75t_L g1033 ( 
.A(n_773),
.Y(n_1033)
);

CKINVDCx20_ASAP7_75t_R g1034 ( 
.A(n_565),
.Y(n_1034)
);

INVx1_ASAP7_75t_L g1035 ( 
.A(n_779),
.Y(n_1035)
);

INVx1_ASAP7_75t_L g1036 ( 
.A(n_779),
.Y(n_1036)
);

INVx1_ASAP7_75t_L g1037 ( 
.A(n_788),
.Y(n_1037)
);

CKINVDCx20_ASAP7_75t_R g1038 ( 
.A(n_569),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_788),
.Y(n_1039)
);

CKINVDCx5p33_ASAP7_75t_R g1040 ( 
.A(n_784),
.Y(n_1040)
);

INVx1_ASAP7_75t_L g1041 ( 
.A(n_822),
.Y(n_1041)
);

INVx2_ASAP7_75t_SL g1042 ( 
.A(n_581),
.Y(n_1042)
);

INVx1_ASAP7_75t_L g1043 ( 
.A(n_822),
.Y(n_1043)
);

CKINVDCx20_ASAP7_75t_R g1044 ( 
.A(n_588),
.Y(n_1044)
);

CKINVDCx16_ASAP7_75t_R g1045 ( 
.A(n_665),
.Y(n_1045)
);

INVx1_ASAP7_75t_L g1046 ( 
.A(n_849),
.Y(n_1046)
);

INVx1_ASAP7_75t_L g1047 ( 
.A(n_849),
.Y(n_1047)
);

CKINVDCx5p33_ASAP7_75t_R g1048 ( 
.A(n_848),
.Y(n_1048)
);

INVx2_ASAP7_75t_L g1049 ( 
.A(n_580),
.Y(n_1049)
);

INVx1_ASAP7_75t_L g1050 ( 
.A(n_858),
.Y(n_1050)
);

INVx1_ASAP7_75t_L g1051 ( 
.A(n_858),
.Y(n_1051)
);

CKINVDCx5p33_ASAP7_75t_R g1052 ( 
.A(n_856),
.Y(n_1052)
);

INVx1_ASAP7_75t_L g1053 ( 
.A(n_884),
.Y(n_1053)
);

CKINVDCx16_ASAP7_75t_R g1054 ( 
.A(n_566),
.Y(n_1054)
);

BUFx6f_ASAP7_75t_L g1055 ( 
.A(n_562),
.Y(n_1055)
);

CKINVDCx16_ASAP7_75t_R g1056 ( 
.A(n_776),
.Y(n_1056)
);

CKINVDCx20_ASAP7_75t_R g1057 ( 
.A(n_624),
.Y(n_1057)
);

INVx1_ASAP7_75t_L g1058 ( 
.A(n_884),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_906),
.Y(n_1059)
);

CKINVDCx5p33_ASAP7_75t_R g1060 ( 
.A(n_557),
.Y(n_1060)
);

CKINVDCx5p33_ASAP7_75t_R g1061 ( 
.A(n_560),
.Y(n_1061)
);

INVx1_ASAP7_75t_L g1062 ( 
.A(n_906),
.Y(n_1062)
);

BUFx3_ASAP7_75t_L g1063 ( 
.A(n_833),
.Y(n_1063)
);

INVx1_ASAP7_75t_L g1064 ( 
.A(n_916),
.Y(n_1064)
);

INVx1_ASAP7_75t_L g1065 ( 
.A(n_916),
.Y(n_1065)
);

CKINVDCx20_ASAP7_75t_R g1066 ( 
.A(n_625),
.Y(n_1066)
);

INVx1_ASAP7_75t_L g1067 ( 
.A(n_927),
.Y(n_1067)
);

INVx1_ASAP7_75t_L g1068 ( 
.A(n_927),
.Y(n_1068)
);

INVxp67_ASAP7_75t_L g1069 ( 
.A(n_667),
.Y(n_1069)
);

INVx1_ASAP7_75t_L g1070 ( 
.A(n_964),
.Y(n_1070)
);

INVx1_ASAP7_75t_L g1071 ( 
.A(n_964),
.Y(n_1071)
);

INVx1_ASAP7_75t_L g1072 ( 
.A(n_974),
.Y(n_1072)
);

CKINVDCx20_ASAP7_75t_R g1073 ( 
.A(n_678),
.Y(n_1073)
);

CKINVDCx5p33_ASAP7_75t_R g1074 ( 
.A(n_561),
.Y(n_1074)
);

INVx1_ASAP7_75t_L g1075 ( 
.A(n_974),
.Y(n_1075)
);

INVx1_ASAP7_75t_L g1076 ( 
.A(n_580),
.Y(n_1076)
);

CKINVDCx5p33_ASAP7_75t_R g1077 ( 
.A(n_563),
.Y(n_1077)
);

INVx2_ASAP7_75t_L g1078 ( 
.A(n_587),
.Y(n_1078)
);

INVx1_ASAP7_75t_L g1079 ( 
.A(n_581),
.Y(n_1079)
);

INVx1_ASAP7_75t_L g1080 ( 
.A(n_582),
.Y(n_1080)
);

INVx1_ASAP7_75t_L g1081 ( 
.A(n_582),
.Y(n_1081)
);

CKINVDCx20_ASAP7_75t_R g1082 ( 
.A(n_683),
.Y(n_1082)
);

INVx1_ASAP7_75t_L g1083 ( 
.A(n_724),
.Y(n_1083)
);

CKINVDCx5p33_ASAP7_75t_R g1084 ( 
.A(n_568),
.Y(n_1084)
);

INVx1_ASAP7_75t_SL g1085 ( 
.A(n_853),
.Y(n_1085)
);

INVx1_ASAP7_75t_L g1086 ( 
.A(n_724),
.Y(n_1086)
);

INVx1_ASAP7_75t_L g1087 ( 
.A(n_826),
.Y(n_1087)
);

INVxp67_ASAP7_75t_SL g1088 ( 
.A(n_621),
.Y(n_1088)
);

CKINVDCx5p33_ASAP7_75t_R g1089 ( 
.A(n_571),
.Y(n_1089)
);

INVx1_ASAP7_75t_L g1090 ( 
.A(n_826),
.Y(n_1090)
);

INVx1_ASAP7_75t_L g1091 ( 
.A(n_871),
.Y(n_1091)
);

CKINVDCx16_ASAP7_75t_R g1092 ( 
.A(n_776),
.Y(n_1092)
);

CKINVDCx5p33_ASAP7_75t_R g1093 ( 
.A(n_1015),
.Y(n_1093)
);

INVx4_ASAP7_75t_L g1094 ( 
.A(n_1008),
.Y(n_1094)
);

INVx3_ASAP7_75t_L g1095 ( 
.A(n_1008),
.Y(n_1095)
);

CKINVDCx20_ASAP7_75t_R g1096 ( 
.A(n_1034),
.Y(n_1096)
);

INVx4_ASAP7_75t_L g1097 ( 
.A(n_1008),
.Y(n_1097)
);

AND2x4_ASAP7_75t_L g1098 ( 
.A(n_1005),
.B(n_621),
.Y(n_1098)
);

CKINVDCx5p33_ASAP7_75t_R g1099 ( 
.A(n_1054),
.Y(n_1099)
);

NAND2xp5_ASAP7_75t_L g1100 ( 
.A(n_1063),
.B(n_567),
.Y(n_1100)
);

INVx2_ASAP7_75t_L g1101 ( 
.A(n_1078),
.Y(n_1101)
);

INVx4_ASAP7_75t_L g1102 ( 
.A(n_1008),
.Y(n_1102)
);

BUFx6f_ASAP7_75t_SL g1103 ( 
.A(n_1063),
.Y(n_1103)
);

INVx4_ASAP7_75t_L g1104 ( 
.A(n_1055),
.Y(n_1104)
);

INVx1_ASAP7_75t_L g1105 ( 
.A(n_1078),
.Y(n_1105)
);

BUFx6f_ASAP7_75t_L g1106 ( 
.A(n_1055),
.Y(n_1106)
);

AND2x2_ASAP7_75t_L g1107 ( 
.A(n_1042),
.B(n_695),
.Y(n_1107)
);

AND2x2_ASAP7_75t_L g1108 ( 
.A(n_1042),
.B(n_695),
.Y(n_1108)
);

INVx1_ASAP7_75t_L g1109 ( 
.A(n_1005),
.Y(n_1109)
);

BUFx2_ASAP7_75t_L g1110 ( 
.A(n_1048),
.Y(n_1110)
);

INVx1_ASAP7_75t_L g1111 ( 
.A(n_1049),
.Y(n_1111)
);

INVx1_ASAP7_75t_L g1112 ( 
.A(n_1049),
.Y(n_1112)
);

CKINVDCx5p33_ASAP7_75t_R g1113 ( 
.A(n_1030),
.Y(n_1113)
);

NAND2xp5_ASAP7_75t_L g1114 ( 
.A(n_1088),
.B(n_833),
.Y(n_1114)
);

NAND2xp5_ASAP7_75t_L g1115 ( 
.A(n_1079),
.B(n_998),
.Y(n_1115)
);

NAND2xp5_ASAP7_75t_L g1116 ( 
.A(n_1080),
.B(n_998),
.Y(n_1116)
);

NAND2xp5_ASAP7_75t_L g1117 ( 
.A(n_1081),
.B(n_594),
.Y(n_1117)
);

BUFx6f_ASAP7_75t_L g1118 ( 
.A(n_1055),
.Y(n_1118)
);

INVxp33_ASAP7_75t_SL g1119 ( 
.A(n_1030),
.Y(n_1119)
);

BUFx6f_ASAP7_75t_L g1120 ( 
.A(n_1055),
.Y(n_1120)
);

CKINVDCx20_ASAP7_75t_R g1121 ( 
.A(n_1034),
.Y(n_1121)
);

INVx4_ASAP7_75t_L g1122 ( 
.A(n_1060),
.Y(n_1122)
);

INVx2_ASAP7_75t_L g1123 ( 
.A(n_1076),
.Y(n_1123)
);

INVx2_ASAP7_75t_L g1124 ( 
.A(n_1006),
.Y(n_1124)
);

CKINVDCx20_ASAP7_75t_R g1125 ( 
.A(n_1038),
.Y(n_1125)
);

INVx1_ASAP7_75t_L g1126 ( 
.A(n_1007),
.Y(n_1126)
);

INVx2_ASAP7_75t_L g1127 ( 
.A(n_1009),
.Y(n_1127)
);

INVx1_ASAP7_75t_L g1128 ( 
.A(n_1011),
.Y(n_1128)
);

NOR2xp33_ASAP7_75t_L g1129 ( 
.A(n_1031),
.B(n_706),
.Y(n_1129)
);

INVx3_ASAP7_75t_L g1130 ( 
.A(n_1012),
.Y(n_1130)
);

INVx4_ASAP7_75t_L g1131 ( 
.A(n_1060),
.Y(n_1131)
);

AND2x2_ASAP7_75t_L g1132 ( 
.A(n_1083),
.B(n_706),
.Y(n_1132)
);

INVx2_ASAP7_75t_L g1133 ( 
.A(n_1013),
.Y(n_1133)
);

INVx1_ASAP7_75t_L g1134 ( 
.A(n_1014),
.Y(n_1134)
);

INVx1_ASAP7_75t_L g1135 ( 
.A(n_1016),
.Y(n_1135)
);

NAND2xp5_ASAP7_75t_L g1136 ( 
.A(n_1086),
.B(n_594),
.Y(n_1136)
);

AND2x2_ASAP7_75t_L g1137 ( 
.A(n_1087),
.B(n_1090),
.Y(n_1137)
);

BUFx6f_ASAP7_75t_L g1138 ( 
.A(n_1017),
.Y(n_1138)
);

HB1xp67_ASAP7_75t_L g1139 ( 
.A(n_1048),
.Y(n_1139)
);

INVxp33_ASAP7_75t_L g1140 ( 
.A(n_1010),
.Y(n_1140)
);

INVx2_ASAP7_75t_L g1141 ( 
.A(n_1018),
.Y(n_1141)
);

INVx1_ASAP7_75t_L g1142 ( 
.A(n_1019),
.Y(n_1142)
);

CKINVDCx5p33_ASAP7_75t_R g1143 ( 
.A(n_1031),
.Y(n_1143)
);

INVx1_ASAP7_75t_L g1144 ( 
.A(n_1020),
.Y(n_1144)
);

NAND2xp5_ASAP7_75t_SL g1145 ( 
.A(n_1040),
.B(n_778),
.Y(n_1145)
);

INVx3_ASAP7_75t_L g1146 ( 
.A(n_1021),
.Y(n_1146)
);

CKINVDCx20_ASAP7_75t_R g1147 ( 
.A(n_1038),
.Y(n_1147)
);

CKINVDCx5p33_ASAP7_75t_R g1148 ( 
.A(n_1040),
.Y(n_1148)
);

INVx1_ASAP7_75t_L g1149 ( 
.A(n_1022),
.Y(n_1149)
);

INVx1_ASAP7_75t_L g1150 ( 
.A(n_1027),
.Y(n_1150)
);

CKINVDCx20_ASAP7_75t_R g1151 ( 
.A(n_1044),
.Y(n_1151)
);

INVx1_ASAP7_75t_L g1152 ( 
.A(n_1029),
.Y(n_1152)
);

INVx1_ASAP7_75t_L g1153 ( 
.A(n_1032),
.Y(n_1153)
);

INVx2_ASAP7_75t_L g1154 ( 
.A(n_1033),
.Y(n_1154)
);

INVx1_ASAP7_75t_L g1155 ( 
.A(n_1035),
.Y(n_1155)
);

INVx1_ASAP7_75t_L g1156 ( 
.A(n_1036),
.Y(n_1156)
);

AND2x4_ASAP7_75t_L g1157 ( 
.A(n_1037),
.B(n_778),
.Y(n_1157)
);

BUFx6f_ASAP7_75t_L g1158 ( 
.A(n_1039),
.Y(n_1158)
);

OAI22xp5_ASAP7_75t_L g1159 ( 
.A1(n_1085),
.A2(n_1069),
.B1(n_1025),
.B2(n_1056),
.Y(n_1159)
);

AND2x4_ASAP7_75t_L g1160 ( 
.A(n_1041),
.B(n_872),
.Y(n_1160)
);

CKINVDCx5p33_ASAP7_75t_R g1161 ( 
.A(n_1092),
.Y(n_1161)
);

INVx1_ASAP7_75t_L g1162 ( 
.A(n_1043),
.Y(n_1162)
);

INVx1_ASAP7_75t_L g1163 ( 
.A(n_1046),
.Y(n_1163)
);

AOI22xp33_ASAP7_75t_L g1164 ( 
.A1(n_1157),
.A2(n_873),
.B1(n_986),
.B2(n_853),
.Y(n_1164)
);

CKINVDCx6p67_ASAP7_75t_R g1165 ( 
.A(n_1103),
.Y(n_1165)
);

BUFx6f_ASAP7_75t_L g1166 ( 
.A(n_1106),
.Y(n_1166)
);

INVx2_ASAP7_75t_L g1167 ( 
.A(n_1101),
.Y(n_1167)
);

NAND2xp5_ASAP7_75t_SL g1168 ( 
.A(n_1129),
.B(n_1045),
.Y(n_1168)
);

INVx2_ASAP7_75t_L g1169 ( 
.A(n_1101),
.Y(n_1169)
);

INVx5_ASAP7_75t_L g1170 ( 
.A(n_1106),
.Y(n_1170)
);

HB1xp67_ASAP7_75t_L g1171 ( 
.A(n_1107),
.Y(n_1171)
);

NOR2xp67_ASAP7_75t_L g1172 ( 
.A(n_1094),
.B(n_774),
.Y(n_1172)
);

CKINVDCx6p67_ASAP7_75t_R g1173 ( 
.A(n_1103),
.Y(n_1173)
);

NAND2xp5_ASAP7_75t_L g1174 ( 
.A(n_1130),
.B(n_1047),
.Y(n_1174)
);

NOR2xp33_ASAP7_75t_L g1175 ( 
.A(n_1100),
.B(n_1061),
.Y(n_1175)
);

AND2x2_ASAP7_75t_L g1176 ( 
.A(n_1107),
.B(n_1050),
.Y(n_1176)
);

INVx2_ASAP7_75t_L g1177 ( 
.A(n_1105),
.Y(n_1177)
);

INVx3_ASAP7_75t_L g1178 ( 
.A(n_1106),
.Y(n_1178)
);

INVx2_ASAP7_75t_L g1179 ( 
.A(n_1105),
.Y(n_1179)
);

INVx4_ASAP7_75t_L g1180 ( 
.A(n_1106),
.Y(n_1180)
);

INVx1_ASAP7_75t_L g1181 ( 
.A(n_1138),
.Y(n_1181)
);

NAND2xp5_ASAP7_75t_L g1182 ( 
.A(n_1130),
.B(n_1146),
.Y(n_1182)
);

INVx2_ASAP7_75t_L g1183 ( 
.A(n_1106),
.Y(n_1183)
);

INVx3_ASAP7_75t_L g1184 ( 
.A(n_1118),
.Y(n_1184)
);

INVx2_ASAP7_75t_L g1185 ( 
.A(n_1118),
.Y(n_1185)
);

CKINVDCx6p67_ASAP7_75t_R g1186 ( 
.A(n_1103),
.Y(n_1186)
);

CKINVDCx20_ASAP7_75t_R g1187 ( 
.A(n_1096),
.Y(n_1187)
);

INVx2_ASAP7_75t_L g1188 ( 
.A(n_1118),
.Y(n_1188)
);

INVx1_ASAP7_75t_L g1189 ( 
.A(n_1138),
.Y(n_1189)
);

INVx3_ASAP7_75t_L g1190 ( 
.A(n_1118),
.Y(n_1190)
);

INVx1_ASAP7_75t_L g1191 ( 
.A(n_1138),
.Y(n_1191)
);

BUFx3_ASAP7_75t_L g1192 ( 
.A(n_1095),
.Y(n_1192)
);

INVx1_ASAP7_75t_L g1193 ( 
.A(n_1138),
.Y(n_1193)
);

AOI22xp33_ASAP7_75t_L g1194 ( 
.A1(n_1157),
.A2(n_1160),
.B1(n_1098),
.B2(n_1132),
.Y(n_1194)
);

INVx2_ASAP7_75t_L g1195 ( 
.A(n_1118),
.Y(n_1195)
);

INVx1_ASAP7_75t_L g1196 ( 
.A(n_1138),
.Y(n_1196)
);

NAND2xp5_ASAP7_75t_L g1197 ( 
.A(n_1130),
.B(n_1051),
.Y(n_1197)
);

INVx2_ASAP7_75t_L g1198 ( 
.A(n_1120),
.Y(n_1198)
);

NOR2xp33_ASAP7_75t_L g1199 ( 
.A(n_1145),
.B(n_1061),
.Y(n_1199)
);

AND2x4_ASAP7_75t_L g1200 ( 
.A(n_1137),
.B(n_872),
.Y(n_1200)
);

NAND2xp33_ASAP7_75t_SL g1201 ( 
.A(n_1140),
.B(n_1025),
.Y(n_1201)
);

NAND2xp5_ASAP7_75t_SL g1202 ( 
.A(n_1122),
.B(n_1074),
.Y(n_1202)
);

AOI22xp33_ASAP7_75t_L g1203 ( 
.A1(n_1157),
.A2(n_986),
.B1(n_873),
.B2(n_1023),
.Y(n_1203)
);

OR2x2_ASAP7_75t_L g1204 ( 
.A(n_1159),
.B(n_1024),
.Y(n_1204)
);

NAND2xp5_ASAP7_75t_SL g1205 ( 
.A(n_1122),
.B(n_1074),
.Y(n_1205)
);

NAND2xp5_ASAP7_75t_SL g1206 ( 
.A(n_1122),
.B(n_1077),
.Y(n_1206)
);

NOR2xp33_ASAP7_75t_L g1207 ( 
.A(n_1114),
.B(n_1077),
.Y(n_1207)
);

NAND3xp33_ASAP7_75t_L g1208 ( 
.A(n_1152),
.B(n_1058),
.C(n_1053),
.Y(n_1208)
);

INVxp67_ASAP7_75t_L g1209 ( 
.A(n_1108),
.Y(n_1209)
);

NAND2xp5_ASAP7_75t_L g1210 ( 
.A(n_1146),
.B(n_1059),
.Y(n_1210)
);

CKINVDCx5p33_ASAP7_75t_R g1211 ( 
.A(n_1093),
.Y(n_1211)
);

INVx1_ASAP7_75t_L g1212 ( 
.A(n_1158),
.Y(n_1212)
);

INVx2_ASAP7_75t_L g1213 ( 
.A(n_1120),
.Y(n_1213)
);

HB1xp67_ASAP7_75t_L g1214 ( 
.A(n_1108),
.Y(n_1214)
);

BUFx3_ASAP7_75t_L g1215 ( 
.A(n_1095),
.Y(n_1215)
);

INVx2_ASAP7_75t_L g1216 ( 
.A(n_1120),
.Y(n_1216)
);

NAND2xp5_ASAP7_75t_L g1217 ( 
.A(n_1146),
.B(n_1062),
.Y(n_1217)
);

INVx2_ASAP7_75t_L g1218 ( 
.A(n_1120),
.Y(n_1218)
);

NAND2xp33_ASAP7_75t_SL g1219 ( 
.A(n_1113),
.B(n_1052),
.Y(n_1219)
);

INVx2_ASAP7_75t_L g1220 ( 
.A(n_1120),
.Y(n_1220)
);

AND2x2_ASAP7_75t_L g1221 ( 
.A(n_1098),
.B(n_1064),
.Y(n_1221)
);

INVx2_ASAP7_75t_L g1222 ( 
.A(n_1095),
.Y(n_1222)
);

INVx1_ASAP7_75t_L g1223 ( 
.A(n_1158),
.Y(n_1223)
);

INVx1_ASAP7_75t_L g1224 ( 
.A(n_1158),
.Y(n_1224)
);

NAND2xp5_ASAP7_75t_L g1225 ( 
.A(n_1098),
.B(n_1065),
.Y(n_1225)
);

INVx4_ASAP7_75t_L g1226 ( 
.A(n_1158),
.Y(n_1226)
);

INVx1_ASAP7_75t_L g1227 ( 
.A(n_1158),
.Y(n_1227)
);

INVx2_ASAP7_75t_SL g1228 ( 
.A(n_1137),
.Y(n_1228)
);

NAND2xp5_ASAP7_75t_SL g1229 ( 
.A(n_1194),
.B(n_1131),
.Y(n_1229)
);

NAND2xp5_ASAP7_75t_SL g1230 ( 
.A(n_1207),
.B(n_1131),
.Y(n_1230)
);

INVx1_ASAP7_75t_L g1231 ( 
.A(n_1182),
.Y(n_1231)
);

NAND2xp5_ASAP7_75t_L g1232 ( 
.A(n_1228),
.B(n_1160),
.Y(n_1232)
);

NAND2xp5_ASAP7_75t_L g1233 ( 
.A(n_1228),
.B(n_1160),
.Y(n_1233)
);

NOR2xp33_ASAP7_75t_L g1234 ( 
.A(n_1209),
.B(n_1131),
.Y(n_1234)
);

INVx2_ASAP7_75t_SL g1235 ( 
.A(n_1176),
.Y(n_1235)
);

INVx2_ASAP7_75t_SL g1236 ( 
.A(n_1176),
.Y(n_1236)
);

NAND2xp5_ASAP7_75t_SL g1237 ( 
.A(n_1209),
.B(n_1093),
.Y(n_1237)
);

INVxp67_ASAP7_75t_L g1238 ( 
.A(n_1201),
.Y(n_1238)
);

AOI22xp5_ASAP7_75t_L g1239 ( 
.A1(n_1175),
.A2(n_1228),
.B1(n_1199),
.B2(n_1214),
.Y(n_1239)
);

INVx1_ASAP7_75t_L g1240 ( 
.A(n_1182),
.Y(n_1240)
);

INVx4_ASAP7_75t_L g1241 ( 
.A(n_1226),
.Y(n_1241)
);

NAND2xp5_ASAP7_75t_SL g1242 ( 
.A(n_1171),
.B(n_1119),
.Y(n_1242)
);

A2O1A1Ixp33_ASAP7_75t_L g1243 ( 
.A1(n_1225),
.A2(n_1132),
.B(n_774),
.C(n_761),
.Y(n_1243)
);

NAND2xp5_ASAP7_75t_L g1244 ( 
.A(n_1171),
.B(n_1126),
.Y(n_1244)
);

INVx2_ASAP7_75t_L g1245 ( 
.A(n_1177),
.Y(n_1245)
);

NAND2xp5_ASAP7_75t_L g1246 ( 
.A(n_1214),
.B(n_1128),
.Y(n_1246)
);

NAND2xp5_ASAP7_75t_L g1247 ( 
.A(n_1221),
.B(n_1134),
.Y(n_1247)
);

INVx2_ASAP7_75t_L g1248 ( 
.A(n_1177),
.Y(n_1248)
);

INVx2_ASAP7_75t_L g1249 ( 
.A(n_1177),
.Y(n_1249)
);

INVx1_ASAP7_75t_L g1250 ( 
.A(n_1174),
.Y(n_1250)
);

INVxp67_ASAP7_75t_SL g1251 ( 
.A(n_1166),
.Y(n_1251)
);

AND2x2_ASAP7_75t_SL g1252 ( 
.A(n_1164),
.B(n_649),
.Y(n_1252)
);

NAND2xp5_ASAP7_75t_L g1253 ( 
.A(n_1221),
.B(n_1135),
.Y(n_1253)
);

INVx1_ASAP7_75t_L g1254 ( 
.A(n_1174),
.Y(n_1254)
);

NAND2xp5_ASAP7_75t_SL g1255 ( 
.A(n_1211),
.B(n_1200),
.Y(n_1255)
);

INVx2_ASAP7_75t_L g1256 ( 
.A(n_1179),
.Y(n_1256)
);

INVx2_ASAP7_75t_L g1257 ( 
.A(n_1179),
.Y(n_1257)
);

AOI22xp5_ASAP7_75t_L g1258 ( 
.A1(n_1225),
.A2(n_600),
.B1(n_748),
.B2(n_730),
.Y(n_1258)
);

NAND2xp5_ASAP7_75t_L g1259 ( 
.A(n_1192),
.B(n_1142),
.Y(n_1259)
);

INVxp67_ASAP7_75t_L g1260 ( 
.A(n_1168),
.Y(n_1260)
);

INVx3_ASAP7_75t_L g1261 ( 
.A(n_1192),
.Y(n_1261)
);

BUFx6f_ASAP7_75t_L g1262 ( 
.A(n_1192),
.Y(n_1262)
);

NAND2xp5_ASAP7_75t_L g1263 ( 
.A(n_1215),
.B(n_1144),
.Y(n_1263)
);

NAND2xp5_ASAP7_75t_L g1264 ( 
.A(n_1215),
.B(n_1149),
.Y(n_1264)
);

AND2x4_ASAP7_75t_L g1265 ( 
.A(n_1200),
.B(n_1163),
.Y(n_1265)
);

INVx2_ASAP7_75t_L g1266 ( 
.A(n_1179),
.Y(n_1266)
);

NOR2xp67_ASAP7_75t_L g1267 ( 
.A(n_1208),
.B(n_1113),
.Y(n_1267)
);

BUFx2_ASAP7_75t_L g1268 ( 
.A(n_1187),
.Y(n_1268)
);

NOR2xp33_ASAP7_75t_L g1269 ( 
.A(n_1202),
.B(n_1119),
.Y(n_1269)
);

INVx1_ASAP7_75t_L g1270 ( 
.A(n_1197),
.Y(n_1270)
);

INVx1_ASAP7_75t_L g1271 ( 
.A(n_1197),
.Y(n_1271)
);

NAND2xp5_ASAP7_75t_SL g1272 ( 
.A(n_1181),
.B(n_562),
.Y(n_1272)
);

INVx1_ASAP7_75t_L g1273 ( 
.A(n_1210),
.Y(n_1273)
);

NOR2xp33_ASAP7_75t_L g1274 ( 
.A(n_1205),
.B(n_1084),
.Y(n_1274)
);

NOR2xp33_ASAP7_75t_L g1275 ( 
.A(n_1206),
.B(n_1084),
.Y(n_1275)
);

NAND2xp5_ASAP7_75t_SL g1276 ( 
.A(n_1200),
.B(n_1143),
.Y(n_1276)
);

NAND2xp5_ASAP7_75t_SL g1277 ( 
.A(n_1200),
.B(n_1143),
.Y(n_1277)
);

INVx2_ASAP7_75t_L g1278 ( 
.A(n_1167),
.Y(n_1278)
);

AOI22xp33_ASAP7_75t_L g1279 ( 
.A1(n_1203),
.A2(n_611),
.B1(n_619),
.B2(n_601),
.Y(n_1279)
);

INVx2_ASAP7_75t_L g1280 ( 
.A(n_1167),
.Y(n_1280)
);

NOR2xp33_ASAP7_75t_L g1281 ( 
.A(n_1204),
.B(n_1089),
.Y(n_1281)
);

INVxp67_ASAP7_75t_L g1282 ( 
.A(n_1204),
.Y(n_1282)
);

NAND2xp5_ASAP7_75t_L g1283 ( 
.A(n_1215),
.B(n_1150),
.Y(n_1283)
);

CKINVDCx5p33_ASAP7_75t_R g1284 ( 
.A(n_1165),
.Y(n_1284)
);

NAND2xp5_ASAP7_75t_L g1285 ( 
.A(n_1181),
.B(n_1089),
.Y(n_1285)
);

INVx2_ASAP7_75t_L g1286 ( 
.A(n_1167),
.Y(n_1286)
);

INVx1_ASAP7_75t_L g1287 ( 
.A(n_1210),
.Y(n_1287)
);

OAI21xp5_ASAP7_75t_L g1288 ( 
.A1(n_1189),
.A2(n_1136),
.B(n_1117),
.Y(n_1288)
);

A2O1A1Ixp33_ASAP7_75t_L g1289 ( 
.A1(n_1217),
.A2(n_761),
.B(n_896),
.C(n_649),
.Y(n_1289)
);

NAND2xp5_ASAP7_75t_L g1290 ( 
.A(n_1189),
.B(n_1152),
.Y(n_1290)
);

NAND2xp5_ASAP7_75t_SL g1291 ( 
.A(n_1217),
.B(n_1148),
.Y(n_1291)
);

NAND2xp5_ASAP7_75t_SL g1292 ( 
.A(n_1172),
.B(n_1148),
.Y(n_1292)
);

NOR2xp67_ASAP7_75t_L g1293 ( 
.A(n_1208),
.B(n_1139),
.Y(n_1293)
);

INVx2_ASAP7_75t_L g1294 ( 
.A(n_1169),
.Y(n_1294)
);

INVxp67_ASAP7_75t_L g1295 ( 
.A(n_1219),
.Y(n_1295)
);

INVxp67_ASAP7_75t_L g1296 ( 
.A(n_1172),
.Y(n_1296)
);

NAND2xp5_ASAP7_75t_L g1297 ( 
.A(n_1191),
.B(n_1153),
.Y(n_1297)
);

NAND2xp5_ASAP7_75t_SL g1298 ( 
.A(n_1191),
.B(n_1161),
.Y(n_1298)
);

NOR2xp33_ASAP7_75t_L g1299 ( 
.A(n_1193),
.B(n_1052),
.Y(n_1299)
);

INVx2_ASAP7_75t_L g1300 ( 
.A(n_1169),
.Y(n_1300)
);

NOR2xp33_ASAP7_75t_R g1301 ( 
.A(n_1165),
.B(n_1099),
.Y(n_1301)
);

INVx2_ASAP7_75t_L g1302 ( 
.A(n_1169),
.Y(n_1302)
);

NAND2xp5_ASAP7_75t_L g1303 ( 
.A(n_1193),
.B(n_1196),
.Y(n_1303)
);

AOI22x1_ASAP7_75t_L g1304 ( 
.A1(n_1183),
.A2(n_896),
.B1(n_1068),
.B2(n_1067),
.Y(n_1304)
);

NAND2xp5_ASAP7_75t_SL g1305 ( 
.A(n_1196),
.B(n_1161),
.Y(n_1305)
);

AND2x6_ASAP7_75t_L g1306 ( 
.A(n_1212),
.B(n_562),
.Y(n_1306)
);

CKINVDCx20_ASAP7_75t_R g1307 ( 
.A(n_1165),
.Y(n_1307)
);

INVx2_ASAP7_75t_L g1308 ( 
.A(n_1222),
.Y(n_1308)
);

NAND2x1_ASAP7_75t_L g1309 ( 
.A(n_1180),
.B(n_1094),
.Y(n_1309)
);

INVxp67_ASAP7_75t_SL g1310 ( 
.A(n_1166),
.Y(n_1310)
);

NAND2xp5_ASAP7_75t_SL g1311 ( 
.A(n_1212),
.B(n_1110),
.Y(n_1311)
);

AOI22xp33_ASAP7_75t_L g1312 ( 
.A1(n_1223),
.A2(n_611),
.B1(n_619),
.B2(n_601),
.Y(n_1312)
);

INVx2_ASAP7_75t_L g1313 ( 
.A(n_1222),
.Y(n_1313)
);

INVx2_ASAP7_75t_L g1314 ( 
.A(n_1222),
.Y(n_1314)
);

NAND2xp5_ASAP7_75t_L g1315 ( 
.A(n_1223),
.B(n_1153),
.Y(n_1315)
);

INVx1_ASAP7_75t_L g1316 ( 
.A(n_1245),
.Y(n_1316)
);

NAND2xp5_ASAP7_75t_SL g1317 ( 
.A(n_1239),
.B(n_1110),
.Y(n_1317)
);

AOI22xp5_ASAP7_75t_L g1318 ( 
.A1(n_1229),
.A2(n_865),
.B1(n_1227),
.B2(n_1224),
.Y(n_1318)
);

INVx1_ASAP7_75t_L g1319 ( 
.A(n_1245),
.Y(n_1319)
);

AND2x2_ASAP7_75t_L g1320 ( 
.A(n_1235),
.B(n_1173),
.Y(n_1320)
);

INVx2_ASAP7_75t_L g1321 ( 
.A(n_1248),
.Y(n_1321)
);

NAND2xp5_ASAP7_75t_L g1322 ( 
.A(n_1231),
.B(n_1224),
.Y(n_1322)
);

NOR2xp33_ASAP7_75t_L g1323 ( 
.A(n_1281),
.B(n_1044),
.Y(n_1323)
);

INVx2_ASAP7_75t_L g1324 ( 
.A(n_1248),
.Y(n_1324)
);

BUFx3_ASAP7_75t_L g1325 ( 
.A(n_1268),
.Y(n_1325)
);

INVx1_ASAP7_75t_L g1326 ( 
.A(n_1249),
.Y(n_1326)
);

NAND2xp5_ASAP7_75t_SL g1327 ( 
.A(n_1236),
.B(n_1099),
.Y(n_1327)
);

OAI22xp5_ASAP7_75t_L g1328 ( 
.A1(n_1252),
.A2(n_558),
.B1(n_570),
.B2(n_564),
.Y(n_1328)
);

AND2x4_ASAP7_75t_L g1329 ( 
.A(n_1265),
.B(n_1155),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_1249),
.Y(n_1330)
);

INVx1_ASAP7_75t_L g1331 ( 
.A(n_1256),
.Y(n_1331)
);

OR2x6_ASAP7_75t_L g1332 ( 
.A(n_1255),
.B(n_556),
.Y(n_1332)
);

NAND2xp5_ASAP7_75t_L g1333 ( 
.A(n_1240),
.B(n_1227),
.Y(n_1333)
);

NAND2xp5_ASAP7_75t_L g1334 ( 
.A(n_1250),
.B(n_1178),
.Y(n_1334)
);

INVx1_ASAP7_75t_SL g1335 ( 
.A(n_1242),
.Y(n_1335)
);

NAND2xp5_ASAP7_75t_SL g1336 ( 
.A(n_1234),
.B(n_1226),
.Y(n_1336)
);

NAND2xp5_ASAP7_75t_L g1337 ( 
.A(n_1254),
.B(n_1178),
.Y(n_1337)
);

BUFx6f_ASAP7_75t_L g1338 ( 
.A(n_1262),
.Y(n_1338)
);

NAND2xp5_ASAP7_75t_SL g1339 ( 
.A(n_1234),
.B(n_1226),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_1256),
.Y(n_1340)
);

NAND2xp5_ASAP7_75t_L g1341 ( 
.A(n_1270),
.B(n_1183),
.Y(n_1341)
);

BUFx6f_ASAP7_75t_L g1342 ( 
.A(n_1262),
.Y(n_1342)
);

INVx1_ASAP7_75t_L g1343 ( 
.A(n_1257),
.Y(n_1343)
);

AO21x1_ASAP7_75t_L g1344 ( 
.A1(n_1230),
.A2(n_1226),
.B(n_576),
.Y(n_1344)
);

NAND2xp5_ASAP7_75t_L g1345 ( 
.A(n_1271),
.B(n_1178),
.Y(n_1345)
);

INVx1_ASAP7_75t_L g1346 ( 
.A(n_1257),
.Y(n_1346)
);

AOI22xp33_ASAP7_75t_L g1347 ( 
.A1(n_1252),
.A2(n_562),
.B1(n_638),
.B2(n_817),
.Y(n_1347)
);

INVx3_ASAP7_75t_L g1348 ( 
.A(n_1262),
.Y(n_1348)
);

INVx2_ASAP7_75t_L g1349 ( 
.A(n_1266),
.Y(n_1349)
);

AOI22xp33_ASAP7_75t_L g1350 ( 
.A1(n_1273),
.A2(n_638),
.B1(n_817),
.B2(n_666),
.Y(n_1350)
);

OR2x2_ASAP7_75t_L g1351 ( 
.A(n_1282),
.B(n_1026),
.Y(n_1351)
);

INVx1_ASAP7_75t_L g1352 ( 
.A(n_1266),
.Y(n_1352)
);

OAI22x1_ASAP7_75t_SL g1353 ( 
.A1(n_1307),
.A2(n_1066),
.B1(n_1073),
.B2(n_1057),
.Y(n_1353)
);

NAND2xp5_ASAP7_75t_L g1354 ( 
.A(n_1287),
.B(n_1183),
.Y(n_1354)
);

INVx2_ASAP7_75t_L g1355 ( 
.A(n_1278),
.Y(n_1355)
);

INVx1_ASAP7_75t_L g1356 ( 
.A(n_1290),
.Y(n_1356)
);

OR2x2_ASAP7_75t_L g1357 ( 
.A(n_1258),
.B(n_1028),
.Y(n_1357)
);

AOI22xp5_ASAP7_75t_L g1358 ( 
.A1(n_1232),
.A2(n_1186),
.B1(n_1173),
.B2(n_1066),
.Y(n_1358)
);

NOR2xp33_ASAP7_75t_L g1359 ( 
.A(n_1281),
.B(n_1057),
.Y(n_1359)
);

AOI22xp5_ASAP7_75t_L g1360 ( 
.A1(n_1233),
.A2(n_1275),
.B1(n_1274),
.B2(n_1238),
.Y(n_1360)
);

CKINVDCx5p33_ASAP7_75t_R g1361 ( 
.A(n_1301),
.Y(n_1361)
);

NAND2xp5_ASAP7_75t_L g1362 ( 
.A(n_1247),
.B(n_1185),
.Y(n_1362)
);

INVx2_ASAP7_75t_L g1363 ( 
.A(n_1278),
.Y(n_1363)
);

AND2x2_ASAP7_75t_SL g1364 ( 
.A(n_1269),
.B(n_967),
.Y(n_1364)
);

AND2x2_ASAP7_75t_L g1365 ( 
.A(n_1260),
.B(n_1173),
.Y(n_1365)
);

INVx1_ASAP7_75t_L g1366 ( 
.A(n_1297),
.Y(n_1366)
);

CKINVDCx5p33_ASAP7_75t_R g1367 ( 
.A(n_1301),
.Y(n_1367)
);

NAND2xp5_ASAP7_75t_L g1368 ( 
.A(n_1253),
.B(n_1185),
.Y(n_1368)
);

INVx2_ASAP7_75t_L g1369 ( 
.A(n_1280),
.Y(n_1369)
);

AND2x6_ASAP7_75t_SL g1370 ( 
.A(n_1269),
.B(n_1274),
.Y(n_1370)
);

INVx2_ASAP7_75t_L g1371 ( 
.A(n_1280),
.Y(n_1371)
);

AOI22xp33_ASAP7_75t_L g1372 ( 
.A1(n_1265),
.A2(n_638),
.B1(n_817),
.B2(n_584),
.Y(n_1372)
);

NAND2xp5_ASAP7_75t_L g1373 ( 
.A(n_1286),
.B(n_1185),
.Y(n_1373)
);

INVx5_ASAP7_75t_L g1374 ( 
.A(n_1241),
.Y(n_1374)
);

NAND2xp5_ASAP7_75t_SL g1375 ( 
.A(n_1275),
.B(n_1124),
.Y(n_1375)
);

NAND2xp5_ASAP7_75t_SL g1376 ( 
.A(n_1267),
.B(n_1124),
.Y(n_1376)
);

NAND2xp5_ASAP7_75t_L g1377 ( 
.A(n_1286),
.B(n_1188),
.Y(n_1377)
);

HB1xp67_ASAP7_75t_L g1378 ( 
.A(n_1244),
.Y(n_1378)
);

BUFx4f_ASAP7_75t_L g1379 ( 
.A(n_1262),
.Y(n_1379)
);

BUFx8_ASAP7_75t_L g1380 ( 
.A(n_1284),
.Y(n_1380)
);

CKINVDCx20_ASAP7_75t_R g1381 ( 
.A(n_1237),
.Y(n_1381)
);

NAND2xp5_ASAP7_75t_L g1382 ( 
.A(n_1294),
.B(n_1188),
.Y(n_1382)
);

NAND2xp5_ASAP7_75t_L g1383 ( 
.A(n_1294),
.B(n_1188),
.Y(n_1383)
);

NAND2xp5_ASAP7_75t_L g1384 ( 
.A(n_1300),
.B(n_1195),
.Y(n_1384)
);

NOR3xp33_ASAP7_75t_SL g1385 ( 
.A(n_1276),
.B(n_1028),
.C(n_593),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_1315),
.Y(n_1386)
);

BUFx6f_ASAP7_75t_L g1387 ( 
.A(n_1261),
.Y(n_1387)
);

INVx1_ASAP7_75t_L g1388 ( 
.A(n_1300),
.Y(n_1388)
);

AOI22xp33_ASAP7_75t_L g1389 ( 
.A1(n_1288),
.A2(n_638),
.B1(n_817),
.B2(n_982),
.Y(n_1389)
);

NAND2xp5_ASAP7_75t_L g1390 ( 
.A(n_1302),
.B(n_1195),
.Y(n_1390)
);

NOR2xp33_ASAP7_75t_L g1391 ( 
.A(n_1291),
.B(n_1073),
.Y(n_1391)
);

AOI22xp33_ASAP7_75t_L g1392 ( 
.A1(n_1261),
.A2(n_638),
.B1(n_817),
.B2(n_1195),
.Y(n_1392)
);

BUFx2_ASAP7_75t_L g1393 ( 
.A(n_1295),
.Y(n_1393)
);

INVx5_ASAP7_75t_L g1394 ( 
.A(n_1241),
.Y(n_1394)
);

INVx2_ASAP7_75t_SL g1395 ( 
.A(n_1246),
.Y(n_1395)
);

AND2x6_ASAP7_75t_SL g1396 ( 
.A(n_1299),
.B(n_558),
.Y(n_1396)
);

AND2x2_ASAP7_75t_L g1397 ( 
.A(n_1299),
.B(n_1186),
.Y(n_1397)
);

AOI22xp33_ASAP7_75t_L g1398 ( 
.A1(n_1259),
.A2(n_817),
.B1(n_1213),
.B2(n_1198),
.Y(n_1398)
);

OAI21xp33_ASAP7_75t_L g1399 ( 
.A1(n_1279),
.A2(n_1277),
.B(n_1285),
.Y(n_1399)
);

AOI22xp33_ASAP7_75t_L g1400 ( 
.A1(n_1263),
.A2(n_817),
.B1(n_1213),
.B2(n_1198),
.Y(n_1400)
);

BUFx2_ASAP7_75t_L g1401 ( 
.A(n_1264),
.Y(n_1401)
);

INVx1_ASAP7_75t_L g1402 ( 
.A(n_1302),
.Y(n_1402)
);

INVx1_ASAP7_75t_L g1403 ( 
.A(n_1308),
.Y(n_1403)
);

HB1xp67_ASAP7_75t_L g1404 ( 
.A(n_1293),
.Y(n_1404)
);

A2O1A1Ixp33_ASAP7_75t_L g1405 ( 
.A1(n_1243),
.A2(n_1156),
.B(n_1162),
.C(n_1155),
.Y(n_1405)
);

AOI22xp5_ASAP7_75t_L g1406 ( 
.A1(n_1283),
.A2(n_1186),
.B1(n_1082),
.B2(n_1184),
.Y(n_1406)
);

NAND2xp5_ASAP7_75t_L g1407 ( 
.A(n_1308),
.B(n_1198),
.Y(n_1407)
);

AND2x2_ASAP7_75t_L g1408 ( 
.A(n_1311),
.B(n_1082),
.Y(n_1408)
);

BUFx3_ASAP7_75t_L g1409 ( 
.A(n_1313),
.Y(n_1409)
);

NOR2xp33_ASAP7_75t_L g1410 ( 
.A(n_1292),
.B(n_1121),
.Y(n_1410)
);

NAND2xp5_ASAP7_75t_SL g1411 ( 
.A(n_1296),
.B(n_1127),
.Y(n_1411)
);

NAND2xp5_ASAP7_75t_L g1412 ( 
.A(n_1313),
.B(n_1213),
.Y(n_1412)
);

INVx1_ASAP7_75t_L g1413 ( 
.A(n_1314),
.Y(n_1413)
);

AND2x2_ASAP7_75t_L g1414 ( 
.A(n_1298),
.B(n_1091),
.Y(n_1414)
);

NAND2xp5_ASAP7_75t_L g1415 ( 
.A(n_1314),
.B(n_1216),
.Y(n_1415)
);

NAND2xp5_ASAP7_75t_L g1416 ( 
.A(n_1251),
.B(n_1216),
.Y(n_1416)
);

INVx1_ASAP7_75t_L g1417 ( 
.A(n_1303),
.Y(n_1417)
);

NAND2xp5_ASAP7_75t_L g1418 ( 
.A(n_1310),
.B(n_1178),
.Y(n_1418)
);

INVx2_ASAP7_75t_SL g1419 ( 
.A(n_1305),
.Y(n_1419)
);

NAND2xp5_ASAP7_75t_L g1420 ( 
.A(n_1312),
.B(n_1216),
.Y(n_1420)
);

INVx2_ASAP7_75t_SL g1421 ( 
.A(n_1272),
.Y(n_1421)
);

AOI22xp5_ASAP7_75t_L g1422 ( 
.A1(n_1272),
.A2(n_1190),
.B1(n_1184),
.B2(n_1218),
.Y(n_1422)
);

INVx1_ASAP7_75t_L g1423 ( 
.A(n_1304),
.Y(n_1423)
);

INVx2_ASAP7_75t_L g1424 ( 
.A(n_1309),
.Y(n_1424)
);

NAND2xp5_ASAP7_75t_SL g1425 ( 
.A(n_1312),
.B(n_1127),
.Y(n_1425)
);

NOR2xp67_ASAP7_75t_L g1426 ( 
.A(n_1279),
.B(n_1115),
.Y(n_1426)
);

INVx1_ASAP7_75t_L g1427 ( 
.A(n_1289),
.Y(n_1427)
);

INVx5_ASAP7_75t_L g1428 ( 
.A(n_1338),
.Y(n_1428)
);

NAND2xp5_ASAP7_75t_SL g1429 ( 
.A(n_1360),
.B(n_1147),
.Y(n_1429)
);

AOI21xp5_ASAP7_75t_L g1430 ( 
.A1(n_1374),
.A2(n_1180),
.B(n_1166),
.Y(n_1430)
);

AOI21xp5_ASAP7_75t_L g1431 ( 
.A1(n_1374),
.A2(n_1180),
.B(n_1166),
.Y(n_1431)
);

NOR2xp33_ASAP7_75t_L g1432 ( 
.A(n_1364),
.B(n_1125),
.Y(n_1432)
);

BUFx6f_ASAP7_75t_L g1433 ( 
.A(n_1338),
.Y(n_1433)
);

O2A1O1Ixp33_ASAP7_75t_L g1434 ( 
.A1(n_1317),
.A2(n_1116),
.B(n_831),
.C(n_586),
.Y(n_1434)
);

NOR2xp33_ASAP7_75t_R g1435 ( 
.A(n_1361),
.B(n_1151),
.Y(n_1435)
);

AOI22xp5_ASAP7_75t_L g1436 ( 
.A1(n_1399),
.A2(n_559),
.B1(n_578),
.B2(n_575),
.Y(n_1436)
);

NAND2xp5_ASAP7_75t_L g1437 ( 
.A(n_1417),
.B(n_1156),
.Y(n_1437)
);

O2A1O1Ixp33_ASAP7_75t_L g1438 ( 
.A1(n_1328),
.A2(n_586),
.B(n_631),
.C(n_556),
.Y(n_1438)
);

OAI22xp5_ASAP7_75t_L g1439 ( 
.A1(n_1328),
.A2(n_701),
.B1(n_737),
.B2(n_711),
.Y(n_1439)
);

AOI22xp33_ASAP7_75t_L g1440 ( 
.A1(n_1426),
.A2(n_817),
.B1(n_962),
.B2(n_1162),
.Y(n_1440)
);

AOI21xp5_ASAP7_75t_L g1441 ( 
.A1(n_1374),
.A2(n_1166),
.B(n_1170),
.Y(n_1441)
);

INVx2_ASAP7_75t_L g1442 ( 
.A(n_1321),
.Y(n_1442)
);

AOI21xp5_ASAP7_75t_L g1443 ( 
.A1(n_1394),
.A2(n_1170),
.B(n_1097),
.Y(n_1443)
);

NAND3xp33_ASAP7_75t_L g1444 ( 
.A(n_1323),
.B(n_595),
.C(n_573),
.Y(n_1444)
);

BUFx3_ASAP7_75t_L g1445 ( 
.A(n_1325),
.Y(n_1445)
);

BUFx6f_ASAP7_75t_L g1446 ( 
.A(n_1338),
.Y(n_1446)
);

AOI21xp5_ASAP7_75t_L g1447 ( 
.A1(n_1394),
.A2(n_1170),
.B(n_1097),
.Y(n_1447)
);

NAND2xp5_ASAP7_75t_L g1448 ( 
.A(n_1356),
.B(n_1133),
.Y(n_1448)
);

OAI21xp5_ASAP7_75t_L g1449 ( 
.A1(n_1427),
.A2(n_1220),
.B(n_1218),
.Y(n_1449)
);

NOR2xp33_ASAP7_75t_L g1450 ( 
.A(n_1359),
.B(n_766),
.Y(n_1450)
);

OAI22xp5_ASAP7_75t_L g1451 ( 
.A1(n_1366),
.A2(n_801),
.B1(n_825),
.B2(n_772),
.Y(n_1451)
);

NOR2xp33_ASAP7_75t_SL g1452 ( 
.A(n_1394),
.B(n_830),
.Y(n_1452)
);

NAND2xp5_ASAP7_75t_L g1453 ( 
.A(n_1386),
.B(n_1133),
.Y(n_1453)
);

AOI22xp5_ASAP7_75t_L g1454 ( 
.A1(n_1391),
.A2(n_630),
.B1(n_637),
.B2(n_583),
.Y(n_1454)
);

A2O1A1Ixp33_ASAP7_75t_L g1455 ( 
.A1(n_1395),
.A2(n_749),
.B(n_888),
.C(n_631),
.Y(n_1455)
);

O2A1O1Ixp33_ASAP7_75t_L g1456 ( 
.A1(n_1378),
.A2(n_888),
.B(n_939),
.C(n_749),
.Y(n_1456)
);

INVx3_ASAP7_75t_L g1457 ( 
.A(n_1342),
.Y(n_1457)
);

AND2x2_ASAP7_75t_SL g1458 ( 
.A(n_1397),
.B(n_636),
.Y(n_1458)
);

AOI21xp5_ASAP7_75t_L g1459 ( 
.A1(n_1394),
.A2(n_1379),
.B(n_1339),
.Y(n_1459)
);

NAND2xp5_ASAP7_75t_L g1460 ( 
.A(n_1401),
.B(n_1141),
.Y(n_1460)
);

AOI21x1_ASAP7_75t_L g1461 ( 
.A1(n_1336),
.A2(n_1220),
.B(n_1218),
.Y(n_1461)
);

NAND2xp5_ASAP7_75t_L g1462 ( 
.A(n_1362),
.B(n_1141),
.Y(n_1462)
);

NAND2xp5_ASAP7_75t_L g1463 ( 
.A(n_1362),
.B(n_1154),
.Y(n_1463)
);

NAND2xp5_ASAP7_75t_L g1464 ( 
.A(n_1368),
.B(n_1154),
.Y(n_1464)
);

NAND2xp5_ASAP7_75t_L g1465 ( 
.A(n_1368),
.B(n_1123),
.Y(n_1465)
);

OAI22xp5_ASAP7_75t_L g1466 ( 
.A1(n_1318),
.A2(n_880),
.B1(n_885),
.B2(n_867),
.Y(n_1466)
);

INVx2_ASAP7_75t_SL g1467 ( 
.A(n_1329),
.Y(n_1467)
);

NOR2xp67_ASAP7_75t_L g1468 ( 
.A(n_1351),
.B(n_1123),
.Y(n_1468)
);

NOR2xp33_ASAP7_75t_L g1469 ( 
.A(n_1370),
.B(n_1335),
.Y(n_1469)
);

OAI22xp5_ASAP7_75t_L g1470 ( 
.A1(n_1322),
.A2(n_900),
.B1(n_955),
.B2(n_890),
.Y(n_1470)
);

INVx1_ASAP7_75t_L g1471 ( 
.A(n_1316),
.Y(n_1471)
);

NAND2xp5_ASAP7_75t_SL g1472 ( 
.A(n_1419),
.B(n_657),
.Y(n_1472)
);

NOR3xp33_ASAP7_75t_L g1473 ( 
.A(n_1327),
.B(n_602),
.C(n_592),
.Y(n_1473)
);

AOI22xp33_ASAP7_75t_L g1474 ( 
.A1(n_1389),
.A2(n_962),
.B1(n_608),
.B2(n_640),
.Y(n_1474)
);

NOR2xp33_ASAP7_75t_L g1475 ( 
.A(n_1393),
.B(n_966),
.Y(n_1475)
);

NOR2xp33_ASAP7_75t_L g1476 ( 
.A(n_1357),
.B(n_978),
.Y(n_1476)
);

NOR3xp33_ASAP7_75t_L g1477 ( 
.A(n_1410),
.B(n_686),
.C(n_664),
.Y(n_1477)
);

INVx2_ASAP7_75t_SL g1478 ( 
.A(n_1329),
.Y(n_1478)
);

BUFx2_ASAP7_75t_L g1479 ( 
.A(n_1381),
.Y(n_1479)
);

AOI21xp5_ASAP7_75t_L g1480 ( 
.A1(n_1379),
.A2(n_1170),
.B(n_1097),
.Y(n_1480)
);

NAND2xp5_ASAP7_75t_L g1481 ( 
.A(n_1322),
.B(n_1184),
.Y(n_1481)
);

OAI22xp5_ASAP7_75t_SL g1482 ( 
.A1(n_1358),
.A2(n_995),
.B1(n_988),
.B2(n_746),
.Y(n_1482)
);

INVx2_ASAP7_75t_L g1483 ( 
.A(n_1324),
.Y(n_1483)
);

NAND2xp5_ASAP7_75t_SL g1484 ( 
.A(n_1365),
.B(n_671),
.Y(n_1484)
);

BUFx12f_ASAP7_75t_L g1485 ( 
.A(n_1380),
.Y(n_1485)
);

OAI21xp33_ASAP7_75t_L g1486 ( 
.A1(n_1414),
.A2(n_847),
.B(n_732),
.Y(n_1486)
);

CKINVDCx14_ASAP7_75t_R g1487 ( 
.A(n_1367),
.Y(n_1487)
);

AOI22xp5_ASAP7_75t_L g1488 ( 
.A1(n_1404),
.A2(n_689),
.B1(n_702),
.B2(n_676),
.Y(n_1488)
);

AOI21xp5_ASAP7_75t_L g1489 ( 
.A1(n_1416),
.A2(n_1170),
.B(n_1104),
.Y(n_1489)
);

NAND2xp5_ASAP7_75t_SL g1490 ( 
.A(n_1406),
.B(n_707),
.Y(n_1490)
);

AND2x4_ASAP7_75t_L g1491 ( 
.A(n_1320),
.B(n_1220),
.Y(n_1491)
);

OAI22x1_ASAP7_75t_L g1492 ( 
.A1(n_1408),
.A2(n_959),
.B1(n_939),
.B2(n_905),
.Y(n_1492)
);

NAND2xp5_ASAP7_75t_SL g1493 ( 
.A(n_1387),
.B(n_715),
.Y(n_1493)
);

AOI22xp33_ASAP7_75t_L g1494 ( 
.A1(n_1375),
.A2(n_962),
.B1(n_608),
.B2(n_640),
.Y(n_1494)
);

AOI21xp5_ASAP7_75t_L g1495 ( 
.A1(n_1416),
.A2(n_1170),
.B(n_1102),
.Y(n_1495)
);

OAI21xp5_ASAP7_75t_L g1496 ( 
.A1(n_1420),
.A2(n_1190),
.B(n_1184),
.Y(n_1496)
);

AOI22xp5_ASAP7_75t_L g1497 ( 
.A1(n_1376),
.A2(n_1332),
.B1(n_1411),
.B2(n_1344),
.Y(n_1497)
);

A2O1A1Ixp33_ASAP7_75t_SL g1498 ( 
.A1(n_1423),
.A2(n_1190),
.B(n_1071),
.C(n_1075),
.Y(n_1498)
);

BUFx12f_ASAP7_75t_L g1499 ( 
.A(n_1380),
.Y(n_1499)
);

AOI21xp5_ASAP7_75t_L g1500 ( 
.A1(n_1333),
.A2(n_1418),
.B(n_1354),
.Y(n_1500)
);

INVx1_ASAP7_75t_L g1501 ( 
.A(n_1319),
.Y(n_1501)
);

O2A1O1Ixp33_ASAP7_75t_L g1502 ( 
.A1(n_1405),
.A2(n_959),
.B(n_570),
.C(n_574),
.Y(n_1502)
);

AOI21xp5_ASAP7_75t_L g1503 ( 
.A1(n_1333),
.A2(n_1354),
.B(n_1341),
.Y(n_1503)
);

A2O1A1Ixp33_ASAP7_75t_L g1504 ( 
.A1(n_1421),
.A2(n_1072),
.B(n_1070),
.C(n_1003),
.Y(n_1504)
);

A2O1A1Ixp33_ASAP7_75t_L g1505 ( 
.A1(n_1341),
.A2(n_1003),
.B(n_871),
.C(n_574),
.Y(n_1505)
);

NAND2xp5_ASAP7_75t_L g1506 ( 
.A(n_1334),
.B(n_1190),
.Y(n_1506)
);

NAND2xp5_ASAP7_75t_L g1507 ( 
.A(n_1337),
.B(n_1109),
.Y(n_1507)
);

NAND2xp5_ASAP7_75t_L g1508 ( 
.A(n_1345),
.B(n_1109),
.Y(n_1508)
);

INVx1_ASAP7_75t_L g1509 ( 
.A(n_1326),
.Y(n_1509)
);

AOI22xp33_ASAP7_75t_L g1510 ( 
.A1(n_1372),
.A2(n_608),
.B1(n_640),
.B2(n_587),
.Y(n_1510)
);

INVx1_ASAP7_75t_L g1511 ( 
.A(n_1330),
.Y(n_1511)
);

INVx1_ASAP7_75t_L g1512 ( 
.A(n_1331),
.Y(n_1512)
);

NAND2xp5_ASAP7_75t_L g1513 ( 
.A(n_1409),
.B(n_1111),
.Y(n_1513)
);

AOI21xp5_ASAP7_75t_L g1514 ( 
.A1(n_1420),
.A2(n_1170),
.B(n_1102),
.Y(n_1514)
);

AOI21xp5_ASAP7_75t_L g1515 ( 
.A1(n_1407),
.A2(n_1102),
.B(n_1094),
.Y(n_1515)
);

INVxp67_ASAP7_75t_L g1516 ( 
.A(n_1332),
.Y(n_1516)
);

AOI21xp5_ASAP7_75t_L g1517 ( 
.A1(n_1407),
.A2(n_1104),
.B(n_720),
.Y(n_1517)
);

INVx2_ASAP7_75t_L g1518 ( 
.A(n_1349),
.Y(n_1518)
);

O2A1O1Ixp33_ASAP7_75t_L g1519 ( 
.A1(n_1332),
.A2(n_579),
.B(n_585),
.C(n_564),
.Y(n_1519)
);

NAND2xp5_ASAP7_75t_L g1520 ( 
.A(n_1340),
.B(n_1343),
.Y(n_1520)
);

A2O1A1Ixp33_ASAP7_75t_L g1521 ( 
.A1(n_1347),
.A2(n_579),
.B(n_590),
.C(n_585),
.Y(n_1521)
);

AOI21xp5_ASAP7_75t_L g1522 ( 
.A1(n_1412),
.A2(n_1104),
.B(n_726),
.Y(n_1522)
);

NAND2xp5_ASAP7_75t_L g1523 ( 
.A(n_1346),
.B(n_1111),
.Y(n_1523)
);

A2O1A1Ixp33_ASAP7_75t_L g1524 ( 
.A1(n_1350),
.A2(n_591),
.B(n_612),
.C(n_590),
.Y(n_1524)
);

INVx2_ASAP7_75t_L g1525 ( 
.A(n_1355),
.Y(n_1525)
);

NOR2xp33_ASAP7_75t_L g1526 ( 
.A(n_1396),
.B(n_904),
.Y(n_1526)
);

NOR2xp33_ASAP7_75t_L g1527 ( 
.A(n_1353),
.B(n_913),
.Y(n_1527)
);

NOR2xp33_ASAP7_75t_R g1528 ( 
.A(n_1348),
.B(n_717),
.Y(n_1528)
);

NAND2xp5_ASAP7_75t_L g1529 ( 
.A(n_1352),
.B(n_1348),
.Y(n_1529)
);

CKINVDCx20_ASAP7_75t_R g1530 ( 
.A(n_1385),
.Y(n_1530)
);

NOR2xp33_ASAP7_75t_L g1531 ( 
.A(n_1387),
.B(n_915),
.Y(n_1531)
);

AOI21xp5_ASAP7_75t_L g1532 ( 
.A1(n_1503),
.A2(n_1415),
.B(n_1412),
.Y(n_1532)
);

AOI21xp5_ASAP7_75t_L g1533 ( 
.A1(n_1500),
.A2(n_1449),
.B(n_1462),
.Y(n_1533)
);

AOI21xp5_ASAP7_75t_L g1534 ( 
.A1(n_1449),
.A2(n_1415),
.B(n_1377),
.Y(n_1534)
);

NAND2xp5_ASAP7_75t_L g1535 ( 
.A(n_1437),
.B(n_1387),
.Y(n_1535)
);

INVx6_ASAP7_75t_SL g1536 ( 
.A(n_1491),
.Y(n_1536)
);

INVx1_ASAP7_75t_L g1537 ( 
.A(n_1471),
.Y(n_1537)
);

OAI21x1_ASAP7_75t_L g1538 ( 
.A1(n_1461),
.A2(n_1377),
.B(n_1373),
.Y(n_1538)
);

INVx1_ASAP7_75t_L g1539 ( 
.A(n_1501),
.Y(n_1539)
);

AND2x2_ASAP7_75t_L g1540 ( 
.A(n_1458),
.B(n_577),
.Y(n_1540)
);

AOI21xp5_ASAP7_75t_L g1541 ( 
.A1(n_1463),
.A2(n_1382),
.B(n_1373),
.Y(n_1541)
);

AOI22xp5_ASAP7_75t_L g1542 ( 
.A1(n_1450),
.A2(n_1425),
.B1(n_1424),
.B2(n_747),
.Y(n_1542)
);

NAND2xp5_ASAP7_75t_L g1543 ( 
.A(n_1448),
.B(n_1363),
.Y(n_1543)
);

A2O1A1Ixp33_ASAP7_75t_L g1544 ( 
.A1(n_1444),
.A2(n_1398),
.B(n_1400),
.C(n_1403),
.Y(n_1544)
);

O2A1O1Ixp33_ASAP7_75t_L g1545 ( 
.A1(n_1477),
.A2(n_921),
.B(n_591),
.C(n_613),
.Y(n_1545)
);

AO31x2_ASAP7_75t_L g1546 ( 
.A1(n_1505),
.A2(n_1402),
.A3(n_1388),
.B(n_1413),
.Y(n_1546)
);

NAND2xp5_ASAP7_75t_L g1547 ( 
.A(n_1453),
.B(n_1369),
.Y(n_1547)
);

BUFx6f_ASAP7_75t_L g1548 ( 
.A(n_1433),
.Y(n_1548)
);

A2O1A1Ixp33_ASAP7_75t_L g1549 ( 
.A1(n_1476),
.A2(n_1392),
.B(n_1371),
.C(n_1422),
.Y(n_1549)
);

AO21x2_ASAP7_75t_L g1550 ( 
.A1(n_1496),
.A2(n_1383),
.B(n_1382),
.Y(n_1550)
);

AOI21xp5_ASAP7_75t_L g1551 ( 
.A1(n_1464),
.A2(n_1384),
.B(n_1383),
.Y(n_1551)
);

AOI21xp5_ASAP7_75t_L g1552 ( 
.A1(n_1465),
.A2(n_1390),
.B(n_1384),
.Y(n_1552)
);

OAI21x1_ASAP7_75t_L g1553 ( 
.A1(n_1514),
.A2(n_1390),
.B(n_1112),
.Y(n_1553)
);

NOR2xp33_ASAP7_75t_L g1554 ( 
.A(n_1475),
.B(n_1342),
.Y(n_1554)
);

NAND2xp5_ASAP7_75t_L g1555 ( 
.A(n_1460),
.B(n_1531),
.Y(n_1555)
);

NAND2xp5_ASAP7_75t_L g1556 ( 
.A(n_1470),
.B(n_1342),
.Y(n_1556)
);

BUFx2_ASAP7_75t_L g1557 ( 
.A(n_1445),
.Y(n_1557)
);

NOR2xp33_ASAP7_75t_L g1558 ( 
.A(n_1429),
.B(n_1466),
.Y(n_1558)
);

OAI21xp5_ASAP7_75t_L g1559 ( 
.A1(n_1521),
.A2(n_1306),
.B(n_1112),
.Y(n_1559)
);

INVx2_ASAP7_75t_L g1560 ( 
.A(n_1442),
.Y(n_1560)
);

NOR2xp33_ASAP7_75t_SL g1561 ( 
.A(n_1452),
.B(n_577),
.Y(n_1561)
);

OAI21xp5_ASAP7_75t_L g1562 ( 
.A1(n_1496),
.A2(n_1306),
.B(n_769),
.Y(n_1562)
);

AOI21xp5_ASAP7_75t_L g1563 ( 
.A1(n_1459),
.A2(n_794),
.B(n_793),
.Y(n_1563)
);

NAND2xp5_ASAP7_75t_L g1564 ( 
.A(n_1486),
.B(n_729),
.Y(n_1564)
);

OAI21xp5_ASAP7_75t_L g1565 ( 
.A1(n_1517),
.A2(n_1306),
.B(n_803),
.Y(n_1565)
);

O2A1O1Ixp33_ASAP7_75t_SL g1566 ( 
.A1(n_1524),
.A2(n_994),
.B(n_613),
.C(n_617),
.Y(n_1566)
);

INVx2_ASAP7_75t_L g1567 ( 
.A(n_1483),
.Y(n_1567)
);

AOI21xp5_ASAP7_75t_L g1568 ( 
.A1(n_1481),
.A2(n_804),
.B(n_802),
.Y(n_1568)
);

O2A1O1Ixp33_ASAP7_75t_SL g1569 ( 
.A1(n_1498),
.A2(n_617),
.B(n_622),
.C(n_612),
.Y(n_1569)
);

NOR2xp33_ASAP7_75t_L g1570 ( 
.A(n_1451),
.B(n_596),
.Y(n_1570)
);

INVx2_ASAP7_75t_SL g1571 ( 
.A(n_1479),
.Y(n_1571)
);

OAI21x1_ASAP7_75t_L g1572 ( 
.A1(n_1430),
.A2(n_646),
.B(n_641),
.Y(n_1572)
);

OAI22xp5_ASAP7_75t_L g1573 ( 
.A1(n_1497),
.A2(n_819),
.B1(n_821),
.B2(n_807),
.Y(n_1573)
);

AND3x2_ASAP7_75t_L g1574 ( 
.A(n_1452),
.B(n_1432),
.C(n_1526),
.Y(n_1574)
);

AO31x2_ASAP7_75t_L g1575 ( 
.A1(n_1504),
.A2(n_628),
.A3(n_629),
.B(n_622),
.Y(n_1575)
);

OAI21xp5_ASAP7_75t_L g1576 ( 
.A1(n_1522),
.A2(n_1306),
.B(n_844),
.Y(n_1576)
);

NOR2xp67_ASAP7_75t_L g1577 ( 
.A(n_1467),
.B(n_467),
.Y(n_1577)
);

AOI21xp5_ASAP7_75t_L g1578 ( 
.A1(n_1431),
.A2(n_846),
.B(n_828),
.Y(n_1578)
);

NOR2xp33_ASAP7_75t_L g1579 ( 
.A(n_1439),
.B(n_597),
.Y(n_1579)
);

NOR2xp33_ASAP7_75t_L g1580 ( 
.A(n_1439),
.B(n_598),
.Y(n_1580)
);

OAI21x1_ASAP7_75t_L g1581 ( 
.A1(n_1489),
.A2(n_647),
.B(n_646),
.Y(n_1581)
);

AOI21xp5_ASAP7_75t_L g1582 ( 
.A1(n_1507),
.A2(n_925),
.B(n_922),
.Y(n_1582)
);

AOI21xp5_ASAP7_75t_L g1583 ( 
.A1(n_1508),
.A2(n_941),
.B(n_934),
.Y(n_1583)
);

NAND2xp5_ASAP7_75t_L g1584 ( 
.A(n_1468),
.B(n_949),
.Y(n_1584)
);

OA21x2_ASAP7_75t_L g1585 ( 
.A1(n_1506),
.A2(n_629),
.B(n_628),
.Y(n_1585)
);

AOI21xp5_ASAP7_75t_SL g1586 ( 
.A1(n_1502),
.A2(n_1441),
.B(n_1520),
.Y(n_1586)
);

OAI21x1_ASAP7_75t_L g1587 ( 
.A1(n_1495),
.A2(n_712),
.B(n_647),
.Y(n_1587)
);

OAI21x1_ASAP7_75t_L g1588 ( 
.A1(n_1515),
.A2(n_721),
.B(n_712),
.Y(n_1588)
);

AO21x2_ASAP7_75t_L g1589 ( 
.A1(n_1529),
.A2(n_1523),
.B(n_1511),
.Y(n_1589)
);

A2O1A1Ixp33_ASAP7_75t_L g1590 ( 
.A1(n_1434),
.A2(n_639),
.B(n_642),
.C(n_632),
.Y(n_1590)
);

A2O1A1Ixp33_ASAP7_75t_L g1591 ( 
.A1(n_1438),
.A2(n_639),
.B(n_642),
.C(n_632),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1509),
.Y(n_1592)
);

BUFx6f_ASAP7_75t_L g1593 ( 
.A(n_1433),
.Y(n_1593)
);

AOI21xp5_ASAP7_75t_L g1594 ( 
.A1(n_1428),
.A2(n_965),
.B(n_951),
.Y(n_1594)
);

A2O1A1Ixp33_ASAP7_75t_L g1595 ( 
.A1(n_1456),
.A2(n_645),
.B(n_650),
.C(n_644),
.Y(n_1595)
);

BUFx3_ASAP7_75t_L g1596 ( 
.A(n_1485),
.Y(n_1596)
);

OAI21x1_ASAP7_75t_L g1597 ( 
.A1(n_1443),
.A2(n_742),
.B(n_721),
.Y(n_1597)
);

AOI21xp5_ASAP7_75t_L g1598 ( 
.A1(n_1428),
.A2(n_980),
.B(n_975),
.Y(n_1598)
);

AND2x2_ASAP7_75t_L g1599 ( 
.A(n_1478),
.B(n_577),
.Y(n_1599)
);

BUFx6f_ASAP7_75t_L g1600 ( 
.A(n_1433),
.Y(n_1600)
);

INVx1_ASAP7_75t_L g1601 ( 
.A(n_1512),
.Y(n_1601)
);

INVx2_ASAP7_75t_L g1602 ( 
.A(n_1518),
.Y(n_1602)
);

NAND2xp5_ASAP7_75t_L g1603 ( 
.A(n_1491),
.B(n_976),
.Y(n_1603)
);

AOI21xp5_ASAP7_75t_L g1604 ( 
.A1(n_1428),
.A2(n_1306),
.B(n_754),
.Y(n_1604)
);

NAND2xp5_ASAP7_75t_L g1605 ( 
.A(n_1513),
.B(n_1484),
.Y(n_1605)
);

BUFx2_ASAP7_75t_L g1606 ( 
.A(n_1516),
.Y(n_1606)
);

INVx3_ASAP7_75t_L g1607 ( 
.A(n_1446),
.Y(n_1607)
);

NAND2xp5_ASAP7_75t_L g1608 ( 
.A(n_1473),
.B(n_604),
.Y(n_1608)
);

OA22x2_ASAP7_75t_L g1609 ( 
.A1(n_1482),
.A2(n_606),
.B1(n_609),
.B2(n_607),
.Y(n_1609)
);

OAI21xp5_ASAP7_75t_L g1610 ( 
.A1(n_1440),
.A2(n_1436),
.B(n_1474),
.Y(n_1610)
);

OAI21xp5_ASAP7_75t_L g1611 ( 
.A1(n_1510),
.A2(n_645),
.B(n_644),
.Y(n_1611)
);

AOI21xp5_ASAP7_75t_L g1612 ( 
.A1(n_1428),
.A2(n_754),
.B(n_742),
.Y(n_1612)
);

AO22x2_ASAP7_75t_L g1613 ( 
.A1(n_1490),
.A2(n_650),
.B1(n_658),
.B2(n_653),
.Y(n_1613)
);

NOR2xp33_ASAP7_75t_L g1614 ( 
.A(n_1469),
.B(n_610),
.Y(n_1614)
);

INVx2_ASAP7_75t_L g1615 ( 
.A(n_1525),
.Y(n_1615)
);

OAI21x1_ASAP7_75t_L g1616 ( 
.A1(n_1447),
.A2(n_823),
.B(n_780),
.Y(n_1616)
);

AOI21xp5_ASAP7_75t_L g1617 ( 
.A1(n_1472),
.A2(n_823),
.B(n_780),
.Y(n_1617)
);

NAND3x1_ASAP7_75t_L g1618 ( 
.A(n_1527),
.B(n_655),
.C(n_653),
.Y(n_1618)
);

AND2x2_ASAP7_75t_L g1619 ( 
.A(n_1492),
.B(n_599),
.Y(n_1619)
);

NAND2xp5_ASAP7_75t_L g1620 ( 
.A(n_1454),
.B(n_614),
.Y(n_1620)
);

BUFx6f_ASAP7_75t_L g1621 ( 
.A(n_1446),
.Y(n_1621)
);

INVx2_ASAP7_75t_SL g1622 ( 
.A(n_1435),
.Y(n_1622)
);

AOI21xp5_ASAP7_75t_L g1623 ( 
.A1(n_1480),
.A2(n_893),
.B(n_859),
.Y(n_1623)
);

AOI21xp5_ASAP7_75t_L g1624 ( 
.A1(n_1493),
.A2(n_893),
.B(n_859),
.Y(n_1624)
);

INVx3_ASAP7_75t_L g1625 ( 
.A(n_1446),
.Y(n_1625)
);

AOI21xp5_ASAP7_75t_L g1626 ( 
.A1(n_1457),
.A2(n_932),
.B(n_923),
.Y(n_1626)
);

INVx6_ASAP7_75t_L g1627 ( 
.A(n_1499),
.Y(n_1627)
);

OAI21x1_ASAP7_75t_L g1628 ( 
.A1(n_1457),
.A2(n_932),
.B(n_923),
.Y(n_1628)
);

INVxp67_ASAP7_75t_SL g1629 ( 
.A(n_1519),
.Y(n_1629)
);

INVx2_ASAP7_75t_L g1630 ( 
.A(n_1488),
.Y(n_1630)
);

NOR2xp33_ASAP7_75t_L g1631 ( 
.A(n_1487),
.B(n_615),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_1455),
.Y(n_1632)
);

INVx1_ASAP7_75t_L g1633 ( 
.A(n_1494),
.Y(n_1633)
);

OAI21x1_ASAP7_75t_L g1634 ( 
.A1(n_1528),
.A2(n_985),
.B(n_968),
.Y(n_1634)
);

OAI21x1_ASAP7_75t_L g1635 ( 
.A1(n_1530),
.A2(n_985),
.B(n_968),
.Y(n_1635)
);

OAI22x1_ASAP7_75t_L g1636 ( 
.A1(n_1450),
.A2(n_690),
.B1(n_713),
.B2(n_677),
.Y(n_1636)
);

A2O1A1Ixp33_ASAP7_75t_L g1637 ( 
.A1(n_1450),
.A2(n_658),
.B(n_663),
.C(n_655),
.Y(n_1637)
);

NAND2xp5_ASAP7_75t_L g1638 ( 
.A(n_1437),
.B(n_616),
.Y(n_1638)
);

NAND2xp5_ASAP7_75t_L g1639 ( 
.A(n_1437),
.B(n_620),
.Y(n_1639)
);

AO32x2_ASAP7_75t_L g1640 ( 
.A1(n_1482),
.A2(n_668),
.A3(n_670),
.B1(n_669),
.B2(n_663),
.Y(n_1640)
);

AND2x4_ASAP7_75t_L g1641 ( 
.A(n_1571),
.B(n_668),
.Y(n_1641)
);

NAND2x1p5_ASAP7_75t_L g1642 ( 
.A(n_1592),
.B(n_669),
.Y(n_1642)
);

INVx2_ASAP7_75t_L g1643 ( 
.A(n_1560),
.Y(n_1643)
);

OAI21x1_ASAP7_75t_L g1644 ( 
.A1(n_1553),
.A2(n_677),
.B(n_674),
.Y(n_1644)
);

INVx1_ASAP7_75t_L g1645 ( 
.A(n_1592),
.Y(n_1645)
);

INVx1_ASAP7_75t_L g1646 ( 
.A(n_1601),
.Y(n_1646)
);

OAI21x1_ASAP7_75t_L g1647 ( 
.A1(n_1538),
.A2(n_687),
.B(n_680),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_1601),
.Y(n_1648)
);

AOI22xp5_ASAP7_75t_L g1649 ( 
.A1(n_1558),
.A2(n_626),
.B1(n_627),
.B2(n_623),
.Y(n_1649)
);

OAI21x1_ASAP7_75t_L g1650 ( 
.A1(n_1532),
.A2(n_687),
.B(n_680),
.Y(n_1650)
);

NOR2xp33_ASAP7_75t_L g1651 ( 
.A(n_1555),
.B(n_633),
.Y(n_1651)
);

NAND2xp5_ASAP7_75t_L g1652 ( 
.A(n_1535),
.B(n_690),
.Y(n_1652)
);

AND2x2_ASAP7_75t_L g1653 ( 
.A(n_1554),
.B(n_1540),
.Y(n_1653)
);

NOR2x1_ASAP7_75t_SL g1654 ( 
.A(n_1589),
.B(n_587),
.Y(n_1654)
);

AOI222xp33_ASAP7_75t_L g1655 ( 
.A1(n_1579),
.A2(n_733),
.B1(n_713),
.B2(n_740),
.C1(n_725),
.C2(n_694),
.Y(n_1655)
);

INVx3_ASAP7_75t_L g1656 ( 
.A(n_1548),
.Y(n_1656)
);

OAI21x1_ASAP7_75t_L g1657 ( 
.A1(n_1572),
.A2(n_740),
.B(n_733),
.Y(n_1657)
);

HB1xp67_ASAP7_75t_L g1658 ( 
.A(n_1589),
.Y(n_1658)
);

OR2x6_ASAP7_75t_L g1659 ( 
.A(n_1586),
.B(n_762),
.Y(n_1659)
);

AND2x6_ASAP7_75t_L g1660 ( 
.A(n_1632),
.B(n_762),
.Y(n_1660)
);

OAI22xp5_ASAP7_75t_L g1661 ( 
.A1(n_1580),
.A2(n_764),
.B1(n_767),
.B2(n_763),
.Y(n_1661)
);

AOI22xp33_ASAP7_75t_SL g1662 ( 
.A1(n_1561),
.A2(n_599),
.B1(n_837),
.B2(n_722),
.Y(n_1662)
);

HB1xp67_ASAP7_75t_L g1663 ( 
.A(n_1546),
.Y(n_1663)
);

OAI21x1_ASAP7_75t_L g1664 ( 
.A1(n_1628),
.A2(n_764),
.B(n_763),
.Y(n_1664)
);

AO31x2_ASAP7_75t_L g1665 ( 
.A1(n_1533),
.A2(n_997),
.A3(n_1002),
.B(n_996),
.Y(n_1665)
);

NOR2xp33_ASAP7_75t_L g1666 ( 
.A(n_1614),
.B(n_634),
.Y(n_1666)
);

OAI21x1_ASAP7_75t_L g1667 ( 
.A1(n_1581),
.A2(n_768),
.B(n_767),
.Y(n_1667)
);

INVx1_ASAP7_75t_SL g1668 ( 
.A(n_1606),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_1537),
.Y(n_1669)
);

AND2x2_ASAP7_75t_L g1670 ( 
.A(n_1613),
.B(n_599),
.Y(n_1670)
);

OAI21x1_ASAP7_75t_L g1671 ( 
.A1(n_1587),
.A2(n_781),
.B(n_768),
.Y(n_1671)
);

INVx2_ASAP7_75t_L g1672 ( 
.A(n_1567),
.Y(n_1672)
);

AOI21xp5_ASAP7_75t_L g1673 ( 
.A1(n_1534),
.A2(n_1551),
.B(n_1541),
.Y(n_1673)
);

OAI21x1_ASAP7_75t_L g1674 ( 
.A1(n_1588),
.A2(n_1616),
.B(n_1597),
.Y(n_1674)
);

NAND2xp5_ASAP7_75t_L g1675 ( 
.A(n_1552),
.B(n_781),
.Y(n_1675)
);

NAND3xp33_ASAP7_75t_L g1676 ( 
.A(n_1570),
.B(n_643),
.C(n_635),
.Y(n_1676)
);

OAI21xp33_ASAP7_75t_SL g1677 ( 
.A1(n_1610),
.A2(n_783),
.B(n_782),
.Y(n_1677)
);

OAI22xp5_ASAP7_75t_L g1678 ( 
.A1(n_1629),
.A2(n_783),
.B1(n_785),
.B2(n_782),
.Y(n_1678)
);

INVx2_ASAP7_75t_L g1679 ( 
.A(n_1602),
.Y(n_1679)
);

INVx5_ASAP7_75t_L g1680 ( 
.A(n_1548),
.Y(n_1680)
);

AO21x2_ASAP7_75t_L g1681 ( 
.A1(n_1562),
.A2(n_787),
.B(n_785),
.Y(n_1681)
);

INVx3_ASAP7_75t_L g1682 ( 
.A(n_1548),
.Y(n_1682)
);

AO21x1_ASAP7_75t_L g1683 ( 
.A1(n_1573),
.A2(n_799),
.B(n_787),
.Y(n_1683)
);

NAND2xp5_ASAP7_75t_L g1684 ( 
.A(n_1539),
.B(n_799),
.Y(n_1684)
);

INVx2_ASAP7_75t_L g1685 ( 
.A(n_1615),
.Y(n_1685)
);

OAI21x1_ASAP7_75t_L g1686 ( 
.A1(n_1623),
.A2(n_815),
.B(n_814),
.Y(n_1686)
);

INVx1_ASAP7_75t_L g1687 ( 
.A(n_1543),
.Y(n_1687)
);

INVx1_ASAP7_75t_L g1688 ( 
.A(n_1547),
.Y(n_1688)
);

AO22x2_ASAP7_75t_L g1689 ( 
.A1(n_1632),
.A2(n_815),
.B1(n_816),
.B2(n_814),
.Y(n_1689)
);

A2O1A1Ixp33_ASAP7_75t_L g1690 ( 
.A1(n_1630),
.A2(n_829),
.B(n_832),
.C(n_816),
.Y(n_1690)
);

OAI21x1_ASAP7_75t_L g1691 ( 
.A1(n_1634),
.A2(n_832),
.B(n_829),
.Y(n_1691)
);

INVx1_ASAP7_75t_L g1692 ( 
.A(n_1626),
.Y(n_1692)
);

CKINVDCx9p33_ASAP7_75t_R g1693 ( 
.A(n_1631),
.Y(n_1693)
);

INVx1_ASAP7_75t_L g1694 ( 
.A(n_1575),
.Y(n_1694)
);

NAND2xp5_ASAP7_75t_L g1695 ( 
.A(n_1556),
.B(n_839),
.Y(n_1695)
);

AND2x2_ASAP7_75t_L g1696 ( 
.A(n_1613),
.B(n_722),
.Y(n_1696)
);

INVx2_ASAP7_75t_L g1697 ( 
.A(n_1546),
.Y(n_1697)
);

OAI21xp5_ASAP7_75t_L g1698 ( 
.A1(n_1549),
.A2(n_841),
.B(n_839),
.Y(n_1698)
);

OAI21x1_ASAP7_75t_L g1699 ( 
.A1(n_1565),
.A2(n_842),
.B(n_841),
.Y(n_1699)
);

AND2x2_ASAP7_75t_L g1700 ( 
.A(n_1636),
.B(n_989),
.Y(n_1700)
);

O2A1O1Ixp33_ASAP7_75t_L g1701 ( 
.A1(n_1545),
.A2(n_845),
.B(n_854),
.C(n_842),
.Y(n_1701)
);

CKINVDCx20_ASAP7_75t_R g1702 ( 
.A(n_1557),
.Y(n_1702)
);

NAND2xp5_ASAP7_75t_L g1703 ( 
.A(n_1605),
.B(n_845),
.Y(n_1703)
);

BUFx2_ASAP7_75t_L g1704 ( 
.A(n_1536),
.Y(n_1704)
);

NAND2xp5_ASAP7_75t_L g1705 ( 
.A(n_1550),
.B(n_854),
.Y(n_1705)
);

O2A1O1Ixp33_ASAP7_75t_L g1706 ( 
.A1(n_1637),
.A2(n_861),
.B(n_862),
.C(n_860),
.Y(n_1706)
);

AOI22xp33_ASAP7_75t_L g1707 ( 
.A1(n_1609),
.A2(n_837),
.B1(n_989),
.B2(n_722),
.Y(n_1707)
);

AO21x1_ASAP7_75t_L g1708 ( 
.A1(n_1620),
.A2(n_861),
.B(n_860),
.Y(n_1708)
);

INVx2_ASAP7_75t_L g1709 ( 
.A(n_1546),
.Y(n_1709)
);

NOR2xp33_ASAP7_75t_L g1710 ( 
.A(n_1574),
.B(n_648),
.Y(n_1710)
);

INVxp67_ASAP7_75t_SL g1711 ( 
.A(n_1585),
.Y(n_1711)
);

INVx2_ASAP7_75t_L g1712 ( 
.A(n_1585),
.Y(n_1712)
);

O2A1O1Ixp33_ASAP7_75t_L g1713 ( 
.A1(n_1595),
.A2(n_869),
.B(n_875),
.C(n_862),
.Y(n_1713)
);

INVx1_ASAP7_75t_L g1714 ( 
.A(n_1575),
.Y(n_1714)
);

AOI221xp5_ASAP7_75t_L g1715 ( 
.A1(n_1608),
.A2(n_891),
.B1(n_901),
.B2(n_875),
.C(n_869),
.Y(n_1715)
);

AO21x2_ASAP7_75t_L g1716 ( 
.A1(n_1576),
.A2(n_901),
.B(n_891),
.Y(n_1716)
);

INVx2_ASAP7_75t_L g1717 ( 
.A(n_1607),
.Y(n_1717)
);

OAI22xp33_ASAP7_75t_L g1718 ( 
.A1(n_1638),
.A2(n_908),
.B1(n_912),
.B2(n_903),
.Y(n_1718)
);

OAI21x1_ASAP7_75t_L g1719 ( 
.A1(n_1604),
.A2(n_1612),
.B(n_1624),
.Y(n_1719)
);

OAI21x1_ASAP7_75t_L g1720 ( 
.A1(n_1559),
.A2(n_908),
.B(n_903),
.Y(n_1720)
);

OAI21x1_ASAP7_75t_L g1721 ( 
.A1(n_1617),
.A2(n_918),
.B(n_912),
.Y(n_1721)
);

AOI21xp33_ASAP7_75t_L g1722 ( 
.A1(n_1564),
.A2(n_929),
.B(n_918),
.Y(n_1722)
);

OAI21x1_ASAP7_75t_L g1723 ( 
.A1(n_1578),
.A2(n_942),
.B(n_929),
.Y(n_1723)
);

AND2x2_ASAP7_75t_L g1724 ( 
.A(n_1635),
.B(n_1599),
.Y(n_1724)
);

OAI21x1_ASAP7_75t_SL g1725 ( 
.A1(n_1633),
.A2(n_1002),
.B(n_943),
.Y(n_1725)
);

BUFx2_ASAP7_75t_SL g1726 ( 
.A(n_1593),
.Y(n_1726)
);

INVx1_ASAP7_75t_L g1727 ( 
.A(n_1575),
.Y(n_1727)
);

AND2x4_ASAP7_75t_L g1728 ( 
.A(n_1607),
.B(n_942),
.Y(n_1728)
);

OAI21x1_ASAP7_75t_L g1729 ( 
.A1(n_1563),
.A2(n_945),
.B(n_943),
.Y(n_1729)
);

AOI22xp33_ASAP7_75t_L g1730 ( 
.A1(n_1619),
.A2(n_840),
.B1(n_874),
.B2(n_837),
.Y(n_1730)
);

CKINVDCx11_ASAP7_75t_R g1731 ( 
.A(n_1596),
.Y(n_1731)
);

AND2x2_ASAP7_75t_L g1732 ( 
.A(n_1653),
.B(n_1640),
.Y(n_1732)
);

NAND2xp5_ASAP7_75t_L g1733 ( 
.A(n_1687),
.B(n_1639),
.Y(n_1733)
);

OR2x2_ASAP7_75t_L g1734 ( 
.A(n_1705),
.B(n_1622),
.Y(n_1734)
);

AND2x2_ASAP7_75t_L g1735 ( 
.A(n_1728),
.B(n_1640),
.Y(n_1735)
);

OA21x2_ASAP7_75t_L g1736 ( 
.A1(n_1673),
.A2(n_1633),
.B(n_1590),
.Y(n_1736)
);

INVx1_ASAP7_75t_L g1737 ( 
.A(n_1645),
.Y(n_1737)
);

OAI22xp5_ASAP7_75t_L g1738 ( 
.A1(n_1666),
.A2(n_1618),
.B1(n_1603),
.B2(n_1542),
.Y(n_1738)
);

OAI22xp5_ASAP7_75t_L g1739 ( 
.A1(n_1662),
.A2(n_1584),
.B1(n_1591),
.B2(n_1536),
.Y(n_1739)
);

NAND2xp5_ASAP7_75t_L g1740 ( 
.A(n_1688),
.B(n_1625),
.Y(n_1740)
);

CKINVDCx5p33_ASAP7_75t_R g1741 ( 
.A(n_1731),
.Y(n_1741)
);

INVxp67_ASAP7_75t_L g1742 ( 
.A(n_1668),
.Y(n_1742)
);

AND2x2_ASAP7_75t_L g1743 ( 
.A(n_1646),
.B(n_1640),
.Y(n_1743)
);

AOI21x1_ASAP7_75t_SL g1744 ( 
.A1(n_1675),
.A2(n_1569),
.B(n_1627),
.Y(n_1744)
);

CKINVDCx20_ASAP7_75t_R g1745 ( 
.A(n_1702),
.Y(n_1745)
);

A2O1A1Ixp33_ASAP7_75t_L g1746 ( 
.A1(n_1722),
.A2(n_1611),
.B(n_1577),
.C(n_1544),
.Y(n_1746)
);

AND2x2_ASAP7_75t_L g1747 ( 
.A(n_1648),
.B(n_1550),
.Y(n_1747)
);

OR2x6_ASAP7_75t_L g1748 ( 
.A(n_1659),
.B(n_1627),
.Y(n_1748)
);

AND2x2_ASAP7_75t_L g1749 ( 
.A(n_1694),
.B(n_1625),
.Y(n_1749)
);

CKINVDCx6p67_ASAP7_75t_R g1750 ( 
.A(n_1680),
.Y(n_1750)
);

AND2x2_ASAP7_75t_L g1751 ( 
.A(n_1714),
.B(n_1593),
.Y(n_1751)
);

AOI21x1_ASAP7_75t_SL g1752 ( 
.A1(n_1675),
.A2(n_1566),
.B(n_1582),
.Y(n_1752)
);

INVx2_ASAP7_75t_L g1753 ( 
.A(n_1697),
.Y(n_1753)
);

BUFx6f_ASAP7_75t_L g1754 ( 
.A(n_1680),
.Y(n_1754)
);

INVx1_ASAP7_75t_L g1755 ( 
.A(n_1669),
.Y(n_1755)
);

AOI21xp5_ASAP7_75t_SL g1756 ( 
.A1(n_1659),
.A2(n_1583),
.B(n_1568),
.Y(n_1756)
);

BUFx4f_ASAP7_75t_L g1757 ( 
.A(n_1660),
.Y(n_1757)
);

CKINVDCx20_ASAP7_75t_R g1758 ( 
.A(n_1693),
.Y(n_1758)
);

OA21x2_ASAP7_75t_L g1759 ( 
.A1(n_1673),
.A2(n_946),
.B(n_945),
.Y(n_1759)
);

AOI21xp5_ASAP7_75t_L g1760 ( 
.A1(n_1659),
.A2(n_1598),
.B(n_1594),
.Y(n_1760)
);

O2A1O1Ixp5_ASAP7_75t_L g1761 ( 
.A1(n_1683),
.A2(n_948),
.B(n_952),
.C(n_946),
.Y(n_1761)
);

INVx1_ASAP7_75t_L g1762 ( 
.A(n_1705),
.Y(n_1762)
);

AOI21xp5_ASAP7_75t_SL g1763 ( 
.A1(n_1710),
.A2(n_1600),
.B(n_1593),
.Y(n_1763)
);

AOI221x1_ASAP7_75t_SL g1764 ( 
.A1(n_1661),
.A2(n_994),
.B1(n_992),
.B2(n_991),
.C(n_954),
.Y(n_1764)
);

O2A1O1Ixp5_ASAP7_75t_L g1765 ( 
.A1(n_1708),
.A2(n_1698),
.B(n_1722),
.C(n_1661),
.Y(n_1765)
);

AND2x4_ASAP7_75t_L g1766 ( 
.A(n_1643),
.B(n_1600),
.Y(n_1766)
);

AOI21xp5_ASAP7_75t_SL g1767 ( 
.A1(n_1701),
.A2(n_1621),
.B(n_1600),
.Y(n_1767)
);

AOI21xp5_ASAP7_75t_L g1768 ( 
.A1(n_1716),
.A2(n_1681),
.B(n_1658),
.Y(n_1768)
);

AND2x2_ASAP7_75t_L g1769 ( 
.A(n_1728),
.B(n_1621),
.Y(n_1769)
);

OR2x2_ASAP7_75t_L g1770 ( 
.A(n_1695),
.B(n_1621),
.Y(n_1770)
);

AND2x4_ASAP7_75t_L g1771 ( 
.A(n_1672),
.B(n_469),
.Y(n_1771)
);

O2A1O1Ixp5_ASAP7_75t_L g1772 ( 
.A1(n_1698),
.A2(n_952),
.B(n_954),
.C(n_948),
.Y(n_1772)
);

NAND2xp5_ASAP7_75t_L g1773 ( 
.A(n_1695),
.B(n_1651),
.Y(n_1773)
);

OA21x2_ASAP7_75t_L g1774 ( 
.A1(n_1644),
.A2(n_957),
.B(n_956),
.Y(n_1774)
);

INVx2_ASAP7_75t_L g1775 ( 
.A(n_1709),
.Y(n_1775)
);

INVx2_ASAP7_75t_L g1776 ( 
.A(n_1665),
.Y(n_1776)
);

OAI22xp5_ASAP7_75t_L g1777 ( 
.A1(n_1662),
.A2(n_1676),
.B1(n_1649),
.B2(n_1668),
.Y(n_1777)
);

AND2x2_ASAP7_75t_L g1778 ( 
.A(n_1727),
.B(n_956),
.Y(n_1778)
);

AOI21x1_ASAP7_75t_SL g1779 ( 
.A1(n_1670),
.A2(n_874),
.B(n_840),
.Y(n_1779)
);

AOI21xp5_ASAP7_75t_SL g1780 ( 
.A1(n_1701),
.A2(n_752),
.B(n_659),
.Y(n_1780)
);

INVx1_ASAP7_75t_L g1781 ( 
.A(n_1679),
.Y(n_1781)
);

AND2x2_ASAP7_75t_L g1782 ( 
.A(n_1689),
.B(n_957),
.Y(n_1782)
);

NAND2xp5_ASAP7_75t_L g1783 ( 
.A(n_1703),
.B(n_1004),
.Y(n_1783)
);

INVx3_ASAP7_75t_L g1784 ( 
.A(n_1665),
.Y(n_1784)
);

AOI21x1_ASAP7_75t_SL g1785 ( 
.A1(n_1696),
.A2(n_874),
.B(n_840),
.Y(n_1785)
);

OAI22xp5_ASAP7_75t_L g1786 ( 
.A1(n_1730),
.A2(n_652),
.B1(n_654),
.B2(n_651),
.Y(n_1786)
);

OA21x2_ASAP7_75t_L g1787 ( 
.A1(n_1647),
.A2(n_969),
.B(n_960),
.Y(n_1787)
);

OAI22xp5_ASAP7_75t_L g1788 ( 
.A1(n_1707),
.A2(n_660),
.B1(n_661),
.B2(n_656),
.Y(n_1788)
);

AND2x2_ASAP7_75t_L g1789 ( 
.A(n_1689),
.B(n_960),
.Y(n_1789)
);

AOI211xp5_ASAP7_75t_L g1790 ( 
.A1(n_1718),
.A2(n_1715),
.B(n_1677),
.C(n_1678),
.Y(n_1790)
);

BUFx3_ASAP7_75t_L g1791 ( 
.A(n_1704),
.Y(n_1791)
);

INVx5_ASAP7_75t_L g1792 ( 
.A(n_1660),
.Y(n_1792)
);

OA21x2_ASAP7_75t_L g1793 ( 
.A1(n_1711),
.A2(n_977),
.B(n_969),
.Y(n_1793)
);

INVx1_ASAP7_75t_L g1794 ( 
.A(n_1685),
.Y(n_1794)
);

AND2x2_ASAP7_75t_L g1795 ( 
.A(n_1642),
.B(n_991),
.Y(n_1795)
);

AND2x2_ASAP7_75t_L g1796 ( 
.A(n_1689),
.B(n_977),
.Y(n_1796)
);

AND2x2_ASAP7_75t_L g1797 ( 
.A(n_1663),
.B(n_979),
.Y(n_1797)
);

OR2x6_ASAP7_75t_L g1798 ( 
.A(n_1776),
.B(n_1663),
.Y(n_1798)
);

INVx1_ASAP7_75t_L g1799 ( 
.A(n_1753),
.Y(n_1799)
);

INVx2_ASAP7_75t_L g1800 ( 
.A(n_1776),
.Y(n_1800)
);

OAI21x1_ASAP7_75t_L g1801 ( 
.A1(n_1784),
.A2(n_1674),
.B(n_1671),
.Y(n_1801)
);

BUFx3_ASAP7_75t_L g1802 ( 
.A(n_1792),
.Y(n_1802)
);

INVx2_ASAP7_75t_L g1803 ( 
.A(n_1753),
.Y(n_1803)
);

OA21x2_ASAP7_75t_L g1804 ( 
.A1(n_1768),
.A2(n_1711),
.B(n_1712),
.Y(n_1804)
);

INVx2_ASAP7_75t_L g1805 ( 
.A(n_1775),
.Y(n_1805)
);

INVx2_ASAP7_75t_L g1806 ( 
.A(n_1775),
.Y(n_1806)
);

AND2x4_ASAP7_75t_L g1807 ( 
.A(n_1784),
.B(n_1747),
.Y(n_1807)
);

OA21x2_ASAP7_75t_L g1808 ( 
.A1(n_1762),
.A2(n_1658),
.B(n_1699),
.Y(n_1808)
);

NOR2xp33_ASAP7_75t_L g1809 ( 
.A(n_1773),
.B(n_1724),
.Y(n_1809)
);

BUFx2_ASAP7_75t_SL g1810 ( 
.A(n_1792),
.Y(n_1810)
);

BUFx3_ASAP7_75t_L g1811 ( 
.A(n_1792),
.Y(n_1811)
);

INVx1_ASAP7_75t_L g1812 ( 
.A(n_1737),
.Y(n_1812)
);

AND2x2_ASAP7_75t_L g1813 ( 
.A(n_1747),
.B(n_1665),
.Y(n_1813)
);

AND2x2_ASAP7_75t_L g1814 ( 
.A(n_1784),
.B(n_1654),
.Y(n_1814)
);

INVx1_ASAP7_75t_L g1815 ( 
.A(n_1755),
.Y(n_1815)
);

OR2x6_ASAP7_75t_L g1816 ( 
.A(n_1756),
.B(n_1719),
.Y(n_1816)
);

INVx1_ASAP7_75t_L g1817 ( 
.A(n_1759),
.Y(n_1817)
);

INVx4_ASAP7_75t_L g1818 ( 
.A(n_1792),
.Y(n_1818)
);

INVx1_ASAP7_75t_L g1819 ( 
.A(n_1759),
.Y(n_1819)
);

INVx1_ASAP7_75t_L g1820 ( 
.A(n_1759),
.Y(n_1820)
);

OAI21x1_ASAP7_75t_L g1821 ( 
.A1(n_1736),
.A2(n_1667),
.B(n_1650),
.Y(n_1821)
);

INVx2_ASAP7_75t_L g1822 ( 
.A(n_1778),
.Y(n_1822)
);

HB1xp67_ASAP7_75t_L g1823 ( 
.A(n_1749),
.Y(n_1823)
);

INVx2_ASAP7_75t_L g1824 ( 
.A(n_1778),
.Y(n_1824)
);

BUFx4f_ASAP7_75t_L g1825 ( 
.A(n_1750),
.Y(n_1825)
);

INVx2_ASAP7_75t_L g1826 ( 
.A(n_1749),
.Y(n_1826)
);

INVx2_ASAP7_75t_L g1827 ( 
.A(n_1736),
.Y(n_1827)
);

AO21x2_ASAP7_75t_L g1828 ( 
.A1(n_1746),
.A2(n_1716),
.B(n_1681),
.Y(n_1828)
);

BUFx6f_ASAP7_75t_L g1829 ( 
.A(n_1792),
.Y(n_1829)
);

OA21x2_ASAP7_75t_L g1830 ( 
.A1(n_1743),
.A2(n_1720),
.B(n_1691),
.Y(n_1830)
);

AND2x2_ASAP7_75t_L g1831 ( 
.A(n_1743),
.B(n_1692),
.Y(n_1831)
);

HB1xp67_ASAP7_75t_L g1832 ( 
.A(n_1797),
.Y(n_1832)
);

AND2x2_ASAP7_75t_L g1833 ( 
.A(n_1797),
.B(n_1660),
.Y(n_1833)
);

BUFx3_ASAP7_75t_L g1834 ( 
.A(n_1751),
.Y(n_1834)
);

HB1xp67_ASAP7_75t_L g1835 ( 
.A(n_1751),
.Y(n_1835)
);

INVx2_ASAP7_75t_L g1836 ( 
.A(n_1736),
.Y(n_1836)
);

HB1xp67_ASAP7_75t_L g1837 ( 
.A(n_1793),
.Y(n_1837)
);

INVx1_ASAP7_75t_L g1838 ( 
.A(n_1793),
.Y(n_1838)
);

AOI22xp5_ASAP7_75t_L g1839 ( 
.A1(n_1790),
.A2(n_1655),
.B1(n_1718),
.B2(n_1715),
.Y(n_1839)
);

AND2x2_ASAP7_75t_L g1840 ( 
.A(n_1732),
.B(n_1660),
.Y(n_1840)
);

INVx2_ASAP7_75t_L g1841 ( 
.A(n_1793),
.Y(n_1841)
);

INVx1_ASAP7_75t_L g1842 ( 
.A(n_1781),
.Y(n_1842)
);

INVx4_ASAP7_75t_L g1843 ( 
.A(n_1750),
.Y(n_1843)
);

INVx1_ASAP7_75t_L g1844 ( 
.A(n_1794),
.Y(n_1844)
);

AND2x2_ASAP7_75t_L g1845 ( 
.A(n_1782),
.B(n_1660),
.Y(n_1845)
);

BUFx2_ASAP7_75t_L g1846 ( 
.A(n_1742),
.Y(n_1846)
);

INVx2_ASAP7_75t_L g1847 ( 
.A(n_1774),
.Y(n_1847)
);

HB1xp67_ASAP7_75t_L g1848 ( 
.A(n_1770),
.Y(n_1848)
);

AND2x2_ASAP7_75t_L g1849 ( 
.A(n_1782),
.B(n_1723),
.Y(n_1849)
);

INVx1_ASAP7_75t_L g1850 ( 
.A(n_1815),
.Y(n_1850)
);

INVx1_ASAP7_75t_L g1851 ( 
.A(n_1815),
.Y(n_1851)
);

INVx1_ASAP7_75t_L g1852 ( 
.A(n_1815),
.Y(n_1852)
);

INVx1_ASAP7_75t_L g1853 ( 
.A(n_1812),
.Y(n_1853)
);

INVx2_ASAP7_75t_L g1854 ( 
.A(n_1800),
.Y(n_1854)
);

NAND2xp5_ASAP7_75t_L g1855 ( 
.A(n_1831),
.B(n_1842),
.Y(n_1855)
);

AND2x2_ASAP7_75t_L g1856 ( 
.A(n_1826),
.B(n_1796),
.Y(n_1856)
);

AND2x4_ASAP7_75t_L g1857 ( 
.A(n_1826),
.B(n_1789),
.Y(n_1857)
);

INVx1_ASAP7_75t_L g1858 ( 
.A(n_1812),
.Y(n_1858)
);

INVx1_ASAP7_75t_L g1859 ( 
.A(n_1799),
.Y(n_1859)
);

NOR2x1_ASAP7_75t_L g1860 ( 
.A(n_1810),
.B(n_1758),
.Y(n_1860)
);

INVx1_ASAP7_75t_L g1861 ( 
.A(n_1799),
.Y(n_1861)
);

NAND2xp5_ASAP7_75t_L g1862 ( 
.A(n_1831),
.B(n_1789),
.Y(n_1862)
);

AND2x2_ASAP7_75t_L g1863 ( 
.A(n_1826),
.B(n_1796),
.Y(n_1863)
);

INVx1_ASAP7_75t_L g1864 ( 
.A(n_1799),
.Y(n_1864)
);

INVx1_ASAP7_75t_L g1865 ( 
.A(n_1842),
.Y(n_1865)
);

BUFx2_ASAP7_75t_L g1866 ( 
.A(n_1807),
.Y(n_1866)
);

INVx1_ASAP7_75t_L g1867 ( 
.A(n_1842),
.Y(n_1867)
);

AND2x2_ASAP7_75t_L g1868 ( 
.A(n_1826),
.B(n_1735),
.Y(n_1868)
);

INVxp67_ASAP7_75t_SL g1869 ( 
.A(n_1837),
.Y(n_1869)
);

INVx2_ASAP7_75t_L g1870 ( 
.A(n_1800),
.Y(n_1870)
);

INVx1_ASAP7_75t_L g1871 ( 
.A(n_1803),
.Y(n_1871)
);

HB1xp67_ASAP7_75t_L g1872 ( 
.A(n_1848),
.Y(n_1872)
);

AND2x2_ASAP7_75t_L g1873 ( 
.A(n_1807),
.B(n_1774),
.Y(n_1873)
);

INVx2_ASAP7_75t_L g1874 ( 
.A(n_1800),
.Y(n_1874)
);

AND2x2_ASAP7_75t_L g1875 ( 
.A(n_1807),
.B(n_1774),
.Y(n_1875)
);

INVx1_ASAP7_75t_L g1876 ( 
.A(n_1803),
.Y(n_1876)
);

BUFx2_ASAP7_75t_L g1877 ( 
.A(n_1807),
.Y(n_1877)
);

INVx2_ASAP7_75t_L g1878 ( 
.A(n_1800),
.Y(n_1878)
);

HB1xp67_ASAP7_75t_L g1879 ( 
.A(n_1848),
.Y(n_1879)
);

NAND3xp33_ASAP7_75t_L g1880 ( 
.A(n_1839),
.B(n_1655),
.C(n_1777),
.Y(n_1880)
);

AND2x4_ASAP7_75t_L g1881 ( 
.A(n_1802),
.B(n_1811),
.Y(n_1881)
);

AND2x2_ASAP7_75t_L g1882 ( 
.A(n_1807),
.B(n_1787),
.Y(n_1882)
);

AND2x2_ASAP7_75t_L g1883 ( 
.A(n_1807),
.B(n_1787),
.Y(n_1883)
);

INVx2_ASAP7_75t_L g1884 ( 
.A(n_1803),
.Y(n_1884)
);

AND2x2_ASAP7_75t_L g1885 ( 
.A(n_1831),
.B(n_1787),
.Y(n_1885)
);

INVx1_ASAP7_75t_L g1886 ( 
.A(n_1803),
.Y(n_1886)
);

INVx2_ASAP7_75t_L g1887 ( 
.A(n_1805),
.Y(n_1887)
);

INVx2_ASAP7_75t_L g1888 ( 
.A(n_1805),
.Y(n_1888)
);

AND2x2_ASAP7_75t_L g1889 ( 
.A(n_1813),
.B(n_1757),
.Y(n_1889)
);

AND2x2_ASAP7_75t_L g1890 ( 
.A(n_1813),
.B(n_1757),
.Y(n_1890)
);

AND2x4_ASAP7_75t_L g1891 ( 
.A(n_1802),
.B(n_1766),
.Y(n_1891)
);

HB1xp67_ASAP7_75t_L g1892 ( 
.A(n_1832),
.Y(n_1892)
);

INVx1_ASAP7_75t_L g1893 ( 
.A(n_1805),
.Y(n_1893)
);

INVx1_ASAP7_75t_L g1894 ( 
.A(n_1805),
.Y(n_1894)
);

INVx2_ASAP7_75t_SL g1895 ( 
.A(n_1802),
.Y(n_1895)
);

INVx1_ASAP7_75t_L g1896 ( 
.A(n_1806),
.Y(n_1896)
);

AND2x2_ASAP7_75t_L g1897 ( 
.A(n_1813),
.B(n_1827),
.Y(n_1897)
);

BUFx2_ASAP7_75t_L g1898 ( 
.A(n_1832),
.Y(n_1898)
);

INVx11_ASAP7_75t_L g1899 ( 
.A(n_1825),
.Y(n_1899)
);

INVx2_ASAP7_75t_L g1900 ( 
.A(n_1806),
.Y(n_1900)
);

INVx1_ASAP7_75t_L g1901 ( 
.A(n_1806),
.Y(n_1901)
);

INVx3_ASAP7_75t_L g1902 ( 
.A(n_1818),
.Y(n_1902)
);

INVx2_ASAP7_75t_L g1903 ( 
.A(n_1806),
.Y(n_1903)
);

AND2x2_ASAP7_75t_L g1904 ( 
.A(n_1827),
.B(n_1757),
.Y(n_1904)
);

NAND2xp5_ASAP7_75t_L g1905 ( 
.A(n_1844),
.B(n_1733),
.Y(n_1905)
);

HB1xp67_ASAP7_75t_L g1906 ( 
.A(n_1872),
.Y(n_1906)
);

AND2x2_ASAP7_75t_L g1907 ( 
.A(n_1866),
.B(n_1835),
.Y(n_1907)
);

BUFx6f_ASAP7_75t_L g1908 ( 
.A(n_1902),
.Y(n_1908)
);

OAI211xp5_ASAP7_75t_L g1909 ( 
.A1(n_1880),
.A2(n_1839),
.B(n_1809),
.C(n_984),
.Y(n_1909)
);

INVx4_ASAP7_75t_L g1910 ( 
.A(n_1899),
.Y(n_1910)
);

INVx5_ASAP7_75t_SL g1911 ( 
.A(n_1899),
.Y(n_1911)
);

BUFx2_ASAP7_75t_L g1912 ( 
.A(n_1881),
.Y(n_1912)
);

AND2x4_ASAP7_75t_L g1913 ( 
.A(n_1866),
.B(n_1802),
.Y(n_1913)
);

OAI21x1_ASAP7_75t_L g1914 ( 
.A1(n_1902),
.A2(n_1836),
.B(n_1827),
.Y(n_1914)
);

AND2x2_ASAP7_75t_L g1915 ( 
.A(n_1877),
.B(n_1897),
.Y(n_1915)
);

OA21x2_ASAP7_75t_L g1916 ( 
.A1(n_1869),
.A2(n_1836),
.B(n_1827),
.Y(n_1916)
);

OAI321xp33_ASAP7_75t_L g1917 ( 
.A1(n_1880),
.A2(n_1738),
.A3(n_1809),
.B1(n_1678),
.B2(n_1746),
.C(n_1748),
.Y(n_1917)
);

INVx2_ASAP7_75t_L g1918 ( 
.A(n_1854),
.Y(n_1918)
);

INVx2_ASAP7_75t_L g1919 ( 
.A(n_1854),
.Y(n_1919)
);

AOI222xp33_ASAP7_75t_L g1920 ( 
.A1(n_1905),
.A2(n_1700),
.B1(n_1783),
.B2(n_984),
.C1(n_992),
.C2(n_979),
.Y(n_1920)
);

INVx2_ASAP7_75t_L g1921 ( 
.A(n_1854),
.Y(n_1921)
);

AND2x2_ASAP7_75t_L g1922 ( 
.A(n_1877),
.B(n_1835),
.Y(n_1922)
);

INVx1_ASAP7_75t_L g1923 ( 
.A(n_1850),
.Y(n_1923)
);

INVx2_ASAP7_75t_SL g1924 ( 
.A(n_1898),
.Y(n_1924)
);

OAI221xp5_ASAP7_75t_L g1925 ( 
.A1(n_1860),
.A2(n_1764),
.B1(n_1765),
.B2(n_1690),
.C(n_1734),
.Y(n_1925)
);

HB1xp67_ASAP7_75t_L g1926 ( 
.A(n_1879),
.Y(n_1926)
);

INVx1_ASAP7_75t_L g1927 ( 
.A(n_1850),
.Y(n_1927)
);

INVx1_ASAP7_75t_L g1928 ( 
.A(n_1851),
.Y(n_1928)
);

INVx1_ASAP7_75t_L g1929 ( 
.A(n_1851),
.Y(n_1929)
);

NOR2x1_ASAP7_75t_L g1930 ( 
.A(n_1860),
.B(n_1846),
.Y(n_1930)
);

INVx1_ASAP7_75t_L g1931 ( 
.A(n_1852),
.Y(n_1931)
);

INVx1_ASAP7_75t_L g1932 ( 
.A(n_1852),
.Y(n_1932)
);

OAI31xp33_ASAP7_75t_L g1933 ( 
.A1(n_1905),
.A2(n_1739),
.A3(n_1795),
.B(n_1845),
.Y(n_1933)
);

AOI22xp33_ASAP7_75t_L g1934 ( 
.A1(n_1889),
.A2(n_1845),
.B1(n_1849),
.B2(n_1828),
.Y(n_1934)
);

AND2x4_ASAP7_75t_L g1935 ( 
.A(n_1881),
.B(n_1811),
.Y(n_1935)
);

INVx1_ASAP7_75t_L g1936 ( 
.A(n_1859),
.Y(n_1936)
);

INVx2_ASAP7_75t_L g1937 ( 
.A(n_1870),
.Y(n_1937)
);

OAI211xp5_ASAP7_75t_L g1938 ( 
.A1(n_1862),
.A2(n_1780),
.B(n_1846),
.C(n_697),
.Y(n_1938)
);

INVx1_ASAP7_75t_L g1939 ( 
.A(n_1936),
.Y(n_1939)
);

INVxp67_ASAP7_75t_SL g1940 ( 
.A(n_1916),
.Y(n_1940)
);

INVx2_ASAP7_75t_L g1941 ( 
.A(n_1916),
.Y(n_1941)
);

INVx2_ASAP7_75t_L g1942 ( 
.A(n_1916),
.Y(n_1942)
);

INVx2_ASAP7_75t_L g1943 ( 
.A(n_1916),
.Y(n_1943)
);

INVx4_ASAP7_75t_SL g1944 ( 
.A(n_1908),
.Y(n_1944)
);

BUFx2_ASAP7_75t_SL g1945 ( 
.A(n_1924),
.Y(n_1945)
);

HB1xp67_ASAP7_75t_L g1946 ( 
.A(n_1936),
.Y(n_1946)
);

AOI21xp33_ASAP7_75t_SL g1947 ( 
.A1(n_1920),
.A2(n_1741),
.B(n_1693),
.Y(n_1947)
);

AND2x6_ASAP7_75t_SL g1948 ( 
.A(n_1935),
.B(n_1741),
.Y(n_1948)
);

INVx1_ASAP7_75t_L g1949 ( 
.A(n_1923),
.Y(n_1949)
);

AND2x2_ASAP7_75t_L g1950 ( 
.A(n_1912),
.B(n_1935),
.Y(n_1950)
);

HB1xp67_ASAP7_75t_L g1951 ( 
.A(n_1906),
.Y(n_1951)
);

BUFx2_ASAP7_75t_L g1952 ( 
.A(n_1930),
.Y(n_1952)
);

INVx3_ASAP7_75t_L g1953 ( 
.A(n_1908),
.Y(n_1953)
);

NOR2x1p5_ASAP7_75t_L g1954 ( 
.A(n_1910),
.B(n_1843),
.Y(n_1954)
);

INVx1_ASAP7_75t_L g1955 ( 
.A(n_1923),
.Y(n_1955)
);

INVx2_ASAP7_75t_L g1956 ( 
.A(n_1918),
.Y(n_1956)
);

OR2x6_ASAP7_75t_L g1957 ( 
.A(n_1930),
.B(n_1810),
.Y(n_1957)
);

INVx2_ASAP7_75t_L g1958 ( 
.A(n_1918),
.Y(n_1958)
);

BUFx3_ASAP7_75t_L g1959 ( 
.A(n_1908),
.Y(n_1959)
);

AND2x6_ASAP7_75t_L g1960 ( 
.A(n_1911),
.B(n_1829),
.Y(n_1960)
);

AND2x2_ASAP7_75t_L g1961 ( 
.A(n_1912),
.B(n_1897),
.Y(n_1961)
);

INVx3_ASAP7_75t_L g1962 ( 
.A(n_1908),
.Y(n_1962)
);

INVx2_ASAP7_75t_L g1963 ( 
.A(n_1918),
.Y(n_1963)
);

INVx1_ASAP7_75t_L g1964 ( 
.A(n_1927),
.Y(n_1964)
);

INVx2_ASAP7_75t_L g1965 ( 
.A(n_1919),
.Y(n_1965)
);

OA21x2_ASAP7_75t_L g1966 ( 
.A1(n_1914),
.A2(n_1869),
.B(n_1836),
.Y(n_1966)
);

INVx2_ASAP7_75t_L g1967 ( 
.A(n_1919),
.Y(n_1967)
);

INVx2_ASAP7_75t_L g1968 ( 
.A(n_1919),
.Y(n_1968)
);

INVx1_ASAP7_75t_SL g1969 ( 
.A(n_1926),
.Y(n_1969)
);

INVx1_ASAP7_75t_L g1970 ( 
.A(n_1927),
.Y(n_1970)
);

NAND2xp5_ASAP7_75t_L g1971 ( 
.A(n_1969),
.B(n_1933),
.Y(n_1971)
);

INVx2_ASAP7_75t_L g1972 ( 
.A(n_1956),
.Y(n_1972)
);

INVx4_ASAP7_75t_L g1973 ( 
.A(n_1948),
.Y(n_1973)
);

INVx2_ASAP7_75t_L g1974 ( 
.A(n_1956),
.Y(n_1974)
);

AND2x2_ASAP7_75t_L g1975 ( 
.A(n_1950),
.B(n_1935),
.Y(n_1975)
);

INVx1_ASAP7_75t_L g1976 ( 
.A(n_1946),
.Y(n_1976)
);

AND2x2_ASAP7_75t_L g1977 ( 
.A(n_1950),
.B(n_1935),
.Y(n_1977)
);

OR2x2_ASAP7_75t_L g1978 ( 
.A(n_1969),
.B(n_1862),
.Y(n_1978)
);

HB1xp67_ASAP7_75t_L g1979 ( 
.A(n_1946),
.Y(n_1979)
);

OR2x2_ASAP7_75t_L g1980 ( 
.A(n_1951),
.B(n_1892),
.Y(n_1980)
);

NOR2xp33_ASAP7_75t_L g1981 ( 
.A(n_1947),
.B(n_1909),
.Y(n_1981)
);

INVx6_ASAP7_75t_L g1982 ( 
.A(n_1948),
.Y(n_1982)
);

INVx4_ASAP7_75t_L g1983 ( 
.A(n_1944),
.Y(n_1983)
);

NAND2xp33_ASAP7_75t_SL g1984 ( 
.A(n_1954),
.B(n_1758),
.Y(n_1984)
);

INVx1_ASAP7_75t_SL g1985 ( 
.A(n_1945),
.Y(n_1985)
);

NAND2x1p5_ASAP7_75t_L g1986 ( 
.A(n_1952),
.B(n_1924),
.Y(n_1986)
);

INVx1_ASAP7_75t_SL g1987 ( 
.A(n_1945),
.Y(n_1987)
);

NAND2xp5_ASAP7_75t_L g1988 ( 
.A(n_1947),
.B(n_1933),
.Y(n_1988)
);

NAND2xp5_ASAP7_75t_L g1989 ( 
.A(n_1961),
.B(n_1846),
.Y(n_1989)
);

INVx4_ASAP7_75t_L g1990 ( 
.A(n_1960),
.Y(n_1990)
);

INVx1_ASAP7_75t_L g1991 ( 
.A(n_1939),
.Y(n_1991)
);

OR2x2_ASAP7_75t_L g1992 ( 
.A(n_1961),
.B(n_1898),
.Y(n_1992)
);

OR2x2_ASAP7_75t_L g1993 ( 
.A(n_1939),
.B(n_1855),
.Y(n_1993)
);

NAND2xp5_ASAP7_75t_L g1994 ( 
.A(n_1952),
.B(n_1907),
.Y(n_1994)
);

NOR2xp33_ASAP7_75t_L g1995 ( 
.A(n_1959),
.B(n_1917),
.Y(n_1995)
);

INVx5_ASAP7_75t_L g1996 ( 
.A(n_1960),
.Y(n_1996)
);

NAND3xp33_ASAP7_75t_SL g1997 ( 
.A(n_1941),
.B(n_1920),
.C(n_1938),
.Y(n_1997)
);

AND2x2_ASAP7_75t_L g1998 ( 
.A(n_1954),
.B(n_1913),
.Y(n_1998)
);

OR2x2_ASAP7_75t_L g1999 ( 
.A(n_1970),
.B(n_1855),
.Y(n_1999)
);

AND2x2_ASAP7_75t_L g2000 ( 
.A(n_1944),
.B(n_1913),
.Y(n_2000)
);

AND2x2_ASAP7_75t_L g2001 ( 
.A(n_1944),
.B(n_1913),
.Y(n_2001)
);

OR2x2_ASAP7_75t_L g2002 ( 
.A(n_1970),
.B(n_1857),
.Y(n_2002)
);

AND2x2_ASAP7_75t_L g2003 ( 
.A(n_1944),
.B(n_1913),
.Y(n_2003)
);

NOR2xp33_ASAP7_75t_L g2004 ( 
.A(n_1959),
.B(n_1917),
.Y(n_2004)
);

AND2x2_ASAP7_75t_L g2005 ( 
.A(n_2000),
.B(n_2001),
.Y(n_2005)
);

AND2x4_ASAP7_75t_L g2006 ( 
.A(n_1983),
.B(n_1944),
.Y(n_2006)
);

NAND2xp5_ASAP7_75t_L g2007 ( 
.A(n_1995),
.B(n_2004),
.Y(n_2007)
);

NAND2x1p5_ASAP7_75t_L g2008 ( 
.A(n_1996),
.B(n_1959),
.Y(n_2008)
);

OR2x2_ASAP7_75t_L g2009 ( 
.A(n_1971),
.B(n_1978),
.Y(n_2009)
);

AND2x2_ASAP7_75t_L g2010 ( 
.A(n_2003),
.B(n_1953),
.Y(n_2010)
);

INVx1_ASAP7_75t_L g2011 ( 
.A(n_1979),
.Y(n_2011)
);

AND2x2_ASAP7_75t_L g2012 ( 
.A(n_1990),
.B(n_1953),
.Y(n_2012)
);

INVxp67_ASAP7_75t_L g2013 ( 
.A(n_1981),
.Y(n_2013)
);

NAND2xp5_ASAP7_75t_L g2014 ( 
.A(n_1995),
.B(n_1949),
.Y(n_2014)
);

OR2x6_ASAP7_75t_L g2015 ( 
.A(n_1973),
.B(n_1957),
.Y(n_2015)
);

INVx1_ASAP7_75t_L g2016 ( 
.A(n_1979),
.Y(n_2016)
);

NOR2x1p5_ASAP7_75t_SL g2017 ( 
.A(n_1972),
.B(n_1956),
.Y(n_2017)
);

OR2x6_ASAP7_75t_L g2018 ( 
.A(n_1973),
.B(n_1957),
.Y(n_2018)
);

OAI21xp5_ASAP7_75t_L g2019 ( 
.A1(n_1997),
.A2(n_1957),
.B(n_1934),
.Y(n_2019)
);

NAND2xp5_ASAP7_75t_L g2020 ( 
.A(n_2004),
.B(n_1949),
.Y(n_2020)
);

AND2x2_ASAP7_75t_L g2021 ( 
.A(n_1990),
.B(n_1953),
.Y(n_2021)
);

AND2x2_ASAP7_75t_L g2022 ( 
.A(n_1990),
.B(n_1953),
.Y(n_2022)
);

AND2x2_ASAP7_75t_L g2023 ( 
.A(n_1975),
.B(n_1962),
.Y(n_2023)
);

NAND2xp5_ASAP7_75t_L g2024 ( 
.A(n_1988),
.B(n_1955),
.Y(n_2024)
);

INVx1_ASAP7_75t_L g2025 ( 
.A(n_1991),
.Y(n_2025)
);

AND2x2_ASAP7_75t_L g2026 ( 
.A(n_1977),
.B(n_1962),
.Y(n_2026)
);

NAND2xp5_ASAP7_75t_L g2027 ( 
.A(n_1981),
.B(n_1955),
.Y(n_2027)
);

INVx1_ASAP7_75t_L g2028 ( 
.A(n_1976),
.Y(n_2028)
);

OR2x2_ASAP7_75t_L g2029 ( 
.A(n_1997),
.B(n_1964),
.Y(n_2029)
);

INVxp67_ASAP7_75t_SL g2030 ( 
.A(n_1986),
.Y(n_2030)
);

AND2x2_ASAP7_75t_L g2031 ( 
.A(n_1985),
.B(n_1962),
.Y(n_2031)
);

INVx1_ASAP7_75t_L g2032 ( 
.A(n_1972),
.Y(n_2032)
);

INVx2_ASAP7_75t_L g2033 ( 
.A(n_1974),
.Y(n_2033)
);

INVx1_ASAP7_75t_L g2034 ( 
.A(n_1974),
.Y(n_2034)
);

AND2x2_ASAP7_75t_L g2035 ( 
.A(n_1987),
.B(n_1962),
.Y(n_2035)
);

INVx1_ASAP7_75t_L g2036 ( 
.A(n_1980),
.Y(n_2036)
);

INVx3_ASAP7_75t_SL g2037 ( 
.A(n_2006),
.Y(n_2037)
);

INVx1_ASAP7_75t_L g2038 ( 
.A(n_2011),
.Y(n_2038)
);

NAND2xp5_ASAP7_75t_L g2039 ( 
.A(n_2007),
.B(n_1982),
.Y(n_2039)
);

OAI21x1_ASAP7_75t_L g2040 ( 
.A1(n_2008),
.A2(n_1986),
.B(n_1994),
.Y(n_2040)
);

INVx2_ASAP7_75t_L g2041 ( 
.A(n_2005),
.Y(n_2041)
);

NAND2xp5_ASAP7_75t_L g2042 ( 
.A(n_2014),
.B(n_1982),
.Y(n_2042)
);

AND2x2_ASAP7_75t_L g2043 ( 
.A(n_2005),
.B(n_1998),
.Y(n_2043)
);

NOR2x1_ASAP7_75t_L g2044 ( 
.A(n_2006),
.B(n_1983),
.Y(n_2044)
);

AND2x2_ASAP7_75t_L g2045 ( 
.A(n_2031),
.B(n_1982),
.Y(n_2045)
);

INVx1_ASAP7_75t_L g2046 ( 
.A(n_2016),
.Y(n_2046)
);

INVx1_ASAP7_75t_L g2047 ( 
.A(n_2025),
.Y(n_2047)
);

INVx1_ASAP7_75t_L g2048 ( 
.A(n_2028),
.Y(n_2048)
);

NAND2xp5_ASAP7_75t_L g2049 ( 
.A(n_2020),
.B(n_1964),
.Y(n_2049)
);

OAI22xp5_ASAP7_75t_L g2050 ( 
.A1(n_2019),
.A2(n_1957),
.B1(n_1925),
.B2(n_1996),
.Y(n_2050)
);

OR2x2_ASAP7_75t_L g2051 ( 
.A(n_2009),
.B(n_1989),
.Y(n_2051)
);

INVxp67_ASAP7_75t_R g2052 ( 
.A(n_2031),
.Y(n_2052)
);

AND2x2_ASAP7_75t_L g2053 ( 
.A(n_2035),
.B(n_1996),
.Y(n_2053)
);

AND2x2_ASAP7_75t_L g2054 ( 
.A(n_2035),
.B(n_1996),
.Y(n_2054)
);

NOR2xp33_ASAP7_75t_L g2055 ( 
.A(n_2013),
.B(n_2027),
.Y(n_2055)
);

INVx1_ASAP7_75t_L g2056 ( 
.A(n_2033),
.Y(n_2056)
);

HB1xp67_ASAP7_75t_L g2057 ( 
.A(n_2029),
.Y(n_2057)
);

NAND3xp33_ASAP7_75t_L g2058 ( 
.A(n_2024),
.B(n_1984),
.C(n_1925),
.Y(n_2058)
);

INVx1_ASAP7_75t_L g2059 ( 
.A(n_2033),
.Y(n_2059)
);

OR2x2_ASAP7_75t_L g2060 ( 
.A(n_2036),
.B(n_1992),
.Y(n_2060)
);

INVx1_ASAP7_75t_L g2061 ( 
.A(n_2032),
.Y(n_2061)
);

AOI22xp33_ASAP7_75t_L g2062 ( 
.A1(n_2015),
.A2(n_1984),
.B1(n_1960),
.B2(n_1957),
.Y(n_2062)
);

NAND2xp5_ASAP7_75t_L g2063 ( 
.A(n_2034),
.B(n_1993),
.Y(n_2063)
);

INVx1_ASAP7_75t_L g2064 ( 
.A(n_2010),
.Y(n_2064)
);

INVx1_ASAP7_75t_L g2065 ( 
.A(n_2010),
.Y(n_2065)
);

INVx2_ASAP7_75t_L g2066 ( 
.A(n_2008),
.Y(n_2066)
);

INVx2_ASAP7_75t_L g2067 ( 
.A(n_2006),
.Y(n_2067)
);

OAI22xp5_ASAP7_75t_L g2068 ( 
.A1(n_2030),
.A2(n_1957),
.B1(n_1940),
.B2(n_1748),
.Y(n_2068)
);

INVx1_ASAP7_75t_SL g2069 ( 
.A(n_2012),
.Y(n_2069)
);

OR2x2_ASAP7_75t_L g2070 ( 
.A(n_2015),
.B(n_2002),
.Y(n_2070)
);

INVx1_ASAP7_75t_L g2071 ( 
.A(n_2017),
.Y(n_2071)
);

INVx1_ASAP7_75t_L g2072 ( 
.A(n_2023),
.Y(n_2072)
);

AND2x4_ASAP7_75t_L g2073 ( 
.A(n_2012),
.B(n_1960),
.Y(n_2073)
);

INVx2_ASAP7_75t_SL g2074 ( 
.A(n_2021),
.Y(n_2074)
);

OR2x2_ASAP7_75t_L g2075 ( 
.A(n_2015),
.B(n_1999),
.Y(n_2075)
);

BUFx3_ASAP7_75t_L g2076 ( 
.A(n_2021),
.Y(n_2076)
);

NAND2xp5_ASAP7_75t_SL g2077 ( 
.A(n_2022),
.B(n_1910),
.Y(n_2077)
);

INVx1_ASAP7_75t_SL g2078 ( 
.A(n_2022),
.Y(n_2078)
);

INVx1_ASAP7_75t_SL g2079 ( 
.A(n_2015),
.Y(n_2079)
);

AND3x1_ASAP7_75t_L g2080 ( 
.A(n_2023),
.B(n_2026),
.C(n_2018),
.Y(n_2080)
);

OR2x2_ASAP7_75t_L g2081 ( 
.A(n_2018),
.B(n_1958),
.Y(n_2081)
);

OAI21xp5_ASAP7_75t_L g2082 ( 
.A1(n_2050),
.A2(n_2018),
.B(n_2026),
.Y(n_2082)
);

AOI22xp5_ASAP7_75t_L g2083 ( 
.A1(n_2050),
.A2(n_2058),
.B1(n_2080),
.B2(n_2055),
.Y(n_2083)
);

OAI21xp5_ASAP7_75t_SL g2084 ( 
.A1(n_2039),
.A2(n_1788),
.B(n_1786),
.Y(n_2084)
);

INVx1_ASAP7_75t_L g2085 ( 
.A(n_2056),
.Y(n_2085)
);

OAI21xp33_ASAP7_75t_L g2086 ( 
.A1(n_2039),
.A2(n_2018),
.B(n_1940),
.Y(n_2086)
);

AND2x2_ASAP7_75t_SL g2087 ( 
.A(n_2057),
.B(n_1910),
.Y(n_2087)
);

OAI322xp33_ASAP7_75t_L g2088 ( 
.A1(n_2057),
.A2(n_734),
.A3(n_698),
.B1(n_751),
.B2(n_770),
.C1(n_710),
.C2(n_682),
.Y(n_2088)
);

OAI21xp33_ASAP7_75t_L g2089 ( 
.A1(n_2042),
.A2(n_1904),
.B(n_1890),
.Y(n_2089)
);

INVx1_ASAP7_75t_L g2090 ( 
.A(n_2059),
.Y(n_2090)
);

AOI322xp5_ASAP7_75t_L g2091 ( 
.A1(n_2042),
.A2(n_1942),
.A3(n_1941),
.B1(n_1943),
.B2(n_1915),
.C1(n_1922),
.C2(n_1907),
.Y(n_2091)
);

NAND2xp5_ASAP7_75t_L g2092 ( 
.A(n_2041),
.B(n_1922),
.Y(n_2092)
);

OAI211xp5_ASAP7_75t_SL g2093 ( 
.A1(n_2079),
.A2(n_1703),
.B(n_1942),
.C(n_1941),
.Y(n_2093)
);

NOR2xp33_ASAP7_75t_SL g2094 ( 
.A(n_2045),
.B(n_1910),
.Y(n_2094)
);

AOI22xp5_ASAP7_75t_L g2095 ( 
.A1(n_2043),
.A2(n_1960),
.B1(n_1881),
.B2(n_1904),
.Y(n_2095)
);

INVx1_ASAP7_75t_L g2096 ( 
.A(n_2061),
.Y(n_2096)
);

AOI22xp5_ASAP7_75t_L g2097 ( 
.A1(n_2052),
.A2(n_1960),
.B1(n_1881),
.B2(n_1904),
.Y(n_2097)
);

OAI322xp33_ASAP7_75t_L g2098 ( 
.A1(n_2038),
.A2(n_741),
.A3(n_700),
.B1(n_757),
.B2(n_791),
.C1(n_718),
.C2(n_684),
.Y(n_2098)
);

INVx1_ASAP7_75t_L g2099 ( 
.A(n_2046),
.Y(n_2099)
);

INVx2_ASAP7_75t_SL g2100 ( 
.A(n_2044),
.Y(n_2100)
);

OAI21xp33_ASAP7_75t_L g2101 ( 
.A1(n_2079),
.A2(n_1890),
.B(n_1889),
.Y(n_2101)
);

INVx1_ASAP7_75t_L g2102 ( 
.A(n_2047),
.Y(n_2102)
);

NOR2x1p5_ASAP7_75t_L g2103 ( 
.A(n_2067),
.B(n_1791),
.Y(n_2103)
);

NAND2xp5_ASAP7_75t_L g2104 ( 
.A(n_2069),
.B(n_2078),
.Y(n_2104)
);

AOI21xp33_ASAP7_75t_L g2105 ( 
.A1(n_2066),
.A2(n_1791),
.B(n_1828),
.Y(n_2105)
);

INVx1_ASAP7_75t_L g2106 ( 
.A(n_2064),
.Y(n_2106)
);

OAI21xp5_ASAP7_75t_L g2107 ( 
.A1(n_2040),
.A2(n_1960),
.B(n_1745),
.Y(n_2107)
);

NAND2xp5_ASAP7_75t_L g2108 ( 
.A(n_2069),
.B(n_1915),
.Y(n_2108)
);

NAND3xp33_ASAP7_75t_L g2109 ( 
.A(n_2074),
.B(n_608),
.C(n_587),
.Y(n_2109)
);

NAND2x1p5_ASAP7_75t_L g2110 ( 
.A(n_2053),
.B(n_1825),
.Y(n_2110)
);

NAND2xp5_ASAP7_75t_L g2111 ( 
.A(n_2078),
.B(n_1958),
.Y(n_2111)
);

NOR2xp33_ASAP7_75t_L g2112 ( 
.A(n_2037),
.B(n_1745),
.Y(n_2112)
);

AND2x2_ASAP7_75t_L g2113 ( 
.A(n_2076),
.B(n_1908),
.Y(n_2113)
);

OAI221xp5_ASAP7_75t_L g2114 ( 
.A1(n_2062),
.A2(n_1908),
.B1(n_1943),
.B2(n_1942),
.C(n_1895),
.Y(n_2114)
);

NOR2xp33_ASAP7_75t_L g2115 ( 
.A(n_2077),
.B(n_1641),
.Y(n_2115)
);

INVx1_ASAP7_75t_L g2116 ( 
.A(n_2065),
.Y(n_2116)
);

NAND3xp33_ASAP7_75t_L g2117 ( 
.A(n_2048),
.B(n_608),
.C(n_587),
.Y(n_2117)
);

AOI22xp33_ASAP7_75t_L g2118 ( 
.A1(n_2051),
.A2(n_1960),
.B1(n_1828),
.B2(n_1845),
.Y(n_2118)
);

NAND2xp5_ASAP7_75t_L g2119 ( 
.A(n_2072),
.B(n_1958),
.Y(n_2119)
);

INVx1_ASAP7_75t_L g2120 ( 
.A(n_2060),
.Y(n_2120)
);

AOI22xp5_ASAP7_75t_L g2121 ( 
.A1(n_2054),
.A2(n_1960),
.B1(n_1890),
.B2(n_1889),
.Y(n_2121)
);

HB1xp67_ASAP7_75t_L g2122 ( 
.A(n_2071),
.Y(n_2122)
);

AOI32xp33_ASAP7_75t_L g2123 ( 
.A1(n_2068),
.A2(n_1943),
.A3(n_1895),
.B1(n_1833),
.B2(n_1902),
.Y(n_2123)
);

AOI22xp5_ASAP7_75t_L g2124 ( 
.A1(n_2073),
.A2(n_1891),
.B1(n_1895),
.B2(n_1748),
.Y(n_2124)
);

NAND2xp5_ASAP7_75t_SL g2125 ( 
.A(n_2073),
.B(n_1911),
.Y(n_2125)
);

AOI22xp5_ASAP7_75t_L g2126 ( 
.A1(n_2068),
.A2(n_1891),
.B1(n_1748),
.B2(n_1902),
.Y(n_2126)
);

OR2x2_ASAP7_75t_L g2127 ( 
.A(n_2075),
.B(n_1968),
.Y(n_2127)
);

NAND3xp33_ASAP7_75t_L g2128 ( 
.A(n_2070),
.B(n_659),
.C(n_640),
.Y(n_2128)
);

AOI22xp5_ASAP7_75t_L g2129 ( 
.A1(n_2049),
.A2(n_1891),
.B1(n_1875),
.B2(n_1882),
.Y(n_2129)
);

OAI21xp5_ASAP7_75t_L g2130 ( 
.A1(n_2049),
.A2(n_2081),
.B(n_2063),
.Y(n_2130)
);

NOR2xp33_ASAP7_75t_L g2131 ( 
.A(n_2063),
.B(n_1641),
.Y(n_2131)
);

AND2x2_ASAP7_75t_L g2132 ( 
.A(n_2052),
.B(n_1963),
.Y(n_2132)
);

INVx1_ASAP7_75t_L g2133 ( 
.A(n_2056),
.Y(n_2133)
);

O2A1O1Ixp5_ASAP7_75t_L g2134 ( 
.A1(n_2050),
.A2(n_1965),
.B(n_1967),
.C(n_1963),
.Y(n_2134)
);

INVx2_ASAP7_75t_L g2135 ( 
.A(n_2076),
.Y(n_2135)
);

NOR2x1_ASAP7_75t_R g2136 ( 
.A(n_2039),
.B(n_691),
.Y(n_2136)
);

NOR3xp33_ASAP7_75t_L g2137 ( 
.A(n_2039),
.B(n_1652),
.C(n_1684),
.Y(n_2137)
);

AOI221xp5_ASAP7_75t_L g2138 ( 
.A1(n_2057),
.A2(n_672),
.B1(n_685),
.B2(n_681),
.C(n_675),
.Y(n_2138)
);

NAND2xp33_ASAP7_75t_L g2139 ( 
.A(n_2057),
.B(n_1829),
.Y(n_2139)
);

OAI21xp5_ASAP7_75t_L g2140 ( 
.A1(n_2050),
.A2(n_1761),
.B(n_1772),
.Y(n_2140)
);

INVx1_ASAP7_75t_L g2141 ( 
.A(n_2056),
.Y(n_2141)
);

AND3x1_ASAP7_75t_L g2142 ( 
.A(n_2055),
.B(n_1785),
.C(n_1779),
.Y(n_2142)
);

A2O1A1Ixp33_ASAP7_75t_L g2143 ( 
.A1(n_2058),
.A2(n_692),
.B(n_693),
.C(n_688),
.Y(n_2143)
);

INVx1_ASAP7_75t_L g2144 ( 
.A(n_2056),
.Y(n_2144)
);

NAND2xp5_ASAP7_75t_L g2145 ( 
.A(n_2041),
.B(n_1963),
.Y(n_2145)
);

INVx2_ASAP7_75t_L g2146 ( 
.A(n_2076),
.Y(n_2146)
);

NAND2xp5_ASAP7_75t_L g2147 ( 
.A(n_2122),
.B(n_2120),
.Y(n_2147)
);

INVx1_ASAP7_75t_SL g2148 ( 
.A(n_2087),
.Y(n_2148)
);

INVx1_ASAP7_75t_L g2149 ( 
.A(n_2104),
.Y(n_2149)
);

OR2x2_ASAP7_75t_L g2150 ( 
.A(n_2135),
.B(n_1967),
.Y(n_2150)
);

NAND2xp5_ASAP7_75t_L g2151 ( 
.A(n_2146),
.B(n_1965),
.Y(n_2151)
);

INVx2_ASAP7_75t_L g2152 ( 
.A(n_2100),
.Y(n_2152)
);

AND2x2_ASAP7_75t_L g2153 ( 
.A(n_2112),
.B(n_1965),
.Y(n_2153)
);

INVx2_ASAP7_75t_SL g2154 ( 
.A(n_2103),
.Y(n_2154)
);

INVx1_ASAP7_75t_L g2155 ( 
.A(n_2106),
.Y(n_2155)
);

OR2x2_ASAP7_75t_L g2156 ( 
.A(n_2116),
.B(n_1967),
.Y(n_2156)
);

BUFx2_ASAP7_75t_L g2157 ( 
.A(n_2136),
.Y(n_2157)
);

AND2x2_ASAP7_75t_L g2158 ( 
.A(n_2082),
.B(n_1968),
.Y(n_2158)
);

INVx1_ASAP7_75t_L g2159 ( 
.A(n_2085),
.Y(n_2159)
);

INVx2_ASAP7_75t_L g2160 ( 
.A(n_2110),
.Y(n_2160)
);

INVxp67_ASAP7_75t_L g2161 ( 
.A(n_2094),
.Y(n_2161)
);

NAND2xp5_ASAP7_75t_L g2162 ( 
.A(n_2083),
.B(n_1968),
.Y(n_2162)
);

INVx1_ASAP7_75t_SL g2163 ( 
.A(n_2139),
.Y(n_2163)
);

NAND2xp5_ASAP7_75t_SL g2164 ( 
.A(n_2107),
.B(n_1911),
.Y(n_2164)
);

AND2x2_ASAP7_75t_L g2165 ( 
.A(n_2131),
.B(n_1891),
.Y(n_2165)
);

INVx1_ASAP7_75t_L g2166 ( 
.A(n_2090),
.Y(n_2166)
);

AND2x2_ASAP7_75t_L g2167 ( 
.A(n_2115),
.B(n_1911),
.Y(n_2167)
);

OR2x2_ASAP7_75t_L g2168 ( 
.A(n_2092),
.B(n_1928),
.Y(n_2168)
);

NAND2xp5_ASAP7_75t_L g2169 ( 
.A(n_2143),
.B(n_1928),
.Y(n_2169)
);

OR2x2_ASAP7_75t_L g2170 ( 
.A(n_2108),
.B(n_1929),
.Y(n_2170)
);

OR2x2_ASAP7_75t_L g2171 ( 
.A(n_2130),
.B(n_1929),
.Y(n_2171)
);

AND2x2_ASAP7_75t_L g2172 ( 
.A(n_2113),
.B(n_1911),
.Y(n_2172)
);

NAND2xp5_ASAP7_75t_L g2173 ( 
.A(n_2137),
.B(n_1931),
.Y(n_2173)
);

AOI22xp33_ASAP7_75t_L g2174 ( 
.A1(n_2101),
.A2(n_1828),
.B1(n_1829),
.B2(n_1811),
.Y(n_2174)
);

NOR2xp33_ASAP7_75t_L g2175 ( 
.A(n_2088),
.B(n_696),
.Y(n_2175)
);

INVxp67_ASAP7_75t_L g2176 ( 
.A(n_2142),
.Y(n_2176)
);

NAND2xp5_ASAP7_75t_L g2177 ( 
.A(n_2138),
.B(n_1932),
.Y(n_2177)
);

AND2x2_ASAP7_75t_L g2178 ( 
.A(n_2125),
.B(n_1856),
.Y(n_2178)
);

AOI22xp33_ASAP7_75t_SL g2179 ( 
.A1(n_2114),
.A2(n_1829),
.B1(n_1966),
.B2(n_1828),
.Y(n_2179)
);

INVx1_ASAP7_75t_L g2180 ( 
.A(n_2133),
.Y(n_2180)
);

AND2x2_ASAP7_75t_L g2181 ( 
.A(n_2132),
.B(n_1856),
.Y(n_2181)
);

INVx2_ASAP7_75t_L g2182 ( 
.A(n_2127),
.Y(n_2182)
);

AND2x2_ASAP7_75t_L g2183 ( 
.A(n_2124),
.B(n_1856),
.Y(n_2183)
);

INVx2_ASAP7_75t_L g2184 ( 
.A(n_2141),
.Y(n_2184)
);

INVx1_ASAP7_75t_SL g2185 ( 
.A(n_2099),
.Y(n_2185)
);

AND2x2_ASAP7_75t_L g2186 ( 
.A(n_2089),
.B(n_1863),
.Y(n_2186)
);

AOI22xp33_ASAP7_75t_L g2187 ( 
.A1(n_2086),
.A2(n_1829),
.B1(n_1811),
.B2(n_1833),
.Y(n_2187)
);

AND2x2_ASAP7_75t_L g2188 ( 
.A(n_2142),
.B(n_1863),
.Y(n_2188)
);

AND2x2_ASAP7_75t_L g2189 ( 
.A(n_2121),
.B(n_1863),
.Y(n_2189)
);

AOI22xp5_ASAP7_75t_L g2190 ( 
.A1(n_2084),
.A2(n_703),
.B1(n_704),
.B2(n_699),
.Y(n_2190)
);

OR2x2_ASAP7_75t_L g2191 ( 
.A(n_2102),
.B(n_1931),
.Y(n_2191)
);

OAI221xp5_ASAP7_75t_L g2192 ( 
.A1(n_2097),
.A2(n_705),
.B1(n_714),
.B2(n_709),
.C(n_708),
.Y(n_2192)
);

INVx1_ASAP7_75t_L g2193 ( 
.A(n_2144),
.Y(n_2193)
);

INVx1_ASAP7_75t_L g2194 ( 
.A(n_2096),
.Y(n_2194)
);

NAND2xp5_ASAP7_75t_SL g2195 ( 
.A(n_2123),
.B(n_1825),
.Y(n_2195)
);

INVx1_ASAP7_75t_L g2196 ( 
.A(n_2111),
.Y(n_2196)
);

NOR2xp33_ASAP7_75t_L g2197 ( 
.A(n_2088),
.B(n_716),
.Y(n_2197)
);

NAND2xp5_ASAP7_75t_L g2198 ( 
.A(n_2128),
.B(n_1932),
.Y(n_2198)
);

NAND2xp5_ASAP7_75t_L g2199 ( 
.A(n_2109),
.B(n_723),
.Y(n_2199)
);

AND2x2_ASAP7_75t_L g2200 ( 
.A(n_2126),
.B(n_1868),
.Y(n_2200)
);

NAND2xp5_ASAP7_75t_L g2201 ( 
.A(n_2091),
.B(n_727),
.Y(n_2201)
);

INVx1_ASAP7_75t_L g2202 ( 
.A(n_2119),
.Y(n_2202)
);

INVx1_ASAP7_75t_L g2203 ( 
.A(n_2145),
.Y(n_2203)
);

INVx1_ASAP7_75t_L g2204 ( 
.A(n_2098),
.Y(n_2204)
);

NAND2xp5_ASAP7_75t_L g2205 ( 
.A(n_2117),
.B(n_728),
.Y(n_2205)
);

NAND2xp5_ASAP7_75t_L g2206 ( 
.A(n_2118),
.B(n_731),
.Y(n_2206)
);

INVxp67_ASAP7_75t_L g2207 ( 
.A(n_2140),
.Y(n_2207)
);

INVxp67_ASAP7_75t_L g2208 ( 
.A(n_2095),
.Y(n_2208)
);

AND2x2_ASAP7_75t_L g2209 ( 
.A(n_2129),
.B(n_1868),
.Y(n_2209)
);

INVx1_ASAP7_75t_L g2210 ( 
.A(n_2098),
.Y(n_2210)
);

HB1xp67_ASAP7_75t_L g2211 ( 
.A(n_2134),
.Y(n_2211)
);

NAND2xp5_ASAP7_75t_L g2212 ( 
.A(n_2105),
.B(n_736),
.Y(n_2212)
);

INVx1_ASAP7_75t_L g2213 ( 
.A(n_2093),
.Y(n_2213)
);

OR2x2_ASAP7_75t_L g2214 ( 
.A(n_2104),
.B(n_1966),
.Y(n_2214)
);

INVx1_ASAP7_75t_L g2215 ( 
.A(n_2104),
.Y(n_2215)
);

OAI22xp5_ASAP7_75t_L g2216 ( 
.A1(n_2083),
.A2(n_1966),
.B1(n_1825),
.B2(n_1767),
.Y(n_2216)
);

NOR2xp33_ASAP7_75t_L g2217 ( 
.A(n_2112),
.B(n_738),
.Y(n_2217)
);

NAND2xp5_ASAP7_75t_L g2218 ( 
.A(n_2135),
.B(n_739),
.Y(n_2218)
);

INVx1_ASAP7_75t_L g2219 ( 
.A(n_2104),
.Y(n_2219)
);

INVx1_ASAP7_75t_L g2220 ( 
.A(n_2104),
.Y(n_2220)
);

INVx1_ASAP7_75t_L g2221 ( 
.A(n_2104),
.Y(n_2221)
);

NAND2xp5_ASAP7_75t_L g2222 ( 
.A(n_2135),
.B(n_743),
.Y(n_2222)
);

INVx3_ASAP7_75t_L g2223 ( 
.A(n_2100),
.Y(n_2223)
);

NAND2xp5_ASAP7_75t_L g2224 ( 
.A(n_2135),
.B(n_744),
.Y(n_2224)
);

NAND2xp5_ASAP7_75t_L g2225 ( 
.A(n_2135),
.B(n_750),
.Y(n_2225)
);

AND2x2_ASAP7_75t_SL g2226 ( 
.A(n_2087),
.B(n_1825),
.Y(n_2226)
);

AND2x4_ASAP7_75t_L g2227 ( 
.A(n_2100),
.B(n_1921),
.Y(n_2227)
);

OR2x2_ASAP7_75t_L g2228 ( 
.A(n_2104),
.B(n_1966),
.Y(n_2228)
);

AOI22xp33_ASAP7_75t_L g2229 ( 
.A1(n_2083),
.A2(n_1829),
.B1(n_1833),
.B2(n_1818),
.Y(n_2229)
);

INVx1_ASAP7_75t_L g2230 ( 
.A(n_2104),
.Y(n_2230)
);

INVx1_ASAP7_75t_SL g2231 ( 
.A(n_2087),
.Y(n_2231)
);

INVx1_ASAP7_75t_L g2232 ( 
.A(n_2104),
.Y(n_2232)
);

NAND2x1_ASAP7_75t_L g2233 ( 
.A(n_2100),
.B(n_1966),
.Y(n_2233)
);

AOI221xp5_ASAP7_75t_L g2234 ( 
.A1(n_2204),
.A2(n_756),
.B1(n_759),
.B2(n_755),
.C(n_753),
.Y(n_2234)
);

INVx1_ASAP7_75t_L g2235 ( 
.A(n_2147),
.Y(n_2235)
);

OAI221xp5_ASAP7_75t_L g2236 ( 
.A1(n_2229),
.A2(n_777),
.B1(n_786),
.B2(n_775),
.C(n_765),
.Y(n_2236)
);

NAND2xp5_ASAP7_75t_L g2237 ( 
.A(n_2223),
.B(n_789),
.Y(n_2237)
);

NAND3xp33_ASAP7_75t_SL g2238 ( 
.A(n_2148),
.B(n_792),
.C(n_790),
.Y(n_2238)
);

OAI21xp33_ASAP7_75t_SL g2239 ( 
.A1(n_2211),
.A2(n_1899),
.B(n_1914),
.Y(n_2239)
);

INVx1_ASAP7_75t_L g2240 ( 
.A(n_2147),
.Y(n_2240)
);

AOI22xp5_ASAP7_75t_L g2241 ( 
.A1(n_2161),
.A2(n_920),
.B1(n_989),
.B2(n_909),
.Y(n_2241)
);

NAND4xp75_ASAP7_75t_L g2242 ( 
.A(n_2226),
.B(n_1652),
.C(n_1684),
.D(n_1760),
.Y(n_2242)
);

NAND2xp5_ASAP7_75t_SL g2243 ( 
.A(n_2148),
.B(n_1829),
.Y(n_2243)
);

NOR2xp33_ASAP7_75t_L g2244 ( 
.A(n_2231),
.B(n_795),
.Y(n_2244)
);

NAND2xp5_ASAP7_75t_L g2245 ( 
.A(n_2223),
.B(n_2152),
.Y(n_2245)
);

NOR4xp25_ASAP7_75t_L g2246 ( 
.A(n_2185),
.B(n_1706),
.C(n_1713),
.D(n_920),
.Y(n_2246)
);

OAI21xp5_ASAP7_75t_L g2247 ( 
.A1(n_2201),
.A2(n_2216),
.B(n_2208),
.Y(n_2247)
);

NAND2xp5_ASAP7_75t_L g2248 ( 
.A(n_2175),
.B(n_796),
.Y(n_2248)
);

AOI21xp5_ASAP7_75t_L g2249 ( 
.A1(n_2201),
.A2(n_1763),
.B(n_1706),
.Y(n_2249)
);

NAND4xp25_ASAP7_75t_L g2250 ( 
.A(n_2149),
.B(n_1769),
.C(n_1843),
.D(n_1740),
.Y(n_2250)
);

AOI211xp5_ASAP7_75t_L g2251 ( 
.A1(n_2216),
.A2(n_798),
.B(n_800),
.C(n_797),
.Y(n_2251)
);

NAND2xp33_ASAP7_75t_R g2252 ( 
.A(n_2157),
.B(n_2),
.Y(n_2252)
);

AOI22xp5_ASAP7_75t_L g2253 ( 
.A1(n_2154),
.A2(n_920),
.B1(n_909),
.B2(n_1829),
.Y(n_2253)
);

AOI221x1_ASAP7_75t_L g2254 ( 
.A1(n_2210),
.A2(n_1725),
.B1(n_752),
.B2(n_806),
.C(n_659),
.Y(n_2254)
);

AOI22xp5_ASAP7_75t_L g2255 ( 
.A1(n_2164),
.A2(n_909),
.B1(n_808),
.B2(n_809),
.Y(n_2255)
);

AOI21xp5_ASAP7_75t_L g2256 ( 
.A1(n_2207),
.A2(n_810),
.B(n_805),
.Y(n_2256)
);

NAND2xp5_ASAP7_75t_L g2257 ( 
.A(n_2197),
.B(n_811),
.Y(n_2257)
);

AOI21xp5_ASAP7_75t_L g2258 ( 
.A1(n_2231),
.A2(n_813),
.B(n_812),
.Y(n_2258)
);

AOI221xp5_ASAP7_75t_L g2259 ( 
.A1(n_2162),
.A2(n_824),
.B1(n_827),
.B2(n_820),
.C(n_818),
.Y(n_2259)
);

OAI21xp33_ASAP7_75t_L g2260 ( 
.A1(n_2215),
.A2(n_1857),
.B(n_1873),
.Y(n_2260)
);

OAI211xp5_ASAP7_75t_L g2261 ( 
.A1(n_2176),
.A2(n_834),
.B(n_836),
.C(n_835),
.Y(n_2261)
);

INVx1_ASAP7_75t_L g2262 ( 
.A(n_2182),
.Y(n_2262)
);

AOI221xp5_ASAP7_75t_L g2263 ( 
.A1(n_2213),
.A2(n_850),
.B1(n_851),
.B2(n_843),
.C(n_838),
.Y(n_2263)
);

INVx1_ASAP7_75t_L g2264 ( 
.A(n_2219),
.Y(n_2264)
);

AOI21xp33_ASAP7_75t_SL g2265 ( 
.A1(n_2220),
.A2(n_1),
.B(n_3),
.Y(n_2265)
);

AOI222xp33_ASAP7_75t_L g2266 ( 
.A1(n_2221),
.A2(n_863),
.B1(n_855),
.B2(n_864),
.C1(n_857),
.C2(n_852),
.Y(n_2266)
);

OAI21xp33_ASAP7_75t_L g2267 ( 
.A1(n_2230),
.A2(n_1857),
.B(n_1873),
.Y(n_2267)
);

NOR2xp33_ASAP7_75t_L g2268 ( 
.A(n_2232),
.B(n_866),
.Y(n_2268)
);

OAI211xp5_ASAP7_75t_SL g2269 ( 
.A1(n_2160),
.A2(n_1713),
.B(n_870),
.C(n_876),
.Y(n_2269)
);

NOR3xp33_ASAP7_75t_L g2270 ( 
.A(n_2192),
.B(n_877),
.C(n_868),
.Y(n_2270)
);

OAI211xp5_ASAP7_75t_SL g2271 ( 
.A1(n_2190),
.A2(n_879),
.B(n_881),
.C(n_878),
.Y(n_2271)
);

OAI221xp5_ASAP7_75t_L g2272 ( 
.A1(n_2187),
.A2(n_886),
.B1(n_887),
.B2(n_883),
.C(n_882),
.Y(n_2272)
);

AOI21xp5_ASAP7_75t_L g2273 ( 
.A1(n_2206),
.A2(n_892),
.B(n_889),
.Y(n_2273)
);

AOI21xp33_ASAP7_75t_L g2274 ( 
.A1(n_2185),
.A2(n_928),
.B(n_907),
.Y(n_2274)
);

NOR3xp33_ASAP7_75t_L g2275 ( 
.A(n_2218),
.B(n_897),
.C(n_895),
.Y(n_2275)
);

AOI22xp33_ASAP7_75t_L g2276 ( 
.A1(n_2172),
.A2(n_1810),
.B1(n_1818),
.B2(n_1843),
.Y(n_2276)
);

OAI21xp33_ASAP7_75t_L g2277 ( 
.A1(n_2178),
.A2(n_1857),
.B(n_1873),
.Y(n_2277)
);

OAI21xp5_ASAP7_75t_SL g2278 ( 
.A1(n_2153),
.A2(n_1849),
.B(n_752),
.Y(n_2278)
);

OAI221xp5_ASAP7_75t_SL g2279 ( 
.A1(n_2163),
.A2(n_1816),
.B1(n_1849),
.B2(n_1882),
.C(n_1875),
.Y(n_2279)
);

NAND4xp25_ASAP7_75t_L g2280 ( 
.A(n_2196),
.B(n_1843),
.C(n_1818),
.D(n_1771),
.Y(n_2280)
);

OAI21xp5_ASAP7_75t_L g2281 ( 
.A1(n_2190),
.A2(n_899),
.B(n_898),
.Y(n_2281)
);

NOR3xp33_ASAP7_75t_L g2282 ( 
.A(n_2222),
.B(n_910),
.C(n_902),
.Y(n_2282)
);

NOR3xp33_ASAP7_75t_L g2283 ( 
.A(n_2224),
.B(n_914),
.C(n_911),
.Y(n_2283)
);

OAI221xp5_ASAP7_75t_SL g2284 ( 
.A1(n_2163),
.A2(n_2174),
.B1(n_2171),
.B2(n_2179),
.C(n_2158),
.Y(n_2284)
);

INVx1_ASAP7_75t_L g2285 ( 
.A(n_2151),
.Y(n_2285)
);

AOI21xp5_ASAP7_75t_L g2286 ( 
.A1(n_2177),
.A2(n_919),
.B(n_917),
.Y(n_2286)
);

AOI211xp5_ASAP7_75t_L g2287 ( 
.A1(n_2155),
.A2(n_926),
.B(n_930),
.C(n_924),
.Y(n_2287)
);

AOI222xp33_ASAP7_75t_L g2288 ( 
.A1(n_2194),
.A2(n_936),
.B1(n_933),
.B2(n_937),
.C1(n_935),
.C2(n_931),
.Y(n_2288)
);

INVx1_ASAP7_75t_L g2289 ( 
.A(n_2191),
.Y(n_2289)
);

AOI211xp5_ASAP7_75t_L g2290 ( 
.A1(n_2202),
.A2(n_940),
.B(n_944),
.C(n_938),
.Y(n_2290)
);

OAI21xp33_ASAP7_75t_L g2291 ( 
.A1(n_2188),
.A2(n_1857),
.B(n_1875),
.Y(n_2291)
);

AOI22xp5_ASAP7_75t_L g2292 ( 
.A1(n_2195),
.A2(n_950),
.B1(n_953),
.B2(n_947),
.Y(n_2292)
);

NAND3xp33_ASAP7_75t_L g2293 ( 
.A(n_2203),
.B(n_659),
.C(n_640),
.Y(n_2293)
);

NAND4xp25_ASAP7_75t_L g2294 ( 
.A(n_2159),
.B(n_1843),
.C(n_1818),
.D(n_1771),
.Y(n_2294)
);

NOR2x1_ASAP7_75t_L g2295 ( 
.A(n_2184),
.B(n_659),
.Y(n_2295)
);

NOR2xp33_ASAP7_75t_L g2296 ( 
.A(n_2225),
.B(n_958),
.Y(n_2296)
);

NAND3xp33_ASAP7_75t_SL g2297 ( 
.A(n_2212),
.B(n_963),
.C(n_961),
.Y(n_2297)
);

NOR3xp33_ASAP7_75t_L g2298 ( 
.A(n_2217),
.B(n_971),
.C(n_970),
.Y(n_2298)
);

AND4x1_ASAP7_75t_L g2299 ( 
.A(n_2166),
.B(n_7),
.C(n_4),
.D(n_5),
.Y(n_2299)
);

AOI221x1_ASAP7_75t_L g2300 ( 
.A1(n_2180),
.A2(n_894),
.B1(n_806),
.B2(n_752),
.C(n_1656),
.Y(n_2300)
);

OR3x1_ASAP7_75t_L g2301 ( 
.A(n_2193),
.B(n_1844),
.C(n_1853),
.Y(n_2301)
);

AOI21xp5_ASAP7_75t_L g2302 ( 
.A1(n_2169),
.A2(n_973),
.B(n_972),
.Y(n_2302)
);

OAI211xp5_ASAP7_75t_SL g2303 ( 
.A1(n_2150),
.A2(n_2205),
.B(n_2199),
.C(n_2198),
.Y(n_2303)
);

A2O1A1Ixp33_ASAP7_75t_L g2304 ( 
.A1(n_2233),
.A2(n_983),
.B(n_987),
.C(n_981),
.Y(n_2304)
);

AOI21xp5_ASAP7_75t_L g2305 ( 
.A1(n_2167),
.A2(n_2173),
.B(n_2214),
.Y(n_2305)
);

AOI221xp5_ASAP7_75t_L g2306 ( 
.A1(n_2227),
.A2(n_2183),
.B1(n_2200),
.B2(n_2168),
.C(n_2228),
.Y(n_2306)
);

NAND3xp33_ASAP7_75t_L g2307 ( 
.A(n_2156),
.B(n_806),
.C(n_752),
.Y(n_2307)
);

NAND2xp5_ASAP7_75t_L g2308 ( 
.A(n_2165),
.B(n_990),
.Y(n_2308)
);

NAND3xp33_ASAP7_75t_L g2309 ( 
.A(n_2227),
.B(n_2170),
.C(n_2181),
.Y(n_2309)
);

AOI221xp5_ASAP7_75t_L g2310 ( 
.A1(n_2189),
.A2(n_993),
.B1(n_1001),
.B2(n_1000),
.C(n_999),
.Y(n_2310)
);

HB1xp67_ASAP7_75t_L g2311 ( 
.A(n_2186),
.Y(n_2311)
);

AOI211xp5_ASAP7_75t_L g2312 ( 
.A1(n_2209),
.A2(n_894),
.B(n_806),
.C(n_1771),
.Y(n_2312)
);

OAI21xp33_ASAP7_75t_L g2313 ( 
.A1(n_2229),
.A2(n_1883),
.B(n_1882),
.Y(n_2313)
);

INVx1_ASAP7_75t_L g2314 ( 
.A(n_2147),
.Y(n_2314)
);

AOI21xp5_ASAP7_75t_L g2315 ( 
.A1(n_2211),
.A2(n_1816),
.B(n_894),
.Y(n_2315)
);

AOI221xp5_ASAP7_75t_L g2316 ( 
.A1(n_2204),
.A2(n_894),
.B1(n_806),
.B2(n_1858),
.C(n_1853),
.Y(n_2316)
);

OAI21xp33_ASAP7_75t_L g2317 ( 
.A1(n_2229),
.A2(n_1883),
.B(n_1897),
.Y(n_2317)
);

NOR2xp33_ASAP7_75t_R g2318 ( 
.A(n_2223),
.B(n_5),
.Y(n_2318)
);

NAND2xp5_ASAP7_75t_SL g2319 ( 
.A(n_2148),
.B(n_1921),
.Y(n_2319)
);

OAI211xp5_ASAP7_75t_SL g2320 ( 
.A1(n_2207),
.A2(n_10),
.B(n_7),
.C(n_9),
.Y(n_2320)
);

INVx1_ASAP7_75t_L g2321 ( 
.A(n_2147),
.Y(n_2321)
);

O2A1O1Ixp33_ASAP7_75t_L g2322 ( 
.A1(n_2201),
.A2(n_1642),
.B(n_1816),
.C(n_1837),
.Y(n_2322)
);

NOR4xp25_ASAP7_75t_L g2323 ( 
.A(n_2185),
.B(n_1717),
.C(n_13),
.D(n_9),
.Y(n_2323)
);

AND4x1_ASAP7_75t_L g2324 ( 
.A(n_2190),
.B(n_15),
.C(n_11),
.D(n_13),
.Y(n_2324)
);

AOI321xp33_ASAP7_75t_L g2325 ( 
.A1(n_2149),
.A2(n_1883),
.A3(n_1885),
.B1(n_1840),
.B2(n_1766),
.C(n_1824),
.Y(n_2325)
);

NAND4xp25_ASAP7_75t_L g2326 ( 
.A(n_2161),
.B(n_1766),
.C(n_1840),
.D(n_1834),
.Y(n_2326)
);

AOI221xp5_ASAP7_75t_L g2327 ( 
.A1(n_2204),
.A2(n_894),
.B1(n_1858),
.B2(n_1937),
.C(n_1921),
.Y(n_2327)
);

AOI221xp5_ASAP7_75t_L g2328 ( 
.A1(n_2204),
.A2(n_1937),
.B1(n_1867),
.B2(n_1865),
.C(n_1864),
.Y(n_2328)
);

AOI22xp33_ASAP7_75t_L g2329 ( 
.A1(n_2204),
.A2(n_1816),
.B1(n_1824),
.B2(n_1822),
.Y(n_2329)
);

NAND2xp5_ASAP7_75t_L g2330 ( 
.A(n_2223),
.B(n_1937),
.Y(n_2330)
);

AOI211xp5_ASAP7_75t_SL g2331 ( 
.A1(n_2161),
.A2(n_1682),
.B(n_1656),
.C(n_18),
.Y(n_2331)
);

AO21x1_ASAP7_75t_L g2332 ( 
.A1(n_2201),
.A2(n_19),
.B(n_17),
.Y(n_2332)
);

AOI22xp5_ASAP7_75t_L g2333 ( 
.A1(n_2161),
.A2(n_1885),
.B1(n_1867),
.B2(n_1865),
.Y(n_2333)
);

AOI21xp5_ASAP7_75t_L g2334 ( 
.A1(n_2211),
.A2(n_1816),
.B(n_1729),
.Y(n_2334)
);

AND3x1_ASAP7_75t_L g2335 ( 
.A(n_2223),
.B(n_1682),
.C(n_1885),
.Y(n_2335)
);

OAI22xp5_ASAP7_75t_L g2336 ( 
.A1(n_2211),
.A2(n_1816),
.B1(n_1754),
.B2(n_1838),
.Y(n_2336)
);

OAI22xp33_ASAP7_75t_L g2337 ( 
.A1(n_2211),
.A2(n_1816),
.B1(n_1754),
.B2(n_1834),
.Y(n_2337)
);

AOI21xp5_ASAP7_75t_L g2338 ( 
.A1(n_2211),
.A2(n_1721),
.B(n_1686),
.Y(n_2338)
);

O2A1O1Ixp33_ASAP7_75t_L g2339 ( 
.A1(n_2201),
.A2(n_19),
.B(n_16),
.C(n_17),
.Y(n_2339)
);

OAI21xp5_ASAP7_75t_SL g2340 ( 
.A1(n_2161),
.A2(n_1840),
.B(n_1754),
.Y(n_2340)
);

AOI221xp5_ASAP7_75t_L g2341 ( 
.A1(n_2204),
.A2(n_1864),
.B1(n_1861),
.B2(n_1859),
.C(n_1871),
.Y(n_2341)
);

NOR3x1_ASAP7_75t_L g2342 ( 
.A(n_2157),
.B(n_16),
.C(n_21),
.Y(n_2342)
);

INVx1_ASAP7_75t_L g2343 ( 
.A(n_2147),
.Y(n_2343)
);

OAI22xp33_ASAP7_75t_L g2344 ( 
.A1(n_2211),
.A2(n_1754),
.B1(n_1834),
.B2(n_1824),
.Y(n_2344)
);

NOR2x1p5_ASAP7_75t_SL g2345 ( 
.A(n_2152),
.B(n_1861),
.Y(n_2345)
);

AOI221xp5_ASAP7_75t_L g2346 ( 
.A1(n_2204),
.A2(n_1886),
.B1(n_1893),
.B2(n_1876),
.C(n_1871),
.Y(n_2346)
);

OAI221xp5_ASAP7_75t_L g2347 ( 
.A1(n_2229),
.A2(n_1824),
.B1(n_1822),
.B2(n_1886),
.C(n_1876),
.Y(n_2347)
);

NAND2xp5_ASAP7_75t_L g2348 ( 
.A(n_2223),
.B(n_1868),
.Y(n_2348)
);

OAI221xp5_ASAP7_75t_L g2349 ( 
.A1(n_2229),
.A2(n_1822),
.B1(n_1894),
.B2(n_1896),
.C(n_1893),
.Y(n_2349)
);

OAI21xp5_ASAP7_75t_SL g2350 ( 
.A1(n_2161),
.A2(n_1822),
.B(n_1836),
.Y(n_2350)
);

OAI21xp5_ASAP7_75t_L g2351 ( 
.A1(n_2211),
.A2(n_1896),
.B(n_1894),
.Y(n_2351)
);

NAND2xp5_ASAP7_75t_L g2352 ( 
.A(n_2223),
.B(n_21),
.Y(n_2352)
);

AOI211xp5_ASAP7_75t_L g2353 ( 
.A1(n_2201),
.A2(n_26),
.B(n_23),
.C(n_25),
.Y(n_2353)
);

NOR3xp33_ASAP7_75t_L g2354 ( 
.A(n_2192),
.B(n_1664),
.C(n_1744),
.Y(n_2354)
);

INVx1_ASAP7_75t_L g2355 ( 
.A(n_2147),
.Y(n_2355)
);

OAI21xp5_ASAP7_75t_L g2356 ( 
.A1(n_2211),
.A2(n_1901),
.B(n_1814),
.Y(n_2356)
);

NOR4xp25_ASAP7_75t_L g2357 ( 
.A(n_2185),
.B(n_28),
.C(n_23),
.D(n_25),
.Y(n_2357)
);

OAI21xp5_ASAP7_75t_SL g2358 ( 
.A1(n_2161),
.A2(n_1823),
.B(n_1814),
.Y(n_2358)
);

NAND2xp5_ASAP7_75t_L g2359 ( 
.A(n_2223),
.B(n_29),
.Y(n_2359)
);

NAND4xp25_ASAP7_75t_L g2360 ( 
.A(n_2161),
.B(n_1834),
.C(n_1814),
.D(n_32),
.Y(n_2360)
);

OAI21xp33_ASAP7_75t_L g2361 ( 
.A1(n_2229),
.A2(n_1823),
.B(n_1901),
.Y(n_2361)
);

NAND2xp5_ASAP7_75t_SL g2362 ( 
.A(n_2148),
.B(n_1680),
.Y(n_2362)
);

OAI322xp33_ASAP7_75t_L g2363 ( 
.A1(n_2201),
.A2(n_1838),
.A3(n_1841),
.B1(n_1819),
.B2(n_1820),
.C1(n_1817),
.C2(n_33),
.Y(n_2363)
);

AOI21xp33_ASAP7_75t_L g2364 ( 
.A1(n_2201),
.A2(n_29),
.B(n_31),
.Y(n_2364)
);

NOR2xp33_ASAP7_75t_L g2365 ( 
.A(n_2148),
.B(n_35),
.Y(n_2365)
);

INVx1_ASAP7_75t_L g2366 ( 
.A(n_2147),
.Y(n_2366)
);

AOI21xp5_ASAP7_75t_L g2367 ( 
.A1(n_2211),
.A2(n_1808),
.B(n_1884),
.Y(n_2367)
);

AOI22xp33_ASAP7_75t_L g2368 ( 
.A1(n_2204),
.A2(n_1838),
.B1(n_1808),
.B2(n_1841),
.Y(n_2368)
);

NAND2xp5_ASAP7_75t_SL g2369 ( 
.A(n_2148),
.B(n_1680),
.Y(n_2369)
);

AOI221x1_ASAP7_75t_L g2370 ( 
.A1(n_2223),
.A2(n_1726),
.B1(n_38),
.B2(n_36),
.C(n_37),
.Y(n_2370)
);

NAND3xp33_ASAP7_75t_SL g2371 ( 
.A(n_2148),
.B(n_36),
.C(n_37),
.Y(n_2371)
);

AOI21xp5_ASAP7_75t_L g2372 ( 
.A1(n_2211),
.A2(n_1808),
.B(n_1884),
.Y(n_2372)
);

NAND2xp5_ASAP7_75t_L g2373 ( 
.A(n_2223),
.B(n_38),
.Y(n_2373)
);

AOI221xp5_ASAP7_75t_L g2374 ( 
.A1(n_2204),
.A2(n_1820),
.B1(n_1819),
.B2(n_1817),
.C(n_1884),
.Y(n_2374)
);

NAND2xp5_ASAP7_75t_L g2375 ( 
.A(n_2223),
.B(n_39),
.Y(n_2375)
);

AOI311xp33_ASAP7_75t_L g2376 ( 
.A1(n_2149),
.A2(n_1820),
.A3(n_1819),
.B(n_1817),
.C(n_42),
.Y(n_2376)
);

NAND2xp5_ASAP7_75t_L g2377 ( 
.A(n_2223),
.B(n_40),
.Y(n_2377)
);

AOI22xp5_ASAP7_75t_L g2378 ( 
.A1(n_2161),
.A2(n_1874),
.B1(n_1878),
.B2(n_1870),
.Y(n_2378)
);

AOI21xp33_ASAP7_75t_SL g2379 ( 
.A1(n_2226),
.A2(n_41),
.B(n_43),
.Y(n_2379)
);

NAND3xp33_ASAP7_75t_SL g2380 ( 
.A(n_2148),
.B(n_43),
.C(n_44),
.Y(n_2380)
);

NAND2xp5_ASAP7_75t_L g2381 ( 
.A(n_2223),
.B(n_45),
.Y(n_2381)
);

AOI221xp5_ASAP7_75t_L g2382 ( 
.A1(n_2204),
.A2(n_1888),
.B1(n_1903),
.B2(n_1900),
.C(n_1887),
.Y(n_2382)
);

NAND2xp5_ASAP7_75t_L g2383 ( 
.A(n_2223),
.B(n_45),
.Y(n_2383)
);

AOI211xp5_ASAP7_75t_L g2384 ( 
.A1(n_2364),
.A2(n_50),
.B(n_48),
.C(n_49),
.Y(n_2384)
);

INVx1_ASAP7_75t_L g2385 ( 
.A(n_2311),
.Y(n_2385)
);

OAI22xp5_ASAP7_75t_SL g2386 ( 
.A1(n_2357),
.A2(n_50),
.B1(n_48),
.B2(n_49),
.Y(n_2386)
);

HB1xp67_ASAP7_75t_L g2387 ( 
.A(n_2318),
.Y(n_2387)
);

AOI221x1_ASAP7_75t_L g2388 ( 
.A1(n_2364),
.A2(n_53),
.B1(n_51),
.B2(n_52),
.C(n_55),
.Y(n_2388)
);

NAND3xp33_ASAP7_75t_L g2389 ( 
.A(n_2331),
.B(n_53),
.C(n_56),
.Y(n_2389)
);

INVx1_ASAP7_75t_L g2390 ( 
.A(n_2352),
.Y(n_2390)
);

O2A1O1Ixp5_ASAP7_75t_L g2391 ( 
.A1(n_2284),
.A2(n_1888),
.B(n_1900),
.C(n_1887),
.Y(n_2391)
);

NOR2x1_ASAP7_75t_L g2392 ( 
.A(n_2371),
.B(n_2380),
.Y(n_2392)
);

O2A1O1Ixp33_ASAP7_75t_L g2393 ( 
.A1(n_2339),
.A2(n_58),
.B(n_56),
.C(n_57),
.Y(n_2393)
);

AOI21xp33_ASAP7_75t_L g2394 ( 
.A1(n_2252),
.A2(n_61),
.B(n_63),
.Y(n_2394)
);

INVx2_ASAP7_75t_L g2395 ( 
.A(n_2245),
.Y(n_2395)
);

INVx2_ASAP7_75t_L g2396 ( 
.A(n_2301),
.Y(n_2396)
);

OAI22xp33_ASAP7_75t_L g2397 ( 
.A1(n_2370),
.A2(n_1841),
.B1(n_1888),
.B2(n_1887),
.Y(n_2397)
);

NAND2xp5_ASAP7_75t_SL g2398 ( 
.A(n_2323),
.B(n_1900),
.Y(n_2398)
);

OAI211xp5_ASAP7_75t_SL g2399 ( 
.A1(n_2247),
.A2(n_65),
.B(n_63),
.C(n_64),
.Y(n_2399)
);

INVx2_ASAP7_75t_L g2400 ( 
.A(n_2335),
.Y(n_2400)
);

OAI211xp5_ASAP7_75t_L g2401 ( 
.A1(n_2376),
.A2(n_67),
.B(n_64),
.C(n_65),
.Y(n_2401)
);

INVx1_ASAP7_75t_L g2402 ( 
.A(n_2359),
.Y(n_2402)
);

INVx1_ASAP7_75t_L g2403 ( 
.A(n_2373),
.Y(n_2403)
);

NAND2xp33_ASAP7_75t_SL g2404 ( 
.A(n_2375),
.B(n_1841),
.Y(n_2404)
);

OA22x2_ASAP7_75t_SL g2405 ( 
.A1(n_2235),
.A2(n_1870),
.B1(n_1878),
.B2(n_1874),
.Y(n_2405)
);

AOI21xp33_ASAP7_75t_L g2406 ( 
.A1(n_2244),
.A2(n_2239),
.B(n_2344),
.Y(n_2406)
);

NAND3xp33_ASAP7_75t_L g2407 ( 
.A(n_2251),
.B(n_2353),
.C(n_2263),
.Y(n_2407)
);

AOI222xp33_ASAP7_75t_L g2408 ( 
.A1(n_2351),
.A2(n_70),
.B1(n_72),
.B2(n_68),
.C1(n_69),
.C2(n_71),
.Y(n_2408)
);

AND2x2_ASAP7_75t_L g2409 ( 
.A(n_2342),
.B(n_70),
.Y(n_2409)
);

CKINVDCx20_ASAP7_75t_R g2410 ( 
.A(n_2332),
.Y(n_2410)
);

NAND2xp5_ASAP7_75t_L g2411 ( 
.A(n_2379),
.B(n_71),
.Y(n_2411)
);

INVx2_ASAP7_75t_L g2412 ( 
.A(n_2377),
.Y(n_2412)
);

OAI221xp5_ASAP7_75t_SL g2413 ( 
.A1(n_2340),
.A2(n_74),
.B1(n_72),
.B2(n_73),
.C(n_75),
.Y(n_2413)
);

AND4x1_ASAP7_75t_L g2414 ( 
.A(n_2365),
.B(n_76),
.C(n_73),
.D(n_75),
.Y(n_2414)
);

OAI211xp5_ASAP7_75t_L g2415 ( 
.A1(n_2315),
.A2(n_80),
.B(n_77),
.C(n_79),
.Y(n_2415)
);

OAI322xp33_ASAP7_75t_L g2416 ( 
.A1(n_2240),
.A2(n_85),
.A3(n_84),
.B1(n_82),
.B2(n_77),
.C1(n_81),
.C2(n_83),
.Y(n_2416)
);

A2O1A1Ixp33_ASAP7_75t_L g2417 ( 
.A1(n_2265),
.A2(n_85),
.B(n_81),
.C(n_84),
.Y(n_2417)
);

A2O1A1Ixp33_ASAP7_75t_L g2418 ( 
.A1(n_2356),
.A2(n_90),
.B(n_87),
.C(n_89),
.Y(n_2418)
);

INVx1_ASAP7_75t_L g2419 ( 
.A(n_2381),
.Y(n_2419)
);

INVx1_ASAP7_75t_L g2420 ( 
.A(n_2383),
.Y(n_2420)
);

INVx1_ASAP7_75t_L g2421 ( 
.A(n_2262),
.Y(n_2421)
);

NOR2xp33_ASAP7_75t_L g2422 ( 
.A(n_2360),
.B(n_90),
.Y(n_2422)
);

OAI22xp5_ASAP7_75t_L g2423 ( 
.A1(n_2255),
.A2(n_1903),
.B1(n_1874),
.B2(n_1878),
.Y(n_2423)
);

A2O1A1Ixp33_ASAP7_75t_SL g2424 ( 
.A1(n_2314),
.A2(n_93),
.B(n_91),
.C(n_92),
.Y(n_2424)
);

AOI221xp5_ASAP7_75t_L g2425 ( 
.A1(n_2363),
.A2(n_93),
.B1(n_91),
.B2(n_92),
.C(n_94),
.Y(n_2425)
);

INVx1_ASAP7_75t_L g2426 ( 
.A(n_2321),
.Y(n_2426)
);

O2A1O1Ixp33_ASAP7_75t_L g2427 ( 
.A1(n_2274),
.A2(n_98),
.B(n_95),
.C(n_96),
.Y(n_2427)
);

NOR2x1p5_ASAP7_75t_L g2428 ( 
.A(n_2238),
.B(n_96),
.Y(n_2428)
);

AOI22xp5_ASAP7_75t_L g2429 ( 
.A1(n_2348),
.A2(n_1903),
.B1(n_1804),
.B2(n_1847),
.Y(n_2429)
);

NAND2xp5_ASAP7_75t_L g2430 ( 
.A(n_2343),
.B(n_99),
.Y(n_2430)
);

NAND2xp5_ASAP7_75t_L g2431 ( 
.A(n_2355),
.B(n_2366),
.Y(n_2431)
);

INVx1_ASAP7_75t_L g2432 ( 
.A(n_2309),
.Y(n_2432)
);

INVx2_ASAP7_75t_L g2433 ( 
.A(n_2295),
.Y(n_2433)
);

INVx1_ASAP7_75t_L g2434 ( 
.A(n_2299),
.Y(n_2434)
);

AOI22xp5_ASAP7_75t_L g2435 ( 
.A1(n_2320),
.A2(n_2326),
.B1(n_2336),
.B2(n_2250),
.Y(n_2435)
);

AOI31xp33_ASAP7_75t_L g2436 ( 
.A1(n_2274),
.A2(n_101),
.A3(n_99),
.B(n_100),
.Y(n_2436)
);

AOI21xp5_ASAP7_75t_L g2437 ( 
.A1(n_2286),
.A2(n_2258),
.B(n_2302),
.Y(n_2437)
);

AOI222xp33_ASAP7_75t_L g2438 ( 
.A1(n_2259),
.A2(n_105),
.B1(n_107),
.B2(n_100),
.C1(n_102),
.C2(n_106),
.Y(n_2438)
);

NAND2xp5_ASAP7_75t_L g2439 ( 
.A(n_2324),
.B(n_102),
.Y(n_2439)
);

HB1xp67_ASAP7_75t_L g2440 ( 
.A(n_2243),
.Y(n_2440)
);

NAND2xp5_ASAP7_75t_L g2441 ( 
.A(n_2296),
.B(n_106),
.Y(n_2441)
);

AND2x4_ASAP7_75t_L g2442 ( 
.A(n_2289),
.B(n_107),
.Y(n_2442)
);

NAND2xp5_ASAP7_75t_L g2443 ( 
.A(n_2268),
.B(n_108),
.Y(n_2443)
);

O2A1O1Ixp5_ASAP7_75t_L g2444 ( 
.A1(n_2319),
.A2(n_1847),
.B(n_111),
.C(n_109),
.Y(n_2444)
);

OAI32xp33_ASAP7_75t_L g2445 ( 
.A1(n_2264),
.A2(n_1847),
.A3(n_113),
.B1(n_110),
.B2(n_112),
.Y(n_2445)
);

OAI21xp5_ASAP7_75t_L g2446 ( 
.A1(n_2305),
.A2(n_1821),
.B(n_110),
.Y(n_2446)
);

INVx1_ASAP7_75t_L g2447 ( 
.A(n_2285),
.Y(n_2447)
);

NOR2xp33_ASAP7_75t_L g2448 ( 
.A(n_2248),
.B(n_112),
.Y(n_2448)
);

A2O1A1Ixp33_ASAP7_75t_L g2449 ( 
.A1(n_2322),
.A2(n_116),
.B(n_114),
.C(n_115),
.Y(n_2449)
);

OAI221xp5_ASAP7_75t_SL g2450 ( 
.A1(n_2306),
.A2(n_116),
.B1(n_114),
.B2(n_115),
.C(n_118),
.Y(n_2450)
);

AOI22xp5_ASAP7_75t_L g2451 ( 
.A1(n_2336),
.A2(n_1804),
.B1(n_1847),
.B2(n_1808),
.Y(n_2451)
);

NOR2x1_ASAP7_75t_SL g2452 ( 
.A(n_2362),
.B(n_120),
.Y(n_2452)
);

INVx2_ASAP7_75t_L g2453 ( 
.A(n_2242),
.Y(n_2453)
);

AOI222xp33_ASAP7_75t_L g2454 ( 
.A1(n_2303),
.A2(n_124),
.B1(n_126),
.B2(n_120),
.C1(n_123),
.C2(n_125),
.Y(n_2454)
);

O2A1O1Ixp33_ASAP7_75t_L g2455 ( 
.A1(n_2369),
.A2(n_126),
.B(n_124),
.C(n_125),
.Y(n_2455)
);

OAI211xp5_ASAP7_75t_L g2456 ( 
.A1(n_2292),
.A2(n_129),
.B(n_127),
.C(n_128),
.Y(n_2456)
);

AOI221xp5_ASAP7_75t_L g2457 ( 
.A1(n_2337),
.A2(n_130),
.B1(n_127),
.B2(n_128),
.C(n_132),
.Y(n_2457)
);

OAI21xp33_ASAP7_75t_L g2458 ( 
.A1(n_2361),
.A2(n_1798),
.B(n_1821),
.Y(n_2458)
);

AOI21xp5_ASAP7_75t_L g2459 ( 
.A1(n_2256),
.A2(n_1808),
.B(n_130),
.Y(n_2459)
);

AOI21xp5_ASAP7_75t_L g2460 ( 
.A1(n_2257),
.A2(n_1808),
.B(n_133),
.Y(n_2460)
);

CKINVDCx5p33_ASAP7_75t_R g2461 ( 
.A(n_2241),
.Y(n_2461)
);

BUFx6f_ASAP7_75t_L g2462 ( 
.A(n_2237),
.Y(n_2462)
);

AOI221xp5_ASAP7_75t_L g2463 ( 
.A1(n_2316),
.A2(n_135),
.B1(n_133),
.B2(n_134),
.C(n_136),
.Y(n_2463)
);

AOI211xp5_ASAP7_75t_L g2464 ( 
.A1(n_2272),
.A2(n_137),
.B(n_134),
.C(n_135),
.Y(n_2464)
);

O2A1O1Ixp33_ASAP7_75t_L g2465 ( 
.A1(n_2304),
.A2(n_141),
.B(n_137),
.C(n_138),
.Y(n_2465)
);

INVx3_ASAP7_75t_L g2466 ( 
.A(n_2330),
.Y(n_2466)
);

OAI22xp5_ASAP7_75t_L g2467 ( 
.A1(n_2276),
.A2(n_1798),
.B1(n_1804),
.B2(n_1830),
.Y(n_2467)
);

AOI22xp5_ASAP7_75t_L g2468 ( 
.A1(n_2280),
.A2(n_1804),
.B1(n_1798),
.B2(n_1830),
.Y(n_2468)
);

NOR4xp25_ASAP7_75t_L g2469 ( 
.A(n_2261),
.B(n_142),
.C(n_138),
.D(n_141),
.Y(n_2469)
);

INVx2_ASAP7_75t_L g2470 ( 
.A(n_2308),
.Y(n_2470)
);

NAND2xp5_ASAP7_75t_L g2471 ( 
.A(n_2266),
.B(n_142),
.Y(n_2471)
);

OAI21xp33_ASAP7_75t_L g2472 ( 
.A1(n_2358),
.A2(n_1798),
.B(n_1821),
.Y(n_2472)
);

AOI21xp5_ASAP7_75t_L g2473 ( 
.A1(n_2367),
.A2(n_143),
.B(n_145),
.Y(n_2473)
);

INVx1_ASAP7_75t_L g2474 ( 
.A(n_2345),
.Y(n_2474)
);

A2O1A1Ixp33_ASAP7_75t_L g2475 ( 
.A1(n_2372),
.A2(n_147),
.B(n_145),
.C(n_146),
.Y(n_2475)
);

INVx1_ASAP7_75t_L g2476 ( 
.A(n_2307),
.Y(n_2476)
);

AOI22xp5_ASAP7_75t_L g2477 ( 
.A1(n_2294),
.A2(n_1804),
.B1(n_1798),
.B2(n_1830),
.Y(n_2477)
);

NAND4xp25_ASAP7_75t_SL g2478 ( 
.A(n_2300),
.B(n_149),
.C(n_146),
.D(n_148),
.Y(n_2478)
);

O2A1O1Ixp33_ASAP7_75t_SL g2479 ( 
.A1(n_2249),
.A2(n_150),
.B(n_148),
.C(n_149),
.Y(n_2479)
);

OAI22xp5_ASAP7_75t_L g2480 ( 
.A1(n_2329),
.A2(n_1798),
.B1(n_1804),
.B2(n_1830),
.Y(n_2480)
);

INVx3_ASAP7_75t_L g2481 ( 
.A(n_2350),
.Y(n_2481)
);

A2O1A1Ixp33_ASAP7_75t_L g2482 ( 
.A1(n_2234),
.A2(n_152),
.B(n_150),
.C(n_151),
.Y(n_2482)
);

OAI311xp33_ASAP7_75t_L g2483 ( 
.A1(n_2278),
.A2(n_154),
.A3(n_151),
.B1(n_153),
.C1(n_155),
.Y(n_2483)
);

OAI22xp33_ASAP7_75t_L g2484 ( 
.A1(n_2254),
.A2(n_1798),
.B1(n_1830),
.B2(n_155),
.Y(n_2484)
);

BUFx2_ASAP7_75t_L g2485 ( 
.A(n_2281),
.Y(n_2485)
);

AOI21xp5_ASAP7_75t_SL g2486 ( 
.A1(n_2297),
.A2(n_153),
.B(n_154),
.Y(n_2486)
);

AOI221xp5_ASAP7_75t_L g2487 ( 
.A1(n_2327),
.A2(n_2374),
.B1(n_2334),
.B2(n_2328),
.C(n_2310),
.Y(n_2487)
);

XOR2xp5_ASAP7_75t_L g2488 ( 
.A(n_2253),
.B(n_156),
.Y(n_2488)
);

OAI21xp5_ASAP7_75t_SL g2489 ( 
.A1(n_2236),
.A2(n_157),
.B(n_158),
.Y(n_2489)
);

OAI21xp33_ASAP7_75t_L g2490 ( 
.A1(n_2317),
.A2(n_2313),
.B(n_2291),
.Y(n_2490)
);

NOR2xp33_ASAP7_75t_L g2491 ( 
.A(n_2271),
.B(n_158),
.Y(n_2491)
);

O2A1O1Ixp33_ASAP7_75t_L g2492 ( 
.A1(n_2290),
.A2(n_161),
.B(n_159),
.C(n_160),
.Y(n_2492)
);

NOR2xp33_ASAP7_75t_L g2493 ( 
.A(n_2273),
.B(n_159),
.Y(n_2493)
);

AOI211xp5_ASAP7_75t_L g2494 ( 
.A1(n_2246),
.A2(n_166),
.B(n_163),
.C(n_164),
.Y(n_2494)
);

AOI221xp5_ASAP7_75t_L g2495 ( 
.A1(n_2293),
.A2(n_168),
.B1(n_163),
.B2(n_164),
.C(n_169),
.Y(n_2495)
);

AOI322xp5_ASAP7_75t_L g2496 ( 
.A1(n_2275),
.A2(n_170),
.A3(n_171),
.B1(n_172),
.B2(n_173),
.C1(n_174),
.C2(n_175),
.Y(n_2496)
);

INVxp67_ASAP7_75t_L g2497 ( 
.A(n_2288),
.Y(n_2497)
);

AOI222xp33_ASAP7_75t_L g2498 ( 
.A1(n_2341),
.A2(n_176),
.B1(n_178),
.B2(n_171),
.C1(n_175),
.C2(n_177),
.Y(n_2498)
);

OR2x2_ASAP7_75t_L g2499 ( 
.A(n_2282),
.B(n_176),
.Y(n_2499)
);

INVxp67_ASAP7_75t_L g2500 ( 
.A(n_2270),
.Y(n_2500)
);

NOR2xp33_ASAP7_75t_L g2501 ( 
.A(n_2283),
.B(n_178),
.Y(n_2501)
);

INVx1_ASAP7_75t_L g2502 ( 
.A(n_2287),
.Y(n_2502)
);

INVx1_ASAP7_75t_L g2503 ( 
.A(n_2387),
.Y(n_2503)
);

INVxp67_ASAP7_75t_L g2504 ( 
.A(n_2392),
.Y(n_2504)
);

NAND2xp5_ASAP7_75t_SL g2505 ( 
.A(n_2386),
.B(n_2382),
.Y(n_2505)
);

AND2x2_ASAP7_75t_L g2506 ( 
.A(n_2434),
.B(n_2298),
.Y(n_2506)
);

INVx1_ASAP7_75t_L g2507 ( 
.A(n_2385),
.Y(n_2507)
);

INVx1_ASAP7_75t_L g2508 ( 
.A(n_2409),
.Y(n_2508)
);

NAND2xp5_ASAP7_75t_L g2509 ( 
.A(n_2414),
.B(n_2312),
.Y(n_2509)
);

AOI21xp5_ASAP7_75t_L g2510 ( 
.A1(n_2401),
.A2(n_2338),
.B(n_2354),
.Y(n_2510)
);

NAND2xp5_ASAP7_75t_SL g2511 ( 
.A(n_2397),
.B(n_2346),
.Y(n_2511)
);

INVx1_ASAP7_75t_L g2512 ( 
.A(n_2442),
.Y(n_2512)
);

OR2x2_ASAP7_75t_L g2513 ( 
.A(n_2389),
.B(n_2333),
.Y(n_2513)
);

OR2x2_ASAP7_75t_L g2514 ( 
.A(n_2469),
.B(n_2260),
.Y(n_2514)
);

NOR2xp33_ASAP7_75t_L g2515 ( 
.A(n_2394),
.B(n_2269),
.Y(n_2515)
);

NAND2xp5_ASAP7_75t_SL g2516 ( 
.A(n_2410),
.B(n_2325),
.Y(n_2516)
);

NAND2xp5_ASAP7_75t_L g2517 ( 
.A(n_2442),
.B(n_2267),
.Y(n_2517)
);

NAND2xp33_ASAP7_75t_SL g2518 ( 
.A(n_2428),
.B(n_2440),
.Y(n_2518)
);

AND2x2_ASAP7_75t_L g2519 ( 
.A(n_2395),
.B(n_2277),
.Y(n_2519)
);

NOR2xp33_ASAP7_75t_L g2520 ( 
.A(n_2439),
.B(n_2349),
.Y(n_2520)
);

OR2x2_ASAP7_75t_L g2521 ( 
.A(n_2432),
.B(n_2450),
.Y(n_2521)
);

BUFx6f_ASAP7_75t_L g2522 ( 
.A(n_2430),
.Y(n_2522)
);

OR2x2_ASAP7_75t_L g2523 ( 
.A(n_2421),
.B(n_2368),
.Y(n_2523)
);

AOI21xp5_ASAP7_75t_L g2524 ( 
.A1(n_2393),
.A2(n_2347),
.B(n_2279),
.Y(n_2524)
);

AND2x2_ASAP7_75t_L g2525 ( 
.A(n_2422),
.B(n_2378),
.Y(n_2525)
);

AND2x2_ASAP7_75t_L g2526 ( 
.A(n_2452),
.B(n_180),
.Y(n_2526)
);

INVx1_ASAP7_75t_L g2527 ( 
.A(n_2396),
.Y(n_2527)
);

INVx1_ASAP7_75t_L g2528 ( 
.A(n_2411),
.Y(n_2528)
);

INVxp67_ASAP7_75t_L g2529 ( 
.A(n_2491),
.Y(n_2529)
);

NAND3xp33_ASAP7_75t_L g2530 ( 
.A(n_2425),
.B(n_181),
.C(n_182),
.Y(n_2530)
);

BUFx6f_ASAP7_75t_L g2531 ( 
.A(n_2462),
.Y(n_2531)
);

INVx1_ASAP7_75t_L g2532 ( 
.A(n_2474),
.Y(n_2532)
);

OR2x2_ASAP7_75t_L g2533 ( 
.A(n_2431),
.B(n_181),
.Y(n_2533)
);

NAND2xp5_ASAP7_75t_L g2534 ( 
.A(n_2417),
.B(n_182),
.Y(n_2534)
);

INVx2_ASAP7_75t_L g2535 ( 
.A(n_2405),
.Y(n_2535)
);

AOI221xp5_ASAP7_75t_L g2536 ( 
.A1(n_2406),
.A2(n_185),
.B1(n_183),
.B2(n_184),
.C(n_186),
.Y(n_2536)
);

INVx1_ASAP7_75t_L g2537 ( 
.A(n_2441),
.Y(n_2537)
);

INVx1_ASAP7_75t_L g2538 ( 
.A(n_2443),
.Y(n_2538)
);

INVx1_ASAP7_75t_L g2539 ( 
.A(n_2426),
.Y(n_2539)
);

NAND2xp5_ASAP7_75t_L g2540 ( 
.A(n_2384),
.B(n_183),
.Y(n_2540)
);

INVx2_ASAP7_75t_SL g2541 ( 
.A(n_2400),
.Y(n_2541)
);

NAND2xp5_ASAP7_75t_L g2542 ( 
.A(n_2388),
.B(n_185),
.Y(n_2542)
);

INVx1_ASAP7_75t_SL g2543 ( 
.A(n_2499),
.Y(n_2543)
);

NAND2xp5_ASAP7_75t_L g2544 ( 
.A(n_2454),
.B(n_187),
.Y(n_2544)
);

INVx1_ASAP7_75t_L g2545 ( 
.A(n_2412),
.Y(n_2545)
);

INVx1_ASAP7_75t_SL g2546 ( 
.A(n_2461),
.Y(n_2546)
);

INVx2_ASAP7_75t_L g2547 ( 
.A(n_2462),
.Y(n_2547)
);

NOR3xp33_ASAP7_75t_L g2548 ( 
.A(n_2407),
.B(n_188),
.C(n_189),
.Y(n_2548)
);

AND2x2_ASAP7_75t_L g2549 ( 
.A(n_2390),
.B(n_188),
.Y(n_2549)
);

NOR2xp33_ASAP7_75t_L g2550 ( 
.A(n_2436),
.B(n_191),
.Y(n_2550)
);

NAND2xp5_ASAP7_75t_L g2551 ( 
.A(n_2424),
.B(n_191),
.Y(n_2551)
);

NAND2xp5_ASAP7_75t_L g2552 ( 
.A(n_2448),
.B(n_2493),
.Y(n_2552)
);

INVx1_ASAP7_75t_L g2553 ( 
.A(n_2402),
.Y(n_2553)
);

NAND2xp5_ASAP7_75t_L g2554 ( 
.A(n_2494),
.B(n_192),
.Y(n_2554)
);

INVx1_ASAP7_75t_L g2555 ( 
.A(n_2403),
.Y(n_2555)
);

AOI21xp5_ASAP7_75t_L g2556 ( 
.A1(n_2479),
.A2(n_193),
.B(n_195),
.Y(n_2556)
);

NAND2xp5_ASAP7_75t_L g2557 ( 
.A(n_2497),
.B(n_195),
.Y(n_2557)
);

INVx1_ASAP7_75t_L g2558 ( 
.A(n_2419),
.Y(n_2558)
);

INVx1_ASAP7_75t_L g2559 ( 
.A(n_2420),
.Y(n_2559)
);

OAI21xp33_ASAP7_75t_L g2560 ( 
.A1(n_2490),
.A2(n_1801),
.B(n_196),
.Y(n_2560)
);

AOI221x1_ASAP7_75t_SL g2561 ( 
.A1(n_2447),
.A2(n_198),
.B1(n_196),
.B2(n_197),
.C(n_200),
.Y(n_2561)
);

OAI21xp33_ASAP7_75t_SL g2562 ( 
.A1(n_2398),
.A2(n_2435),
.B(n_2481),
.Y(n_2562)
);

NOR2xp33_ASAP7_75t_L g2563 ( 
.A(n_2399),
.B(n_202),
.Y(n_2563)
);

INVxp67_ASAP7_75t_SL g2564 ( 
.A(n_2455),
.Y(n_2564)
);

AND2x2_ASAP7_75t_L g2565 ( 
.A(n_2470),
.B(n_203),
.Y(n_2565)
);

NAND2xp5_ASAP7_75t_L g2566 ( 
.A(n_2462),
.B(n_206),
.Y(n_2566)
);

INVxp67_ASAP7_75t_L g2567 ( 
.A(n_2501),
.Y(n_2567)
);

INVx1_ASAP7_75t_L g2568 ( 
.A(n_2466),
.Y(n_2568)
);

OR2x2_ASAP7_75t_L g2569 ( 
.A(n_2413),
.B(n_209),
.Y(n_2569)
);

OR2x2_ASAP7_75t_L g2570 ( 
.A(n_2471),
.B(n_209),
.Y(n_2570)
);

OAI31xp33_ASAP7_75t_L g2571 ( 
.A1(n_2483),
.A2(n_213),
.A3(n_210),
.B(n_211),
.Y(n_2571)
);

NAND2x1_ASAP7_75t_SL g2572 ( 
.A(n_2481),
.B(n_211),
.Y(n_2572)
);

INVx1_ASAP7_75t_L g2573 ( 
.A(n_2466),
.Y(n_2573)
);

OAI221xp5_ASAP7_75t_L g2574 ( 
.A1(n_2391),
.A2(n_215),
.B1(n_213),
.B2(n_214),
.C(n_216),
.Y(n_2574)
);

NOR2x1_ASAP7_75t_L g2575 ( 
.A(n_2478),
.B(n_215),
.Y(n_2575)
);

INVx2_ASAP7_75t_L g2576 ( 
.A(n_2433),
.Y(n_2576)
);

NOR2x1_ASAP7_75t_L g2577 ( 
.A(n_2486),
.B(n_217),
.Y(n_2577)
);

NOR2x1_ASAP7_75t_L g2578 ( 
.A(n_2416),
.B(n_218),
.Y(n_2578)
);

INVx1_ASAP7_75t_L g2579 ( 
.A(n_2453),
.Y(n_2579)
);

INVx1_ASAP7_75t_L g2580 ( 
.A(n_2502),
.Y(n_2580)
);

AND2x2_ASAP7_75t_L g2581 ( 
.A(n_2485),
.B(n_219),
.Y(n_2581)
);

CKINVDCx5p33_ASAP7_75t_R g2582 ( 
.A(n_2500),
.Y(n_2582)
);

AND2x2_ASAP7_75t_L g2583 ( 
.A(n_2446),
.B(n_221),
.Y(n_2583)
);

NAND2xp5_ASAP7_75t_L g2584 ( 
.A(n_2464),
.B(n_223),
.Y(n_2584)
);

INVx1_ASAP7_75t_L g2585 ( 
.A(n_2488),
.Y(n_2585)
);

NOR2x1_ASAP7_75t_L g2586 ( 
.A(n_2456),
.B(n_223),
.Y(n_2586)
);

NOR2xp33_ASAP7_75t_L g2587 ( 
.A(n_2489),
.B(n_224),
.Y(n_2587)
);

INVx1_ASAP7_75t_L g2588 ( 
.A(n_2427),
.Y(n_2588)
);

AOI21xp5_ASAP7_75t_L g2589 ( 
.A1(n_2473),
.A2(n_225),
.B(n_226),
.Y(n_2589)
);

AOI21xp33_ASAP7_75t_L g2590 ( 
.A1(n_2484),
.A2(n_227),
.B(n_228),
.Y(n_2590)
);

NAND2xp5_ASAP7_75t_L g2591 ( 
.A(n_2437),
.B(n_228),
.Y(n_2591)
);

NAND2xp5_ASAP7_75t_L g2592 ( 
.A(n_2438),
.B(n_229),
.Y(n_2592)
);

NAND2xp5_ASAP7_75t_L g2593 ( 
.A(n_2482),
.B(n_229),
.Y(n_2593)
);

INVx1_ASAP7_75t_L g2594 ( 
.A(n_2476),
.Y(n_2594)
);

INVxp67_ASAP7_75t_L g2595 ( 
.A(n_2408),
.Y(n_2595)
);

INVx1_ASAP7_75t_L g2596 ( 
.A(n_2445),
.Y(n_2596)
);

NAND2xp5_ASAP7_75t_L g2597 ( 
.A(n_2496),
.B(n_230),
.Y(n_2597)
);

INVx2_ASAP7_75t_SL g2598 ( 
.A(n_2423),
.Y(n_2598)
);

NOR2x1_ASAP7_75t_L g2599 ( 
.A(n_2415),
.B(n_230),
.Y(n_2599)
);

AND2x2_ASAP7_75t_L g2600 ( 
.A(n_2449),
.B(n_2418),
.Y(n_2600)
);

NOR2xp67_ASAP7_75t_L g2601 ( 
.A(n_2460),
.B(n_231),
.Y(n_2601)
);

NAND2xp5_ASAP7_75t_SL g2602 ( 
.A(n_2444),
.B(n_231),
.Y(n_2602)
);

OAI221xp5_ASAP7_75t_L g2603 ( 
.A1(n_2457),
.A2(n_2487),
.B1(n_2463),
.B2(n_2475),
.C(n_2459),
.Y(n_2603)
);

AND2x2_ASAP7_75t_L g2604 ( 
.A(n_2498),
.B(n_233),
.Y(n_2604)
);

INVx1_ASAP7_75t_SL g2605 ( 
.A(n_2404),
.Y(n_2605)
);

OAI32xp33_ASAP7_75t_L g2606 ( 
.A1(n_2458),
.A2(n_235),
.A3(n_233),
.B1(n_234),
.B2(n_236),
.Y(n_2606)
);

AOI221xp5_ASAP7_75t_L g2607 ( 
.A1(n_2492),
.A2(n_236),
.B1(n_234),
.B2(n_235),
.C(n_239),
.Y(n_2607)
);

NAND2xp5_ASAP7_75t_L g2608 ( 
.A(n_2495),
.B(n_239),
.Y(n_2608)
);

AND2x2_ASAP7_75t_L g2609 ( 
.A(n_2472),
.B(n_240),
.Y(n_2609)
);

OAI21xp33_ASAP7_75t_SL g2610 ( 
.A1(n_2477),
.A2(n_240),
.B(n_241),
.Y(n_2610)
);

AND2x2_ASAP7_75t_L g2611 ( 
.A(n_2468),
.B(n_243),
.Y(n_2611)
);

INVx1_ASAP7_75t_L g2612 ( 
.A(n_2465),
.Y(n_2612)
);

INVx1_ASAP7_75t_L g2613 ( 
.A(n_2429),
.Y(n_2613)
);

INVx2_ASAP7_75t_SL g2614 ( 
.A(n_2467),
.Y(n_2614)
);

OA21x2_ASAP7_75t_L g2615 ( 
.A1(n_2451),
.A2(n_243),
.B(n_244),
.Y(n_2615)
);

AND2x2_ASAP7_75t_L g2616 ( 
.A(n_2480),
.B(n_244),
.Y(n_2616)
);

INVx1_ASAP7_75t_L g2617 ( 
.A(n_2387),
.Y(n_2617)
);

INVx1_ASAP7_75t_L g2618 ( 
.A(n_2387),
.Y(n_2618)
);

OR2x2_ASAP7_75t_L g2619 ( 
.A(n_2387),
.B(n_245),
.Y(n_2619)
);

NAND2xp5_ASAP7_75t_SL g2620 ( 
.A(n_2392),
.B(n_245),
.Y(n_2620)
);

INVxp33_ASAP7_75t_L g2621 ( 
.A(n_2392),
.Y(n_2621)
);

AOI22xp5_ASAP7_75t_L g2622 ( 
.A1(n_2410),
.A2(n_1830),
.B1(n_1801),
.B2(n_248),
.Y(n_2622)
);

NOR2x1_ASAP7_75t_L g2623 ( 
.A(n_2478),
.B(n_246),
.Y(n_2623)
);

INVx1_ASAP7_75t_L g2624 ( 
.A(n_2387),
.Y(n_2624)
);

INVx2_ASAP7_75t_L g2625 ( 
.A(n_2452),
.Y(n_2625)
);

NOR3xp33_ASAP7_75t_L g2626 ( 
.A(n_2450),
.B(n_247),
.C(n_248),
.Y(n_2626)
);

OAI221xp5_ASAP7_75t_L g2627 ( 
.A1(n_2392),
.A2(n_251),
.B1(n_247),
.B2(n_250),
.C(n_253),
.Y(n_2627)
);

NOR3xp33_ASAP7_75t_L g2628 ( 
.A(n_2450),
.B(n_250),
.C(n_254),
.Y(n_2628)
);

INVx2_ASAP7_75t_SL g2629 ( 
.A(n_2387),
.Y(n_2629)
);

OR2x2_ASAP7_75t_L g2630 ( 
.A(n_2387),
.B(n_254),
.Y(n_2630)
);

AND2x4_ASAP7_75t_L g2631 ( 
.A(n_2387),
.B(n_255),
.Y(n_2631)
);

NAND2xp5_ASAP7_75t_L g2632 ( 
.A(n_2387),
.B(n_257),
.Y(n_2632)
);

INVx1_ASAP7_75t_L g2633 ( 
.A(n_2387),
.Y(n_2633)
);

AND2x2_ASAP7_75t_L g2634 ( 
.A(n_2387),
.B(n_257),
.Y(n_2634)
);

INVx1_ASAP7_75t_L g2635 ( 
.A(n_2387),
.Y(n_2635)
);

NAND2xp5_ASAP7_75t_L g2636 ( 
.A(n_2387),
.B(n_258),
.Y(n_2636)
);

OR2x2_ASAP7_75t_L g2637 ( 
.A(n_2387),
.B(n_258),
.Y(n_2637)
);

NOR2x1_ASAP7_75t_L g2638 ( 
.A(n_2478),
.B(n_259),
.Y(n_2638)
);

OR2x2_ASAP7_75t_L g2639 ( 
.A(n_2387),
.B(n_259),
.Y(n_2639)
);

INVx1_ASAP7_75t_SL g2640 ( 
.A(n_2387),
.Y(n_2640)
);

NAND3xp33_ASAP7_75t_L g2641 ( 
.A(n_2392),
.B(n_260),
.C(n_261),
.Y(n_2641)
);

INVx1_ASAP7_75t_L g2642 ( 
.A(n_2387),
.Y(n_2642)
);

INVx1_ASAP7_75t_L g2643 ( 
.A(n_2387),
.Y(n_2643)
);

HB1xp67_ASAP7_75t_L g2644 ( 
.A(n_2387),
.Y(n_2644)
);

INVx1_ASAP7_75t_L g2645 ( 
.A(n_2387),
.Y(n_2645)
);

INVx1_ASAP7_75t_L g2646 ( 
.A(n_2387),
.Y(n_2646)
);

AND2x2_ASAP7_75t_L g2647 ( 
.A(n_2387),
.B(n_260),
.Y(n_2647)
);

INVx1_ASAP7_75t_L g2648 ( 
.A(n_2387),
.Y(n_2648)
);

INVx2_ASAP7_75t_SL g2649 ( 
.A(n_2387),
.Y(n_2649)
);

NOR2x1_ASAP7_75t_L g2650 ( 
.A(n_2478),
.B(n_261),
.Y(n_2650)
);

NAND2xp5_ASAP7_75t_L g2651 ( 
.A(n_2387),
.B(n_262),
.Y(n_2651)
);

AND2x2_ASAP7_75t_L g2652 ( 
.A(n_2508),
.B(n_263),
.Y(n_2652)
);

NAND2xp33_ASAP7_75t_SL g2653 ( 
.A(n_2572),
.B(n_263),
.Y(n_2653)
);

AOI32xp33_ASAP7_75t_L g2654 ( 
.A1(n_2621),
.A2(n_266),
.A3(n_264),
.B1(n_265),
.B2(n_267),
.Y(n_2654)
);

NOR2xp33_ASAP7_75t_R g2655 ( 
.A(n_2518),
.B(n_264),
.Y(n_2655)
);

NAND4xp75_ASAP7_75t_L g2656 ( 
.A(n_2562),
.B(n_2578),
.C(n_2620),
.D(n_2577),
.Y(n_2656)
);

AOI22xp5_ASAP7_75t_L g2657 ( 
.A1(n_2504),
.A2(n_1801),
.B1(n_271),
.B2(n_267),
.Y(n_2657)
);

OAI221xp5_ASAP7_75t_SL g2658 ( 
.A1(n_2571),
.A2(n_274),
.B1(n_269),
.B2(n_272),
.C(n_276),
.Y(n_2658)
);

AND3x1_ASAP7_75t_L g2659 ( 
.A(n_2626),
.B(n_272),
.C(n_274),
.Y(n_2659)
);

AOI22xp5_ASAP7_75t_L g2660 ( 
.A1(n_2629),
.A2(n_2649),
.B1(n_2640),
.B2(n_2541),
.Y(n_2660)
);

OAI21x1_ASAP7_75t_L g2661 ( 
.A1(n_2556),
.A2(n_1752),
.B(n_1657),
.Y(n_2661)
);

INVx1_ASAP7_75t_L g2662 ( 
.A(n_2644),
.Y(n_2662)
);

AOI32xp33_ASAP7_75t_L g2663 ( 
.A1(n_2575),
.A2(n_280),
.A3(n_277),
.B1(n_279),
.B2(n_282),
.Y(n_2663)
);

NOR2xp33_ASAP7_75t_L g2664 ( 
.A(n_2512),
.B(n_277),
.Y(n_2664)
);

INVxp67_ASAP7_75t_L g2665 ( 
.A(n_2531),
.Y(n_2665)
);

O2A1O1Ixp33_ASAP7_75t_L g2666 ( 
.A1(n_2542),
.A2(n_284),
.B(n_282),
.C(n_283),
.Y(n_2666)
);

AND2x2_ASAP7_75t_L g2667 ( 
.A(n_2623),
.B(n_283),
.Y(n_2667)
);

AOI221xp5_ASAP7_75t_L g2668 ( 
.A1(n_2536),
.A2(n_286),
.B1(n_284),
.B2(n_285),
.C(n_287),
.Y(n_2668)
);

AOI21xp5_ASAP7_75t_L g2669 ( 
.A1(n_2516),
.A2(n_287),
.B(n_289),
.Y(n_2669)
);

NAND2xp5_ASAP7_75t_L g2670 ( 
.A(n_2631),
.B(n_2634),
.Y(n_2670)
);

NOR2xp67_ASAP7_75t_L g2671 ( 
.A(n_2625),
.B(n_2526),
.Y(n_2671)
);

BUFx2_ASAP7_75t_L g2672 ( 
.A(n_2531),
.Y(n_2672)
);

OAI221xp5_ASAP7_75t_L g2673 ( 
.A1(n_2560),
.A2(n_292),
.B1(n_293),
.B2(n_294),
.C(n_295),
.Y(n_2673)
);

INVx1_ASAP7_75t_L g2674 ( 
.A(n_2531),
.Y(n_2674)
);

INVxp67_ASAP7_75t_SL g2675 ( 
.A(n_2638),
.Y(n_2675)
);

AOI221x1_ASAP7_75t_L g2676 ( 
.A1(n_2548),
.A2(n_293),
.B1(n_294),
.B2(n_295),
.C(n_296),
.Y(n_2676)
);

INVxp67_ASAP7_75t_SL g2677 ( 
.A(n_2650),
.Y(n_2677)
);

INVx1_ASAP7_75t_L g2678 ( 
.A(n_2647),
.Y(n_2678)
);

NAND2xp33_ASAP7_75t_R g2679 ( 
.A(n_2551),
.B(n_297),
.Y(n_2679)
);

NOR2xp33_ASAP7_75t_L g2680 ( 
.A(n_2546),
.B(n_297),
.Y(n_2680)
);

INVx1_ASAP7_75t_L g2681 ( 
.A(n_2619),
.Y(n_2681)
);

NAND4xp25_ASAP7_75t_SL g2682 ( 
.A(n_2510),
.B(n_301),
.C(n_298),
.D(n_300),
.Y(n_2682)
);

INVx1_ASAP7_75t_L g2683 ( 
.A(n_2630),
.Y(n_2683)
);

OR2x2_ASAP7_75t_L g2684 ( 
.A(n_2637),
.B(n_302),
.Y(n_2684)
);

NAND2xp5_ASAP7_75t_L g2685 ( 
.A(n_2631),
.B(n_303),
.Y(n_2685)
);

NAND2xp5_ASAP7_75t_L g2686 ( 
.A(n_2561),
.B(n_303),
.Y(n_2686)
);

XOR2xp5_ASAP7_75t_L g2687 ( 
.A(n_2521),
.B(n_305),
.Y(n_2687)
);

HB1xp67_ASAP7_75t_L g2688 ( 
.A(n_2639),
.Y(n_2688)
);

NAND2xp5_ASAP7_75t_L g2689 ( 
.A(n_2503),
.B(n_2617),
.Y(n_2689)
);

OAI22xp5_ASAP7_75t_L g2690 ( 
.A1(n_2530),
.A2(n_2527),
.B1(n_2596),
.B2(n_2618),
.Y(n_2690)
);

AOI322xp5_ASAP7_75t_L g2691 ( 
.A1(n_2564),
.A2(n_305),
.A3(n_306),
.B1(n_307),
.B2(n_308),
.C1(n_309),
.C2(n_310),
.Y(n_2691)
);

NAND2xp33_ASAP7_75t_L g2692 ( 
.A(n_2628),
.B(n_307),
.Y(n_2692)
);

HB1xp67_ASAP7_75t_L g2693 ( 
.A(n_2581),
.Y(n_2693)
);

INVx1_ASAP7_75t_L g2694 ( 
.A(n_2532),
.Y(n_2694)
);

AND2x4_ASAP7_75t_L g2695 ( 
.A(n_2547),
.B(n_310),
.Y(n_2695)
);

AOI221xp5_ASAP7_75t_L g2696 ( 
.A1(n_2590),
.A2(n_311),
.B1(n_312),
.B2(n_313),
.C(n_314),
.Y(n_2696)
);

NAND2xp5_ASAP7_75t_L g2697 ( 
.A(n_2624),
.B(n_311),
.Y(n_2697)
);

AND2x4_ASAP7_75t_L g2698 ( 
.A(n_2633),
.B(n_313),
.Y(n_2698)
);

INVx1_ASAP7_75t_SL g2699 ( 
.A(n_2566),
.Y(n_2699)
);

INVx1_ASAP7_75t_L g2700 ( 
.A(n_2635),
.Y(n_2700)
);

NOR2xp33_ASAP7_75t_L g2701 ( 
.A(n_2642),
.B(n_314),
.Y(n_2701)
);

NOR2x1_ASAP7_75t_L g2702 ( 
.A(n_2641),
.B(n_315),
.Y(n_2702)
);

CKINVDCx5p33_ASAP7_75t_R g2703 ( 
.A(n_2582),
.Y(n_2703)
);

O2A1O1Ixp5_ASAP7_75t_L g2704 ( 
.A1(n_2505),
.A2(n_318),
.B(n_316),
.C(n_317),
.Y(n_2704)
);

NAND2xp5_ASAP7_75t_L g2705 ( 
.A(n_2643),
.B(n_317),
.Y(n_2705)
);

INVx1_ASAP7_75t_L g2706 ( 
.A(n_2645),
.Y(n_2706)
);

AOI211xp5_ASAP7_75t_L g2707 ( 
.A1(n_2606),
.A2(n_320),
.B(n_318),
.C(n_319),
.Y(n_2707)
);

AOI21xp5_ASAP7_75t_L g2708 ( 
.A1(n_2591),
.A2(n_319),
.B(n_321),
.Y(n_2708)
);

INVx3_ASAP7_75t_SL g2709 ( 
.A(n_2522),
.Y(n_2709)
);

NAND2xp33_ASAP7_75t_SL g2710 ( 
.A(n_2602),
.B(n_322),
.Y(n_2710)
);

A2O1A1Ixp33_ASAP7_75t_SL g2711 ( 
.A1(n_2646),
.A2(n_327),
.B(n_325),
.C(n_326),
.Y(n_2711)
);

INVx1_ASAP7_75t_L g2712 ( 
.A(n_2648),
.Y(n_2712)
);

A2O1A1Ixp33_ASAP7_75t_SL g2713 ( 
.A1(n_2507),
.A2(n_327),
.B(n_325),
.C(n_326),
.Y(n_2713)
);

AOI21xp5_ASAP7_75t_L g2714 ( 
.A1(n_2589),
.A2(n_328),
.B(n_330),
.Y(n_2714)
);

INVx1_ASAP7_75t_SL g2715 ( 
.A(n_2565),
.Y(n_2715)
);

INVx1_ASAP7_75t_L g2716 ( 
.A(n_2632),
.Y(n_2716)
);

AOI21xp33_ASAP7_75t_SL g2717 ( 
.A1(n_2627),
.A2(n_328),
.B(n_331),
.Y(n_2717)
);

NOR2xp33_ASAP7_75t_R g2718 ( 
.A(n_2588),
.B(n_331),
.Y(n_2718)
);

NAND2xp5_ASAP7_75t_L g2719 ( 
.A(n_2550),
.B(n_332),
.Y(n_2719)
);

INVx3_ASAP7_75t_L g2720 ( 
.A(n_2522),
.Y(n_2720)
);

INVx1_ASAP7_75t_L g2721 ( 
.A(n_2636),
.Y(n_2721)
);

NOR2xp33_ASAP7_75t_R g2722 ( 
.A(n_2568),
.B(n_332),
.Y(n_2722)
);

AO22x2_ASAP7_75t_L g2723 ( 
.A1(n_2569),
.A2(n_335),
.B1(n_333),
.B2(n_334),
.Y(n_2723)
);

INVx2_ASAP7_75t_L g2724 ( 
.A(n_2535),
.Y(n_2724)
);

AOI21xp5_ASAP7_75t_L g2725 ( 
.A1(n_2592),
.A2(n_333),
.B(n_334),
.Y(n_2725)
);

NAND2xp5_ASAP7_75t_L g2726 ( 
.A(n_2563),
.B(n_335),
.Y(n_2726)
);

OAI211xp5_ASAP7_75t_L g2727 ( 
.A1(n_2599),
.A2(n_338),
.B(n_336),
.C(n_337),
.Y(n_2727)
);

NAND2xp33_ASAP7_75t_R g2728 ( 
.A(n_2604),
.B(n_337),
.Y(n_2728)
);

CKINVDCx20_ASAP7_75t_R g2729 ( 
.A(n_2595),
.Y(n_2729)
);

NAND2xp5_ASAP7_75t_L g2730 ( 
.A(n_2549),
.B(n_338),
.Y(n_2730)
);

INVx1_ASAP7_75t_L g2731 ( 
.A(n_2651),
.Y(n_2731)
);

OAI221xp5_ASAP7_75t_L g2732 ( 
.A1(n_2610),
.A2(n_339),
.B1(n_340),
.B2(n_341),
.C(n_342),
.Y(n_2732)
);

NOR2xp33_ASAP7_75t_L g2733 ( 
.A(n_2514),
.B(n_339),
.Y(n_2733)
);

INVx1_ASAP7_75t_L g2734 ( 
.A(n_2533),
.Y(n_2734)
);

INVx2_ASAP7_75t_SL g2735 ( 
.A(n_2573),
.Y(n_2735)
);

AND2x4_ASAP7_75t_L g2736 ( 
.A(n_2576),
.B(n_340),
.Y(n_2736)
);

OAI221xp5_ASAP7_75t_L g2737 ( 
.A1(n_2603),
.A2(n_341),
.B1(n_342),
.B2(n_344),
.C(n_345),
.Y(n_2737)
);

OAI22xp5_ASAP7_75t_L g2738 ( 
.A1(n_2513),
.A2(n_347),
.B1(n_344),
.B2(n_346),
.Y(n_2738)
);

INVx1_ASAP7_75t_L g2739 ( 
.A(n_2519),
.Y(n_2739)
);

OAI22xp5_ASAP7_75t_L g2740 ( 
.A1(n_2660),
.A2(n_2579),
.B1(n_2597),
.B2(n_2612),
.Y(n_2740)
);

AND2x2_ASAP7_75t_L g2741 ( 
.A(n_2675),
.B(n_2586),
.Y(n_2741)
);

OR2x2_ASAP7_75t_L g2742 ( 
.A(n_2670),
.B(n_2544),
.Y(n_2742)
);

NAND4xp75_ASAP7_75t_L g2743 ( 
.A(n_2671),
.B(n_2669),
.C(n_2702),
.D(n_2662),
.Y(n_2743)
);

INVx1_ASAP7_75t_L g2744 ( 
.A(n_2667),
.Y(n_2744)
);

NOR2xp33_ASAP7_75t_L g2745 ( 
.A(n_2658),
.B(n_2529),
.Y(n_2745)
);

NOR2xp33_ASAP7_75t_R g2746 ( 
.A(n_2653),
.B(n_2585),
.Y(n_2746)
);

AO21x1_ASAP7_75t_L g2747 ( 
.A1(n_2710),
.A2(n_2557),
.B(n_2554),
.Y(n_2747)
);

NAND2xp5_ASAP7_75t_L g2748 ( 
.A(n_2677),
.B(n_2600),
.Y(n_2748)
);

NAND2xp5_ASAP7_75t_SL g2749 ( 
.A(n_2720),
.B(n_2655),
.Y(n_2749)
);

OR2x2_ASAP7_75t_L g2750 ( 
.A(n_2709),
.B(n_2517),
.Y(n_2750)
);

OAI22xp5_ASAP7_75t_SL g2751 ( 
.A1(n_2659),
.A2(n_2587),
.B1(n_2515),
.B2(n_2509),
.Y(n_2751)
);

NOR3xp33_ASAP7_75t_L g2752 ( 
.A(n_2656),
.B(n_2528),
.C(n_2567),
.Y(n_2752)
);

INVxp67_ASAP7_75t_L g2753 ( 
.A(n_2672),
.Y(n_2753)
);

AND2x4_ASAP7_75t_SL g2754 ( 
.A(n_2720),
.B(n_2522),
.Y(n_2754)
);

INVx4_ASAP7_75t_L g2755 ( 
.A(n_2703),
.Y(n_2755)
);

OR5x1_ASAP7_75t_L g2756 ( 
.A(n_2682),
.B(n_2523),
.C(n_2614),
.D(n_2605),
.E(n_2598),
.Y(n_2756)
);

AND2x2_ASAP7_75t_L g2757 ( 
.A(n_2693),
.B(n_2525),
.Y(n_2757)
);

AOI22xp5_ASAP7_75t_L g2758 ( 
.A1(n_2729),
.A2(n_2520),
.B1(n_2506),
.B2(n_2580),
.Y(n_2758)
);

INVx2_ASAP7_75t_SL g2759 ( 
.A(n_2698),
.Y(n_2759)
);

CKINVDCx5p33_ASAP7_75t_R g2760 ( 
.A(n_2728),
.Y(n_2760)
);

NOR2x1_ASAP7_75t_L g2761 ( 
.A(n_2727),
.B(n_2540),
.Y(n_2761)
);

INVx2_ASAP7_75t_L g2762 ( 
.A(n_2695),
.Y(n_2762)
);

INVx1_ASAP7_75t_L g2763 ( 
.A(n_2652),
.Y(n_2763)
);

NOR2x1_ASAP7_75t_L g2764 ( 
.A(n_2684),
.B(n_2539),
.Y(n_2764)
);

NAND4xp75_ASAP7_75t_L g2765 ( 
.A(n_2733),
.B(n_2545),
.C(n_2594),
.D(n_2555),
.Y(n_2765)
);

NAND4xp75_ASAP7_75t_L g2766 ( 
.A(n_2739),
.B(n_2558),
.C(n_2559),
.D(n_2553),
.Y(n_2766)
);

NOR2xp33_ASAP7_75t_R g2767 ( 
.A(n_2679),
.B(n_2534),
.Y(n_2767)
);

HB1xp67_ASAP7_75t_L g2768 ( 
.A(n_2722),
.Y(n_2768)
);

OR2x2_ASAP7_75t_L g2769 ( 
.A(n_2686),
.B(n_2570),
.Y(n_2769)
);

NOR2xp33_ASAP7_75t_L g2770 ( 
.A(n_2665),
.B(n_2543),
.Y(n_2770)
);

NAND2x1p5_ASAP7_75t_SL g2771 ( 
.A(n_2735),
.B(n_2609),
.Y(n_2771)
);

OAI211xp5_ASAP7_75t_L g2772 ( 
.A1(n_2718),
.A2(n_2607),
.B(n_2552),
.C(n_2601),
.Y(n_2772)
);

NOR2x1_ASAP7_75t_L g2773 ( 
.A(n_2685),
.B(n_2584),
.Y(n_2773)
);

AOI211xp5_ASAP7_75t_L g2774 ( 
.A1(n_2690),
.A2(n_2574),
.B(n_2583),
.C(n_2538),
.Y(n_2774)
);

NAND2x1p5_ASAP7_75t_L g2775 ( 
.A(n_2715),
.B(n_2681),
.Y(n_2775)
);

NAND2xp5_ASAP7_75t_L g2776 ( 
.A(n_2691),
.B(n_2537),
.Y(n_2776)
);

NAND4xp75_ASAP7_75t_L g2777 ( 
.A(n_2689),
.B(n_2616),
.C(n_2608),
.D(n_2593),
.Y(n_2777)
);

INVx1_ASAP7_75t_L g2778 ( 
.A(n_2688),
.Y(n_2778)
);

XOR2x1_ASAP7_75t_L g2779 ( 
.A(n_2736),
.B(n_2695),
.Y(n_2779)
);

NOR2x1_ASAP7_75t_L g2780 ( 
.A(n_2736),
.B(n_2683),
.Y(n_2780)
);

NOR3xp33_ASAP7_75t_SL g2781 ( 
.A(n_2700),
.B(n_2511),
.C(n_2524),
.Y(n_2781)
);

NOR2xp33_ASAP7_75t_R g2782 ( 
.A(n_2678),
.B(n_2692),
.Y(n_2782)
);

OAI211xp5_ASAP7_75t_SL g2783 ( 
.A1(n_2706),
.A2(n_2613),
.B(n_2622),
.C(n_2615),
.Y(n_2783)
);

INVx1_ASAP7_75t_L g2784 ( 
.A(n_2723),
.Y(n_2784)
);

AND3x2_ASAP7_75t_L g2785 ( 
.A(n_2674),
.B(n_2611),
.C(n_2615),
.Y(n_2785)
);

NOR2x1_ASAP7_75t_SL g2786 ( 
.A(n_2712),
.B(n_346),
.Y(n_2786)
);

INVx1_ASAP7_75t_L g2787 ( 
.A(n_2723),
.Y(n_2787)
);

NAND4xp75_ASAP7_75t_L g2788 ( 
.A(n_2725),
.B(n_351),
.C(n_347),
.D(n_350),
.Y(n_2788)
);

BUFx2_ASAP7_75t_L g2789 ( 
.A(n_2698),
.Y(n_2789)
);

NAND2xp5_ASAP7_75t_L g2790 ( 
.A(n_2663),
.B(n_351),
.Y(n_2790)
);

INVxp67_ASAP7_75t_L g2791 ( 
.A(n_2664),
.Y(n_2791)
);

NAND4xp75_ASAP7_75t_L g2792 ( 
.A(n_2704),
.B(n_354),
.C(n_352),
.D(n_353),
.Y(n_2792)
);

AOI221xp5_ASAP7_75t_SL g2793 ( 
.A1(n_2717),
.A2(n_352),
.B1(n_354),
.B2(n_355),
.C(n_357),
.Y(n_2793)
);

INVx3_ASAP7_75t_L g2794 ( 
.A(n_2734),
.Y(n_2794)
);

INVx3_ASAP7_75t_L g2795 ( 
.A(n_2724),
.Y(n_2795)
);

NOR3xp33_ASAP7_75t_L g2796 ( 
.A(n_2666),
.B(n_355),
.C(n_357),
.Y(n_2796)
);

INVxp33_ASAP7_75t_L g2797 ( 
.A(n_2687),
.Y(n_2797)
);

INVxp67_ASAP7_75t_SL g2798 ( 
.A(n_2779),
.Y(n_2798)
);

NOR2xp33_ASAP7_75t_L g2799 ( 
.A(n_2789),
.B(n_2737),
.Y(n_2799)
);

NOR2x1p5_ASAP7_75t_L g2800 ( 
.A(n_2792),
.B(n_2719),
.Y(n_2800)
);

NAND4xp75_ASAP7_75t_L g2801 ( 
.A(n_2780),
.B(n_2764),
.C(n_2773),
.D(n_2741),
.Y(n_2801)
);

XNOR2x1_ASAP7_75t_L g2802 ( 
.A(n_2750),
.B(n_2699),
.Y(n_2802)
);

HB1xp67_ASAP7_75t_L g2803 ( 
.A(n_2784),
.Y(n_2803)
);

OR2x2_ASAP7_75t_L g2804 ( 
.A(n_2759),
.B(n_2697),
.Y(n_2804)
);

XNOR2xp5_ASAP7_75t_L g2805 ( 
.A(n_2740),
.B(n_2707),
.Y(n_2805)
);

NAND4xp75_ASAP7_75t_L g2806 ( 
.A(n_2761),
.B(n_2787),
.C(n_2749),
.D(n_2747),
.Y(n_2806)
);

NAND2xp5_ASAP7_75t_SL g2807 ( 
.A(n_2760),
.B(n_2654),
.Y(n_2807)
);

INVxp67_ASAP7_75t_SL g2808 ( 
.A(n_2786),
.Y(n_2808)
);

INVx1_ASAP7_75t_L g2809 ( 
.A(n_2754),
.Y(n_2809)
);

INVx2_ASAP7_75t_L g2810 ( 
.A(n_2775),
.Y(n_2810)
);

INVx2_ASAP7_75t_L g2811 ( 
.A(n_2762),
.Y(n_2811)
);

AND2x2_ASAP7_75t_L g2812 ( 
.A(n_2757),
.B(n_2680),
.Y(n_2812)
);

INVx2_ASAP7_75t_L g2813 ( 
.A(n_2771),
.Y(n_2813)
);

OAI22xp5_ASAP7_75t_L g2814 ( 
.A1(n_2753),
.A2(n_2732),
.B1(n_2673),
.B2(n_2726),
.Y(n_2814)
);

NAND4xp75_ASAP7_75t_L g2815 ( 
.A(n_2781),
.B(n_2694),
.C(n_2676),
.D(n_2716),
.Y(n_2815)
);

INVx2_ASAP7_75t_L g2816 ( 
.A(n_2795),
.Y(n_2816)
);

NAND4xp75_ASAP7_75t_L g2817 ( 
.A(n_2748),
.B(n_2731),
.C(n_2721),
.D(n_2705),
.Y(n_2817)
);

NAND2xp5_ASAP7_75t_L g2818 ( 
.A(n_2785),
.B(n_2701),
.Y(n_2818)
);

INVx2_ASAP7_75t_L g2819 ( 
.A(n_2795),
.Y(n_2819)
);

AND2x4_ASAP7_75t_L g2820 ( 
.A(n_2794),
.B(n_2730),
.Y(n_2820)
);

INVx1_ASAP7_75t_L g2821 ( 
.A(n_2768),
.Y(n_2821)
);

CKINVDCx20_ASAP7_75t_R g2822 ( 
.A(n_2751),
.Y(n_2822)
);

INVx1_ASAP7_75t_L g2823 ( 
.A(n_2794),
.Y(n_2823)
);

NAND2xp5_ASAP7_75t_L g2824 ( 
.A(n_2778),
.B(n_2711),
.Y(n_2824)
);

NOR3x1_ASAP7_75t_L g2825 ( 
.A(n_2743),
.B(n_2713),
.C(n_2738),
.Y(n_2825)
);

XNOR2xp5_ASAP7_75t_L g2826 ( 
.A(n_2756),
.B(n_2696),
.Y(n_2826)
);

A2O1A1Ixp33_ASAP7_75t_L g2827 ( 
.A1(n_2770),
.A2(n_2714),
.B(n_2708),
.C(n_2668),
.Y(n_2827)
);

INVx2_ASAP7_75t_L g2828 ( 
.A(n_2755),
.Y(n_2828)
);

NOR4xp25_ASAP7_75t_L g2829 ( 
.A(n_2783),
.B(n_2657),
.C(n_2661),
.D(n_360),
.Y(n_2829)
);

AND3x4_ASAP7_75t_L g2830 ( 
.A(n_2752),
.B(n_358),
.C(n_359),
.Y(n_2830)
);

NOR4xp25_ASAP7_75t_L g2831 ( 
.A(n_2772),
.B(n_360),
.C(n_358),
.D(n_359),
.Y(n_2831)
);

OR2x6_ASAP7_75t_L g2832 ( 
.A(n_2765),
.B(n_361),
.Y(n_2832)
);

NAND3xp33_ASAP7_75t_L g2833 ( 
.A(n_2774),
.B(n_362),
.C(n_363),
.Y(n_2833)
);

AOI322xp5_ASAP7_75t_L g2834 ( 
.A1(n_2798),
.A2(n_2745),
.A3(n_2776),
.B1(n_2744),
.B2(n_2763),
.C1(n_2796),
.C2(n_2758),
.Y(n_2834)
);

INVx1_ASAP7_75t_L g2835 ( 
.A(n_2803),
.Y(n_2835)
);

AOI322xp5_ASAP7_75t_L g2836 ( 
.A1(n_2799),
.A2(n_2791),
.A3(n_2793),
.B1(n_2790),
.B2(n_2777),
.C1(n_2746),
.C2(n_2782),
.Y(n_2836)
);

OAI322xp33_ASAP7_75t_L g2837 ( 
.A1(n_2823),
.A2(n_2742),
.A3(n_2769),
.B1(n_2755),
.B2(n_2766),
.C1(n_2767),
.C2(n_2797),
.Y(n_2837)
);

XNOR2xp5_ASAP7_75t_L g2838 ( 
.A(n_2802),
.B(n_2788),
.Y(n_2838)
);

OAI211xp5_ASAP7_75t_SL g2839 ( 
.A1(n_2807),
.A2(n_366),
.B(n_363),
.C(n_365),
.Y(n_2839)
);

XNOR2xp5_ASAP7_75t_L g2840 ( 
.A(n_2805),
.B(n_367),
.Y(n_2840)
);

OAI221xp5_ASAP7_75t_L g2841 ( 
.A1(n_2808),
.A2(n_2831),
.B1(n_2810),
.B2(n_2818),
.C(n_2813),
.Y(n_2841)
);

AOI322xp5_ASAP7_75t_L g2842 ( 
.A1(n_2809),
.A2(n_368),
.A3(n_369),
.B1(n_370),
.B2(n_373),
.C1(n_375),
.C2(n_379),
.Y(n_2842)
);

HB1xp67_ASAP7_75t_L g2843 ( 
.A(n_2801),
.Y(n_2843)
);

INVx1_ASAP7_75t_L g2844 ( 
.A(n_2823),
.Y(n_2844)
);

OAI221xp5_ASAP7_75t_L g2845 ( 
.A1(n_2826),
.A2(n_368),
.B1(n_380),
.B2(n_381),
.C(n_382),
.Y(n_2845)
);

NAND2xp5_ASAP7_75t_L g2846 ( 
.A(n_2811),
.B(n_380),
.Y(n_2846)
);

AOI221xp5_ASAP7_75t_L g2847 ( 
.A1(n_2829),
.A2(n_383),
.B1(n_384),
.B2(n_385),
.C(n_386),
.Y(n_2847)
);

AOI31xp33_ASAP7_75t_L g2848 ( 
.A1(n_2824),
.A2(n_2809),
.A3(n_2812),
.B(n_2833),
.Y(n_2848)
);

INVx2_ASAP7_75t_L g2849 ( 
.A(n_2832),
.Y(n_2849)
);

AOI221xp5_ASAP7_75t_L g2850 ( 
.A1(n_2814),
.A2(n_383),
.B1(n_384),
.B2(n_385),
.C(n_386),
.Y(n_2850)
);

AOI32xp33_ASAP7_75t_L g2851 ( 
.A1(n_2821),
.A2(n_387),
.A3(n_388),
.B1(n_389),
.B2(n_390),
.Y(n_2851)
);

HB1xp67_ASAP7_75t_L g2852 ( 
.A(n_2840),
.Y(n_2852)
);

OAI21xp5_ASAP7_75t_L g2853 ( 
.A1(n_2835),
.A2(n_2806),
.B(n_2827),
.Y(n_2853)
);

OAI22xp5_ASAP7_75t_SL g2854 ( 
.A1(n_2841),
.A2(n_2822),
.B1(n_2830),
.B2(n_2832),
.Y(n_2854)
);

AOI22x1_ASAP7_75t_L g2855 ( 
.A1(n_2843),
.A2(n_2816),
.B1(n_2819),
.B2(n_2800),
.Y(n_2855)
);

OAI22xp5_ASAP7_75t_L g2856 ( 
.A1(n_2845),
.A2(n_2821),
.B1(n_2828),
.B2(n_2804),
.Y(n_2856)
);

OAI21xp5_ASAP7_75t_L g2857 ( 
.A1(n_2834),
.A2(n_2838),
.B(n_2815),
.Y(n_2857)
);

INVx1_ASAP7_75t_L g2858 ( 
.A(n_2846),
.Y(n_2858)
);

INVx1_ASAP7_75t_L g2859 ( 
.A(n_2844),
.Y(n_2859)
);

NAND2xp5_ASAP7_75t_L g2860 ( 
.A(n_2851),
.B(n_2820),
.Y(n_2860)
);

OAI22xp5_ASAP7_75t_SL g2861 ( 
.A1(n_2849),
.A2(n_2820),
.B1(n_2825),
.B2(n_2817),
.Y(n_2861)
);

XNOR2x1_ASAP7_75t_L g2862 ( 
.A(n_2837),
.B(n_387),
.Y(n_2862)
);

AOI22xp5_ASAP7_75t_L g2863 ( 
.A1(n_2839),
.A2(n_388),
.B1(n_391),
.B2(n_392),
.Y(n_2863)
);

INVx2_ASAP7_75t_L g2864 ( 
.A(n_2842),
.Y(n_2864)
);

INVx1_ASAP7_75t_SL g2865 ( 
.A(n_2848),
.Y(n_2865)
);

AOI21xp5_ASAP7_75t_L g2866 ( 
.A1(n_2847),
.A2(n_391),
.B(n_393),
.Y(n_2866)
);

INVx1_ASAP7_75t_L g2867 ( 
.A(n_2854),
.Y(n_2867)
);

AOI21xp5_ASAP7_75t_SL g2868 ( 
.A1(n_2862),
.A2(n_2850),
.B(n_2836),
.Y(n_2868)
);

OAI211xp5_ASAP7_75t_L g2869 ( 
.A1(n_2853),
.A2(n_393),
.B(n_394),
.C(n_395),
.Y(n_2869)
);

OAI22xp5_ASAP7_75t_L g2870 ( 
.A1(n_2863),
.A2(n_395),
.B1(n_396),
.B2(n_397),
.Y(n_2870)
);

AO221x1_ASAP7_75t_L g2871 ( 
.A1(n_2861),
.A2(n_2856),
.B1(n_2859),
.B2(n_2864),
.C(n_2858),
.Y(n_2871)
);

OAI22xp5_ASAP7_75t_L g2872 ( 
.A1(n_2865),
.A2(n_397),
.B1(n_399),
.B2(n_400),
.Y(n_2872)
);

HB1xp67_ASAP7_75t_L g2873 ( 
.A(n_2860),
.Y(n_2873)
);

AOI21xp33_ASAP7_75t_L g2874 ( 
.A1(n_2855),
.A2(n_399),
.B(n_400),
.Y(n_2874)
);

AOI21xp5_ASAP7_75t_L g2875 ( 
.A1(n_2857),
.A2(n_401),
.B(n_402),
.Y(n_2875)
);

AOI21xp5_ASAP7_75t_L g2876 ( 
.A1(n_2866),
.A2(n_401),
.B(n_402),
.Y(n_2876)
);

HB1xp67_ASAP7_75t_L g2877 ( 
.A(n_2852),
.Y(n_2877)
);

INVx3_ASAP7_75t_L g2878 ( 
.A(n_2859),
.Y(n_2878)
);

OAI22xp33_ASAP7_75t_SL g2879 ( 
.A1(n_2865),
.A2(n_403),
.B1(n_404),
.B2(n_405),
.Y(n_2879)
);

NAND2xp5_ASAP7_75t_L g2880 ( 
.A(n_2865),
.B(n_405),
.Y(n_2880)
);

INVx2_ASAP7_75t_L g2881 ( 
.A(n_2855),
.Y(n_2881)
);

A2O1A1Ixp33_ASAP7_75t_L g2882 ( 
.A1(n_2853),
.A2(n_406),
.B(n_407),
.C(n_408),
.Y(n_2882)
);

NOR2xp67_ASAP7_75t_L g2883 ( 
.A(n_2869),
.B(n_407),
.Y(n_2883)
);

NAND2xp5_ASAP7_75t_SL g2884 ( 
.A(n_2879),
.B(n_408),
.Y(n_2884)
);

HB1xp67_ASAP7_75t_L g2885 ( 
.A(n_2878),
.Y(n_2885)
);

OAI22xp5_ASAP7_75t_SL g2886 ( 
.A1(n_2881),
.A2(n_409),
.B1(n_411),
.B2(n_412),
.Y(n_2886)
);

OAI22xp5_ASAP7_75t_L g2887 ( 
.A1(n_2867),
.A2(n_409),
.B1(n_411),
.B2(n_412),
.Y(n_2887)
);

NOR2xp33_ASAP7_75t_L g2888 ( 
.A(n_2874),
.B(n_414),
.Y(n_2888)
);

AOI21xp5_ASAP7_75t_L g2889 ( 
.A1(n_2868),
.A2(n_414),
.B(n_415),
.Y(n_2889)
);

INVx3_ASAP7_75t_L g2890 ( 
.A(n_2878),
.Y(n_2890)
);

BUFx2_ASAP7_75t_L g2891 ( 
.A(n_2882),
.Y(n_2891)
);

INVx1_ASAP7_75t_L g2892 ( 
.A(n_2880),
.Y(n_2892)
);

INVx1_ASAP7_75t_SL g2893 ( 
.A(n_2877),
.Y(n_2893)
);

CKINVDCx20_ASAP7_75t_R g2894 ( 
.A(n_2893),
.Y(n_2894)
);

HB1xp67_ASAP7_75t_L g2895 ( 
.A(n_2885),
.Y(n_2895)
);

INVx1_ASAP7_75t_L g2896 ( 
.A(n_2890),
.Y(n_2896)
);

OAI221xp5_ASAP7_75t_L g2897 ( 
.A1(n_2890),
.A2(n_2873),
.B1(n_2875),
.B2(n_2876),
.C(n_2870),
.Y(n_2897)
);

INVx1_ASAP7_75t_L g2898 ( 
.A(n_2886),
.Y(n_2898)
);

AOI22xp5_ASAP7_75t_L g2899 ( 
.A1(n_2888),
.A2(n_2871),
.B1(n_2872),
.B2(n_418),
.Y(n_2899)
);

AOI31xp33_ASAP7_75t_L g2900 ( 
.A1(n_2889),
.A2(n_416),
.A3(n_417),
.B(n_418),
.Y(n_2900)
);

XOR2xp5_ASAP7_75t_L g2901 ( 
.A(n_2894),
.B(n_2892),
.Y(n_2901)
);

AOI22xp33_ASAP7_75t_SL g2902 ( 
.A1(n_2895),
.A2(n_2891),
.B1(n_2887),
.B2(n_2883),
.Y(n_2902)
);

AOI221xp5_ASAP7_75t_L g2903 ( 
.A1(n_2897),
.A2(n_2884),
.B1(n_419),
.B2(n_420),
.C(n_421),
.Y(n_2903)
);

AOI22xp5_ASAP7_75t_L g2904 ( 
.A1(n_2899),
.A2(n_417),
.B1(n_422),
.B2(n_423),
.Y(n_2904)
);

OR2x2_ASAP7_75t_L g2905 ( 
.A(n_2896),
.B(n_423),
.Y(n_2905)
);

HB1xp67_ASAP7_75t_L g2906 ( 
.A(n_2898),
.Y(n_2906)
);

INVx1_ASAP7_75t_SL g2907 ( 
.A(n_2900),
.Y(n_2907)
);

AOI21xp33_ASAP7_75t_L g2908 ( 
.A1(n_2901),
.A2(n_424),
.B(n_425),
.Y(n_2908)
);

AOI22xp33_ASAP7_75t_L g2909 ( 
.A1(n_2906),
.A2(n_424),
.B1(n_425),
.B2(n_426),
.Y(n_2909)
);

OA22x2_ASAP7_75t_L g2910 ( 
.A1(n_2904),
.A2(n_2907),
.B1(n_2903),
.B2(n_2902),
.Y(n_2910)
);

AOI322xp5_ASAP7_75t_L g2911 ( 
.A1(n_2908),
.A2(n_2909),
.A3(n_2910),
.B1(n_2905),
.B2(n_431),
.C1(n_432),
.C2(n_433),
.Y(n_2911)
);

OAI22xp5_ASAP7_75t_L g2912 ( 
.A1(n_2911),
.A2(n_426),
.B1(n_427),
.B2(n_430),
.Y(n_2912)
);

AOI211xp5_ASAP7_75t_L g2913 ( 
.A1(n_2912),
.A2(n_427),
.B(n_430),
.C(n_433),
.Y(n_2913)
);


endmodule