module fake_jpeg_30704_n_35 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_35);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_35;

wire n_13;
wire n_21;
wire n_33;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_34;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_12;
wire n_32;
wire n_15;

NOR2xp33_ASAP7_75t_L g10 ( 
.A(n_7),
.B(n_9),
.Y(n_10)
);

BUFx6f_ASAP7_75t_L g11 ( 
.A(n_2),
.Y(n_11)
);

NAND2xp5_ASAP7_75t_L g12 ( 
.A(n_6),
.B(n_7),
.Y(n_12)
);

INVx4_ASAP7_75t_L g13 ( 
.A(n_8),
.Y(n_13)
);

INVx3_ASAP7_75t_L g14 ( 
.A(n_2),
.Y(n_14)
);

AOI22xp5_ASAP7_75t_SL g15 ( 
.A1(n_14),
.A2(n_13),
.B1(n_12),
.B2(n_11),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_15),
.B(n_16),
.Y(n_22)
);

INVxp33_ASAP7_75t_L g16 ( 
.A(n_13),
.Y(n_16)
);

AND2x6_ASAP7_75t_L g17 ( 
.A(n_12),
.B(n_0),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g24 ( 
.A(n_17),
.B(n_18),
.Y(n_24)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_19),
.B(n_20),
.Y(n_25)
);

INVx2_ASAP7_75t_SL g20 ( 
.A(n_13),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_20),
.B(n_11),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_21),
.B(n_10),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_16),
.Y(n_23)
);

AND2x2_ASAP7_75t_SL g26 ( 
.A(n_23),
.B(n_0),
.Y(n_26)
);

INVxp67_ASAP7_75t_L g32 ( 
.A(n_26),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_L g27 ( 
.A1(n_22),
.A2(n_10),
.B1(n_3),
.B2(n_4),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_27),
.B(n_29),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_SL g31 ( 
.A(n_28),
.B(n_25),
.Y(n_31)
);

AOI21xp5_ASAP7_75t_SL g29 ( 
.A1(n_21),
.A2(n_1),
.B(n_3),
.Y(n_29)
);

AND2x2_ASAP7_75t_L g34 ( 
.A(n_31),
.B(n_5),
.Y(n_34)
);

AOI322xp5_ASAP7_75t_L g33 ( 
.A1(n_30),
.A2(n_24),
.A3(n_28),
.B1(n_5),
.B2(n_6),
.C1(n_1),
.C2(n_4),
.Y(n_33)
);

OAI21xp5_ASAP7_75t_SL g35 ( 
.A1(n_33),
.A2(n_34),
.B(n_32),
.Y(n_35)
);


endmodule