module real_jpeg_22569_n_17 (n_8, n_0, n_2, n_341, n_10, n_9, n_12, n_6, n_340, n_11, n_14, n_7, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_17);

input n_8;
input n_0;
input n_2;
input n_341;
input n_10;
input n_9;
input n_12;
input n_6;
input n_340;
input n_11;
input n_14;
input n_7;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_17;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_338;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_18;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_330;
wire n_298;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_0),
.A2(n_64),
.B1(n_65),
.B2(n_126),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_0),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_L g164 ( 
.A1(n_0),
.A2(n_46),
.B1(n_48),
.B2(n_126),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_SL g220 ( 
.A1(n_0),
.A2(n_31),
.B1(n_32),
.B2(n_126),
.Y(n_220)
);

AOI22xp33_ASAP7_75t_SL g263 ( 
.A1(n_0),
.A2(n_23),
.B1(n_25),
.B2(n_126),
.Y(n_263)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_1),
.A2(n_23),
.B1(n_25),
.B2(n_57),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_1),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_1),
.A2(n_31),
.B1(n_32),
.B2(n_57),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g210 ( 
.A1(n_1),
.A2(n_57),
.B1(n_64),
.B2(n_65),
.Y(n_210)
);

AOI22xp33_ASAP7_75t_L g254 ( 
.A1(n_1),
.A2(n_46),
.B1(n_48),
.B2(n_57),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_L g33 ( 
.A1(n_2),
.A2(n_23),
.B1(n_25),
.B2(n_34),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_2),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_2),
.A2(n_31),
.B1(n_32),
.B2(n_34),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_2),
.A2(n_34),
.B1(n_46),
.B2(n_48),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g252 ( 
.A1(n_2),
.A2(n_34),
.B1(n_64),
.B2(n_65),
.Y(n_252)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_3),
.A2(n_46),
.B1(n_48),
.B2(n_121),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_3),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_3),
.A2(n_64),
.B1(n_65),
.B2(n_121),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_SL g185 ( 
.A1(n_3),
.A2(n_31),
.B1(n_32),
.B2(n_121),
.Y(n_185)
);

AOI22xp33_ASAP7_75t_SL g234 ( 
.A1(n_3),
.A2(n_23),
.B1(n_25),
.B2(n_121),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g21 ( 
.A1(n_4),
.A2(n_22),
.B1(n_23),
.B2(n_25),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_4),
.Y(n_22)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_4),
.A2(n_22),
.B1(n_31),
.B2(n_32),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_4),
.A2(n_22),
.B1(n_64),
.B2(n_65),
.Y(n_243)
);

AOI22xp33_ASAP7_75t_SL g286 ( 
.A1(n_4),
.A2(n_22),
.B1(n_46),
.B2(n_48),
.Y(n_286)
);

BUFx16f_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_6),
.A2(n_23),
.B1(n_25),
.B2(n_90),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_6),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_6),
.A2(n_64),
.B1(n_65),
.B2(n_90),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_L g217 ( 
.A1(n_6),
.A2(n_46),
.B1(n_48),
.B2(n_90),
.Y(n_217)
);

OAI22xp33_ASAP7_75t_SL g260 ( 
.A1(n_6),
.A2(n_31),
.B1(n_32),
.B2(n_90),
.Y(n_260)
);

A2O1A1O1Ixp25_ASAP7_75t_L g105 ( 
.A1(n_7),
.A2(n_48),
.B(n_60),
.C(n_106),
.D(n_107),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_7),
.B(n_48),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_7),
.B(n_45),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_7),
.Y(n_145)
);

OAI21xp33_ASAP7_75t_L g151 ( 
.A1(n_7),
.A2(n_127),
.B(n_129),
.Y(n_151)
);

A2O1A1O1Ixp25_ASAP7_75t_L g165 ( 
.A1(n_7),
.A2(n_31),
.B(n_42),
.C(n_166),
.D(n_167),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_7),
.B(n_31),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_7),
.B(n_35),
.Y(n_189)
);

AOI21xp33_ASAP7_75t_L g205 ( 
.A1(n_7),
.A2(n_32),
.B(n_206),
.Y(n_205)
);

OAI22xp33_ASAP7_75t_SL g223 ( 
.A1(n_7),
.A2(n_23),
.B1(n_25),
.B2(n_145),
.Y(n_223)
);

INVx6_ASAP7_75t_L g128 ( 
.A(n_8),
.Y(n_128)
);

INVx8_ASAP7_75t_L g147 ( 
.A(n_8),
.Y(n_147)
);

BUFx10_ASAP7_75t_L g64 ( 
.A(n_9),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_10),
.A2(n_23),
.B1(n_25),
.B2(n_55),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_10),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_10),
.A2(n_55),
.B1(n_64),
.B2(n_65),
.Y(n_191)
);

AOI22xp33_ASAP7_75t_SL g245 ( 
.A1(n_10),
.A2(n_46),
.B1(n_48),
.B2(n_55),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_L g279 ( 
.A1(n_10),
.A2(n_31),
.B1(n_32),
.B2(n_55),
.Y(n_279)
);

BUFx12_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

AOI22xp33_ASAP7_75t_L g108 ( 
.A1(n_12),
.A2(n_46),
.B1(n_48),
.B2(n_109),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_12),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_12),
.A2(n_64),
.B1(n_65),
.B2(n_109),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_L g168 ( 
.A1(n_12),
.A2(n_31),
.B1(n_32),
.B2(n_109),
.Y(n_168)
);

OAI22xp33_ASAP7_75t_SL g226 ( 
.A1(n_12),
.A2(n_23),
.B1(n_25),
.B2(n_109),
.Y(n_226)
);

INVx13_ASAP7_75t_L g43 ( 
.A(n_13),
.Y(n_43)
);

INVx13_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_L g30 ( 
.A1(n_14),
.A2(n_28),
.B1(n_31),
.B2(n_32),
.Y(n_30)
);

INVx11_ASAP7_75t_L g61 ( 
.A(n_15),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_16),
.Y(n_46)
);

XNOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_76),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_74),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_36),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_20),
.B(n_36),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_26),
.B1(n_33),
.B2(n_35),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_21),
.A2(n_26),
.B1(n_35),
.B2(n_70),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_23),
.Y(n_25)
);

A2O1A1Ixp33_ASAP7_75t_L g27 ( 
.A1(n_23),
.A2(n_28),
.B(n_29),
.C(n_30),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_23),
.B(n_28),
.Y(n_29)
);

A2O1A1Ixp33_ASAP7_75t_L g204 ( 
.A1(n_23),
.A2(n_28),
.B(n_145),
.C(n_205),
.Y(n_204)
);

BUFx2_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

AOI21xp5_ASAP7_75t_L g222 ( 
.A1(n_26),
.A2(n_223),
.B(n_224),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_26),
.B(n_226),
.Y(n_235)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_27),
.A2(n_30),
.B1(n_54),
.B2(n_56),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_27),
.A2(n_30),
.B1(n_54),
.B2(n_89),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_27),
.A2(n_30),
.B1(n_234),
.B2(n_263),
.Y(n_262)
);

OAI21xp5_ASAP7_75t_SL g281 ( 
.A1(n_27),
.A2(n_225),
.B(n_263),
.Y(n_281)
);

INVx4_ASAP7_75t_L g206 ( 
.A(n_28),
.Y(n_206)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_30),
.Y(n_35)
);

OAI21xp33_ASAP7_75t_L g233 ( 
.A1(n_30),
.A2(n_234),
.B(n_235),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_L g305 ( 
.A1(n_30),
.A2(n_89),
.B(n_235),
.Y(n_305)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

O2A1O1Ixp33_ASAP7_75t_SL g42 ( 
.A1(n_32),
.A2(n_43),
.B(n_44),
.C(n_45),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_32),
.B(n_43),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_35),
.B(n_226),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g36 ( 
.A(n_37),
.B(n_69),
.C(n_71),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_37),
.A2(n_38),
.B1(n_79),
.B2(n_81),
.Y(n_78)
);

CKINVDCx14_ASAP7_75t_R g37 ( 
.A(n_38),
.Y(n_37)
);

MAJIxp5_ASAP7_75t_L g38 ( 
.A(n_39),
.B(n_52),
.C(n_58),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_39),
.A2(n_40),
.B1(n_58),
.B2(n_87),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_40),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_SL g40 ( 
.A1(n_41),
.A2(n_49),
.B1(n_50),
.B2(n_51),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_41),
.A2(n_49),
.B1(n_50),
.B2(n_94),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_41),
.A2(n_50),
.B1(n_185),
.B2(n_220),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_L g237 ( 
.A1(n_41),
.A2(n_220),
.B(n_238),
.Y(n_237)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

OAI21xp5_ASAP7_75t_SL g72 ( 
.A1(n_42),
.A2(n_45),
.B(n_73),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_42),
.B(n_187),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_42),
.A2(n_45),
.B1(n_260),
.B2(n_279),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_42),
.A2(n_45),
.B1(n_95),
.B2(n_279),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_L g45 ( 
.A1(n_43),
.A2(n_46),
.B1(n_47),
.B2(n_48),
.Y(n_45)
);

INVx11_ASAP7_75t_L g47 ( 
.A(n_43),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_44),
.Y(n_174)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_45),
.Y(n_50)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_46),
.Y(n_48)
);

O2A1O1Ixp33_ASAP7_75t_L g60 ( 
.A1(n_46),
.A2(n_61),
.B(n_62),
.C(n_63),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_46),
.B(n_61),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_46),
.B(n_47),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_48),
.A2(n_166),
.B1(n_173),
.B2(n_174),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_50),
.B(n_168),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_L g184 ( 
.A1(n_50),
.A2(n_185),
.B(n_186),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_L g258 ( 
.A1(n_50),
.A2(n_186),
.B(n_259),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_51),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_52),
.A2(n_53),
.B1(n_85),
.B2(n_86),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_53),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_56),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_58),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g326 ( 
.A1(n_58),
.A2(n_87),
.B1(n_92),
.B2(n_93),
.Y(n_326)
);

AOI21xp5_ASAP7_75t_SL g58 ( 
.A1(n_59),
.A2(n_67),
.B(n_68),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_59),
.A2(n_67),
.B1(n_120),
.B2(n_164),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_SL g195 ( 
.A1(n_59),
.A2(n_164),
.B(n_196),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g244 ( 
.A1(n_59),
.A2(n_67),
.B1(n_217),
.B2(n_245),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_L g253 ( 
.A1(n_59),
.A2(n_67),
.B1(n_245),
.B2(n_254),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_59),
.A2(n_67),
.B1(n_254),
.B2(n_286),
.Y(n_285)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_60),
.B(n_123),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_60),
.A2(n_63),
.B1(n_295),
.B2(n_296),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_61),
.A2(n_64),
.B1(n_65),
.B2(n_66),
.Y(n_63)
);

CKINVDCx9p33_ASAP7_75t_R g66 ( 
.A(n_61),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_61),
.B(n_65),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_62),
.A2(n_64),
.B1(n_112),
.B2(n_113),
.Y(n_111)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_63),
.Y(n_67)
);

INVx13_ASAP7_75t_L g65 ( 
.A(n_64),
.Y(n_65)
);

NAND2x1_ASAP7_75t_SL g127 ( 
.A(n_64),
.B(n_128),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_65),
.B(n_153),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_67),
.B(n_108),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_L g119 ( 
.A1(n_67),
.A2(n_120),
.B(n_122),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g144 ( 
.A(n_67),
.B(n_145),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_L g216 ( 
.A1(n_67),
.A2(n_122),
.B(n_217),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_68),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_69),
.A2(n_71),
.B1(n_72),
.B2(n_80),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_69),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_72),
.Y(n_71)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

AOI21xp5_ASAP7_75t_L g76 ( 
.A1(n_77),
.A2(n_96),
.B(n_338),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_82),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_78),
.B(n_82),
.Y(n_338)
);

CKINVDCx16_ASAP7_75t_R g81 ( 
.A(n_79),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_88),
.C(n_91),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g330 ( 
.A1(n_83),
.A2(n_84),
.B1(n_88),
.B2(n_324),
.Y(n_330)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_87),
.B(n_88),
.C(n_92),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g323 ( 
.A1(n_88),
.A2(n_324),
.B1(n_325),
.B2(n_326),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_88),
.Y(n_324)
);

XOR2xp5_ASAP7_75t_L g329 ( 
.A(n_91),
.B(n_330),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_93),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_95),
.Y(n_94)
);

OAI321xp33_ASAP7_75t_L g96 ( 
.A1(n_97),
.A2(n_321),
.A3(n_331),
.B1(n_336),
.B2(n_337),
.C(n_340),
.Y(n_96)
);

AOI321xp33_ASAP7_75t_L g97 ( 
.A1(n_98),
.A2(n_271),
.A3(n_309),
.B1(n_315),
.B2(n_320),
.C(n_341),
.Y(n_97)
);

NOR3xp33_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_228),
.C(n_267),
.Y(n_98)
);

AOI21x1_ASAP7_75t_L g99 ( 
.A1(n_100),
.A2(n_198),
.B(n_227),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_SL g100 ( 
.A1(n_101),
.A2(n_179),
.B(n_197),
.Y(n_100)
);

AOI21xp5_ASAP7_75t_L g101 ( 
.A1(n_102),
.A2(n_158),
.B(n_178),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_SL g102 ( 
.A1(n_103),
.A2(n_133),
.B(n_157),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_114),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_104),
.B(n_114),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_105),
.B(n_110),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_105),
.A2(n_110),
.B1(n_111),
.B2(n_141),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_105),
.Y(n_141)
);

CKINVDCx16_ASAP7_75t_R g113 ( 
.A(n_106),
.Y(n_113)
);

CKINVDCx14_ASAP7_75t_R g196 ( 
.A(n_107),
.Y(n_196)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_108),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_111),
.Y(n_110)
);

XNOR2xp5_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_124),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_116),
.A2(n_117),
.B1(n_118),
.B2(n_119),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_116),
.B(n_119),
.C(n_124),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_117),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_119),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_SL g124 ( 
.A1(n_125),
.A2(n_127),
.B(n_129),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_125),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_127),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_127),
.B(n_131),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_127),
.A2(n_128),
.B1(n_209),
.B2(n_210),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g242 ( 
.A1(n_127),
.A2(n_154),
.B1(n_210),
.B2(n_243),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_L g251 ( 
.A1(n_127),
.A2(n_147),
.B1(n_243),
.B2(n_252),
.Y(n_251)
);

AOI21xp5_ASAP7_75t_L g284 ( 
.A1(n_127),
.A2(n_128),
.B(n_252),
.Y(n_284)
);

INVx5_ASAP7_75t_L g132 ( 
.A(n_128),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_130),
.B(n_132),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_131),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_132),
.A2(n_136),
.B1(n_138),
.B2(n_139),
.Y(n_135)
);

INVx4_ASAP7_75t_L g154 ( 
.A(n_132),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_L g175 ( 
.A1(n_132),
.A2(n_149),
.B(n_176),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_132),
.A2(n_138),
.B1(n_176),
.B2(n_191),
.Y(n_190)
);

AOI21xp5_ASAP7_75t_L g133 ( 
.A1(n_134),
.A2(n_142),
.B(n_156),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_140),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g156 ( 
.A(n_135),
.B(n_140),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_137),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_L g146 ( 
.A1(n_137),
.A2(n_147),
.B(n_148),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_SL g142 ( 
.A1(n_143),
.A2(n_150),
.B(n_155),
.Y(n_142)
);

NOR2x1_ASAP7_75t_R g143 ( 
.A(n_144),
.B(n_146),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_144),
.B(n_146),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_145),
.B(n_154),
.Y(n_153)
);

INVxp67_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_151),
.B(n_152),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_160),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_SL g178 ( 
.A(n_159),
.B(n_160),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_161),
.A2(n_162),
.B1(n_171),
.B2(n_177),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_163),
.A2(n_165),
.B1(n_169),
.B2(n_170),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_163),
.Y(n_170)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_165),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_165),
.B(n_170),
.C(n_177),
.Y(n_180)
);

CKINVDCx16_ASAP7_75t_R g238 ( 
.A(n_167),
.Y(n_238)
);

INVxp67_ASAP7_75t_L g187 ( 
.A(n_168),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_171),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_175),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_172),
.B(n_175),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_181),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_180),
.B(n_181),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_193),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_182),
.B(n_194),
.C(n_195),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_183),
.A2(n_184),
.B1(n_188),
.B2(n_192),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_183),
.B(n_189),
.C(n_190),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_184),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_188),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_190),
.Y(n_188)
);

INVxp67_ASAP7_75t_L g209 ( 
.A(n_191),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_195),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_200),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_199),
.B(n_200),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_214),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_202),
.A2(n_211),
.B1(n_212),
.B2(n_213),
.Y(n_201)
);

CKINVDCx16_ASAP7_75t_R g212 ( 
.A(n_202),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_202),
.B(n_213),
.C(n_214),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_203),
.A2(n_204),
.B1(n_207),
.B2(n_208),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_203),
.B(n_208),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_204),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_208),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_211),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_222),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_216),
.A2(n_218),
.B1(n_219),
.B2(n_221),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_216),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_218),
.B(n_221),
.C(n_222),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_219),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_225),
.Y(n_224)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

AOI21xp33_ASAP7_75t_L g316 ( 
.A1(n_229),
.A2(n_317),
.B(n_318),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_247),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_230),
.B(n_247),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_241),
.C(n_246),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_231),
.B(n_270),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_240),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_233),
.A2(n_236),
.B1(n_237),
.B2(n_239),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_233),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_236),
.B(n_239),
.C(n_240),
.Y(n_265)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_241),
.B(n_246),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_244),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_242),
.B(n_244),
.Y(n_256)
);

AOI22xp33_ASAP7_75t_SL g247 ( 
.A1(n_248),
.A2(n_249),
.B1(n_265),
.B2(n_266),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_255),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_250),
.B(n_255),
.C(n_266),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_253),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_251),
.B(n_253),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_257),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_256),
.B(n_261),
.C(n_264),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_258),
.A2(n_261),
.B1(n_262),
.B2(n_264),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_258),
.Y(n_264)
);

CKINVDCx16_ASAP7_75t_R g259 ( 
.A(n_260),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_262),
.Y(n_261)
);

CKINVDCx16_ASAP7_75t_R g266 ( 
.A(n_265),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_268),
.B(n_269),
.Y(n_267)
);

AND2x2_ASAP7_75t_L g317 ( 
.A(n_268),
.B(n_269),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_289),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_SL g320 ( 
.A(n_272),
.B(n_289),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_273),
.B(n_282),
.C(n_288),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_SL g313 ( 
.A1(n_273),
.A2(n_274),
.B1(n_282),
.B2(n_314),
.Y(n_313)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_275),
.B(n_276),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_275),
.B(n_278),
.C(n_280),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_L g276 ( 
.A1(n_277),
.A2(n_278),
.B1(n_280),
.B2(n_281),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_278),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_281),
.Y(n_280)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_282),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_L g282 ( 
.A1(n_283),
.A2(n_284),
.B1(n_285),
.B2(n_287),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_283),
.A2(n_284),
.B1(n_304),
.B2(n_305),
.Y(n_303)
);

OAI21xp5_ASAP7_75t_L g328 ( 
.A1(n_283),
.A2(n_301),
.B(n_305),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_284),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_284),
.B(n_285),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_285),
.Y(n_287)
);

CKINVDCx16_ASAP7_75t_R g295 ( 
.A(n_286),
.Y(n_295)
);

XOR2xp5_ASAP7_75t_L g312 ( 
.A(n_288),
.B(n_313),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_290),
.A2(n_291),
.B1(n_307),
.B2(n_308),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_L g291 ( 
.A1(n_292),
.A2(n_293),
.B1(n_299),
.B2(n_300),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_292),
.B(n_300),
.C(n_308),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_293),
.Y(n_292)
);

OAI21xp5_ASAP7_75t_L g293 ( 
.A1(n_294),
.A2(n_297),
.B(n_298),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_294),
.B(n_297),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_298),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_SL g334 ( 
.A1(n_298),
.A2(n_323),
.B1(n_327),
.B2(n_335),
.Y(n_334)
);

CKINVDCx16_ASAP7_75t_R g299 ( 
.A(n_300),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_301),
.A2(n_302),
.B1(n_303),
.B2(n_306),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_303),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_305),
.Y(n_304)
);

CKINVDCx16_ASAP7_75t_R g308 ( 
.A(n_307),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

OAI21xp5_ASAP7_75t_SL g315 ( 
.A1(n_310),
.A2(n_316),
.B(n_319),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_311),
.B(n_312),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_SL g319 ( 
.A(n_311),
.B(n_312),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_322),
.B(n_329),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_322),
.B(n_329),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_323),
.B(n_327),
.C(n_328),
.Y(n_322)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_323),
.Y(n_335)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

XNOR2xp5_ASAP7_75t_L g333 ( 
.A(n_328),
.B(n_334),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_332),
.B(n_333),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_SL g336 ( 
.A(n_332),
.B(n_333),
.Y(n_336)
);


endmodule