module fake_jpeg_10725_n_392 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_392);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_392;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_19;
wire n_182;
wire n_385;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_11),
.Y(n_16)
);

INVx6_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_5),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

BUFx10_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_13),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_15),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_12),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_1),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_0),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_13),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_4),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_7),
.Y(n_36)
);

INVx1_ASAP7_75t_SL g37 ( 
.A(n_8),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_7),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_9),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_12),
.Y(n_40)
);

INVx13_ASAP7_75t_L g41 ( 
.A(n_1),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_7),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_3),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_9),
.B(n_10),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_31),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_45),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_44),
.B(n_16),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_46),
.B(n_73),
.Y(n_104)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_38),
.Y(n_47)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_47),
.Y(n_100)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_38),
.Y(n_48)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_48),
.Y(n_107)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_21),
.Y(n_49)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_49),
.Y(n_95)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_50),
.Y(n_109)
);

BUFx4f_ASAP7_75t_L g51 ( 
.A(n_23),
.Y(n_51)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_51),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_23),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_52),
.B(n_56),
.Y(n_108)
);

INVx11_ASAP7_75t_L g53 ( 
.A(n_23),
.Y(n_53)
);

CKINVDCx16_ASAP7_75t_R g118 ( 
.A(n_53),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_31),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_54),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_31),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_55),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g56 ( 
.A(n_44),
.B(n_14),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_22),
.Y(n_57)
);

BUFx12f_ASAP7_75t_L g93 ( 
.A(n_57),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_23),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_58),
.B(n_69),
.Y(n_110)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_27),
.Y(n_59)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_59),
.Y(n_106)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_22),
.Y(n_60)
);

INVx1_ASAP7_75t_SL g123 ( 
.A(n_60),
.Y(n_123)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_43),
.Y(n_61)
);

INVx6_ASAP7_75t_L g98 ( 
.A(n_61),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_17),
.B(n_0),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_62),
.B(n_71),
.Y(n_115)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_22),
.Y(n_63)
);

INVx5_ASAP7_75t_L g89 ( 
.A(n_63),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_31),
.Y(n_64)
);

INVx6_ASAP7_75t_L g128 ( 
.A(n_64),
.Y(n_128)
);

INVx11_ASAP7_75t_L g65 ( 
.A(n_23),
.Y(n_65)
);

INVx5_ASAP7_75t_L g91 ( 
.A(n_65),
.Y(n_91)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_27),
.Y(n_66)
);

INVx2_ASAP7_75t_SL g99 ( 
.A(n_66),
.Y(n_99)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_35),
.Y(n_67)
);

INVx5_ASAP7_75t_L g114 ( 
.A(n_67),
.Y(n_114)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_35),
.Y(n_68)
);

INVx5_ASAP7_75t_L g119 ( 
.A(n_68),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_23),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_39),
.Y(n_70)
);

INVx5_ASAP7_75t_L g121 ( 
.A(n_70),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_17),
.B(n_0),
.Y(n_71)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_36),
.Y(n_72)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_72),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_16),
.B(n_14),
.Y(n_73)
);

BUFx10_ASAP7_75t_L g74 ( 
.A(n_41),
.Y(n_74)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_74),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_39),
.Y(n_75)
);

INVx5_ASAP7_75t_L g122 ( 
.A(n_75),
.Y(n_122)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_35),
.Y(n_76)
);

HB1xp67_ASAP7_75t_L g85 ( 
.A(n_76),
.Y(n_85)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_39),
.Y(n_77)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_77),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_24),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_78),
.B(n_25),
.Y(n_90)
);

BUFx12f_ASAP7_75t_L g79 ( 
.A(n_27),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g112 ( 
.A(n_79),
.B(n_81),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_39),
.Y(n_80)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_80),
.Y(n_124)
);

BUFx12f_ASAP7_75t_L g81 ( 
.A(n_28),
.Y(n_81)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_21),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_82),
.B(n_25),
.Y(n_127)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_36),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_83),
.B(n_36),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_63),
.A2(n_37),
.B1(n_28),
.B2(n_17),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g173 ( 
.A1(n_86),
.A2(n_97),
.B1(n_102),
.B2(n_2),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_62),
.A2(n_71),
.B1(n_47),
.B2(n_48),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_87),
.A2(n_103),
.B1(n_113),
.B2(n_125),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_90),
.B(n_101),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_61),
.A2(n_19),
.B1(n_42),
.B2(n_43),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_92),
.A2(n_96),
.B1(n_129),
.B2(n_32),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_L g96 ( 
.A1(n_45),
.A2(n_19),
.B1(n_18),
.B2(n_32),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_67),
.A2(n_37),
.B1(n_28),
.B2(n_43),
.Y(n_97)
);

OR2x2_ASAP7_75t_L g101 ( 
.A(n_74),
.B(n_29),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_68),
.A2(n_37),
.B1(n_42),
.B2(n_43),
.Y(n_102)
);

OAI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_54),
.A2(n_19),
.B1(n_42),
.B2(n_29),
.Y(n_103)
);

HAxp5_ASAP7_75t_SL g111 ( 
.A(n_74),
.B(n_41),
.CON(n_111),
.SN(n_111)
);

OR2x4_ASAP7_75t_L g154 ( 
.A(n_111),
.B(n_105),
.Y(n_154)
);

OAI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_55),
.A2(n_19),
.B1(n_42),
.B2(n_26),
.Y(n_113)
);

OAI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_64),
.A2(n_20),
.B1(n_26),
.B2(n_30),
.Y(n_125)
);

AND2x2_ASAP7_75t_L g152 ( 
.A(n_126),
.B(n_81),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_127),
.B(n_34),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_70),
.A2(n_30),
.B1(n_40),
.B2(n_24),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_50),
.B(n_40),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_130),
.B(n_34),
.Y(n_144)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_94),
.Y(n_131)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_131),
.Y(n_200)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_112),
.Y(n_132)
);

CKINVDCx11_ASAP7_75t_R g191 ( 
.A(n_132),
.Y(n_191)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_94),
.Y(n_133)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_133),
.Y(n_213)
);

BUFx3_ASAP7_75t_L g134 ( 
.A(n_93),
.Y(n_134)
);

INVx5_ASAP7_75t_L g196 ( 
.A(n_134),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_115),
.B(n_20),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_135),
.B(n_145),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_87),
.B(n_83),
.C(n_72),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_136),
.B(n_138),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_92),
.A2(n_102),
.B1(n_97),
.B2(n_86),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_L g197 ( 
.A1(n_137),
.A2(n_114),
.B1(n_89),
.B2(n_122),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_95),
.B(n_66),
.C(n_59),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_109),
.Y(n_139)
);

INVx1_ASAP7_75t_SL g214 ( 
.A(n_139),
.Y(n_214)
);

CKINVDCx16_ASAP7_75t_R g141 ( 
.A(n_112),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_141),
.B(n_143),
.Y(n_179)
);

OAI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_101),
.A2(n_80),
.B1(n_75),
.B2(n_74),
.Y(n_142)
);

OAI22xp33_ASAP7_75t_SL g185 ( 
.A1(n_142),
.A2(n_88),
.B1(n_120),
.B2(n_91),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_144),
.B(n_150),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_100),
.B(n_18),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_116),
.Y(n_146)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_146),
.Y(n_211)
);

A2O1A1Ixp33_ASAP7_75t_L g147 ( 
.A1(n_108),
.A2(n_65),
.B(n_53),
.C(n_41),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_147),
.B(n_149),
.Y(n_188)
);

AND2x2_ASAP7_75t_L g205 ( 
.A(n_148),
.B(n_152),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_107),
.B(n_33),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_104),
.B(n_81),
.Y(n_150)
);

A2O1A1Ixp33_ASAP7_75t_L g151 ( 
.A1(n_111),
.A2(n_33),
.B(n_13),
.C(n_14),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_151),
.B(n_161),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_110),
.B(n_79),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_153),
.B(n_158),
.Y(n_212)
);

CKINVDCx16_ASAP7_75t_R g189 ( 
.A(n_154),
.Y(n_189)
);

AOI32xp33_ASAP7_75t_L g155 ( 
.A1(n_99),
.A2(n_60),
.A3(n_79),
.B1(n_36),
.B2(n_51),
.Y(n_155)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_155),
.B(n_174),
.Y(n_199)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_106),
.Y(n_156)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_156),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_85),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_157),
.B(n_170),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_126),
.B(n_11),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_99),
.B(n_10),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_159),
.B(n_163),
.Y(n_217)
);

INVx13_ASAP7_75t_L g160 ( 
.A(n_105),
.Y(n_160)
);

INVx3_ASAP7_75t_SL g182 ( 
.A(n_160),
.Y(n_182)
);

A2O1A1Ixp33_ASAP7_75t_L g161 ( 
.A1(n_124),
.A2(n_10),
.B(n_51),
.C(n_60),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_98),
.B(n_0),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_162),
.B(n_164),
.Y(n_193)
);

NOR2x1_ASAP7_75t_L g163 ( 
.A(n_93),
.B(n_76),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_98),
.B(n_1),
.Y(n_164)
);

BUFx2_ASAP7_75t_L g165 ( 
.A(n_89),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g201 ( 
.A(n_165),
.Y(n_201)
);

INVx5_ASAP7_75t_L g166 ( 
.A(n_93),
.Y(n_166)
);

INVx3_ASAP7_75t_L g183 ( 
.A(n_166),
.Y(n_183)
);

INVx8_ASAP7_75t_L g167 ( 
.A(n_84),
.Y(n_167)
);

INVx4_ASAP7_75t_L g180 ( 
.A(n_167),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_128),
.A2(n_77),
.B1(n_57),
.B2(n_3),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_168),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_117),
.B(n_106),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_169),
.B(n_175),
.Y(n_195)
);

BUFx12_ASAP7_75t_L g170 ( 
.A(n_123),
.Y(n_170)
);

BUFx12_ASAP7_75t_L g171 ( 
.A(n_123),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_171),
.B(n_119),
.Y(n_184)
);

AND2x6_ASAP7_75t_L g172 ( 
.A(n_118),
.B(n_1),
.Y(n_172)
);

AND2x6_ASAP7_75t_L g198 ( 
.A(n_172),
.B(n_2),
.Y(n_198)
);

AOI21xp5_ASAP7_75t_L g215 ( 
.A1(n_173),
.A2(n_8),
.B(n_9),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_84),
.B(n_2),
.C(n_3),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_121),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_176),
.A2(n_128),
.B1(n_120),
.B2(n_88),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_177),
.A2(n_185),
.B1(n_187),
.B2(n_210),
.Y(n_226)
);

INVxp67_ASAP7_75t_L g251 ( 
.A(n_184),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_176),
.A2(n_121),
.B1(n_122),
.B2(n_119),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_140),
.B(n_114),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_SL g234 ( 
.A(n_190),
.B(n_202),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_197),
.A2(n_132),
.B1(n_169),
.B2(n_138),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_198),
.B(n_206),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_135),
.B(n_91),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_162),
.B(n_3),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_203),
.B(n_204),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_164),
.B(n_4),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_157),
.B(n_4),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_145),
.B(n_6),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_207),
.B(n_208),
.Y(n_235)
);

AND2x6_ASAP7_75t_L g208 ( 
.A(n_147),
.B(n_6),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_149),
.B(n_6),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_209),
.B(n_194),
.Y(n_236)
);

AND2x2_ASAP7_75t_L g252 ( 
.A(n_215),
.B(n_192),
.Y(n_252)
);

OA22x2_ASAP7_75t_L g218 ( 
.A1(n_189),
.A2(n_154),
.B1(n_137),
.B2(n_172),
.Y(n_218)
);

AND2x2_ASAP7_75t_L g257 ( 
.A(n_218),
.B(n_233),
.Y(n_257)
);

AO22x1_ASAP7_75t_L g219 ( 
.A1(n_189),
.A2(n_163),
.B1(n_161),
.B2(n_155),
.Y(n_219)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_219),
.Y(n_258)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_195),
.Y(n_220)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_220),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_221),
.A2(n_243),
.B1(n_224),
.B2(n_220),
.Y(n_278)
);

FAx1_ASAP7_75t_SL g222 ( 
.A(n_178),
.B(n_136),
.CI(n_151),
.CON(n_222),
.SN(n_222)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_222),
.B(n_230),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_186),
.B(n_152),
.C(n_139),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_223),
.B(n_199),
.C(n_178),
.Y(n_255)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_195),
.Y(n_224)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_224),
.Y(n_270)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_200),
.Y(n_225)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_225),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_205),
.A2(n_148),
.B1(n_168),
.B2(n_152),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_227),
.A2(n_232),
.B1(n_247),
.B2(n_188),
.Y(n_254)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_200),
.Y(n_230)
);

INVx3_ASAP7_75t_L g231 ( 
.A(n_180),
.Y(n_231)
);

HB1xp67_ASAP7_75t_L g269 ( 
.A(n_231),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_205),
.A2(n_174),
.B1(n_146),
.B2(n_156),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_213),
.Y(n_233)
);

INVxp67_ASAP7_75t_L g276 ( 
.A(n_236),
.Y(n_276)
);

OR2x2_ASAP7_75t_L g237 ( 
.A(n_188),
.B(n_131),
.Y(n_237)
);

OAI21xp5_ASAP7_75t_L g268 ( 
.A1(n_237),
.A2(n_252),
.B(n_204),
.Y(n_268)
);

AO22x1_ASAP7_75t_SL g238 ( 
.A1(n_205),
.A2(n_133),
.B1(n_175),
.B2(n_167),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_238),
.B(n_242),
.Y(n_262)
);

AOI21xp5_ASAP7_75t_L g239 ( 
.A1(n_192),
.A2(n_166),
.B(n_165),
.Y(n_239)
);

AOI21xp5_ASAP7_75t_L g253 ( 
.A1(n_239),
.A2(n_201),
.B(n_191),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_179),
.B(n_134),
.Y(n_240)
);

CKINVDCx14_ASAP7_75t_R g260 ( 
.A(n_240),
.Y(n_260)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_213),
.Y(n_241)
);

AND2x2_ASAP7_75t_L g267 ( 
.A(n_241),
.B(n_244),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_193),
.B(n_160),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_181),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_243),
.B(n_245),
.Y(n_280)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_211),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_211),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_212),
.B(n_170),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_246),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_177),
.A2(n_170),
.B1(n_171),
.B2(n_187),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_216),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_248),
.B(n_249),
.Y(n_282)
);

NOR2x1_ASAP7_75t_R g249 ( 
.A(n_186),
.B(n_171),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_216),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_250),
.B(n_214),
.Y(n_283)
);

OAI21xp5_ASAP7_75t_SL g295 ( 
.A1(n_253),
.A2(n_256),
.B(n_263),
.Y(n_295)
);

INVxp67_ASAP7_75t_L g289 ( 
.A(n_254),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_255),
.B(n_259),
.C(n_251),
.Y(n_293)
);

AOI21xp5_ASAP7_75t_L g256 ( 
.A1(n_239),
.A2(n_215),
.B(n_199),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_223),
.B(n_193),
.Y(n_259)
);

AND2x2_ASAP7_75t_SL g261 ( 
.A(n_249),
.B(n_191),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_SL g291 ( 
.A(n_261),
.B(n_268),
.Y(n_291)
);

AOI21xp5_ASAP7_75t_L g263 ( 
.A1(n_252),
.A2(n_217),
.B(n_208),
.Y(n_263)
);

AOI21xp5_ASAP7_75t_L g264 ( 
.A1(n_252),
.A2(n_196),
.B(n_201),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_SL g305 ( 
.A(n_264),
.B(n_273),
.C(n_238),
.Y(n_305)
);

AOI21xp5_ASAP7_75t_L g273 ( 
.A1(n_237),
.A2(n_196),
.B(n_183),
.Y(n_273)
);

BUFx6f_ASAP7_75t_L g274 ( 
.A(n_231),
.Y(n_274)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_274),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_242),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_275),
.B(n_279),
.Y(n_298)
);

AOI22xp33_ASAP7_75t_L g277 ( 
.A1(n_226),
.A2(n_214),
.B1(n_180),
.B2(n_210),
.Y(n_277)
);

AOI22xp33_ASAP7_75t_SL g300 ( 
.A1(n_277),
.A2(n_233),
.B1(n_244),
.B2(n_245),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_278),
.A2(n_227),
.B1(n_226),
.B2(n_247),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_225),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_230),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_281),
.B(n_241),
.Y(n_294)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_283),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_259),
.B(n_229),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_286),
.B(n_293),
.C(n_304),
.Y(n_311)
);

BUFx12_ASAP7_75t_L g287 ( 
.A(n_269),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_287),
.B(n_302),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_SL g288 ( 
.A(n_276),
.B(n_234),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_288),
.B(n_290),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_271),
.B(n_251),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_267),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_292),
.B(n_301),
.Y(n_310)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_294),
.Y(n_315)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_280),
.Y(n_296)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_296),
.Y(n_318)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_280),
.Y(n_297)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_297),
.Y(n_314)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_272),
.Y(n_299)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_299),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_SL g319 ( 
.A1(n_300),
.A2(n_253),
.B1(n_273),
.B2(n_264),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_275),
.B(n_229),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_265),
.B(n_203),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_272),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_303),
.A2(n_306),
.B1(n_254),
.B2(n_262),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_255),
.B(n_232),
.C(n_218),
.Y(n_304)
);

XNOR2x1_ASAP7_75t_L g328 ( 
.A(n_305),
.B(n_307),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_265),
.B(n_238),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_262),
.B(n_228),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_SL g313 ( 
.A(n_308),
.B(n_278),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_SL g344 ( 
.A1(n_312),
.A2(n_321),
.B1(n_323),
.B2(n_325),
.Y(n_344)
);

XNOR2xp5_ASAP7_75t_SL g337 ( 
.A(n_313),
.B(n_295),
.Y(n_337)
);

OA21x2_ASAP7_75t_SL g316 ( 
.A1(n_301),
.A2(n_271),
.B(n_282),
.Y(n_316)
);

NOR3xp33_ASAP7_75t_SL g333 ( 
.A(n_316),
.B(n_308),
.C(n_270),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_293),
.B(n_261),
.C(n_282),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_317),
.B(n_329),
.C(n_291),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_L g343 ( 
.A1(n_319),
.A2(n_322),
.B1(n_219),
.B2(n_303),
.Y(n_343)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_289),
.A2(n_257),
.B1(n_258),
.B2(n_270),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_SL g322 ( 
.A1(n_296),
.A2(n_258),
.B1(n_256),
.B2(n_266),
.Y(n_322)
);

AOI22xp5_ASAP7_75t_L g323 ( 
.A1(n_306),
.A2(n_297),
.B1(n_285),
.B2(n_257),
.Y(n_323)
);

XOR2xp5_ASAP7_75t_L g324 ( 
.A(n_304),
.B(n_261),
.Y(n_324)
);

XOR2xp5_ASAP7_75t_L g330 ( 
.A(n_324),
.B(n_327),
.Y(n_330)
);

AOI22xp5_ASAP7_75t_L g325 ( 
.A1(n_285),
.A2(n_257),
.B1(n_307),
.B2(n_292),
.Y(n_325)
);

XOR2xp5_ASAP7_75t_L g327 ( 
.A(n_286),
.B(n_261),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_291),
.B(n_266),
.C(n_268),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_L g354 ( 
.A(n_331),
.B(n_337),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_309),
.B(n_288),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_332),
.B(n_333),
.Y(n_352)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_320),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_334),
.B(n_335),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_310),
.B(n_298),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_326),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_336),
.B(n_338),
.Y(n_351)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_310),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_313),
.B(n_260),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_SL g349 ( 
.A(n_339),
.B(n_346),
.Y(n_349)
);

XNOR2x1_ASAP7_75t_L g340 ( 
.A(n_324),
.B(n_295),
.Y(n_340)
);

XOR2xp5_ASAP7_75t_L g359 ( 
.A(n_340),
.B(n_343),
.Y(n_359)
);

OAI21xp5_ASAP7_75t_L g341 ( 
.A1(n_319),
.A2(n_305),
.B(n_294),
.Y(n_341)
);

AND2x2_ASAP7_75t_L g347 ( 
.A(n_341),
.B(n_342),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_315),
.B(n_281),
.Y(n_342)
);

AOI21xp5_ASAP7_75t_L g345 ( 
.A1(n_323),
.A2(n_263),
.B(n_235),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_L g356 ( 
.A(n_345),
.B(n_327),
.Y(n_356)
);

OR2x2_ASAP7_75t_L g346 ( 
.A(n_318),
.B(n_222),
.Y(n_346)
);

AOI22xp5_ASAP7_75t_SL g348 ( 
.A1(n_344),
.A2(n_329),
.B1(n_322),
.B2(n_317),
.Y(n_348)
);

XNOR2xp5_ASAP7_75t_L g363 ( 
.A(n_348),
.B(n_355),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_SL g350 ( 
.A(n_331),
.B(n_311),
.Y(n_350)
);

AOI21xp5_ASAP7_75t_L g368 ( 
.A1(n_350),
.A2(n_356),
.B(n_343),
.Y(n_368)
);

XNOR2xp5_ASAP7_75t_L g355 ( 
.A(n_330),
.B(n_311),
.Y(n_355)
);

MAJIxp5_ASAP7_75t_L g357 ( 
.A(n_330),
.B(n_328),
.C(n_314),
.Y(n_357)
);

MAJIxp5_ASAP7_75t_L g360 ( 
.A(n_357),
.B(n_358),
.C(n_354),
.Y(n_360)
);

XNOR2xp5_ASAP7_75t_L g358 ( 
.A(n_340),
.B(n_328),
.Y(n_358)
);

XNOR2xp5_ASAP7_75t_L g374 ( 
.A(n_360),
.B(n_361),
.Y(n_374)
);

XOR2xp5_ASAP7_75t_L g361 ( 
.A(n_357),
.B(n_341),
.Y(n_361)
);

AOI22xp5_ASAP7_75t_L g362 ( 
.A1(n_347),
.A2(n_344),
.B1(n_338),
.B2(n_335),
.Y(n_362)
);

AND2x2_ASAP7_75t_L g375 ( 
.A(n_362),
.B(n_365),
.Y(n_375)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_348),
.B(n_359),
.C(n_347),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_364),
.B(n_366),
.Y(n_371)
);

AOI22xp5_ASAP7_75t_L g365 ( 
.A1(n_359),
.A2(n_314),
.B1(n_342),
.B2(n_333),
.Y(n_365)
);

AOI22xp5_ASAP7_75t_L g366 ( 
.A1(n_353),
.A2(n_326),
.B1(n_299),
.B2(n_279),
.Y(n_366)
);

OAI21xp5_ASAP7_75t_SL g367 ( 
.A1(n_352),
.A2(n_345),
.B(n_346),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_367),
.B(n_369),
.Y(n_372)
);

XOR2xp5_ASAP7_75t_L g373 ( 
.A(n_368),
.B(n_337),
.Y(n_373)
);

AOI22xp5_ASAP7_75t_L g369 ( 
.A1(n_349),
.A2(n_302),
.B1(n_312),
.B2(n_284),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_SL g370 ( 
.A(n_360),
.B(n_351),
.Y(n_370)
);

AOI21xp5_ASAP7_75t_L g381 ( 
.A1(n_370),
.A2(n_376),
.B(n_377),
.Y(n_381)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_373),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_SL g376 ( 
.A(n_363),
.B(n_274),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_L g377 ( 
.A(n_365),
.B(n_274),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_L g378 ( 
.A(n_362),
.B(n_321),
.Y(n_378)
);

OAI21xp5_ASAP7_75t_L g380 ( 
.A1(n_378),
.A2(n_364),
.B(n_283),
.Y(n_380)
);

XNOR2xp5_ASAP7_75t_SL g379 ( 
.A(n_375),
.B(n_361),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_L g386 ( 
.A(n_379),
.B(n_380),
.Y(n_386)
);

AOI22xp5_ASAP7_75t_L g382 ( 
.A1(n_372),
.A2(n_284),
.B1(n_363),
.B2(n_267),
.Y(n_382)
);

OAI22xp5_ASAP7_75t_L g385 ( 
.A1(n_382),
.A2(n_384),
.B1(n_378),
.B2(n_371),
.Y(n_385)
);

XOR2xp5_ASAP7_75t_L g384 ( 
.A(n_374),
.B(n_325),
.Y(n_384)
);

AOI322xp5_ASAP7_75t_L g388 ( 
.A1(n_385),
.A2(n_387),
.A3(n_287),
.B1(n_381),
.B2(n_218),
.C1(n_379),
.C2(n_219),
.Y(n_388)
);

AOI322xp5_ASAP7_75t_L g387 ( 
.A1(n_383),
.A2(n_375),
.A3(n_198),
.B1(n_287),
.B2(n_218),
.C1(n_222),
.C2(n_267),
.Y(n_387)
);

AOI21xp5_ASAP7_75t_L g390 ( 
.A1(n_388),
.A2(n_389),
.B(n_183),
.Y(n_390)
);

AOI31xp67_ASAP7_75t_SL g389 ( 
.A1(n_386),
.A2(n_287),
.A3(n_248),
.B(n_250),
.Y(n_389)
);

AOI21xp5_ASAP7_75t_L g391 ( 
.A1(n_390),
.A2(n_182),
.B(n_352),
.Y(n_391)
);

XNOR2xp5_ASAP7_75t_L g392 ( 
.A(n_391),
.B(n_182),
.Y(n_392)
);


endmodule