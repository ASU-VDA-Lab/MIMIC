module fake_netlist_5_2300_n_627 (n_16, n_0, n_12, n_9, n_25, n_18, n_22, n_1, n_8, n_10, n_24, n_21, n_4, n_11, n_17, n_19, n_7, n_15, n_26, n_20, n_5, n_14, n_2, n_23, n_13, n_3, n_6, n_627);

input n_16;
input n_0;
input n_12;
input n_9;
input n_25;
input n_18;
input n_22;
input n_1;
input n_8;
input n_10;
input n_24;
input n_21;
input n_4;
input n_11;
input n_17;
input n_19;
input n_7;
input n_15;
input n_26;
input n_20;
input n_5;
input n_14;
input n_2;
input n_23;
input n_13;
input n_3;
input n_6;

output n_627;

wire n_137;
wire n_294;
wire n_431;
wire n_318;
wire n_419;
wire n_380;
wire n_611;
wire n_444;
wire n_469;
wire n_615;
wire n_82;
wire n_194;
wire n_316;
wire n_389;
wire n_549;
wire n_418;
wire n_248;
wire n_124;
wire n_86;
wire n_136;
wire n_146;
wire n_315;
wire n_268;
wire n_523;
wire n_451;
wire n_532;
wire n_619;
wire n_408;
wire n_61;
wire n_376;
wire n_503;
wire n_127;
wire n_75;
wire n_235;
wire n_226;
wire n_605;
wire n_74;
wire n_515;
wire n_57;
wire n_353;
wire n_351;
wire n_367;
wire n_620;
wire n_452;
wire n_397;
wire n_493;
wire n_111;
wire n_525;
wire n_483;
wire n_544;
wire n_155;
wire n_552;
wire n_547;
wire n_43;
wire n_116;
wire n_467;
wire n_564;
wire n_423;
wire n_501;
wire n_46;
wire n_245;
wire n_284;
wire n_139;
wire n_38;
wire n_105;
wire n_280;
wire n_590;
wire n_378;
wire n_551;
wire n_581;
wire n_382;
wire n_554;
wire n_254;
wire n_33;
wire n_583;
wire n_302;
wire n_265;
wire n_526;
wire n_372;
wire n_443;
wire n_293;
wire n_244;
wire n_47;
wire n_173;
wire n_198;
wire n_447;
wire n_247;
wire n_368;
wire n_314;
wire n_433;
wire n_604;
wire n_321;
wire n_292;
wire n_625;
wire n_621;
wire n_100;
wire n_455;
wire n_417;
wire n_612;
wire n_212;
wire n_385;
wire n_498;
wire n_516;
wire n_507;
wire n_119;
wire n_497;
wire n_606;
wire n_559;
wire n_275;
wire n_252;
wire n_624;
wire n_295;
wire n_133;
wire n_330;
wire n_508;
wire n_506;
wire n_610;
wire n_509;
wire n_568;
wire n_39;
wire n_147;
wire n_373;
wire n_67;
wire n_307;
wire n_439;
wire n_87;
wire n_150;
wire n_530;
wire n_556;
wire n_106;
wire n_209;
wire n_259;
wire n_448;
wire n_375;
wire n_301;
wire n_576;
wire n_68;
wire n_93;
wire n_186;
wire n_537;
wire n_134;
wire n_191;
wire n_587;
wire n_51;
wire n_63;
wire n_492;
wire n_563;
wire n_171;
wire n_153;
wire n_524;
wire n_399;
wire n_341;
wire n_204;
wire n_394;
wire n_250;
wire n_579;
wire n_548;
wire n_543;
wire n_260;
wire n_298;
wire n_320;
wire n_518;
wire n_505;
wire n_286;
wire n_122;
wire n_282;
wire n_331;
wire n_406;
wire n_519;
wire n_470;
wire n_325;
wire n_449;
wire n_132;
wire n_90;
wire n_546;
wire n_101;
wire n_281;
wire n_240;
wire n_381;
wire n_189;
wire n_220;
wire n_291;
wire n_231;
wire n_257;
wire n_390;
wire n_31;
wire n_456;
wire n_371;
wire n_481;
wire n_535;
wire n_152;
wire n_540;
wire n_317;
wire n_618;
wire n_323;
wire n_569;
wire n_195;
wire n_42;
wire n_356;
wire n_227;
wire n_592;
wire n_45;
wire n_271;
wire n_94;
wire n_335;
wire n_123;
wire n_370;
wire n_167;
wire n_234;
wire n_343;
wire n_379;
wire n_428;
wire n_308;
wire n_267;
wire n_514;
wire n_457;
wire n_570;
wire n_297;
wire n_156;
wire n_603;
wire n_225;
wire n_377;
wire n_484;
wire n_219;
wire n_442;
wire n_157;
wire n_131;
wire n_192;
wire n_600;
wire n_223;
wire n_392;
wire n_158;
wire n_138;
wire n_264;
wire n_109;
wire n_472;
wire n_454;
wire n_387;
wire n_374;
wire n_163;
wire n_276;
wire n_339;
wire n_95;
wire n_185;
wire n_183;
wire n_243;
wire n_398;
wire n_396;
wire n_347;
wire n_169;
wire n_59;
wire n_522;
wire n_550;
wire n_255;
wire n_215;
wire n_350;
wire n_196;
wire n_459;
wire n_211;
wire n_218;
wire n_400;
wire n_181;
wire n_436;
wire n_290;
wire n_580;
wire n_221;
wire n_178;
wire n_622;
wire n_386;
wire n_578;
wire n_287;
wire n_344;
wire n_555;
wire n_473;
wire n_422;
wire n_475;
wire n_72;
wire n_104;
wire n_41;
wire n_415;
wire n_56;
wire n_141;
wire n_485;
wire n_496;
wire n_355;
wire n_486;
wire n_336;
wire n_584;
wire n_591;
wire n_145;
wire n_48;
wire n_521;
wire n_614;
wire n_50;
wire n_337;
wire n_430;
wire n_313;
wire n_88;
wire n_479;
wire n_528;
wire n_510;
wire n_216;
wire n_168;
wire n_395;
wire n_164;
wire n_432;
wire n_553;
wire n_311;
wire n_208;
wire n_142;
wire n_214;
wire n_328;
wire n_140;
wire n_299;
wire n_303;
wire n_369;
wire n_296;
wire n_613;
wire n_241;
wire n_357;
wire n_598;
wire n_608;
wire n_184;
wire n_446;
wire n_445;
wire n_65;
wire n_78;
wire n_144;
wire n_114;
wire n_96;
wire n_165;
wire n_468;
wire n_499;
wire n_213;
wire n_129;
wire n_342;
wire n_482;
wire n_517;
wire n_98;
wire n_588;
wire n_361;
wire n_464;
wire n_363;
wire n_402;
wire n_413;
wire n_197;
wire n_107;
wire n_573;
wire n_69;
wire n_236;
wire n_388;
wire n_249;
wire n_304;
wire n_329;
wire n_203;
wire n_274;
wire n_577;
wire n_384;
wire n_582;
wire n_460;
wire n_80;
wire n_35;
wire n_73;
wire n_277;
wire n_92;
wire n_338;
wire n_149;
wire n_477;
wire n_461;
wire n_571;
wire n_333;
wire n_309;
wire n_30;
wire n_512;
wire n_84;
wire n_462;
wire n_130;
wire n_322;
wire n_567;
wire n_258;
wire n_29;
wire n_79;
wire n_151;
wire n_306;
wire n_458;
wire n_288;
wire n_188;
wire n_190;
wire n_201;
wire n_263;
wire n_471;
wire n_609;
wire n_44;
wire n_224;
wire n_40;
wire n_34;
wire n_228;
wire n_283;
wire n_383;
wire n_474;
wire n_112;
wire n_542;
wire n_85;
wire n_463;
wire n_488;
wire n_595;
wire n_502;
wire n_239;
wire n_466;
wire n_420;
wire n_489;
wire n_55;
wire n_617;
wire n_49;
wire n_310;
wire n_54;
wire n_593;
wire n_504;
wire n_511;
wire n_586;
wire n_465;
wire n_76;
wire n_358;
wire n_362;
wire n_170;
wire n_332;
wire n_27;
wire n_77;
wire n_102;
wire n_161;
wire n_273;
wire n_349;
wire n_585;
wire n_270;
wire n_616;
wire n_230;
wire n_81;
wire n_118;
wire n_601;
wire n_279;
wire n_70;
wire n_253;
wire n_261;
wire n_174;
wire n_289;
wire n_206;
wire n_172;
wire n_217;
wire n_440;
wire n_478;
wire n_545;
wire n_441;
wire n_450;
wire n_312;
wire n_476;
wire n_429;
wire n_534;
wire n_345;
wire n_210;
wire n_494;
wire n_365;
wire n_91;
wire n_176;
wire n_557;
wire n_182;
wire n_143;
wire n_83;
wire n_354;
wire n_575;
wire n_607;
wire n_480;
wire n_237;
wire n_425;
wire n_513;
wire n_407;
wire n_527;
wire n_180;
wire n_560;
wire n_340;
wire n_207;
wire n_561;
wire n_37;
wire n_346;
wire n_393;
wire n_229;
wire n_108;
wire n_495;
wire n_487;
wire n_602;
wire n_574;
wire n_437;
wire n_66;
wire n_177;
wire n_60;
wire n_403;
wire n_453;
wire n_421;
wire n_58;
wire n_623;
wire n_405;
wire n_359;
wire n_490;
wire n_117;
wire n_326;
wire n_233;
wire n_404;
wire n_205;
wire n_366;
wire n_572;
wire n_113;
wire n_246;
wire n_596;
wire n_179;
wire n_125;
wire n_410;
wire n_558;
wire n_269;
wire n_529;
wire n_128;
wire n_285;
wire n_412;
wire n_120;
wire n_232;
wire n_327;
wire n_135;
wire n_126;
wire n_202;
wire n_266;
wire n_272;
wire n_491;
wire n_427;
wire n_193;
wire n_251;
wire n_352;
wire n_53;
wire n_160;
wire n_566;
wire n_426;
wire n_520;
wire n_565;
wire n_409;
wire n_589;
wire n_597;
wire n_500;
wire n_562;
wire n_154;
wire n_62;
wire n_148;
wire n_71;
wire n_300;
wire n_435;
wire n_159;
wire n_334;
wire n_599;
wire n_541;
wire n_391;
wire n_434;
wire n_539;
wire n_175;
wire n_538;
wire n_262;
wire n_238;
wire n_99;
wire n_411;
wire n_414;
wire n_319;
wire n_364;
wire n_536;
wire n_531;
wire n_121;
wire n_242;
wire n_360;
wire n_36;
wire n_594;
wire n_200;
wire n_162;
wire n_64;
wire n_222;
wire n_28;
wire n_89;
wire n_438;
wire n_115;
wire n_324;
wire n_416;
wire n_199;
wire n_187;
wire n_32;
wire n_401;
wire n_103;
wire n_348;
wire n_97;
wire n_166;
wire n_626;
wire n_424;
wire n_256;
wire n_305;
wire n_533;
wire n_52;
wire n_278;
wire n_110;

INVx1_ASAP7_75t_L g27 ( 
.A(n_23),
.Y(n_27)
);

INVxp67_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_26),
.B(n_2),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_20),
.Y(n_32)
);

BUFx10_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

INVx2_ASAP7_75t_SL g34 ( 
.A(n_3),
.Y(n_34)
);

XOR2xp5_ASAP7_75t_L g35 ( 
.A(n_22),
.B(n_6),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_5),
.Y(n_36)
);

NOR2xp67_ASAP7_75t_L g37 ( 
.A(n_14),
.B(n_0),
.Y(n_37)
);

CKINVDCx5p33_ASAP7_75t_R g38 ( 
.A(n_13),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_2),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_24),
.Y(n_40)
);

BUFx2_ASAP7_75t_L g41 ( 
.A(n_16),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_7),
.Y(n_42)
);

BUFx10_ASAP7_75t_L g43 ( 
.A(n_18),
.Y(n_43)
);

INVx1_ASAP7_75t_SL g44 ( 
.A(n_7),
.Y(n_44)
);

OR2x2_ASAP7_75t_L g45 ( 
.A(n_16),
.B(n_8),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_0),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_25),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_19),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_9),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_4),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_14),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_10),
.Y(n_52)
);

INVx1_ASAP7_75t_SL g53 ( 
.A(n_11),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

OA21x2_ASAP7_75t_L g56 ( 
.A1(n_42),
.A2(n_1),
.B(n_3),
.Y(n_56)
);

OA21x2_ASAP7_75t_L g57 ( 
.A1(n_42),
.A2(n_1),
.B(n_5),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_36),
.Y(n_59)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_27),
.Y(n_60)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_27),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_48),
.Y(n_62)
);

AND2x4_ASAP7_75t_L g63 ( 
.A(n_48),
.B(n_32),
.Y(n_63)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_36),
.Y(n_64)
);

BUFx8_ASAP7_75t_L g65 ( 
.A(n_41),
.Y(n_65)
);

AND2x4_ASAP7_75t_L g66 ( 
.A(n_48),
.B(n_21),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_63),
.B(n_36),
.Y(n_67)
);

NAND2xp33_ASAP7_75t_L g68 ( 
.A(n_62),
.B(n_36),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_60),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_63),
.B(n_36),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_60),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_60),
.Y(n_72)
);

BUFx2_ASAP7_75t_L g73 ( 
.A(n_65),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_60),
.Y(n_74)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_64),
.Y(n_75)
);

AND2x4_ASAP7_75t_L g76 ( 
.A(n_66),
.B(n_32),
.Y(n_76)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_64),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_65),
.B(n_43),
.Y(n_78)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_59),
.Y(n_79)
);

INVx8_ASAP7_75t_L g80 ( 
.A(n_66),
.Y(n_80)
);

CKINVDCx5p33_ASAP7_75t_R g81 ( 
.A(n_65),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_63),
.B(n_36),
.Y(n_82)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_64),
.Y(n_83)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_64),
.Y(n_84)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_64),
.Y(n_85)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_59),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_78),
.A2(n_35),
.B1(n_41),
.B2(n_53),
.Y(n_87)
);

INVx2_ASAP7_75t_SL g88 ( 
.A(n_67),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_75),
.B(n_65),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_75),
.B(n_77),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_81),
.A2(n_35),
.B1(n_44),
.B2(n_38),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_75),
.B(n_66),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_L g93 ( 
.A1(n_78),
.A2(n_65),
.B1(n_63),
.B2(n_56),
.Y(n_93)
);

BUFx6f_ASAP7_75t_SL g94 ( 
.A(n_76),
.Y(n_94)
);

INVx1_ASAP7_75t_SL g95 ( 
.A(n_76),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_75),
.B(n_66),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_75),
.B(n_66),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_83),
.Y(n_98)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_83),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_73),
.B(n_65),
.Y(n_100)
);

OR2x6_ASAP7_75t_L g101 ( 
.A(n_76),
.B(n_66),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_77),
.B(n_66),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_77),
.B(n_66),
.Y(n_103)
);

OR2x6_ASAP7_75t_L g104 ( 
.A(n_76),
.B(n_45),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_77),
.B(n_63),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_77),
.B(n_63),
.Y(n_106)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_69),
.Y(n_107)
);

BUFx3_ASAP7_75t_L g108 ( 
.A(n_67),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_83),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_84),
.B(n_65),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_73),
.A2(n_45),
.B1(n_28),
.B2(n_31),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_84),
.B(n_63),
.Y(n_112)
);

BUFx3_ASAP7_75t_L g113 ( 
.A(n_67),
.Y(n_113)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_84),
.Y(n_114)
);

OAI221xp5_ASAP7_75t_L g115 ( 
.A1(n_70),
.A2(n_42),
.B1(n_34),
.B2(n_46),
.C(n_39),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_73),
.B(n_43),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_85),
.B(n_63),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_85),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_85),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_82),
.B(n_62),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_76),
.B(n_34),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_82),
.B(n_62),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_82),
.B(n_43),
.Y(n_123)
);

NAND2xp33_ASAP7_75t_L g124 ( 
.A(n_80),
.B(n_62),
.Y(n_124)
);

INVx2_ASAP7_75t_SL g125 ( 
.A(n_123),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_L g126 ( 
.A1(n_93),
.A2(n_56),
.B1(n_57),
.B2(n_61),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_88),
.B(n_70),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_88),
.B(n_80),
.Y(n_128)
);

NAND2x1_ASAP7_75t_L g129 ( 
.A(n_101),
.B(n_64),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_108),
.B(n_80),
.Y(n_130)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_108),
.Y(n_131)
);

AOI21xp5_ASAP7_75t_L g132 ( 
.A1(n_124),
.A2(n_80),
.B(n_68),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_113),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_95),
.B(n_80),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_113),
.Y(n_135)
);

OR2x2_ASAP7_75t_L g136 ( 
.A(n_87),
.B(n_44),
.Y(n_136)
);

AOI21xp5_ASAP7_75t_L g137 ( 
.A1(n_124),
.A2(n_80),
.B(n_68),
.Y(n_137)
);

A2O1A1Ixp33_ASAP7_75t_L g138 ( 
.A1(n_121),
.A2(n_80),
.B(n_47),
.C(n_37),
.Y(n_138)
);

A2O1A1Ixp33_ASAP7_75t_L g139 ( 
.A1(n_87),
.A2(n_47),
.B(n_37),
.C(n_60),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_104),
.A2(n_62),
.B1(n_57),
.B2(n_56),
.Y(n_140)
);

AOI21xp5_ASAP7_75t_L g141 ( 
.A1(n_105),
.A2(n_86),
.B(n_79),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_98),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_104),
.A2(n_62),
.B1(n_57),
.B2(n_56),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_120),
.B(n_62),
.Y(n_144)
);

AND2x2_ASAP7_75t_L g145 ( 
.A(n_104),
.B(n_33),
.Y(n_145)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_107),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_98),
.B(n_62),
.Y(n_147)
);

O2A1O1Ixp5_ASAP7_75t_L g148 ( 
.A1(n_90),
.A2(n_61),
.B(n_64),
.C(n_58),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_104),
.A2(n_62),
.B1(n_56),
.B2(n_57),
.Y(n_149)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_107),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_111),
.A2(n_62),
.B1(n_56),
.B2(n_57),
.Y(n_151)
);

AOI21xp5_ASAP7_75t_L g152 ( 
.A1(n_106),
.A2(n_86),
.B(n_79),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_L g153 ( 
.A1(n_92),
.A2(n_102),
.B(n_103),
.Y(n_153)
);

CKINVDCx10_ASAP7_75t_R g154 ( 
.A(n_91),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_L g155 ( 
.A1(n_112),
.A2(n_86),
.B(n_79),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_116),
.B(n_33),
.Y(n_156)
);

NOR2x1p5_ASAP7_75t_SL g157 ( 
.A(n_99),
.B(n_86),
.Y(n_157)
);

AOI21xp5_ASAP7_75t_L g158 ( 
.A1(n_117),
.A2(n_79),
.B(n_74),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_101),
.A2(n_57),
.B1(n_56),
.B2(n_61),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_122),
.B(n_62),
.Y(n_160)
);

AOI21x1_ASAP7_75t_L g161 ( 
.A1(n_99),
.A2(n_74),
.B(n_72),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_101),
.A2(n_57),
.B1(n_56),
.B2(n_61),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_101),
.A2(n_57),
.B1(n_43),
.B2(n_61),
.Y(n_163)
);

AOI21xp5_ASAP7_75t_L g164 ( 
.A1(n_96),
.A2(n_72),
.B(n_71),
.Y(n_164)
);

BUFx12f_ASAP7_75t_L g165 ( 
.A(n_115),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_109),
.Y(n_166)
);

BUFx12f_ASAP7_75t_L g167 ( 
.A(n_94),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_109),
.B(n_71),
.Y(n_168)
);

OR2x2_ASAP7_75t_L g169 ( 
.A(n_114),
.B(n_39),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_114),
.B(n_69),
.Y(n_170)
);

NAND2x1p5_ASAP7_75t_L g171 ( 
.A(n_118),
.B(n_55),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_119),
.B(n_33),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_118),
.B(n_55),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_119),
.Y(n_174)
);

OAI21x1_ASAP7_75t_L g175 ( 
.A1(n_97),
.A2(n_58),
.B(n_54),
.Y(n_175)
);

AOI21xp5_ASAP7_75t_L g176 ( 
.A1(n_110),
.A2(n_58),
.B(n_59),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_89),
.B(n_55),
.Y(n_177)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_94),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_100),
.B(n_33),
.Y(n_179)
);

O2A1O1Ixp33_ASAP7_75t_SL g180 ( 
.A1(n_94),
.A2(n_30),
.B(n_46),
.C(n_29),
.Y(n_180)
);

OR2x2_ASAP7_75t_L g181 ( 
.A(n_136),
.B(n_30),
.Y(n_181)
);

BUFx10_ASAP7_75t_L g182 ( 
.A(n_179),
.Y(n_182)
);

OAI21x1_ASAP7_75t_L g183 ( 
.A1(n_161),
.A2(n_175),
.B(n_148),
.Y(n_183)
);

CKINVDCx8_ASAP7_75t_R g184 ( 
.A(n_154),
.Y(n_184)
);

A2O1A1Ixp33_ASAP7_75t_L g185 ( 
.A1(n_179),
.A2(n_156),
.B(n_172),
.C(n_153),
.Y(n_185)
);

AO21x2_ASAP7_75t_L g186 ( 
.A1(n_177),
.A2(n_54),
.B(n_58),
.Y(n_186)
);

INVxp67_ASAP7_75t_SL g187 ( 
.A(n_131),
.Y(n_187)
);

CKINVDCx11_ASAP7_75t_R g188 ( 
.A(n_167),
.Y(n_188)
);

AOI21xp5_ASAP7_75t_L g189 ( 
.A1(n_132),
.A2(n_137),
.B(n_130),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_131),
.B(n_54),
.Y(n_190)
);

OAI21x1_ASAP7_75t_L g191 ( 
.A1(n_148),
.A2(n_58),
.B(n_29),
.Y(n_191)
);

AO31x2_ASAP7_75t_L g192 ( 
.A1(n_159),
.A2(n_52),
.A3(n_51),
.B(n_50),
.Y(n_192)
);

OAI21x1_ASAP7_75t_L g193 ( 
.A1(n_162),
.A2(n_52),
.B(n_51),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_133),
.Y(n_194)
);

OAI21x1_ASAP7_75t_SL g195 ( 
.A1(n_126),
.A2(n_50),
.B(n_49),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_135),
.Y(n_196)
);

BUFx12f_ASAP7_75t_L g197 ( 
.A(n_165),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_145),
.Y(n_198)
);

INVx2_ASAP7_75t_SL g199 ( 
.A(n_166),
.Y(n_199)
);

NAND2xp33_ASAP7_75t_R g200 ( 
.A(n_156),
.B(n_6),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_127),
.B(n_49),
.Y(n_201)
);

OA21x2_ASAP7_75t_L g202 ( 
.A1(n_126),
.A2(n_59),
.B(n_9),
.Y(n_202)
);

NAND2xp33_ASAP7_75t_L g203 ( 
.A(n_166),
.B(n_59),
.Y(n_203)
);

AOI21xp5_ASAP7_75t_L g204 ( 
.A1(n_128),
.A2(n_134),
.B(n_129),
.Y(n_204)
);

AOI21xp5_ASAP7_75t_L g205 ( 
.A1(n_134),
.A2(n_59),
.B(n_10),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_142),
.Y(n_206)
);

BUFx6f_ASAP7_75t_L g207 ( 
.A(n_166),
.Y(n_207)
);

INVx3_ASAP7_75t_L g208 ( 
.A(n_166),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_172),
.B(n_59),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_125),
.A2(n_59),
.B1(n_12),
.B2(n_15),
.Y(n_210)
);

HB1xp67_ASAP7_75t_L g211 ( 
.A(n_169),
.Y(n_211)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_174),
.Y(n_212)
);

AOI21xp5_ASAP7_75t_L g213 ( 
.A1(n_144),
.A2(n_160),
.B(n_152),
.Y(n_213)
);

AOI221x1_ASAP7_75t_L g214 ( 
.A1(n_138),
.A2(n_8),
.B1(n_15),
.B2(n_17),
.C(n_59),
.Y(n_214)
);

BUFx2_ASAP7_75t_L g215 ( 
.A(n_178),
.Y(n_215)
);

OAI21x1_ASAP7_75t_L g216 ( 
.A1(n_164),
.A2(n_59),
.B(n_17),
.Y(n_216)
);

HB1xp67_ASAP7_75t_L g217 ( 
.A(n_139),
.Y(n_217)
);

OAI21x1_ASAP7_75t_L g218 ( 
.A1(n_147),
.A2(n_59),
.B(n_140),
.Y(n_218)
);

INVx1_ASAP7_75t_SL g219 ( 
.A(n_146),
.Y(n_219)
);

HB1xp67_ASAP7_75t_L g220 ( 
.A(n_150),
.Y(n_220)
);

AOI21xp5_ASAP7_75t_SL g221 ( 
.A1(n_143),
.A2(n_59),
.B(n_149),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_L g222 ( 
.A1(n_141),
.A2(n_151),
.B(n_155),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_L g223 ( 
.A1(n_163),
.A2(n_158),
.B(n_144),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_168),
.B(n_170),
.Y(n_224)
);

NOR2xp67_ASAP7_75t_L g225 ( 
.A(n_173),
.B(n_160),
.Y(n_225)
);

A2O1A1Ixp33_ASAP7_75t_L g226 ( 
.A1(n_157),
.A2(n_176),
.B(n_180),
.C(n_171),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_L g227 ( 
.A1(n_171),
.A2(n_153),
.B(n_148),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_180),
.Y(n_228)
);

OR2x2_ASAP7_75t_L g229 ( 
.A(n_211),
.B(n_181),
.Y(n_229)
);

INVx3_ASAP7_75t_L g230 ( 
.A(n_207),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_212),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_185),
.B(n_217),
.Y(n_232)
);

OAI21xp5_ASAP7_75t_L g233 ( 
.A1(n_227),
.A2(n_222),
.B(n_218),
.Y(n_233)
);

OAI21x1_ASAP7_75t_L g234 ( 
.A1(n_183),
.A2(n_189),
.B(n_218),
.Y(n_234)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_202),
.Y(n_235)
);

BUFx8_ASAP7_75t_L g236 ( 
.A(n_197),
.Y(n_236)
);

BUFx12f_ASAP7_75t_L g237 ( 
.A(n_188),
.Y(n_237)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_202),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_212),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_219),
.B(n_201),
.Y(n_240)
);

AO21x2_ASAP7_75t_L g241 ( 
.A1(n_193),
.A2(n_216),
.B(n_223),
.Y(n_241)
);

OAI21x1_ASAP7_75t_L g242 ( 
.A1(n_183),
.A2(n_204),
.B(n_191),
.Y(n_242)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_202),
.Y(n_243)
);

HB1xp67_ASAP7_75t_L g244 ( 
.A(n_215),
.Y(n_244)
);

AO21x2_ASAP7_75t_L g245 ( 
.A1(n_193),
.A2(n_216),
.B(n_195),
.Y(n_245)
);

INVx3_ASAP7_75t_L g246 ( 
.A(n_207),
.Y(n_246)
);

A2O1A1Ixp33_ASAP7_75t_L g247 ( 
.A1(n_206),
.A2(n_228),
.B(n_213),
.C(n_225),
.Y(n_247)
);

OAI21x1_ASAP7_75t_L g248 ( 
.A1(n_191),
.A2(n_195),
.B(n_221),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_207),
.Y(n_249)
);

OAI21x1_ASAP7_75t_L g250 ( 
.A1(n_221),
.A2(n_205),
.B(n_208),
.Y(n_250)
);

OR2x2_ASAP7_75t_L g251 ( 
.A(n_181),
.B(n_194),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_187),
.B(n_224),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_207),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_207),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_L g255 ( 
.A1(n_226),
.A2(n_209),
.B(n_214),
.Y(n_255)
);

AND2x2_ASAP7_75t_L g256 ( 
.A(n_182),
.B(n_192),
.Y(n_256)
);

BUFx3_ASAP7_75t_L g257 ( 
.A(n_208),
.Y(n_257)
);

OA21x2_ASAP7_75t_L g258 ( 
.A1(n_214),
.A2(n_190),
.B(n_196),
.Y(n_258)
);

BUFx2_ASAP7_75t_L g259 ( 
.A(n_208),
.Y(n_259)
);

INVx6_ASAP7_75t_L g260 ( 
.A(n_182),
.Y(n_260)
);

OAI21xp5_ASAP7_75t_L g261 ( 
.A1(n_199),
.A2(n_220),
.B(n_210),
.Y(n_261)
);

BUFx2_ASAP7_75t_R g262 ( 
.A(n_184),
.Y(n_262)
);

OAI21x1_ASAP7_75t_L g263 ( 
.A1(n_192),
.A2(n_186),
.B(n_199),
.Y(n_263)
);

OR2x6_ASAP7_75t_L g264 ( 
.A(n_215),
.B(n_197),
.Y(n_264)
);

AOI21xp5_ASAP7_75t_L g265 ( 
.A1(n_203),
.A2(n_186),
.B(n_198),
.Y(n_265)
);

OAI21x1_ASAP7_75t_L g266 ( 
.A1(n_192),
.A2(n_186),
.B(n_203),
.Y(n_266)
);

OAI21x1_ASAP7_75t_L g267 ( 
.A1(n_192),
.A2(n_182),
.B(n_200),
.Y(n_267)
);

OA21x2_ASAP7_75t_L g268 ( 
.A1(n_192),
.A2(n_198),
.B(n_188),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_184),
.B(n_185),
.Y(n_269)
);

OAI21x1_ASAP7_75t_L g270 ( 
.A1(n_183),
.A2(n_189),
.B(n_218),
.Y(n_270)
);

NOR2x1_ASAP7_75t_R g271 ( 
.A(n_188),
.B(n_167),
.Y(n_271)
);

NAND2x1p5_ASAP7_75t_L g272 ( 
.A(n_207),
.B(n_208),
.Y(n_272)
);

AND2x2_ASAP7_75t_L g273 ( 
.A(n_185),
.B(n_217),
.Y(n_273)
);

INVx2_ASAP7_75t_SL g274 ( 
.A(n_207),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_185),
.B(n_131),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_185),
.B(n_127),
.Y(n_276)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_202),
.Y(n_277)
);

OAI21x1_ASAP7_75t_L g278 ( 
.A1(n_183),
.A2(n_189),
.B(n_218),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_185),
.B(n_127),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_231),
.Y(n_280)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_235),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_231),
.Y(n_282)
);

BUFx6f_ASAP7_75t_L g283 ( 
.A(n_248),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_239),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_273),
.B(n_232),
.Y(n_285)
);

AO21x2_ASAP7_75t_L g286 ( 
.A1(n_255),
.A2(n_233),
.B(n_241),
.Y(n_286)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_235),
.Y(n_287)
);

AOI22xp33_ASAP7_75t_L g288 ( 
.A1(n_273),
.A2(n_269),
.B1(n_232),
.B2(n_276),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_239),
.Y(n_289)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_235),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_238),
.Y(n_291)
);

AND2x4_ASAP7_75t_L g292 ( 
.A(n_257),
.B(n_246),
.Y(n_292)
);

INVx2_ASAP7_75t_SL g293 ( 
.A(n_257),
.Y(n_293)
);

INVxp67_ASAP7_75t_L g294 ( 
.A(n_229),
.Y(n_294)
);

OA21x2_ASAP7_75t_L g295 ( 
.A1(n_255),
.A2(n_233),
.B(n_242),
.Y(n_295)
);

OR2x2_ASAP7_75t_L g296 ( 
.A(n_276),
.B(n_279),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_243),
.Y(n_297)
);

AND2x2_ASAP7_75t_L g298 ( 
.A(n_279),
.B(n_275),
.Y(n_298)
);

AO21x2_ASAP7_75t_L g299 ( 
.A1(n_241),
.A2(n_245),
.B(n_270),
.Y(n_299)
);

OR2x2_ASAP7_75t_L g300 ( 
.A(n_256),
.B(n_267),
.Y(n_300)
);

AND2x4_ASAP7_75t_L g301 ( 
.A(n_257),
.B(n_230),
.Y(n_301)
);

AO21x2_ASAP7_75t_L g302 ( 
.A1(n_241),
.A2(n_245),
.B(n_278),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_243),
.Y(n_303)
);

OR2x2_ASAP7_75t_L g304 ( 
.A(n_256),
.B(n_267),
.Y(n_304)
);

AND2x4_ASAP7_75t_L g305 ( 
.A(n_230),
.B(n_246),
.Y(n_305)
);

OR2x2_ASAP7_75t_L g306 ( 
.A(n_251),
.B(n_229),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_277),
.Y(n_307)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_242),
.Y(n_308)
);

HB1xp67_ASAP7_75t_L g309 ( 
.A(n_244),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_252),
.Y(n_310)
);

AND2x2_ASAP7_75t_L g311 ( 
.A(n_249),
.B(n_254),
.Y(n_311)
);

OAI21xp5_ASAP7_75t_L g312 ( 
.A1(n_247),
.A2(n_266),
.B(n_263),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_252),
.Y(n_313)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_248),
.Y(n_314)
);

AOI21x1_ASAP7_75t_L g315 ( 
.A1(n_234),
.A2(n_278),
.B(n_270),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_272),
.Y(n_316)
);

AND2x2_ASAP7_75t_L g317 ( 
.A(n_249),
.B(n_254),
.Y(n_317)
);

BUFx2_ASAP7_75t_L g318 ( 
.A(n_259),
.Y(n_318)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_263),
.Y(n_319)
);

CKINVDCx11_ASAP7_75t_R g320 ( 
.A(n_237),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_291),
.Y(n_321)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_281),
.Y(n_322)
);

AND2x2_ASAP7_75t_L g323 ( 
.A(n_288),
.B(n_268),
.Y(n_323)
);

NOR2xp67_ASAP7_75t_L g324 ( 
.A(n_310),
.B(n_240),
.Y(n_324)
);

AND2x2_ASAP7_75t_L g325 ( 
.A(n_288),
.B(n_268),
.Y(n_325)
);

AND2x4_ASAP7_75t_L g326 ( 
.A(n_292),
.B(n_230),
.Y(n_326)
);

HB1xp67_ASAP7_75t_L g327 ( 
.A(n_306),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_285),
.B(n_259),
.Y(n_328)
);

HB1xp67_ASAP7_75t_L g329 ( 
.A(n_306),
.Y(n_329)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_281),
.Y(n_330)
);

BUFx3_ASAP7_75t_L g331 ( 
.A(n_318),
.Y(n_331)
);

INVx2_ASAP7_75t_L g332 ( 
.A(n_281),
.Y(n_332)
);

INVx2_ASAP7_75t_L g333 ( 
.A(n_281),
.Y(n_333)
);

OAI22xp5_ASAP7_75t_L g334 ( 
.A1(n_285),
.A2(n_251),
.B1(n_265),
.B2(n_260),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_291),
.Y(n_335)
);

INVx2_ASAP7_75t_L g336 ( 
.A(n_287),
.Y(n_336)
);

BUFx5_ASAP7_75t_L g337 ( 
.A(n_298),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_297),
.Y(n_338)
);

INVx2_ASAP7_75t_L g339 ( 
.A(n_287),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_297),
.Y(n_340)
);

HB1xp67_ASAP7_75t_L g341 ( 
.A(n_306),
.Y(n_341)
);

INVxp67_ASAP7_75t_L g342 ( 
.A(n_309),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_303),
.Y(n_343)
);

HB1xp67_ASAP7_75t_L g344 ( 
.A(n_318),
.Y(n_344)
);

AND2x2_ASAP7_75t_L g345 ( 
.A(n_311),
.B(n_268),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_303),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_307),
.Y(n_347)
);

INVx2_ASAP7_75t_L g348 ( 
.A(n_287),
.Y(n_348)
);

AND2x2_ASAP7_75t_L g349 ( 
.A(n_311),
.B(n_268),
.Y(n_349)
);

NOR2x1_ASAP7_75t_SL g350 ( 
.A(n_310),
.B(n_245),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_307),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_287),
.Y(n_352)
);

AND2x2_ASAP7_75t_L g353 ( 
.A(n_311),
.B(n_258),
.Y(n_353)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_290),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_321),
.Y(n_355)
);

AND2x2_ASAP7_75t_L g356 ( 
.A(n_353),
.B(n_304),
.Y(n_356)
);

INVxp67_ASAP7_75t_L g357 ( 
.A(n_327),
.Y(n_357)
);

BUFx3_ASAP7_75t_L g358 ( 
.A(n_331),
.Y(n_358)
);

INVx2_ASAP7_75t_L g359 ( 
.A(n_337),
.Y(n_359)
);

INVxp67_ASAP7_75t_L g360 ( 
.A(n_329),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_321),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_335),
.Y(n_362)
);

OR2x2_ASAP7_75t_L g363 ( 
.A(n_341),
.B(n_300),
.Y(n_363)
);

INVxp67_ASAP7_75t_SL g364 ( 
.A(n_344),
.Y(n_364)
);

AND2x2_ASAP7_75t_L g365 ( 
.A(n_353),
.B(n_304),
.Y(n_365)
);

AND2x2_ASAP7_75t_L g366 ( 
.A(n_337),
.B(n_304),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_328),
.B(n_313),
.Y(n_367)
);

OR2x2_ASAP7_75t_L g368 ( 
.A(n_323),
.B(n_300),
.Y(n_368)
);

BUFx2_ASAP7_75t_L g369 ( 
.A(n_331),
.Y(n_369)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_337),
.Y(n_370)
);

INVx2_ASAP7_75t_SL g371 ( 
.A(n_331),
.Y(n_371)
);

INVx2_ASAP7_75t_L g372 ( 
.A(n_337),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_335),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_338),
.Y(n_374)
);

AND2x2_ASAP7_75t_L g375 ( 
.A(n_337),
.B(n_300),
.Y(n_375)
);

AND2x2_ASAP7_75t_L g376 ( 
.A(n_337),
.B(n_323),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_338),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_340),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_340),
.Y(n_379)
);

INVx5_ASAP7_75t_SL g380 ( 
.A(n_326),
.Y(n_380)
);

BUFx2_ASAP7_75t_L g381 ( 
.A(n_344),
.Y(n_381)
);

HB1xp67_ASAP7_75t_L g382 ( 
.A(n_337),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_343),
.Y(n_383)
);

NOR2x1_ASAP7_75t_L g384 ( 
.A(n_324),
.B(n_313),
.Y(n_384)
);

HB1xp67_ASAP7_75t_L g385 ( 
.A(n_342),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_343),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_346),
.Y(n_387)
);

HB1xp67_ASAP7_75t_L g388 ( 
.A(n_342),
.Y(n_388)
);

AND2x2_ASAP7_75t_L g389 ( 
.A(n_337),
.B(n_286),
.Y(n_389)
);

INVxp67_ASAP7_75t_L g390 ( 
.A(n_385),
.Y(n_390)
);

OR2x2_ASAP7_75t_L g391 ( 
.A(n_368),
.B(n_286),
.Y(n_391)
);

NOR4xp25_ASAP7_75t_L g392 ( 
.A(n_357),
.B(n_334),
.C(n_294),
.D(n_325),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_355),
.Y(n_393)
);

AND2x2_ASAP7_75t_L g394 ( 
.A(n_356),
.B(n_325),
.Y(n_394)
);

INVxp33_ASAP7_75t_L g395 ( 
.A(n_388),
.Y(n_395)
);

NOR2xp67_ASAP7_75t_L g396 ( 
.A(n_357),
.B(n_294),
.Y(n_396)
);

AND2x2_ASAP7_75t_L g397 ( 
.A(n_356),
.B(n_345),
.Y(n_397)
);

AND2x4_ASAP7_75t_L g398 ( 
.A(n_358),
.B(n_345),
.Y(n_398)
);

AND2x2_ASAP7_75t_L g399 ( 
.A(n_356),
.B(n_349),
.Y(n_399)
);

OR2x2_ASAP7_75t_L g400 ( 
.A(n_368),
.B(n_337),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_355),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_361),
.Y(n_402)
);

INVx2_ASAP7_75t_L g403 ( 
.A(n_361),
.Y(n_403)
);

OR2x2_ASAP7_75t_L g404 ( 
.A(n_376),
.B(n_286),
.Y(n_404)
);

AND2x2_ASAP7_75t_L g405 ( 
.A(n_365),
.B(n_349),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_360),
.B(n_328),
.Y(n_406)
);

AOI22xp5_ASAP7_75t_L g407 ( 
.A1(n_384),
.A2(n_334),
.B1(n_324),
.B2(n_264),
.Y(n_407)
);

OR2x2_ASAP7_75t_L g408 ( 
.A(n_365),
.B(n_337),
.Y(n_408)
);

AND2x4_ASAP7_75t_L g409 ( 
.A(n_358),
.B(n_350),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_362),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_362),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_373),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_373),
.Y(n_413)
);

OR2x2_ASAP7_75t_L g414 ( 
.A(n_376),
.B(n_286),
.Y(n_414)
);

OR2x2_ASAP7_75t_L g415 ( 
.A(n_376),
.B(n_286),
.Y(n_415)
);

OR2x2_ASAP7_75t_L g416 ( 
.A(n_365),
.B(n_295),
.Y(n_416)
);

AND2x2_ASAP7_75t_L g417 ( 
.A(n_366),
.B(n_350),
.Y(n_417)
);

AND2x2_ASAP7_75t_L g418 ( 
.A(n_366),
.B(n_295),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_360),
.B(n_298),
.Y(n_419)
);

AND2x4_ASAP7_75t_L g420 ( 
.A(n_358),
.B(n_314),
.Y(n_420)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_374),
.Y(n_421)
);

AND2x4_ASAP7_75t_L g422 ( 
.A(n_371),
.B(n_314),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_367),
.B(n_298),
.Y(n_423)
);

AND2x2_ASAP7_75t_L g424 ( 
.A(n_394),
.B(n_389),
.Y(n_424)
);

OR2x2_ASAP7_75t_L g425 ( 
.A(n_404),
.B(n_389),
.Y(n_425)
);

OR2x2_ASAP7_75t_L g426 ( 
.A(n_404),
.B(n_389),
.Y(n_426)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_403),
.Y(n_427)
);

AND2x4_ASAP7_75t_L g428 ( 
.A(n_409),
.B(n_371),
.Y(n_428)
);

AND2x2_ASAP7_75t_L g429 ( 
.A(n_394),
.B(n_366),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_403),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_421),
.Y(n_431)
);

INVx2_ASAP7_75t_SL g432 ( 
.A(n_421),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_393),
.Y(n_433)
);

NAND2x1p5_ASAP7_75t_L g434 ( 
.A(n_407),
.B(n_384),
.Y(n_434)
);

OR2x2_ASAP7_75t_L g435 ( 
.A(n_414),
.B(n_415),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_390),
.B(n_381),
.Y(n_436)
);

INVx2_ASAP7_75t_L g437 ( 
.A(n_401),
.Y(n_437)
);

NAND2x1_ASAP7_75t_L g438 ( 
.A(n_409),
.B(n_420),
.Y(n_438)
);

INVxp67_ASAP7_75t_L g439 ( 
.A(n_396),
.Y(n_439)
);

INVx3_ASAP7_75t_L g440 ( 
.A(n_409),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_402),
.Y(n_441)
);

AND2x2_ASAP7_75t_L g442 ( 
.A(n_417),
.B(n_375),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_406),
.B(n_381),
.Y(n_443)
);

INVx2_ASAP7_75t_L g444 ( 
.A(n_410),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_411),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_412),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_413),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_395),
.Y(n_448)
);

NOR2x1_ASAP7_75t_L g449 ( 
.A(n_419),
.B(n_369),
.Y(n_449)
);

NAND3xp33_ASAP7_75t_L g450 ( 
.A(n_392),
.B(n_367),
.C(n_309),
.Y(n_450)
);

NOR2xp33_ASAP7_75t_L g451 ( 
.A(n_395),
.B(n_320),
.Y(n_451)
);

AND2x2_ASAP7_75t_L g452 ( 
.A(n_417),
.B(n_375),
.Y(n_452)
);

OR2x2_ASAP7_75t_L g453 ( 
.A(n_414),
.B(n_363),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_391),
.Y(n_454)
);

AND2x2_ASAP7_75t_L g455 ( 
.A(n_418),
.B(n_375),
.Y(n_455)
);

AND2x2_ASAP7_75t_L g456 ( 
.A(n_418),
.B(n_397),
.Y(n_456)
);

OR2x2_ASAP7_75t_L g457 ( 
.A(n_415),
.B(n_363),
.Y(n_457)
);

INVxp67_ASAP7_75t_SL g458 ( 
.A(n_400),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_423),
.B(n_364),
.Y(n_459)
);

INVx2_ASAP7_75t_SL g460 ( 
.A(n_448),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_433),
.Y(n_461)
);

AND2x4_ASAP7_75t_L g462 ( 
.A(n_440),
.B(n_398),
.Y(n_462)
);

AND2x2_ASAP7_75t_L g463 ( 
.A(n_429),
.B(n_397),
.Y(n_463)
);

OAI221xp5_ASAP7_75t_L g464 ( 
.A1(n_434),
.A2(n_264),
.B1(n_391),
.B2(n_408),
.C(n_371),
.Y(n_464)
);

AND2x2_ASAP7_75t_L g465 ( 
.A(n_429),
.B(n_399),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_433),
.Y(n_466)
);

OAI221xp5_ASAP7_75t_L g467 ( 
.A1(n_434),
.A2(n_264),
.B1(n_416),
.B2(n_370),
.C(n_372),
.Y(n_467)
);

OAI22xp33_ASAP7_75t_L g468 ( 
.A1(n_450),
.A2(n_382),
.B1(n_359),
.B2(n_372),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_437),
.Y(n_469)
);

AO21x2_ASAP7_75t_L g470 ( 
.A1(n_454),
.A2(n_312),
.B(n_315),
.Y(n_470)
);

AOI22xp33_ASAP7_75t_L g471 ( 
.A1(n_451),
.A2(n_434),
.B1(n_436),
.B2(n_439),
.Y(n_471)
);

NAND2x1p5_ASAP7_75t_L g472 ( 
.A(n_449),
.B(n_369),
.Y(n_472)
);

NOR2xp33_ASAP7_75t_L g473 ( 
.A(n_443),
.B(n_399),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_437),
.Y(n_474)
);

OA21x2_ASAP7_75t_L g475 ( 
.A1(n_454),
.A2(n_379),
.B(n_387),
.Y(n_475)
);

OA21x2_ASAP7_75t_L g476 ( 
.A1(n_427),
.A2(n_379),
.B(n_387),
.Y(n_476)
);

OAI21xp5_ASAP7_75t_SL g477 ( 
.A1(n_440),
.A2(n_320),
.B(n_398),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_SL g478 ( 
.A(n_459),
.B(n_398),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_444),
.Y(n_479)
);

AOI21xp33_ASAP7_75t_SL g480 ( 
.A1(n_435),
.A2(n_264),
.B(n_262),
.Y(n_480)
);

INVx2_ASAP7_75t_L g481 ( 
.A(n_427),
.Y(n_481)
);

OAI22xp33_ASAP7_75t_L g482 ( 
.A1(n_458),
.A2(n_382),
.B1(n_359),
.B2(n_370),
.Y(n_482)
);

AOI22xp5_ASAP7_75t_L g483 ( 
.A1(n_428),
.A2(n_260),
.B1(n_380),
.B2(n_326),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_444),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_441),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g486 ( 
.A(n_424),
.B(n_405),
.Y(n_486)
);

AND2x4_ASAP7_75t_L g487 ( 
.A(n_440),
.B(n_420),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g488 ( 
.A(n_424),
.B(n_456),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_445),
.Y(n_489)
);

HB1xp67_ASAP7_75t_L g490 ( 
.A(n_432),
.Y(n_490)
);

AOI222xp33_ASAP7_75t_L g491 ( 
.A1(n_446),
.A2(n_271),
.B1(n_237),
.B2(n_236),
.C1(n_405),
.C2(n_364),
.Y(n_491)
);

NOR2xp33_ASAP7_75t_L g492 ( 
.A(n_435),
.B(n_260),
.Y(n_492)
);

NOR4xp25_ASAP7_75t_L g493 ( 
.A(n_447),
.B(n_377),
.C(n_386),
.D(n_383),
.Y(n_493)
);

NOR2xp33_ASAP7_75t_L g494 ( 
.A(n_480),
.B(n_237),
.Y(n_494)
);

OAI211xp5_ASAP7_75t_L g495 ( 
.A1(n_471),
.A2(n_438),
.B(n_426),
.C(n_425),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_461),
.Y(n_496)
);

O2A1O1Ixp33_ASAP7_75t_L g497 ( 
.A1(n_468),
.A2(n_264),
.B(n_438),
.C(n_430),
.Y(n_497)
);

AND2x2_ASAP7_75t_L g498 ( 
.A(n_462),
.B(n_442),
.Y(n_498)
);

NAND3xp33_ASAP7_75t_SL g499 ( 
.A(n_471),
.B(n_491),
.C(n_464),
.Y(n_499)
);

AOI221xp5_ASAP7_75t_L g500 ( 
.A1(n_468),
.A2(n_431),
.B1(n_442),
.B2(n_452),
.C(n_432),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_SL g501 ( 
.A(n_472),
.B(n_428),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_466),
.Y(n_502)
);

AOI22xp5_ASAP7_75t_L g503 ( 
.A1(n_492),
.A2(n_428),
.B1(n_380),
.B2(n_457),
.Y(n_503)
);

OAI32xp33_ASAP7_75t_L g504 ( 
.A1(n_472),
.A2(n_425),
.A3(n_426),
.B1(n_457),
.B2(n_453),
.Y(n_504)
);

OAI222xp33_ASAP7_75t_L g505 ( 
.A1(n_467),
.A2(n_453),
.B1(n_452),
.B2(n_455),
.C1(n_456),
.C2(n_372),
.Y(n_505)
);

AOI22xp5_ASAP7_75t_L g506 ( 
.A1(n_492),
.A2(n_380),
.B1(n_260),
.B2(n_359),
.Y(n_506)
);

AND2x2_ASAP7_75t_L g507 ( 
.A(n_462),
.B(n_455),
.Y(n_507)
);

AOI22xp5_ASAP7_75t_L g508 ( 
.A1(n_477),
.A2(n_380),
.B1(n_260),
.B2(n_370),
.Y(n_508)
);

AOI221xp5_ASAP7_75t_L g509 ( 
.A1(n_493),
.A2(n_377),
.B1(n_374),
.B2(n_386),
.C(n_383),
.Y(n_509)
);

NOR2x1_ASAP7_75t_L g510 ( 
.A(n_478),
.B(n_378),
.Y(n_510)
);

OR2x6_ASAP7_75t_L g511 ( 
.A(n_460),
.B(n_420),
.Y(n_511)
);

OAI21xp5_ASAP7_75t_SL g512 ( 
.A1(n_483),
.A2(n_236),
.B(n_271),
.Y(n_512)
);

OAI22xp33_ASAP7_75t_L g513 ( 
.A1(n_478),
.A2(n_378),
.B1(n_296),
.B2(n_283),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_473),
.B(n_422),
.Y(n_514)
);

AOI22xp5_ASAP7_75t_L g515 ( 
.A1(n_473),
.A2(n_380),
.B1(n_326),
.B2(n_422),
.Y(n_515)
);

AOI21xp33_ASAP7_75t_SL g516 ( 
.A1(n_482),
.A2(n_236),
.B(n_296),
.Y(n_516)
);

XOR2xp5_ASAP7_75t_L g517 ( 
.A(n_486),
.B(n_326),
.Y(n_517)
);

AOI211xp5_ASAP7_75t_L g518 ( 
.A1(n_482),
.A2(n_261),
.B(n_422),
.C(n_312),
.Y(n_518)
);

AOI32xp33_ASAP7_75t_L g519 ( 
.A1(n_463),
.A2(n_301),
.A3(n_292),
.B1(n_318),
.B2(n_316),
.Y(n_519)
);

NAND3xp33_ASAP7_75t_L g520 ( 
.A(n_485),
.B(n_296),
.C(n_261),
.Y(n_520)
);

OAI221xp5_ASAP7_75t_L g521 ( 
.A1(n_489),
.A2(n_316),
.B1(n_346),
.B2(n_347),
.C(n_351),
.Y(n_521)
);

OAI32xp33_ASAP7_75t_L g522 ( 
.A1(n_501),
.A2(n_490),
.A3(n_488),
.B1(n_474),
.B2(n_484),
.Y(n_522)
);

NOR2x1p5_ASAP7_75t_SL g523 ( 
.A(n_496),
.B(n_481),
.Y(n_523)
);

NOR2xp33_ASAP7_75t_L g524 ( 
.A(n_494),
.B(n_236),
.Y(n_524)
);

XOR2x2_ASAP7_75t_L g525 ( 
.A(n_499),
.B(n_465),
.Y(n_525)
);

INVx2_ASAP7_75t_L g526 ( 
.A(n_498),
.Y(n_526)
);

OAI221xp5_ASAP7_75t_L g527 ( 
.A1(n_495),
.A2(n_479),
.B1(n_469),
.B2(n_490),
.C(n_475),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_510),
.B(n_500),
.Y(n_528)
);

AOI221xp5_ASAP7_75t_L g529 ( 
.A1(n_504),
.A2(n_487),
.B1(n_470),
.B2(n_284),
.C(n_289),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_SL g530 ( 
.A(n_513),
.B(n_487),
.Y(n_530)
);

OAI22xp5_ASAP7_75t_L g531 ( 
.A1(n_508),
.A2(n_380),
.B1(n_475),
.B2(n_476),
.Y(n_531)
);

NAND4xp25_ASAP7_75t_L g532 ( 
.A(n_497),
.B(n_284),
.C(n_282),
.D(n_280),
.Y(n_532)
);

AOI21xp5_ASAP7_75t_L g533 ( 
.A1(n_512),
.A2(n_470),
.B(n_475),
.Y(n_533)
);

OAI22xp5_ASAP7_75t_SL g534 ( 
.A1(n_503),
.A2(n_515),
.B1(n_511),
.B2(n_517),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_514),
.B(n_476),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_502),
.Y(n_536)
);

AOI21xp5_ASAP7_75t_L g537 ( 
.A1(n_505),
.A2(n_476),
.B(n_351),
.Y(n_537)
);

OAI211xp5_ASAP7_75t_L g538 ( 
.A1(n_516),
.A2(n_347),
.B(n_280),
.C(n_289),
.Y(n_538)
);

OAI221xp5_ASAP7_75t_L g539 ( 
.A1(n_506),
.A2(n_519),
.B1(n_518),
.B2(n_521),
.C(n_509),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_SL g540 ( 
.A(n_507),
.B(n_283),
.Y(n_540)
);

NAND3xp33_ASAP7_75t_L g541 ( 
.A(n_520),
.B(n_283),
.C(n_305),
.Y(n_541)
);

NOR2xp33_ASAP7_75t_SL g542 ( 
.A(n_511),
.B(n_314),
.Y(n_542)
);

NAND3xp33_ASAP7_75t_L g543 ( 
.A(n_511),
.B(n_283),
.C(n_305),
.Y(n_543)
);

AOI32xp33_ASAP7_75t_L g544 ( 
.A1(n_500),
.A2(n_301),
.A3(n_292),
.B1(n_317),
.B2(n_305),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_L g545 ( 
.A(n_510),
.B(n_295),
.Y(n_545)
);

NAND4xp25_ASAP7_75t_L g546 ( 
.A(n_499),
.B(n_282),
.C(n_317),
.D(n_305),
.Y(n_546)
);

AOI222xp33_ASAP7_75t_L g547 ( 
.A1(n_525),
.A2(n_528),
.B1(n_539),
.B2(n_529),
.C1(n_534),
.C2(n_527),
.Y(n_547)
);

NAND5xp2_ASAP7_75t_L g548 ( 
.A(n_544),
.B(n_317),
.C(n_272),
.D(n_253),
.E(n_352),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_536),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_L g550 ( 
.A(n_546),
.B(n_301),
.Y(n_550)
);

NOR3xp33_ASAP7_75t_L g551 ( 
.A(n_546),
.B(n_250),
.C(n_293),
.Y(n_551)
);

NOR4xp25_ASAP7_75t_L g552 ( 
.A(n_530),
.B(n_293),
.C(n_253),
.D(n_314),
.Y(n_552)
);

NOR2x1_ASAP7_75t_L g553 ( 
.A(n_524),
.B(n_258),
.Y(n_553)
);

OAI211xp5_ASAP7_75t_L g554 ( 
.A1(n_522),
.A2(n_295),
.B(n_283),
.C(n_258),
.Y(n_554)
);

NOR2xp33_ASAP7_75t_L g555 ( 
.A(n_526),
.B(n_305),
.Y(n_555)
);

NAND3xp33_ASAP7_75t_L g556 ( 
.A(n_541),
.B(n_283),
.C(n_292),
.Y(n_556)
);

AOI21xp5_ASAP7_75t_SL g557 ( 
.A1(n_538),
.A2(n_293),
.B(n_258),
.Y(n_557)
);

NOR3xp33_ASAP7_75t_L g558 ( 
.A(n_532),
.B(n_250),
.C(n_301),
.Y(n_558)
);

AOI21xp5_ASAP7_75t_L g559 ( 
.A1(n_533),
.A2(n_292),
.B(n_301),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_L g560 ( 
.A(n_537),
.B(n_295),
.Y(n_560)
);

NOR2x1_ASAP7_75t_L g561 ( 
.A(n_543),
.B(n_302),
.Y(n_561)
);

OAI21xp5_ASAP7_75t_L g562 ( 
.A1(n_531),
.A2(n_266),
.B(n_234),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_L g563 ( 
.A(n_535),
.B(n_295),
.Y(n_563)
);

NAND4xp75_ASAP7_75t_L g564 ( 
.A(n_561),
.B(n_553),
.C(n_559),
.D(n_547),
.Y(n_564)
);

AND2x2_ASAP7_75t_L g565 ( 
.A(n_555),
.B(n_540),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_549),
.Y(n_566)
);

AND3x2_ASAP7_75t_L g567 ( 
.A(n_552),
.B(n_542),
.C(n_523),
.Y(n_567)
);

NAND4xp25_ASAP7_75t_L g568 ( 
.A(n_551),
.B(n_545),
.C(n_352),
.D(n_230),
.Y(n_568)
);

NOR3x1_ASAP7_75t_L g569 ( 
.A(n_554),
.B(n_274),
.C(n_283),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_L g570 ( 
.A(n_555),
.B(n_283),
.Y(n_570)
);

NOR3xp33_ASAP7_75t_L g571 ( 
.A(n_562),
.B(n_246),
.C(n_274),
.Y(n_571)
);

INVx2_ASAP7_75t_L g572 ( 
.A(n_550),
.Y(n_572)
);

NOR3x1_ASAP7_75t_L g573 ( 
.A(n_556),
.B(n_272),
.C(n_302),
.Y(n_573)
);

NOR2x1_ASAP7_75t_L g574 ( 
.A(n_548),
.B(n_246),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_560),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_563),
.Y(n_576)
);

NAND3xp33_ASAP7_75t_L g577 ( 
.A(n_558),
.B(n_319),
.C(n_348),
.Y(n_577)
);

AOI211x1_ASAP7_75t_L g578 ( 
.A1(n_557),
.A2(n_315),
.B(n_241),
.C(n_245),
.Y(n_578)
);

NOR2xp67_ASAP7_75t_L g579 ( 
.A(n_554),
.B(n_354),
.Y(n_579)
);

NAND4xp25_ASAP7_75t_L g580 ( 
.A(n_547),
.B(n_319),
.C(n_348),
.D(n_339),
.Y(n_580)
);

AND2x4_ASAP7_75t_L g581 ( 
.A(n_549),
.B(n_302),
.Y(n_581)
);

INVx2_ASAP7_75t_L g582 ( 
.A(n_566),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_565),
.Y(n_583)
);

NOR2x1_ASAP7_75t_L g584 ( 
.A(n_564),
.B(n_302),
.Y(n_584)
);

AO22x2_ASAP7_75t_L g585 ( 
.A1(n_572),
.A2(n_319),
.B1(n_308),
.B2(n_354),
.Y(n_585)
);

INVx1_ASAP7_75t_SL g586 ( 
.A(n_574),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_L g587 ( 
.A(n_580),
.B(n_302),
.Y(n_587)
);

NAND3xp33_ASAP7_75t_L g588 ( 
.A(n_567),
.B(n_319),
.C(n_308),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_581),
.Y(n_589)
);

INVx3_ASAP7_75t_L g590 ( 
.A(n_581),
.Y(n_590)
);

NOR4xp75_ASAP7_75t_SL g591 ( 
.A(n_570),
.B(n_299),
.C(n_315),
.D(n_354),
.Y(n_591)
);

BUFx6f_ASAP7_75t_L g592 ( 
.A(n_577),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_576),
.Y(n_593)
);

AOI22xp5_ASAP7_75t_L g594 ( 
.A1(n_568),
.A2(n_299),
.B1(n_339),
.B2(n_336),
.Y(n_594)
);

NOR2xp33_ASAP7_75t_L g595 ( 
.A(n_575),
.B(n_299),
.Y(n_595)
);

NOR2x1_ASAP7_75t_L g596 ( 
.A(n_579),
.B(n_573),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_582),
.Y(n_597)
);

INVx2_ASAP7_75t_L g598 ( 
.A(n_583),
.Y(n_598)
);

OAI22xp5_ASAP7_75t_L g599 ( 
.A1(n_588),
.A2(n_584),
.B1(n_586),
.B2(n_596),
.Y(n_599)
);

AND2x4_ASAP7_75t_L g600 ( 
.A(n_593),
.B(n_571),
.Y(n_600)
);

AND2x4_ASAP7_75t_L g601 ( 
.A(n_589),
.B(n_569),
.Y(n_601)
);

AOI21xp5_ASAP7_75t_L g602 ( 
.A1(n_592),
.A2(n_578),
.B(n_299),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_585),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_L g604 ( 
.A(n_592),
.B(n_578),
.Y(n_604)
);

XNOR2x1_ASAP7_75t_L g605 ( 
.A(n_594),
.B(n_592),
.Y(n_605)
);

AOI21xp5_ASAP7_75t_L g606 ( 
.A1(n_599),
.A2(n_595),
.B(n_587),
.Y(n_606)
);

AOI21xp5_ASAP7_75t_L g607 ( 
.A1(n_604),
.A2(n_590),
.B(n_585),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_598),
.Y(n_608)
);

XOR2x1_ASAP7_75t_L g609 ( 
.A(n_597),
.B(n_591),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_601),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_601),
.Y(n_611)
);

AO22x2_ASAP7_75t_L g612 ( 
.A1(n_605),
.A2(n_308),
.B1(n_348),
.B2(n_322),
.Y(n_612)
);

OAI21xp33_ASAP7_75t_L g613 ( 
.A1(n_610),
.A2(n_600),
.B(n_602),
.Y(n_613)
);

XOR2xp5_ASAP7_75t_L g614 ( 
.A(n_611),
.B(n_608),
.Y(n_614)
);

XNOR2xp5_ASAP7_75t_L g615 ( 
.A(n_606),
.B(n_603),
.Y(n_615)
);

OA22x2_ASAP7_75t_L g616 ( 
.A1(n_609),
.A2(n_339),
.B1(n_336),
.B2(n_333),
.Y(n_616)
);

OAI22xp5_ASAP7_75t_L g617 ( 
.A1(n_607),
.A2(n_333),
.B1(n_332),
.B2(n_330),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_612),
.Y(n_618)
);

AND2x2_ASAP7_75t_L g619 ( 
.A(n_610),
.B(n_299),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_614),
.Y(n_620)
);

XOR2xp5_ASAP7_75t_L g621 ( 
.A(n_615),
.B(n_308),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_613),
.Y(n_622)
);

INVx2_ASAP7_75t_L g623 ( 
.A(n_620),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_L g624 ( 
.A(n_622),
.B(n_619),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_623),
.B(n_621),
.Y(n_625)
);

OAI21xp5_ASAP7_75t_L g626 ( 
.A1(n_625),
.A2(n_624),
.B(n_617),
.Y(n_626)
);

OAI22xp33_ASAP7_75t_L g627 ( 
.A1(n_626),
.A2(n_618),
.B1(n_616),
.B2(n_322),
.Y(n_627)
);


endmodule