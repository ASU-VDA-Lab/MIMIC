module fake_jpeg_10756_n_613 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_613);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_613;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_543;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_170;
wire n_602;
wire n_313;
wire n_574;
wire n_542;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_292;
wire n_213;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_539;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_384;
wire n_296;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_599;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_17),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_16),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_9),
.Y(n_23)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_4),
.Y(n_25)
);

INVx11_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_12),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

INVx11_ASAP7_75t_SL g31 ( 
.A(n_8),
.Y(n_31)
);

BUFx12_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_10),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_2),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_12),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_7),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_3),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_4),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_16),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_2),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_15),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_12),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_1),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_1),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_1),
.Y(n_46)
);

CKINVDCx16_ASAP7_75t_R g47 ( 
.A(n_6),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_11),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_5),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_8),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_9),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_9),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_8),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_14),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_14),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_10),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_5),
.Y(n_57)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_13),
.Y(n_58)
);

INVx11_ASAP7_75t_L g59 ( 
.A(n_26),
.Y(n_59)
);

INVx8_ASAP7_75t_L g143 ( 
.A(n_59),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_32),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_60),
.B(n_68),
.Y(n_142)
);

INVx2_ASAP7_75t_SL g61 ( 
.A(n_22),
.Y(n_61)
);

HB1xp67_ASAP7_75t_L g135 ( 
.A(n_61),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_19),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_62),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_19),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_63),
.Y(n_131)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_48),
.Y(n_64)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_64),
.Y(n_128)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_18),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_65),
.Y(n_148)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_46),
.Y(n_66)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_66),
.Y(n_126)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_58),
.Y(n_67)
);

INVx5_ASAP7_75t_L g123 ( 
.A(n_67),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_20),
.B(n_17),
.Y(n_68)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_21),
.Y(n_69)
);

INVx5_ASAP7_75t_L g158 ( 
.A(n_69),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_19),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_70),
.Y(n_163)
);

OR2x2_ASAP7_75t_L g71 ( 
.A(n_28),
.B(n_17),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_71),
.B(n_87),
.Y(n_177)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_21),
.Y(n_72)
);

BUFx12f_ASAP7_75t_L g179 ( 
.A(n_72),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_19),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_73),
.Y(n_167)
);

BUFx3_ASAP7_75t_L g74 ( 
.A(n_21),
.Y(n_74)
);

BUFx12f_ASAP7_75t_L g192 ( 
.A(n_74),
.Y(n_192)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_36),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g178 ( 
.A(n_75),
.Y(n_178)
);

BUFx5_ASAP7_75t_L g76 ( 
.A(n_18),
.Y(n_76)
);

BUFx12f_ASAP7_75t_L g169 ( 
.A(n_76),
.Y(n_169)
);

BUFx5_ASAP7_75t_L g77 ( 
.A(n_18),
.Y(n_77)
);

INVx4_ASAP7_75t_L g138 ( 
.A(n_77),
.Y(n_138)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_46),
.Y(n_78)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_78),
.Y(n_127)
);

BUFx12f_ASAP7_75t_L g79 ( 
.A(n_48),
.Y(n_79)
);

INVx5_ASAP7_75t_L g159 ( 
.A(n_79),
.Y(n_159)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_28),
.Y(n_80)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_80),
.Y(n_134)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_39),
.Y(n_81)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_81),
.Y(n_140)
);

INVx5_ASAP7_75t_L g82 ( 
.A(n_58),
.Y(n_82)
);

INVx5_ASAP7_75t_L g184 ( 
.A(n_82),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_36),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g180 ( 
.A(n_83),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_36),
.Y(n_84)
);

INVx6_ASAP7_75t_L g146 ( 
.A(n_84),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_36),
.Y(n_85)
);

INVx6_ASAP7_75t_L g168 ( 
.A(n_85),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_18),
.Y(n_86)
);

INVx8_ASAP7_75t_L g194 ( 
.A(n_86),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_32),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_30),
.Y(n_88)
);

INVx3_ASAP7_75t_L g156 ( 
.A(n_88),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_30),
.Y(n_89)
);

INVx3_ASAP7_75t_L g172 ( 
.A(n_89),
.Y(n_172)
);

INVx8_ASAP7_75t_L g90 ( 
.A(n_30),
.Y(n_90)
);

INVx3_ASAP7_75t_L g173 ( 
.A(n_90),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_30),
.Y(n_91)
);

INVx3_ASAP7_75t_L g199 ( 
.A(n_91),
.Y(n_199)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_48),
.Y(n_92)
);

INVx3_ASAP7_75t_L g200 ( 
.A(n_92),
.Y(n_200)
);

INVx6_ASAP7_75t_L g93 ( 
.A(n_43),
.Y(n_93)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_93),
.Y(n_129)
);

INVx8_ASAP7_75t_L g94 ( 
.A(n_43),
.Y(n_94)
);

INVx4_ASAP7_75t_L g139 ( 
.A(n_94),
.Y(n_139)
);

HAxp5_ASAP7_75t_SL g95 ( 
.A(n_26),
.B(n_0),
.CON(n_95),
.SN(n_95)
);

OAI21xp33_ASAP7_75t_L g137 ( 
.A1(n_95),
.A2(n_0),
.B(n_1),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_43),
.Y(n_96)
);

INVx4_ASAP7_75t_L g141 ( 
.A(n_96),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_20),
.B(n_17),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g160 ( 
.A(n_97),
.B(n_98),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_29),
.B(n_16),
.Y(n_98)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_57),
.Y(n_99)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_99),
.Y(n_150)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_39),
.Y(n_100)
);

INVx4_ASAP7_75t_L g145 ( 
.A(n_100),
.Y(n_145)
);

BUFx3_ASAP7_75t_L g101 ( 
.A(n_42),
.Y(n_101)
);

INVx4_ASAP7_75t_L g149 ( 
.A(n_101),
.Y(n_149)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_39),
.Y(n_102)
);

INVx4_ASAP7_75t_L g155 ( 
.A(n_102),
.Y(n_155)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_57),
.Y(n_103)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_103),
.Y(n_154)
);

INVx8_ASAP7_75t_L g104 ( 
.A(n_43),
.Y(n_104)
);

INVx4_ASAP7_75t_L g171 ( 
.A(n_104),
.Y(n_171)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_57),
.Y(n_105)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_105),
.Y(n_176)
);

BUFx3_ASAP7_75t_L g106 ( 
.A(n_42),
.Y(n_106)
);

INVx4_ASAP7_75t_L g183 ( 
.A(n_106),
.Y(n_183)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_55),
.Y(n_107)
);

INVx4_ASAP7_75t_L g185 ( 
.A(n_107),
.Y(n_185)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_27),
.Y(n_108)
);

INVx4_ASAP7_75t_L g186 ( 
.A(n_108),
.Y(n_186)
);

BUFx5_ASAP7_75t_L g109 ( 
.A(n_55),
.Y(n_109)
);

INVx4_ASAP7_75t_L g190 ( 
.A(n_109),
.Y(n_190)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_42),
.Y(n_110)
);

INVx4_ASAP7_75t_L g202 ( 
.A(n_110),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_55),
.Y(n_111)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_111),
.Y(n_181)
);

BUFx5_ASAP7_75t_L g112 ( 
.A(n_55),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g162 ( 
.A(n_112),
.B(n_114),
.Y(n_162)
);

BUFx3_ASAP7_75t_L g113 ( 
.A(n_42),
.Y(n_113)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_113),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_29),
.B(n_15),
.Y(n_114)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_27),
.Y(n_115)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_115),
.Y(n_201)
);

INVx8_ASAP7_75t_L g116 ( 
.A(n_26),
.Y(n_116)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_116),
.Y(n_188)
);

BUFx3_ASAP7_75t_L g117 ( 
.A(n_42),
.Y(n_117)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_117),
.Y(n_191)
);

INVx4_ASAP7_75t_L g118 ( 
.A(n_54),
.Y(n_118)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_118),
.Y(n_136)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_27),
.Y(n_119)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_119),
.Y(n_147)
);

BUFx12f_ASAP7_75t_L g120 ( 
.A(n_49),
.Y(n_120)
);

INVx4_ASAP7_75t_SL g133 ( 
.A(n_120),
.Y(n_133)
);

INVx8_ASAP7_75t_L g121 ( 
.A(n_31),
.Y(n_121)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_121),
.Y(n_198)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_49),
.Y(n_122)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_122),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_71),
.B(n_35),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_125),
.B(n_164),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_65),
.A2(n_40),
.B1(n_24),
.B2(n_22),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_130),
.A2(n_152),
.B1(n_157),
.B2(n_175),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_93),
.A2(n_40),
.B1(n_24),
.B2(n_22),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_132),
.A2(n_144),
.B1(n_151),
.B2(n_153),
.Y(n_219)
);

OAI21xp33_ASAP7_75t_L g232 ( 
.A1(n_137),
.A2(n_0),
.B(n_1),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_86),
.A2(n_40),
.B1(n_24),
.B2(n_58),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_88),
.A2(n_49),
.B1(n_33),
.B2(n_35),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_69),
.A2(n_54),
.B1(n_38),
.B2(n_41),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_89),
.A2(n_56),
.B1(n_33),
.B2(n_38),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_SL g157 ( 
.A1(n_95),
.A2(n_54),
.B1(n_41),
.B2(n_44),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_59),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_SL g253 ( 
.A(n_161),
.B(n_2),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_61),
.B(n_56),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_81),
.B(n_44),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g255 ( 
.A(n_165),
.B(n_195),
.Y(n_255)
);

OAI22xp33_ASAP7_75t_L g166 ( 
.A1(n_62),
.A2(n_45),
.B1(n_53),
.B2(n_52),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_166),
.A2(n_174),
.B1(n_197),
.B2(n_199),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_100),
.B(n_23),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_170),
.B(n_182),
.Y(n_213)
);

OAI22xp33_ASAP7_75t_L g174 ( 
.A1(n_63),
.A2(n_45),
.B1(n_53),
.B2(n_52),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_91),
.A2(n_37),
.B1(n_25),
.B2(n_34),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_102),
.B(n_37),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_110),
.B(n_34),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_193),
.B(n_54),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_118),
.B(n_51),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_90),
.Y(n_196)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_196),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_96),
.A2(n_54),
.B1(n_25),
.B2(n_23),
.Y(n_197)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_129),
.Y(n_203)
);

INVx2_ASAP7_75t_L g288 ( 
.A(n_203),
.Y(n_288)
);

AOI22xp33_ASAP7_75t_L g204 ( 
.A1(n_166),
.A2(n_94),
.B1(n_104),
.B2(n_47),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_204),
.A2(n_224),
.B1(n_163),
.B2(n_167),
.Y(n_284)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_181),
.Y(n_205)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_205),
.Y(n_298)
);

OA22x2_ASAP7_75t_SL g209 ( 
.A1(n_137),
.A2(n_47),
.B1(n_120),
.B2(n_31),
.Y(n_209)
);

AO21x1_ASAP7_75t_L g325 ( 
.A1(n_209),
.A2(n_268),
.B(n_9),
.Y(n_325)
);

AOI22xp33_ASAP7_75t_SL g210 ( 
.A1(n_135),
.A2(n_121),
.B1(n_74),
.B2(n_72),
.Y(n_210)
);

INVxp67_ASAP7_75t_L g303 ( 
.A(n_210),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_142),
.B(n_79),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g315 ( 
.A(n_211),
.B(n_216),
.Y(n_315)
);

INVx6_ASAP7_75t_L g212 ( 
.A(n_124),
.Y(n_212)
);

INVx5_ASAP7_75t_L g331 ( 
.A(n_212),
.Y(n_331)
);

HB1xp67_ASAP7_75t_L g214 ( 
.A(n_135),
.Y(n_214)
);

INVxp67_ASAP7_75t_SL g304 ( 
.A(n_214),
.Y(n_304)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_150),
.Y(n_215)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_215),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_165),
.B(n_50),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_217),
.B(n_260),
.Y(n_278)
);

BUFx3_ASAP7_75t_L g218 ( 
.A(n_179),
.Y(n_218)
);

INVx4_ASAP7_75t_L g291 ( 
.A(n_218),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_157),
.A2(n_85),
.B1(n_73),
.B2(n_75),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_220),
.A2(n_225),
.B1(n_236),
.B2(n_251),
.Y(n_277)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_134),
.Y(n_221)
);

INVx1_ASAP7_75t_SL g305 ( 
.A(n_221),
.Y(n_305)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_198),
.Y(n_222)
);

INVx1_ASAP7_75t_SL g311 ( 
.A(n_222),
.Y(n_311)
);

CKINVDCx16_ASAP7_75t_R g223 ( 
.A(n_133),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g322 ( 
.A(n_223),
.B(n_229),
.Y(n_322)
);

AOI22xp33_ASAP7_75t_L g224 ( 
.A1(n_174),
.A2(n_107),
.B1(n_111),
.B2(n_70),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_195),
.A2(n_84),
.B1(n_83),
.B2(n_113),
.Y(n_225)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_154),
.Y(n_226)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_226),
.Y(n_283)
);

AND2x2_ASAP7_75t_L g227 ( 
.A(n_126),
.B(n_117),
.Y(n_227)
);

CKINVDCx16_ASAP7_75t_R g318 ( 
.A(n_227),
.Y(n_318)
);

BUFx12f_ASAP7_75t_L g228 ( 
.A(n_133),
.Y(n_228)
);

INVx4_ASAP7_75t_L g316 ( 
.A(n_228),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_142),
.B(n_79),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_160),
.B(n_50),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_230),
.B(n_246),
.Y(n_287)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_136),
.Y(n_231)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_231),
.Y(n_293)
);

AND2x2_ASAP7_75t_L g306 ( 
.A(n_232),
.B(n_241),
.Y(n_306)
);

BUFx3_ASAP7_75t_L g233 ( 
.A(n_179),
.Y(n_233)
);

INVx3_ASAP7_75t_L g276 ( 
.A(n_233),
.Y(n_276)
);

AND2x2_ASAP7_75t_L g234 ( 
.A(n_127),
.B(n_106),
.Y(n_234)
);

CKINVDCx16_ASAP7_75t_R g320 ( 
.A(n_234),
.Y(n_320)
);

INVx5_ASAP7_75t_L g235 ( 
.A(n_179),
.Y(n_235)
);

INVx3_ASAP7_75t_L g295 ( 
.A(n_235),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_177),
.A2(n_101),
.B1(n_120),
.B2(n_51),
.Y(n_236)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_176),
.Y(n_237)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_237),
.Y(n_309)
);

BUFx12f_ASAP7_75t_L g238 ( 
.A(n_124),
.Y(n_238)
);

INVx3_ASAP7_75t_L g296 ( 
.A(n_238),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_162),
.B(n_189),
.C(n_147),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_239),
.B(n_247),
.C(n_261),
.Y(n_286)
);

INVx3_ASAP7_75t_L g240 ( 
.A(n_139),
.Y(n_240)
);

INVx3_ASAP7_75t_L g313 ( 
.A(n_240),
.Y(n_313)
);

OAI21xp33_ASAP7_75t_L g241 ( 
.A1(n_162),
.A2(n_15),
.B(n_14),
.Y(n_241)
);

INVx2_ASAP7_75t_SL g242 ( 
.A(n_173),
.Y(n_242)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_242),
.Y(n_310)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_201),
.Y(n_243)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_243),
.Y(n_323)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_128),
.Y(n_244)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_244),
.Y(n_327)
);

OAI22xp33_ASAP7_75t_SL g245 ( 
.A1(n_152),
.A2(n_116),
.B1(n_32),
.B2(n_15),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_245),
.A2(n_274),
.B1(n_169),
.B2(n_192),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_177),
.Y(n_246)
);

AND2x2_ASAP7_75t_L g247 ( 
.A(n_140),
.B(n_0),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_160),
.B(n_14),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_248),
.B(n_253),
.Y(n_294)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_200),
.Y(n_249)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_249),
.Y(n_330)
);

BUFx6f_ASAP7_75t_L g250 ( 
.A(n_131),
.Y(n_250)
);

INVx3_ASAP7_75t_L g333 ( 
.A(n_250),
.Y(n_333)
);

OAI22xp5_ASAP7_75t_L g251 ( 
.A1(n_146),
.A2(n_32),
.B1(n_13),
.B2(n_12),
.Y(n_251)
);

BUFx6f_ASAP7_75t_L g252 ( 
.A(n_131),
.Y(n_252)
);

INVx11_ASAP7_75t_L g324 ( 
.A(n_252),
.Y(n_324)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_187),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_254),
.B(n_256),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_202),
.B(n_155),
.Y(n_256)
);

INVx3_ASAP7_75t_L g257 ( 
.A(n_171),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_257),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_145),
.B(n_13),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_258),
.B(n_259),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_194),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_186),
.B(n_11),
.Y(n_260)
);

AND2x2_ASAP7_75t_L g261 ( 
.A(n_191),
.B(n_2),
.Y(n_261)
);

AND2x2_ASAP7_75t_L g262 ( 
.A(n_149),
.B(n_2),
.Y(n_262)
);

OAI21xp5_ASAP7_75t_SL g285 ( 
.A1(n_262),
.A2(n_247),
.B(n_261),
.Y(n_285)
);

INVx5_ASAP7_75t_L g263 ( 
.A(n_192),
.Y(n_263)
);

INVxp67_ASAP7_75t_L g307 ( 
.A(n_263),
.Y(n_307)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_156),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_264),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_194),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_265),
.Y(n_314)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_172),
.Y(n_266)
);

INVxp67_ASAP7_75t_L g329 ( 
.A(n_266),
.Y(n_329)
);

AOI22xp33_ASAP7_75t_SL g267 ( 
.A1(n_158),
.A2(n_32),
.B1(n_11),
.B2(n_5),
.Y(n_267)
);

AOI22xp33_ASAP7_75t_SL g280 ( 
.A1(n_267),
.A2(n_269),
.B1(n_272),
.B2(n_273),
.Y(n_280)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_148),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_141),
.Y(n_270)
);

OR2x2_ASAP7_75t_L g302 ( 
.A(n_270),
.B(n_143),
.Y(n_302)
);

OAI22xp33_ASAP7_75t_L g271 ( 
.A1(n_185),
.A2(n_11),
.B1(n_4),
.B2(n_5),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g319 ( 
.A1(n_271),
.A2(n_167),
.B1(n_178),
.B2(n_143),
.Y(n_319)
);

AOI22xp33_ASAP7_75t_SL g272 ( 
.A1(n_123),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_272)
);

INVx3_ASAP7_75t_L g273 ( 
.A(n_159),
.Y(n_273)
);

CKINVDCx14_ASAP7_75t_R g274 ( 
.A(n_192),
.Y(n_274)
);

BUFx12f_ASAP7_75t_L g275 ( 
.A(n_163),
.Y(n_275)
);

AOI22xp33_ASAP7_75t_SL g299 ( 
.A1(n_275),
.A2(n_169),
.B1(n_190),
.B2(n_138),
.Y(n_299)
);

AOI21xp5_ASAP7_75t_L g279 ( 
.A1(n_206),
.A2(n_184),
.B(n_183),
.Y(n_279)
);

OAI21xp5_ASAP7_75t_SL g349 ( 
.A1(n_279),
.A2(n_328),
.B(n_335),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_217),
.B(n_168),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_281),
.B(n_290),
.Y(n_340)
);

OAI22xp5_ASAP7_75t_L g336 ( 
.A1(n_282),
.A2(n_319),
.B1(n_325),
.B2(n_334),
.Y(n_336)
);

AOI22xp33_ASAP7_75t_SL g338 ( 
.A1(n_284),
.A2(n_292),
.B1(n_225),
.B2(n_303),
.Y(n_338)
);

AND2x2_ASAP7_75t_L g353 ( 
.A(n_285),
.B(n_227),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_255),
.B(n_146),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_268),
.A2(n_148),
.B1(n_168),
.B2(n_180),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g344 ( 
.A1(n_292),
.A2(n_321),
.B1(n_271),
.B2(n_212),
.Y(n_344)
);

INVxp67_ASAP7_75t_L g362 ( 
.A(n_299),
.Y(n_362)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_213),
.B(n_188),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_300),
.B(n_262),
.C(n_234),
.Y(n_341)
);

INVx1_ASAP7_75t_SL g346 ( 
.A(n_302),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_261),
.B(n_239),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_312),
.B(n_326),
.Y(n_352)
);

OAI21xp5_ASAP7_75t_L g317 ( 
.A1(n_232),
.A2(n_180),
.B(n_178),
.Y(n_317)
);

OAI21xp5_ASAP7_75t_L g365 ( 
.A1(n_317),
.A2(n_218),
.B(n_233),
.Y(n_365)
);

OAI22xp5_ASAP7_75t_SL g321 ( 
.A1(n_219),
.A2(n_3),
.B1(n_4),
.B2(n_6),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_208),
.B(n_3),
.Y(n_326)
);

AOI21xp5_ASAP7_75t_L g328 ( 
.A1(n_209),
.A2(n_262),
.B(n_247),
.Y(n_328)
);

AOI22xp33_ASAP7_75t_L g334 ( 
.A1(n_220),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_334)
);

AOI22xp5_ASAP7_75t_SL g335 ( 
.A1(n_236),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_335)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_310),
.Y(n_337)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_337),
.Y(n_415)
);

OAI22xp5_ASAP7_75t_L g388 ( 
.A1(n_338),
.A2(n_344),
.B1(n_345),
.B2(n_348),
.Y(n_388)
);

XOR2xp5_ASAP7_75t_L g339 ( 
.A(n_312),
.B(n_241),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g401 ( 
.A(n_339),
.B(n_360),
.C(n_370),
.Y(n_401)
);

XNOR2xp5_ASAP7_75t_L g397 ( 
.A(n_341),
.B(n_371),
.Y(n_397)
);

OAI22xp5_ASAP7_75t_SL g342 ( 
.A1(n_325),
.A2(n_219),
.B1(n_209),
.B2(n_269),
.Y(n_342)
);

AOI22xp5_ASAP7_75t_L g404 ( 
.A1(n_342),
.A2(n_350),
.B1(n_380),
.B2(n_323),
.Y(n_404)
);

BUFx12f_ASAP7_75t_L g343 ( 
.A(n_289),
.Y(n_343)
);

BUFx6f_ASAP7_75t_L g410 ( 
.A(n_343),
.Y(n_410)
);

AOI22xp5_ASAP7_75t_L g345 ( 
.A1(n_321),
.A2(n_242),
.B1(n_234),
.B2(n_227),
.Y(n_345)
);

AOI22xp33_ASAP7_75t_SL g347 ( 
.A1(n_303),
.A2(n_242),
.B1(n_264),
.B2(n_266),
.Y(n_347)
);

INVxp67_ASAP7_75t_L g406 ( 
.A(n_347),
.Y(n_406)
);

AOI22xp5_ASAP7_75t_L g348 ( 
.A1(n_284),
.A2(n_277),
.B1(n_325),
.B2(n_281),
.Y(n_348)
);

OAI22xp5_ASAP7_75t_SL g350 ( 
.A1(n_277),
.A2(n_237),
.B1(n_226),
.B2(n_215),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_310),
.Y(n_351)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_351),
.Y(n_416)
);

XNOR2x1_ASAP7_75t_SL g386 ( 
.A(n_353),
.B(n_364),
.Y(n_386)
);

INVx2_ASAP7_75t_SL g354 ( 
.A(n_331),
.Y(n_354)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_354),
.Y(n_408)
);

AO22x1_ASAP7_75t_SL g355 ( 
.A1(n_328),
.A2(n_203),
.B1(n_205),
.B2(n_243),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_355),
.B(n_356),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_278),
.B(n_207),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_283),
.Y(n_357)
);

BUFx2_ASAP7_75t_L g413 ( 
.A(n_357),
.Y(n_413)
);

CKINVDCx20_ASAP7_75t_R g358 ( 
.A(n_301),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_SL g396 ( 
.A(n_358),
.B(n_359),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_SL g359 ( 
.A(n_287),
.B(n_254),
.Y(n_359)
);

XNOR2xp5_ASAP7_75t_L g360 ( 
.A(n_286),
.B(n_257),
.Y(n_360)
);

AOI22xp33_ASAP7_75t_SL g361 ( 
.A1(n_314),
.A2(n_304),
.B1(n_289),
.B2(n_313),
.Y(n_361)
);

INVxp67_ASAP7_75t_L g417 ( 
.A(n_361),
.Y(n_417)
);

AOI22xp5_ASAP7_75t_L g363 ( 
.A1(n_279),
.A2(n_240),
.B1(n_252),
.B2(n_250),
.Y(n_363)
);

OAI22xp5_ASAP7_75t_L g414 ( 
.A1(n_363),
.A2(n_368),
.B1(n_382),
.B2(n_316),
.Y(n_414)
);

AND2x2_ASAP7_75t_L g364 ( 
.A(n_317),
.B(n_228),
.Y(n_364)
);

AO21x1_ASAP7_75t_L g395 ( 
.A1(n_365),
.A2(n_307),
.B(n_329),
.Y(n_395)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_283),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_SL g383 ( 
.A(n_366),
.B(n_378),
.Y(n_383)
);

AND2x2_ASAP7_75t_L g367 ( 
.A(n_332),
.B(n_228),
.Y(n_367)
);

OAI21xp5_ASAP7_75t_SL g412 ( 
.A1(n_367),
.A2(n_374),
.B(n_298),
.Y(n_412)
);

AOI22xp5_ASAP7_75t_L g368 ( 
.A1(n_290),
.A2(n_273),
.B1(n_263),
.B2(n_235),
.Y(n_368)
);

NAND3xp33_ASAP7_75t_L g369 ( 
.A(n_294),
.B(n_238),
.C(n_275),
.Y(n_369)
);

HAxp5_ASAP7_75t_SL g405 ( 
.A(n_369),
.B(n_372),
.CON(n_405),
.SN(n_405)
);

MAJIxp5_ASAP7_75t_L g370 ( 
.A(n_286),
.B(n_238),
.C(n_275),
.Y(n_370)
);

MAJIxp5_ASAP7_75t_L g371 ( 
.A(n_300),
.B(n_315),
.C(n_278),
.Y(n_371)
);

NAND3xp33_ASAP7_75t_L g372 ( 
.A(n_322),
.B(n_326),
.C(n_285),
.Y(n_372)
);

INVx2_ASAP7_75t_L g373 ( 
.A(n_288),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_373),
.B(n_381),
.Y(n_387)
);

OAI21xp5_ASAP7_75t_SL g374 ( 
.A1(n_306),
.A2(n_320),
.B(n_318),
.Y(n_374)
);

XOR2xp5_ASAP7_75t_L g375 ( 
.A(n_306),
.B(n_320),
.Y(n_375)
);

XNOR2xp5_ASAP7_75t_L g403 ( 
.A(n_375),
.B(n_376),
.Y(n_403)
);

XOR2xp5_ASAP7_75t_L g376 ( 
.A(n_306),
.B(n_318),
.Y(n_376)
);

CKINVDCx20_ASAP7_75t_R g377 ( 
.A(n_324),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_SL g392 ( 
.A(n_377),
.B(n_329),
.Y(n_392)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_309),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_309),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_SL g399 ( 
.A(n_379),
.B(n_327),
.Y(n_399)
);

OAI22xp5_ASAP7_75t_L g380 ( 
.A1(n_335),
.A2(n_319),
.B1(n_282),
.B2(n_314),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_302),
.B(n_297),
.Y(n_381)
);

AOI22xp5_ASAP7_75t_L g382 ( 
.A1(n_305),
.A2(n_311),
.B1(n_293),
.B2(n_330),
.Y(n_382)
);

OAI22xp5_ASAP7_75t_SL g384 ( 
.A1(n_348),
.A2(n_344),
.B1(n_340),
.B2(n_346),
.Y(n_384)
);

AOI22xp5_ASAP7_75t_L g445 ( 
.A1(n_384),
.A2(n_389),
.B1(n_391),
.B2(n_393),
.Y(n_445)
);

OAI22xp5_ASAP7_75t_SL g389 ( 
.A1(n_340),
.A2(n_280),
.B1(n_302),
.B2(n_305),
.Y(n_389)
);

CKINVDCx20_ASAP7_75t_R g390 ( 
.A(n_382),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_L g438 ( 
.A(n_390),
.B(n_392),
.Y(n_438)
);

OAI22xp5_ASAP7_75t_SL g391 ( 
.A1(n_346),
.A2(n_311),
.B1(n_293),
.B2(n_333),
.Y(n_391)
);

OAI22xp5_ASAP7_75t_SL g393 ( 
.A1(n_342),
.A2(n_333),
.B1(n_331),
.B2(n_330),
.Y(n_393)
);

CKINVDCx20_ASAP7_75t_R g394 ( 
.A(n_381),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_394),
.B(n_399),
.Y(n_425)
);

INVx1_ASAP7_75t_SL g428 ( 
.A(n_395),
.Y(n_428)
);

OAI22xp5_ASAP7_75t_SL g398 ( 
.A1(n_345),
.A2(n_327),
.B1(n_297),
.B2(n_323),
.Y(n_398)
);

AOI22xp5_ASAP7_75t_L g459 ( 
.A1(n_398),
.A2(n_407),
.B1(n_411),
.B2(n_419),
.Y(n_459)
);

CKINVDCx20_ASAP7_75t_R g400 ( 
.A(n_367),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_400),
.B(n_409),
.Y(n_434)
);

AOI22xp5_ASAP7_75t_SL g402 ( 
.A1(n_364),
.A2(n_307),
.B1(n_295),
.B2(n_316),
.Y(n_402)
);

AOI21xp5_ASAP7_75t_L g454 ( 
.A1(n_402),
.A2(n_354),
.B(n_291),
.Y(n_454)
);

OAI22xp5_ASAP7_75t_L g448 ( 
.A1(n_404),
.A2(n_357),
.B1(n_378),
.B2(n_366),
.Y(n_448)
);

OAI22xp5_ASAP7_75t_SL g407 ( 
.A1(n_356),
.A2(n_313),
.B1(n_308),
.B2(n_324),
.Y(n_407)
);

CKINVDCx20_ASAP7_75t_R g409 ( 
.A(n_367),
.Y(n_409)
);

OAI22xp5_ASAP7_75t_SL g411 ( 
.A1(n_352),
.A2(n_308),
.B1(n_298),
.B2(n_288),
.Y(n_411)
);

AND2x2_ASAP7_75t_L g441 ( 
.A(n_412),
.B(n_414),
.Y(n_441)
);

INVx4_ASAP7_75t_SL g418 ( 
.A(n_365),
.Y(n_418)
);

INVx4_ASAP7_75t_L g453 ( 
.A(n_418),
.Y(n_453)
);

OAI22xp5_ASAP7_75t_SL g419 ( 
.A1(n_352),
.A2(n_295),
.B1(n_276),
.B2(n_296),
.Y(n_419)
);

XNOR2xp5_ASAP7_75t_SL g420 ( 
.A(n_360),
.B(n_291),
.Y(n_420)
);

XNOR2xp5_ASAP7_75t_L g424 ( 
.A(n_420),
.B(n_376),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_371),
.B(n_276),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_421),
.B(n_422),
.Y(n_439)
);

CKINVDCx16_ASAP7_75t_R g422 ( 
.A(n_364),
.Y(n_422)
);

OAI32xp33_ASAP7_75t_L g423 ( 
.A1(n_355),
.A2(n_349),
.A3(n_350),
.B1(n_374),
.B2(n_337),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_423),
.B(n_385),
.Y(n_443)
);

XOR2xp5_ASAP7_75t_L g460 ( 
.A(n_424),
.B(n_403),
.Y(n_460)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_383),
.Y(n_426)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_426),
.Y(n_484)
);

CKINVDCx20_ASAP7_75t_R g427 ( 
.A(n_383),
.Y(n_427)
);

CKINVDCx20_ASAP7_75t_R g461 ( 
.A(n_427),
.Y(n_461)
);

XNOR2xp5_ASAP7_75t_L g429 ( 
.A(n_397),
.B(n_339),
.Y(n_429)
);

MAJIxp5_ASAP7_75t_L g469 ( 
.A(n_429),
.B(n_430),
.C(n_440),
.Y(n_469)
);

MAJIxp5_ASAP7_75t_L g430 ( 
.A(n_401),
.B(n_370),
.C(n_375),
.Y(n_430)
);

AOI22xp33_ASAP7_75t_L g431 ( 
.A1(n_393),
.A2(n_362),
.B1(n_336),
.B2(n_351),
.Y(n_431)
);

OAI22xp5_ASAP7_75t_L g472 ( 
.A1(n_431),
.A2(n_443),
.B1(n_455),
.B2(n_395),
.Y(n_472)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_387),
.Y(n_432)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_432),
.Y(n_463)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_387),
.Y(n_433)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_433),
.Y(n_473)
);

OAI22xp5_ASAP7_75t_SL g435 ( 
.A1(n_404),
.A2(n_349),
.B1(n_363),
.B2(n_362),
.Y(n_435)
);

AOI22xp5_ASAP7_75t_L g465 ( 
.A1(n_435),
.A2(n_436),
.B1(n_437),
.B2(n_448),
.Y(n_465)
);

OAI22xp5_ASAP7_75t_SL g436 ( 
.A1(n_394),
.A2(n_368),
.B1(n_341),
.B2(n_355),
.Y(n_436)
);

OAI22x1_ASAP7_75t_SL g437 ( 
.A1(n_388),
.A2(n_384),
.B1(n_418),
.B2(n_423),
.Y(n_437)
);

XNOR2xp5_ASAP7_75t_L g440 ( 
.A(n_397),
.B(n_353),
.Y(n_440)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_399),
.Y(n_442)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_442),
.Y(n_477)
);

CKINVDCx20_ASAP7_75t_R g444 ( 
.A(n_396),
.Y(n_444)
);

CKINVDCx20_ASAP7_75t_R g466 ( 
.A(n_444),
.Y(n_466)
);

CKINVDCx20_ASAP7_75t_R g446 ( 
.A(n_419),
.Y(n_446)
);

CKINVDCx20_ASAP7_75t_R g474 ( 
.A(n_446),
.Y(n_474)
);

CKINVDCx20_ASAP7_75t_R g447 ( 
.A(n_407),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_447),
.B(n_450),
.Y(n_468)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_415),
.Y(n_449)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_449),
.Y(n_480)
);

OA21x2_ASAP7_75t_L g450 ( 
.A1(n_385),
.A2(n_353),
.B(n_354),
.Y(n_450)
);

XNOR2xp5_ASAP7_75t_L g451 ( 
.A(n_401),
.B(n_379),
.Y(n_451)
);

MAJIxp5_ASAP7_75t_L g481 ( 
.A(n_451),
.B(n_457),
.C(n_386),
.Y(n_481)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_415),
.Y(n_452)
);

INVx1_ASAP7_75t_SL g464 ( 
.A(n_452),
.Y(n_464)
);

AND2x2_ASAP7_75t_L g483 ( 
.A(n_454),
.B(n_412),
.Y(n_483)
);

OAI22xp5_ASAP7_75t_L g455 ( 
.A1(n_390),
.A2(n_417),
.B1(n_395),
.B2(n_388),
.Y(n_455)
);

OAI32xp33_ASAP7_75t_L g456 ( 
.A1(n_421),
.A2(n_296),
.A3(n_343),
.B1(n_373),
.B2(n_398),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_456),
.B(n_409),
.Y(n_471)
);

XNOR2xp5_ASAP7_75t_L g457 ( 
.A(n_403),
.B(n_343),
.Y(n_457)
);

CKINVDCx20_ASAP7_75t_R g458 ( 
.A(n_411),
.Y(n_458)
);

CKINVDCx20_ASAP7_75t_R g479 ( 
.A(n_458),
.Y(n_479)
);

XNOR2xp5_ASAP7_75t_SL g507 ( 
.A(n_460),
.B(n_459),
.Y(n_507)
);

INVxp67_ASAP7_75t_L g462 ( 
.A(n_439),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g511 ( 
.A(n_462),
.B(n_453),
.Y(n_511)
);

NOR2xp67_ASAP7_75t_SL g467 ( 
.A(n_457),
.B(n_420),
.Y(n_467)
);

OAI21xp5_ASAP7_75t_SL g505 ( 
.A1(n_467),
.A2(n_483),
.B(n_481),
.Y(n_505)
);

NOR2xp67_ASAP7_75t_L g470 ( 
.A(n_442),
.B(n_405),
.Y(n_470)
);

NOR2xp33_ASAP7_75t_L g514 ( 
.A(n_470),
.B(n_489),
.Y(n_514)
);

AO21x1_ASAP7_75t_L g513 ( 
.A1(n_471),
.A2(n_459),
.B(n_449),
.Y(n_513)
);

AOI22xp5_ASAP7_75t_L g501 ( 
.A1(n_472),
.A2(n_476),
.B1(n_441),
.B2(n_450),
.Y(n_501)
);

AOI22xp5_ASAP7_75t_L g475 ( 
.A1(n_437),
.A2(n_389),
.B1(n_414),
.B2(n_422),
.Y(n_475)
);

OAI22xp5_ASAP7_75t_SL g497 ( 
.A1(n_475),
.A2(n_482),
.B1(n_445),
.B2(n_428),
.Y(n_497)
);

OAI22xp5_ASAP7_75t_SL g476 ( 
.A1(n_445),
.A2(n_406),
.B1(n_418),
.B2(n_400),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_425),
.B(n_426),
.Y(n_478)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_478),
.Y(n_492)
);

MAJIxp5_ASAP7_75t_L g503 ( 
.A(n_481),
.B(n_491),
.C(n_436),
.Y(n_503)
);

AOI22xp5_ASAP7_75t_L g482 ( 
.A1(n_441),
.A2(n_391),
.B1(n_416),
.B2(n_392),
.Y(n_482)
);

XOR2xp5_ASAP7_75t_L g485 ( 
.A(n_429),
.B(n_386),
.Y(n_485)
);

XOR2xp5_ASAP7_75t_L g493 ( 
.A(n_485),
.B(n_486),
.Y(n_493)
);

XNOR2xp5_ASAP7_75t_L g486 ( 
.A(n_440),
.B(n_402),
.Y(n_486)
);

XNOR2x2_ASAP7_75t_SL g487 ( 
.A(n_424),
.B(n_416),
.Y(n_487)
);

OAI211xp5_ASAP7_75t_SL g506 ( 
.A1(n_487),
.A2(n_456),
.B(n_441),
.C(n_454),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g488 ( 
.A(n_425),
.B(n_413),
.Y(n_488)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_488),
.Y(n_495)
);

NAND3xp33_ASAP7_75t_L g489 ( 
.A(n_439),
.B(n_343),
.C(n_413),
.Y(n_489)
);

XNOR2xp5_ASAP7_75t_L g490 ( 
.A(n_451),
.B(n_408),
.Y(n_490)
);

XOR2xp5_ASAP7_75t_L g504 ( 
.A(n_490),
.B(n_491),
.Y(n_504)
);

MAJIxp5_ASAP7_75t_L g491 ( 
.A(n_430),
.B(n_434),
.C(n_450),
.Y(n_491)
);

AOI22xp33_ASAP7_75t_L g494 ( 
.A1(n_461),
.A2(n_435),
.B1(n_447),
.B2(n_438),
.Y(n_494)
);

OAI22xp5_ASAP7_75t_L g526 ( 
.A1(n_494),
.A2(n_499),
.B1(n_512),
.B2(n_513),
.Y(n_526)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_488),
.Y(n_496)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_496),
.Y(n_523)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_497),
.Y(n_520)
);

NOR3xp33_ASAP7_75t_SL g498 ( 
.A(n_466),
.B(n_434),
.C(n_428),
.Y(n_498)
);

CKINVDCx14_ASAP7_75t_R g522 ( 
.A(n_498),
.Y(n_522)
);

CKINVDCx20_ASAP7_75t_R g499 ( 
.A(n_478),
.Y(n_499)
);

OAI22xp5_ASAP7_75t_L g500 ( 
.A1(n_465),
.A2(n_433),
.B1(n_432),
.B2(n_443),
.Y(n_500)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_500),
.Y(n_527)
);

OAI22xp5_ASAP7_75t_SL g533 ( 
.A1(n_501),
.A2(n_475),
.B1(n_471),
.B2(n_482),
.Y(n_533)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_480),
.Y(n_502)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_502),
.Y(n_528)
);

XNOR2xp5_ASAP7_75t_L g524 ( 
.A(n_503),
.B(n_504),
.Y(n_524)
);

XOR2xp5_ASAP7_75t_L g535 ( 
.A(n_505),
.B(n_516),
.Y(n_535)
);

XNOR2xp5_ASAP7_75t_SL g539 ( 
.A(n_506),
.B(n_507),
.Y(n_539)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_480),
.Y(n_508)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_508),
.Y(n_529)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_477),
.Y(n_509)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_509),
.Y(n_537)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_477),
.Y(n_510)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_510),
.Y(n_542)
);

CKINVDCx16_ASAP7_75t_R g521 ( 
.A(n_511),
.Y(n_521)
);

CKINVDCx20_ASAP7_75t_R g512 ( 
.A(n_468),
.Y(n_512)
);

MAJIxp5_ASAP7_75t_L g515 ( 
.A(n_469),
.B(n_452),
.C(n_453),
.Y(n_515)
);

MAJIxp5_ASAP7_75t_L g525 ( 
.A(n_515),
.B(n_490),
.C(n_486),
.Y(n_525)
);

XOR2xp5_ASAP7_75t_L g516 ( 
.A(n_469),
.B(n_460),
.Y(n_516)
);

NOR2xp33_ASAP7_75t_SL g517 ( 
.A(n_484),
.B(n_410),
.Y(n_517)
);

CKINVDCx14_ASAP7_75t_R g534 ( 
.A(n_517),
.Y(n_534)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_464),
.Y(n_518)
);

OAI22xp5_ASAP7_75t_L g531 ( 
.A1(n_518),
.A2(n_519),
.B1(n_462),
.B2(n_512),
.Y(n_531)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_464),
.Y(n_519)
);

MAJIxp5_ASAP7_75t_L g557 ( 
.A(n_525),
.B(n_540),
.C(n_518),
.Y(n_557)
);

MAJIxp5_ASAP7_75t_L g530 ( 
.A(n_515),
.B(n_485),
.C(n_487),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_SL g551 ( 
.A(n_530),
.B(n_532),
.Y(n_551)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_531),
.Y(n_546)
);

MAJIxp5_ASAP7_75t_L g532 ( 
.A(n_504),
.B(n_476),
.C(n_465),
.Y(n_532)
);

AOI22xp33_ASAP7_75t_SL g545 ( 
.A1(n_533),
.A2(n_497),
.B1(n_492),
.B2(n_506),
.Y(n_545)
);

XOR2xp5_ASAP7_75t_L g536 ( 
.A(n_493),
.B(n_483),
.Y(n_536)
);

XOR2xp5_ASAP7_75t_L g558 ( 
.A(n_536),
.B(n_541),
.Y(n_558)
);

XNOR2xp5_ASAP7_75t_L g538 ( 
.A(n_503),
.B(n_483),
.Y(n_538)
);

XNOR2xp5_ASAP7_75t_L g553 ( 
.A(n_538),
.B(n_507),
.Y(n_553)
);

MAJIxp5_ASAP7_75t_L g540 ( 
.A(n_516),
.B(n_473),
.C(n_463),
.Y(n_540)
);

XOR2xp5_ASAP7_75t_L g541 ( 
.A(n_493),
.B(n_468),
.Y(n_541)
);

FAx1_ASAP7_75t_SL g543 ( 
.A(n_539),
.B(n_532),
.CI(n_500),
.CON(n_543),
.SN(n_543)
);

OR2x2_ASAP7_75t_L g577 ( 
.A(n_543),
.B(n_554),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_L g544 ( 
.A(n_528),
.B(n_519),
.Y(n_544)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_544),
.Y(n_576)
);

OAI22xp5_ASAP7_75t_SL g563 ( 
.A1(n_545),
.A2(n_520),
.B1(n_521),
.B2(n_539),
.Y(n_563)
);

AOI21xp5_ASAP7_75t_L g547 ( 
.A1(n_526),
.A2(n_514),
.B(n_513),
.Y(n_547)
);

AOI21xp5_ASAP7_75t_L g566 ( 
.A1(n_547),
.A2(n_550),
.B(n_556),
.Y(n_566)
);

OAI22xp5_ASAP7_75t_SL g548 ( 
.A1(n_527),
.A2(n_513),
.B1(n_501),
.B2(n_492),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_L g574 ( 
.A(n_548),
.B(n_549),
.Y(n_574)
);

CKINVDCx14_ASAP7_75t_R g549 ( 
.A(n_522),
.Y(n_549)
);

OR2x2_ASAP7_75t_L g550 ( 
.A(n_523),
.B(n_463),
.Y(n_550)
);

NOR2xp33_ASAP7_75t_L g552 ( 
.A(n_540),
.B(n_479),
.Y(n_552)
);

NOR2xp33_ASAP7_75t_SL g567 ( 
.A(n_552),
.B(n_538),
.Y(n_567)
);

XNOR2xp5_ASAP7_75t_L g573 ( 
.A(n_553),
.B(n_555),
.Y(n_573)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_528),
.Y(n_554)
);

XNOR2xp5_ASAP7_75t_L g555 ( 
.A(n_524),
.B(n_505),
.Y(n_555)
);

OAI21xp5_ASAP7_75t_L g556 ( 
.A1(n_533),
.A2(n_499),
.B(n_495),
.Y(n_556)
);

NOR2xp33_ASAP7_75t_L g569 ( 
.A(n_557),
.B(n_559),
.Y(n_569)
);

OAI22xp5_ASAP7_75t_SL g559 ( 
.A1(n_527),
.A2(n_496),
.B1(n_495),
.B2(n_511),
.Y(n_559)
);

OAI22xp5_ASAP7_75t_L g560 ( 
.A1(n_520),
.A2(n_474),
.B1(n_473),
.B2(n_498),
.Y(n_560)
);

XOR2xp5_ASAP7_75t_L g565 ( 
.A(n_560),
.B(n_510),
.Y(n_565)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_529),
.Y(n_561)
);

NOR2xp33_ASAP7_75t_L g570 ( 
.A(n_561),
.B(n_517),
.Y(n_570)
);

MAJIxp5_ASAP7_75t_L g562 ( 
.A(n_557),
.B(n_524),
.C(n_525),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_L g581 ( 
.A(n_562),
.B(n_570),
.Y(n_581)
);

AND2x2_ASAP7_75t_L g586 ( 
.A(n_563),
.B(n_548),
.Y(n_586)
);

OAI21xp5_ASAP7_75t_SL g564 ( 
.A1(n_547),
.A2(n_534),
.B(n_530),
.Y(n_564)
);

AOI21xp5_ASAP7_75t_L g579 ( 
.A1(n_564),
.A2(n_568),
.B(n_571),
.Y(n_579)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_565),
.Y(n_578)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_567),
.Y(n_589)
);

OAI21xp5_ASAP7_75t_SL g568 ( 
.A1(n_546),
.A2(n_509),
.B(n_529),
.Y(n_568)
);

AOI21xp5_ASAP7_75t_L g571 ( 
.A1(n_546),
.A2(n_541),
.B(n_536),
.Y(n_571)
);

MAJIxp5_ASAP7_75t_L g572 ( 
.A(n_555),
.B(n_535),
.C(n_537),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_L g584 ( 
.A(n_572),
.B(n_575),
.Y(n_584)
);

MAJIxp5_ASAP7_75t_L g575 ( 
.A(n_558),
.B(n_535),
.C(n_537),
.Y(n_575)
);

NOR2xp33_ASAP7_75t_SL g580 ( 
.A(n_569),
.B(n_562),
.Y(n_580)
);

NOR2xp33_ASAP7_75t_SL g597 ( 
.A(n_580),
.B(n_572),
.Y(n_597)
);

OAI22xp5_ASAP7_75t_SL g582 ( 
.A1(n_566),
.A2(n_556),
.B1(n_550),
.B2(n_560),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_L g593 ( 
.A(n_582),
.B(n_583),
.Y(n_593)
);

NOR2xp33_ASAP7_75t_L g583 ( 
.A(n_574),
.B(n_543),
.Y(n_583)
);

NOR2xp33_ASAP7_75t_L g585 ( 
.A(n_574),
.B(n_543),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_L g596 ( 
.A(n_585),
.B(n_586),
.Y(n_596)
);

HB1xp67_ASAP7_75t_L g587 ( 
.A(n_566),
.Y(n_587)
);

HB1xp67_ASAP7_75t_L g591 ( 
.A(n_587),
.Y(n_591)
);

OAI22xp5_ASAP7_75t_SL g588 ( 
.A1(n_577),
.A2(n_551),
.B1(n_561),
.B2(n_554),
.Y(n_588)
);

INVxp67_ASAP7_75t_L g590 ( 
.A(n_588),
.Y(n_590)
);

NOR2xp33_ASAP7_75t_L g592 ( 
.A(n_581),
.B(n_584),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_SL g603 ( 
.A(n_592),
.B(n_594),
.Y(n_603)
);

XOR2xp5_ASAP7_75t_L g594 ( 
.A(n_588),
.B(n_573),
.Y(n_594)
);

AOI21xp5_ASAP7_75t_L g595 ( 
.A1(n_579),
.A2(n_564),
.B(n_577),
.Y(n_595)
);

AOI21xp5_ASAP7_75t_L g599 ( 
.A1(n_595),
.A2(n_597),
.B(n_598),
.Y(n_599)
);

OAI21xp5_ASAP7_75t_SL g598 ( 
.A1(n_579),
.A2(n_575),
.B(n_571),
.Y(n_598)
);

AOI21xp5_ASAP7_75t_L g600 ( 
.A1(n_593),
.A2(n_589),
.B(n_586),
.Y(n_600)
);

OAI21x1_ASAP7_75t_L g606 ( 
.A1(n_600),
.A2(n_602),
.B(n_604),
.Y(n_606)
);

MAJIxp5_ASAP7_75t_L g601 ( 
.A(n_596),
.B(n_578),
.C(n_576),
.Y(n_601)
);

MAJIxp5_ASAP7_75t_L g605 ( 
.A(n_601),
.B(n_573),
.C(n_565),
.Y(n_605)
);

AOI21xp5_ASAP7_75t_L g602 ( 
.A1(n_590),
.A2(n_591),
.B(n_568),
.Y(n_602)
);

O2A1O1Ixp33_ASAP7_75t_SL g604 ( 
.A1(n_591),
.A2(n_582),
.B(n_559),
.C(n_563),
.Y(n_604)
);

MAJIxp5_ASAP7_75t_L g608 ( 
.A(n_605),
.B(n_607),
.C(n_599),
.Y(n_608)
);

MAJIxp5_ASAP7_75t_L g607 ( 
.A(n_603),
.B(n_544),
.C(n_558),
.Y(n_607)
);

MAJIxp5_ASAP7_75t_L g610 ( 
.A(n_608),
.B(n_609),
.C(n_542),
.Y(n_610)
);

AOI321xp33_ASAP7_75t_L g609 ( 
.A1(n_606),
.A2(n_542),
.A3(n_502),
.B1(n_508),
.B2(n_553),
.C(n_410),
.Y(n_609)
);

MAJIxp5_ASAP7_75t_L g611 ( 
.A(n_610),
.B(n_410),
.C(n_413),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_611),
.Y(n_612)
);

NOR2xp33_ASAP7_75t_L g613 ( 
.A(n_612),
.B(n_408),
.Y(n_613)
);


endmodule