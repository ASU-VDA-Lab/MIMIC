module fake_jpeg_8233_n_256 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_256);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_256;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_192;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_14),
.Y(n_15)
);

BUFx5_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

INVx4_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_5),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

INVx6_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

BUFx16f_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_0),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

INVx11_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

INVx2_ASAP7_75t_SL g28 ( 
.A(n_10),
.Y(n_28)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_13),
.B(n_4),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

INVx11_ASAP7_75t_L g32 ( 
.A(n_26),
.Y(n_32)
);

INVx11_ASAP7_75t_L g46 ( 
.A(n_32),
.Y(n_46)
);

OR2x2_ASAP7_75t_L g33 ( 
.A(n_20),
.B(n_0),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_33),
.B(n_36),
.Y(n_45)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_23),
.Y(n_34)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_34),
.Y(n_57)
);

AOI21xp33_ASAP7_75t_L g35 ( 
.A1(n_23),
.A2(n_0),
.B(n_1),
.Y(n_35)
);

AND2x2_ASAP7_75t_L g52 ( 
.A(n_35),
.B(n_3),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_30),
.B(n_2),
.Y(n_36)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_31),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_37),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_26),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_27),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_39),
.B(n_40),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_23),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_23),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_41),
.B(n_25),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_26),
.Y(n_42)
);

INVx2_ASAP7_75t_SL g50 ( 
.A(n_42),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g43 ( 
.A1(n_39),
.A2(n_22),
.B1(n_27),
.B2(n_29),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_43),
.A2(n_44),
.B1(n_54),
.B2(n_55),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g44 ( 
.A1(n_39),
.A2(n_22),
.B1(n_27),
.B2(n_29),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_33),
.B(n_25),
.Y(n_48)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_48),
.B(n_58),
.Y(n_72)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_32),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_49),
.B(n_51),
.Y(n_75)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_32),
.Y(n_51)
);

A2O1A1Ixp33_ASAP7_75t_L g71 ( 
.A1(n_52),
.A2(n_63),
.B(n_36),
.C(n_24),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_35),
.A2(n_22),
.B1(n_28),
.B2(n_29),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_37),
.A2(n_28),
.B1(n_18),
.B2(n_16),
.Y(n_55)
);

AND2x2_ASAP7_75t_SL g58 ( 
.A(n_34),
.B(n_16),
.Y(n_58)
);

INVx2_ASAP7_75t_SL g59 ( 
.A(n_34),
.Y(n_59)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_59),
.Y(n_70)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_38),
.Y(n_60)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_60),
.Y(n_74)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_61),
.Y(n_78)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_38),
.Y(n_62)
);

INVx1_ASAP7_75t_SL g69 ( 
.A(n_62),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_33),
.B(n_30),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_L g64 ( 
.A1(n_37),
.A2(n_28),
.B1(n_18),
.B2(n_24),
.Y(n_64)
);

OAI22xp33_ASAP7_75t_L g81 ( 
.A1(n_64),
.A2(n_18),
.B1(n_20),
.B2(n_21),
.Y(n_81)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_38),
.Y(n_65)
);

HAxp5_ASAP7_75t_SL g67 ( 
.A(n_65),
.B(n_42),
.CON(n_67),
.SN(n_67)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_46),
.Y(n_66)
);

INVx11_ASAP7_75t_L g109 ( 
.A(n_66),
.Y(n_109)
);

OAI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_67),
.A2(n_85),
.B1(n_86),
.B2(n_51),
.Y(n_91)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_56),
.Y(n_68)
);

BUFx2_ASAP7_75t_SL g92 ( 
.A(n_68),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_71),
.B(n_63),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_53),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_73),
.B(n_76),
.Y(n_105)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_46),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_53),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_77),
.B(n_83),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_46),
.Y(n_79)
);

INVxp33_ASAP7_75t_L g108 ( 
.A(n_79),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_56),
.Y(n_80)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_80),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_L g93 ( 
.A1(n_81),
.A2(n_47),
.B1(n_50),
.B2(n_49),
.Y(n_93)
);

INVx13_ASAP7_75t_L g83 ( 
.A(n_59),
.Y(n_83)
);

BUFx12f_ASAP7_75t_L g84 ( 
.A(n_59),
.Y(n_84)
);

CKINVDCx16_ASAP7_75t_R g90 ( 
.A(n_84),
.Y(n_90)
);

INVx8_ASAP7_75t_L g85 ( 
.A(n_56),
.Y(n_85)
);

INVx8_ASAP7_75t_L g86 ( 
.A(n_50),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_72),
.B(n_52),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_87),
.B(n_98),
.Y(n_123)
);

INVx13_ASAP7_75t_L g88 ( 
.A(n_84),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_88),
.B(n_97),
.Y(n_116)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_72),
.B(n_54),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g113 ( 
.A(n_89),
.B(n_58),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_L g111 ( 
.A1(n_91),
.A2(n_93),
.B1(n_68),
.B2(n_85),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_82),
.A2(n_52),
.B1(n_47),
.B2(n_62),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_94),
.A2(n_57),
.B1(n_69),
.B2(n_17),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_78),
.A2(n_65),
.B1(n_60),
.B2(n_50),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_95),
.A2(n_96),
.B1(n_104),
.B2(n_83),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_78),
.A2(n_71),
.B1(n_72),
.B2(n_66),
.Y(n_96)
);

INVx13_ASAP7_75t_L g97 ( 
.A(n_84),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_75),
.B(n_48),
.Y(n_98)
);

INVx13_ASAP7_75t_L g99 ( 
.A(n_84),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_99),
.B(n_100),
.Y(n_119)
);

BUFx24_ASAP7_75t_SL g100 ( 
.A(n_70),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g120 ( 
.A(n_101),
.B(n_106),
.Y(n_120)
);

NOR3xp33_ASAP7_75t_L g102 ( 
.A(n_81),
.B(n_45),
.C(n_67),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_102),
.B(n_19),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_76),
.A2(n_61),
.B1(n_57),
.B2(n_58),
.Y(n_104)
);

OR2x2_ASAP7_75t_L g106 ( 
.A(n_86),
.B(n_45),
.Y(n_106)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_105),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_110),
.B(n_115),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_111),
.B(n_125),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_87),
.B(n_58),
.C(n_70),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_112),
.B(n_114),
.C(n_122),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_SL g144 ( 
.A(n_113),
.B(n_129),
.Y(n_144)
);

XOR2xp5_ASAP7_75t_L g114 ( 
.A(n_96),
.B(n_41),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_109),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_101),
.B(n_33),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_117),
.B(n_124),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_118),
.A2(n_130),
.B1(n_92),
.B2(n_57),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_SL g121 ( 
.A(n_106),
.B(n_98),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_121),
.B(n_126),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_89),
.B(n_74),
.C(n_69),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_109),
.Y(n_124)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_105),
.Y(n_125)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_109),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_127),
.B(n_128),
.Y(n_147)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_95),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_SL g129 ( 
.A1(n_94),
.A2(n_74),
.B(n_41),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_89),
.B(n_41),
.C(n_40),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_131),
.B(n_112),
.C(n_129),
.Y(n_152)
);

CKINVDCx14_ASAP7_75t_R g132 ( 
.A(n_107),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_132),
.B(n_99),
.Y(n_149)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_116),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_133),
.B(n_135),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_L g134 ( 
.A1(n_120),
.A2(n_107),
.B(n_106),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_SL g158 ( 
.A1(n_134),
.A2(n_143),
.B(n_110),
.Y(n_158)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_121),
.Y(n_135)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_115),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_137),
.B(n_140),
.Y(n_159)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_124),
.Y(n_140)
);

XOR2xp5_ASAP7_75t_L g141 ( 
.A(n_114),
.B(n_104),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_141),
.B(n_152),
.C(n_154),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_L g143 ( 
.A1(n_120),
.A2(n_17),
.B(n_21),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_127),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_145),
.B(n_155),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_146),
.A2(n_130),
.B1(n_99),
.B2(n_97),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_123),
.B(n_79),
.Y(n_148)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_148),
.Y(n_157)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_149),
.Y(n_162)
);

OR2x2_ASAP7_75t_L g150 ( 
.A(n_128),
.B(n_15),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_150),
.B(n_15),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_123),
.B(n_90),
.Y(n_153)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_153),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_131),
.B(n_90),
.C(n_92),
.Y(n_154)
);

CKINVDCx16_ASAP7_75t_R g155 ( 
.A(n_118),
.Y(n_155)
);

CKINVDCx14_ASAP7_75t_R g179 ( 
.A(n_158),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_L g160 ( 
.A1(n_134),
.A2(n_122),
.B(n_125),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_SL g193 ( 
.A(n_160),
.B(n_25),
.Y(n_193)
);

INVx8_ASAP7_75t_L g161 ( 
.A(n_145),
.Y(n_161)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_161),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_164),
.A2(n_170),
.B1(n_146),
.B2(n_142),
.Y(n_182)
);

HB1xp67_ASAP7_75t_L g165 ( 
.A(n_137),
.Y(n_165)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_165),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_166),
.B(n_172),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_135),
.B(n_113),
.Y(n_167)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_167),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_147),
.A2(n_113),
.B1(n_103),
.B2(n_88),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_153),
.B(n_148),
.Y(n_171)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_171),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_136),
.Y(n_172)
);

CKINVDCx16_ASAP7_75t_R g173 ( 
.A(n_139),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_173),
.B(n_174),
.Y(n_186)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_140),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_133),
.B(n_108),
.Y(n_175)
);

INVxp67_ASAP7_75t_L g184 ( 
.A(n_175),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_141),
.B(n_119),
.Y(n_176)
);

FAx1_ASAP7_75t_L g194 ( 
.A(n_176),
.B(n_19),
.CI(n_25),
.CON(n_194),
.SN(n_194)
);

BUFx6f_ASAP7_75t_L g177 ( 
.A(n_161),
.Y(n_177)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_177),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_168),
.B(n_138),
.C(n_152),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_180),
.B(n_185),
.C(n_188),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_182),
.A2(n_192),
.B1(n_195),
.B2(n_184),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_168),
.B(n_138),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_160),
.B(n_144),
.Y(n_188)
);

AO22x1_ASAP7_75t_L g190 ( 
.A1(n_158),
.A2(n_144),
.B1(n_151),
.B2(n_150),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_190),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_176),
.B(n_154),
.C(n_151),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_191),
.B(n_156),
.C(n_172),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_169),
.A2(n_143),
.B1(n_97),
.B2(n_88),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_SL g199 ( 
.A(n_193),
.B(n_195),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_194),
.B(n_170),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_SL g195 ( 
.A(n_167),
.B(n_3),
.Y(n_195)
);

AOI21xp5_ASAP7_75t_L g198 ( 
.A1(n_179),
.A2(n_159),
.B(n_156),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_SL g211 ( 
.A1(n_198),
.A2(n_203),
.B(n_206),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_200),
.B(n_205),
.C(n_209),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_202),
.A2(n_162),
.B1(n_31),
.B2(n_19),
.Y(n_219)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_186),
.Y(n_203)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_204),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_185),
.B(n_157),
.C(n_171),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_187),
.Y(n_206)
);

OAI321xp33_ASAP7_75t_L g207 ( 
.A1(n_190),
.A2(n_194),
.A3(n_173),
.B1(n_164),
.B2(n_163),
.C(n_193),
.Y(n_207)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_207),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_178),
.B(n_161),
.Y(n_208)
);

BUFx24_ASAP7_75t_SL g214 ( 
.A(n_208),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_188),
.B(n_157),
.C(n_159),
.Y(n_209)
);

BUFx2_ASAP7_75t_L g210 ( 
.A(n_177),
.Y(n_210)
);

BUFx10_ASAP7_75t_L g217 ( 
.A(n_210),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_L g213 ( 
.A1(n_205),
.A2(n_174),
.B(n_184),
.Y(n_213)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_213),
.Y(n_230)
);

A2O1A1Ixp33_ASAP7_75t_L g215 ( 
.A1(n_201),
.A2(n_183),
.B(n_189),
.C(n_163),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_215),
.B(n_199),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_197),
.B(n_194),
.C(n_181),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_216),
.B(n_218),
.C(n_221),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_197),
.B(n_162),
.C(n_166),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_219),
.A2(n_220),
.B1(n_25),
.B2(n_19),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_196),
.A2(n_31),
.B1(n_42),
.B2(n_80),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_209),
.B(n_41),
.Y(n_221)
);

INVx11_ASAP7_75t_L g224 ( 
.A(n_217),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_224),
.B(n_214),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_218),
.B(n_200),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_225),
.B(n_231),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_226),
.B(n_227),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_223),
.B(n_210),
.Y(n_227)
);

A2O1A1Ixp33_ASAP7_75t_SL g228 ( 
.A1(n_222),
.A2(n_199),
.B(n_42),
.C(n_41),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_228),
.A2(n_233),
.B1(n_6),
.B2(n_7),
.Y(n_234)
);

FAx1_ASAP7_75t_SL g232 ( 
.A(n_215),
.B(n_40),
.CI(n_13),
.CON(n_232),
.SN(n_232)
);

BUFx24_ASAP7_75t_SL g240 ( 
.A(n_232),
.Y(n_240)
);

AO22x1_ASAP7_75t_L g233 ( 
.A1(n_211),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_233)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_234),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_235),
.B(n_238),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_224),
.B(n_212),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_237),
.B(n_230),
.Y(n_243)
);

INVxp33_ASAP7_75t_L g238 ( 
.A(n_232),
.Y(n_238)
);

OAI21xp5_ASAP7_75t_L g239 ( 
.A1(n_229),
.A2(n_212),
.B(n_216),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_239),
.B(n_229),
.C(n_236),
.Y(n_242)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_242),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_243),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_241),
.B(n_221),
.Y(n_244)
);

AOI322xp5_ASAP7_75t_L g248 ( 
.A1(n_244),
.A2(n_246),
.A3(n_228),
.B1(n_217),
.B2(n_40),
.C1(n_12),
.C2(n_7),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_240),
.A2(n_228),
.B1(n_233),
.B2(n_217),
.Y(n_246)
);

BUFx24_ASAP7_75t_SL g252 ( 
.A(n_248),
.Y(n_252)
);

AOI322xp5_ASAP7_75t_L g251 ( 
.A1(n_245),
.A2(n_12),
.A3(n_9),
.B1(n_10),
.B2(n_11),
.C1(n_8),
.C2(n_40),
.Y(n_251)
);

A2O1A1O1Ixp25_ASAP7_75t_L g253 ( 
.A1(n_251),
.A2(n_245),
.B(n_247),
.C(n_10),
.D(n_11),
.Y(n_253)
);

NAND3xp33_ASAP7_75t_L g254 ( 
.A(n_253),
.B(n_8),
.C(n_9),
.Y(n_254)
);

O2A1O1Ixp33_ASAP7_75t_SL g255 ( 
.A1(n_254),
.A2(n_252),
.B(n_250),
.C(n_8),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_SL g256 ( 
.A(n_255),
.B(n_249),
.Y(n_256)
);


endmodule