module fake_jpeg_9682_n_103 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_103);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_103;

wire n_10;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_9;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g9 ( 
.A(n_7),
.Y(n_9)
);

INVx1_ASAP7_75t_L g10 ( 
.A(n_5),
.Y(n_10)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_8),
.Y(n_11)
);

BUFx12f_ASAP7_75t_L g12 ( 
.A(n_2),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_0),
.Y(n_13)
);

INVx6_ASAP7_75t_L g14 ( 
.A(n_0),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_5),
.Y(n_15)
);

BUFx10_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_5),
.B(n_4),
.Y(n_18)
);

BUFx16f_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_18),
.B(n_1),
.Y(n_20)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_20),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_18),
.B(n_1),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_21),
.B(n_22),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_10),
.B(n_1),
.Y(n_22)
);

BUFx24_ASAP7_75t_L g23 ( 
.A(n_19),
.Y(n_23)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_23),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_24),
.Y(n_34)
);

INVx3_ASAP7_75t_SL g25 ( 
.A(n_19),
.Y(n_25)
);

CKINVDCx14_ASAP7_75t_R g33 ( 
.A(n_25),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_19),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_26),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_9),
.B(n_2),
.Y(n_27)
);

AND2x2_ASAP7_75t_L g31 ( 
.A(n_27),
.B(n_10),
.Y(n_31)
);

NAND3xp33_ASAP7_75t_L g42 ( 
.A(n_31),
.B(n_35),
.C(n_36),
.Y(n_42)
);

AND2x2_ASAP7_75t_L g35 ( 
.A(n_25),
.B(n_19),
.Y(n_35)
);

AOI32xp33_ASAP7_75t_L g36 ( 
.A1(n_25),
.A2(n_14),
.A3(n_19),
.B1(n_15),
.B2(n_13),
.Y(n_36)
);

CKINVDCx12_ASAP7_75t_R g37 ( 
.A(n_23),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_37),
.B(n_26),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_31),
.B(n_22),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_38),
.B(n_44),
.Y(n_50)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_39),
.B(n_40),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_35),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_L g41 ( 
.A1(n_36),
.A2(n_14),
.B1(n_10),
.B2(n_13),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_41),
.A2(n_14),
.B1(n_11),
.B2(n_9),
.Y(n_57)
);

HB1xp67_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_43),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_32),
.B(n_20),
.Y(n_44)
);

INVxp67_ASAP7_75t_L g53 ( 
.A(n_45),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_29),
.B(n_27),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_46),
.B(n_47),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_29),
.B(n_21),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_28),
.B(n_15),
.Y(n_48)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_48),
.Y(n_51)
);

OAI21xp5_ASAP7_75t_L g49 ( 
.A1(n_39),
.A2(n_32),
.B(n_28),
.Y(n_49)
);

AOI21xp5_ASAP7_75t_L g62 ( 
.A1(n_49),
.A2(n_54),
.B(n_38),
.Y(n_62)
);

OAI21xp5_ASAP7_75t_L g54 ( 
.A1(n_40),
.A2(n_33),
.B(n_35),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_57),
.B(n_58),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_41),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_42),
.A2(n_30),
.B1(n_11),
.B2(n_24),
.Y(n_59)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_59),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g60 ( 
.A(n_50),
.B(n_54),
.C(n_49),
.Y(n_60)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_60),
.B(n_63),
.C(n_59),
.Y(n_72)
);

OAI21xp5_ASAP7_75t_L g76 ( 
.A1(n_62),
.A2(n_16),
.B(n_17),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g63 ( 
.A(n_50),
.B(n_44),
.C(n_26),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_56),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_64),
.B(n_65),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_55),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_51),
.B(n_34),
.Y(n_67)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_67),
.Y(n_78)
);

AND2x2_ASAP7_75t_L g68 ( 
.A(n_52),
.B(n_23),
.Y(n_68)
);

AOI21xp5_ASAP7_75t_L g71 ( 
.A1(n_68),
.A2(n_53),
.B(n_23),
.Y(n_71)
);

OAI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_58),
.A2(n_30),
.B1(n_16),
.B2(n_17),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_69),
.A2(n_55),
.B1(n_57),
.B2(n_37),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_61),
.B(n_51),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_70),
.B(n_74),
.Y(n_82)
);

XOR2xp5_ASAP7_75t_L g85 ( 
.A(n_71),
.B(n_76),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_72),
.B(n_73),
.C(n_66),
.Y(n_79)
);

XNOR2xp5_ASAP7_75t_L g73 ( 
.A(n_60),
.B(n_62),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_63),
.B(n_53),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_75),
.B(n_26),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_79),
.B(n_80),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_73),
.B(n_66),
.C(n_68),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_78),
.B(n_77),
.Y(n_81)
);

OAI21xp5_ASAP7_75t_SL g89 ( 
.A1(n_81),
.A2(n_84),
.B(n_16),
.Y(n_89)
);

OR2x2_ASAP7_75t_L g91 ( 
.A(n_83),
.B(n_2),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_75),
.Y(n_84)
);

AOI31xp33_ASAP7_75t_L g86 ( 
.A1(n_72),
.A2(n_68),
.A3(n_76),
.B(n_26),
.Y(n_86)
);

OAI221xp5_ASAP7_75t_L g90 ( 
.A1(n_86),
.A2(n_17),
.B1(n_12),
.B2(n_16),
.C(n_24),
.Y(n_90)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_82),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_87),
.B(n_89),
.Y(n_93)
);

NAND3xp33_ASAP7_75t_L g94 ( 
.A(n_90),
.B(n_3),
.C(n_4),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_91),
.B(n_3),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_85),
.A2(n_3),
.B1(n_4),
.B2(n_6),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_95),
.B(n_96),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_88),
.B(n_79),
.C(n_80),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_L g97 ( 
.A1(n_93),
.A2(n_92),
.B(n_91),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_SL g100 ( 
.A1(n_97),
.A2(n_17),
.B(n_12),
.Y(n_100)
);

AOI321xp33_ASAP7_75t_L g99 ( 
.A1(n_98),
.A2(n_12),
.A3(n_16),
.B1(n_17),
.B2(n_94),
.C(n_96),
.Y(n_99)
);

NOR2x1_ASAP7_75t_L g102 ( 
.A(n_99),
.B(n_12),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_100),
.B(n_16),
.Y(n_101)
);

XOR2xp5_ASAP7_75t_L g103 ( 
.A(n_101),
.B(n_102),
.Y(n_103)
);


endmodule