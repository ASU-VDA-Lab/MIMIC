module fake_netlist_1_3018_n_926 (n_117, n_219, n_44, n_133, n_149, n_220, n_81, n_69, n_214, n_204, n_221, n_185, n_22, n_203, n_57, n_88, n_52, n_26, n_50, n_33, n_102, n_73, n_49, n_119, n_141, n_115, n_97, n_80, n_167, n_107, n_158, n_60, n_114, n_121, n_41, n_35, n_94, n_65, n_171, n_196, n_125, n_192, n_9, n_161, n_10, n_177, n_130, n_189, n_103, n_19, n_87, n_137, n_180, n_104, n_160, n_98, n_74, n_206, n_154, n_7, n_29, n_195, n_165, n_146, n_45, n_85, n_181, n_101, n_62, n_36, n_47, n_215, n_37, n_34, n_5, n_23, n_8, n_91, n_108, n_116, n_155, n_209, n_217, n_139, n_16, n_13, n_198, n_169, n_193, n_152, n_113, n_95, n_124, n_156, n_128, n_120, n_129, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_135, n_42, n_188, n_24, n_78, n_197, n_201, n_6, n_4, n_127, n_170, n_40, n_111, n_157, n_79, n_202, n_210, n_38, n_64, n_142, n_184, n_191, n_200, n_46, n_31, n_208, n_211, n_58, n_122, n_187, n_138, n_126, n_178, n_118, n_32, n_0, n_179, n_84, n_131, n_112, n_55, n_205, n_12, n_86, n_143, n_213, n_182, n_166, n_162, n_186, n_75, n_163, n_226, n_105, n_159, n_174, n_227, n_72, n_136, n_43, n_76, n_89, n_176, n_68, n_144, n_27, n_53, n_183, n_67, n_77, n_216, n_20, n_2, n_147, n_199, n_54, n_148, n_123, n_83, n_172, n_28, n_48, n_100, n_212, n_92, n_11, n_223, n_25, n_30, n_59, n_150, n_218, n_168, n_194, n_3, n_18, n_110, n_66, n_134, n_222, n_1, n_164, n_82, n_106, n_175, n_15, n_173, n_190, n_145, n_153, n_61, n_21, n_99, n_109, n_93, n_132, n_151, n_51, n_140, n_207, n_224, n_96, n_225, n_39, n_926);
input n_117;
input n_219;
input n_44;
input n_133;
input n_149;
input n_220;
input n_81;
input n_69;
input n_214;
input n_204;
input n_221;
input n_185;
input n_22;
input n_203;
input n_57;
input n_88;
input n_52;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_119;
input n_141;
input n_115;
input n_97;
input n_80;
input n_167;
input n_107;
input n_158;
input n_60;
input n_114;
input n_121;
input n_41;
input n_35;
input n_94;
input n_65;
input n_171;
input n_196;
input n_125;
input n_192;
input n_9;
input n_161;
input n_10;
input n_177;
input n_130;
input n_189;
input n_103;
input n_19;
input n_87;
input n_137;
input n_180;
input n_104;
input n_160;
input n_98;
input n_74;
input n_206;
input n_154;
input n_7;
input n_29;
input n_195;
input n_165;
input n_146;
input n_45;
input n_85;
input n_181;
input n_101;
input n_62;
input n_36;
input n_47;
input n_215;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_108;
input n_116;
input n_155;
input n_209;
input n_217;
input n_139;
input n_16;
input n_13;
input n_198;
input n_169;
input n_193;
input n_152;
input n_113;
input n_95;
input n_124;
input n_156;
input n_128;
input n_120;
input n_129;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_135;
input n_42;
input n_188;
input n_24;
input n_78;
input n_197;
input n_201;
input n_6;
input n_4;
input n_127;
input n_170;
input n_40;
input n_111;
input n_157;
input n_79;
input n_202;
input n_210;
input n_38;
input n_64;
input n_142;
input n_184;
input n_191;
input n_200;
input n_46;
input n_31;
input n_208;
input n_211;
input n_58;
input n_122;
input n_187;
input n_138;
input n_126;
input n_178;
input n_118;
input n_32;
input n_0;
input n_179;
input n_84;
input n_131;
input n_112;
input n_55;
input n_205;
input n_12;
input n_86;
input n_143;
input n_213;
input n_182;
input n_166;
input n_162;
input n_186;
input n_75;
input n_163;
input n_226;
input n_105;
input n_159;
input n_174;
input n_227;
input n_72;
input n_136;
input n_43;
input n_76;
input n_89;
input n_176;
input n_68;
input n_144;
input n_27;
input n_53;
input n_183;
input n_67;
input n_77;
input n_216;
input n_20;
input n_2;
input n_147;
input n_199;
input n_54;
input n_148;
input n_123;
input n_83;
input n_172;
input n_28;
input n_48;
input n_100;
input n_212;
input n_92;
input n_11;
input n_223;
input n_25;
input n_30;
input n_59;
input n_150;
input n_218;
input n_168;
input n_194;
input n_3;
input n_18;
input n_110;
input n_66;
input n_134;
input n_222;
input n_1;
input n_164;
input n_82;
input n_106;
input n_175;
input n_15;
input n_173;
input n_190;
input n_145;
input n_153;
input n_61;
input n_21;
input n_99;
input n_109;
input n_93;
input n_132;
input n_151;
input n_51;
input n_140;
input n_207;
input n_224;
input n_96;
input n_225;
input n_39;
output n_926;
wire n_663;
wire n_707;
wire n_791;
wire n_361;
wire n_513;
wire n_838;
wire n_705;
wire n_603;
wire n_604;
wire n_858;
wire n_590;
wire n_407;
wire n_885;
wire n_755;
wire n_646;
wire n_792;
wire n_284;
wire n_278;
wire n_500;
wire n_925;
wire n_848;
wire n_607;
wire n_808;
wire n_829;
wire n_431;
wire n_484;
wire n_862;
wire n_852;
wire n_496;
wire n_667;
wire n_311;
wire n_801;
wire n_292;
wire n_309;
wire n_701;
wire n_612;
wire n_328;
wire n_655;
wire n_468;
wire n_743;
wire n_917;
wire n_523;
wire n_903;
wire n_920;
wire n_229;
wire n_757;
wire n_750;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_770;
wire n_918;
wire n_252;
wire n_878;
wire n_814;
wire n_911;
wire n_637;
wire n_817;
wire n_802;
wire n_856;
wire n_353;
wire n_564;
wire n_779;
wire n_528;
wire n_288;
wire n_383;
wire n_904;
wire n_661;
wire n_850;
wire n_762;
wire n_672;
wire n_532;
wire n_627;
wire n_758;
wire n_544;
wire n_890;
wire n_400;
wire n_787;
wire n_853;
wire n_296;
wire n_765;
wire n_386;
wire n_432;
wire n_659;
wire n_807;
wire n_877;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_896;
wire n_334;
wire n_783;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_715;
wire n_463;
wire n_789;
wire n_330;
wire n_587;
wire n_662;
wire n_678;
wire n_387;
wire n_476;
wire n_434;
wire n_384;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_812;
wire n_598;
wire n_489;
wire n_777;
wire n_732;
wire n_752;
wire n_351;
wire n_860;
wire n_401;
wire n_461;
wire n_305;
wire n_599;
wire n_228;
wire n_786;
wire n_724;
wire n_857;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_922;
wire n_234;
wire n_465;
wire n_796;
wire n_609;
wire n_636;
wire n_914;
wire n_909;
wire n_366;
wire n_596;
wire n_286;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_773;
wire n_847;
wire n_840;
wire n_392;
wire n_668;
wire n_846;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_563;
wire n_540;
wire n_638;
wire n_830;
wire n_560;
wire n_517;
wire n_479;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_726;
wire n_780;
wire n_712;
wire n_447;
wire n_872;
wire n_608;
wire n_897;
wire n_567;
wire n_809;
wire n_888;
wire n_580;
wire n_502;
wire n_921;
wire n_543;
wire n_854;
wire n_455;
wire n_312;
wire n_529;
wire n_630;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_865;
wire n_915;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_764;
wire n_314;
wire n_237;
wire n_255;
wire n_426;
wire n_624;
wire n_725;
wire n_769;
wire n_818;
wire n_844;
wire n_230;
wire n_274;
wire n_738;
wire n_282;
wire n_319;
wire n_499;
wire n_895;
wire n_417;
wire n_798;
wire n_241;
wire n_575;
wire n_238;
wire n_711;
wire n_318;
wire n_884;
wire n_887;
wire n_471;
wire n_632;
wire n_767;
wire n_828;
wire n_293;
wire n_506;
wire n_533;
wire n_393;
wire n_490;
wire n_247;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_826;
wire n_304;
wire n_399;
wire n_892;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_863;
wire n_322;
wire n_310;
wire n_907;
wire n_708;
wire n_307;
wire n_634;
wire n_610;
wire n_730;
wire n_696;
wire n_735;
wire n_771;
wire n_784;
wire n_474;
wire n_354;
wire n_402;
wire n_893;
wire n_413;
wire n_676;
wire n_391;
wire n_910;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_813;
wire n_352;
wire n_746;
wire n_619;
wire n_882;
wire n_268;
wire n_501;
wire n_248;
wire n_871;
wire n_803;
wire n_299;
wire n_338;
wire n_519;
wire n_699;
wire n_729;
wire n_805;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_849;
wire n_864;
wire n_810;
wire n_329;
wire n_251;
wire n_747;
wire n_635;
wire n_889;
wire n_731;
wire n_689;
wire n_905;
wire n_902;
wire n_525;
wire n_876;
wire n_886;
wire n_507;
wire n_605;
wire n_719;
wire n_704;
wire n_611;
wire n_633;
wire n_873;
wire n_271;
wire n_760;
wire n_751;
wire n_800;
wire n_626;
wire n_302;
wire n_466;
wire n_900;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_259;
wire n_308;
wire n_546;
wire n_412;
wire n_664;
wire n_827;
wire n_565;
wire n_788;
wire n_475;
wire n_578;
wire n_542;
wire n_537;
wire n_660;
wire n_430;
wire n_839;
wire n_450;
wire n_579;
wire n_776;
wire n_879;
wire n_403;
wire n_557;
wire n_516;
wire n_842;
wire n_254;
wire n_549;
wire n_622;
wire n_832;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_768;
wire n_869;
wire n_797;
wire n_285;
wire n_420;
wire n_446;
wire n_423;
wire n_342;
wire n_621;
wire n_666;
wire n_880;
wire n_799;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_874;
wire n_388;
wire n_454;
wire n_687;
wire n_273;
wire n_505;
wire n_706;
wire n_822;
wire n_823;
wire n_390;
wire n_682;
wire n_514;
wire n_486;
wire n_906;
wire n_720;
wire n_568;
wire n_245;
wire n_357;
wire n_653;
wire n_716;
wire n_881;
wire n_260;
wire n_806;
wire n_539;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_718;
wire n_536;
wire n_816;
wire n_265;
wire n_264;
wire n_522;
wire n_883;
wire n_573;
wire n_898;
wire n_673;
wire n_669;
wire n_754;
wire n_775;
wire n_616;
wire n_365;
wire n_717;
wire n_541;
wire n_409;
wire n_315;
wire n_363;
wire n_733;
wire n_861;
wire n_899;
wire n_295;
wire n_654;
wire n_263;
wire n_894;
wire n_495;
wire n_428;
wire n_364;
wire n_566;
wire n_794;
wire n_376;
wire n_639;
wire n_552;
wire n_744;
wire n_677;
wire n_344;
wire n_503;
wire n_283;
wire n_756;
wire n_520;
wire n_681;
wire n_435;
wire n_577;
wire n_870;
wire n_790;
wire n_761;
wire n_615;
wire n_472;
wire n_419;
wire n_851;
wire n_825;
wire n_396;
wire n_804;
wire n_477;
wire n_815;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_721;
wire n_640;
wire n_908;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_821;
wire n_745;
wire n_684;
wire n_440;
wire n_553;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_723;
wire n_811;
wire n_749;
wire n_835;
wire n_535;
wire n_530;
wire n_737;
wire n_778;
wire n_358;
wire n_795;
wire n_267;
wire n_456;
wire n_782;
wire n_449;
wire n_300;
wire n_734;
wire n_524;
wire n_584;
wire n_919;
wire n_763;
wire n_497;
wire n_728;
wire n_339;
wire n_657;
wire n_583;
wire n_875;
wire n_620;
wire n_240;
wire n_841;
wire n_912;
wire n_924;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_441;
wire n_836;
wire n_923;
wire n_561;
wire n_335;
wire n_272;
wire n_741;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_397;
wire n_306;
wire n_242;
wire n_766;
wire n_602;
wire n_831;
wire n_859;
wire n_424;
wire n_714;
wire n_629;
wire n_569;
wire n_297;
wire n_837;
wire n_410;
wire n_774;
wire n_867;
wire n_377;
wire n_510;
wire n_343;
wire n_675;
wire n_291;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_855;
wire n_722;
wire n_618;
wire n_834;
wire n_901;
wire n_727;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_785;
wire n_375;
wire n_451;
wire n_487;
wire n_748;
wire n_371;
wire n_688;
wire n_868;
wire n_323;
wire n_473;
wire n_347;
wire n_820;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_843;
wire n_266;
wire n_683;
wire n_824;
wire n_538;
wire n_793;
wire n_492;
wire n_592;
wire n_753;
wire n_368;
wire n_355;
wire n_382;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_521;
wire n_695;
wire n_625;
wire n_650;
wire n_469;
wire n_742;
wire n_585;
wire n_913;
wire n_845;
wire n_713;
wire n_891;
wire n_457;
wire n_595;
wire n_759;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_833;
wire n_866;
wire n_736;
wire n_287;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_781;
wire n_916;
wire n_421;
wire n_709;
wire n_739;
wire n_740;
wire n_483;
wire n_408;
wire n_772;
wire n_290;
wire n_405;
wire n_819;
wire n_280;
wire n_395;
wire n_406;
wire n_491;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g228 ( .A(n_151), .Y(n_228) );
CKINVDCx20_ASAP7_75t_R g229 ( .A(n_224), .Y(n_229) );
INVx2_ASAP7_75t_L g230 ( .A(n_38), .Y(n_230) );
INVx1_ASAP7_75t_L g231 ( .A(n_225), .Y(n_231) );
CKINVDCx20_ASAP7_75t_R g232 ( .A(n_134), .Y(n_232) );
INVxp67_ASAP7_75t_L g233 ( .A(n_108), .Y(n_233) );
INVxp67_ASAP7_75t_SL g234 ( .A(n_43), .Y(n_234) );
INVx1_ASAP7_75t_L g235 ( .A(n_53), .Y(n_235) );
INVx1_ASAP7_75t_L g236 ( .A(n_179), .Y(n_236) );
OR2x2_ASAP7_75t_L g237 ( .A(n_101), .B(n_85), .Y(n_237) );
CKINVDCx5p33_ASAP7_75t_R g238 ( .A(n_199), .Y(n_238) );
CKINVDCx5p33_ASAP7_75t_R g239 ( .A(n_128), .Y(n_239) );
INVx1_ASAP7_75t_L g240 ( .A(n_89), .Y(n_240) );
CKINVDCx5p33_ASAP7_75t_R g241 ( .A(n_192), .Y(n_241) );
INVx1_ASAP7_75t_L g242 ( .A(n_215), .Y(n_242) );
BUFx2_ASAP7_75t_L g243 ( .A(n_95), .Y(n_243) );
INVx1_ASAP7_75t_L g244 ( .A(n_68), .Y(n_244) );
INVx1_ASAP7_75t_L g245 ( .A(n_94), .Y(n_245) );
CKINVDCx5p33_ASAP7_75t_R g246 ( .A(n_218), .Y(n_246) );
INVx1_ASAP7_75t_L g247 ( .A(n_137), .Y(n_247) );
INVx1_ASAP7_75t_L g248 ( .A(n_129), .Y(n_248) );
CKINVDCx20_ASAP7_75t_R g249 ( .A(n_83), .Y(n_249) );
INVx1_ASAP7_75t_L g250 ( .A(n_23), .Y(n_250) );
CKINVDCx16_ASAP7_75t_R g251 ( .A(n_213), .Y(n_251) );
INVxp33_ASAP7_75t_L g252 ( .A(n_135), .Y(n_252) );
CKINVDCx5p33_ASAP7_75t_R g253 ( .A(n_161), .Y(n_253) );
INVx1_ASAP7_75t_L g254 ( .A(n_184), .Y(n_254) );
INVx1_ASAP7_75t_L g255 ( .A(n_159), .Y(n_255) );
NOR2xp67_ASAP7_75t_L g256 ( .A(n_66), .B(n_73), .Y(n_256) );
INVx1_ASAP7_75t_L g257 ( .A(n_12), .Y(n_257) );
INVx1_ASAP7_75t_L g258 ( .A(n_118), .Y(n_258) );
CKINVDCx16_ASAP7_75t_R g259 ( .A(n_181), .Y(n_259) );
BUFx2_ASAP7_75t_L g260 ( .A(n_91), .Y(n_260) );
INVx1_ASAP7_75t_L g261 ( .A(n_205), .Y(n_261) );
INVx2_ASAP7_75t_L g262 ( .A(n_73), .Y(n_262) );
INVx1_ASAP7_75t_L g263 ( .A(n_87), .Y(n_263) );
INVx1_ASAP7_75t_L g264 ( .A(n_126), .Y(n_264) );
INVx1_ASAP7_75t_L g265 ( .A(n_142), .Y(n_265) );
INVx2_ASAP7_75t_L g266 ( .A(n_119), .Y(n_266) );
CKINVDCx20_ASAP7_75t_R g267 ( .A(n_19), .Y(n_267) );
INVx1_ASAP7_75t_L g268 ( .A(n_34), .Y(n_268) );
INVx1_ASAP7_75t_L g269 ( .A(n_33), .Y(n_269) );
INVx2_ASAP7_75t_L g270 ( .A(n_227), .Y(n_270) );
XNOR2xp5_ASAP7_75t_L g271 ( .A(n_203), .B(n_147), .Y(n_271) );
INVx1_ASAP7_75t_L g272 ( .A(n_1), .Y(n_272) );
CKINVDCx5p33_ASAP7_75t_R g273 ( .A(n_24), .Y(n_273) );
CKINVDCx5p33_ASAP7_75t_R g274 ( .A(n_115), .Y(n_274) );
INVx1_ASAP7_75t_L g275 ( .A(n_138), .Y(n_275) );
INVx1_ASAP7_75t_L g276 ( .A(n_197), .Y(n_276) );
CKINVDCx5p33_ASAP7_75t_R g277 ( .A(n_169), .Y(n_277) );
INVxp67_ASAP7_75t_SL g278 ( .A(n_198), .Y(n_278) );
INVx1_ASAP7_75t_L g279 ( .A(n_32), .Y(n_279) );
INVxp67_ASAP7_75t_L g280 ( .A(n_110), .Y(n_280) );
INVx1_ASAP7_75t_L g281 ( .A(n_23), .Y(n_281) );
CKINVDCx5p33_ASAP7_75t_R g282 ( .A(n_36), .Y(n_282) );
INVxp33_ASAP7_75t_L g283 ( .A(n_154), .Y(n_283) );
INVx1_ASAP7_75t_L g284 ( .A(n_28), .Y(n_284) );
CKINVDCx14_ASAP7_75t_R g285 ( .A(n_168), .Y(n_285) );
INVx1_ASAP7_75t_L g286 ( .A(n_70), .Y(n_286) );
INVx1_ASAP7_75t_L g287 ( .A(n_155), .Y(n_287) );
INVx2_ASAP7_75t_L g288 ( .A(n_208), .Y(n_288) );
INVx1_ASAP7_75t_L g289 ( .A(n_219), .Y(n_289) );
CKINVDCx20_ASAP7_75t_R g290 ( .A(n_1), .Y(n_290) );
INVx1_ASAP7_75t_L g291 ( .A(n_171), .Y(n_291) );
INVx1_ASAP7_75t_L g292 ( .A(n_93), .Y(n_292) );
BUFx3_ASAP7_75t_L g293 ( .A(n_25), .Y(n_293) );
NOR2xp67_ASAP7_75t_L g294 ( .A(n_123), .B(n_188), .Y(n_294) );
INVx2_ASAP7_75t_L g295 ( .A(n_121), .Y(n_295) );
INVx1_ASAP7_75t_L g296 ( .A(n_79), .Y(n_296) );
INVx1_ASAP7_75t_L g297 ( .A(n_114), .Y(n_297) );
INVx1_ASAP7_75t_L g298 ( .A(n_56), .Y(n_298) );
CKINVDCx20_ASAP7_75t_R g299 ( .A(n_28), .Y(n_299) );
OR2x2_ASAP7_75t_L g300 ( .A(n_88), .B(n_125), .Y(n_300) );
INVx1_ASAP7_75t_L g301 ( .A(n_141), .Y(n_301) );
INVx1_ASAP7_75t_L g302 ( .A(n_36), .Y(n_302) );
INVx1_ASAP7_75t_L g303 ( .A(n_212), .Y(n_303) );
INVx1_ASAP7_75t_L g304 ( .A(n_66), .Y(n_304) );
INVxp33_ASAP7_75t_L g305 ( .A(n_209), .Y(n_305) );
INVx1_ASAP7_75t_L g306 ( .A(n_74), .Y(n_306) );
CKINVDCx5p33_ASAP7_75t_R g307 ( .A(n_193), .Y(n_307) );
INVx1_ASAP7_75t_L g308 ( .A(n_70), .Y(n_308) );
CKINVDCx5p33_ASAP7_75t_R g309 ( .A(n_116), .Y(n_309) );
INVx1_ASAP7_75t_L g310 ( .A(n_194), .Y(n_310) );
CKINVDCx20_ASAP7_75t_R g311 ( .A(n_15), .Y(n_311) );
INVx2_ASAP7_75t_L g312 ( .A(n_157), .Y(n_312) );
BUFx6f_ASAP7_75t_L g313 ( .A(n_24), .Y(n_313) );
INVx1_ASAP7_75t_L g314 ( .A(n_136), .Y(n_314) );
BUFx5_ASAP7_75t_L g315 ( .A(n_201), .Y(n_315) );
CKINVDCx16_ASAP7_75t_R g316 ( .A(n_148), .Y(n_316) );
INVx2_ASAP7_75t_L g317 ( .A(n_86), .Y(n_317) );
INVx4_ASAP7_75t_R g318 ( .A(n_19), .Y(n_318) );
CKINVDCx5p33_ASAP7_75t_R g319 ( .A(n_56), .Y(n_319) );
INVx1_ASAP7_75t_L g320 ( .A(n_124), .Y(n_320) );
INVx1_ASAP7_75t_L g321 ( .A(n_180), .Y(n_321) );
INVx1_ASAP7_75t_L g322 ( .A(n_178), .Y(n_322) );
INVx1_ASAP7_75t_L g323 ( .A(n_189), .Y(n_323) );
INVx1_ASAP7_75t_L g324 ( .A(n_117), .Y(n_324) );
INVx1_ASAP7_75t_L g325 ( .A(n_52), .Y(n_325) );
INVx1_ASAP7_75t_L g326 ( .A(n_206), .Y(n_326) );
INVx1_ASAP7_75t_L g327 ( .A(n_211), .Y(n_327) );
CKINVDCx20_ASAP7_75t_R g328 ( .A(n_202), .Y(n_328) );
INVx1_ASAP7_75t_L g329 ( .A(n_47), .Y(n_329) );
INVx1_ASAP7_75t_L g330 ( .A(n_40), .Y(n_330) );
INVx1_ASAP7_75t_SL g331 ( .A(n_150), .Y(n_331) );
BUFx2_ASAP7_75t_SL g332 ( .A(n_216), .Y(n_332) );
INVx1_ASAP7_75t_L g333 ( .A(n_158), .Y(n_333) );
INVx1_ASAP7_75t_L g334 ( .A(n_11), .Y(n_334) );
CKINVDCx16_ASAP7_75t_R g335 ( .A(n_21), .Y(n_335) );
INVxp67_ASAP7_75t_L g336 ( .A(n_153), .Y(n_336) );
OR2x2_ASAP7_75t_L g337 ( .A(n_44), .B(n_45), .Y(n_337) );
CKINVDCx5p33_ASAP7_75t_R g338 ( .A(n_96), .Y(n_338) );
CKINVDCx5p33_ASAP7_75t_R g339 ( .A(n_65), .Y(n_339) );
CKINVDCx5p33_ASAP7_75t_R g340 ( .A(n_71), .Y(n_340) );
INVx1_ASAP7_75t_L g341 ( .A(n_195), .Y(n_341) );
INVx1_ASAP7_75t_L g342 ( .A(n_46), .Y(n_342) );
BUFx2_ASAP7_75t_L g343 ( .A(n_223), .Y(n_343) );
HB1xp67_ASAP7_75t_L g344 ( .A(n_120), .Y(n_344) );
INVx1_ASAP7_75t_L g345 ( .A(n_204), .Y(n_345) );
NOR2xp67_ASAP7_75t_L g346 ( .A(n_210), .B(n_222), .Y(n_346) );
INVx2_ASAP7_75t_L g347 ( .A(n_30), .Y(n_347) );
INVx3_ASAP7_75t_L g348 ( .A(n_13), .Y(n_348) );
INVx1_ASAP7_75t_L g349 ( .A(n_90), .Y(n_349) );
CKINVDCx5p33_ASAP7_75t_R g350 ( .A(n_92), .Y(n_350) );
INVx1_ASAP7_75t_L g351 ( .A(n_146), .Y(n_351) );
INVx1_ASAP7_75t_L g352 ( .A(n_54), .Y(n_352) );
CKINVDCx14_ASAP7_75t_R g353 ( .A(n_68), .Y(n_353) );
INVx1_ASAP7_75t_L g354 ( .A(n_47), .Y(n_354) );
INVx1_ASAP7_75t_L g355 ( .A(n_133), .Y(n_355) );
CKINVDCx5p33_ASAP7_75t_R g356 ( .A(n_112), .Y(n_356) );
INVx1_ASAP7_75t_L g357 ( .A(n_106), .Y(n_357) );
HB1xp67_ASAP7_75t_L g358 ( .A(n_72), .Y(n_358) );
INVx1_ASAP7_75t_L g359 ( .A(n_172), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_200), .Y(n_360) );
INVx1_ASAP7_75t_L g361 ( .A(n_45), .Y(n_361) );
BUFx2_ASAP7_75t_L g362 ( .A(n_139), .Y(n_362) );
INVx1_ASAP7_75t_L g363 ( .A(n_53), .Y(n_363) );
INVx1_ASAP7_75t_L g364 ( .A(n_107), .Y(n_364) );
BUFx3_ASAP7_75t_L g365 ( .A(n_84), .Y(n_365) );
NOR2xp33_ASAP7_75t_L g366 ( .A(n_252), .B(n_0), .Y(n_366) );
AND2x6_ASAP7_75t_L g367 ( .A(n_365), .B(n_80), .Y(n_367) );
INVx3_ASAP7_75t_L g368 ( .A(n_348), .Y(n_368) );
INVx2_ASAP7_75t_L g369 ( .A(n_315), .Y(n_369) );
NOR2xp33_ASAP7_75t_L g370 ( .A(n_252), .B(n_283), .Y(n_370) );
CKINVDCx5p33_ASAP7_75t_R g371 ( .A(n_251), .Y(n_371) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_243), .B(n_0), .Y(n_372) );
AOI22xp5_ASAP7_75t_SL g373 ( .A1(n_267), .A2(n_2), .B1(n_3), .B2(n_4), .Y(n_373) );
INVx2_ASAP7_75t_L g374 ( .A(n_315), .Y(n_374) );
INVx1_ASAP7_75t_L g375 ( .A(n_348), .Y(n_375) );
AND2x4_ASAP7_75t_L g376 ( .A(n_348), .B(n_2), .Y(n_376) );
BUFx12f_ASAP7_75t_L g377 ( .A(n_238), .Y(n_377) );
AND2x2_ASAP7_75t_L g378 ( .A(n_283), .B(n_3), .Y(n_378) );
OAI22xp5_ASAP7_75t_SL g379 ( .A1(n_267), .A2(n_4), .B1(n_5), .B2(n_6), .Y(n_379) );
BUFx2_ASAP7_75t_L g380 ( .A(n_353), .Y(n_380) );
AOI22xp5_ASAP7_75t_L g381 ( .A1(n_353), .A2(n_5), .B1(n_6), .B2(n_7), .Y(n_381) );
INVx2_ASAP7_75t_L g382 ( .A(n_315), .Y(n_382) );
INVx2_ASAP7_75t_L g383 ( .A(n_315), .Y(n_383) );
INVx3_ASAP7_75t_L g384 ( .A(n_293), .Y(n_384) );
OAI22xp5_ASAP7_75t_SL g385 ( .A1(n_290), .A2(n_7), .B1(n_8), .B2(n_9), .Y(n_385) );
OAI22xp5_ASAP7_75t_SL g386 ( .A1(n_290), .A2(n_8), .B1(n_9), .B2(n_10), .Y(n_386) );
BUFx8_ASAP7_75t_L g387 ( .A(n_260), .Y(n_387) );
OAI21x1_ASAP7_75t_L g388 ( .A1(n_266), .A2(n_82), .B(n_81), .Y(n_388) );
INVx3_ASAP7_75t_L g389 ( .A(n_293), .Y(n_389) );
INVx4_ASAP7_75t_L g390 ( .A(n_313), .Y(n_390) );
INVx3_ASAP7_75t_L g391 ( .A(n_266), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_230), .Y(n_392) );
INVx2_ASAP7_75t_L g393 ( .A(n_315), .Y(n_393) );
INVx1_ASAP7_75t_L g394 ( .A(n_230), .Y(n_394) );
AOI22xp5_ASAP7_75t_L g395 ( .A1(n_335), .A2(n_10), .B1(n_11), .B2(n_12), .Y(n_395) );
INVx1_ASAP7_75t_L g396 ( .A(n_262), .Y(n_396) );
HB1xp67_ASAP7_75t_L g397 ( .A(n_358), .Y(n_397) );
INVx2_ASAP7_75t_L g398 ( .A(n_315), .Y(n_398) );
BUFx2_ASAP7_75t_L g399 ( .A(n_285), .Y(n_399) );
INVx1_ASAP7_75t_L g400 ( .A(n_262), .Y(n_400) );
INVx1_ASAP7_75t_L g401 ( .A(n_369), .Y(n_401) );
NAND2xp5_ASAP7_75t_L g402 ( .A(n_370), .B(n_343), .Y(n_402) );
INVx1_ASAP7_75t_L g403 ( .A(n_369), .Y(n_403) );
INVx1_ASAP7_75t_L g404 ( .A(n_369), .Y(n_404) );
NAND2xp5_ASAP7_75t_L g405 ( .A(n_370), .B(n_362), .Y(n_405) );
NAND2xp5_ASAP7_75t_SL g406 ( .A(n_399), .B(n_259), .Y(n_406) );
INVx1_ASAP7_75t_SL g407 ( .A(n_380), .Y(n_407) );
NAND2xp5_ASAP7_75t_SL g408 ( .A(n_399), .B(n_316), .Y(n_408) );
INVx1_ASAP7_75t_L g409 ( .A(n_374), .Y(n_409) );
INVx2_ASAP7_75t_L g410 ( .A(n_374), .Y(n_410) );
INVx2_ASAP7_75t_L g411 ( .A(n_374), .Y(n_411) );
NAND2xp5_ASAP7_75t_L g412 ( .A(n_368), .B(n_344), .Y(n_412) );
INVx3_ASAP7_75t_L g413 ( .A(n_376), .Y(n_413) );
AOI22xp5_ASAP7_75t_L g414 ( .A1(n_378), .A2(n_381), .B1(n_376), .B2(n_395), .Y(n_414) );
INVx1_ASAP7_75t_L g415 ( .A(n_382), .Y(n_415) );
AND2x2_ASAP7_75t_L g416 ( .A(n_397), .B(n_305), .Y(n_416) );
NOR2xp33_ASAP7_75t_L g417 ( .A(n_371), .B(n_233), .Y(n_417) );
CKINVDCx20_ASAP7_75t_R g418 ( .A(n_387), .Y(n_418) );
AND2x2_ASAP7_75t_L g419 ( .A(n_397), .B(n_285), .Y(n_419) );
BUFx6f_ASAP7_75t_L g420 ( .A(n_388), .Y(n_420) );
NOR3xp33_ASAP7_75t_L g421 ( .A(n_379), .B(n_234), .C(n_273), .Y(n_421) );
INVx4_ASAP7_75t_L g422 ( .A(n_376), .Y(n_422) );
INVx1_ASAP7_75t_L g423 ( .A(n_382), .Y(n_423) );
NOR2xp33_ASAP7_75t_L g424 ( .A(n_377), .B(n_280), .Y(n_424) );
OR2x2_ASAP7_75t_L g425 ( .A(n_372), .B(n_273), .Y(n_425) );
INVx2_ASAP7_75t_L g426 ( .A(n_382), .Y(n_426) );
NAND2xp5_ASAP7_75t_L g427 ( .A(n_378), .B(n_282), .Y(n_427) );
NAND2xp5_ASAP7_75t_SL g428 ( .A(n_387), .B(n_238), .Y(n_428) );
NAND3x1_ASAP7_75t_L g429 ( .A(n_381), .B(n_244), .C(n_235), .Y(n_429) );
BUFx3_ASAP7_75t_L g430 ( .A(n_376), .Y(n_430) );
OR2x2_ASAP7_75t_L g431 ( .A(n_372), .B(n_282), .Y(n_431) );
AND2x2_ASAP7_75t_L g432 ( .A(n_378), .B(n_347), .Y(n_432) );
BUFx6f_ASAP7_75t_L g433 ( .A(n_388), .Y(n_433) );
NAND2xp5_ASAP7_75t_L g434 ( .A(n_368), .B(n_270), .Y(n_434) );
INVx1_ASAP7_75t_L g435 ( .A(n_383), .Y(n_435) );
NAND2xp5_ASAP7_75t_L g436 ( .A(n_368), .B(n_319), .Y(n_436) );
NOR2xp33_ASAP7_75t_L g437 ( .A(n_377), .B(n_336), .Y(n_437) );
NAND2xp5_ASAP7_75t_SL g438 ( .A(n_387), .B(n_239), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_383), .Y(n_439) );
INVx4_ASAP7_75t_L g440 ( .A(n_376), .Y(n_440) );
INVx2_ASAP7_75t_SL g441 ( .A(n_368), .Y(n_441) );
INVx2_ASAP7_75t_L g442 ( .A(n_383), .Y(n_442) );
INVx2_ASAP7_75t_L g443 ( .A(n_393), .Y(n_443) );
BUFx10_ASAP7_75t_L g444 ( .A(n_367), .Y(n_444) );
NAND2xp5_ASAP7_75t_L g445 ( .A(n_412), .B(n_387), .Y(n_445) );
NAND2xp5_ASAP7_75t_SL g446 ( .A(n_422), .B(n_387), .Y(n_446) );
AOI22xp5_ASAP7_75t_L g447 ( .A1(n_414), .A2(n_377), .B1(n_366), .B2(n_395), .Y(n_447) );
NAND2xp5_ASAP7_75t_L g448 ( .A(n_412), .B(n_366), .Y(n_448) );
OAI22xp5_ASAP7_75t_SL g449 ( .A1(n_418), .A2(n_385), .B1(n_386), .B2(n_379), .Y(n_449) );
NAND2xp5_ASAP7_75t_SL g450 ( .A(n_422), .B(n_393), .Y(n_450) );
INVx2_ASAP7_75t_SL g451 ( .A(n_407), .Y(n_451) );
OAI22xp5_ASAP7_75t_L g452 ( .A1(n_414), .A2(n_232), .B1(n_249), .B2(n_229), .Y(n_452) );
INVx3_ASAP7_75t_L g453 ( .A(n_422), .Y(n_453) );
NAND2xp5_ASAP7_75t_L g454 ( .A(n_432), .B(n_375), .Y(n_454) );
HB1xp67_ASAP7_75t_L g455 ( .A(n_407), .Y(n_455) );
NAND2xp5_ASAP7_75t_L g456 ( .A(n_432), .B(n_384), .Y(n_456) );
NAND2xp5_ASAP7_75t_SL g457 ( .A(n_440), .B(n_393), .Y(n_457) );
AOI22xp33_ASAP7_75t_SL g458 ( .A1(n_419), .A2(n_373), .B1(n_386), .B2(n_385), .Y(n_458) );
AOI22xp33_ASAP7_75t_L g459 ( .A1(n_430), .A2(n_391), .B1(n_367), .B2(n_398), .Y(n_459) );
AOI22xp5_ASAP7_75t_L g460 ( .A1(n_419), .A2(n_232), .B1(n_249), .B2(n_229), .Y(n_460) );
NOR2xp33_ASAP7_75t_L g461 ( .A(n_402), .B(n_392), .Y(n_461) );
OAI21xp5_ASAP7_75t_L g462 ( .A1(n_401), .A2(n_388), .B(n_398), .Y(n_462) );
NAND2xp5_ASAP7_75t_SL g463 ( .A(n_440), .B(n_239), .Y(n_463) );
INVx1_ASAP7_75t_L g464 ( .A(n_441), .Y(n_464) );
NOR2x1p5_ASAP7_75t_L g465 ( .A(n_416), .B(n_339), .Y(n_465) );
BUFx6f_ASAP7_75t_L g466 ( .A(n_444), .Y(n_466) );
NAND2xp5_ASAP7_75t_L g467 ( .A(n_405), .B(n_384), .Y(n_467) );
BUFx3_ASAP7_75t_L g468 ( .A(n_416), .Y(n_468) );
INVx1_ASAP7_75t_L g469 ( .A(n_441), .Y(n_469) );
NAND2xp5_ASAP7_75t_SL g470 ( .A(n_440), .B(n_398), .Y(n_470) );
NAND2xp5_ASAP7_75t_SL g471 ( .A(n_440), .B(n_228), .Y(n_471) );
NAND2xp5_ASAP7_75t_SL g472 ( .A(n_427), .B(n_241), .Y(n_472) );
AND2x6_ASAP7_75t_L g473 ( .A(n_413), .B(n_384), .Y(n_473) );
INVx1_ASAP7_75t_L g474 ( .A(n_434), .Y(n_474) );
O2A1O1Ixp5_ASAP7_75t_L g475 ( .A1(n_436), .A2(n_389), .B(n_278), .C(n_231), .Y(n_475) );
AOI22xp5_ASAP7_75t_L g476 ( .A1(n_425), .A2(n_328), .B1(n_339), .B2(n_340), .Y(n_476) );
INVx2_ASAP7_75t_SL g477 ( .A(n_425), .Y(n_477) );
NAND2xp5_ASAP7_75t_SL g478 ( .A(n_431), .B(n_246), .Y(n_478) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_431), .B(n_389), .Y(n_479) );
NAND2xp5_ASAP7_75t_L g480 ( .A(n_413), .B(n_389), .Y(n_480) );
NAND2xp5_ASAP7_75t_L g481 ( .A(n_406), .B(n_389), .Y(n_481) );
NAND2xp5_ASAP7_75t_L g482 ( .A(n_408), .B(n_246), .Y(n_482) );
INVx2_ASAP7_75t_SL g483 ( .A(n_428), .Y(n_483) );
NOR2xp33_ASAP7_75t_L g484 ( .A(n_424), .B(n_392), .Y(n_484) );
AOI22xp33_ASAP7_75t_L g485 ( .A1(n_420), .A2(n_391), .B1(n_367), .B2(n_394), .Y(n_485) );
AOI22xp5_ASAP7_75t_L g486 ( .A1(n_438), .A2(n_257), .B1(n_268), .B2(n_250), .Y(n_486) );
NAND3xp33_ASAP7_75t_SL g487 ( .A(n_421), .B(n_311), .C(n_299), .Y(n_487) );
AND2x6_ASAP7_75t_SL g488 ( .A(n_417), .B(n_373), .Y(n_488) );
AOI22xp33_ASAP7_75t_L g489 ( .A1(n_420), .A2(n_391), .B1(n_367), .B2(n_394), .Y(n_489) );
A2O1A1Ixp33_ASAP7_75t_L g490 ( .A1(n_401), .A2(n_391), .B(n_400), .C(n_396), .Y(n_490) );
INVx2_ASAP7_75t_L g491 ( .A(n_410), .Y(n_491) );
INVx2_ASAP7_75t_L g492 ( .A(n_410), .Y(n_492) );
BUFx3_ASAP7_75t_L g493 ( .A(n_403), .Y(n_493) );
AOI22xp5_ASAP7_75t_L g494 ( .A1(n_429), .A2(n_269), .B1(n_279), .B2(n_272), .Y(n_494) );
NAND3xp33_ASAP7_75t_L g495 ( .A(n_437), .B(n_274), .C(n_253), .Y(n_495) );
INVxp67_ASAP7_75t_SL g496 ( .A(n_404), .Y(n_496) );
OR2x6_ASAP7_75t_L g497 ( .A(n_429), .B(n_337), .Y(n_497) );
INVx2_ASAP7_75t_L g498 ( .A(n_410), .Y(n_498) );
NAND2xp5_ASAP7_75t_SL g499 ( .A(n_444), .B(n_236), .Y(n_499) );
NAND2xp5_ASAP7_75t_SL g500 ( .A(n_420), .B(n_240), .Y(n_500) );
NAND2xp5_ASAP7_75t_SL g501 ( .A(n_420), .B(n_242), .Y(n_501) );
AOI22xp5_ASAP7_75t_L g502 ( .A1(n_404), .A2(n_284), .B1(n_286), .B2(n_281), .Y(n_502) );
NOR2xp33_ASAP7_75t_L g503 ( .A(n_409), .B(n_396), .Y(n_503) );
OAI22xp5_ASAP7_75t_SL g504 ( .A1(n_420), .A2(n_311), .B1(n_299), .B2(n_271), .Y(n_504) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_409), .B(n_253), .Y(n_505) );
AND2x6_ASAP7_75t_SL g506 ( .A(n_415), .B(n_298), .Y(n_506) );
INVx2_ASAP7_75t_L g507 ( .A(n_411), .Y(n_507) );
OAI22xp5_ASAP7_75t_L g508 ( .A1(n_433), .A2(n_302), .B1(n_306), .B2(n_304), .Y(n_508) );
AOI22xp33_ASAP7_75t_L g509 ( .A1(n_433), .A2(n_391), .B1(n_367), .B2(n_400), .Y(n_509) );
INVx2_ASAP7_75t_L g510 ( .A(n_426), .Y(n_510) );
AND2x4_ASAP7_75t_L g511 ( .A(n_433), .B(n_256), .Y(n_511) );
NAND2xp5_ASAP7_75t_SL g512 ( .A(n_433), .B(n_245), .Y(n_512) );
NAND2xp5_ASAP7_75t_SL g513 ( .A(n_433), .B(n_247), .Y(n_513) );
INVx2_ASAP7_75t_SL g514 ( .A(n_415), .Y(n_514) );
AOI22xp5_ASAP7_75t_L g515 ( .A1(n_423), .A2(n_325), .B1(n_329), .B2(n_308), .Y(n_515) );
AOI22xp5_ASAP7_75t_L g516 ( .A1(n_435), .A2(n_334), .B1(n_342), .B2(n_330), .Y(n_516) );
NAND2xp5_ASAP7_75t_SL g517 ( .A(n_451), .B(n_277), .Y(n_517) );
A2O1A1Ixp33_ASAP7_75t_L g518 ( .A1(n_461), .A2(n_439), .B(n_442), .C(n_426), .Y(n_518) );
AND2x6_ASAP7_75t_L g519 ( .A(n_474), .B(n_365), .Y(n_519) );
BUFx3_ASAP7_75t_L g520 ( .A(n_455), .Y(n_520) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_477), .B(n_443), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_445), .B(n_448), .Y(n_522) );
INVx6_ASAP7_75t_L g523 ( .A(n_506), .Y(n_523) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_461), .B(n_443), .Y(n_524) );
INVx1_ASAP7_75t_L g525 ( .A(n_454), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g526 ( .A(n_496), .B(n_352), .Y(n_526) );
BUFx6f_ASAP7_75t_L g527 ( .A(n_493), .Y(n_527) );
NOR2xp33_ASAP7_75t_L g528 ( .A(n_468), .B(n_354), .Y(n_528) );
AOI21xp5_ASAP7_75t_L g529 ( .A1(n_500), .A2(n_254), .B(n_248), .Y(n_529) );
OAI21xp5_ASAP7_75t_L g530 ( .A1(n_462), .A2(n_367), .B(n_258), .Y(n_530) );
NAND3xp33_ASAP7_75t_SL g531 ( .A(n_458), .B(n_309), .C(n_307), .Y(n_531) );
NOR2xp33_ASAP7_75t_L g532 ( .A(n_478), .B(n_361), .Y(n_532) );
BUFx6f_ASAP7_75t_L g533 ( .A(n_466), .Y(n_533) );
NAND2x1p5_ASAP7_75t_L g534 ( .A(n_446), .B(n_347), .Y(n_534) );
INVx1_ASAP7_75t_L g535 ( .A(n_479), .Y(n_535) );
NAND2xp33_ASAP7_75t_L g536 ( .A(n_473), .B(n_367), .Y(n_536) );
A2O1A1Ixp33_ASAP7_75t_L g537 ( .A1(n_484), .A2(n_363), .B(n_255), .C(n_263), .Y(n_537) );
AOI21xp5_ASAP7_75t_L g538 ( .A1(n_501), .A2(n_264), .B(n_261), .Y(n_538) );
AOI21xp5_ASAP7_75t_L g539 ( .A1(n_512), .A2(n_275), .B(n_265), .Y(n_539) );
INVx3_ASAP7_75t_L g540 ( .A(n_453), .Y(n_540) );
HB1xp67_ASAP7_75t_L g541 ( .A(n_452), .Y(n_541) );
O2A1O1Ixp33_ASAP7_75t_L g542 ( .A1(n_508), .A2(n_287), .B(n_289), .C(n_276), .Y(n_542) );
BUFx4f_ASAP7_75t_L g543 ( .A(n_497), .Y(n_543) );
AOI21xp5_ASAP7_75t_L g544 ( .A1(n_513), .A2(n_292), .B(n_291), .Y(n_544) );
AOI21x1_ASAP7_75t_L g545 ( .A1(n_513), .A2(n_346), .B(n_294), .Y(n_545) );
AND2x6_ASAP7_75t_L g546 ( .A(n_453), .B(n_296), .Y(n_546) );
INVx1_ASAP7_75t_SL g547 ( .A(n_514), .Y(n_547) );
INVx3_ASAP7_75t_L g548 ( .A(n_473), .Y(n_548) );
AOI21xp5_ASAP7_75t_L g549 ( .A1(n_450), .A2(n_301), .B(n_297), .Y(n_549) );
AO32x1_ASAP7_75t_L g550 ( .A1(n_483), .A2(n_390), .A3(n_326), .B1(n_364), .B2(n_360), .Y(n_550) );
A2O1A1Ixp33_ASAP7_75t_L g551 ( .A1(n_475), .A2(n_310), .B(n_314), .C(n_303), .Y(n_551) );
AOI21xp5_ASAP7_75t_L g552 ( .A1(n_450), .A2(n_321), .B(n_320), .Y(n_552) );
AOI21xp5_ASAP7_75t_L g553 ( .A1(n_457), .A2(n_323), .B(n_322), .Y(n_553) );
INVx3_ASAP7_75t_L g554 ( .A(n_473), .Y(n_554) );
INVx1_ASAP7_75t_L g555 ( .A(n_503), .Y(n_555) );
INVx3_ASAP7_75t_L g556 ( .A(n_473), .Y(n_556) );
NOR2xp33_ASAP7_75t_L g557 ( .A(n_482), .B(n_338), .Y(n_557) );
AOI21xp5_ASAP7_75t_L g558 ( .A1(n_457), .A2(n_327), .B(n_324), .Y(n_558) );
INVx4_ASAP7_75t_L g559 ( .A(n_473), .Y(n_559) );
INVx2_ASAP7_75t_SL g560 ( .A(n_465), .Y(n_560) );
A2O1A1Ixp33_ASAP7_75t_L g561 ( .A1(n_503), .A2(n_341), .B(n_345), .C(n_333), .Y(n_561) );
NOR2xp33_ASAP7_75t_L g562 ( .A(n_476), .B(n_338), .Y(n_562) );
CKINVDCx5p33_ASAP7_75t_R g563 ( .A(n_460), .Y(n_563) );
OAI22x1_ASAP7_75t_L g564 ( .A1(n_494), .A2(n_356), .B1(n_350), .B2(n_318), .Y(n_564) );
HB1xp67_ASAP7_75t_L g565 ( .A(n_504), .Y(n_565) );
OR2x2_ASAP7_75t_L g566 ( .A(n_497), .B(n_13), .Y(n_566) );
AOI21xp5_ASAP7_75t_L g567 ( .A1(n_470), .A2(n_351), .B(n_349), .Y(n_567) );
HB1xp67_ASAP7_75t_L g568 ( .A(n_497), .Y(n_568) );
AOI22xp5_ASAP7_75t_L g569 ( .A1(n_486), .A2(n_367), .B1(n_355), .B2(n_359), .Y(n_569) );
AOI21xp5_ASAP7_75t_L g570 ( .A1(n_471), .A2(n_357), .B(n_295), .Y(n_570) );
INVx1_ASAP7_75t_SL g571 ( .A(n_491), .Y(n_571) );
O2A1O1Ixp33_ASAP7_75t_L g572 ( .A1(n_467), .A2(n_317), .B(n_312), .C(n_288), .Y(n_572) );
NOR2xp33_ASAP7_75t_L g573 ( .A(n_472), .B(n_331), .Y(n_573) );
AOI21xp5_ASAP7_75t_L g574 ( .A1(n_471), .A2(n_317), .B(n_312), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g575 ( .A(n_492), .B(n_390), .Y(n_575) );
HB1xp67_ASAP7_75t_L g576 ( .A(n_505), .Y(n_576) );
AOI22xp33_ASAP7_75t_L g577 ( .A1(n_511), .A2(n_390), .B1(n_313), .B2(n_332), .Y(n_577) );
AOI22xp5_ASAP7_75t_L g578 ( .A1(n_487), .A2(n_313), .B1(n_390), .B2(n_315), .Y(n_578) );
AOI21xp5_ASAP7_75t_L g579 ( .A1(n_480), .A2(n_300), .B(n_237), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g580 ( .A(n_498), .B(n_390), .Y(n_580) );
AOI22xp5_ASAP7_75t_L g581 ( .A1(n_463), .A2(n_14), .B1(n_15), .B2(n_16), .Y(n_581) );
OAI22xp5_ASAP7_75t_L g582 ( .A1(n_490), .A2(n_14), .B1(n_16), .B2(n_17), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g583 ( .A(n_481), .B(n_17), .Y(n_583) );
OAI22xp33_ASAP7_75t_L g584 ( .A1(n_502), .A2(n_18), .B1(n_20), .B2(n_21), .Y(n_584) );
NOR2xp33_ASAP7_75t_L g585 ( .A(n_515), .B(n_18), .Y(n_585) );
BUFx3_ASAP7_75t_L g586 ( .A(n_511), .Y(n_586) );
AND2x2_ASAP7_75t_L g587 ( .A(n_516), .B(n_20), .Y(n_587) );
OAI22xp5_ASAP7_75t_SL g588 ( .A1(n_488), .A2(n_22), .B1(n_25), .B2(n_26), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g589 ( .A(n_507), .B(n_22), .Y(n_589) );
HB1xp67_ASAP7_75t_L g590 ( .A(n_510), .Y(n_590) );
NOR2xp33_ASAP7_75t_L g591 ( .A(n_464), .B(n_26), .Y(n_591) );
INVx2_ASAP7_75t_L g592 ( .A(n_469), .Y(n_592) );
BUFx2_ASAP7_75t_L g593 ( .A(n_466), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g594 ( .A(n_459), .B(n_27), .Y(n_594) );
NOR2xp33_ASAP7_75t_L g595 ( .A(n_499), .B(n_29), .Y(n_595) );
OAI22x1_ASAP7_75t_SL g596 ( .A1(n_485), .A2(n_31), .B1(n_32), .B2(n_33), .Y(n_596) );
AOI21xp5_ASAP7_75t_L g597 ( .A1(n_485), .A2(n_489), .B(n_509), .Y(n_597) );
AOI22xp33_ASAP7_75t_L g598 ( .A1(n_489), .A2(n_31), .B1(n_35), .B2(n_37), .Y(n_598) );
O2A1O1Ixp33_ASAP7_75t_SL g599 ( .A1(n_500), .A2(n_145), .B(n_221), .C(n_220), .Y(n_599) );
HB1xp67_ASAP7_75t_L g600 ( .A(n_455), .Y(n_600) );
HB1xp67_ASAP7_75t_L g601 ( .A(n_455), .Y(n_601) );
NOR2x1_ASAP7_75t_L g602 ( .A(n_495), .B(n_39), .Y(n_602) );
AND2x2_ASAP7_75t_L g603 ( .A(n_455), .B(n_39), .Y(n_603) );
AND2x2_ASAP7_75t_L g604 ( .A(n_455), .B(n_40), .Y(n_604) );
A2O1A1Ixp33_ASAP7_75t_L g605 ( .A1(n_461), .A2(n_41), .B(n_42), .C(n_43), .Y(n_605) );
AND2x2_ASAP7_75t_L g606 ( .A(n_455), .B(n_41), .Y(n_606) );
NAND2xp5_ASAP7_75t_SL g607 ( .A(n_451), .B(n_42), .Y(n_607) );
INVx3_ASAP7_75t_L g608 ( .A(n_493), .Y(n_608) );
AOI21xp5_ASAP7_75t_L g609 ( .A1(n_500), .A2(n_149), .B(n_217), .Y(n_609) );
INVx1_ASAP7_75t_L g610 ( .A(n_456), .Y(n_610) );
OAI22xp5_ASAP7_75t_L g611 ( .A1(n_522), .A2(n_48), .B1(n_49), .B2(n_50), .Y(n_611) );
BUFx10_ASAP7_75t_L g612 ( .A(n_600), .Y(n_612) );
BUFx12f_ASAP7_75t_L g613 ( .A(n_523), .Y(n_613) );
AO31x2_ASAP7_75t_L g614 ( .A1(n_551), .A2(n_48), .A3(n_49), .B(n_50), .Y(n_614) );
INVx1_ASAP7_75t_L g615 ( .A(n_521), .Y(n_615) );
AND2x2_ASAP7_75t_L g616 ( .A(n_601), .B(n_51), .Y(n_616) );
AND2x4_ASAP7_75t_L g617 ( .A(n_525), .B(n_51), .Y(n_617) );
AOI22xp33_ASAP7_75t_L g618 ( .A1(n_541), .A2(n_52), .B1(n_54), .B2(n_55), .Y(n_618) );
A2O1A1Ixp33_ASAP7_75t_L g619 ( .A1(n_522), .A2(n_55), .B(n_57), .C(n_58), .Y(n_619) );
O2A1O1Ixp33_ASAP7_75t_L g620 ( .A1(n_537), .A2(n_57), .B(n_58), .C(n_59), .Y(n_620) );
AOI21xp5_ASAP7_75t_L g621 ( .A1(n_530), .A2(n_152), .B(n_214), .Y(n_621) );
INVxp67_ASAP7_75t_SL g622 ( .A(n_547), .Y(n_622) );
AOI22xp33_ASAP7_75t_L g623 ( .A1(n_565), .A2(n_59), .B1(n_60), .B2(n_61), .Y(n_623) );
O2A1O1Ixp33_ASAP7_75t_L g624 ( .A1(n_561), .A2(n_60), .B(n_61), .C(n_62), .Y(n_624) );
INVx1_ASAP7_75t_SL g625 ( .A(n_603), .Y(n_625) );
AND2x2_ASAP7_75t_L g626 ( .A(n_543), .B(n_62), .Y(n_626) );
OAI21xp5_ASAP7_75t_L g627 ( .A1(n_530), .A2(n_156), .B(n_207), .Y(n_627) );
A2O1A1Ixp33_ASAP7_75t_L g628 ( .A1(n_579), .A2(n_63), .B(n_64), .C(n_65), .Y(n_628) );
BUFx8_ASAP7_75t_L g629 ( .A(n_566), .Y(n_629) );
A2O1A1Ixp33_ASAP7_75t_L g630 ( .A1(n_591), .A2(n_63), .B(n_64), .C(n_67), .Y(n_630) );
A2O1A1Ixp33_ASAP7_75t_L g631 ( .A1(n_555), .A2(n_67), .B(n_69), .C(n_71), .Y(n_631) );
A2O1A1Ixp33_ASAP7_75t_L g632 ( .A1(n_595), .A2(n_69), .B(n_72), .C(n_74), .Y(n_632) );
AND2x2_ASAP7_75t_L g633 ( .A(n_543), .B(n_75), .Y(n_633) );
AO31x2_ASAP7_75t_L g634 ( .A1(n_605), .A2(n_75), .A3(n_76), .B(n_77), .Y(n_634) );
AO31x2_ASAP7_75t_L g635 ( .A1(n_582), .A2(n_76), .A3(n_77), .B(n_78), .Y(n_635) );
AOI22xp5_ASAP7_75t_L g636 ( .A1(n_563), .A2(n_78), .B1(n_97), .B2(n_98), .Y(n_636) );
AOI21xp5_ASAP7_75t_L g637 ( .A1(n_575), .A2(n_99), .B(n_100), .Y(n_637) );
INVx3_ASAP7_75t_L g638 ( .A(n_527), .Y(n_638) );
INVx4_ASAP7_75t_L g639 ( .A(n_559), .Y(n_639) );
O2A1O1Ixp33_ASAP7_75t_L g640 ( .A1(n_584), .A2(n_102), .B(n_103), .C(n_104), .Y(n_640) );
OR2x2_ASAP7_75t_L g641 ( .A(n_568), .B(n_105), .Y(n_641) );
A2O1A1Ixp33_ASAP7_75t_L g642 ( .A1(n_535), .A2(n_109), .B(n_111), .C(n_113), .Y(n_642) );
NOR2xp33_ASAP7_75t_L g643 ( .A(n_562), .B(n_122), .Y(n_643) );
NOR2xp33_ASAP7_75t_SL g644 ( .A(n_559), .B(n_127), .Y(n_644) );
AOI22xp5_ASAP7_75t_L g645 ( .A1(n_531), .A2(n_130), .B1(n_131), .B2(n_132), .Y(n_645) );
INVx2_ASAP7_75t_SL g646 ( .A(n_604), .Y(n_646) );
O2A1O1Ixp33_ASAP7_75t_L g647 ( .A1(n_542), .A2(n_140), .B(n_143), .C(n_144), .Y(n_647) );
BUFx2_ASAP7_75t_L g648 ( .A(n_546), .Y(n_648) );
INVx2_ASAP7_75t_L g649 ( .A(n_592), .Y(n_649) );
O2A1O1Ixp33_ASAP7_75t_L g650 ( .A1(n_585), .A2(n_160), .B(n_162), .C(n_163), .Y(n_650) );
AO31x2_ASAP7_75t_L g651 ( .A1(n_582), .A2(n_164), .A3(n_165), .B(n_166), .Y(n_651) );
AOI21xp5_ASAP7_75t_L g652 ( .A1(n_580), .A2(n_167), .B(n_170), .Y(n_652) );
INVx1_ASAP7_75t_L g653 ( .A(n_606), .Y(n_653) );
AOI21xp5_ASAP7_75t_L g654 ( .A1(n_580), .A2(n_173), .B(n_174), .Y(n_654) );
NOR2xp33_ASAP7_75t_L g655 ( .A(n_560), .B(n_175), .Y(n_655) );
AO31x2_ASAP7_75t_L g656 ( .A1(n_589), .A2(n_176), .A3(n_177), .B(n_182), .Y(n_656) );
AO31x2_ASAP7_75t_L g657 ( .A1(n_589), .A2(n_183), .A3(n_185), .B(n_186), .Y(n_657) );
A2O1A1Ixp33_ASAP7_75t_L g658 ( .A1(n_572), .A2(n_187), .B(n_190), .C(n_191), .Y(n_658) );
AO21x1_ASAP7_75t_L g659 ( .A1(n_534), .A2(n_545), .B(n_536), .Y(n_659) );
NOR2xp33_ASAP7_75t_L g660 ( .A(n_576), .B(n_196), .Y(n_660) );
OR2x6_ASAP7_75t_L g661 ( .A(n_588), .B(n_226), .Y(n_661) );
CKINVDCx12_ASAP7_75t_R g662 ( .A(n_587), .Y(n_662) );
AO31x2_ASAP7_75t_L g663 ( .A1(n_594), .A2(n_574), .A3(n_570), .B(n_609), .Y(n_663) );
O2A1O1Ixp33_ASAP7_75t_SL g664 ( .A1(n_571), .A2(n_594), .B(n_583), .C(n_607), .Y(n_664) );
INVx1_ASAP7_75t_L g665 ( .A(n_526), .Y(n_665) );
BUFx3_ASAP7_75t_L g666 ( .A(n_608), .Y(n_666) );
CKINVDCx5p33_ASAP7_75t_R g667 ( .A(n_564), .Y(n_667) );
NOR2xp33_ASAP7_75t_L g668 ( .A(n_532), .B(n_517), .Y(n_668) );
AND2x4_ASAP7_75t_L g669 ( .A(n_610), .B(n_548), .Y(n_669) );
BUFx6f_ASAP7_75t_L g670 ( .A(n_533), .Y(n_670) );
BUFx8_ASAP7_75t_SL g671 ( .A(n_586), .Y(n_671) );
INVx4_ASAP7_75t_L g672 ( .A(n_546), .Y(n_672) );
OAI221xp5_ASAP7_75t_L g673 ( .A1(n_578), .A2(n_528), .B1(n_557), .B2(n_573), .C(n_581), .Y(n_673) );
AND2x4_ASAP7_75t_L g674 ( .A(n_548), .B(n_554), .Y(n_674) );
INVx3_ASAP7_75t_L g675 ( .A(n_546), .Y(n_675) );
INVx2_ASAP7_75t_SL g676 ( .A(n_546), .Y(n_676) );
AND2x4_ASAP7_75t_L g677 ( .A(n_554), .B(n_556), .Y(n_677) );
INVx1_ASAP7_75t_L g678 ( .A(n_590), .Y(n_678) );
INVx1_ASAP7_75t_SL g679 ( .A(n_519), .Y(n_679) );
BUFx12f_ASAP7_75t_L g680 ( .A(n_593), .Y(n_680) );
OAI22xp5_ASAP7_75t_L g681 ( .A1(n_556), .A2(n_598), .B1(n_569), .B2(n_577), .Y(n_681) );
INVx5_ASAP7_75t_L g682 ( .A(n_533), .Y(n_682) );
OAI21x1_ASAP7_75t_L g683 ( .A1(n_529), .A2(n_544), .B(n_538), .Y(n_683) );
INVx2_ASAP7_75t_SL g684 ( .A(n_602), .Y(n_684) );
AO31x2_ASAP7_75t_L g685 ( .A1(n_539), .A2(n_553), .A3(n_567), .B(n_549), .Y(n_685) );
OAI21xp5_ASAP7_75t_L g686 ( .A1(n_552), .A2(n_558), .B(n_540), .Y(n_686) );
INVx1_ASAP7_75t_L g687 ( .A(n_596), .Y(n_687) );
AOI22xp33_ASAP7_75t_L g688 ( .A1(n_550), .A2(n_541), .B1(n_449), .B2(n_565), .Y(n_688) );
OAI21xp5_ASAP7_75t_L g689 ( .A1(n_599), .A2(n_522), .B(n_518), .Y(n_689) );
AO31x2_ASAP7_75t_L g690 ( .A1(n_550), .A2(n_518), .A3(n_551), .B(n_597), .Y(n_690) );
O2A1O1Ixp33_ASAP7_75t_L g691 ( .A1(n_550), .A2(n_522), .B(n_537), .C(n_561), .Y(n_691) );
OAI222xp33_ASAP7_75t_L g692 ( .A1(n_541), .A2(n_452), .B1(n_458), .B2(n_373), .C1(n_381), .C2(n_460), .Y(n_692) );
A2O1A1Ixp33_ASAP7_75t_L g693 ( .A1(n_522), .A2(n_461), .B(n_579), .C(n_484), .Y(n_693) );
NOR2xp33_ASAP7_75t_SL g694 ( .A(n_543), .B(n_452), .Y(n_694) );
AO22x2_ASAP7_75t_L g695 ( .A1(n_566), .A2(n_452), .B1(n_451), .B2(n_531), .Y(n_695) );
INVx1_ASAP7_75t_L g696 ( .A(n_521), .Y(n_696) );
AOI22xp5_ASAP7_75t_L g697 ( .A1(n_547), .A2(n_452), .B1(n_451), .B2(n_455), .Y(n_697) );
AO31x2_ASAP7_75t_L g698 ( .A1(n_518), .A2(n_551), .A3(n_597), .B(n_561), .Y(n_698) );
OAI22xp5_ASAP7_75t_L g699 ( .A1(n_522), .A2(n_547), .B1(n_524), .B2(n_525), .Y(n_699) );
CKINVDCx20_ASAP7_75t_R g700 ( .A(n_520), .Y(n_700) );
A2O1A1Ixp33_ASAP7_75t_L g701 ( .A1(n_522), .A2(n_461), .B(n_579), .C(n_484), .Y(n_701) );
AO31x2_ASAP7_75t_L g702 ( .A1(n_518), .A2(n_551), .A3(n_597), .B(n_561), .Y(n_702) );
INVx1_ASAP7_75t_L g703 ( .A(n_521), .Y(n_703) );
AND2x2_ASAP7_75t_L g704 ( .A(n_600), .B(n_455), .Y(n_704) );
NAND2xp5_ASAP7_75t_L g705 ( .A(n_525), .B(n_477), .Y(n_705) );
NOR2xp33_ASAP7_75t_L g706 ( .A(n_541), .B(n_460), .Y(n_706) );
O2A1O1Ixp33_ASAP7_75t_L g707 ( .A1(n_522), .A2(n_537), .B(n_561), .C(n_541), .Y(n_707) );
NAND2xp5_ASAP7_75t_L g708 ( .A(n_665), .B(n_615), .Y(n_708) );
NAND2xp5_ASAP7_75t_L g709 ( .A(n_696), .B(n_703), .Y(n_709) );
INVx1_ASAP7_75t_L g710 ( .A(n_705), .Y(n_710) );
INVx8_ASAP7_75t_L g711 ( .A(n_700), .Y(n_711) );
INVx3_ASAP7_75t_L g712 ( .A(n_672), .Y(n_712) );
AOI21xp33_ASAP7_75t_L g713 ( .A1(n_691), .A2(n_707), .B(n_695), .Y(n_713) );
INVx1_ASAP7_75t_L g714 ( .A(n_678), .Y(n_714) );
AOI222xp33_ASAP7_75t_L g715 ( .A1(n_692), .A2(n_706), .B1(n_687), .B2(n_694), .C1(n_629), .C2(n_704), .Y(n_715) );
AOI221xp5_ASAP7_75t_L g716 ( .A1(n_695), .A2(n_653), .B1(n_668), .B2(n_688), .C(n_673), .Y(n_716) );
AO31x2_ASAP7_75t_L g717 ( .A1(n_659), .A2(n_658), .A3(n_621), .B(n_628), .Y(n_717) );
BUFx12f_ASAP7_75t_L g718 ( .A(n_613), .Y(n_718) );
INVx1_ASAP7_75t_L g719 ( .A(n_617), .Y(n_719) );
NAND2xp5_ASAP7_75t_L g720 ( .A(n_649), .B(n_697), .Y(n_720) );
AOI221xp5_ASAP7_75t_L g721 ( .A1(n_620), .A2(n_625), .B1(n_624), .B2(n_667), .C(n_646), .Y(n_721) );
OAI21xp5_ASAP7_75t_L g722 ( .A1(n_686), .A2(n_681), .B(n_683), .Y(n_722) );
OR2x6_ASAP7_75t_L g723 ( .A(n_672), .B(n_617), .Y(n_723) );
NOR2xp33_ASAP7_75t_L g724 ( .A(n_662), .B(n_629), .Y(n_724) );
HB1xp67_ASAP7_75t_L g725 ( .A(n_622), .Y(n_725) );
AOI22xp33_ASAP7_75t_L g726 ( .A1(n_661), .A2(n_616), .B1(n_643), .B2(n_660), .Y(n_726) );
A2O1A1Ixp33_ASAP7_75t_L g727 ( .A1(n_640), .A2(n_647), .B(n_650), .C(n_684), .Y(n_727) );
OR2x6_ASAP7_75t_L g728 ( .A(n_648), .B(n_676), .Y(n_728) );
AND2x2_ASAP7_75t_L g729 ( .A(n_612), .B(n_633), .Y(n_729) );
HB1xp67_ASAP7_75t_L g730 ( .A(n_680), .Y(n_730) );
NOR2xp33_ASAP7_75t_L g731 ( .A(n_671), .B(n_661), .Y(n_731) );
OA21x2_ASAP7_75t_L g732 ( .A1(n_642), .A2(n_637), .B(n_652), .Y(n_732) );
NAND2xp5_ASAP7_75t_L g733 ( .A(n_698), .B(n_702), .Y(n_733) );
AND2x2_ASAP7_75t_L g734 ( .A(n_626), .B(n_666), .Y(n_734) );
NAND2xp5_ASAP7_75t_L g735 ( .A(n_698), .B(n_702), .Y(n_735) );
INVx1_ASAP7_75t_L g736 ( .A(n_611), .Y(n_736) );
OA21x2_ASAP7_75t_L g737 ( .A1(n_654), .A2(n_619), .B(n_630), .Y(n_737) );
AOI21xp5_ASAP7_75t_L g738 ( .A1(n_644), .A2(n_669), .B(n_679), .Y(n_738) );
AOI22xp33_ASAP7_75t_L g739 ( .A1(n_669), .A2(n_675), .B1(n_618), .B2(n_623), .Y(n_739) );
AO21x2_ASAP7_75t_L g740 ( .A1(n_645), .A2(n_631), .B(n_632), .Y(n_740) );
OAI21x1_ASAP7_75t_L g741 ( .A1(n_638), .A2(n_641), .B(n_670), .Y(n_741) );
AND2x2_ASAP7_75t_L g742 ( .A(n_635), .B(n_634), .Y(n_742) );
BUFx4f_ASAP7_75t_L g743 ( .A(n_674), .Y(n_743) );
OR2x2_ASAP7_75t_L g744 ( .A(n_635), .B(n_614), .Y(n_744) );
AND2x4_ASAP7_75t_L g745 ( .A(n_639), .B(n_682), .Y(n_745) );
AOI21xp5_ASAP7_75t_L g746 ( .A1(n_677), .A2(n_639), .B(n_655), .Y(n_746) );
AOI21xp5_ASAP7_75t_L g747 ( .A1(n_636), .A2(n_663), .B(n_690), .Y(n_747) );
OAI22xp5_ASAP7_75t_L g748 ( .A1(n_635), .A2(n_634), .B1(n_614), .B2(n_651), .Y(n_748) );
AOI21xp5_ASAP7_75t_L g749 ( .A1(n_663), .A2(n_690), .B(n_685), .Y(n_749) );
NAND2xp5_ASAP7_75t_L g750 ( .A(n_690), .B(n_685), .Y(n_750) );
OR2x6_ASAP7_75t_L g751 ( .A(n_656), .B(n_657), .Y(n_751) );
OR2x2_ASAP7_75t_L g752 ( .A(n_685), .B(n_656), .Y(n_752) );
INVx1_ASAP7_75t_L g753 ( .A(n_656), .Y(n_753) );
A2O1A1Ixp33_ASAP7_75t_L g754 ( .A1(n_663), .A2(n_701), .B(n_693), .C(n_707), .Y(n_754) );
OAI221xp5_ASAP7_75t_L g755 ( .A1(n_657), .A2(n_458), .B1(n_447), .B2(n_414), .C(n_688), .Y(n_755) );
OAI221xp5_ASAP7_75t_L g756 ( .A1(n_688), .A2(n_458), .B1(n_447), .B2(n_414), .C(n_694), .Y(n_756) );
NAND2xp5_ASAP7_75t_L g757 ( .A(n_665), .B(n_522), .Y(n_757) );
INVx1_ASAP7_75t_L g758 ( .A(n_705), .Y(n_758) );
AND2x2_ASAP7_75t_L g759 ( .A(n_704), .B(n_455), .Y(n_759) );
NAND2xp5_ASAP7_75t_L g760 ( .A(n_665), .B(n_522), .Y(n_760) );
CKINVDCx20_ASAP7_75t_R g761 ( .A(n_700), .Y(n_761) );
AOI22xp33_ASAP7_75t_L g762 ( .A1(n_695), .A2(n_565), .B1(n_541), .B2(n_449), .Y(n_762) );
AND2x2_ASAP7_75t_L g763 ( .A(n_704), .B(n_455), .Y(n_763) );
HB1xp67_ASAP7_75t_L g764 ( .A(n_700), .Y(n_764) );
AOI22xp33_ASAP7_75t_L g765 ( .A1(n_695), .A2(n_565), .B1(n_541), .B2(n_449), .Y(n_765) );
OAI21xp5_ASAP7_75t_SL g766 ( .A1(n_692), .A2(n_452), .B(n_458), .Y(n_766) );
INVx1_ASAP7_75t_L g767 ( .A(n_705), .Y(n_767) );
AND2x2_ASAP7_75t_L g768 ( .A(n_704), .B(n_455), .Y(n_768) );
INVx1_ASAP7_75t_L g769 ( .A(n_705), .Y(n_769) );
OAI221xp5_ASAP7_75t_L g770 ( .A1(n_706), .A2(n_458), .B1(n_447), .B2(n_414), .C(n_451), .Y(n_770) );
AOI21xp5_ASAP7_75t_L g771 ( .A1(n_664), .A2(n_689), .B(n_699), .Y(n_771) );
INVx1_ASAP7_75t_L g772 ( .A(n_705), .Y(n_772) );
CKINVDCx5p33_ASAP7_75t_R g773 ( .A(n_613), .Y(n_773) );
AOI22xp33_ASAP7_75t_L g774 ( .A1(n_695), .A2(n_565), .B1(n_541), .B2(n_449), .Y(n_774) );
AND2x2_ASAP7_75t_L g775 ( .A(n_704), .B(n_455), .Y(n_775) );
AOI22xp33_ASAP7_75t_L g776 ( .A1(n_695), .A2(n_565), .B1(n_541), .B2(n_449), .Y(n_776) );
AOI222xp33_ASAP7_75t_L g777 ( .A1(n_692), .A2(n_449), .B1(n_386), .B2(n_379), .C1(n_385), .C2(n_541), .Y(n_777) );
NAND2xp5_ASAP7_75t_L g778 ( .A(n_665), .B(n_522), .Y(n_778) );
A2O1A1Ixp33_ASAP7_75t_L g779 ( .A1(n_693), .A2(n_701), .B(n_707), .C(n_691), .Y(n_779) );
CKINVDCx6p67_ASAP7_75t_R g780 ( .A(n_613), .Y(n_780) );
OR2x2_ASAP7_75t_L g781 ( .A(n_705), .B(n_455), .Y(n_781) );
OAI21x1_ASAP7_75t_SL g782 ( .A1(n_672), .A2(n_699), .B(n_627), .Y(n_782) );
NAND2x1p5_ASAP7_75t_L g783 ( .A(n_672), .B(n_547), .Y(n_783) );
A2O1A1Ixp33_ASAP7_75t_L g784 ( .A1(n_693), .A2(n_701), .B(n_707), .C(n_691), .Y(n_784) );
BUFx8_ASAP7_75t_L g785 ( .A(n_613), .Y(n_785) );
NAND2xp5_ASAP7_75t_L g786 ( .A(n_665), .B(n_522), .Y(n_786) );
OAI22xp5_ASAP7_75t_L g787 ( .A1(n_699), .A2(n_701), .B1(n_693), .B2(n_696), .Y(n_787) );
A2O1A1Ixp33_ASAP7_75t_L g788 ( .A1(n_693), .A2(n_701), .B(n_707), .C(n_691), .Y(n_788) );
NAND2xp5_ASAP7_75t_L g789 ( .A(n_665), .B(n_522), .Y(n_789) );
OR2x2_ASAP7_75t_L g790 ( .A(n_757), .B(n_760), .Y(n_790) );
NAND2xp5_ASAP7_75t_L g791 ( .A(n_766), .B(n_759), .Y(n_791) );
AND2x2_ASAP7_75t_L g792 ( .A(n_757), .B(n_760), .Y(n_792) );
OR2x2_ASAP7_75t_L g793 ( .A(n_778), .B(n_786), .Y(n_793) );
INVx2_ASAP7_75t_SL g794 ( .A(n_745), .Y(n_794) );
AND2x2_ASAP7_75t_L g795 ( .A(n_778), .B(n_786), .Y(n_795) );
AND2x2_ASAP7_75t_L g796 ( .A(n_789), .B(n_709), .Y(n_796) );
AND2x2_ASAP7_75t_L g797 ( .A(n_709), .B(n_708), .Y(n_797) );
NAND2xp5_ASAP7_75t_L g798 ( .A(n_763), .B(n_768), .Y(n_798) );
OR2x2_ASAP7_75t_L g799 ( .A(n_781), .B(n_723), .Y(n_799) );
AOI221xp5_ASAP7_75t_L g800 ( .A1(n_770), .A2(n_756), .B1(n_755), .B2(n_774), .C(n_765), .Y(n_800) );
NOR2xp33_ASAP7_75t_L g801 ( .A(n_756), .B(n_710), .Y(n_801) );
NAND4xp25_ASAP7_75t_L g802 ( .A(n_777), .B(n_715), .C(n_776), .D(n_762), .Y(n_802) );
AND2x4_ASAP7_75t_L g803 ( .A(n_722), .B(n_723), .Y(n_803) );
OR2x2_ASAP7_75t_L g804 ( .A(n_723), .B(n_775), .Y(n_804) );
AOI22xp33_ASAP7_75t_SL g805 ( .A1(n_755), .A2(n_731), .B1(n_782), .B2(n_711), .Y(n_805) );
NAND3xp33_ASAP7_75t_L g806 ( .A(n_754), .B(n_713), .C(n_788), .Y(n_806) );
HB1xp67_ASAP7_75t_L g807 ( .A(n_725), .Y(n_807) );
NAND2xp5_ASAP7_75t_L g808 ( .A(n_758), .B(n_767), .Y(n_808) );
OR2x2_ASAP7_75t_L g809 ( .A(n_720), .B(n_744), .Y(n_809) );
INVx1_ASAP7_75t_L g810 ( .A(n_742), .Y(n_810) );
OA21x2_ASAP7_75t_L g811 ( .A1(n_747), .A2(n_713), .B(n_753), .Y(n_811) );
INVx2_ASAP7_75t_L g812 ( .A(n_750), .Y(n_812) );
INVx1_ASAP7_75t_L g813 ( .A(n_787), .Y(n_813) );
OR2x6_ASAP7_75t_L g814 ( .A(n_783), .B(n_738), .Y(n_814) );
INVx1_ASAP7_75t_L g815 ( .A(n_787), .Y(n_815) );
AOI22xp33_ASAP7_75t_L g816 ( .A1(n_715), .A2(n_777), .B1(n_716), .B2(n_721), .Y(n_816) );
INVx1_ASAP7_75t_L g817 ( .A(n_748), .Y(n_817) );
INVx1_ASAP7_75t_L g818 ( .A(n_748), .Y(n_818) );
NOR2xp33_ASAP7_75t_L g819 ( .A(n_769), .B(n_772), .Y(n_819) );
NAND2xp5_ASAP7_75t_L g820 ( .A(n_714), .B(n_726), .Y(n_820) );
AND2x4_ASAP7_75t_L g821 ( .A(n_712), .B(n_784), .Y(n_821) );
OR2x6_ASAP7_75t_L g822 ( .A(n_783), .B(n_728), .Y(n_822) );
AND2x2_ASAP7_75t_L g823 ( .A(n_736), .B(n_719), .Y(n_823) );
OR2x2_ASAP7_75t_L g824 ( .A(n_733), .B(n_735), .Y(n_824) );
OR2x6_ASAP7_75t_L g825 ( .A(n_728), .B(n_741), .Y(n_825) );
OAI22xp5_ASAP7_75t_L g826 ( .A1(n_739), .A2(n_743), .B1(n_728), .B2(n_779), .Y(n_826) );
NAND2xp5_ASAP7_75t_L g827 ( .A(n_729), .B(n_734), .Y(n_827) );
OAI221xp5_ASAP7_75t_SL g828 ( .A1(n_771), .A2(n_751), .B1(n_780), .B2(n_724), .C(n_727), .Y(n_828) );
AOI211xp5_ASAP7_75t_SL g829 ( .A1(n_761), .A2(n_764), .B(n_746), .C(n_730), .Y(n_829) );
NAND2xp5_ASAP7_75t_L g830 ( .A(n_711), .B(n_743), .Y(n_830) );
INVx2_ASAP7_75t_L g831 ( .A(n_751), .Y(n_831) );
HB1xp67_ASAP7_75t_L g832 ( .A(n_711), .Y(n_832) );
AND2x2_ASAP7_75t_L g833 ( .A(n_737), .B(n_740), .Y(n_833) );
INVx2_ASAP7_75t_SL g834 ( .A(n_785), .Y(n_834) );
INVx1_ASAP7_75t_L g835 ( .A(n_717), .Y(n_835) );
OA21x2_ASAP7_75t_L g836 ( .A1(n_732), .A2(n_773), .B(n_785), .Y(n_836) );
AND2x2_ASAP7_75t_L g837 ( .A(n_732), .B(n_718), .Y(n_837) );
AND2x2_ASAP7_75t_L g838 ( .A(n_757), .B(n_760), .Y(n_838) );
NAND2xp5_ASAP7_75t_L g839 ( .A(n_766), .B(n_541), .Y(n_839) );
AND2x2_ASAP7_75t_L g840 ( .A(n_757), .B(n_760), .Y(n_840) );
AND2x2_ASAP7_75t_L g841 ( .A(n_757), .B(n_760), .Y(n_841) );
OA21x2_ASAP7_75t_L g842 ( .A1(n_722), .A2(n_754), .B(n_749), .Y(n_842) );
INVx2_ASAP7_75t_L g843 ( .A(n_752), .Y(n_843) );
AND2x2_ASAP7_75t_L g844 ( .A(n_810), .B(n_797), .Y(n_844) );
INVx5_ASAP7_75t_L g845 ( .A(n_822), .Y(n_845) );
AND2x2_ASAP7_75t_L g846 ( .A(n_810), .B(n_797), .Y(n_846) );
OR2x2_ASAP7_75t_L g847 ( .A(n_824), .B(n_809), .Y(n_847) );
AND2x4_ASAP7_75t_L g848 ( .A(n_803), .B(n_831), .Y(n_848) );
AND2x2_ASAP7_75t_L g849 ( .A(n_796), .B(n_792), .Y(n_849) );
NOR2x1_ASAP7_75t_SL g850 ( .A(n_822), .B(n_814), .Y(n_850) );
AND2x2_ASAP7_75t_SL g851 ( .A(n_803), .B(n_836), .Y(n_851) );
AND2x2_ASAP7_75t_L g852 ( .A(n_796), .B(n_792), .Y(n_852) );
AND2x2_ASAP7_75t_L g853 ( .A(n_795), .B(n_838), .Y(n_853) );
AND2x2_ASAP7_75t_L g854 ( .A(n_795), .B(n_838), .Y(n_854) );
NAND2x1p5_ASAP7_75t_SL g855 ( .A(n_837), .B(n_794), .Y(n_855) );
AND2x2_ASAP7_75t_L g856 ( .A(n_840), .B(n_841), .Y(n_856) );
HB1xp67_ASAP7_75t_L g857 ( .A(n_807), .Y(n_857) );
AND2x2_ASAP7_75t_L g858 ( .A(n_813), .B(n_815), .Y(n_858) );
AND2x2_ASAP7_75t_L g859 ( .A(n_813), .B(n_815), .Y(n_859) );
OR2x6_ASAP7_75t_L g860 ( .A(n_825), .B(n_822), .Y(n_860) );
AOI22xp33_ASAP7_75t_L g861 ( .A1(n_802), .A2(n_816), .B1(n_800), .B2(n_801), .Y(n_861) );
HB1xp67_ASAP7_75t_L g862 ( .A(n_812), .Y(n_862) );
AND2x2_ASAP7_75t_L g863 ( .A(n_823), .B(n_817), .Y(n_863) );
AOI22xp33_ASAP7_75t_L g864 ( .A1(n_839), .A2(n_826), .B1(n_791), .B2(n_805), .Y(n_864) );
NAND2xp5_ASAP7_75t_L g865 ( .A(n_790), .B(n_793), .Y(n_865) );
OR2x2_ASAP7_75t_L g866 ( .A(n_820), .B(n_843), .Y(n_866) );
BUFx2_ASAP7_75t_L g867 ( .A(n_843), .Y(n_867) );
AND2x2_ASAP7_75t_L g868 ( .A(n_818), .B(n_833), .Y(n_868) );
NAND3xp33_ASAP7_75t_L g869 ( .A(n_861), .B(n_829), .C(n_828), .Y(n_869) );
AND2x2_ASAP7_75t_L g870 ( .A(n_863), .B(n_833), .Y(n_870) );
AND2x2_ASAP7_75t_L g871 ( .A(n_863), .B(n_842), .Y(n_871) );
NAND2xp5_ASAP7_75t_L g872 ( .A(n_858), .B(n_806), .Y(n_872) );
OR2x2_ASAP7_75t_L g873 ( .A(n_847), .B(n_835), .Y(n_873) );
INVx2_ASAP7_75t_SL g874 ( .A(n_845), .Y(n_874) );
NOR3xp33_ASAP7_75t_SL g875 ( .A(n_865), .B(n_830), .C(n_819), .Y(n_875) );
NAND2xp5_ASAP7_75t_L g876 ( .A(n_859), .B(n_806), .Y(n_876) );
NOR2xp33_ASAP7_75t_L g877 ( .A(n_853), .B(n_834), .Y(n_877) );
INVxp67_ASAP7_75t_SL g878 ( .A(n_862), .Y(n_878) );
NOR3xp33_ASAP7_75t_SL g879 ( .A(n_865), .B(n_827), .C(n_798), .Y(n_879) );
INVxp67_ASAP7_75t_L g880 ( .A(n_857), .Y(n_880) );
AND2x2_ASAP7_75t_L g881 ( .A(n_868), .B(n_811), .Y(n_881) );
NOR2xp33_ASAP7_75t_L g882 ( .A(n_854), .B(n_832), .Y(n_882) );
AND2x2_ASAP7_75t_L g883 ( .A(n_844), .B(n_811), .Y(n_883) );
AND2x2_ASAP7_75t_L g884 ( .A(n_846), .B(n_811), .Y(n_884) );
AND2x2_ASAP7_75t_L g885 ( .A(n_846), .B(n_835), .Y(n_885) );
AOI22xp33_ASAP7_75t_L g886 ( .A1(n_869), .A2(n_864), .B1(n_851), .B2(n_821), .Y(n_886) );
CKINVDCx16_ASAP7_75t_R g887 ( .A(n_877), .Y(n_887) );
NAND2xp5_ASAP7_75t_L g888 ( .A(n_885), .B(n_849), .Y(n_888) );
INVx2_ASAP7_75t_SL g889 ( .A(n_874), .Y(n_889) );
AND2x2_ASAP7_75t_L g890 ( .A(n_883), .B(n_851), .Y(n_890) );
OR2x2_ASAP7_75t_L g891 ( .A(n_883), .B(n_866), .Y(n_891) );
AND2x2_ASAP7_75t_L g892 ( .A(n_884), .B(n_848), .Y(n_892) );
OR2x2_ASAP7_75t_L g893 ( .A(n_884), .B(n_866), .Y(n_893) );
BUFx2_ASAP7_75t_L g894 ( .A(n_878), .Y(n_894) );
OR2x2_ASAP7_75t_L g895 ( .A(n_872), .B(n_867), .Y(n_895) );
INVx1_ASAP7_75t_L g896 ( .A(n_880), .Y(n_896) );
NAND2xp5_ASAP7_75t_L g897 ( .A(n_885), .B(n_849), .Y(n_897) );
NAND2xp5_ASAP7_75t_L g898 ( .A(n_870), .B(n_852), .Y(n_898) );
NAND2xp5_ASAP7_75t_L g899 ( .A(n_876), .B(n_856), .Y(n_899) );
AOI22xp5_ASAP7_75t_L g900 ( .A1(n_886), .A2(n_869), .B1(n_879), .B2(n_875), .Y(n_900) );
AND2x2_ASAP7_75t_L g901 ( .A(n_892), .B(n_881), .Y(n_901) );
HB1xp67_ASAP7_75t_L g902 ( .A(n_894), .Y(n_902) );
INVxp67_ASAP7_75t_SL g903 ( .A(n_894), .Y(n_903) );
NAND2xp5_ASAP7_75t_L g904 ( .A(n_899), .B(n_871), .Y(n_904) );
OR2x2_ASAP7_75t_L g905 ( .A(n_891), .B(n_873), .Y(n_905) );
CKINVDCx16_ASAP7_75t_R g906 ( .A(n_887), .Y(n_906) );
INVx1_ASAP7_75t_SL g907 ( .A(n_893), .Y(n_907) );
INVx2_ASAP7_75t_SL g908 ( .A(n_889), .Y(n_908) );
INVx1_ASAP7_75t_L g909 ( .A(n_905), .Y(n_909) );
INVx2_ASAP7_75t_SL g910 ( .A(n_908), .Y(n_910) );
NAND2xp5_ASAP7_75t_L g911 ( .A(n_907), .B(n_896), .Y(n_911) );
AOI322xp5_ASAP7_75t_L g912 ( .A1(n_906), .A2(n_879), .A3(n_898), .B1(n_897), .B2(n_888), .C1(n_882), .C2(n_890), .Y(n_912) );
HB1xp67_ASAP7_75t_L g913 ( .A(n_902), .Y(n_913) );
OAI21xp5_ASAP7_75t_L g914 ( .A1(n_912), .A2(n_900), .B(n_903), .Y(n_914) );
AND2x2_ASAP7_75t_L g915 ( .A(n_910), .B(n_901), .Y(n_915) );
NAND2xp5_ASAP7_75t_L g916 ( .A(n_909), .B(n_904), .Y(n_916) );
NAND3xp33_ASAP7_75t_L g917 ( .A(n_914), .B(n_913), .C(n_911), .Y(n_917) );
O2A1O1Ixp33_ASAP7_75t_L g918 ( .A1(n_917), .A2(n_808), .B(n_915), .C(n_916), .Y(n_918) );
INVx1_ASAP7_75t_L g919 ( .A(n_918), .Y(n_919) );
INVx1_ASAP7_75t_L g920 ( .A(n_919), .Y(n_920) );
INVx2_ASAP7_75t_L g921 ( .A(n_920), .Y(n_921) );
INVx2_ASAP7_75t_L g922 ( .A(n_921), .Y(n_922) );
AOI21xp33_ASAP7_75t_SL g923 ( .A1(n_922), .A2(n_855), .B(n_799), .Y(n_923) );
AOI22xp5_ASAP7_75t_L g924 ( .A1(n_923), .A2(n_821), .B1(n_845), .B2(n_860), .Y(n_924) );
AO21x2_ASAP7_75t_L g925 ( .A1(n_924), .A2(n_855), .B(n_850), .Y(n_925) );
AOI21xp33_ASAP7_75t_L g926 ( .A1(n_925), .A2(n_804), .B(n_895), .Y(n_926) );
endmodule