module fake_netlist_6_3065_n_1265 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_166, n_28, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_173, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_171, n_31, n_57, n_169, n_53, n_51, n_44, n_56, n_1265);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_173;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_171;
input n_31;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1265;

wire n_992;
wire n_801;
wire n_1234;
wire n_1199;
wire n_741;
wire n_1027;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1038;
wire n_578;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_783;
wire n_798;
wire n_188;
wire n_509;
wire n_245;
wire n_1209;
wire n_677;
wire n_805;
wire n_1151;
wire n_396;
wire n_350;
wire n_442;
wire n_480;
wire n_1009;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1032;
wire n_1247;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_200;
wire n_447;
wire n_1172;
wire n_852;
wire n_229;
wire n_1078;
wire n_250;
wire n_544;
wire n_1140;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1143;
wire n_1232;
wire n_658;
wire n_616;
wire n_1119;
wire n_428;
wire n_641;
wire n_822;
wire n_693;
wire n_1056;
wire n_758;
wire n_516;
wire n_1163;
wire n_1180;
wire n_943;
wire n_491;
wire n_772;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_343;
wire n_953;
wire n_1094;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_638;
wire n_1211;
wire n_381;
wire n_887;
wire n_713;
wire n_976;
wire n_224;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_659;
wire n_407;
wire n_913;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_577;
wire n_619;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_323;
wire n_606;
wire n_818;
wire n_1123;
wire n_513;
wire n_645;
wire n_331;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_788;
wire n_939;
wire n_821;
wire n_938;
wire n_1068;
wire n_329;
wire n_982;
wire n_549;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_243;
wire n_979;
wire n_905;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_547;
wire n_558;
wire n_1064;
wire n_634;
wire n_966;
wire n_764;
wire n_692;
wire n_733;
wire n_1233;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_882;
wire n_586;
wire n_423;
wire n_318;
wire n_1111;
wire n_715;
wire n_1251;
wire n_530;
wire n_277;
wire n_618;
wire n_199;
wire n_1167;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_210;
wire n_1069;
wire n_612;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_429;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_286;
wire n_254;
wire n_242;
wire n_835;
wire n_1214;
wire n_928;
wire n_690;
wire n_850;
wire n_816;
wire n_1157;
wire n_1188;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_267;
wire n_1124;
wire n_515;
wire n_598;
wire n_696;
wire n_961;
wire n_437;
wire n_1082;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_891;
wire n_949;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_881;
wire n_1008;
wire n_760;
wire n_590;
wire n_362;
wire n_1033;
wire n_462;
wire n_1052;
wire n_304;
wire n_694;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_342;
wire n_1044;
wire n_449;
wire n_1208;
wire n_1164;
wire n_1072;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_840;
wire n_874;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_615;
wire n_1249;
wire n_1127;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_353;
wire n_605;
wire n_826;
wire n_872;
wire n_1139;
wire n_718;
wire n_1018;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_622;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_631;
wire n_720;
wire n_842;
wire n_843;
wire n_656;
wire n_989;
wire n_797;
wire n_1246;
wire n_899;
wire n_189;
wire n_738;
wire n_1035;
wire n_294;
wire n_499;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_648;
wire n_657;
wire n_1049;
wire n_803;
wire n_290;
wire n_926;
wire n_927;
wire n_919;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_777;
wire n_272;
wire n_526;
wire n_1183;
wire n_293;
wire n_1070;
wire n_458;
wire n_998;
wire n_717;
wire n_1178;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_184;
wire n_552;
wire n_216;
wire n_912;
wire n_745;
wire n_1142;
wire n_716;
wire n_623;
wire n_1048;
wire n_1201;
wire n_884;
wire n_731;
wire n_755;
wire n_931;
wire n_1021;
wire n_527;
wire n_683;
wire n_811;
wire n_1207;
wire n_474;
wire n_312;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_589;
wire n_819;
wire n_767;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_399;
wire n_211;
wire n_231;
wire n_505;
wire n_319;
wire n_537;
wire n_311;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_386;
wire n_1220;
wire n_556;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1053;
wire n_416;
wire n_520;
wire n_418;
wire n_1093;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_217;
wire n_518;
wire n_1185;
wire n_453;
wire n_215;
wire n_914;
wire n_759;
wire n_426;
wire n_317;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1224;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_335;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_983;
wire n_427;
wire n_496;
wire n_906;
wire n_688;
wire n_1077;
wire n_351;
wire n_259;
wire n_385;
wire n_858;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_664;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_580;
wire n_762;
wire n_1202;
wire n_1030;
wire n_465;
wire n_1079;
wire n_341;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_485;
wire n_443;
wire n_892;
wire n_768;
wire n_421;
wire n_238;
wire n_1095;
wire n_202;
wire n_597;
wire n_280;
wire n_1187;
wire n_610;
wire n_1024;
wire n_198;
wire n_179;
wire n_248;
wire n_517;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1115;
wire n_750;
wire n_901;
wire n_468;
wire n_923;
wire n_504;
wire n_183;
wire n_1015;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1182;
wire n_785;
wire n_746;
wire n_609;
wire n_1168;
wire n_1216;
wire n_302;
wire n_380;
wire n_1190;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_239;
wire n_782;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_986;
wire n_1081;
wire n_402;
wire n_352;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_662;
wire n_374;
wire n_1152;
wire n_450;
wire n_921;
wire n_711;
wire n_579;
wire n_937;
wire n_370;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_258;
wire n_456;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_936;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_227;
wire n_204;
wire n_482;
wire n_934;
wire n_420;
wire n_394;
wire n_942;
wire n_543;
wire n_1225;
wire n_325;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_548;
wire n_282;
wire n_833;
wire n_523;
wire n_707;
wire n_345;
wire n_799;
wire n_1155;
wire n_273;
wire n_787;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1241;
wire n_569;
wire n_737;
wire n_1235;
wire n_1229;
wire n_306;
wire n_346;
wire n_1029;
wire n_790;
wire n_1210;
wire n_299;
wire n_1248;
wire n_902;
wire n_333;
wire n_1047;
wire n_431;
wire n_459;
wire n_502;
wire n_672;
wire n_1257;
wire n_285;
wire n_655;
wire n_706;
wire n_1045;
wire n_786;
wire n_1236;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1002;
wire n_545;
wire n_489;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_660;
wire n_438;
wire n_1200;
wire n_479;
wire n_869;
wire n_1154;
wire n_1113;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1177;
wire n_332;
wire n_1150;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_194;
wire n_1007;
wire n_855;
wire n_591;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_661;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1217;
wire n_751;
wire n_749;
wire n_310;
wire n_969;
wire n_988;
wire n_1065;
wire n_1255;
wire n_568;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_214;
wire n_246;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1130;
wire n_181;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_555;
wire n_389;
wire n_814;
wire n_669;
wire n_300;
wire n_222;
wire n_747;
wire n_1105;
wire n_721;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_378;
wire n_1196;
wire n_377;
wire n_863;
wire n_601;
wire n_338;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1147;
wire n_360;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1205;
wire n_1258;
wire n_1173;
wire n_525;
wire n_1116;
wire n_611;
wire n_1219;
wire n_1174;
wire n_1016;
wire n_795;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_911;
wire n_653;
wire n_236;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_779;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_366;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_719;
wire n_228;
wire n_455;
wire n_363;
wire n_1090;
wire n_592;
wire n_829;
wire n_1156;
wire n_393;
wire n_984;
wire n_503;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_981;
wire n_714;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_802;
wire n_561;
wire n_980;
wire n_1198;
wire n_436;
wire n_409;
wire n_1244;
wire n_240;
wire n_756;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1034;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_553;
wire n_849;
wire n_753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1055;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_271;
wire n_404;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_534;
wire n_1006;
wire n_373;
wire n_257;
wire n_730;
wire n_670;
wire n_203;
wire n_207;
wire n_1089;
wire n_205;
wire n_1242;
wire n_681;
wire n_1226;
wire n_412;
wire n_640;
wire n_965;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_457;
wire n_364;
wire n_629;
wire n_900;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_192;
wire n_649;
wire n_1240;

INVx2_ASAP7_75t_L g179 ( 
.A(n_125),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_133),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_11),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_46),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_56),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_82),
.Y(n_184)
);

BUFx2_ASAP7_75t_L g185 ( 
.A(n_129),
.Y(n_185)
);

BUFx3_ASAP7_75t_L g186 ( 
.A(n_149),
.Y(n_186)
);

BUFx10_ASAP7_75t_L g187 ( 
.A(n_114),
.Y(n_187)
);

CKINVDCx16_ASAP7_75t_R g188 ( 
.A(n_53),
.Y(n_188)
);

BUFx6f_ASAP7_75t_L g189 ( 
.A(n_168),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_40),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_20),
.Y(n_191)
);

BUFx10_ASAP7_75t_L g192 ( 
.A(n_98),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_106),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_7),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_6),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_69),
.Y(n_196)
);

INVx2_ASAP7_75t_SL g197 ( 
.A(n_14),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_22),
.Y(n_198)
);

BUFx3_ASAP7_75t_L g199 ( 
.A(n_64),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_111),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_134),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_150),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_65),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_32),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_25),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_131),
.Y(n_206)
);

BUFx8_ASAP7_75t_SL g207 ( 
.A(n_97),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_124),
.Y(n_208)
);

INVxp67_ASAP7_75t_L g209 ( 
.A(n_119),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_79),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_57),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_71),
.Y(n_212)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_72),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_171),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_107),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_19),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_137),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_96),
.Y(n_218)
);

INVx2_ASAP7_75t_SL g219 ( 
.A(n_0),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_123),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_30),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_172),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_50),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_63),
.Y(n_224)
);

INVx2_ASAP7_75t_SL g225 ( 
.A(n_10),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_61),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_116),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_120),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_105),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_100),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_14),
.Y(n_231)
);

BUFx6f_ASAP7_75t_L g232 ( 
.A(n_27),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_164),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_10),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_142),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_38),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_191),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_194),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_195),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_182),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_183),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_184),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_190),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_193),
.Y(n_244)
);

BUFx10_ASAP7_75t_L g245 ( 
.A(n_232),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_196),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_232),
.Y(n_247)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_232),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_200),
.Y(n_249)
);

BUFx10_ASAP7_75t_L g250 ( 
.A(n_232),
.Y(n_250)
);

INVx1_ASAP7_75t_SL g251 ( 
.A(n_198),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_181),
.Y(n_252)
);

BUFx10_ASAP7_75t_L g253 ( 
.A(n_204),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_201),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_214),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_202),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_203),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_206),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_216),
.Y(n_259)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_189),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_186),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_208),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_215),
.Y(n_263)
);

INVx2_ASAP7_75t_SL g264 ( 
.A(n_197),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_211),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_218),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_240),
.Y(n_267)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_248),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_241),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_242),
.Y(n_270)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_248),
.Y(n_271)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_260),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_260),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_243),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_244),
.Y(n_275)
);

BUFx3_ASAP7_75t_L g276 ( 
.A(n_245),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_247),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_249),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_252),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_246),
.Y(n_280)
);

BUFx3_ASAP7_75t_L g281 ( 
.A(n_245),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_259),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_256),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_257),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_245),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_254),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_250),
.Y(n_287)
);

INVxp33_ASAP7_75t_SL g288 ( 
.A(n_258),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_262),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_265),
.B(n_186),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_237),
.Y(n_291)
);

HB1xp67_ASAP7_75t_L g292 ( 
.A(n_237),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_250),
.Y(n_293)
);

INVxp33_ASAP7_75t_L g294 ( 
.A(n_261),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_250),
.Y(n_295)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_264),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_264),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_238),
.Y(n_298)
);

INVxp33_ASAP7_75t_L g299 ( 
.A(n_251),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_238),
.Y(n_300)
);

NOR2xp67_ASAP7_75t_L g301 ( 
.A(n_239),
.B(n_209),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_239),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_255),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_266),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_253),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_253),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_253),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_263),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_240),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_248),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_240),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_248),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_248),
.Y(n_313)
);

HB1xp67_ASAP7_75t_L g314 ( 
.A(n_237),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_240),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_248),
.Y(n_316)
);

BUFx6f_ASAP7_75t_L g317 ( 
.A(n_248),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_240),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_277),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_279),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_267),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_277),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_269),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_272),
.Y(n_324)
);

INVxp33_ASAP7_75t_SL g325 ( 
.A(n_303),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_270),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_272),
.Y(n_327)
);

INVxp67_ASAP7_75t_SL g328 ( 
.A(n_317),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_268),
.Y(n_329)
);

INVxp33_ASAP7_75t_SL g330 ( 
.A(n_304),
.Y(n_330)
);

INVxp67_ASAP7_75t_SL g331 ( 
.A(n_317),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_274),
.Y(n_332)
);

INVxp67_ASAP7_75t_SL g333 ( 
.A(n_317),
.Y(n_333)
);

INVxp33_ASAP7_75t_SL g334 ( 
.A(n_275),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_268),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_271),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_271),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_278),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_273),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_273),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_279),
.Y(n_341)
);

BUFx3_ASAP7_75t_L g342 ( 
.A(n_276),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_280),
.Y(n_343)
);

BUFx2_ASAP7_75t_SL g344 ( 
.A(n_301),
.Y(n_344)
);

XNOR2xp5_ASAP7_75t_L g345 ( 
.A(n_299),
.B(n_198),
.Y(n_345)
);

INVxp33_ASAP7_75t_SL g346 ( 
.A(n_283),
.Y(n_346)
);

INVxp67_ASAP7_75t_SL g347 ( 
.A(n_317),
.Y(n_347)
);

INVx2_ASAP7_75t_L g348 ( 
.A(n_310),
.Y(n_348)
);

CKINVDCx16_ASAP7_75t_R g349 ( 
.A(n_286),
.Y(n_349)
);

INVxp33_ASAP7_75t_SL g350 ( 
.A(n_284),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_310),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_312),
.Y(n_352)
);

INVx2_ASAP7_75t_L g353 ( 
.A(n_312),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_313),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_282),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_282),
.Y(n_356)
);

INVxp67_ASAP7_75t_L g357 ( 
.A(n_292),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_317),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_313),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_316),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_316),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_289),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_296),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_309),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_296),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_297),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_297),
.Y(n_367)
);

INVxp33_ASAP7_75t_L g368 ( 
.A(n_314),
.Y(n_368)
);

HB1xp67_ASAP7_75t_L g369 ( 
.A(n_285),
.Y(n_369)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_348),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_320),
.B(n_290),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_344),
.B(n_288),
.Y(n_372)
);

INVx4_ASAP7_75t_L g373 ( 
.A(n_348),
.Y(n_373)
);

INVx2_ASAP7_75t_L g374 ( 
.A(n_353),
.Y(n_374)
);

BUFx3_ASAP7_75t_L g375 ( 
.A(n_342),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_341),
.B(n_298),
.Y(n_376)
);

AND2x4_ASAP7_75t_L g377 ( 
.A(n_355),
.B(n_199),
.Y(n_377)
);

HB1xp67_ASAP7_75t_L g378 ( 
.A(n_345),
.Y(n_378)
);

AND2x4_ASAP7_75t_L g379 ( 
.A(n_356),
.B(n_199),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_319),
.B(n_298),
.Y(n_380)
);

BUFx6f_ASAP7_75t_L g381 ( 
.A(n_319),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_322),
.B(n_300),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_353),
.Y(n_383)
);

BUFx6f_ASAP7_75t_L g384 ( 
.A(n_322),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_L g385 ( 
.A(n_344),
.B(n_300),
.Y(n_385)
);

INVx3_ASAP7_75t_L g386 ( 
.A(n_339),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_339),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_366),
.B(n_302),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_366),
.B(n_302),
.Y(n_389)
);

NOR2xp33_ASAP7_75t_L g390 ( 
.A(n_369),
.B(n_291),
.Y(n_390)
);

BUFx6f_ASAP7_75t_L g391 ( 
.A(n_358),
.Y(n_391)
);

AND2x2_ASAP7_75t_L g392 ( 
.A(n_367),
.B(n_294),
.Y(n_392)
);

AND2x4_ASAP7_75t_L g393 ( 
.A(n_367),
.B(n_180),
.Y(n_393)
);

BUFx2_ASAP7_75t_L g394 ( 
.A(n_345),
.Y(n_394)
);

BUFx6f_ASAP7_75t_L g395 ( 
.A(n_340),
.Y(n_395)
);

AND2x4_ASAP7_75t_L g396 ( 
.A(n_363),
.B(n_220),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_351),
.Y(n_397)
);

INVx5_ASAP7_75t_L g398 ( 
.A(n_342),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_351),
.Y(n_399)
);

AND2x6_ASAP7_75t_L g400 ( 
.A(n_352),
.B(n_179),
.Y(n_400)
);

INVx5_ASAP7_75t_L g401 ( 
.A(n_328),
.Y(n_401)
);

INVx4_ASAP7_75t_L g402 ( 
.A(n_324),
.Y(n_402)
);

AND2x4_ASAP7_75t_L g403 ( 
.A(n_363),
.B(n_233),
.Y(n_403)
);

AND2x2_ASAP7_75t_L g404 ( 
.A(n_365),
.B(n_352),
.Y(n_404)
);

NOR2xp33_ASAP7_75t_L g405 ( 
.A(n_368),
.B(n_311),
.Y(n_405)
);

AND2x4_ASAP7_75t_L g406 ( 
.A(n_365),
.B(n_185),
.Y(n_406)
);

HB1xp67_ASAP7_75t_L g407 ( 
.A(n_357),
.Y(n_407)
);

INVx4_ASAP7_75t_L g408 ( 
.A(n_324),
.Y(n_408)
);

AND2x4_ASAP7_75t_L g409 ( 
.A(n_354),
.B(n_179),
.Y(n_409)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_354),
.Y(n_410)
);

INVx5_ASAP7_75t_L g411 ( 
.A(n_331),
.Y(n_411)
);

AND2x4_ASAP7_75t_L g412 ( 
.A(n_359),
.B(n_213),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_359),
.Y(n_413)
);

AND2x2_ASAP7_75t_L g414 ( 
.A(n_360),
.B(n_285),
.Y(n_414)
);

BUFx12f_ASAP7_75t_L g415 ( 
.A(n_321),
.Y(n_415)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_410),
.Y(n_416)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_410),
.Y(n_417)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_370),
.Y(n_418)
);

NOR2xp33_ASAP7_75t_L g419 ( 
.A(n_385),
.B(n_334),
.Y(n_419)
);

INVx4_ASAP7_75t_L g420 ( 
.A(n_381),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_371),
.B(n_315),
.Y(n_421)
);

BUFx6f_ASAP7_75t_L g422 ( 
.A(n_381),
.Y(n_422)
);

BUFx12f_ASAP7_75t_L g423 ( 
.A(n_415),
.Y(n_423)
);

BUFx6f_ASAP7_75t_L g424 ( 
.A(n_381),
.Y(n_424)
);

OAI21x1_ASAP7_75t_L g425 ( 
.A1(n_386),
.A2(n_361),
.B(n_360),
.Y(n_425)
);

OA21x2_ASAP7_75t_L g426 ( 
.A1(n_387),
.A2(n_361),
.B(n_329),
.Y(n_426)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_370),
.Y(n_427)
);

INVx3_ASAP7_75t_L g428 ( 
.A(n_381),
.Y(n_428)
);

INVx2_ASAP7_75t_SL g429 ( 
.A(n_392),
.Y(n_429)
);

INVx3_ASAP7_75t_L g430 ( 
.A(n_381),
.Y(n_430)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_374),
.Y(n_431)
);

INVx3_ASAP7_75t_L g432 ( 
.A(n_384),
.Y(n_432)
);

INVx2_ASAP7_75t_L g433 ( 
.A(n_374),
.Y(n_433)
);

AOI22xp5_ASAP7_75t_L g434 ( 
.A1(n_384),
.A2(n_318),
.B1(n_350),
.B2(n_346),
.Y(n_434)
);

OAI22x1_ASAP7_75t_SL g435 ( 
.A1(n_394),
.A2(n_325),
.B1(n_330),
.B2(n_338),
.Y(n_435)
);

NAND2xp33_ASAP7_75t_SL g436 ( 
.A(n_384),
.B(n_210),
.Y(n_436)
);

OAI22xp5_ASAP7_75t_SL g437 ( 
.A1(n_394),
.A2(n_349),
.B1(n_308),
.B2(n_362),
.Y(n_437)
);

OA21x2_ASAP7_75t_L g438 ( 
.A1(n_387),
.A2(n_329),
.B(n_327),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_404),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_380),
.B(n_333),
.Y(n_440)
);

CKINVDCx20_ASAP7_75t_R g441 ( 
.A(n_378),
.Y(n_441)
);

AOI22xp5_ASAP7_75t_L g442 ( 
.A1(n_384),
.A2(n_227),
.B1(n_210),
.B2(n_224),
.Y(n_442)
);

BUFx6f_ASAP7_75t_L g443 ( 
.A(n_395),
.Y(n_443)
);

OAI22xp5_ASAP7_75t_L g444 ( 
.A1(n_382),
.A2(n_226),
.B1(n_224),
.B2(n_343),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_404),
.B(n_347),
.Y(n_445)
);

CKINVDCx20_ASAP7_75t_R g446 ( 
.A(n_415),
.Y(n_446)
);

BUFx6f_ASAP7_75t_L g447 ( 
.A(n_395),
.Y(n_447)
);

NOR2xp33_ASAP7_75t_L g448 ( 
.A(n_372),
.B(n_390),
.Y(n_448)
);

AOI22xp5_ASAP7_75t_L g449 ( 
.A1(n_414),
.A2(n_226),
.B1(n_364),
.B2(n_332),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_397),
.Y(n_450)
);

INVx2_ASAP7_75t_L g451 ( 
.A(n_397),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_399),
.Y(n_452)
);

XNOR2x2_ASAP7_75t_L g453 ( 
.A(n_405),
.B(n_308),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_399),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_414),
.B(n_305),
.Y(n_455)
);

AND2x2_ASAP7_75t_SL g456 ( 
.A(n_393),
.B(n_213),
.Y(n_456)
);

INVx2_ASAP7_75t_L g457 ( 
.A(n_413),
.Y(n_457)
);

BUFx6f_ASAP7_75t_L g458 ( 
.A(n_395),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_413),
.Y(n_459)
);

OAI21x1_ASAP7_75t_L g460 ( 
.A1(n_383),
.A2(n_335),
.B(n_327),
.Y(n_460)
);

AND2x2_ASAP7_75t_L g461 ( 
.A(n_392),
.B(n_305),
.Y(n_461)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_383),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_388),
.B(n_306),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_395),
.Y(n_464)
);

INVx3_ASAP7_75t_L g465 ( 
.A(n_373),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_389),
.B(n_306),
.Y(n_466)
);

OAI22xp5_ASAP7_75t_SL g467 ( 
.A1(n_407),
.A2(n_323),
.B1(n_326),
.B2(n_307),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_376),
.B(n_307),
.Y(n_468)
);

AND2x4_ASAP7_75t_L g469 ( 
.A(n_375),
.B(n_398),
.Y(n_469)
);

CKINVDCx20_ASAP7_75t_R g470 ( 
.A(n_375),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_395),
.Y(n_471)
);

BUFx8_ASAP7_75t_SL g472 ( 
.A(n_406),
.Y(n_472)
);

BUFx6f_ASAP7_75t_L g473 ( 
.A(n_391),
.Y(n_473)
);

INVx5_ASAP7_75t_L g474 ( 
.A(n_400),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_402),
.Y(n_475)
);

HB1xp67_ASAP7_75t_L g476 ( 
.A(n_377),
.Y(n_476)
);

AOI22xp5_ASAP7_75t_L g477 ( 
.A1(n_393),
.A2(n_188),
.B1(n_295),
.B2(n_293),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_402),
.Y(n_478)
);

AND2x2_ASAP7_75t_L g479 ( 
.A(n_406),
.B(n_287),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_402),
.Y(n_480)
);

OAI21x1_ASAP7_75t_L g481 ( 
.A1(n_373),
.A2(n_337),
.B(n_336),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_393),
.B(n_373),
.Y(n_482)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_373),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_402),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_393),
.B(n_337),
.Y(n_485)
);

OR2x2_ASAP7_75t_L g486 ( 
.A(n_406),
.B(n_287),
.Y(n_486)
);

INVx3_ASAP7_75t_L g487 ( 
.A(n_408),
.Y(n_487)
);

OA21x2_ASAP7_75t_L g488 ( 
.A1(n_412),
.A2(n_295),
.B(n_293),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_412),
.B(n_276),
.Y(n_489)
);

INVx2_ASAP7_75t_SL g490 ( 
.A(n_406),
.Y(n_490)
);

AND2x4_ASAP7_75t_L g491 ( 
.A(n_398),
.B(n_396),
.Y(n_491)
);

OAI22xp5_ASAP7_75t_SL g492 ( 
.A1(n_398),
.A2(n_221),
.B1(n_205),
.B2(n_234),
.Y(n_492)
);

INVx3_ASAP7_75t_L g493 ( 
.A(n_408),
.Y(n_493)
);

INVx2_ASAP7_75t_L g494 ( 
.A(n_408),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_409),
.B(n_281),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_408),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_409),
.Y(n_497)
);

BUFx6f_ASAP7_75t_L g498 ( 
.A(n_391),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_409),
.Y(n_499)
);

OA21x2_ASAP7_75t_L g500 ( 
.A1(n_412),
.A2(n_217),
.B(n_212),
.Y(n_500)
);

INVx2_ASAP7_75t_L g501 ( 
.A(n_391),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_412),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_451),
.Y(n_503)
);

AND2x4_ASAP7_75t_L g504 ( 
.A(n_469),
.B(n_398),
.Y(n_504)
);

INVxp67_ASAP7_75t_L g505 ( 
.A(n_461),
.Y(n_505)
);

CKINVDCx5p33_ASAP7_75t_R g506 ( 
.A(n_423),
.Y(n_506)
);

BUFx6f_ASAP7_75t_L g507 ( 
.A(n_422),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_451),
.Y(n_508)
);

AND2x2_ASAP7_75t_SL g509 ( 
.A(n_456),
.B(n_396),
.Y(n_509)
);

BUFx3_ASAP7_75t_L g510 ( 
.A(n_470),
.Y(n_510)
);

CKINVDCx5p33_ASAP7_75t_R g511 ( 
.A(n_423),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_457),
.Y(n_512)
);

CKINVDCx5p33_ASAP7_75t_R g513 ( 
.A(n_446),
.Y(n_513)
);

CKINVDCx5p33_ASAP7_75t_R g514 ( 
.A(n_446),
.Y(n_514)
);

CKINVDCx5p33_ASAP7_75t_R g515 ( 
.A(n_435),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_457),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_448),
.B(n_439),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_462),
.Y(n_518)
);

NOR2xp33_ASAP7_75t_L g519 ( 
.A(n_448),
.B(n_398),
.Y(n_519)
);

INVx2_ASAP7_75t_L g520 ( 
.A(n_416),
.Y(n_520)
);

BUFx2_ASAP7_75t_L g521 ( 
.A(n_470),
.Y(n_521)
);

NOR2xp33_ASAP7_75t_R g522 ( 
.A(n_436),
.B(n_398),
.Y(n_522)
);

CKINVDCx5p33_ASAP7_75t_R g523 ( 
.A(n_472),
.Y(n_523)
);

NAND2xp33_ASAP7_75t_SL g524 ( 
.A(n_422),
.B(n_391),
.Y(n_524)
);

CKINVDCx5p33_ASAP7_75t_R g525 ( 
.A(n_472),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_462),
.Y(n_526)
);

INVx4_ASAP7_75t_L g527 ( 
.A(n_422),
.Y(n_527)
);

CKINVDCx5p33_ASAP7_75t_R g528 ( 
.A(n_437),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_416),
.Y(n_529)
);

BUFx2_ASAP7_75t_L g530 ( 
.A(n_441),
.Y(n_530)
);

INVx2_ASAP7_75t_L g531 ( 
.A(n_417),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_417),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_419),
.B(n_377),
.Y(n_533)
);

INVx2_ASAP7_75t_L g534 ( 
.A(n_483),
.Y(n_534)
);

BUFx3_ASAP7_75t_L g535 ( 
.A(n_441),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_L g536 ( 
.A(n_419),
.B(n_377),
.Y(n_536)
);

CKINVDCx5p33_ASAP7_75t_R g537 ( 
.A(n_434),
.Y(n_537)
);

AND2x4_ASAP7_75t_L g538 ( 
.A(n_469),
.B(n_377),
.Y(n_538)
);

INVx2_ASAP7_75t_L g539 ( 
.A(n_483),
.Y(n_539)
);

INVx2_ASAP7_75t_L g540 ( 
.A(n_418),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_L g541 ( 
.A(n_421),
.B(n_379),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_450),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_452),
.Y(n_543)
);

INVx2_ASAP7_75t_L g544 ( 
.A(n_418),
.Y(n_544)
);

CKINVDCx5p33_ASAP7_75t_R g545 ( 
.A(n_467),
.Y(n_545)
);

CKINVDCx16_ASAP7_75t_R g546 ( 
.A(n_449),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_454),
.Y(n_547)
);

NOR2xp33_ASAP7_75t_L g548 ( 
.A(n_444),
.B(n_379),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_459),
.Y(n_549)
);

INVx3_ASAP7_75t_L g550 ( 
.A(n_465),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_427),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_427),
.Y(n_552)
);

BUFx6f_ASAP7_75t_L g553 ( 
.A(n_422),
.Y(n_553)
);

CKINVDCx20_ASAP7_75t_R g554 ( 
.A(n_442),
.Y(n_554)
);

CKINVDCx20_ASAP7_75t_R g555 ( 
.A(n_436),
.Y(n_555)
);

INVx3_ASAP7_75t_L g556 ( 
.A(n_465),
.Y(n_556)
);

CKINVDCx20_ASAP7_75t_R g557 ( 
.A(n_492),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_431),
.Y(n_558)
);

CKINVDCx20_ASAP7_75t_R g559 ( 
.A(n_477),
.Y(n_559)
);

CKINVDCx5p33_ASAP7_75t_R g560 ( 
.A(n_453),
.Y(n_560)
);

INVx3_ASAP7_75t_L g561 ( 
.A(n_420),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_431),
.Y(n_562)
);

INVxp67_ASAP7_75t_L g563 ( 
.A(n_429),
.Y(n_563)
);

HB1xp67_ASAP7_75t_L g564 ( 
.A(n_476),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_433),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_L g566 ( 
.A(n_463),
.B(n_379),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_433),
.Y(n_567)
);

CKINVDCx20_ASAP7_75t_R g568 ( 
.A(n_486),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_476),
.Y(n_569)
);

INVx2_ASAP7_75t_SL g570 ( 
.A(n_507),
.Y(n_570)
);

INVx2_ASAP7_75t_L g571 ( 
.A(n_540),
.Y(n_571)
);

BUFx6f_ASAP7_75t_L g572 ( 
.A(n_507),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_540),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_520),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_SL g575 ( 
.A(n_537),
.B(n_468),
.Y(n_575)
);

INVx2_ASAP7_75t_L g576 ( 
.A(n_544),
.Y(n_576)
);

INVx2_ASAP7_75t_L g577 ( 
.A(n_544),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_SL g578 ( 
.A(n_546),
.B(n_466),
.Y(n_578)
);

INVx2_ASAP7_75t_L g579 ( 
.A(n_520),
.Y(n_579)
);

BUFx3_ASAP7_75t_L g580 ( 
.A(n_504),
.Y(n_580)
);

INVx2_ASAP7_75t_L g581 ( 
.A(n_531),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_531),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_534),
.Y(n_583)
);

BUFx6f_ASAP7_75t_SL g584 ( 
.A(n_504),
.Y(n_584)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_534),
.Y(n_585)
);

BUFx10_ASAP7_75t_L g586 ( 
.A(n_504),
.Y(n_586)
);

INVx3_ASAP7_75t_L g587 ( 
.A(n_561),
.Y(n_587)
);

AO21x2_ASAP7_75t_L g588 ( 
.A1(n_541),
.A2(n_481),
.B(n_482),
.Y(n_588)
);

AND2x6_ASAP7_75t_L g589 ( 
.A(n_561),
.B(n_487),
.Y(n_589)
);

INVx2_ASAP7_75t_L g590 ( 
.A(n_539),
.Y(n_590)
);

INVx2_ASAP7_75t_L g591 ( 
.A(n_539),
.Y(n_591)
);

BUFx6f_ASAP7_75t_SL g592 ( 
.A(n_509),
.Y(n_592)
);

INVx3_ASAP7_75t_L g593 ( 
.A(n_561),
.Y(n_593)
);

OAI22xp33_ASAP7_75t_L g594 ( 
.A1(n_560),
.A2(n_455),
.B1(n_490),
.B2(n_489),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_503),
.Y(n_595)
);

INVx2_ASAP7_75t_L g596 ( 
.A(n_508),
.Y(n_596)
);

INVx2_ASAP7_75t_L g597 ( 
.A(n_512),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_516),
.Y(n_598)
);

CKINVDCx6p67_ASAP7_75t_R g599 ( 
.A(n_510),
.Y(n_599)
);

INVx2_ASAP7_75t_L g600 ( 
.A(n_518),
.Y(n_600)
);

INVx2_ASAP7_75t_L g601 ( 
.A(n_526),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_SL g602 ( 
.A(n_533),
.B(n_456),
.Y(n_602)
);

INVx2_ASAP7_75t_L g603 ( 
.A(n_551),
.Y(n_603)
);

BUFx10_ASAP7_75t_L g604 ( 
.A(n_538),
.Y(n_604)
);

INVx3_ASAP7_75t_L g605 ( 
.A(n_550),
.Y(n_605)
);

INVx2_ASAP7_75t_L g606 ( 
.A(n_552),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_L g607 ( 
.A(n_517),
.B(n_445),
.Y(n_607)
);

INVxp67_ASAP7_75t_L g608 ( 
.A(n_530),
.Y(n_608)
);

BUFx3_ASAP7_75t_L g609 ( 
.A(n_599),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_SL g610 ( 
.A(n_594),
.B(n_509),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_595),
.Y(n_611)
);

INVx2_ASAP7_75t_L g612 ( 
.A(n_571),
.Y(n_612)
);

AND3x1_ASAP7_75t_L g613 ( 
.A(n_599),
.B(n_545),
.C(n_557),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_L g614 ( 
.A(n_607),
.B(n_505),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_595),
.Y(n_615)
);

INVx2_ASAP7_75t_L g616 ( 
.A(n_571),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_L g617 ( 
.A(n_607),
.B(n_575),
.Y(n_617)
);

NOR2xp33_ASAP7_75t_L g618 ( 
.A(n_578),
.B(n_554),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_SL g619 ( 
.A(n_602),
.B(n_536),
.Y(n_619)
);

NAND2xp33_ASAP7_75t_L g620 ( 
.A(n_589),
.B(n_528),
.Y(n_620)
);

INVx2_ASAP7_75t_L g621 ( 
.A(n_571),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_598),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_598),
.Y(n_623)
);

NOR2xp33_ASAP7_75t_L g624 ( 
.A(n_608),
.B(n_554),
.Y(n_624)
);

INVx3_ASAP7_75t_L g625 ( 
.A(n_586),
.Y(n_625)
);

AND2x6_ASAP7_75t_L g626 ( 
.A(n_587),
.B(n_550),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_596),
.Y(n_627)
);

INVx4_ASAP7_75t_L g628 ( 
.A(n_584),
.Y(n_628)
);

INVx2_ASAP7_75t_L g629 ( 
.A(n_573),
.Y(n_629)
);

AOI22xp33_ASAP7_75t_L g630 ( 
.A1(n_592),
.A2(n_559),
.B1(n_548),
.B2(n_555),
.Y(n_630)
);

OAI22xp33_ASAP7_75t_L g631 ( 
.A1(n_596),
.A2(n_559),
.B1(n_555),
.B2(n_557),
.Y(n_631)
);

INVx2_ASAP7_75t_L g632 ( 
.A(n_573),
.Y(n_632)
);

INVx2_ASAP7_75t_L g633 ( 
.A(n_573),
.Y(n_633)
);

AND2x6_ASAP7_75t_L g634 ( 
.A(n_587),
.B(n_550),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_596),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_597),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_L g637 ( 
.A(n_580),
.B(n_563),
.Y(n_637)
);

BUFx10_ASAP7_75t_L g638 ( 
.A(n_584),
.Y(n_638)
);

INVxp67_ASAP7_75t_SL g639 ( 
.A(n_597),
.Y(n_639)
);

INVx3_ASAP7_75t_L g640 ( 
.A(n_586),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_597),
.Y(n_641)
);

AOI22xp33_ASAP7_75t_L g642 ( 
.A1(n_592),
.A2(n_566),
.B1(n_568),
.B2(n_543),
.Y(n_642)
);

INVx2_ASAP7_75t_L g643 ( 
.A(n_576),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_600),
.Y(n_644)
);

BUFx4f_ASAP7_75t_L g645 ( 
.A(n_572),
.Y(n_645)
);

INVx6_ASAP7_75t_L g646 ( 
.A(n_586),
.Y(n_646)
);

BUFx6f_ASAP7_75t_L g647 ( 
.A(n_572),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_600),
.Y(n_648)
);

INVxp33_ASAP7_75t_L g649 ( 
.A(n_600),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_601),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_601),
.Y(n_651)
);

INVx1_ASAP7_75t_SL g652 ( 
.A(n_580),
.Y(n_652)
);

INVxp67_ASAP7_75t_L g653 ( 
.A(n_601),
.Y(n_653)
);

OR2x6_ASAP7_75t_L g654 ( 
.A(n_603),
.B(n_494),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_580),
.B(n_479),
.Y(n_655)
);

INVx1_ASAP7_75t_SL g656 ( 
.A(n_586),
.Y(n_656)
);

BUFx6f_ASAP7_75t_L g657 ( 
.A(n_572),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_L g658 ( 
.A(n_603),
.B(n_564),
.Y(n_658)
);

INVx3_ASAP7_75t_L g659 ( 
.A(n_584),
.Y(n_659)
);

INVx2_ASAP7_75t_L g660 ( 
.A(n_576),
.Y(n_660)
);

AOI22xp33_ASAP7_75t_L g661 ( 
.A1(n_592),
.A2(n_568),
.B1(n_547),
.B2(n_549),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_603),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_606),
.Y(n_663)
);

NAND2xp33_ASAP7_75t_L g664 ( 
.A(n_589),
.B(n_522),
.Y(n_664)
);

AND2x2_ASAP7_75t_L g665 ( 
.A(n_606),
.B(n_510),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_606),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_574),
.Y(n_667)
);

INVx2_ASAP7_75t_L g668 ( 
.A(n_576),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_SL g669 ( 
.A(n_587),
.B(n_519),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_574),
.Y(n_670)
);

INVx4_ASAP7_75t_SL g671 ( 
.A(n_584),
.Y(n_671)
);

BUFx3_ASAP7_75t_L g672 ( 
.A(n_572),
.Y(n_672)
);

AOI22xp33_ASAP7_75t_L g673 ( 
.A1(n_592),
.A2(n_542),
.B1(n_225),
.B2(n_219),
.Y(n_673)
);

INVx2_ASAP7_75t_L g674 ( 
.A(n_577),
.Y(n_674)
);

INVx2_ASAP7_75t_L g675 ( 
.A(n_577),
.Y(n_675)
);

CKINVDCx20_ASAP7_75t_R g676 ( 
.A(n_604),
.Y(n_676)
);

INVx4_ASAP7_75t_L g677 ( 
.A(n_572),
.Y(n_677)
);

INVx2_ASAP7_75t_L g678 ( 
.A(n_577),
.Y(n_678)
);

NOR2xp33_ASAP7_75t_L g679 ( 
.A(n_605),
.B(n_569),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_582),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_SL g681 ( 
.A(n_587),
.B(n_487),
.Y(n_681)
);

INVx2_ASAP7_75t_L g682 ( 
.A(n_579),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_582),
.Y(n_683)
);

OR2x6_ASAP7_75t_L g684 ( 
.A(n_605),
.B(n_494),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_579),
.Y(n_685)
);

AOI22xp33_ASAP7_75t_L g686 ( 
.A1(n_583),
.A2(n_396),
.B1(n_403),
.B2(n_379),
.Y(n_686)
);

INVx2_ASAP7_75t_L g687 ( 
.A(n_579),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_581),
.Y(n_688)
);

CKINVDCx11_ASAP7_75t_R g689 ( 
.A(n_604),
.Y(n_689)
);

INVx2_ASAP7_75t_SL g690 ( 
.A(n_604),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_L g691 ( 
.A(n_583),
.B(n_538),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_581),
.Y(n_692)
);

INVx8_ASAP7_75t_L g693 ( 
.A(n_572),
.Y(n_693)
);

NOR2xp33_ASAP7_75t_L g694 ( 
.A(n_605),
.B(n_535),
.Y(n_694)
);

AND2x2_ASAP7_75t_L g695 ( 
.A(n_665),
.B(n_521),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_611),
.Y(n_696)
);

NOR2xp33_ASAP7_75t_L g697 ( 
.A(n_617),
.B(n_535),
.Y(n_697)
);

INVx2_ASAP7_75t_L g698 ( 
.A(n_615),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_622),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_623),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_SL g701 ( 
.A(n_630),
.B(n_631),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_639),
.Y(n_702)
);

INVx2_ASAP7_75t_L g703 ( 
.A(n_627),
.Y(n_703)
);

NOR2xp33_ASAP7_75t_L g704 ( 
.A(n_624),
.B(n_513),
.Y(n_704)
);

INVx2_ASAP7_75t_L g705 ( 
.A(n_635),
.Y(n_705)
);

NOR2xp33_ASAP7_75t_L g706 ( 
.A(n_631),
.B(n_605),
.Y(n_706)
);

INVx2_ASAP7_75t_L g707 ( 
.A(n_636),
.Y(n_707)
);

NOR2xp33_ASAP7_75t_L g708 ( 
.A(n_624),
.B(n_513),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_639),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_641),
.Y(n_710)
);

AOI21xp5_ASAP7_75t_L g711 ( 
.A1(n_664),
.A2(n_524),
.B(n_493),
.Y(n_711)
);

CKINVDCx5p33_ASAP7_75t_R g712 ( 
.A(n_609),
.Y(n_712)
);

BUFx6f_ASAP7_75t_L g713 ( 
.A(n_609),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_644),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_SL g715 ( 
.A(n_630),
.B(n_604),
.Y(n_715)
);

NAND2x1p5_ASAP7_75t_L g716 ( 
.A(n_628),
.B(n_593),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_648),
.Y(n_717)
);

OR2x2_ASAP7_75t_L g718 ( 
.A(n_614),
.B(n_583),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_650),
.Y(n_719)
);

XOR2xp5_ASAP7_75t_L g720 ( 
.A(n_613),
.B(n_514),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_651),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_662),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_663),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_666),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_667),
.Y(n_725)
);

AND2x2_ASAP7_75t_L g726 ( 
.A(n_618),
.B(n_585),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_670),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_680),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_683),
.Y(n_729)
);

INVx3_ASAP7_75t_L g730 ( 
.A(n_638),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_653),
.Y(n_731)
);

CKINVDCx5p33_ASAP7_75t_R g732 ( 
.A(n_689),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_653),
.Y(n_733)
);

AOI22xp5_ASAP7_75t_L g734 ( 
.A1(n_618),
.A2(n_642),
.B1(n_661),
.B2(n_610),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_685),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_688),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_692),
.Y(n_737)
);

INVx2_ASAP7_75t_SL g738 ( 
.A(n_693),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_619),
.B(n_585),
.Y(n_739)
);

NOR2xp33_ASAP7_75t_L g740 ( 
.A(n_637),
.B(n_514),
.Y(n_740)
);

INVxp67_ASAP7_75t_SL g741 ( 
.A(n_658),
.Y(n_741)
);

CKINVDCx16_ASAP7_75t_R g742 ( 
.A(n_676),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_612),
.Y(n_743)
);

AND2x2_ASAP7_75t_SL g744 ( 
.A(n_620),
.B(n_527),
.Y(n_744)
);

INVx2_ASAP7_75t_L g745 ( 
.A(n_616),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_621),
.Y(n_746)
);

NOR2xp33_ASAP7_75t_L g747 ( 
.A(n_655),
.B(n_529),
.Y(n_747)
);

OAI21xp5_ASAP7_75t_L g748 ( 
.A1(n_619),
.A2(n_440),
.B(n_425),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_629),
.Y(n_749)
);

AOI21xp5_ASAP7_75t_L g750 ( 
.A1(n_669),
.A2(n_524),
.B(n_493),
.Y(n_750)
);

NOR2xp33_ASAP7_75t_L g751 ( 
.A(n_694),
.B(n_515),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_632),
.Y(n_752)
);

XOR2xp5_ASAP7_75t_L g753 ( 
.A(n_676),
.B(n_523),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_633),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_643),
.Y(n_755)
);

AND2x2_ASAP7_75t_SL g756 ( 
.A(n_642),
.B(n_527),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_660),
.Y(n_757)
);

CKINVDCx5p33_ASAP7_75t_R g758 ( 
.A(n_689),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_649),
.B(n_585),
.Y(n_759)
);

INVxp67_ASAP7_75t_SL g760 ( 
.A(n_649),
.Y(n_760)
);

INVx2_ASAP7_75t_L g761 ( 
.A(n_668),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_674),
.Y(n_762)
);

AOI21x1_ASAP7_75t_L g763 ( 
.A1(n_669),
.A2(n_610),
.B(n_681),
.Y(n_763)
);

AND2x2_ASAP7_75t_L g764 ( 
.A(n_694),
.B(n_590),
.Y(n_764)
);

AND2x2_ASAP7_75t_L g765 ( 
.A(n_652),
.B(n_590),
.Y(n_765)
);

NOR2xp33_ASAP7_75t_L g766 ( 
.A(n_673),
.B(n_532),
.Y(n_766)
);

AND2x4_ASAP7_75t_L g767 ( 
.A(n_671),
.B(n_659),
.Y(n_767)
);

INVxp67_ASAP7_75t_L g768 ( 
.A(n_679),
.Y(n_768)
);

AND2x2_ASAP7_75t_L g769 ( 
.A(n_661),
.B(n_590),
.Y(n_769)
);

XOR2xp5_ASAP7_75t_L g770 ( 
.A(n_673),
.B(n_525),
.Y(n_770)
);

NOR2xp33_ASAP7_75t_L g771 ( 
.A(n_691),
.B(n_495),
.Y(n_771)
);

NAND2xp33_ASAP7_75t_SL g772 ( 
.A(n_628),
.B(n_506),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_675),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_678),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_682),
.Y(n_775)
);

INVx2_ASAP7_75t_L g776 ( 
.A(n_687),
.Y(n_776)
);

XOR2xp5_ASAP7_75t_L g777 ( 
.A(n_659),
.B(n_511),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_654),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_654),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_654),
.Y(n_780)
);

AND2x2_ASAP7_75t_L g781 ( 
.A(n_679),
.B(n_656),
.Y(n_781)
);

INVxp67_ASAP7_75t_L g782 ( 
.A(n_672),
.Y(n_782)
);

OAI22xp5_ASAP7_75t_L g783 ( 
.A1(n_734),
.A2(n_686),
.B1(n_646),
.B2(n_645),
.Y(n_783)
);

CKINVDCx5p33_ASAP7_75t_R g784 ( 
.A(n_732),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_696),
.Y(n_785)
);

OAI21xp33_ASAP7_75t_L g786 ( 
.A1(n_701),
.A2(n_231),
.B(n_396),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_L g787 ( 
.A(n_741),
.B(n_588),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_L g788 ( 
.A(n_741),
.B(n_768),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_768),
.B(n_588),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_699),
.Y(n_790)
);

OR2x2_ASAP7_75t_L g791 ( 
.A(n_760),
.B(n_684),
.Y(n_791)
);

NOR2xp33_ASAP7_75t_L g792 ( 
.A(n_740),
.B(n_207),
.Y(n_792)
);

NAND2xp33_ASAP7_75t_L g793 ( 
.A(n_758),
.B(n_690),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_SL g794 ( 
.A(n_742),
.B(n_638),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_SL g795 ( 
.A(n_713),
.B(n_625),
.Y(n_795)
);

INVx2_ASAP7_75t_SL g796 ( 
.A(n_713),
.Y(n_796)
);

INVx2_ASAP7_75t_SL g797 ( 
.A(n_713),
.Y(n_797)
);

INVx1_ASAP7_75t_SL g798 ( 
.A(n_695),
.Y(n_798)
);

NOR2xp33_ASAP7_75t_L g799 ( 
.A(n_704),
.B(n_207),
.Y(n_799)
);

INVx2_ASAP7_75t_L g800 ( 
.A(n_698),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_SL g801 ( 
.A(n_697),
.B(n_625),
.Y(n_801)
);

INVx2_ASAP7_75t_SL g802 ( 
.A(n_712),
.Y(n_802)
);

INVx2_ASAP7_75t_L g803 ( 
.A(n_700),
.Y(n_803)
);

AND2x2_ASAP7_75t_L g804 ( 
.A(n_781),
.B(n_672),
.Y(n_804)
);

INVx2_ASAP7_75t_SL g805 ( 
.A(n_777),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_L g806 ( 
.A(n_726),
.B(n_640),
.Y(n_806)
);

NOR2xp33_ASAP7_75t_L g807 ( 
.A(n_708),
.B(n_187),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_L g808 ( 
.A(n_764),
.B(n_640),
.Y(n_808)
);

OAI22xp33_ASAP7_75t_L g809 ( 
.A1(n_715),
.A2(n_646),
.B1(n_684),
.B2(n_645),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_725),
.Y(n_810)
);

AOI22xp33_ASAP7_75t_L g811 ( 
.A1(n_706),
.A2(n_192),
.B1(n_187),
.B2(n_538),
.Y(n_811)
);

INVx2_ASAP7_75t_L g812 ( 
.A(n_727),
.Y(n_812)
);

AND2x2_ASAP7_75t_SL g813 ( 
.A(n_744),
.B(n_671),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_L g814 ( 
.A(n_697),
.B(n_684),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_L g815 ( 
.A(n_718),
.B(n_591),
.Y(n_815)
);

BUFx12f_ASAP7_75t_L g816 ( 
.A(n_738),
.Y(n_816)
);

BUFx3_ASAP7_75t_L g817 ( 
.A(n_753),
.Y(n_817)
);

AND2x2_ASAP7_75t_L g818 ( 
.A(n_760),
.B(n_647),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_L g819 ( 
.A(n_702),
.B(n_588),
.Y(n_819)
);

AO22x1_ASAP7_75t_L g820 ( 
.A1(n_751),
.A2(n_634),
.B1(n_626),
.B2(n_677),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_728),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_729),
.Y(n_822)
);

AOI22xp33_ASAP7_75t_L g823 ( 
.A1(n_706),
.A2(n_192),
.B1(n_187),
.B2(n_403),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_L g824 ( 
.A(n_709),
.B(n_588),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_SL g825 ( 
.A(n_730),
.B(n_671),
.Y(n_825)
);

OAI22xp5_ASAP7_75t_L g826 ( 
.A1(n_756),
.A2(n_686),
.B1(n_646),
.B2(n_471),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_710),
.Y(n_827)
);

BUFx6f_ASAP7_75t_L g828 ( 
.A(n_767),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_L g829 ( 
.A(n_731),
.B(n_581),
.Y(n_829)
);

AOI22xp5_ASAP7_75t_L g830 ( 
.A1(n_772),
.A2(n_192),
.B1(n_403),
.B2(n_497),
.Y(n_830)
);

INVx2_ASAP7_75t_SL g831 ( 
.A(n_730),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_L g832 ( 
.A(n_733),
.B(n_591),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_714),
.Y(n_833)
);

NOR2xp67_ASAP7_75t_L g834 ( 
.A(n_782),
.B(n_677),
.Y(n_834)
);

OR2x2_ASAP7_75t_L g835 ( 
.A(n_717),
.B(n_681),
.Y(n_835)
);

INVx2_ASAP7_75t_L g836 ( 
.A(n_703),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_L g837 ( 
.A(n_719),
.B(n_591),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_721),
.B(n_647),
.Y(n_838)
);

AOI22xp5_ASAP7_75t_L g839 ( 
.A1(n_770),
.A2(n_403),
.B1(n_502),
.B2(n_499),
.Y(n_839)
);

OAI21xp5_ASAP7_75t_L g840 ( 
.A1(n_771),
.A2(n_485),
.B(n_500),
.Y(n_840)
);

O2A1O1Ixp33_ASAP7_75t_L g841 ( 
.A1(n_766),
.A2(n_570),
.B(n_558),
.C(n_565),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_SL g842 ( 
.A(n_744),
.B(n_647),
.Y(n_842)
);

NAND2xp33_ASAP7_75t_L g843 ( 
.A(n_720),
.B(n_626),
.Y(n_843)
);

AND2x2_ASAP7_75t_L g844 ( 
.A(n_769),
.B(n_647),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_722),
.Y(n_845)
);

NOR2xp33_ASAP7_75t_L g846 ( 
.A(n_747),
.B(n_222),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_723),
.Y(n_847)
);

NOR2xp33_ASAP7_75t_L g848 ( 
.A(n_747),
.B(n_223),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_724),
.Y(n_849)
);

INVx2_ASAP7_75t_L g850 ( 
.A(n_705),
.Y(n_850)
);

INVx2_ASAP7_75t_SL g851 ( 
.A(n_767),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_L g852 ( 
.A(n_735),
.B(n_736),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_L g853 ( 
.A(n_737),
.B(n_657),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_707),
.B(n_657),
.Y(n_854)
);

NOR3xp33_ASAP7_75t_L g855 ( 
.A(n_771),
.B(n_570),
.C(n_229),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_L g856 ( 
.A(n_759),
.B(n_657),
.Y(n_856)
);

NAND3xp33_ASAP7_75t_L g857 ( 
.A(n_766),
.B(n_230),
.C(n_228),
.Y(n_857)
);

CKINVDCx5p33_ASAP7_75t_R g858 ( 
.A(n_784),
.Y(n_858)
);

AOI22xp33_ASAP7_75t_L g859 ( 
.A1(n_786),
.A2(n_756),
.B1(n_189),
.B2(n_748),
.Y(n_859)
);

HB1xp67_ASAP7_75t_L g860 ( 
.A(n_788),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_SL g861 ( 
.A(n_813),
.B(n_716),
.Y(n_861)
);

NOR2xp33_ASAP7_75t_L g862 ( 
.A(n_807),
.B(n_782),
.Y(n_862)
);

AOI22xp33_ASAP7_75t_L g863 ( 
.A1(n_855),
.A2(n_848),
.B1(n_846),
.B2(n_811),
.Y(n_863)
);

INVx3_ASAP7_75t_L g864 ( 
.A(n_828),
.Y(n_864)
);

AOI22xp5_ASAP7_75t_L g865 ( 
.A1(n_809),
.A2(n_779),
.B1(n_780),
.B2(n_778),
.Y(n_865)
);

AND2x2_ASAP7_75t_L g866 ( 
.A(n_818),
.B(n_716),
.Y(n_866)
);

O2A1O1Ixp33_ASAP7_75t_L g867 ( 
.A1(n_823),
.A2(n_739),
.B(n_750),
.C(n_748),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_788),
.B(n_739),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_785),
.Y(n_869)
);

INVx2_ASAP7_75t_SL g870 ( 
.A(n_796),
.Y(n_870)
);

AOI21xp5_ASAP7_75t_L g871 ( 
.A1(n_857),
.A2(n_711),
.B(n_750),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_790),
.Y(n_872)
);

AOI22xp33_ASAP7_75t_L g873 ( 
.A1(n_801),
.A2(n_189),
.B1(n_634),
.B2(n_626),
.Y(n_873)
);

INVx2_ASAP7_75t_L g874 ( 
.A(n_803),
.Y(n_874)
);

NOR2xp33_ASAP7_75t_SL g875 ( 
.A(n_802),
.B(n_765),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_808),
.B(n_763),
.Y(n_876)
);

BUFx3_ASAP7_75t_L g877 ( 
.A(n_816),
.Y(n_877)
);

BUFx3_ASAP7_75t_L g878 ( 
.A(n_817),
.Y(n_878)
);

AOI22xp33_ASAP7_75t_L g879 ( 
.A1(n_792),
.A2(n_189),
.B1(n_746),
.B2(n_743),
.Y(n_879)
);

AOI22xp5_ASAP7_75t_L g880 ( 
.A1(n_783),
.A2(n_843),
.B1(n_830),
.B2(n_826),
.Y(n_880)
);

NOR2x2_ASAP7_75t_L g881 ( 
.A(n_812),
.B(n_745),
.Y(n_881)
);

AOI22xp33_ASAP7_75t_L g882 ( 
.A1(n_799),
.A2(n_634),
.B1(n_626),
.B2(n_711),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_L g883 ( 
.A(n_806),
.B(n_759),
.Y(n_883)
);

NOR2xp33_ASAP7_75t_L g884 ( 
.A(n_794),
.B(n_749),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_SL g885 ( 
.A(n_828),
.B(n_761),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_810),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_L g887 ( 
.A(n_856),
.B(n_752),
.Y(n_887)
);

INVx3_ASAP7_75t_L g888 ( 
.A(n_828),
.Y(n_888)
);

INVx4_ASAP7_75t_L g889 ( 
.A(n_797),
.Y(n_889)
);

INVxp67_ASAP7_75t_L g890 ( 
.A(n_789),
.Y(n_890)
);

AND2x6_ASAP7_75t_SL g891 ( 
.A(n_814),
.B(n_754),
.Y(n_891)
);

INVx2_ASAP7_75t_L g892 ( 
.A(n_800),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_821),
.Y(n_893)
);

NAND2xp33_ASAP7_75t_L g894 ( 
.A(n_805),
.B(n_626),
.Y(n_894)
);

A2O1A1Ixp33_ASAP7_75t_L g895 ( 
.A1(n_839),
.A2(n_693),
.B(n_236),
.C(n_235),
.Y(n_895)
);

AND2x2_ASAP7_75t_SL g896 ( 
.A(n_793),
.B(n_787),
.Y(n_896)
);

INVx2_ASAP7_75t_L g897 ( 
.A(n_822),
.Y(n_897)
);

O2A1O1Ixp5_ASAP7_75t_L g898 ( 
.A1(n_820),
.A2(n_776),
.B(n_755),
.C(n_762),
.Y(n_898)
);

A2O1A1Ixp33_ASAP7_75t_L g899 ( 
.A1(n_841),
.A2(n_842),
.B(n_840),
.C(n_825),
.Y(n_899)
);

NOR2xp33_ASAP7_75t_L g900 ( 
.A(n_798),
.B(n_757),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_827),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_833),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_L g903 ( 
.A(n_836),
.B(n_773),
.Y(n_903)
);

CKINVDCx5p33_ASAP7_75t_R g904 ( 
.A(n_831),
.Y(n_904)
);

NOR2xp33_ASAP7_75t_L g905 ( 
.A(n_804),
.B(n_774),
.Y(n_905)
);

INVx2_ASAP7_75t_L g906 ( 
.A(n_850),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_L g907 ( 
.A(n_845),
.B(n_775),
.Y(n_907)
);

NOR2x1_ASAP7_75t_R g908 ( 
.A(n_795),
.B(n_281),
.Y(n_908)
);

INVx2_ASAP7_75t_L g909 ( 
.A(n_847),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_L g910 ( 
.A(n_849),
.B(n_657),
.Y(n_910)
);

AOI22xp33_ASAP7_75t_L g911 ( 
.A1(n_789),
.A2(n_500),
.B1(n_488),
.B2(n_567),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_SL g912 ( 
.A(n_851),
.B(n_693),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_L g913 ( 
.A(n_844),
.B(n_852),
.Y(n_913)
);

AOI22xp33_ASAP7_75t_L g914 ( 
.A1(n_791),
.A2(n_634),
.B1(n_400),
.B2(n_500),
.Y(n_914)
);

HB1xp67_ASAP7_75t_L g915 ( 
.A(n_819),
.Y(n_915)
);

OAI21xp5_ASAP7_75t_L g916 ( 
.A1(n_787),
.A2(n_634),
.B(n_488),
.Y(n_916)
);

INVx2_ASAP7_75t_L g917 ( 
.A(n_852),
.Y(n_917)
);

NOR2xp33_ASAP7_75t_L g918 ( 
.A(n_854),
.B(n_0),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_L g919 ( 
.A(n_815),
.B(n_1),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_L g920 ( 
.A(n_838),
.B(n_1),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_L g921 ( 
.A(n_838),
.B(n_2),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_L g922 ( 
.A(n_853),
.B(n_2),
.Y(n_922)
);

AOI22xp5_ASAP7_75t_L g923 ( 
.A1(n_834),
.A2(n_488),
.B1(n_469),
.B2(n_464),
.Y(n_923)
);

AND2x6_ASAP7_75t_SL g924 ( 
.A(n_854),
.B(n_562),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_L g925 ( 
.A(n_853),
.B(n_3),
.Y(n_925)
);

INVx2_ASAP7_75t_L g926 ( 
.A(n_835),
.Y(n_926)
);

AOI22xp5_ASAP7_75t_L g927 ( 
.A1(n_819),
.A2(n_400),
.B1(n_593),
.B2(n_589),
.Y(n_927)
);

AOI22xp5_ASAP7_75t_L g928 ( 
.A1(n_824),
.A2(n_400),
.B1(n_593),
.B2(n_589),
.Y(n_928)
);

OR2x6_ASAP7_75t_L g929 ( 
.A(n_824),
.B(n_593),
.Y(n_929)
);

INVx2_ASAP7_75t_L g930 ( 
.A(n_829),
.Y(n_930)
);

NOR2xp33_ASAP7_75t_SL g931 ( 
.A(n_829),
.B(n_527),
.Y(n_931)
);

BUFx6f_ASAP7_75t_L g932 ( 
.A(n_832),
.Y(n_932)
);

INVx1_ASAP7_75t_L g933 ( 
.A(n_837),
.Y(n_933)
);

INVx3_ASAP7_75t_L g934 ( 
.A(n_832),
.Y(n_934)
);

INVx1_ASAP7_75t_L g935 ( 
.A(n_837),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_L g936 ( 
.A(n_788),
.B(n_3),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_869),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_L g938 ( 
.A(n_860),
.B(n_890),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_872),
.Y(n_939)
);

HB1xp67_ASAP7_75t_L g940 ( 
.A(n_860),
.Y(n_940)
);

INVx3_ASAP7_75t_L g941 ( 
.A(n_889),
.Y(n_941)
);

BUFx6f_ASAP7_75t_L g942 ( 
.A(n_877),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_L g943 ( 
.A(n_876),
.B(n_4),
.Y(n_943)
);

OR2x2_ASAP7_75t_L g944 ( 
.A(n_913),
.B(n_4),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_L g945 ( 
.A(n_868),
.B(n_5),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_L g946 ( 
.A(n_926),
.B(n_5),
.Y(n_946)
);

INVx2_ASAP7_75t_L g947 ( 
.A(n_881),
.Y(n_947)
);

NOR2xp33_ASAP7_75t_L g948 ( 
.A(n_862),
.B(n_6),
.Y(n_948)
);

INVx1_ASAP7_75t_SL g949 ( 
.A(n_891),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_SL g950 ( 
.A(n_896),
.B(n_507),
.Y(n_950)
);

NOR2xp33_ASAP7_75t_L g951 ( 
.A(n_878),
.B(n_7),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_886),
.Y(n_952)
);

INVx2_ASAP7_75t_SL g953 ( 
.A(n_904),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_893),
.Y(n_954)
);

INVx1_ASAP7_75t_L g955 ( 
.A(n_901),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_L g956 ( 
.A(n_890),
.B(n_8),
.Y(n_956)
);

NAND2x1p5_ASAP7_75t_L g957 ( 
.A(n_896),
.B(n_507),
.Y(n_957)
);

INVx1_ASAP7_75t_L g958 ( 
.A(n_902),
.Y(n_958)
);

NAND3xp33_ASAP7_75t_SL g959 ( 
.A(n_863),
.B(n_880),
.C(n_879),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_L g960 ( 
.A(n_883),
.B(n_8),
.Y(n_960)
);

AOI22xp5_ASAP7_75t_L g961 ( 
.A1(n_863),
.A2(n_589),
.B1(n_400),
.B2(n_553),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_897),
.Y(n_962)
);

AND2x2_ASAP7_75t_L g963 ( 
.A(n_866),
.B(n_9),
.Y(n_963)
);

INVx1_ASAP7_75t_L g964 ( 
.A(n_909),
.Y(n_964)
);

INVx2_ASAP7_75t_L g965 ( 
.A(n_917),
.Y(n_965)
);

CKINVDCx5p33_ASAP7_75t_R g966 ( 
.A(n_858),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_874),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_SL g968 ( 
.A(n_875),
.B(n_553),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_892),
.Y(n_969)
);

AOI22xp33_ASAP7_75t_L g970 ( 
.A1(n_859),
.A2(n_882),
.B1(n_879),
.B2(n_861),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_L g971 ( 
.A(n_934),
.B(n_9),
.Y(n_971)
);

AOI22xp5_ASAP7_75t_L g972 ( 
.A1(n_859),
.A2(n_589),
.B1(n_400),
.B2(n_553),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_L g973 ( 
.A(n_934),
.B(n_11),
.Y(n_973)
);

AND2x2_ASAP7_75t_L g974 ( 
.A(n_932),
.B(n_12),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_L g975 ( 
.A(n_915),
.B(n_12),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_L g976 ( 
.A(n_932),
.B(n_933),
.Y(n_976)
);

OAI21xp33_ASAP7_75t_L g977 ( 
.A1(n_899),
.A2(n_501),
.B(n_478),
.Y(n_977)
);

OR2x6_ASAP7_75t_L g978 ( 
.A(n_871),
.B(n_929),
.Y(n_978)
);

NAND2xp5_ASAP7_75t_L g979 ( 
.A(n_932),
.B(n_13),
.Y(n_979)
);

AOI22xp33_ASAP7_75t_L g980 ( 
.A1(n_871),
.A2(n_400),
.B1(n_491),
.B2(n_391),
.Y(n_980)
);

NAND2x1p5_ASAP7_75t_L g981 ( 
.A(n_889),
.B(n_553),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_L g982 ( 
.A(n_935),
.B(n_13),
.Y(n_982)
);

AOI22xp33_ASAP7_75t_L g983 ( 
.A1(n_918),
.A2(n_491),
.B1(n_589),
.B2(n_501),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_SL g984 ( 
.A(n_865),
.B(n_424),
.Y(n_984)
);

AOI22xp33_ASAP7_75t_L g985 ( 
.A1(n_884),
.A2(n_491),
.B1(n_589),
.B2(n_424),
.Y(n_985)
);

INVx1_ASAP7_75t_L g986 ( 
.A(n_906),
.Y(n_986)
);

INVx2_ASAP7_75t_L g987 ( 
.A(n_930),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_L g988 ( 
.A(n_887),
.B(n_15),
.Y(n_988)
);

INVx1_ASAP7_75t_L g989 ( 
.A(n_907),
.Y(n_989)
);

NAND3xp33_ASAP7_75t_SL g990 ( 
.A(n_895),
.B(n_480),
.C(n_475),
.Y(n_990)
);

INVx1_ASAP7_75t_L g991 ( 
.A(n_903),
.Y(n_991)
);

AOI22xp5_ASAP7_75t_L g992 ( 
.A1(n_894),
.A2(n_428),
.B1(n_432),
.B2(n_430),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_915),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_L g994 ( 
.A(n_929),
.B(n_15),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_L g995 ( 
.A(n_905),
.B(n_16),
.Y(n_995)
);

BUFx6f_ASAP7_75t_L g996 ( 
.A(n_942),
.Y(n_996)
);

NOR2xp33_ASAP7_75t_L g997 ( 
.A(n_949),
.B(n_936),
.Y(n_997)
);

OR2x6_ASAP7_75t_L g998 ( 
.A(n_957),
.B(n_950),
.Y(n_998)
);

INVx2_ASAP7_75t_SL g999 ( 
.A(n_942),
.Y(n_999)
);

AND2x6_ASAP7_75t_L g1000 ( 
.A(n_949),
.B(n_923),
.Y(n_1000)
);

INVx2_ASAP7_75t_L g1001 ( 
.A(n_947),
.Y(n_1001)
);

AOI22xp33_ASAP7_75t_L g1002 ( 
.A1(n_959),
.A2(n_916),
.B1(n_873),
.B2(n_928),
.Y(n_1002)
);

INVx1_ASAP7_75t_L g1003 ( 
.A(n_937),
.Y(n_1003)
);

INVx3_ASAP7_75t_L g1004 ( 
.A(n_941),
.Y(n_1004)
);

INVx2_ASAP7_75t_SL g1005 ( 
.A(n_942),
.Y(n_1005)
);

NOR2xp33_ASAP7_75t_L g1006 ( 
.A(n_943),
.B(n_900),
.Y(n_1006)
);

INVx3_ASAP7_75t_L g1007 ( 
.A(n_941),
.Y(n_1007)
);

INVx1_ASAP7_75t_L g1008 ( 
.A(n_939),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_952),
.Y(n_1009)
);

INVx2_ASAP7_75t_L g1010 ( 
.A(n_954),
.Y(n_1010)
);

INVxp67_ASAP7_75t_L g1011 ( 
.A(n_975),
.Y(n_1011)
);

BUFx6f_ASAP7_75t_L g1012 ( 
.A(n_974),
.Y(n_1012)
);

INVx3_ASAP7_75t_L g1013 ( 
.A(n_981),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_L g1014 ( 
.A(n_989),
.B(n_924),
.Y(n_1014)
);

OAI22xp5_ASAP7_75t_L g1015 ( 
.A1(n_970),
.A2(n_927),
.B1(n_920),
.B2(n_925),
.Y(n_1015)
);

BUFx2_ASAP7_75t_L g1016 ( 
.A(n_957),
.Y(n_1016)
);

INVx1_ASAP7_75t_L g1017 ( 
.A(n_955),
.Y(n_1017)
);

AND2x6_ASAP7_75t_L g1018 ( 
.A(n_992),
.B(n_921),
.Y(n_1018)
);

INVx1_ASAP7_75t_L g1019 ( 
.A(n_958),
.Y(n_1019)
);

BUFx10_ASAP7_75t_L g1020 ( 
.A(n_951),
.Y(n_1020)
);

INVx3_ASAP7_75t_L g1021 ( 
.A(n_981),
.Y(n_1021)
);

AOI22xp5_ASAP7_75t_L g1022 ( 
.A1(n_977),
.A2(n_912),
.B1(n_931),
.B2(n_922),
.Y(n_1022)
);

NAND3xp33_ASAP7_75t_L g1023 ( 
.A(n_948),
.B(n_978),
.C(n_984),
.Y(n_1023)
);

O2A1O1Ixp33_ASAP7_75t_L g1024 ( 
.A1(n_956),
.A2(n_919),
.B(n_898),
.C(n_867),
.Y(n_1024)
);

INVx1_ASAP7_75t_L g1025 ( 
.A(n_962),
.Y(n_1025)
);

CKINVDCx20_ASAP7_75t_R g1026 ( 
.A(n_966),
.Y(n_1026)
);

INVx2_ASAP7_75t_L g1027 ( 
.A(n_993),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_L g1028 ( 
.A(n_991),
.B(n_929),
.Y(n_1028)
);

NOR2x1p5_ASAP7_75t_L g1029 ( 
.A(n_995),
.B(n_864),
.Y(n_1029)
);

INVx2_ASAP7_75t_L g1030 ( 
.A(n_964),
.Y(n_1030)
);

INVx1_ASAP7_75t_L g1031 ( 
.A(n_940),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_L g1032 ( 
.A(n_975),
.B(n_870),
.Y(n_1032)
);

BUFx6f_ASAP7_75t_L g1033 ( 
.A(n_979),
.Y(n_1033)
);

OR2x2_ASAP7_75t_L g1034 ( 
.A(n_938),
.B(n_976),
.Y(n_1034)
);

CKINVDCx5p33_ASAP7_75t_R g1035 ( 
.A(n_953),
.Y(n_1035)
);

INVx2_ASAP7_75t_L g1036 ( 
.A(n_965),
.Y(n_1036)
);

NAND2xp5_ASAP7_75t_L g1037 ( 
.A(n_938),
.B(n_910),
.Y(n_1037)
);

INVx1_ASAP7_75t_L g1038 ( 
.A(n_967),
.Y(n_1038)
);

INVx5_ASAP7_75t_L g1039 ( 
.A(n_978),
.Y(n_1039)
);

INVx2_ASAP7_75t_L g1040 ( 
.A(n_987),
.Y(n_1040)
);

INVx2_ASAP7_75t_SL g1041 ( 
.A(n_969),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_986),
.Y(n_1042)
);

AOI22x1_ASAP7_75t_L g1043 ( 
.A1(n_944),
.A2(n_864),
.B1(n_888),
.B2(n_908),
.Y(n_1043)
);

INVx2_ASAP7_75t_L g1044 ( 
.A(n_978),
.Y(n_1044)
);

BUFx6f_ASAP7_75t_SL g1045 ( 
.A(n_960),
.Y(n_1045)
);

INVx2_ASAP7_75t_L g1046 ( 
.A(n_971),
.Y(n_1046)
);

AND2x4_ASAP7_75t_L g1047 ( 
.A(n_968),
.B(n_888),
.Y(n_1047)
);

INVx2_ASAP7_75t_SL g1048 ( 
.A(n_963),
.Y(n_1048)
);

AOI22xp5_ASAP7_75t_L g1049 ( 
.A1(n_961),
.A2(n_885),
.B1(n_914),
.B2(n_911),
.Y(n_1049)
);

INVx2_ASAP7_75t_L g1050 ( 
.A(n_973),
.Y(n_1050)
);

NAND2xp5_ASAP7_75t_L g1051 ( 
.A(n_945),
.B(n_867),
.Y(n_1051)
);

AND2x6_ASAP7_75t_SL g1052 ( 
.A(n_946),
.B(n_16),
.Y(n_1052)
);

INVx5_ASAP7_75t_L g1053 ( 
.A(n_994),
.Y(n_1053)
);

AOI22xp5_ASAP7_75t_L g1054 ( 
.A1(n_990),
.A2(n_972),
.B1(n_994),
.B2(n_983),
.Y(n_1054)
);

INVx4_ASAP7_75t_L g1055 ( 
.A(n_982),
.Y(n_1055)
);

CKINVDCx5p33_ASAP7_75t_R g1056 ( 
.A(n_988),
.Y(n_1056)
);

INVx1_ASAP7_75t_L g1057 ( 
.A(n_980),
.Y(n_1057)
);

INVx1_ASAP7_75t_L g1058 ( 
.A(n_985),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_937),
.Y(n_1059)
);

AOI22x1_ASAP7_75t_L g1060 ( 
.A1(n_949),
.A2(n_898),
.B1(n_18),
.B2(n_19),
.Y(n_1060)
);

NAND2xp5_ASAP7_75t_L g1061 ( 
.A(n_989),
.B(n_911),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_SL g1062 ( 
.A(n_1039),
.B(n_424),
.Y(n_1062)
);

AOI21xp5_ASAP7_75t_L g1063 ( 
.A1(n_1051),
.A2(n_496),
.B(n_484),
.Y(n_1063)
);

INVx4_ASAP7_75t_L g1064 ( 
.A(n_996),
.Y(n_1064)
);

INVx2_ASAP7_75t_L g1065 ( 
.A(n_1001),
.Y(n_1065)
);

NOR2xp33_ASAP7_75t_L g1066 ( 
.A(n_1055),
.B(n_17),
.Y(n_1066)
);

INVx2_ASAP7_75t_L g1067 ( 
.A(n_1033),
.Y(n_1067)
);

O2A1O1Ixp33_ASAP7_75t_L g1068 ( 
.A1(n_1024),
.A2(n_17),
.B(n_18),
.C(n_20),
.Y(n_1068)
);

AOI21xp5_ASAP7_75t_L g1069 ( 
.A1(n_1023),
.A2(n_1060),
.B(n_1014),
.Y(n_1069)
);

OAI22xp5_ASAP7_75t_L g1070 ( 
.A1(n_1002),
.A2(n_426),
.B1(n_556),
.B2(n_438),
.Y(n_1070)
);

BUFx6f_ASAP7_75t_L g1071 ( 
.A(n_996),
.Y(n_1071)
);

AND2x2_ASAP7_75t_L g1072 ( 
.A(n_1044),
.B(n_21),
.Y(n_1072)
);

AOI21xp5_ASAP7_75t_L g1073 ( 
.A1(n_1015),
.A2(n_460),
.B(n_21),
.Y(n_1073)
);

NOR2xp33_ASAP7_75t_L g1074 ( 
.A(n_1055),
.B(n_22),
.Y(n_1074)
);

INVx1_ASAP7_75t_L g1075 ( 
.A(n_1003),
.Y(n_1075)
);

NAND2xp5_ASAP7_75t_L g1076 ( 
.A(n_1053),
.B(n_23),
.Y(n_1076)
);

OAI22xp5_ASAP7_75t_L g1077 ( 
.A1(n_1054),
.A2(n_426),
.B1(n_556),
.B2(n_438),
.Y(n_1077)
);

NAND2xp5_ASAP7_75t_L g1078 ( 
.A(n_1053),
.B(n_23),
.Y(n_1078)
);

NOR2xp67_ASAP7_75t_L g1079 ( 
.A(n_1039),
.B(n_24),
.Y(n_1079)
);

O2A1O1Ixp5_ASAP7_75t_L g1080 ( 
.A1(n_1069),
.A2(n_1061),
.B(n_997),
.C(n_1031),
.Y(n_1080)
);

OAI21x1_ASAP7_75t_L g1081 ( 
.A1(n_1065),
.A2(n_1007),
.B(n_1004),
.Y(n_1081)
);

OA22x2_ASAP7_75t_L g1082 ( 
.A1(n_1076),
.A2(n_1011),
.B1(n_999),
.B2(n_1005),
.Y(n_1082)
);

NAND2xp5_ASAP7_75t_L g1083 ( 
.A(n_1075),
.B(n_1053),
.Y(n_1083)
);

INVx2_ASAP7_75t_L g1084 ( 
.A(n_1071),
.Y(n_1084)
);

INVx2_ASAP7_75t_L g1085 ( 
.A(n_1071),
.Y(n_1085)
);

O2A1O1Ixp5_ASAP7_75t_L g1086 ( 
.A1(n_1062),
.A2(n_1028),
.B(n_1050),
.C(n_1046),
.Y(n_1086)
);

NAND2xp5_ASAP7_75t_L g1087 ( 
.A(n_1067),
.B(n_1008),
.Y(n_1087)
);

INVx1_ASAP7_75t_L g1088 ( 
.A(n_1078),
.Y(n_1088)
);

A2O1A1Ixp33_ASAP7_75t_L g1089 ( 
.A1(n_1068),
.A2(n_1039),
.B(n_1006),
.C(n_1029),
.Y(n_1089)
);

AOI21x1_ASAP7_75t_L g1090 ( 
.A1(n_1079),
.A2(n_1032),
.B(n_1016),
.Y(n_1090)
);

OAI21x1_ASAP7_75t_L g1091 ( 
.A1(n_1072),
.A2(n_1007),
.B(n_1004),
.Y(n_1091)
);

NAND2xp5_ASAP7_75t_L g1092 ( 
.A(n_1064),
.B(n_1009),
.Y(n_1092)
);

AO31x2_ASAP7_75t_L g1093 ( 
.A1(n_1064),
.A2(n_1059),
.A3(n_1019),
.B(n_1017),
.Y(n_1093)
);

AOI21xp5_ASAP7_75t_L g1094 ( 
.A1(n_1073),
.A2(n_1043),
.B(n_1057),
.Y(n_1094)
);

AOI21xp33_ASAP7_75t_L g1095 ( 
.A1(n_1066),
.A2(n_1074),
.B(n_1077),
.Y(n_1095)
);

A2O1A1Ixp33_ASAP7_75t_L g1096 ( 
.A1(n_1063),
.A2(n_1058),
.B(n_1022),
.C(n_1052),
.Y(n_1096)
);

INVx1_ASAP7_75t_L g1097 ( 
.A(n_1071),
.Y(n_1097)
);

INVx2_ASAP7_75t_L g1098 ( 
.A(n_1070),
.Y(n_1098)
);

AOI21xp5_ASAP7_75t_L g1099 ( 
.A1(n_1068),
.A2(n_1056),
.B(n_1026),
.Y(n_1099)
);

OAI21x1_ASAP7_75t_L g1100 ( 
.A1(n_1065),
.A2(n_1021),
.B(n_1013),
.Y(n_1100)
);

OAI21x1_ASAP7_75t_L g1101 ( 
.A1(n_1065),
.A2(n_1021),
.B(n_1013),
.Y(n_1101)
);

AND2x2_ASAP7_75t_L g1102 ( 
.A(n_1067),
.B(n_1033),
.Y(n_1102)
);

AOI21xp5_ASAP7_75t_L g1103 ( 
.A1(n_1068),
.A2(n_1037),
.B(n_1048),
.Y(n_1103)
);

NAND2xp5_ASAP7_75t_L g1104 ( 
.A(n_1075),
.B(n_1010),
.Y(n_1104)
);

BUFx2_ASAP7_75t_L g1105 ( 
.A(n_1082),
.Y(n_1105)
);

INVx2_ASAP7_75t_L g1106 ( 
.A(n_1093),
.Y(n_1106)
);

OAI22xp5_ASAP7_75t_L g1107 ( 
.A1(n_1096),
.A2(n_1045),
.B1(n_998),
.B2(n_1049),
.Y(n_1107)
);

BUFx2_ASAP7_75t_L g1108 ( 
.A(n_1082),
.Y(n_1108)
);

NAND2xp5_ASAP7_75t_L g1109 ( 
.A(n_1088),
.B(n_1000),
.Y(n_1109)
);

NAND2xp5_ASAP7_75t_L g1110 ( 
.A(n_1103),
.B(n_1000),
.Y(n_1110)
);

INVx2_ASAP7_75t_L g1111 ( 
.A(n_1093),
.Y(n_1111)
);

O2A1O1Ixp33_ASAP7_75t_L g1112 ( 
.A1(n_1107),
.A2(n_1080),
.B(n_1089),
.C(n_1095),
.Y(n_1112)
);

AND2x4_ASAP7_75t_L g1113 ( 
.A(n_1105),
.B(n_1102),
.Y(n_1113)
);

OAI22xp5_ASAP7_75t_L g1114 ( 
.A1(n_1112),
.A2(n_1107),
.B1(n_1110),
.B2(n_1108),
.Y(n_1114)
);

AOI21x1_ASAP7_75t_L g1115 ( 
.A1(n_1113),
.A2(n_1106),
.B(n_1111),
.Y(n_1115)
);

CKINVDCx20_ASAP7_75t_R g1116 ( 
.A(n_1114),
.Y(n_1116)
);

INVx1_ASAP7_75t_L g1117 ( 
.A(n_1115),
.Y(n_1117)
);

INVx1_ASAP7_75t_L g1118 ( 
.A(n_1115),
.Y(n_1118)
);

OAI21x1_ASAP7_75t_L g1119 ( 
.A1(n_1117),
.A2(n_1090),
.B(n_1085),
.Y(n_1119)
);

HB1xp67_ASAP7_75t_L g1120 ( 
.A(n_1118),
.Y(n_1120)
);

AO31x2_ASAP7_75t_L g1121 ( 
.A1(n_1116),
.A2(n_1109),
.A3(n_1097),
.B(n_1084),
.Y(n_1121)
);

INVx2_ASAP7_75t_L g1122 ( 
.A(n_1119),
.Y(n_1122)
);

BUFx2_ASAP7_75t_L g1123 ( 
.A(n_1121),
.Y(n_1123)
);

INVx1_ASAP7_75t_L g1124 ( 
.A(n_1123),
.Y(n_1124)
);

INVx1_ASAP7_75t_L g1125 ( 
.A(n_1122),
.Y(n_1125)
);

INVx1_ASAP7_75t_L g1126 ( 
.A(n_1124),
.Y(n_1126)
);

OA21x2_ASAP7_75t_L g1127 ( 
.A1(n_1125),
.A2(n_1120),
.B(n_1083),
.Y(n_1127)
);

INVx2_ASAP7_75t_L g1128 ( 
.A(n_1127),
.Y(n_1128)
);

OR2x2_ASAP7_75t_L g1129 ( 
.A(n_1127),
.B(n_1121),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_1129),
.Y(n_1130)
);

BUFx2_ASAP7_75t_L g1131 ( 
.A(n_1128),
.Y(n_1131)
);

INVx4_ASAP7_75t_L g1132 ( 
.A(n_1131),
.Y(n_1132)
);

AND2x2_ASAP7_75t_L g1133 ( 
.A(n_1130),
.B(n_1126),
.Y(n_1133)
);

OAI22xp5_ASAP7_75t_L g1134 ( 
.A1(n_1132),
.A2(n_1127),
.B1(n_1083),
.B2(n_1092),
.Y(n_1134)
);

INVx1_ASAP7_75t_L g1135 ( 
.A(n_1133),
.Y(n_1135)
);

INVx2_ASAP7_75t_L g1136 ( 
.A(n_1132),
.Y(n_1136)
);

AOI22xp5_ASAP7_75t_L g1137 ( 
.A1(n_1136),
.A2(n_1135),
.B1(n_1134),
.B2(n_1092),
.Y(n_1137)
);

OR2x2_ASAP7_75t_L g1138 ( 
.A(n_1134),
.B(n_1087),
.Y(n_1138)
);

INVx2_ASAP7_75t_L g1139 ( 
.A(n_1136),
.Y(n_1139)
);

BUFx2_ASAP7_75t_SL g1140 ( 
.A(n_1139),
.Y(n_1140)
);

AOI22xp33_ASAP7_75t_L g1141 ( 
.A1(n_1138),
.A2(n_1095),
.B1(n_1098),
.B2(n_996),
.Y(n_1141)
);

AND2x2_ASAP7_75t_L g1142 ( 
.A(n_1140),
.B(n_1137),
.Y(n_1142)
);

AOI22xp33_ASAP7_75t_L g1143 ( 
.A1(n_1141),
.A2(n_1094),
.B1(n_1000),
.B2(n_1087),
.Y(n_1143)
);

INVx1_ASAP7_75t_L g1144 ( 
.A(n_1142),
.Y(n_1144)
);

INVx1_ASAP7_75t_L g1145 ( 
.A(n_1143),
.Y(n_1145)
);

NAND2xp5_ASAP7_75t_L g1146 ( 
.A(n_1144),
.B(n_1099),
.Y(n_1146)
);

INVx1_ASAP7_75t_L g1147 ( 
.A(n_1145),
.Y(n_1147)
);

CKINVDCx20_ASAP7_75t_R g1148 ( 
.A(n_1147),
.Y(n_1148)
);

NAND2xp33_ASAP7_75t_SL g1149 ( 
.A(n_1146),
.B(n_1035),
.Y(n_1149)
);

INVx1_ASAP7_75t_L g1150 ( 
.A(n_1149),
.Y(n_1150)
);

OR2x2_ASAP7_75t_L g1151 ( 
.A(n_1148),
.B(n_1091),
.Y(n_1151)
);

OR2x2_ASAP7_75t_L g1152 ( 
.A(n_1151),
.B(n_1093),
.Y(n_1152)
);

INVx1_ASAP7_75t_L g1153 ( 
.A(n_1150),
.Y(n_1153)
);

INVx2_ASAP7_75t_SL g1154 ( 
.A(n_1151),
.Y(n_1154)
);

AND2x2_ASAP7_75t_L g1155 ( 
.A(n_1154),
.B(n_1081),
.Y(n_1155)
);

INVx1_ASAP7_75t_SL g1156 ( 
.A(n_1153),
.Y(n_1156)
);

NOR2xp67_ASAP7_75t_SL g1157 ( 
.A(n_1152),
.B(n_1033),
.Y(n_1157)
);

INVx1_ASAP7_75t_L g1158 ( 
.A(n_1157),
.Y(n_1158)
);

INVxp67_ASAP7_75t_L g1159 ( 
.A(n_1156),
.Y(n_1159)
);

OAI221xp5_ASAP7_75t_L g1160 ( 
.A1(n_1159),
.A2(n_1155),
.B1(n_1094),
.B2(n_26),
.C(n_27),
.Y(n_1160)
);

HB1xp67_ASAP7_75t_L g1161 ( 
.A(n_1158),
.Y(n_1161)
);

AOI211x1_ASAP7_75t_L g1162 ( 
.A1(n_1160),
.A2(n_1104),
.B(n_25),
.C(n_26),
.Y(n_1162)
);

INVx1_ASAP7_75t_L g1163 ( 
.A(n_1161),
.Y(n_1163)
);

AND2x2_ASAP7_75t_L g1164 ( 
.A(n_1163),
.B(n_1020),
.Y(n_1164)
);

OR2x2_ASAP7_75t_L g1165 ( 
.A(n_1162),
.B(n_24),
.Y(n_1165)
);

INVxp67_ASAP7_75t_L g1166 ( 
.A(n_1165),
.Y(n_1166)
);

AOI221xp5_ASAP7_75t_L g1167 ( 
.A1(n_1164),
.A2(n_28),
.B1(n_29),
.B2(n_30),
.C(n_31),
.Y(n_1167)
);

NOR2xp33_ASAP7_75t_SL g1168 ( 
.A(n_1166),
.B(n_1020),
.Y(n_1168)
);

INVx1_ASAP7_75t_L g1169 ( 
.A(n_1167),
.Y(n_1169)
);

INVx1_ASAP7_75t_SL g1170 ( 
.A(n_1169),
.Y(n_1170)
);

INVx2_ASAP7_75t_L g1171 ( 
.A(n_1168),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_1169),
.Y(n_1172)
);

OAI21xp5_ASAP7_75t_SL g1173 ( 
.A1(n_1170),
.A2(n_28),
.B(n_29),
.Y(n_1173)
);

NAND4xp75_ASAP7_75t_L g1174 ( 
.A(n_1172),
.B(n_31),
.C(n_32),
.D(n_33),
.Y(n_1174)
);

NAND2xp5_ASAP7_75t_L g1175 ( 
.A(n_1171),
.B(n_33),
.Y(n_1175)
);

NOR2x1_ASAP7_75t_L g1176 ( 
.A(n_1173),
.B(n_34),
.Y(n_1176)
);

OAI322xp33_ASAP7_75t_L g1177 ( 
.A1(n_1175),
.A2(n_34),
.A3(n_35),
.B1(n_36),
.B2(n_1104),
.C1(n_39),
.C2(n_41),
.Y(n_1177)
);

AOI221xp5_ASAP7_75t_L g1178 ( 
.A1(n_1176),
.A2(n_1177),
.B1(n_1174),
.B2(n_35),
.C(n_36),
.Y(n_1178)
);

AOI222xp33_ASAP7_75t_L g1179 ( 
.A1(n_1176),
.A2(n_1000),
.B1(n_1012),
.B2(n_1101),
.C1(n_1100),
.C2(n_45),
.Y(n_1179)
);

INVx1_ASAP7_75t_L g1180 ( 
.A(n_1178),
.Y(n_1180)
);

AOI32xp33_ASAP7_75t_L g1181 ( 
.A1(n_1179),
.A2(n_37),
.A3(n_42),
.B1(n_43),
.B2(n_44),
.Y(n_1181)
);

OAI221xp5_ASAP7_75t_SL g1182 ( 
.A1(n_1180),
.A2(n_47),
.B1(n_48),
.B2(n_49),
.C(n_51),
.Y(n_1182)
);

OAI22xp5_ASAP7_75t_L g1183 ( 
.A1(n_1181),
.A2(n_1012),
.B1(n_54),
.B2(n_55),
.Y(n_1183)
);

NOR3xp33_ASAP7_75t_L g1184 ( 
.A(n_1183),
.B(n_52),
.C(n_58),
.Y(n_1184)
);

AOI221xp5_ASAP7_75t_L g1185 ( 
.A1(n_1182),
.A2(n_1086),
.B1(n_1012),
.B2(n_62),
.C(n_66),
.Y(n_1185)
);

INVx2_ASAP7_75t_L g1186 ( 
.A(n_1184),
.Y(n_1186)
);

INVx2_ASAP7_75t_L g1187 ( 
.A(n_1185),
.Y(n_1187)
);

OAI22xp33_ASAP7_75t_SL g1188 ( 
.A1(n_1187),
.A2(n_1186),
.B1(n_60),
.B2(n_67),
.Y(n_1188)
);

AND3x4_ASAP7_75t_L g1189 ( 
.A(n_1186),
.B(n_59),
.C(n_68),
.Y(n_1189)
);

INVx1_ASAP7_75t_L g1190 ( 
.A(n_1186),
.Y(n_1190)
);

NAND3xp33_ASAP7_75t_SL g1191 ( 
.A(n_1190),
.B(n_70),
.C(n_73),
.Y(n_1191)
);

NOR3xp33_ASAP7_75t_L g1192 ( 
.A(n_1188),
.B(n_74),
.C(n_75),
.Y(n_1192)
);

NAND2xp5_ASAP7_75t_L g1193 ( 
.A(n_1189),
.B(n_76),
.Y(n_1193)
);

OR3x1_ASAP7_75t_L g1194 ( 
.A(n_1191),
.B(n_77),
.C(n_78),
.Y(n_1194)
);

NAND2xp5_ASAP7_75t_L g1195 ( 
.A(n_1193),
.B(n_80),
.Y(n_1195)
);

INVx2_ASAP7_75t_L g1196 ( 
.A(n_1194),
.Y(n_1196)
);

XOR2xp5_ASAP7_75t_L g1197 ( 
.A(n_1195),
.B(n_1192),
.Y(n_1197)
);

XNOR2xp5_ASAP7_75t_L g1198 ( 
.A(n_1197),
.B(n_81),
.Y(n_1198)
);

INVx1_ASAP7_75t_L g1199 ( 
.A(n_1196),
.Y(n_1199)
);

INVx1_ASAP7_75t_L g1200 ( 
.A(n_1199),
.Y(n_1200)
);

INVx2_ASAP7_75t_SL g1201 ( 
.A(n_1198),
.Y(n_1201)
);

HB1xp67_ASAP7_75t_L g1202 ( 
.A(n_1200),
.Y(n_1202)
);

OAI22xp5_ASAP7_75t_L g1203 ( 
.A1(n_1201),
.A2(n_83),
.B1(n_84),
.B2(n_85),
.Y(n_1203)
);

INVxp67_ASAP7_75t_SL g1204 ( 
.A(n_1202),
.Y(n_1204)
);

OAI222xp33_ASAP7_75t_L g1205 ( 
.A1(n_1203),
.A2(n_86),
.B1(n_87),
.B2(n_88),
.C1(n_89),
.C2(n_90),
.Y(n_1205)
);

OAI21xp5_ASAP7_75t_L g1206 ( 
.A1(n_1204),
.A2(n_91),
.B(n_92),
.Y(n_1206)
);

INVx1_ASAP7_75t_L g1207 ( 
.A(n_1205),
.Y(n_1207)
);

INVx2_ASAP7_75t_L g1208 ( 
.A(n_1204),
.Y(n_1208)
);

OR2x2_ASAP7_75t_L g1209 ( 
.A(n_1208),
.B(n_93),
.Y(n_1209)
);

O2A1O1Ixp33_ASAP7_75t_L g1210 ( 
.A1(n_1207),
.A2(n_94),
.B(n_95),
.C(n_99),
.Y(n_1210)
);

OAI222xp33_ASAP7_75t_L g1211 ( 
.A1(n_1206),
.A2(n_101),
.B1(n_102),
.B2(n_103),
.C1(n_104),
.C2(n_108),
.Y(n_1211)
);

AOI221x1_ASAP7_75t_L g1212 ( 
.A1(n_1210),
.A2(n_109),
.B1(n_110),
.B2(n_112),
.C(n_113),
.Y(n_1212)
);

BUFx3_ASAP7_75t_L g1213 ( 
.A(n_1209),
.Y(n_1213)
);

NAND2xp5_ASAP7_75t_L g1214 ( 
.A(n_1213),
.B(n_1211),
.Y(n_1214)
);

OAI211xp5_ASAP7_75t_SL g1215 ( 
.A1(n_1212),
.A2(n_115),
.B(n_117),
.C(n_118),
.Y(n_1215)
);

INVx2_ASAP7_75t_L g1216 ( 
.A(n_1214),
.Y(n_1216)
);

INVx1_ASAP7_75t_L g1217 ( 
.A(n_1215),
.Y(n_1217)
);

OAI22xp5_ASAP7_75t_SL g1218 ( 
.A1(n_1216),
.A2(n_121),
.B1(n_122),
.B2(n_126),
.Y(n_1218)
);

CKINVDCx20_ASAP7_75t_R g1219 ( 
.A(n_1217),
.Y(n_1219)
);

AOI21xp5_ASAP7_75t_L g1220 ( 
.A1(n_1219),
.A2(n_127),
.B(n_128),
.Y(n_1220)
);

AOI21xp33_ASAP7_75t_SL g1221 ( 
.A1(n_1218),
.A2(n_130),
.B(n_132),
.Y(n_1221)
);

HB1xp67_ASAP7_75t_L g1222 ( 
.A(n_1219),
.Y(n_1222)
);

OAI21xp5_ASAP7_75t_L g1223 ( 
.A1(n_1222),
.A2(n_135),
.B(n_136),
.Y(n_1223)
);

OAI22xp5_ASAP7_75t_L g1224 ( 
.A1(n_1221),
.A2(n_138),
.B1(n_139),
.B2(n_140),
.Y(n_1224)
);

AOI221xp5_ASAP7_75t_L g1225 ( 
.A1(n_1220),
.A2(n_141),
.B1(n_143),
.B2(n_144),
.C(n_145),
.Y(n_1225)
);

OAI22xp33_ASAP7_75t_L g1226 ( 
.A1(n_1224),
.A2(n_146),
.B1(n_147),
.B2(n_148),
.Y(n_1226)
);

AOI22xp5_ASAP7_75t_L g1227 ( 
.A1(n_1225),
.A2(n_151),
.B1(n_152),
.B2(n_153),
.Y(n_1227)
);

AOI22xp5_ASAP7_75t_L g1228 ( 
.A1(n_1223),
.A2(n_154),
.B1(n_155),
.B2(n_156),
.Y(n_1228)
);

AOI22xp5_ASAP7_75t_L g1229 ( 
.A1(n_1224),
.A2(n_157),
.B1(n_158),
.B2(n_159),
.Y(n_1229)
);

XOR2xp5_ASAP7_75t_L g1230 ( 
.A(n_1226),
.B(n_160),
.Y(n_1230)
);

OAI211xp5_ASAP7_75t_L g1231 ( 
.A1(n_1227),
.A2(n_161),
.B(n_162),
.C(n_163),
.Y(n_1231)
);

NOR2xp33_ASAP7_75t_L g1232 ( 
.A(n_1229),
.B(n_1228),
.Y(n_1232)
);

OAI21xp5_ASAP7_75t_L g1233 ( 
.A1(n_1226),
.A2(n_165),
.B(n_166),
.Y(n_1233)
);

OAI211xp5_ASAP7_75t_L g1234 ( 
.A1(n_1227),
.A2(n_167),
.B(n_169),
.C(n_170),
.Y(n_1234)
);

AOI22x1_ASAP7_75t_L g1235 ( 
.A1(n_1226),
.A2(n_173),
.B1(n_174),
.B2(n_175),
.Y(n_1235)
);

INVx1_ASAP7_75t_L g1236 ( 
.A(n_1226),
.Y(n_1236)
);

OAI21xp33_ASAP7_75t_L g1237 ( 
.A1(n_1226),
.A2(n_176),
.B(n_177),
.Y(n_1237)
);

AOI21xp5_ASAP7_75t_L g1238 ( 
.A1(n_1226),
.A2(n_178),
.B(n_401),
.Y(n_1238)
);

AO21x2_ASAP7_75t_L g1239 ( 
.A1(n_1226),
.A2(n_460),
.B(n_1047),
.Y(n_1239)
);

NAND2xp5_ASAP7_75t_SL g1240 ( 
.A(n_1226),
.B(n_498),
.Y(n_1240)
);

NAND2xp5_ASAP7_75t_L g1241 ( 
.A(n_1226),
.B(n_498),
.Y(n_1241)
);

AND2x2_ASAP7_75t_L g1242 ( 
.A(n_1236),
.B(n_498),
.Y(n_1242)
);

INVx1_ASAP7_75t_L g1243 ( 
.A(n_1232),
.Y(n_1243)
);

NAND2xp5_ASAP7_75t_L g1244 ( 
.A(n_1241),
.B(n_498),
.Y(n_1244)
);

BUFx3_ASAP7_75t_L g1245 ( 
.A(n_1240),
.Y(n_1245)
);

AND2x2_ASAP7_75t_SL g1246 ( 
.A(n_1230),
.B(n_1047),
.Y(n_1246)
);

OAI21x1_ASAP7_75t_L g1247 ( 
.A1(n_1238),
.A2(n_432),
.B(n_430),
.Y(n_1247)
);

OR2x2_ASAP7_75t_L g1248 ( 
.A(n_1233),
.B(n_473),
.Y(n_1248)
);

AOI21xp5_ASAP7_75t_L g1249 ( 
.A1(n_1237),
.A2(n_401),
.B(n_411),
.Y(n_1249)
);

CKINVDCx14_ASAP7_75t_R g1250 ( 
.A(n_1243),
.Y(n_1250)
);

AOI22xp33_ASAP7_75t_L g1251 ( 
.A1(n_1245),
.A2(n_1235),
.B1(n_1239),
.B2(n_1234),
.Y(n_1251)
);

NAND3xp33_ASAP7_75t_L g1252 ( 
.A(n_1248),
.B(n_1231),
.C(n_1239),
.Y(n_1252)
);

AOI22xp33_ASAP7_75t_SL g1253 ( 
.A1(n_1247),
.A2(n_473),
.B1(n_447),
.B2(n_443),
.Y(n_1253)
);

INVx1_ASAP7_75t_L g1254 ( 
.A(n_1244),
.Y(n_1254)
);

INVx1_ASAP7_75t_L g1255 ( 
.A(n_1249),
.Y(n_1255)
);

OAI21xp5_ASAP7_75t_L g1256 ( 
.A1(n_1250),
.A2(n_1254),
.B(n_1255),
.Y(n_1256)
);

AO21x2_ASAP7_75t_L g1257 ( 
.A1(n_1252),
.A2(n_1246),
.B(n_1242),
.Y(n_1257)
);

AO21x2_ASAP7_75t_L g1258 ( 
.A1(n_1251),
.A2(n_1042),
.B(n_1038),
.Y(n_1258)
);

OA22x2_ASAP7_75t_L g1259 ( 
.A1(n_1253),
.A2(n_1041),
.B1(n_1025),
.B2(n_1036),
.Y(n_1259)
);

AOI221xp5_ASAP7_75t_L g1260 ( 
.A1(n_1256),
.A2(n_1040),
.B1(n_1030),
.B2(n_1027),
.C(n_473),
.Y(n_1260)
);

AOI221x1_ASAP7_75t_L g1261 ( 
.A1(n_1257),
.A2(n_473),
.B1(n_458),
.B2(n_447),
.C(n_424),
.Y(n_1261)
);

AOI22xp33_ASAP7_75t_L g1262 ( 
.A1(n_1260),
.A2(n_1259),
.B1(n_1258),
.B2(n_998),
.Y(n_1262)
);

AOI21xp33_ASAP7_75t_L g1263 ( 
.A1(n_1262),
.A2(n_1261),
.B(n_1034),
.Y(n_1263)
);

AOI211xp5_ASAP7_75t_L g1264 ( 
.A1(n_1263),
.A2(n_1018),
.B(n_458),
.C(n_447),
.Y(n_1264)
);

AOI211xp5_ASAP7_75t_L g1265 ( 
.A1(n_1264),
.A2(n_1018),
.B(n_474),
.C(n_458),
.Y(n_1265)
);


endmodule