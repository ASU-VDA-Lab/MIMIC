module real_aes_3114_n_282 (n_17, n_28, n_226, n_76, n_202, n_255, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_257, n_261, n_262, n_238, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_263, n_230, n_165, n_51, n_195, n_246, n_248, n_252, n_176, n_27, n_163, n_222, n_249, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_254, n_18, n_207, n_104, n_21, n_31, n_8, n_251, n_183, n_266, n_205, n_220, n_211, n_10, n_281, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_234, n_153, n_75, n_178, n_219, n_256, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_239, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_253, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_274, n_95, n_131, n_144, n_164, n_231, n_169, n_242, n_44, n_102, n_188, n_269, n_152, n_198, n_201, n_122, n_7, n_228, n_272, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_275, n_69, n_279, n_46, n_109, n_59, n_25, n_203, n_236, n_278, n_73, n_77, n_218, n_81, n_133, n_48, n_267, n_270, n_260, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_273, n_138, n_50, n_114, n_276, n_89, n_170, n_277, n_26, n_235, n_265, n_86, n_93, n_182, n_154, n_127, n_199, n_245, n_161, n_189, n_13, n_24, n_271, n_217, n_2, n_142, n_55, n_168, n_175, n_241, n_145, n_62, n_105, n_223, n_84, n_227, n_67, n_92, n_33, n_206, n_258, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_250, n_116, n_94, n_229, n_39, n_5, n_45, n_60, n_233, n_240, n_247, n_280, n_38, n_259, n_155, n_243, n_118, n_143, n_139, n_244, n_192, n_213, n_268, n_136, n_87, n_171, n_0, n_157, n_78, n_264, n_101, n_63, n_1, n_146, n_237, n_107, n_184, n_53, n_36, n_282);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_255;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_257;
input n_261;
input n_262;
input n_238;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_263;
input n_230;
input n_165;
input n_51;
input n_195;
input n_246;
input n_248;
input n_252;
input n_176;
input n_27;
input n_163;
input n_222;
input n_249;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_254;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_251;
input n_183;
input n_266;
input n_205;
input n_220;
input n_211;
input n_10;
input n_281;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_234;
input n_153;
input n_75;
input n_178;
input n_219;
input n_256;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_239;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_253;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_274;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_242;
input n_44;
input n_102;
input n_188;
input n_269;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_272;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_275;
input n_69;
input n_279;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_236;
input n_278;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_267;
input n_270;
input n_260;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_273;
input n_138;
input n_50;
input n_114;
input n_276;
input n_89;
input n_170;
input n_277;
input n_26;
input n_235;
input n_265;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_245;
input n_161;
input n_189;
input n_13;
input n_24;
input n_271;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_241;
input n_145;
input n_62;
input n_105;
input n_223;
input n_84;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_258;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_250;
input n_116;
input n_94;
input n_229;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_240;
input n_247;
input n_280;
input n_38;
input n_259;
input n_155;
input n_243;
input n_118;
input n_143;
input n_139;
input n_244;
input n_192;
input n_213;
input n_268;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_264;
input n_101;
input n_63;
input n_1;
input n_146;
input n_237;
input n_107;
input n_184;
input n_53;
input n_36;
output n_282;
wire n_480;
wire n_476;
wire n_758;
wire n_599;
wire n_436;
wire n_887;
wire n_684;
wire n_390;
wire n_821;
wire n_830;
wire n_285;
wire n_624;
wire n_980;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_838;
wire n_933;
wire n_485;
wire n_822;
wire n_846;
wire n_750;
wire n_631;
wire n_977;
wire n_943;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_905;
wire n_518;
wire n_792;
wire n_878;
wire n_665;
wire n_667;
wire n_991;
wire n_1004;
wire n_580;
wire n_577;
wire n_469;
wire n_987;
wire n_362;
wire n_759;
wire n_979;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_900;
wire n_328;
wire n_718;
wire n_318;
wire n_841;
wire n_355;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_329;
wire n_766;
wire n_852;
wire n_974;
wire n_857;
wire n_919;
wire n_461;
wire n_908;
wire n_571;
wire n_376;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_894;
wire n_923;
wire n_952;
wire n_429;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_460;
wire n_937;
wire n_989;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_963;
wire n_865;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_884;
wire n_560;
wire n_660;
wire n_814;
wire n_944;
wire n_886;
wire n_594;
wire n_856;
wire n_983;
wire n_767;
wire n_696;
wire n_889;
wire n_955;
wire n_975;
wire n_704;
wire n_941;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_932;
wire n_399;
wire n_948;
wire n_700;
wire n_958;
wire n_677;
wire n_378;
wire n_591;
wire n_775;
wire n_763;
wire n_870;
wire n_961;
wire n_489;
wire n_427;
wire n_678;
wire n_548;
wire n_415;
wire n_572;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_625;
wire n_953;
wire n_462;
wire n_289;
wire n_615;
wire n_990;
wire n_550;
wire n_966;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_883;
wire n_478;
wire n_356;
wire n_918;
wire n_584;
wire n_896;
wire n_408;
wire n_553;
wire n_578;
wire n_994;
wire n_372;
wire n_528;
wire n_495;
wire n_892;
wire n_370;
wire n_384;
wire n_744;
wire n_938;
wire n_352;
wire n_935;
wire n_824;
wire n_951;
wire n_467;
wire n_875;
wire n_327;
wire n_992;
wire n_774;
wire n_813;
wire n_791;
wire n_981;
wire n_559;
wire n_466;
wire n_636;
wire n_872;
wire n_976;
wire n_906;
wire n_477;
wire n_515;
wire n_984;
wire n_680;
wire n_595;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_904;
wire n_840;
wire n_570;
wire n_675;
wire n_931;
wire n_920;
wire n_530;
wire n_835;
wire n_535;
wire n_732;
wire n_834;
wire n_882;
wire n_784;
wire n_496;
wire n_693;
wire n_962;
wire n_468;
wire n_746;
wire n_284;
wire n_656;
wire n_316;
wire n_532;
wire n_755;
wire n_409;
wire n_781;
wire n_748;
wire n_860;
wire n_996;
wire n_523;
wire n_298;
wire n_909;
wire n_439;
wire n_576;
wire n_924;
wire n_956;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_874;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_455;
wire n_504;
wire n_725;
wire n_973;
wire n_310;
wire n_671;
wire n_960;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_903;
wire n_454;
wire n_812;
wire n_782;
wire n_443;
wire n_565;
wire n_817;
wire n_760;
wire n_608;
wire n_925;
wire n_534;
wire n_708;
wire n_457;
wire n_345;
wire n_304;
wire n_885;
wire n_950;
wire n_381;
wire n_993;
wire n_493;
wire n_311;
wire n_324;
wire n_664;
wire n_367;
wire n_819;
wire n_737;
wire n_581;
wire n_610;
wire n_936;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_940;
wire n_722;
wire n_745;
wire n_867;
wire n_339;
wire n_398;
wire n_688;
wire n_425;
wire n_609;
wire n_879;
wire n_331;
wire n_363;
wire n_417;
wire n_754;
wire n_607;
wire n_449;
wire n_1006;
wire n_323;
wire n_690;
wire n_629;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_901;
wire n_561;
wire n_970;
wire n_947;
wire n_876;
wire n_437;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_527;
wire n_434;
wire n_505;
wire n_502;
wire n_769;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_672;
wire n_567;
wire n_916;
wire n_406;
wire n_426;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_658;
wire n_676;
wire n_986;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_880;
wire n_1008;
wire n_807;
wire n_286;
wire n_416;
wire n_790;
wire n_895;
wire n_832;
wire n_410;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_913;
wire n_999;
wire n_619;
wire n_391;
wire n_360;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_361;
wire n_917;
wire n_632;
wire n_768;
wire n_412;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_985;
wire n_777;
wire n_501;
wire n_488;
wire n_910;
wire n_642;
wire n_613;
wire n_869;
wire n_387;
wire n_957;
wire n_995;
wire n_296;
wire n_702;
wire n_954;
wire n_969;
wire n_912;
wire n_1009;
wire n_1007;
wire n_302;
wire n_464;
wire n_351;
wire n_945;
wire n_604;
wire n_734;
wire n_898;
wire n_848;
wire n_392;
wire n_562;
wire n_288;
wire n_713;
wire n_404;
wire n_598;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_303;
wire n_569;
wire n_997;
wire n_563;
wire n_785;
wire n_891;
wire n_430;
wire n_568;
wire n_413;
wire n_471;
wire n_902;
wire n_853;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_699;
wire n_533;
wire n_1000;
wire n_1003;
wire n_366;
wire n_346;
wire n_727;
wire n_397;
wire n_293;
wire n_358;
wire n_385;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_536;
wire n_914;
wire n_707;
wire n_622;
wire n_470;
wire n_915;
wire n_851;
wire n_1002;
wire n_934;
wire n_494;
wire n_1001;
wire n_711;
wire n_864;
wire n_377;
wire n_927;
wire n_965;
wire n_723;
wire n_662;
wire n_295;
wire n_382;
wire n_845;
wire n_850;
wire n_720;
wire n_354;
wire n_972;
wire n_435;
wire n_511;
wire n_484;
wire n_326;
wire n_893;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_930;
wire n_411;
wire n_697;
wire n_291;
wire n_978;
wire n_847;
wire n_907;
wire n_779;
wire n_498;
wire n_481;
wire n_691;
wire n_765;
wire n_826;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_1005;
wire n_939;
wire n_487;
wire n_831;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_928;
wire n_899;
wire n_692;
wire n_544;
wire n_789;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_827;
wire n_809;
wire n_482;
wire n_633;
wire n_679;
wire n_520;
wire n_922;
wire n_926;
wire n_942;
wire n_472;
wire n_971;
wire n_866;
wire n_452;
wire n_787;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_959;
wire n_946;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_858;
wire n_873;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_753;
wire n_283;
wire n_314;
wire n_741;
wire n_623;
wire n_721;
wire n_446;
wire n_681;
wire n_982;
wire n_359;
wire n_717;
wire n_456;
wire n_312;
wire n_712;
wire n_433;
wire n_516;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_524;
wire n_861;
wire n_705;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_541;
wire n_839;
wire n_639;
wire n_546;
wire n_587;
wire n_811;
wire n_459;
wire n_558;
wire n_863;
wire n_998;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_836;
wire n_888;
wire n_793;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_929;
wire n_686;
wire n_776;
wire n_803;
wire n_890;
wire n_543;
wire n_497;
wire n_514;
wire n_949;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_911;
wire n_772;
wire n_450;
wire n_788;
wire n_441;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_967;
wire n_837;
wire n_871;
wire n_474;
wire n_829;
wire n_988;
wire n_921;
wire n_375;
wire n_597;
wire n_640;
wire n_340;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_729;
wire n_687;
wire n_844;
wire n_968;
wire n_650;
wire n_646;
wire n_710;
wire n_743;
wire n_393;
wire n_294;
wire n_652;
wire n_703;
wire n_823;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_854;
wire n_424;
wire n_877;
wire n_802;
wire n_868;
wire n_574;
wire n_337;
wire n_842;
wire n_849;
wire n_475;
wire n_554;
wire n_897;
wire n_855;
wire n_798;
wire n_668;
wire n_797;
wire n_862;
AOI22xp33_ASAP7_75t_L g625 ( .A1(n_0), .A2(n_254), .B1(n_420), .B2(n_421), .Y(n_625) );
AO22x2_ASAP7_75t_L g606 ( .A1(n_1), .A2(n_607), .B1(n_627), .B2(n_628), .Y(n_606) );
INVxp67_ASAP7_75t_SL g627 ( .A(n_1), .Y(n_627) );
AOI22xp5_ASAP7_75t_L g752 ( .A1(n_1), .A2(n_62), .B1(n_753), .B2(n_754), .Y(n_752) );
AOI22xp33_ASAP7_75t_L g647 ( .A1(n_2), .A2(n_71), .B1(n_455), .B2(n_509), .Y(n_647) );
HB1xp67_ASAP7_75t_L g293 ( .A(n_3), .Y(n_293) );
AND2x4_ASAP7_75t_L g716 ( .A(n_3), .B(n_274), .Y(n_716) );
AND2x4_ASAP7_75t_L g721 ( .A(n_3), .B(n_722), .Y(n_721) );
AOI22xp33_ASAP7_75t_L g654 ( .A1(n_4), .A2(n_25), .B1(n_368), .B2(n_388), .Y(n_654) );
INVx1_ASAP7_75t_L g702 ( .A(n_5), .Y(n_702) );
AOI22xp33_ASAP7_75t_L g596 ( .A1(n_6), .A2(n_128), .B1(n_424), .B2(n_568), .Y(n_596) );
AOI22xp33_ASAP7_75t_L g500 ( .A1(n_7), .A2(n_187), .B1(n_388), .B2(n_501), .Y(n_500) );
AOI22xp33_ASAP7_75t_L g544 ( .A1(n_8), .A2(n_244), .B1(n_503), .B2(n_504), .Y(n_544) );
AOI22xp33_ASAP7_75t_L g655 ( .A1(n_9), .A2(n_49), .B1(n_373), .B2(n_656), .Y(n_655) );
AOI22xp33_ASAP7_75t_L g624 ( .A1(n_10), .A2(n_15), .B1(n_484), .B2(n_485), .Y(n_624) );
AOI22xp33_ASAP7_75t_L g684 ( .A1(n_11), .A2(n_104), .B1(n_420), .B2(n_421), .Y(n_684) );
AOI22xp5_ASAP7_75t_L g538 ( .A1(n_12), .A2(n_16), .B1(n_380), .B2(n_539), .Y(n_538) );
AOI22xp33_ASAP7_75t_L g648 ( .A1(n_13), .A2(n_224), .B1(n_380), .B2(n_382), .Y(n_648) );
AOI22xp33_ASAP7_75t_L g689 ( .A1(n_14), .A2(n_86), .B1(n_454), .B2(n_690), .Y(n_689) );
AOI22xp33_ASAP7_75t_L g649 ( .A1(n_17), .A2(n_93), .B1(n_373), .B2(n_543), .Y(n_649) );
AOI22xp33_ASAP7_75t_L g483 ( .A1(n_18), .A2(n_133), .B1(n_484), .B2(n_485), .Y(n_483) );
INVx1_ASAP7_75t_L g525 ( .A(n_19), .Y(n_525) );
AOI22xp5_ASAP7_75t_L g581 ( .A1(n_20), .A2(n_228), .B1(n_458), .B2(n_582), .Y(n_581) );
AOI22xp5_ASAP7_75t_L g749 ( .A1(n_21), .A2(n_92), .B1(n_725), .B2(n_750), .Y(n_749) );
AOI22xp33_ASAP7_75t_L g948 ( .A1(n_22), .A2(n_146), .B1(n_463), .B2(n_949), .Y(n_948) );
CKINVDCx20_ASAP7_75t_R g440 ( .A(n_23), .Y(n_440) );
AOI22xp33_ASAP7_75t_L g664 ( .A1(n_24), .A2(n_131), .B1(n_306), .B2(n_345), .Y(n_664) );
INVx1_ASAP7_75t_L g743 ( .A(n_26), .Y(n_743) );
AOI221xp5_ASAP7_75t_L g697 ( .A1(n_27), .A2(n_34), .B1(n_391), .B2(n_698), .C(n_700), .Y(n_697) );
INVx1_ASAP7_75t_L g341 ( .A(n_28), .Y(n_341) );
AOI22xp33_ASAP7_75t_L g506 ( .A1(n_29), .A2(n_159), .B1(n_380), .B2(n_507), .Y(n_506) );
INVx1_ASAP7_75t_L g445 ( .A(n_30), .Y(n_445) );
AOI22xp33_ASAP7_75t_L g461 ( .A1(n_31), .A2(n_115), .B1(n_462), .B2(n_463), .Y(n_461) );
AOI21x1_ASAP7_75t_L g518 ( .A1(n_32), .A2(n_519), .B(n_524), .Y(n_518) );
AOI21xp5_ASAP7_75t_L g573 ( .A1(n_33), .A2(n_431), .B(n_574), .Y(n_573) );
AOI22xp33_ASAP7_75t_L g712 ( .A1(n_35), .A2(n_91), .B1(n_713), .B2(n_717), .Y(n_712) );
AOI22xp33_ASAP7_75t_L g430 ( .A1(n_36), .A2(n_149), .B1(n_431), .B2(n_432), .Y(n_430) );
AOI22xp33_ASAP7_75t_L g666 ( .A1(n_37), .A2(n_231), .B1(n_527), .B2(n_667), .Y(n_666) );
INVx1_ASAP7_75t_SL g827 ( .A(n_38), .Y(n_827) );
XNOR2x1_ASAP7_75t_L g301 ( .A(n_39), .B(n_302), .Y(n_301) );
AOI22xp33_ASAP7_75t_L g979 ( .A1(n_40), .A2(n_85), .B1(n_503), .B2(n_980), .Y(n_979) );
INVx1_ASAP7_75t_L g641 ( .A(n_41), .Y(n_641) );
NOR2xp33_ASAP7_75t_L g291 ( .A(n_42), .B(n_210), .Y(n_291) );
INVx1_ASAP7_75t_L g317 ( .A(n_42), .Y(n_317) );
INVxp67_ASAP7_75t_L g358 ( .A(n_42), .Y(n_358) );
AOI22xp33_ASAP7_75t_L g688 ( .A1(n_43), .A2(n_168), .B1(n_373), .B2(n_568), .Y(n_688) );
INVx1_ASAP7_75t_L g593 ( .A(n_44), .Y(n_593) );
AOI22xp5_ASAP7_75t_L g695 ( .A1(n_45), .A2(n_95), .B1(n_330), .B2(n_458), .Y(n_695) );
AOI22xp33_ASAP7_75t_L g758 ( .A1(n_46), .A2(n_99), .B1(n_720), .B2(n_732), .Y(n_758) );
AOI22xp33_ASAP7_75t_L g945 ( .A1(n_47), .A2(n_66), .B1(n_509), .B2(n_543), .Y(n_945) );
AOI22xp33_ASAP7_75t_L g542 ( .A1(n_48), .A2(n_111), .B1(n_509), .B2(n_543), .Y(n_542) );
AOI22xp33_ASAP7_75t_L g665 ( .A1(n_50), .A2(n_166), .B1(n_391), .B2(n_463), .Y(n_665) );
AOI22xp5_ASAP7_75t_L g427 ( .A1(n_51), .A2(n_82), .B1(n_428), .B2(n_429), .Y(n_427) );
XNOR2x1_ASAP7_75t_L g562 ( .A(n_52), .B(n_563), .Y(n_562) );
NAND2xp5_ASAP7_75t_SL g313 ( .A(n_53), .B(n_312), .Y(n_313) );
AOI22xp33_ASAP7_75t_L g588 ( .A1(n_54), .A2(n_125), .B1(n_330), .B2(n_578), .Y(n_588) );
AOI22xp33_ASAP7_75t_L g950 ( .A1(n_55), .A2(n_117), .B1(n_951), .B2(n_953), .Y(n_950) );
AOI21xp33_ASAP7_75t_SL g609 ( .A1(n_56), .A2(n_476), .B(n_610), .Y(n_609) );
AOI22xp33_ASAP7_75t_L g657 ( .A1(n_57), .A2(n_260), .B1(n_382), .B2(n_658), .Y(n_657) );
AOI22xp33_ASAP7_75t_L g660 ( .A1(n_58), .A2(n_127), .B1(n_361), .B2(n_468), .Y(n_660) );
INVx1_ASAP7_75t_L g417 ( .A(n_59), .Y(n_417) );
INVx1_ASAP7_75t_L g493 ( .A(n_60), .Y(n_493) );
AOI22xp33_ASAP7_75t_L g676 ( .A1(n_61), .A2(n_265), .B1(n_432), .B2(n_435), .Y(n_676) );
AOI22xp33_ASAP7_75t_L g728 ( .A1(n_63), .A2(n_165), .B1(n_729), .B2(n_730), .Y(n_728) );
CKINVDCx20_ASAP7_75t_R g778 ( .A(n_64), .Y(n_778) );
AOI22xp33_ASAP7_75t_L g569 ( .A1(n_65), .A2(n_234), .B1(n_361), .B2(n_375), .Y(n_569) );
BUFx2_ASAP7_75t_L g615 ( .A(n_67), .Y(n_615) );
INVxp67_ASAP7_75t_R g745 ( .A(n_68), .Y(n_745) );
XNOR2x1_ASAP7_75t_L g585 ( .A(n_69), .B(n_586), .Y(n_585) );
AOI22xp33_ASAP7_75t_L g682 ( .A1(n_70), .A2(n_110), .B1(n_484), .B2(n_485), .Y(n_682) );
INVx1_ASAP7_75t_L g701 ( .A(n_72), .Y(n_701) );
INVx2_ASAP7_75t_L g288 ( .A(n_73), .Y(n_288) );
INVx1_ASAP7_75t_L g983 ( .A(n_74), .Y(n_983) );
INVx1_ASAP7_75t_L g715 ( .A(n_75), .Y(n_715) );
AND2x4_ASAP7_75t_L g718 ( .A(n_75), .B(n_288), .Y(n_718) );
INVx1_ASAP7_75t_SL g751 ( .A(n_75), .Y(n_751) );
OAI22xp5_ASAP7_75t_L g971 ( .A1(n_76), .A2(n_972), .B1(n_973), .B2(n_1004), .Y(n_971) );
CKINVDCx5p33_ASAP7_75t_R g972 ( .A(n_76), .Y(n_972) );
AOI22xp33_ASAP7_75t_L g475 ( .A1(n_77), .A2(n_248), .B1(n_330), .B2(n_476), .Y(n_475) );
INVx1_ASAP7_75t_L g985 ( .A(n_78), .Y(n_985) );
AOI22xp33_ASAP7_75t_L g635 ( .A1(n_79), .A2(n_164), .B1(n_330), .B2(n_636), .Y(n_635) );
AOI22xp5_ASAP7_75t_L g422 ( .A1(n_80), .A2(n_190), .B1(n_423), .B2(n_424), .Y(n_422) );
AOI22xp33_ASAP7_75t_L g991 ( .A1(n_81), .A2(n_249), .B1(n_992), .B2(n_994), .Y(n_991) );
NAND2xp5_ASAP7_75t_L g555 ( .A(n_83), .B(n_556), .Y(n_555) );
AOI22xp33_ASAP7_75t_L g598 ( .A1(n_84), .A2(n_174), .B1(n_375), .B2(n_454), .Y(n_598) );
AOI22xp5_ASAP7_75t_L g761 ( .A1(n_87), .A2(n_201), .B1(n_725), .B2(n_750), .Y(n_761) );
AOI22xp33_ASAP7_75t_L g508 ( .A1(n_88), .A2(n_242), .B1(n_509), .B2(n_510), .Y(n_508) );
AOI22xp33_ASAP7_75t_SL g545 ( .A1(n_89), .A2(n_258), .B1(n_388), .B2(n_455), .Y(n_545) );
BUFx6f_ASAP7_75t_L g312 ( .A(n_90), .Y(n_312) );
AOI22xp33_ASAP7_75t_L g683 ( .A1(n_94), .A2(n_212), .B1(n_437), .B2(n_438), .Y(n_683) );
INVx1_ASAP7_75t_L g398 ( .A(n_96), .Y(n_398) );
INVx1_ASAP7_75t_L g488 ( .A(n_97), .Y(n_488) );
AOI21xp5_ASAP7_75t_L g637 ( .A1(n_98), .A2(n_638), .B(n_640), .Y(n_637) );
CKINVDCx16_ASAP7_75t_R g741 ( .A(n_100), .Y(n_741) );
AOI22xp33_ASAP7_75t_L g719 ( .A1(n_101), .A2(n_170), .B1(n_720), .B2(n_723), .Y(n_719) );
AOI22xp5_ASAP7_75t_L g552 ( .A1(n_102), .A2(n_223), .B1(n_463), .B2(n_553), .Y(n_552) );
AOI22xp33_ASAP7_75t_L g632 ( .A1(n_103), .A2(n_158), .B1(n_458), .B2(n_633), .Y(n_632) );
AOI22xp33_ASAP7_75t_L g512 ( .A1(n_105), .A2(n_281), .B1(n_345), .B2(n_513), .Y(n_512) );
INVx1_ASAP7_75t_L g323 ( .A(n_106), .Y(n_323) );
NAND2xp5_ASAP7_75t_L g355 ( .A(n_106), .B(n_209), .Y(n_355) );
AOI22xp5_ASAP7_75t_L g693 ( .A1(n_107), .A2(n_157), .B1(n_388), .B2(n_501), .Y(n_693) );
AOI22xp33_ASAP7_75t_L g565 ( .A1(n_108), .A2(n_182), .B1(n_451), .B2(n_501), .Y(n_565) );
AOI22xp33_ASAP7_75t_L g589 ( .A1(n_109), .A2(n_178), .B1(n_306), .B2(n_582), .Y(n_589) );
AOI21xp5_ASAP7_75t_L g955 ( .A1(n_112), .A2(n_956), .B(n_958), .Y(n_955) );
AOI22xp33_ASAP7_75t_L g675 ( .A1(n_113), .A2(n_225), .B1(n_431), .B2(n_434), .Y(n_675) );
AOI22xp33_ASAP7_75t_L g942 ( .A1(n_114), .A2(n_202), .B1(n_388), .B2(n_455), .Y(n_942) );
INVx1_ASAP7_75t_L g773 ( .A(n_116), .Y(n_773) );
AOI22xp33_ASAP7_75t_L g757 ( .A1(n_118), .A2(n_171), .B1(n_713), .B2(n_730), .Y(n_757) );
AOI22xp33_ASAP7_75t_L g557 ( .A1(n_119), .A2(n_186), .B1(n_558), .B2(n_559), .Y(n_557) );
INVx1_ASAP7_75t_L g1001 ( .A(n_120), .Y(n_1001) );
INVx1_ASAP7_75t_L g535 ( .A(n_121), .Y(n_535) );
AOI22xp33_ASAP7_75t_L g646 ( .A1(n_122), .A2(n_216), .B1(n_388), .B2(n_504), .Y(n_646) );
INVx1_ASAP7_75t_L g988 ( .A(n_123), .Y(n_988) );
AOI22xp33_ASAP7_75t_L g502 ( .A1(n_124), .A2(n_163), .B1(n_503), .B2(n_504), .Y(n_502) );
AOI22xp33_ASAP7_75t_L g623 ( .A1(n_126), .A2(n_276), .B1(n_428), .B2(n_429), .Y(n_623) );
AOI22xp5_ASAP7_75t_L g995 ( .A1(n_129), .A2(n_238), .B1(n_996), .B2(n_998), .Y(n_995) );
NAND2xp5_ASAP7_75t_L g594 ( .A(n_130), .B(n_580), .Y(n_594) );
INVx1_ASAP7_75t_L g611 ( .A(n_132), .Y(n_611) );
AOI22xp33_ASAP7_75t_L g829 ( .A1(n_134), .A2(n_177), .B1(n_717), .B2(n_729), .Y(n_829) );
AOI22xp33_ASAP7_75t_L g486 ( .A1(n_135), .A2(n_257), .B1(n_420), .B2(n_421), .Y(n_486) );
AOI22xp5_ASAP7_75t_L g480 ( .A1(n_136), .A2(n_245), .B1(n_437), .B2(n_438), .Y(n_480) );
INVx1_ASAP7_75t_L g343 ( .A(n_137), .Y(n_343) );
AOI22xp33_ASAP7_75t_L g450 ( .A1(n_138), .A2(n_192), .B1(n_385), .B2(n_451), .Y(n_450) );
INVx1_ASAP7_75t_L g961 ( .A(n_139), .Y(n_961) );
AOI22xp33_ASAP7_75t_L g566 ( .A1(n_140), .A2(n_169), .B1(n_567), .B2(n_568), .Y(n_566) );
XOR2x2_ASAP7_75t_L g409 ( .A(n_141), .B(n_410), .Y(n_409) );
AOI22xp33_ASAP7_75t_SL g621 ( .A1(n_142), .A2(n_241), .B1(n_432), .B2(n_578), .Y(n_621) );
AOI21xp33_ASAP7_75t_L g590 ( .A1(n_143), .A2(n_591), .B(n_592), .Y(n_590) );
AOI22xp33_ASAP7_75t_L g457 ( .A1(n_144), .A2(n_147), .B1(n_458), .B2(n_459), .Y(n_457) );
AOI22xp33_ASAP7_75t_L g599 ( .A1(n_145), .A2(n_155), .B1(n_451), .B2(n_600), .Y(n_599) );
AOI22xp5_ASAP7_75t_L g597 ( .A1(n_148), .A2(n_214), .B1(n_382), .B2(n_466), .Y(n_597) );
AOI22xp33_ASAP7_75t_L g372 ( .A1(n_150), .A2(n_152), .B1(n_373), .B2(n_375), .Y(n_372) );
AOI22xp5_ASAP7_75t_L g976 ( .A1(n_151), .A2(n_243), .B1(n_504), .B2(n_977), .Y(n_976) );
AOI22xp5_ASAP7_75t_L g477 ( .A1(n_153), .A2(n_184), .B1(n_306), .B2(n_478), .Y(n_477) );
AOI22xp33_ASAP7_75t_L g577 ( .A1(n_154), .A2(n_196), .B1(n_330), .B2(n_578), .Y(n_577) );
AOI22xp5_ASAP7_75t_L g762 ( .A1(n_156), .A2(n_252), .B1(n_753), .B2(n_754), .Y(n_762) );
INVx1_ASAP7_75t_L g575 ( .A(n_160), .Y(n_575) );
INVx1_ASAP7_75t_L g774 ( .A(n_161), .Y(n_774) );
INVx1_ASAP7_75t_L g776 ( .A(n_162), .Y(n_776) );
INVx1_ASAP7_75t_L g987 ( .A(n_167), .Y(n_987) );
INVxp67_ASAP7_75t_SL g938 ( .A(n_170), .Y(n_938) );
AOI22xp33_ASAP7_75t_L g970 ( .A1(n_170), .A2(n_971), .B1(n_1005), .B2(n_1007), .Y(n_970) );
AOI22xp33_ASAP7_75t_L g360 ( .A1(n_172), .A2(n_219), .B1(n_361), .B2(n_368), .Y(n_360) );
AOI22xp33_ASAP7_75t_L g570 ( .A1(n_173), .A2(n_262), .B1(n_466), .B2(n_571), .Y(n_570) );
INVx1_ASAP7_75t_L g671 ( .A(n_175), .Y(n_671) );
NAND2xp5_ASAP7_75t_L g962 ( .A(n_176), .B(n_963), .Y(n_962) );
XOR2xp5_ASAP7_75t_L g629 ( .A(n_177), .B(n_630), .Y(n_629) );
AOI22xp5_ASAP7_75t_L g453 ( .A1(n_179), .A2(n_251), .B1(n_454), .B2(n_455), .Y(n_453) );
AOI22xp33_ASAP7_75t_L g943 ( .A1(n_180), .A2(n_264), .B1(n_503), .B2(n_656), .Y(n_943) );
OA22x2_ASAP7_75t_L g327 ( .A1(n_181), .A2(n_210), .B1(n_312), .B2(n_326), .Y(n_327) );
INVx1_ASAP7_75t_L g336 ( .A(n_181), .Y(n_336) );
AOI22xp33_ASAP7_75t_L g384 ( .A1(n_183), .A2(n_278), .B1(n_385), .B2(n_388), .Y(n_384) );
AOI22xp5_ASAP7_75t_L g692 ( .A1(n_185), .A2(n_236), .B1(n_382), .B2(n_466), .Y(n_692) );
AOI22xp33_ASAP7_75t_L g436 ( .A1(n_188), .A2(n_191), .B1(n_437), .B2(n_438), .Y(n_436) );
INVx1_ASAP7_75t_SL g668 ( .A(n_189), .Y(n_668) );
AOI22xp33_ASAP7_75t_L g467 ( .A1(n_193), .A2(n_267), .B1(n_373), .B2(n_468), .Y(n_467) );
AOI22xp5_ASAP7_75t_L g419 ( .A1(n_194), .A2(n_261), .B1(n_420), .B2(n_421), .Y(n_419) );
AOI22xp33_ASAP7_75t_L g515 ( .A1(n_195), .A2(n_272), .B1(n_391), .B2(n_516), .Y(n_515) );
AOI22xp5_ASAP7_75t_L g481 ( .A1(n_197), .A2(n_208), .B1(n_428), .B2(n_429), .Y(n_481) );
XOR2x2_ASAP7_75t_L g497 ( .A(n_198), .B(n_498), .Y(n_497) );
AOI22xp33_ASAP7_75t_L g433 ( .A1(n_199), .A2(n_230), .B1(n_434), .B2(n_435), .Y(n_433) );
AOI22xp33_ASAP7_75t_L g696 ( .A1(n_200), .A2(n_237), .B1(n_350), .B2(n_591), .Y(n_696) );
AOI22xp33_ASAP7_75t_L g944 ( .A1(n_203), .A2(n_255), .B1(n_380), .B2(n_539), .Y(n_944) );
INVx1_ASAP7_75t_L g495 ( .A(n_204), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g642 ( .A(n_205), .B(n_643), .Y(n_642) );
BUFx2_ASAP7_75t_L g619 ( .A(n_206), .Y(n_619) );
AOI22xp33_ASAP7_75t_L g626 ( .A1(n_207), .A2(n_240), .B1(n_437), .B2(n_438), .Y(n_626) );
INVx1_ASAP7_75t_L g319 ( .A(n_209), .Y(n_319) );
NAND2xp5_ASAP7_75t_L g406 ( .A(n_209), .B(n_334), .Y(n_406) );
OAI21xp33_ASAP7_75t_L g337 ( .A1(n_210), .A2(n_227), .B(n_338), .Y(n_337) );
NAND2xp5_ASAP7_75t_L g674 ( .A(n_211), .B(n_639), .Y(n_674) );
CKINVDCx6p67_ASAP7_75t_R g739 ( .A(n_213), .Y(n_739) );
AOI22xp33_ASAP7_75t_L g731 ( .A1(n_215), .A2(n_279), .B1(n_720), .B2(n_732), .Y(n_731) );
INVx1_ASAP7_75t_L g328 ( .A(n_217), .Y(n_328) );
AOI22xp33_ASAP7_75t_L g681 ( .A1(n_218), .A2(n_263), .B1(n_428), .B2(n_429), .Y(n_681) );
AOI221x1_ASAP7_75t_SL g442 ( .A1(n_220), .A2(n_221), .B1(n_345), .B2(n_443), .C(n_444), .Y(n_442) );
INVx1_ASAP7_75t_L g551 ( .A(n_222), .Y(n_551) );
AOI221xp5_ASAP7_75t_L g411 ( .A1(n_226), .A2(n_275), .B1(n_412), .B2(n_414), .C(n_416), .Y(n_411) );
NOR2xp33_ASAP7_75t_L g292 ( .A(n_227), .B(n_266), .Y(n_292) );
INVx1_ASAP7_75t_L g325 ( .A(n_227), .Y(n_325) );
AOI21xp33_ASAP7_75t_L g549 ( .A1(n_229), .A2(n_345), .B(n_550), .Y(n_549) );
AOI22xp33_ASAP7_75t_L g1003 ( .A1(n_232), .A2(n_246), .B1(n_350), .B2(n_400), .Y(n_1003) );
AOI221xp5_ASAP7_75t_L g390 ( .A1(n_233), .A2(n_270), .B1(n_391), .B2(n_393), .C(n_397), .Y(n_390) );
AOI21xp5_ASAP7_75t_L g490 ( .A1(n_235), .A2(n_491), .B(n_492), .Y(n_490) );
INVx1_ASAP7_75t_L g828 ( .A(n_239), .Y(n_828) );
INVx1_ASAP7_75t_L g679 ( .A(n_247), .Y(n_679) );
AOI22xp33_ASAP7_75t_L g465 ( .A1(n_250), .A2(n_269), .B1(n_382), .B2(n_466), .Y(n_465) );
AOI21xp33_ASAP7_75t_L g677 ( .A1(n_253), .A2(n_415), .B(n_678), .Y(n_677) );
AOI21xp5_ASAP7_75t_L g612 ( .A1(n_256), .A2(n_523), .B(n_613), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g662 ( .A(n_259), .B(n_663), .Y(n_662) );
NAND2xp5_ASAP7_75t_L g310 ( .A(n_266), .B(n_311), .Y(n_310) );
NAND2xp5_ASAP7_75t_L g579 ( .A(n_268), .B(n_580), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g349 ( .A(n_271), .B(n_350), .Y(n_349) );
INVx1_ASAP7_75t_L g528 ( .A(n_273), .Y(n_528) );
INVx1_ASAP7_75t_L g722 ( .A(n_274), .Y(n_722) );
AOI22xp33_ASAP7_75t_L g379 ( .A1(n_277), .A2(n_280), .B1(n_380), .B2(n_382), .Y(n_379) );
AOI21xp5_ASAP7_75t_L g282 ( .A1(n_283), .A2(n_294), .B(n_706), .Y(n_282) );
INVx1_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
BUFx4_ASAP7_75t_SL g284 ( .A(n_285), .Y(n_284) );
NAND3xp33_ASAP7_75t_L g285 ( .A(n_286), .B(n_289), .C(n_293), .Y(n_285) );
AND2x2_ASAP7_75t_L g967 ( .A(n_286), .B(n_968), .Y(n_967) );
AND2x2_ASAP7_75t_L g1006 ( .A(n_286), .B(n_969), .Y(n_1006) );
INVx1_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
OA21x2_ASAP7_75t_L g1008 ( .A1(n_287), .A2(n_751), .B(n_1009), .Y(n_1008) );
HB1xp67_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
AND2x2_ASAP7_75t_L g714 ( .A(n_288), .B(n_715), .Y(n_714) );
AND3x4_ASAP7_75t_L g750 ( .A(n_288), .B(n_721), .C(n_751), .Y(n_750) );
NOR2xp33_ASAP7_75t_L g968 ( .A(n_289), .B(n_969), .Y(n_968) );
HB1xp67_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
AO21x2_ASAP7_75t_L g403 ( .A1(n_290), .A2(n_404), .B(n_405), .Y(n_403) );
NAND2xp5_ASAP7_75t_L g290 ( .A(n_291), .B(n_292), .Y(n_290) );
INVx1_ASAP7_75t_L g969 ( .A(n_293), .Y(n_969) );
XNOR2xp5_ASAP7_75t_L g294 ( .A(n_295), .B(n_529), .Y(n_294) );
XNOR2x1_ASAP7_75t_L g295 ( .A(n_296), .B(n_470), .Y(n_295) );
INVx2_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
OA22x2_ASAP7_75t_L g297 ( .A1(n_298), .A2(n_407), .B1(n_408), .B2(n_469), .Y(n_297) );
INVx1_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
INVx1_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
INVx1_ASAP7_75t_L g469 ( .A(n_300), .Y(n_469) );
INVx2_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
NAND4xp75_ASAP7_75t_L g302 ( .A(n_303), .B(n_359), .C(n_378), .D(n_390), .Y(n_302) );
NOR2xp67_ASAP7_75t_L g303 ( .A(n_304), .B(n_342), .Y(n_303) );
OAI22xp5_ASAP7_75t_L g304 ( .A1(n_305), .A2(n_328), .B1(n_329), .B2(n_341), .Y(n_304) );
INVx3_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
BUFx6f_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
BUFx3_ASAP7_75t_L g458 ( .A(n_307), .Y(n_458) );
INVx2_ASAP7_75t_L g514 ( .A(n_307), .Y(n_514) );
AND2x2_ASAP7_75t_L g307 ( .A(n_308), .B(n_320), .Y(n_307) );
AND2x4_ASAP7_75t_L g346 ( .A(n_308), .B(n_347), .Y(n_346) );
AND2x4_ASAP7_75t_L g381 ( .A(n_308), .B(n_363), .Y(n_381) );
AND2x4_ASAP7_75t_L g431 ( .A(n_308), .B(n_347), .Y(n_431) );
AND2x4_ASAP7_75t_L g434 ( .A(n_308), .B(n_320), .Y(n_434) );
AND2x4_ASAP7_75t_L g437 ( .A(n_308), .B(n_363), .Y(n_437) );
AND2x4_ASAP7_75t_L g308 ( .A(n_309), .B(n_314), .Y(n_308) );
INVx2_ASAP7_75t_L g340 ( .A(n_309), .Y(n_340) );
AND2x2_ASAP7_75t_L g352 ( .A(n_309), .B(n_353), .Y(n_352) );
AND2x4_ASAP7_75t_L g365 ( .A(n_309), .B(n_366), .Y(n_365) );
OR2x2_ASAP7_75t_L g371 ( .A(n_309), .B(n_367), .Y(n_371) );
AND2x4_ASAP7_75t_L g309 ( .A(n_310), .B(n_313), .Y(n_309) );
NAND2xp5_ASAP7_75t_L g316 ( .A(n_311), .B(n_317), .Y(n_316) );
INVxp67_ASAP7_75t_L g334 ( .A(n_311), .Y(n_334) );
INVx3_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
NAND2xp33_ASAP7_75t_L g318 ( .A(n_312), .B(n_319), .Y(n_318) );
NAND2xp33_ASAP7_75t_L g322 ( .A(n_312), .B(n_323), .Y(n_322) );
INVx2_ASAP7_75t_L g326 ( .A(n_312), .Y(n_326) );
INVx1_ASAP7_75t_L g338 ( .A(n_312), .Y(n_338) );
HB1xp67_ASAP7_75t_L g354 ( .A(n_312), .Y(n_354) );
NAND3xp33_ASAP7_75t_L g405 ( .A(n_313), .B(n_333), .C(n_406), .Y(n_405) );
AND2x4_ASAP7_75t_L g339 ( .A(n_314), .B(n_340), .Y(n_339) );
INVx1_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
INVx1_ASAP7_75t_L g367 ( .A(n_315), .Y(n_367) );
AND2x2_ASAP7_75t_L g315 ( .A(n_316), .B(n_318), .Y(n_315) );
AND2x2_ASAP7_75t_L g374 ( .A(n_320), .B(n_365), .Y(n_374) );
AND2x4_ASAP7_75t_L g386 ( .A(n_320), .B(n_387), .Y(n_386) );
AND2x2_ASAP7_75t_L g396 ( .A(n_320), .B(n_339), .Y(n_396) );
AND2x2_ASAP7_75t_L g425 ( .A(n_320), .B(n_365), .Y(n_425) );
AND2x4_ASAP7_75t_L g484 ( .A(n_320), .B(n_365), .Y(n_484) );
AND2x4_ASAP7_75t_L g485 ( .A(n_320), .B(n_370), .Y(n_485) );
AND2x2_ASAP7_75t_L g491 ( .A(n_320), .B(n_339), .Y(n_491) );
AND2x2_ASAP7_75t_L g320 ( .A(n_321), .B(n_327), .Y(n_320) );
INVx1_ASAP7_75t_L g348 ( .A(n_321), .Y(n_348) );
NAND2xp5_ASAP7_75t_L g321 ( .A(n_322), .B(n_324), .Y(n_321) );
NAND2xp5_ASAP7_75t_L g335 ( .A(n_323), .B(n_336), .Y(n_335) );
NAND2xp5_ASAP7_75t_L g324 ( .A(n_325), .B(n_326), .Y(n_324) );
OAI21xp5_ASAP7_75t_L g357 ( .A1(n_325), .A2(n_338), .B(n_358), .Y(n_357) );
AND2x2_ASAP7_75t_L g347 ( .A(n_327), .B(n_348), .Y(n_347) );
AND2x2_ASAP7_75t_L g356 ( .A(n_327), .B(n_357), .Y(n_356) );
INVx1_ASAP7_75t_L g364 ( .A(n_327), .Y(n_364) );
OAI22xp5_ASAP7_75t_L g982 ( .A1(n_329), .A2(n_983), .B1(n_984), .B2(n_985), .Y(n_982) );
INVx3_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
BUFx6f_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
BUFx6f_ASAP7_75t_L g463 ( .A(n_331), .Y(n_463) );
INVx3_ASAP7_75t_L g517 ( .A(n_331), .Y(n_517) );
AND2x4_ASAP7_75t_L g331 ( .A(n_332), .B(n_339), .Y(n_331) );
AND2x4_ASAP7_75t_L g377 ( .A(n_332), .B(n_365), .Y(n_377) );
AND2x4_ASAP7_75t_L g389 ( .A(n_332), .B(n_370), .Y(n_389) );
AND2x4_ASAP7_75t_L g421 ( .A(n_332), .B(n_365), .Y(n_421) );
AND2x4_ASAP7_75t_L g429 ( .A(n_332), .B(n_370), .Y(n_429) );
AND2x4_ASAP7_75t_L g432 ( .A(n_332), .B(n_339), .Y(n_432) );
AND2x2_ASAP7_75t_L g332 ( .A(n_333), .B(n_337), .Y(n_332) );
NAND2xp5_ASAP7_75t_L g333 ( .A(n_334), .B(n_335), .Y(n_333) );
AND2x2_ASAP7_75t_L g383 ( .A(n_339), .B(n_363), .Y(n_383) );
AND2x4_ASAP7_75t_L g392 ( .A(n_339), .B(n_347), .Y(n_392) );
AND2x2_ASAP7_75t_L g415 ( .A(n_339), .B(n_347), .Y(n_415) );
AND2x4_ASAP7_75t_L g438 ( .A(n_339), .B(n_363), .Y(n_438) );
OAI21xp5_ASAP7_75t_L g342 ( .A1(n_343), .A2(n_344), .B(n_349), .Y(n_342) );
OAI22xp5_ASAP7_75t_L g986 ( .A1(n_344), .A2(n_987), .B1(n_988), .B2(n_989), .Y(n_986) );
INVx4_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
BUFx6f_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
BUFx3_ASAP7_75t_L g476 ( .A(n_346), .Y(n_476) );
BUFx3_ASAP7_75t_L g591 ( .A(n_346), .Y(n_591) );
INVx1_ASAP7_75t_L g634 ( .A(n_346), .Y(n_634) );
AND2x4_ASAP7_75t_L g363 ( .A(n_348), .B(n_364), .Y(n_363) );
BUFx4f_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
INVx5_ASAP7_75t_L g460 ( .A(n_351), .Y(n_460) );
BUFx2_ASAP7_75t_L g582 ( .A(n_351), .Y(n_582) );
BUFx2_ASAP7_75t_L g960 ( .A(n_351), .Y(n_960) );
AND2x4_ASAP7_75t_L g351 ( .A(n_352), .B(n_356), .Y(n_351) );
AND2x2_ASAP7_75t_L g435 ( .A(n_352), .B(n_356), .Y(n_435) );
AND2x4_ASAP7_75t_L g617 ( .A(n_352), .B(n_356), .Y(n_617) );
NAND2xp5_ASAP7_75t_L g353 ( .A(n_354), .B(n_355), .Y(n_353) );
INVx1_ASAP7_75t_L g404 ( .A(n_354), .Y(n_404) );
AND2x2_ASAP7_75t_L g359 ( .A(n_360), .B(n_372), .Y(n_359) );
INVx1_ASAP7_75t_L g993 ( .A(n_361), .Y(n_993) );
BUFx12f_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
BUFx6f_ASAP7_75t_L g454 ( .A(n_362), .Y(n_454) );
BUFx6f_ASAP7_75t_L g509 ( .A(n_362), .Y(n_509) );
AND2x4_ASAP7_75t_L g362 ( .A(n_363), .B(n_365), .Y(n_362) );
AND2x4_ASAP7_75t_L g369 ( .A(n_363), .B(n_370), .Y(n_369) );
AND2x4_ASAP7_75t_L g420 ( .A(n_363), .B(n_365), .Y(n_420) );
AND2x4_ASAP7_75t_L g428 ( .A(n_363), .B(n_387), .Y(n_428) );
INVx1_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
BUFx6f_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
BUFx6f_ASAP7_75t_L g455 ( .A(n_369), .Y(n_455) );
BUFx6f_ASAP7_75t_L g501 ( .A(n_369), .Y(n_501) );
BUFx6f_ASAP7_75t_L g600 ( .A(n_369), .Y(n_600) );
INVx2_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
INVx2_ASAP7_75t_L g387 ( .A(n_371), .Y(n_387) );
BUFx6f_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
BUFx8_ASAP7_75t_L g503 ( .A(n_374), .Y(n_503) );
INVx2_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
INVx2_ASAP7_75t_L g468 ( .A(n_376), .Y(n_468) );
INVx1_ASAP7_75t_L g510 ( .A(n_376), .Y(n_510) );
INVx4_ASAP7_75t_L g543 ( .A(n_376), .Y(n_543) );
INVx4_ASAP7_75t_L g690 ( .A(n_376), .Y(n_690) );
INVx1_ASAP7_75t_L g980 ( .A(n_376), .Y(n_980) );
INVx8_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
AND2x2_ASAP7_75t_L g378 ( .A(n_379), .B(n_384), .Y(n_378) );
BUFx6f_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
BUFx12f_ASAP7_75t_L g466 ( .A(n_381), .Y(n_466) );
INVx3_ASAP7_75t_L g659 ( .A(n_381), .Y(n_659) );
BUFx6f_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
BUFx5_ASAP7_75t_L g507 ( .A(n_383), .Y(n_507) );
INVx1_ASAP7_75t_L g541 ( .A(n_383), .Y(n_541) );
BUFx3_ASAP7_75t_L g571 ( .A(n_383), .Y(n_571) );
BUFx12f_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
BUFx6f_ASAP7_75t_L g423 ( .A(n_386), .Y(n_423) );
BUFx3_ASAP7_75t_L g504 ( .A(n_386), .Y(n_504) );
BUFx6f_ASAP7_75t_L g568 ( .A(n_386), .Y(n_568) );
BUFx6f_ASAP7_75t_L g656 ( .A(n_386), .Y(n_656) );
BUFx12f_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
INVx6_ASAP7_75t_L g452 ( .A(n_389), .Y(n_452) );
BUFx3_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
BUFx8_ASAP7_75t_SL g462 ( .A(n_392), .Y(n_462) );
INVx2_ASAP7_75t_L g554 ( .A(n_392), .Y(n_554) );
BUFx6f_ASAP7_75t_L g578 ( .A(n_392), .Y(n_578) );
INVx2_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
INVx1_ASAP7_75t_L g443 ( .A(n_394), .Y(n_443) );
INVx2_ASAP7_75t_L g663 ( .A(n_394), .Y(n_663) );
BUFx6f_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
INVx2_ASAP7_75t_L g639 ( .A(n_395), .Y(n_639) );
INVx2_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
INVx3_ASAP7_75t_L g413 ( .A(n_396), .Y(n_413) );
BUFx3_ASAP7_75t_L g523 ( .A(n_396), .Y(n_523) );
NOR2xp33_ASAP7_75t_L g397 ( .A(n_398), .B(n_399), .Y(n_397) );
INVx2_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
INVx4_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
NOR2xp33_ASAP7_75t_L g416 ( .A(n_401), .B(n_417), .Y(n_416) );
NOR2xp33_ASAP7_75t_L g678 ( .A(n_401), .B(n_679), .Y(n_678) );
INVx4_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
INVx3_ASAP7_75t_L g494 ( .A(n_402), .Y(n_494) );
INVx3_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
BUFx6f_ASAP7_75t_L g448 ( .A(n_403), .Y(n_448) );
INVx1_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
XNOR2xp5_ASAP7_75t_L g408 ( .A(n_409), .B(n_439), .Y(n_408) );
NAND3x1_ASAP7_75t_L g410 ( .A(n_411), .B(n_418), .C(n_426), .Y(n_410) );
HB1xp67_ASAP7_75t_L g556 ( .A(n_412), .Y(n_556) );
INVx2_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
INVx2_ASAP7_75t_L g580 ( .A(n_413), .Y(n_580) );
HB1xp67_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
AND2x2_ASAP7_75t_L g418 ( .A(n_419), .B(n_422), .Y(n_418) );
BUFx6f_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
BUFx4f_ASAP7_75t_L g567 ( .A(n_425), .Y(n_567) );
AND4x1_ASAP7_75t_L g426 ( .A(n_427), .B(n_430), .C(n_433), .D(n_436), .Y(n_426) );
INVx2_ASAP7_75t_L g620 ( .A(n_434), .Y(n_620) );
XOR2xp5_ASAP7_75t_L g439 ( .A(n_440), .B(n_441), .Y(n_439) );
NAND4xp75_ASAP7_75t_L g441 ( .A(n_442), .B(n_449), .C(n_456), .D(n_464), .Y(n_441) );
NOR2xp33_ASAP7_75t_L g444 ( .A(n_445), .B(n_446), .Y(n_444) );
OAI22xp5_ASAP7_75t_L g524 ( .A1(n_446), .A2(n_525), .B1(n_526), .B2(n_528), .Y(n_524) );
INVx2_ASAP7_75t_SL g446 ( .A(n_447), .Y(n_446) );
INVx2_ASAP7_75t_SL g447 ( .A(n_448), .Y(n_447) );
BUFx6f_ASAP7_75t_L g576 ( .A(n_448), .Y(n_576) );
BUFx6f_ASAP7_75t_L g644 ( .A(n_448), .Y(n_644) );
INVx1_ASAP7_75t_L g667 ( .A(n_448), .Y(n_667) );
AND2x2_ASAP7_75t_L g449 ( .A(n_450), .B(n_453), .Y(n_449) );
INVx5_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
INVx2_ASAP7_75t_L g978 ( .A(n_452), .Y(n_978) );
AND2x2_ASAP7_75t_L g456 ( .A(n_457), .B(n_461), .Y(n_456) );
INVx2_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
INVx3_ASAP7_75t_L g478 ( .A(n_460), .Y(n_478) );
INVx4_ASAP7_75t_L g527 ( .A(n_460), .Y(n_527) );
INVx2_ASAP7_75t_L g558 ( .A(n_460), .Y(n_558) );
INVx1_ASAP7_75t_L g489 ( .A(n_462), .Y(n_489) );
AND2x2_ASAP7_75t_L g464 ( .A(n_465), .B(n_467), .Y(n_464) );
AOI22xp5_ASAP7_75t_L g470 ( .A1(n_471), .A2(n_472), .B1(n_496), .B2(n_497), .Y(n_470) );
INVx1_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
XOR2x2_ASAP7_75t_L g472 ( .A(n_473), .B(n_495), .Y(n_472) );
NOR4xp75_ASAP7_75t_L g473 ( .A(n_474), .B(n_479), .C(n_482), .D(n_487), .Y(n_473) );
NAND2xp5_ASAP7_75t_L g474 ( .A(n_475), .B(n_477), .Y(n_474) );
INVx2_ASAP7_75t_L g952 ( .A(n_476), .Y(n_952) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_480), .B(n_481), .Y(n_479) );
NAND2xp5_ASAP7_75t_SL g482 ( .A(n_483), .B(n_486), .Y(n_482) );
OAI21x1_ASAP7_75t_SL g487 ( .A1(n_488), .A2(n_489), .B(n_490), .Y(n_487) );
INVx2_ASAP7_75t_L g699 ( .A(n_491), .Y(n_699) );
NOR2xp33_ASAP7_75t_L g492 ( .A(n_493), .B(n_494), .Y(n_492) );
NOR2xp33_ASAP7_75t_L g550 ( .A(n_494), .B(n_551), .Y(n_550) );
NOR2xp33_ASAP7_75t_L g592 ( .A(n_494), .B(n_593), .Y(n_592) );
NOR2xp33_ASAP7_75t_L g610 ( .A(n_494), .B(n_611), .Y(n_610) );
NOR2xp33_ASAP7_75t_L g700 ( .A(n_494), .B(n_701), .Y(n_700) );
INVx2_ASAP7_75t_SL g496 ( .A(n_497), .Y(n_496) );
NAND4xp75_ASAP7_75t_SL g498 ( .A(n_499), .B(n_505), .C(n_511), .D(n_518), .Y(n_498) );
AND2x2_ASAP7_75t_L g499 ( .A(n_500), .B(n_502), .Y(n_499) );
AND2x2_ASAP7_75t_L g505 ( .A(n_506), .B(n_508), .Y(n_505) );
AND2x2_ASAP7_75t_L g511 ( .A(n_512), .B(n_515), .Y(n_511) );
INVx1_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
BUFx6f_ASAP7_75t_L g560 ( .A(n_514), .Y(n_560) );
INVx2_ASAP7_75t_L g954 ( .A(n_514), .Y(n_954) );
INVx2_ASAP7_75t_L g516 ( .A(n_517), .Y(n_516) );
INVx1_ASAP7_75t_L g519 ( .A(n_520), .Y(n_519) );
INVx1_ASAP7_75t_L g520 ( .A(n_521), .Y(n_520) );
INVx2_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
INVx2_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
INVx1_ASAP7_75t_L g957 ( .A(n_523), .Y(n_957) );
INVx2_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
XNOR2xp5_ASAP7_75t_L g529 ( .A(n_530), .B(n_602), .Y(n_529) );
AOI22xp5_ASAP7_75t_L g530 ( .A1(n_531), .A2(n_583), .B1(n_584), .B2(n_601), .Y(n_530) );
HB1xp67_ASAP7_75t_L g531 ( .A(n_532), .Y(n_531) );
INVx1_ASAP7_75t_L g601 ( .A(n_532), .Y(n_601) );
AO22x2_ASAP7_75t_L g532 ( .A1(n_533), .A2(n_534), .B1(n_561), .B2(n_562), .Y(n_532) );
INVx2_ASAP7_75t_SL g533 ( .A(n_534), .Y(n_533) );
XNOR2x1_ASAP7_75t_L g534 ( .A(n_535), .B(n_536), .Y(n_534) );
NOR2x1_ASAP7_75t_L g536 ( .A(n_537), .B(n_546), .Y(n_536) );
NAND4xp25_ASAP7_75t_L g537 ( .A(n_538), .B(n_542), .C(n_544), .D(n_545), .Y(n_537) );
BUFx6f_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
INVx2_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
NAND3xp33_ASAP7_75t_L g546 ( .A(n_547), .B(n_555), .C(n_557), .Y(n_546) );
INVx1_ASAP7_75t_L g547 ( .A(n_548), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_549), .B(n_552), .Y(n_548) );
INVx3_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
INVx2_ASAP7_75t_L g636 ( .A(n_554), .Y(n_636) );
INVx2_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
HB1xp67_ASAP7_75t_L g989 ( .A(n_560), .Y(n_989) );
INVx1_ASAP7_75t_SL g561 ( .A(n_562), .Y(n_561) );
NOR2x1_ASAP7_75t_L g563 ( .A(n_564), .B(n_572), .Y(n_563) );
NAND4xp25_ASAP7_75t_L g564 ( .A(n_565), .B(n_566), .C(n_569), .D(n_570), .Y(n_564) );
BUFx2_ASAP7_75t_L g998 ( .A(n_571), .Y(n_998) );
NAND4xp25_ASAP7_75t_SL g572 ( .A(n_573), .B(n_577), .C(n_579), .D(n_581), .Y(n_572) );
NOR2xp33_ASAP7_75t_L g574 ( .A(n_575), .B(n_576), .Y(n_574) );
BUFx3_ASAP7_75t_L g949 ( .A(n_578), .Y(n_949) );
INVx2_ASAP7_75t_L g984 ( .A(n_578), .Y(n_984) );
INVx1_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
HB1xp67_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
NOR2x1_ASAP7_75t_L g586 ( .A(n_587), .B(n_595), .Y(n_586) );
NAND4xp25_ASAP7_75t_L g587 ( .A(n_588), .B(n_589), .C(n_590), .D(n_594), .Y(n_587) );
NAND4xp25_ASAP7_75t_SL g595 ( .A(n_596), .B(n_597), .C(n_598), .D(n_599), .Y(n_595) );
BUFx3_ASAP7_75t_L g994 ( .A(n_600), .Y(n_994) );
AOI22xp5_ASAP7_75t_L g602 ( .A1(n_603), .A2(n_604), .B1(n_650), .B2(n_705), .Y(n_602) );
INVx1_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
BUFx2_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
XNOR2xp5_ASAP7_75t_SL g605 ( .A(n_606), .B(n_629), .Y(n_605) );
INVx1_ASAP7_75t_L g628 ( .A(n_607), .Y(n_628) );
NOR2x1_ASAP7_75t_L g607 ( .A(n_608), .B(n_622), .Y(n_607) );
NAND3xp33_ASAP7_75t_L g608 ( .A(n_609), .B(n_612), .C(n_621), .Y(n_608) );
OAI22xp5_ASAP7_75t_L g613 ( .A1(n_614), .A2(n_616), .B1(n_618), .B2(n_620), .Y(n_613) );
CKINVDCx16_ASAP7_75t_R g614 ( .A(n_615), .Y(n_614) );
OAI21xp5_ASAP7_75t_L g640 ( .A1(n_616), .A2(n_641), .B(n_642), .Y(n_640) );
INVx4_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
CKINVDCx9p33_ASAP7_75t_R g618 ( .A(n_619), .Y(n_618) );
NAND4xp25_ASAP7_75t_L g622 ( .A(n_623), .B(n_624), .C(n_625), .D(n_626), .Y(n_622) );
NOR2x1_ASAP7_75t_SL g630 ( .A(n_631), .B(n_645), .Y(n_630) );
NAND3xp33_ASAP7_75t_L g631 ( .A(n_632), .B(n_635), .C(n_637), .Y(n_631) );
INVx2_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
BUFx3_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
INVx1_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
INVx2_ASAP7_75t_L g963 ( .A(n_644), .Y(n_963) );
NAND4xp25_ASAP7_75t_SL g645 ( .A(n_646), .B(n_647), .C(n_648), .D(n_649), .Y(n_645) );
INVx2_ASAP7_75t_L g705 ( .A(n_650), .Y(n_705) );
OA22x2_ASAP7_75t_L g650 ( .A1(n_651), .A2(n_669), .B1(n_703), .B2(n_704), .Y(n_650) );
INVx1_ASAP7_75t_SL g703 ( .A(n_651), .Y(n_703) );
XOR2x2_ASAP7_75t_L g651 ( .A(n_652), .B(n_668), .Y(n_651) );
NOR2x1_ASAP7_75t_L g652 ( .A(n_653), .B(n_661), .Y(n_652) );
NAND4xp25_ASAP7_75t_L g653 ( .A(n_654), .B(n_655), .C(n_657), .D(n_660), .Y(n_653) );
INVx1_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
INVx2_ASAP7_75t_L g997 ( .A(n_659), .Y(n_997) );
NAND4xp25_ASAP7_75t_L g661 ( .A(n_662), .B(n_664), .C(n_665), .D(n_666), .Y(n_661) );
INVx1_ASAP7_75t_L g704 ( .A(n_669), .Y(n_704) );
XNOR2x1_ASAP7_75t_L g669 ( .A(n_670), .B(n_685), .Y(n_669) );
XNOR2x1_ASAP7_75t_L g670 ( .A(n_671), .B(n_672), .Y(n_670) );
OR2x2_ASAP7_75t_L g672 ( .A(n_673), .B(n_680), .Y(n_672) );
NAND4xp25_ASAP7_75t_L g673 ( .A(n_674), .B(n_675), .C(n_676), .D(n_677), .Y(n_673) );
NAND4xp25_ASAP7_75t_L g680 ( .A(n_681), .B(n_682), .C(n_683), .D(n_684), .Y(n_680) );
XNOR2x1_ASAP7_75t_L g685 ( .A(n_686), .B(n_702), .Y(n_685) );
NAND4xp75_ASAP7_75t_L g686 ( .A(n_687), .B(n_691), .C(n_694), .D(n_697), .Y(n_686) );
AND2x2_ASAP7_75t_L g687 ( .A(n_688), .B(n_689), .Y(n_687) );
AND2x2_ASAP7_75t_L g691 ( .A(n_692), .B(n_693), .Y(n_691) );
AND2x2_ASAP7_75t_L g694 ( .A(n_695), .B(n_696), .Y(n_694) );
INVx2_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
OAI221xp5_ASAP7_75t_SL g706 ( .A1(n_707), .A2(n_933), .B1(n_936), .B2(n_965), .C(n_970), .Y(n_706) );
O2A1O1Ixp33_ASAP7_75t_L g707 ( .A1(n_708), .A2(n_799), .B(n_824), .C(n_830), .Y(n_707) );
OAI211xp5_ASAP7_75t_L g708 ( .A1(n_709), .A2(n_733), .B(n_763), .C(n_782), .Y(n_708) );
INVx1_ASAP7_75t_L g884 ( .A(n_709), .Y(n_884) );
NAND2xp5_ASAP7_75t_L g709 ( .A(n_710), .B(n_726), .Y(n_709) );
AND2x2_ASAP7_75t_L g780 ( .A(n_710), .B(n_781), .Y(n_780) );
INVx2_ASAP7_75t_L g810 ( .A(n_710), .Y(n_810) );
NOR2xp33_ASAP7_75t_L g832 ( .A(n_710), .B(n_825), .Y(n_832) );
NAND2xp5_ASAP7_75t_L g910 ( .A(n_710), .B(n_825), .Y(n_910) );
NOR3xp33_ASAP7_75t_L g929 ( .A(n_710), .B(n_815), .C(n_930), .Y(n_929) );
INVx3_ASAP7_75t_L g710 ( .A(n_711), .Y(n_710) );
OR2x2_ASAP7_75t_L g793 ( .A(n_711), .B(n_726), .Y(n_793) );
NOR2xp33_ASAP7_75t_L g854 ( .A(n_711), .B(n_786), .Y(n_854) );
AND2x2_ASAP7_75t_L g890 ( .A(n_711), .B(n_891), .Y(n_890) );
NAND2xp5_ASAP7_75t_L g915 ( .A(n_711), .B(n_726), .Y(n_915) );
NAND2xp5_ASAP7_75t_L g916 ( .A(n_711), .B(n_818), .Y(n_916) );
AND2x2_ASAP7_75t_L g927 ( .A(n_711), .B(n_727), .Y(n_927) );
AND2x4_ASAP7_75t_L g711 ( .A(n_712), .B(n_719), .Y(n_711) );
AND2x2_ASAP7_75t_L g713 ( .A(n_714), .B(n_716), .Y(n_713) );
AND2x4_ASAP7_75t_L g720 ( .A(n_714), .B(n_721), .Y(n_720) );
AND2x4_ASAP7_75t_L g729 ( .A(n_714), .B(n_716), .Y(n_729) );
AND2x2_ASAP7_75t_L g753 ( .A(n_714), .B(n_716), .Y(n_753) );
AND2x4_ASAP7_75t_L g717 ( .A(n_716), .B(n_718), .Y(n_717) );
AND2x2_ASAP7_75t_L g730 ( .A(n_716), .B(n_718), .Y(n_730) );
AND2x2_ASAP7_75t_L g754 ( .A(n_716), .B(n_718), .Y(n_754) );
INVx2_ASAP7_75t_L g746 ( .A(n_717), .Y(n_746) );
AND2x4_ASAP7_75t_L g725 ( .A(n_718), .B(n_721), .Y(n_725) );
AND2x4_ASAP7_75t_L g732 ( .A(n_718), .B(n_721), .Y(n_732) );
NAND2xp5_ASAP7_75t_L g740 ( .A(n_718), .B(n_721), .Y(n_740) );
INVx3_ASAP7_75t_L g738 ( .A(n_720), .Y(n_738) );
CKINVDCx5p33_ASAP7_75t_R g1009 ( .A(n_721), .Y(n_1009) );
INVx2_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
INVx2_ASAP7_75t_SL g724 ( .A(n_725), .Y(n_724) );
INVx3_ASAP7_75t_L g807 ( .A(n_726), .Y(n_807) );
AND2x2_ASAP7_75t_L g811 ( .A(n_726), .B(n_736), .Y(n_811) );
INVx2_ASAP7_75t_L g726 ( .A(n_727), .Y(n_726) );
AND2x2_ASAP7_75t_L g818 ( .A(n_727), .B(n_736), .Y(n_818) );
AND2x2_ASAP7_75t_L g849 ( .A(n_727), .B(n_781), .Y(n_849) );
OR2x2_ASAP7_75t_L g859 ( .A(n_727), .B(n_736), .Y(n_859) );
AND2x2_ASAP7_75t_L g727 ( .A(n_728), .B(n_731), .Y(n_727) );
INVx3_ASAP7_75t_L g744 ( .A(n_729), .Y(n_744) );
NAND2xp5_ASAP7_75t_L g733 ( .A(n_734), .B(n_747), .Y(n_733) );
INVx2_ASAP7_75t_L g837 ( .A(n_734), .Y(n_837) );
O2A1O1Ixp33_ASAP7_75t_SL g894 ( .A1(n_734), .A2(n_765), .B(n_895), .C(n_897), .Y(n_894) );
BUFx2_ASAP7_75t_L g734 ( .A(n_735), .Y(n_734) );
NOR2xp33_ASAP7_75t_L g783 ( .A(n_735), .B(n_784), .Y(n_783) );
NOR2xp33_ASAP7_75t_L g794 ( .A(n_735), .B(n_795), .Y(n_794) );
INVx1_ASAP7_75t_L g844 ( .A(n_735), .Y(n_844) );
AND2x2_ASAP7_75t_L g877 ( .A(n_735), .B(n_855), .Y(n_877) );
O2A1O1Ixp33_ASAP7_75t_L g881 ( .A1(n_735), .A2(n_882), .B(n_883), .C(n_884), .Y(n_881) );
INVx2_ASAP7_75t_L g735 ( .A(n_736), .Y(n_735) );
INVx3_ASAP7_75t_L g781 ( .A(n_736), .Y(n_781) );
NOR2xp33_ASAP7_75t_L g823 ( .A(n_736), .B(n_770), .Y(n_823) );
OR2x2_ASAP7_75t_L g736 ( .A(n_737), .B(n_742), .Y(n_736) );
OAI22xp5_ASAP7_75t_L g737 ( .A1(n_738), .A2(n_739), .B1(n_740), .B2(n_741), .Y(n_737) );
OAI221xp5_ASAP7_75t_L g826 ( .A1(n_738), .A2(n_740), .B1(n_827), .B2(n_828), .C(n_829), .Y(n_826) );
OAI22xp5_ASAP7_75t_L g771 ( .A1(n_740), .A2(n_772), .B1(n_773), .B2(n_774), .Y(n_771) );
BUFx2_ASAP7_75t_L g935 ( .A(n_740), .Y(n_935) );
OAI22xp5_ASAP7_75t_L g742 ( .A1(n_743), .A2(n_744), .B1(n_745), .B2(n_746), .Y(n_742) );
AND2x2_ASAP7_75t_L g769 ( .A(n_747), .B(n_770), .Y(n_769) );
INVx1_ASAP7_75t_L g847 ( .A(n_747), .Y(n_847) );
AND2x2_ASAP7_75t_L g747 ( .A(n_748), .B(n_755), .Y(n_747) );
CKINVDCx6p67_ASAP7_75t_R g766 ( .A(n_748), .Y(n_766) );
NAND2xp5_ASAP7_75t_L g784 ( .A(n_748), .B(n_760), .Y(n_784) );
INVx1_ASAP7_75t_L g791 ( .A(n_748), .Y(n_791) );
AND2x2_ASAP7_75t_L g803 ( .A(n_748), .B(n_804), .Y(n_803) );
OR2x2_ASAP7_75t_L g874 ( .A(n_748), .B(n_760), .Y(n_874) );
AND2x2_ASAP7_75t_L g748 ( .A(n_749), .B(n_752), .Y(n_748) );
INVx1_ASAP7_75t_L g772 ( .A(n_750), .Y(n_772) );
INVx1_ASAP7_75t_L g779 ( .A(n_753), .Y(n_779) );
INVx1_ASAP7_75t_L g777 ( .A(n_754), .Y(n_777) );
AND2x2_ASAP7_75t_SL g900 ( .A(n_755), .B(n_766), .Y(n_900) );
AND2x2_ASAP7_75t_L g907 ( .A(n_755), .B(n_836), .Y(n_907) );
OR2x2_ASAP7_75t_L g913 ( .A(n_755), .B(n_804), .Y(n_913) );
INVxp33_ASAP7_75t_L g920 ( .A(n_755), .Y(n_920) );
AND2x2_ASAP7_75t_L g755 ( .A(n_756), .B(n_759), .Y(n_755) );
INVx1_ASAP7_75t_L g768 ( .A(n_756), .Y(n_768) );
AND2x2_ASAP7_75t_L g796 ( .A(n_756), .B(n_760), .Y(n_796) );
NAND2xp5_ASAP7_75t_L g756 ( .A(n_757), .B(n_758), .Y(n_756) );
AND2x2_ASAP7_75t_L g767 ( .A(n_759), .B(n_768), .Y(n_767) );
NAND2xp5_ASAP7_75t_L g871 ( .A(n_759), .B(n_790), .Y(n_871) );
OAI222xp33_ASAP7_75t_L g904 ( .A1(n_759), .A2(n_888), .B1(n_893), .B2(n_905), .C1(n_906), .C2(n_908), .Y(n_904) );
CKINVDCx5p33_ASAP7_75t_R g759 ( .A(n_760), .Y(n_759) );
AND2x2_ASAP7_75t_L g804 ( .A(n_760), .B(n_768), .Y(n_804) );
AOI322xp5_ASAP7_75t_L g853 ( .A1(n_760), .A2(n_807), .A3(n_809), .B1(n_844), .B2(n_854), .C1(n_855), .C2(n_857), .Y(n_853) );
AND2x4_ASAP7_75t_SL g760 ( .A(n_761), .B(n_762), .Y(n_760) );
OAI21xp5_ASAP7_75t_L g763 ( .A1(n_764), .A2(n_769), .B(n_780), .Y(n_763) );
INVx1_ASAP7_75t_L g764 ( .A(n_765), .Y(n_764) );
NAND2xp5_ASAP7_75t_L g765 ( .A(n_766), .B(n_767), .Y(n_765) );
AND2x2_ASAP7_75t_L g797 ( .A(n_766), .B(n_798), .Y(n_797) );
NAND2xp5_ASAP7_75t_L g805 ( .A(n_766), .B(n_796), .Y(n_805) );
NAND2xp5_ASAP7_75t_L g816 ( .A(n_766), .B(n_770), .Y(n_816) );
NOR2xp33_ASAP7_75t_L g817 ( .A(n_766), .B(n_812), .Y(n_817) );
AND2x2_ASAP7_75t_L g840 ( .A(n_766), .B(n_768), .Y(n_840) );
OAI22xp5_ASAP7_75t_L g845 ( .A1(n_766), .A2(n_846), .B1(n_847), .B2(n_848), .Y(n_845) );
AND2x2_ASAP7_75t_L g865 ( .A(n_766), .B(n_804), .Y(n_865) );
NAND2xp5_ASAP7_75t_L g885 ( .A(n_766), .B(n_843), .Y(n_885) );
AND2x2_ASAP7_75t_L g835 ( .A(n_767), .B(n_836), .Y(n_835) );
AND2x2_ASAP7_75t_L g843 ( .A(n_767), .B(n_770), .Y(n_843) );
INVx1_ASAP7_75t_L g858 ( .A(n_767), .Y(n_858) );
NOR2xp33_ASAP7_75t_L g789 ( .A(n_768), .B(n_790), .Y(n_789) );
AND2x2_ASAP7_75t_L g822 ( .A(n_768), .B(n_790), .Y(n_822) );
INVx1_ASAP7_75t_L g852 ( .A(n_768), .Y(n_852) );
INVx1_ASAP7_75t_L g787 ( .A(n_770), .Y(n_787) );
CKINVDCx6p67_ASAP7_75t_R g798 ( .A(n_770), .Y(n_798) );
AND2x2_ASAP7_75t_L g861 ( .A(n_770), .B(n_781), .Y(n_861) );
NAND2xp5_ASAP7_75t_L g893 ( .A(n_770), .B(n_789), .Y(n_893) );
NOR2xp33_ASAP7_75t_L g925 ( .A(n_770), .B(n_781), .Y(n_925) );
OR2x6_ASAP7_75t_SL g770 ( .A(n_771), .B(n_775), .Y(n_770) );
OAI22xp5_ASAP7_75t_L g775 ( .A1(n_776), .A2(n_777), .B1(n_778), .B2(n_779), .Y(n_775) );
NOR2xp33_ASAP7_75t_L g868 ( .A(n_781), .B(n_793), .Y(n_868) );
NAND2xp5_ASAP7_75t_L g883 ( .A(n_781), .B(n_810), .Y(n_883) );
NAND2xp5_ASAP7_75t_L g895 ( .A(n_781), .B(n_896), .Y(n_895) );
NOR2xp33_ASAP7_75t_L g931 ( .A(n_781), .B(n_798), .Y(n_931) );
O2A1O1Ixp33_ASAP7_75t_L g782 ( .A1(n_783), .A2(n_785), .B(n_792), .C(n_794), .Y(n_782) );
NOR2xp33_ASAP7_75t_L g785 ( .A(n_786), .B(n_788), .Y(n_785) );
NAND2xp5_ASAP7_75t_L g879 ( .A(n_786), .B(n_803), .Y(n_879) );
NAND2xp5_ASAP7_75t_L g905 ( .A(n_786), .B(n_849), .Y(n_905) );
NOR2xp33_ASAP7_75t_L g919 ( .A(n_786), .B(n_920), .Y(n_919) );
INVx3_ASAP7_75t_L g786 ( .A(n_787), .Y(n_786) );
INVx1_ASAP7_75t_L g788 ( .A(n_789), .Y(n_788) );
AND2x2_ASAP7_75t_L g836 ( .A(n_790), .B(n_798), .Y(n_836) );
AND2x2_ASAP7_75t_L g842 ( .A(n_790), .B(n_843), .Y(n_842) );
NAND2xp5_ASAP7_75t_L g851 ( .A(n_790), .B(n_852), .Y(n_851) );
INVx1_ASAP7_75t_L g790 ( .A(n_791), .Y(n_790) );
AOI221xp5_ASAP7_75t_L g876 ( .A1(n_792), .A2(n_825), .B1(n_877), .B2(n_878), .C(n_880), .Y(n_876) );
INVx1_ASAP7_75t_L g792 ( .A(n_793), .Y(n_792) );
NAND2xp5_ASAP7_75t_L g795 ( .A(n_796), .B(n_797), .Y(n_795) );
INVx1_ASAP7_75t_L g812 ( .A(n_796), .Y(n_812) );
AND2x2_ASAP7_75t_L g855 ( .A(n_796), .B(n_856), .Y(n_855) );
AND2x2_ASAP7_75t_L g896 ( .A(n_796), .B(n_836), .Y(n_896) );
INVxp67_ASAP7_75t_L g914 ( .A(n_797), .Y(n_914) );
NAND2xp5_ASAP7_75t_L g806 ( .A(n_798), .B(n_807), .Y(n_806) );
NAND2xp5_ASAP7_75t_L g838 ( .A(n_798), .B(n_818), .Y(n_838) );
NAND2xp5_ASAP7_75t_L g848 ( .A(n_798), .B(n_849), .Y(n_848) );
NAND2xp5_ASAP7_75t_L g864 ( .A(n_798), .B(n_865), .Y(n_864) );
NOR2xp33_ASAP7_75t_L g870 ( .A(n_798), .B(n_871), .Y(n_870) );
NOR2xp33_ASAP7_75t_L g875 ( .A(n_798), .B(n_859), .Y(n_875) );
OAI221xp5_ASAP7_75t_L g799 ( .A1(n_800), .A2(n_806), .B1(n_808), .B2(n_812), .C(n_813), .Y(n_799) );
INVx1_ASAP7_75t_L g800 ( .A(n_801), .Y(n_800) );
NAND2xp5_ASAP7_75t_L g801 ( .A(n_802), .B(n_805), .Y(n_801) );
OAI221xp5_ASAP7_75t_L g921 ( .A1(n_802), .A2(n_915), .B1(n_922), .B2(n_926), .C(n_928), .Y(n_921) );
INVx1_ASAP7_75t_L g802 ( .A(n_803), .Y(n_802) );
OAI21xp33_ASAP7_75t_L g872 ( .A1(n_803), .A2(n_873), .B(n_875), .Y(n_872) );
INVx1_ASAP7_75t_L g815 ( .A(n_804), .Y(n_815) );
NAND2xp5_ASAP7_75t_L g860 ( .A(n_804), .B(n_861), .Y(n_860) );
OAI321xp33_ASAP7_75t_L g911 ( .A1(n_805), .A2(n_912), .A3(n_914), .B1(n_915), .B2(n_916), .C(n_917), .Y(n_911) );
INVx3_ASAP7_75t_L g820 ( .A(n_807), .Y(n_820) );
INVx1_ASAP7_75t_L g908 ( .A(n_807), .Y(n_908) );
O2A1O1Ixp33_ASAP7_75t_SL g850 ( .A1(n_808), .A2(n_851), .B(n_853), .C(n_862), .Y(n_850) );
NAND2xp5_ASAP7_75t_L g808 ( .A(n_809), .B(n_811), .Y(n_808) );
NOR2xp33_ASAP7_75t_L g898 ( .A(n_809), .B(n_899), .Y(n_898) );
INVx3_ASAP7_75t_L g809 ( .A(n_810), .Y(n_809) );
INVx1_ASAP7_75t_L g846 ( .A(n_811), .Y(n_846) );
NAND3xp33_ASAP7_75t_L g917 ( .A(n_811), .B(n_822), .C(n_854), .Y(n_917) );
O2A1O1Ixp33_ASAP7_75t_L g813 ( .A1(n_814), .A2(n_817), .B(n_818), .C(n_819), .Y(n_813) );
NOR2xp33_ASAP7_75t_L g814 ( .A(n_815), .B(n_816), .Y(n_814) );
INVx1_ASAP7_75t_L g856 ( .A(n_816), .Y(n_856) );
NOR2xp33_ASAP7_75t_L g834 ( .A(n_817), .B(n_835), .Y(n_834) );
NOR2xp33_ASAP7_75t_L g819 ( .A(n_820), .B(n_821), .Y(n_819) );
NAND2xp5_ASAP7_75t_L g866 ( .A(n_820), .B(n_862), .Y(n_866) );
NAND2xp5_ASAP7_75t_L g897 ( .A(n_820), .B(n_825), .Y(n_897) );
NAND2xp5_ASAP7_75t_L g821 ( .A(n_822), .B(n_823), .Y(n_821) );
CKINVDCx16_ASAP7_75t_R g932 ( .A(n_824), .Y(n_932) );
INVx1_ASAP7_75t_L g824 ( .A(n_825), .Y(n_824) );
BUFx3_ASAP7_75t_L g825 ( .A(n_826), .Y(n_825) );
INVx2_ASAP7_75t_L g862 ( .A(n_826), .Y(n_862) );
NAND5xp2_ASAP7_75t_L g830 ( .A(n_831), .B(n_876), .C(n_889), .D(n_901), .E(n_918), .Y(n_830) );
AOI211xp5_ASAP7_75t_L g831 ( .A1(n_832), .A2(n_833), .B(n_850), .C(n_863), .Y(n_831) );
OAI221xp5_ASAP7_75t_L g833 ( .A1(n_834), .A2(n_837), .B1(n_838), .B2(n_839), .C(n_841), .Y(n_833) );
INVx1_ASAP7_75t_L g839 ( .A(n_840), .Y(n_839) );
AOI21xp5_ASAP7_75t_L g841 ( .A1(n_842), .A2(n_844), .B(n_845), .Y(n_841) );
NOR2xp33_ASAP7_75t_L g878 ( .A(n_844), .B(n_879), .Y(n_878) );
INVx1_ASAP7_75t_L g888 ( .A(n_849), .Y(n_888) );
INVx1_ASAP7_75t_L g924 ( .A(n_852), .Y(n_924) );
OAI21xp33_ASAP7_75t_SL g857 ( .A1(n_858), .A2(n_859), .B(n_860), .Y(n_857) );
INVx1_ASAP7_75t_L g891 ( .A(n_859), .Y(n_891) );
NAND2xp5_ASAP7_75t_L g899 ( .A(n_861), .B(n_900), .Y(n_899) );
CKINVDCx16_ASAP7_75t_R g882 ( .A(n_862), .Y(n_882) );
NOR2xp33_ASAP7_75t_L g887 ( .A(n_862), .B(n_888), .Y(n_887) );
OAI221xp5_ASAP7_75t_L g863 ( .A1(n_864), .A2(n_866), .B1(n_867), .B2(n_869), .C(n_872), .Y(n_863) );
NAND2xp5_ASAP7_75t_L g886 ( .A(n_865), .B(n_887), .Y(n_886) );
INVx1_ASAP7_75t_L g867 ( .A(n_868), .Y(n_867) );
INVx1_ASAP7_75t_L g869 ( .A(n_870), .Y(n_869) );
INVx1_ASAP7_75t_L g873 ( .A(n_874), .Y(n_873) );
INVx1_ASAP7_75t_L g902 ( .A(n_879), .Y(n_902) );
OAI21xp33_ASAP7_75t_L g880 ( .A1(n_881), .A2(n_885), .B(n_886), .Y(n_880) );
AOI211xp5_ASAP7_75t_L g889 ( .A1(n_890), .A2(n_892), .B(n_894), .C(n_898), .Y(n_889) );
A2O1A1Ixp33_ASAP7_75t_L g918 ( .A1(n_890), .A2(n_919), .B(n_921), .C(n_932), .Y(n_918) );
INVx1_ASAP7_75t_L g892 ( .A(n_893), .Y(n_892) );
INVx1_ASAP7_75t_L g903 ( .A(n_897), .Y(n_903) );
AOI221xp5_ASAP7_75t_L g901 ( .A1(n_902), .A2(n_903), .B1(n_904), .B2(n_909), .C(n_911), .Y(n_901) );
INVx1_ASAP7_75t_L g906 ( .A(n_907), .Y(n_906) );
INVx1_ASAP7_75t_L g909 ( .A(n_910), .Y(n_909) );
INVxp67_ASAP7_75t_L g912 ( .A(n_913), .Y(n_912) );
NAND2xp5_ASAP7_75t_L g922 ( .A(n_923), .B(n_925), .Y(n_922) );
INVx1_ASAP7_75t_L g923 ( .A(n_924), .Y(n_923) );
INVx1_ASAP7_75t_L g926 ( .A(n_927), .Y(n_926) );
INVx1_ASAP7_75t_L g928 ( .A(n_929), .Y(n_928) );
INVx1_ASAP7_75t_L g930 ( .A(n_931), .Y(n_930) );
CKINVDCx5p33_ASAP7_75t_R g933 ( .A(n_934), .Y(n_933) );
INVx1_ASAP7_75t_L g934 ( .A(n_935), .Y(n_934) );
INVx2_ASAP7_75t_L g936 ( .A(n_937), .Y(n_936) );
AO21x2_ASAP7_75t_L g937 ( .A1(n_938), .A2(n_939), .B(n_964), .Y(n_937) );
NOR3xp33_ASAP7_75t_L g964 ( .A(n_938), .B(n_941), .C(n_947), .Y(n_964) );
NAND2xp5_ASAP7_75t_L g939 ( .A(n_940), .B(n_946), .Y(n_939) );
INVx1_ASAP7_75t_L g940 ( .A(n_941), .Y(n_940) );
NAND4xp25_ASAP7_75t_SL g941 ( .A(n_942), .B(n_943), .C(n_944), .D(n_945), .Y(n_941) );
INVx1_ASAP7_75t_L g946 ( .A(n_947), .Y(n_946) );
NAND3xp33_ASAP7_75t_L g947 ( .A(n_948), .B(n_950), .C(n_955), .Y(n_947) );
INVx2_ASAP7_75t_L g951 ( .A(n_952), .Y(n_951) );
BUFx3_ASAP7_75t_L g953 ( .A(n_954), .Y(n_953) );
INVx1_ASAP7_75t_L g1002 ( .A(n_956), .Y(n_1002) );
INVx2_ASAP7_75t_L g956 ( .A(n_957), .Y(n_956) );
OAI21xp5_ASAP7_75t_SL g958 ( .A1(n_959), .A2(n_961), .B(n_962), .Y(n_958) );
INVxp67_ASAP7_75t_L g959 ( .A(n_960), .Y(n_959) );
INVx1_ASAP7_75t_L g965 ( .A(n_966), .Y(n_965) );
HB1xp67_ASAP7_75t_L g966 ( .A(n_967), .Y(n_966) );
INVx1_ASAP7_75t_L g1004 ( .A(n_973), .Y(n_1004) );
HB1xp67_ASAP7_75t_L g973 ( .A(n_974), .Y(n_973) );
NAND4xp75_ASAP7_75t_L g974 ( .A(n_975), .B(n_981), .C(n_990), .D(n_999), .Y(n_974) );
AND2x2_ASAP7_75t_L g975 ( .A(n_976), .B(n_979), .Y(n_975) );
BUFx2_ASAP7_75t_L g977 ( .A(n_978), .Y(n_977) );
NOR2x1_ASAP7_75t_L g981 ( .A(n_982), .B(n_986), .Y(n_981) );
AND2x2_ASAP7_75t_L g990 ( .A(n_991), .B(n_995), .Y(n_990) );
INVx1_ASAP7_75t_L g992 ( .A(n_993), .Y(n_992) );
BUFx4f_ASAP7_75t_L g996 ( .A(n_997), .Y(n_996) );
INVx1_ASAP7_75t_L g999 ( .A(n_1000), .Y(n_999) );
OAI21xp33_ASAP7_75t_L g1000 ( .A1(n_1001), .A2(n_1002), .B(n_1003), .Y(n_1000) );
HB1xp67_ASAP7_75t_L g1005 ( .A(n_1006), .Y(n_1005) );
HB1xp67_ASAP7_75t_L g1007 ( .A(n_1008), .Y(n_1007) );
endmodule