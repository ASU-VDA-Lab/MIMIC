module real_jpeg_1900_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_384;
wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_128;
wire n_216;
wire n_202;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_393;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_372;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_286;
wire n_166;
wire n_215;
wire n_176;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_330;
wire n_298;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;
wire n_364;

INVx2_ASAP7_75t_L g111 ( 
.A(n_0),
.Y(n_111)
);

BUFx3_ASAP7_75t_L g133 ( 
.A(n_1),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_2),
.B(n_29),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_2),
.B(n_36),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_2),
.B(n_47),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_2),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_2),
.B(n_59),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_2),
.B(n_78),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_3),
.B(n_36),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_3),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_3),
.B(n_29),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_3),
.B(n_47),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_3),
.B(n_59),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_4),
.B(n_29),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_4),
.B(n_47),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_4),
.B(n_59),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_4),
.B(n_36),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_4),
.B(n_78),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_4),
.B(n_109),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_4),
.B(n_133),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_4),
.B(n_24),
.Y(n_318)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_5),
.Y(n_47)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

BUFx10_ASAP7_75t_L g78 ( 
.A(n_7),
.Y(n_78)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_9),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_9),
.B(n_59),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_9),
.B(n_109),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_9),
.B(n_78),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_9),
.B(n_133),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_9),
.B(n_24),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_10),
.B(n_29),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_10),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_10),
.B(n_47),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_10),
.B(n_59),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_10),
.B(n_78),
.Y(n_77)
);

AND2x2_ASAP7_75t_SL g108 ( 
.A(n_10),
.B(n_109),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_10),
.B(n_133),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_10),
.B(n_24),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_11),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_12),
.B(n_24),
.Y(n_23)
);

CKINVDCx14_ASAP7_75t_R g44 ( 
.A(n_12),
.Y(n_44)
);

AND2x2_ASAP7_75t_L g68 ( 
.A(n_12),
.B(n_29),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_12),
.B(n_47),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_12),
.B(n_59),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_12),
.B(n_78),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_12),
.B(n_109),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_12),
.B(n_133),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_13),
.B(n_24),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_13),
.B(n_36),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_13),
.B(n_29),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_13),
.B(n_47),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_13),
.B(n_59),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_13),
.B(n_133),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_13),
.B(n_109),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_13),
.B(n_78),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_14),
.B(n_24),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_14),
.B(n_36),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_14),
.B(n_29),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_14),
.B(n_47),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_14),
.B(n_109),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_14),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_15),
.Y(n_60)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_87),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_86),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_61),
.Y(n_18)
);

OR2x2_ASAP7_75t_L g86 ( 
.A(n_19),
.B(n_61),
.Y(n_86)
);

XOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_48),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_SL g20 ( 
.A1(n_21),
.A2(n_22),
.B1(n_40),
.B2(n_41),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_26),
.B1(n_27),
.B2(n_39),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_23),
.Y(n_39)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_23),
.B(n_72),
.C(n_73),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_23),
.A2(n_39),
.B1(n_126),
.B2(n_128),
.Y(n_125)
);

INVx4_ASAP7_75t_L g158 ( 
.A(n_24),
.Y(n_158)
);

INVx6_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_27),
.Y(n_26)
);

OAI21xp5_ASAP7_75t_L g27 ( 
.A1(n_28),
.A2(n_32),
.B(n_38),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_28),
.B(n_32),
.Y(n_38)
);

MAJIxp5_ASAP7_75t_L g41 ( 
.A(n_28),
.B(n_42),
.C(n_45),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_L g51 ( 
.A1(n_28),
.A2(n_45),
.B1(n_46),
.B2(n_52),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_28),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g328 ( 
.A1(n_28),
.A2(n_52),
.B1(n_329),
.B2(n_330),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_28),
.B(n_330),
.C(n_331),
.Y(n_342)
);

INVx4_ASAP7_75t_L g203 ( 
.A(n_29),
.Y(n_203)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_SL g352 ( 
.A1(n_32),
.A2(n_33),
.B1(n_353),
.B2(n_354),
.Y(n_352)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_33),
.B(n_108),
.C(n_132),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_34),
.B(n_35),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_SL g43 ( 
.A(n_35),
.B(n_44),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_35),
.B(n_166),
.Y(n_314)
);

INVx6_ASAP7_75t_SL g35 ( 
.A(n_36),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_41),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_42),
.A2(n_43),
.B1(n_50),
.B2(n_51),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_42),
.A2(n_43),
.B1(n_123),
.B2(n_124),
.Y(n_122)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_43),
.B(n_100),
.C(n_102),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_45),
.A2(n_46),
.B1(n_57),
.B2(n_58),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_45),
.A2(n_46),
.B1(n_210),
.B2(n_211),
.Y(n_209)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

MAJIxp5_ASAP7_75t_L g54 ( 
.A(n_46),
.B(n_55),
.C(n_57),
.Y(n_54)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_46),
.B(n_101),
.C(n_210),
.Y(n_315)
);

INVx3_ASAP7_75t_SL g165 ( 
.A(n_47),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g48 ( 
.A(n_49),
.B(n_53),
.C(n_54),
.Y(n_48)
);

XNOR2xp5_ASAP7_75t_L g84 ( 
.A(n_49),
.B(n_85),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_51),
.Y(n_50)
);

XNOR2xp5_ASAP7_75t_L g85 ( 
.A(n_53),
.B(n_54),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_55),
.A2(n_56),
.B1(n_81),
.B2(n_82),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_56),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_57),
.A2(n_58),
.B1(n_76),
.B2(n_77),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_L g159 ( 
.A1(n_57),
.A2(n_58),
.B1(n_120),
.B2(n_160),
.Y(n_159)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_58),
.B(n_76),
.C(n_79),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_58),
.B(n_120),
.C(n_156),
.Y(n_200)
);

INVx4_ASAP7_75t_L g311 ( 
.A(n_59),
.Y(n_311)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

MAJIxp5_ASAP7_75t_L g61 ( 
.A(n_62),
.B(n_83),
.C(n_84),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_62),
.A2(n_63),
.B1(n_136),
.B2(n_137),
.Y(n_135)
);

CKINVDCx16_ASAP7_75t_R g62 ( 
.A(n_63),
.Y(n_62)
);

MAJIxp5_ASAP7_75t_L g63 ( 
.A(n_64),
.B(n_75),
.C(n_80),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_64),
.A2(n_65),
.B1(n_93),
.B2(n_94),
.Y(n_92)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

XOR2xp5_ASAP7_75t_L g65 ( 
.A(n_66),
.B(n_71),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_67),
.A2(n_68),
.B1(n_69),
.B2(n_70),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_67),
.B(n_70),
.C(n_71),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g345 ( 
.A1(n_67),
.A2(n_68),
.B1(n_346),
.B2(n_347),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_SL g371 ( 
.A1(n_67),
.A2(n_68),
.B1(n_134),
.B2(n_372),
.Y(n_371)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_68),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_68),
.B(n_130),
.C(n_134),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g368 ( 
.A(n_68),
.B(n_344),
.C(n_347),
.Y(n_368)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_70),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_72),
.A2(n_73),
.B1(n_74),
.B2(n_127),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_72),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_72),
.A2(n_127),
.B1(n_313),
.B2(n_314),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_72),
.B(n_310),
.C(n_314),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_74),
.Y(n_73)
);

XNOR2xp5_ASAP7_75t_SL g93 ( 
.A(n_75),
.B(n_80),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_SL g104 ( 
.A(n_76),
.B(n_105),
.C(n_107),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_76),
.A2(n_77),
.B1(n_107),
.B2(n_108),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_76),
.A2(n_77),
.B1(n_181),
.B2(n_187),
.Y(n_186)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_77),
.B(n_181),
.C(n_182),
.Y(n_180)
);

INVx13_ASAP7_75t_L g205 ( 
.A(n_78),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g97 ( 
.A(n_79),
.B(n_98),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_82),
.Y(n_81)
);

XNOR2xp5_ASAP7_75t_SL g136 ( 
.A(n_83),
.B(n_84),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_L g87 ( 
.A1(n_88),
.A2(n_138),
.B(n_402),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_135),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g403 ( 
.A(n_90),
.B(n_135),
.Y(n_403)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_95),
.C(n_112),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g387 ( 
.A1(n_91),
.A2(n_92),
.B1(n_95),
.B2(n_388),
.Y(n_387)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_93),
.Y(n_94)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_95),
.Y(n_388)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_99),
.C(n_104),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g392 ( 
.A1(n_96),
.A2(n_97),
.B1(n_393),
.B2(n_394),
.Y(n_392)
);

CKINVDCx16_ASAP7_75t_R g96 ( 
.A(n_97),
.Y(n_96)
);

XNOR2xp5_ASAP7_75t_SL g393 ( 
.A(n_99),
.B(n_104),
.Y(n_393)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_100),
.A2(n_101),
.B1(n_102),
.B2(n_103),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_100),
.A2(n_101),
.B1(n_208),
.B2(n_209),
.Y(n_207)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_105),
.A2(n_106),
.B1(n_116),
.B2(n_117),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_106),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_107),
.A2(n_108),
.B1(n_220),
.B2(n_223),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g353 ( 
.A1(n_107),
.A2(n_108),
.B1(n_132),
.B2(n_244),
.Y(n_353)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_108),
.Y(n_107)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_110),
.B(n_225),
.Y(n_266)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

XNOR2xp5_ASAP7_75t_L g386 ( 
.A(n_112),
.B(n_387),
.Y(n_386)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_125),
.C(n_129),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_SL g390 ( 
.A(n_113),
.B(n_391),
.Y(n_390)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_118),
.C(n_122),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g363 ( 
.A1(n_114),
.A2(n_115),
.B1(n_364),
.B2(n_365),
.Y(n_363)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

CKINVDCx14_ASAP7_75t_R g116 ( 
.A(n_117),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_SL g364 ( 
.A(n_118),
.B(n_122),
.Y(n_364)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_120),
.C(n_121),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_SL g358 ( 
.A(n_119),
.B(n_121),
.Y(n_358)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_120),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g357 ( 
.A1(n_120),
.A2(n_160),
.B1(n_358),
.B2(n_359),
.Y(n_357)
);

CKINVDCx16_ASAP7_75t_R g123 ( 
.A(n_124),
.Y(n_123)
);

XNOR2xp5_ASAP7_75t_L g391 ( 
.A(n_125),
.B(n_129),
.Y(n_391)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_126),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g369 ( 
.A1(n_130),
.A2(n_131),
.B1(n_370),
.B2(n_371),
.Y(n_369)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_132),
.B(n_148),
.Y(n_147)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_132),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_132),
.A2(n_242),
.B1(n_243),
.B2(n_244),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_132),
.A2(n_148),
.B1(n_178),
.B2(n_244),
.Y(n_317)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_133),
.Y(n_176)
);

CKINVDCx16_ASAP7_75t_R g372 ( 
.A(n_134),
.Y(n_372)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_136),
.Y(n_137)
);

AOI21xp5_ASAP7_75t_L g138 ( 
.A1(n_139),
.A2(n_384),
.B(n_399),
.Y(n_138)
);

OAI31xp33_ASAP7_75t_L g139 ( 
.A1(n_140),
.A2(n_334),
.A3(n_373),
.B(n_378),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_141),
.B(n_302),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_226),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_194),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_143),
.B(n_194),
.Y(n_380)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_161),
.C(n_184),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_144),
.B(n_299),
.Y(n_298)
);

BUFx24_ASAP7_75t_SL g407 ( 
.A(n_144),
.Y(n_407)
);

FAx1_ASAP7_75t_SL g144 ( 
.A(n_145),
.B(n_151),
.CI(n_155),
.CON(n_144),
.SN(n_144)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_145),
.B(n_151),
.C(n_155),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_149),
.C(n_150),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_146),
.A2(n_147),
.B1(n_294),
.B2(n_295),
.Y(n_293)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

O2A1O1Ixp33_ASAP7_75t_L g356 ( 
.A1(n_147),
.A2(n_178),
.B(n_244),
.C(n_318),
.Y(n_356)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_148),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_148),
.A2(n_175),
.B1(n_178),
.B2(n_193),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_SL g295 ( 
.A(n_149),
.B(n_150),
.Y(n_295)
);

OAI21xp5_ASAP7_75t_L g151 ( 
.A1(n_152),
.A2(n_153),
.B(n_154),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_152),
.B(n_153),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_154),
.A2(n_215),
.B1(n_216),
.B2(n_217),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_154),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_159),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_158),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_157),
.B(n_176),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_157),
.B(n_205),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_158),
.B(n_225),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_161),
.B(n_184),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_162),
.A2(n_163),
.B1(n_172),
.B2(n_183),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_162),
.B(n_173),
.C(n_180),
.Y(n_196)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_167),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_164),
.B(n_169),
.C(n_171),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_166),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_166),
.B(n_203),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_168),
.A2(n_169),
.B1(n_170),
.B2(n_171),
.Y(n_167)
);

CKINVDCx16_ASAP7_75t_R g171 ( 
.A(n_168),
.Y(n_171)
);

CKINVDCx14_ASAP7_75t_R g169 ( 
.A(n_170),
.Y(n_169)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_172),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_173),
.A2(n_174),
.B1(n_179),
.B2(n_180),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_178),
.Y(n_174)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_175),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_177),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_177),
.B(n_205),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_177),
.B(n_311),
.Y(n_310)
);

CKINVDCx16_ASAP7_75t_R g179 ( 
.A(n_180),
.Y(n_179)
);

INVxp67_ASAP7_75t_L g187 ( 
.A(n_181),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_182),
.B(n_186),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_188),
.C(n_192),
.Y(n_184)
);

FAx1_ASAP7_75t_SL g289 ( 
.A(n_185),
.B(n_188),
.CI(n_192),
.CON(n_289),
.SN(n_289)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_190),
.C(n_191),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_189),
.B(n_191),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_190),
.B(n_237),
.Y(n_236)
);

BUFx24_ASAP7_75t_SL g410 ( 
.A(n_194),
.Y(n_410)
);

FAx1_ASAP7_75t_SL g194 ( 
.A(n_195),
.B(n_212),
.CI(n_213),
.CON(n_194),
.SN(n_194)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_195),
.B(n_212),
.C(n_213),
.Y(n_333)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_197),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_196),
.B(n_199),
.C(n_206),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_198),
.A2(n_199),
.B1(n_206),
.B2(n_207),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_201),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_200),
.B(n_202),
.C(n_204),
.Y(n_325)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_204),
.Y(n_201)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

CKINVDCx16_ASAP7_75t_R g211 ( 
.A(n_210),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_218),
.Y(n_213)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_215),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_215),
.B(n_216),
.C(n_218),
.Y(n_322)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_224),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_220),
.A2(n_221),
.B1(n_222),
.B2(n_223),
.Y(n_219)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_220),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_220),
.B(n_222),
.C(n_224),
.Y(n_332)
);

CKINVDCx16_ASAP7_75t_R g221 ( 
.A(n_222),
.Y(n_221)
);

AOI21xp5_ASAP7_75t_SL g226 ( 
.A1(n_227),
.A2(n_297),
.B(n_301),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_SL g227 ( 
.A1(n_228),
.A2(n_285),
.B(n_296),
.Y(n_227)
);

AOI21xp5_ASAP7_75t_L g228 ( 
.A1(n_229),
.A2(n_257),
.B(n_284),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_230),
.B(n_248),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_230),
.B(n_248),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_240),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_232),
.A2(n_236),
.B1(n_238),
.B2(n_239),
.Y(n_231)
);

CKINVDCx14_ASAP7_75t_R g238 ( 
.A(n_232),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_234),
.C(n_235),
.Y(n_232)
);

FAx1_ASAP7_75t_SL g249 ( 
.A(n_233),
.B(n_234),
.CI(n_235),
.CON(n_249),
.SN(n_249)
);

CKINVDCx16_ASAP7_75t_R g239 ( 
.A(n_236),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_236),
.B(n_238),
.C(n_240),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_SL g240 ( 
.A(n_241),
.B(n_245),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_241),
.B(n_246),
.C(n_247),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_242),
.B(n_244),
.Y(n_241)
);

CKINVDCx16_ASAP7_75t_R g242 ( 
.A(n_243),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_247),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_250),
.C(n_256),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_249),
.B(n_281),
.Y(n_280)
);

BUFx24_ASAP7_75t_SL g405 ( 
.A(n_249),
.Y(n_405)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_250),
.A2(n_251),
.B1(n_256),
.B2(n_282),
.Y(n_281)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_254),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_252),
.A2(n_253),
.B1(n_254),
.B2(n_255),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_253),
.Y(n_252)
);

CKINVDCx16_ASAP7_75t_R g254 ( 
.A(n_255),
.Y(n_254)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_256),
.Y(n_282)
);

OAI21xp5_ASAP7_75t_L g257 ( 
.A1(n_258),
.A2(n_278),
.B(n_283),
.Y(n_257)
);

AOI21xp5_ASAP7_75t_L g258 ( 
.A1(n_259),
.A2(n_269),
.B(n_277),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_260),
.B(n_265),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_260),
.B(n_265),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_264),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_263),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_262),
.B(n_263),
.C(n_264),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_266),
.B(n_267),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_266),
.B(n_271),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_L g274 ( 
.A1(n_266),
.A2(n_267),
.B1(n_268),
.B2(n_275),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_266),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_268),
.Y(n_267)
);

OAI21xp5_ASAP7_75t_L g269 ( 
.A1(n_270),
.A2(n_272),
.B(n_276),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_273),
.B(n_274),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_273),
.B(n_274),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_279),
.B(n_280),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_279),
.B(n_280),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_286),
.B(n_287),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_SL g296 ( 
.A(n_286),
.B(n_287),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_288),
.A2(n_289),
.B1(n_290),
.B2(n_291),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_288),
.B(n_292),
.C(n_293),
.Y(n_300)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

BUFx24_ASAP7_75t_SL g409 ( 
.A(n_289),
.Y(n_409)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

XOR2xp5_ASAP7_75t_L g291 ( 
.A(n_292),
.B(n_293),
.Y(n_291)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_SL g297 ( 
.A(n_298),
.B(n_300),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_298),
.B(n_300),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

OAI21xp5_ASAP7_75t_L g379 ( 
.A1(n_303),
.A2(n_380),
.B(n_381),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_SL g303 ( 
.A(n_304),
.B(n_333),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_304),
.B(n_333),
.Y(n_381)
);

XNOR2xp5_ASAP7_75t_L g304 ( 
.A(n_305),
.B(n_306),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g377 ( 
.A(n_305),
.B(n_307),
.C(n_320),
.Y(n_377)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_307),
.A2(n_308),
.B1(n_319),
.B2(n_320),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

BUFx24_ASAP7_75t_SL g406 ( 
.A(n_308),
.Y(n_406)
);

FAx1_ASAP7_75t_SL g308 ( 
.A(n_309),
.B(n_315),
.CI(n_316),
.CON(n_308),
.SN(n_308)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_309),
.B(n_315),
.C(n_316),
.Y(n_340)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_310),
.B(n_312),
.Y(n_309)
);

INVxp67_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_SL g316 ( 
.A(n_317),
.B(n_318),
.Y(n_316)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_L g320 ( 
.A1(n_321),
.A2(n_322),
.B1(n_323),
.B2(n_324),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g349 ( 
.A(n_321),
.B(n_325),
.C(n_326),
.Y(n_349)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_SL g324 ( 
.A(n_325),
.B(n_326),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_L g326 ( 
.A1(n_327),
.A2(n_328),
.B1(n_331),
.B2(n_332),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_330),
.Y(n_329)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_332),
.Y(n_331)
);

INVxp33_ASAP7_75t_L g334 ( 
.A(n_335),
.Y(n_334)
);

A2O1A1O1Ixp25_ASAP7_75t_SL g378 ( 
.A1(n_335),
.A2(n_374),
.B(n_379),
.C(n_382),
.D(n_383),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_336),
.B(n_360),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g383 ( 
.A(n_336),
.B(n_360),
.Y(n_383)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_337),
.B(n_349),
.C(n_350),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_L g376 ( 
.A1(n_337),
.A2(n_338),
.B1(n_350),
.B2(n_351),
.Y(n_376)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_338),
.Y(n_337)
);

AOI22xp5_ASAP7_75t_L g338 ( 
.A1(n_339),
.A2(n_340),
.B1(n_341),
.B2(n_348),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g361 ( 
.A(n_339),
.B(n_342),
.C(n_343),
.Y(n_361)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_340),
.Y(n_339)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_341),
.Y(n_348)
);

XNOR2xp5_ASAP7_75t_SL g341 ( 
.A(n_342),
.B(n_343),
.Y(n_341)
);

XOR2xp5_ASAP7_75t_L g343 ( 
.A(n_344),
.B(n_345),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g347 ( 
.A(n_346),
.Y(n_347)
);

XOR2xp5_ASAP7_75t_L g375 ( 
.A(n_349),
.B(n_376),
.Y(n_375)
);

CKINVDCx14_ASAP7_75t_R g350 ( 
.A(n_351),
.Y(n_350)
);

XNOR2xp5_ASAP7_75t_SL g351 ( 
.A(n_352),
.B(n_355),
.Y(n_351)
);

MAJIxp5_ASAP7_75t_L g367 ( 
.A(n_352),
.B(n_356),
.C(n_357),
.Y(n_367)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_353),
.Y(n_354)
);

XNOR2xp5_ASAP7_75t_L g355 ( 
.A(n_356),
.B(n_357),
.Y(n_355)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_358),
.Y(n_359)
);

XNOR2xp5_ASAP7_75t_L g360 ( 
.A(n_361),
.B(n_362),
.Y(n_360)
);

MAJIxp5_ASAP7_75t_L g398 ( 
.A(n_361),
.B(n_363),
.C(n_366),
.Y(n_398)
);

XNOR2xp5_ASAP7_75t_L g362 ( 
.A(n_363),
.B(n_366),
.Y(n_362)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_364),
.Y(n_365)
);

BUFx24_ASAP7_75t_SL g411 ( 
.A(n_366),
.Y(n_411)
);

FAx1_ASAP7_75t_SL g366 ( 
.A(n_367),
.B(n_368),
.CI(n_369),
.CON(n_366),
.SN(n_366)
);

MAJIxp5_ASAP7_75t_L g395 ( 
.A(n_367),
.B(n_368),
.C(n_369),
.Y(n_395)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_371),
.Y(n_370)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_374),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_SL g374 ( 
.A(n_375),
.B(n_377),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_L g382 ( 
.A(n_375),
.B(n_377),
.Y(n_382)
);

NOR2xp33_ASAP7_75t_L g384 ( 
.A(n_385),
.B(n_396),
.Y(n_384)
);

OAI21xp5_ASAP7_75t_L g399 ( 
.A1(n_385),
.A2(n_400),
.B(n_401),
.Y(n_399)
);

NOR2xp33_ASAP7_75t_SL g385 ( 
.A(n_386),
.B(n_389),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_386),
.B(n_389),
.Y(n_401)
);

MAJIxp5_ASAP7_75t_L g389 ( 
.A(n_390),
.B(n_392),
.C(n_395),
.Y(n_389)
);

FAx1_ASAP7_75t_SL g397 ( 
.A(n_390),
.B(n_392),
.CI(n_395),
.CON(n_397),
.SN(n_397)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_393),
.Y(n_394)
);

NOR2xp33_ASAP7_75t_SL g396 ( 
.A(n_397),
.B(n_398),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_397),
.B(n_398),
.Y(n_400)
);

BUFx24_ASAP7_75t_SL g404 ( 
.A(n_397),
.Y(n_404)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_403),
.Y(n_402)
);


endmodule