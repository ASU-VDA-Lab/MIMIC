module fake_netlist_5_1719_n_1110 (n_137, n_210, n_168, n_260, n_164, n_191, n_91, n_208, n_82, n_122, n_194, n_142, n_176, n_10, n_214, n_140, n_24, n_248, n_124, n_86, n_136, n_146, n_268, n_182, n_143, n_83, n_132, n_61, n_237, n_90, n_241, n_127, n_75, n_101, n_180, n_184, n_226, n_235, n_65, n_78, n_74, n_144, n_207, n_240, n_114, n_57, n_96, n_37, n_189, n_220, n_165, n_111, n_229, n_108, n_231, n_257, n_213, n_129, n_31, n_13, n_66, n_98, n_177, n_60, n_155, n_152, n_197, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_236, n_18, n_116, n_195, n_42, n_22, n_227, n_1, n_45, n_117, n_249, n_271, n_46, n_233, n_21, n_94, n_203, n_245, n_205, n_113, n_38, n_123, n_139, n_105, n_246, n_80, n_4, n_179, n_125, n_35, n_269, n_167, n_128, n_73, n_234, n_17, n_92, n_19, n_267, n_149, n_120, n_232, n_135, n_30, n_156, n_5, n_33, n_126, n_254, n_14, n_225, n_84, n_23, n_202, n_130, n_266, n_272, n_219, n_157, n_258, n_265, n_29, n_79, n_193, n_131, n_151, n_47, n_173, n_192, n_244, n_251, n_25, n_53, n_160, n_198, n_223, n_247, n_188, n_190, n_8, n_201, n_158, n_263, n_44, n_224, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_228, n_264, n_109, n_112, n_212, n_85, n_159, n_163, n_95, n_119, n_183, n_185, n_243, n_239, n_175, n_252, n_169, n_59, n_262, n_26, n_255, n_133, n_238, n_215, n_55, n_196, n_99, n_2, n_211, n_218, n_181, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_178, n_221, n_12, n_67, n_121, n_242, n_36, n_76, n_200, n_87, n_150, n_162, n_27, n_170, n_64, n_77, n_102, n_106, n_161, n_209, n_259, n_273, n_270, n_222, n_230, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_253, n_261, n_72, n_174, n_186, n_199, n_134, n_187, n_32, n_41, n_104, n_172, n_103, n_56, n_51, n_63, n_97, n_141, n_166, n_11, n_206, n_217, n_171, n_153, n_7, n_15, n_145, n_256, n_48, n_204, n_50, n_250, n_52, n_88, n_110, n_216, n_1110);

input n_137;
input n_210;
input n_168;
input n_260;
input n_164;
input n_191;
input n_91;
input n_208;
input n_82;
input n_122;
input n_194;
input n_142;
input n_176;
input n_10;
input n_214;
input n_140;
input n_24;
input n_248;
input n_124;
input n_86;
input n_136;
input n_146;
input n_268;
input n_182;
input n_143;
input n_83;
input n_132;
input n_61;
input n_237;
input n_90;
input n_241;
input n_127;
input n_75;
input n_101;
input n_180;
input n_184;
input n_226;
input n_235;
input n_65;
input n_78;
input n_74;
input n_144;
input n_207;
input n_240;
input n_114;
input n_57;
input n_96;
input n_37;
input n_189;
input n_220;
input n_165;
input n_111;
input n_229;
input n_108;
input n_231;
input n_257;
input n_213;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_177;
input n_60;
input n_155;
input n_152;
input n_197;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_236;
input n_18;
input n_116;
input n_195;
input n_42;
input n_22;
input n_227;
input n_1;
input n_45;
input n_117;
input n_249;
input n_271;
input n_46;
input n_233;
input n_21;
input n_94;
input n_203;
input n_245;
input n_205;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_246;
input n_80;
input n_4;
input n_179;
input n_125;
input n_35;
input n_269;
input n_167;
input n_128;
input n_73;
input n_234;
input n_17;
input n_92;
input n_19;
input n_267;
input n_149;
input n_120;
input n_232;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_254;
input n_14;
input n_225;
input n_84;
input n_23;
input n_202;
input n_130;
input n_266;
input n_272;
input n_219;
input n_157;
input n_258;
input n_265;
input n_29;
input n_79;
input n_193;
input n_131;
input n_151;
input n_47;
input n_173;
input n_192;
input n_244;
input n_251;
input n_25;
input n_53;
input n_160;
input n_198;
input n_223;
input n_247;
input n_188;
input n_190;
input n_8;
input n_201;
input n_158;
input n_263;
input n_44;
input n_224;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_228;
input n_264;
input n_109;
input n_112;
input n_212;
input n_85;
input n_159;
input n_163;
input n_95;
input n_119;
input n_183;
input n_185;
input n_243;
input n_239;
input n_175;
input n_252;
input n_169;
input n_59;
input n_262;
input n_26;
input n_255;
input n_133;
input n_238;
input n_215;
input n_55;
input n_196;
input n_99;
input n_2;
input n_211;
input n_218;
input n_181;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_178;
input n_221;
input n_12;
input n_67;
input n_121;
input n_242;
input n_36;
input n_76;
input n_200;
input n_87;
input n_150;
input n_162;
input n_27;
input n_170;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_209;
input n_259;
input n_273;
input n_270;
input n_222;
input n_230;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_253;
input n_261;
input n_72;
input n_174;
input n_186;
input n_199;
input n_134;
input n_187;
input n_32;
input n_41;
input n_104;
input n_172;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_166;
input n_11;
input n_206;
input n_217;
input n_171;
input n_153;
input n_7;
input n_15;
input n_145;
input n_256;
input n_48;
input n_204;
input n_50;
input n_250;
input n_52;
input n_88;
input n_110;
input n_216;

output n_1110;

wire n_924;
wire n_676;
wire n_294;
wire n_431;
wire n_318;
wire n_380;
wire n_419;
wire n_977;
wire n_653;
wire n_611;
wire n_444;
wire n_642;
wire n_469;
wire n_615;
wire n_851;
wire n_1060;
wire n_316;
wire n_785;
wire n_389;
wire n_843;
wire n_855;
wire n_549;
wire n_684;
wire n_850;
wire n_418;
wire n_523;
wire n_315;
wire n_451;
wire n_532;
wire n_705;
wire n_619;
wire n_408;
wire n_865;
wire n_913;
wire n_678;
wire n_664;
wire n_376;
wire n_697;
wire n_503;
wire n_967;
wire n_605;
wire n_776;
wire n_928;
wire n_667;
wire n_515;
wire n_790;
wire n_353;
wire n_351;
wire n_367;
wire n_620;
wire n_643;
wire n_1055;
wire n_916;
wire n_452;
wire n_885;
wire n_1081;
wire n_525;
wire n_397;
wire n_493;
wire n_880;
wire n_703;
wire n_698;
wire n_980;
wire n_483;
wire n_544;
wire n_683;
wire n_1007;
wire n_780;
wire n_649;
wire n_552;
wire n_1057;
wire n_1051;
wire n_547;
wire n_1066;
wire n_1085;
wire n_721;
wire n_998;
wire n_841;
wire n_1050;
wire n_1099;
wire n_956;
wire n_564;
wire n_467;
wire n_802;
wire n_423;
wire n_840;
wire n_501;
wire n_284;
wire n_823;
wire n_725;
wire n_983;
wire n_280;
wire n_744;
wire n_1021;
wire n_629;
wire n_590;
wire n_672;
wire n_873;
wire n_378;
wire n_551;
wire n_762;
wire n_581;
wire n_688;
wire n_382;
wire n_554;
wire n_800;
wire n_898;
wire n_690;
wire n_1013;
wire n_583;
wire n_671;
wire n_718;
wire n_819;
wire n_302;
wire n_1022;
wire n_526;
wire n_915;
wire n_719;
wire n_293;
wire n_443;
wire n_372;
wire n_677;
wire n_859;
wire n_864;
wire n_951;
wire n_821;
wire n_714;
wire n_447;
wire n_368;
wire n_433;
wire n_314;
wire n_604;
wire n_321;
wire n_292;
wire n_909;
wire n_625;
wire n_854;
wire n_949;
wire n_621;
wire n_753;
wire n_997;
wire n_455;
wire n_674;
wire n_1048;
wire n_932;
wire n_417;
wire n_946;
wire n_1008;
wire n_612;
wire n_1001;
wire n_385;
wire n_498;
wire n_516;
wire n_933;
wire n_788;
wire n_507;
wire n_497;
wire n_689;
wire n_738;
wire n_912;
wire n_606;
wire n_559;
wire n_275;
wire n_640;
wire n_968;
wire n_624;
wire n_825;
wire n_295;
wire n_1010;
wire n_330;
wire n_877;
wire n_508;
wire n_739;
wire n_506;
wire n_737;
wire n_610;
wire n_972;
wire n_692;
wire n_986;
wire n_755;
wire n_509;
wire n_568;
wire n_936;
wire n_373;
wire n_820;
wire n_757;
wire n_947;
wire n_1090;
wire n_307;
wire n_633;
wire n_439;
wire n_530;
wire n_1024;
wire n_556;
wire n_1063;
wire n_1107;
wire n_448;
wire n_758;
wire n_999;
wire n_668;
wire n_733;
wire n_991;
wire n_375;
wire n_301;
wire n_828;
wire n_779;
wire n_576;
wire n_1032;
wire n_929;
wire n_981;
wire n_941;
wire n_804;
wire n_867;
wire n_537;
wire n_902;
wire n_587;
wire n_945;
wire n_659;
wire n_492;
wire n_792;
wire n_1104;
wire n_563;
wire n_756;
wire n_878;
wire n_524;
wire n_943;
wire n_399;
wire n_579;
wire n_394;
wire n_341;
wire n_992;
wire n_1049;
wire n_938;
wire n_1098;
wire n_741;
wire n_548;
wire n_543;
wire n_1068;
wire n_812;
wire n_842;
wire n_298;
wire n_650;
wire n_984;
wire n_320;
wire n_694;
wire n_518;
wire n_505;
wire n_286;
wire n_883;
wire n_282;
wire n_752;
wire n_331;
wire n_906;
wire n_905;
wire n_519;
wire n_406;
wire n_470;
wire n_919;
wire n_782;
wire n_908;
wire n_1108;
wire n_449;
wire n_325;
wire n_1073;
wire n_1100;
wire n_862;
wire n_900;
wire n_724;
wire n_856;
wire n_546;
wire n_1016;
wire n_760;
wire n_658;
wire n_281;
wire n_918;
wire n_942;
wire n_381;
wire n_291;
wire n_390;
wire n_731;
wire n_456;
wire n_371;
wire n_1077;
wire n_959;
wire n_481;
wire n_535;
wire n_709;
wire n_540;
wire n_317;
wire n_618;
wire n_940;
wire n_896;
wire n_323;
wire n_569;
wire n_769;
wire n_356;
wire n_592;
wire n_920;
wire n_894;
wire n_1046;
wire n_934;
wire n_1017;
wire n_831;
wire n_826;
wire n_335;
wire n_886;
wire n_978;
wire n_964;
wire n_1054;
wire n_654;
wire n_370;
wire n_976;
wire n_1095;
wire n_1096;
wire n_343;
wire n_308;
wire n_379;
wire n_428;
wire n_514;
wire n_457;
wire n_570;
wire n_833;
wire n_297;
wire n_1045;
wire n_1079;
wire n_853;
wire n_603;
wire n_377;
wire n_1078;
wire n_751;
wire n_484;
wire n_775;
wire n_1033;
wire n_988;
wire n_442;
wire n_814;
wire n_636;
wire n_786;
wire n_1083;
wire n_600;
wire n_660;
wire n_392;
wire n_655;
wire n_704;
wire n_787;
wire n_1009;
wire n_669;
wire n_472;
wire n_750;
wire n_742;
wire n_454;
wire n_961;
wire n_995;
wire n_955;
wire n_387;
wire n_771;
wire n_374;
wire n_276;
wire n_339;
wire n_882;
wire n_398;
wire n_396;
wire n_1036;
wire n_635;
wire n_1097;
wire n_347;
wire n_763;
wire n_522;
wire n_550;
wire n_696;
wire n_897;
wire n_350;
wire n_798;
wire n_662;
wire n_459;
wire n_1020;
wire n_646;
wire n_1062;
wire n_400;
wire n_930;
wire n_436;
wire n_962;
wire n_290;
wire n_580;
wire n_622;
wire n_1040;
wire n_1087;
wire n_723;
wire n_1065;
wire n_1035;
wire n_386;
wire n_578;
wire n_994;
wire n_926;
wire n_287;
wire n_344;
wire n_848;
wire n_555;
wire n_783;
wire n_473;
wire n_422;
wire n_475;
wire n_777;
wire n_1070;
wire n_1030;
wire n_661;
wire n_682;
wire n_415;
wire n_485;
wire n_1043;
wire n_1071;
wire n_496;
wire n_355;
wire n_958;
wire n_849;
wire n_1034;
wire n_486;
wire n_670;
wire n_816;
wire n_336;
wire n_584;
wire n_681;
wire n_591;
wire n_922;
wire n_521;
wire n_614;
wire n_663;
wire n_845;
wire n_430;
wire n_337;
wire n_313;
wire n_631;
wire n_673;
wire n_837;
wire n_528;
wire n_479;
wire n_510;
wire n_680;
wire n_974;
wire n_432;
wire n_553;
wire n_395;
wire n_727;
wire n_839;
wire n_901;
wire n_311;
wire n_813;
wire n_957;
wire n_830;
wire n_773;
wire n_743;
wire n_328;
wire n_801;
wire n_299;
wire n_303;
wire n_369;
wire n_675;
wire n_888;
wire n_296;
wire n_613;
wire n_871;
wire n_637;
wire n_357;
wire n_875;
wire n_598;
wire n_685;
wire n_608;
wire n_446;
wire n_445;
wire n_749;
wire n_829;
wire n_858;
wire n_1064;
wire n_923;
wire n_772;
wire n_691;
wire n_881;
wire n_717;
wire n_468;
wire n_499;
wire n_939;
wire n_342;
wire n_517;
wire n_482;
wire n_1088;
wire n_588;
wire n_361;
wire n_464;
wire n_789;
wire n_363;
wire n_402;
wire n_413;
wire n_734;
wire n_638;
wire n_1086;
wire n_700;
wire n_796;
wire n_573;
wire n_866;
wire n_1069;
wire n_1075;
wire n_969;
wire n_388;
wire n_761;
wire n_1012;
wire n_1019;
wire n_1105;
wire n_903;
wire n_1006;
wire n_740;
wire n_304;
wire n_329;
wire n_274;
wire n_577;
wire n_384;
wire n_582;
wire n_460;
wire n_889;
wire n_973;
wire n_277;
wire n_1061;
wire n_477;
wire n_571;
wire n_461;
wire n_338;
wire n_333;
wire n_693;
wire n_309;
wire n_512;
wire n_836;
wire n_990;
wire n_462;
wire n_975;
wire n_322;
wire n_567;
wire n_652;
wire n_778;
wire n_306;
wire n_907;
wire n_722;
wire n_1093;
wire n_458;
wire n_288;
wire n_770;
wire n_844;
wire n_1031;
wire n_471;
wire n_609;
wire n_852;
wire n_989;
wire n_1041;
wire n_1039;
wire n_1102;
wire n_283;
wire n_1028;
wire n_383;
wire n_711;
wire n_781;
wire n_834;
wire n_474;
wire n_765;
wire n_542;
wire n_488;
wire n_463;
wire n_595;
wire n_736;
wire n_502;
wire n_892;
wire n_893;
wire n_1015;
wire n_1000;
wire n_891;
wire n_466;
wire n_420;
wire n_630;
wire n_489;
wire n_632;
wire n_699;
wire n_979;
wire n_1002;
wire n_617;
wire n_310;
wire n_593;
wire n_504;
wire n_511;
wire n_748;
wire n_586;
wire n_846;
wire n_874;
wire n_465;
wire n_838;
wire n_358;
wire n_1058;
wire n_362;
wire n_876;
wire n_332;
wire n_1053;
wire n_1101;
wire n_585;
wire n_349;
wire n_1106;
wire n_616;
wire n_953;
wire n_601;
wire n_279;
wire n_917;
wire n_1014;
wire n_966;
wire n_987;
wire n_289;
wire n_745;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_767;
wire n_993;
wire n_440;
wire n_726;
wire n_478;
wire n_793;
wire n_545;
wire n_982;
wire n_441;
wire n_860;
wire n_1103;
wire n_450;
wire n_648;
wire n_312;
wire n_476;
wire n_818;
wire n_429;
wire n_861;
wire n_534;
wire n_948;
wire n_1076;
wire n_884;
wire n_899;
wire n_345;
wire n_944;
wire n_1091;
wire n_494;
wire n_641;
wire n_628;
wire n_365;
wire n_774;
wire n_730;
wire n_729;
wire n_1059;
wire n_1084;
wire n_970;
wire n_911;
wire n_557;
wire n_1005;
wire n_354;
wire n_575;
wire n_647;
wire n_480;
wire n_607;
wire n_425;
wire n_513;
wire n_407;
wire n_527;
wire n_679;
wire n_707;
wire n_710;
wire n_795;
wire n_695;
wire n_832;
wire n_857;
wire n_560;
wire n_656;
wire n_340;
wire n_1094;
wire n_561;
wire n_1044;
wire n_346;
wire n_937;
wire n_393;
wire n_495;
wire n_487;
wire n_602;
wire n_665;
wire n_574;
wire n_437;
wire n_453;
wire n_403;
wire n_421;
wire n_879;
wire n_1072;
wire n_720;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_863;
wire n_910;
wire n_971;
wire n_490;
wire n_805;
wire n_1027;
wire n_326;
wire n_794;
wire n_768;
wire n_921;
wire n_996;
wire n_404;
wire n_686;
wire n_572;
wire n_366;
wire n_712;
wire n_847;
wire n_754;
wire n_815;
wire n_596;
wire n_410;
wire n_1042;
wire n_558;
wire n_708;
wire n_529;
wire n_735;
wire n_702;
wire n_285;
wire n_822;
wire n_412;
wire n_327;
wire n_1109;
wire n_657;
wire n_644;
wire n_728;
wire n_895;
wire n_1037;
wire n_1080;
wire n_491;
wire n_1074;
wire n_427;
wire n_791;
wire n_732;
wire n_352;
wire n_566;
wire n_565;
wire n_426;
wire n_520;
wire n_808;
wire n_409;
wire n_797;
wire n_1038;
wire n_1025;
wire n_1082;
wire n_887;
wire n_589;
wire n_716;
wire n_597;
wire n_500;
wire n_562;
wire n_1067;
wire n_300;
wire n_651;
wire n_435;
wire n_809;
wire n_870;
wire n_952;
wire n_334;
wire n_599;
wire n_766;
wire n_811;
wire n_931;
wire n_541;
wire n_807;
wire n_391;
wire n_701;
wire n_434;
wire n_1023;
wire n_645;
wire n_539;
wire n_835;
wire n_538;
wire n_666;
wire n_803;
wire n_868;
wire n_1092;
wire n_639;
wire n_799;
wire n_914;
wire n_687;
wire n_715;
wire n_411;
wire n_414;
wire n_1026;
wire n_319;
wire n_364;
wire n_965;
wire n_927;
wire n_1089;
wire n_536;
wire n_531;
wire n_1004;
wire n_935;
wire n_817;
wire n_872;
wire n_360;
wire n_594;
wire n_764;
wire n_890;
wire n_1056;
wire n_960;
wire n_759;
wire n_1018;
wire n_438;
wire n_806;
wire n_713;
wire n_1011;
wire n_904;
wire n_985;
wire n_1047;
wire n_869;
wire n_324;
wire n_810;
wire n_634;
wire n_416;
wire n_827;
wire n_401;
wire n_348;
wire n_1029;
wire n_626;
wire n_925;
wire n_424;
wire n_1003;
wire n_706;
wire n_746;
wire n_305;
wire n_533;
wire n_950;
wire n_747;
wire n_278;
wire n_784;

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_259),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_18),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_26),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_172),
.Y(n_277)
);

BUFx10_ASAP7_75t_L g278 ( 
.A(n_271),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_157),
.Y(n_279)
);

BUFx6f_ASAP7_75t_L g280 ( 
.A(n_122),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_218),
.Y(n_281)
);

OR2x2_ASAP7_75t_L g282 ( 
.A(n_156),
.B(n_185),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_26),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_202),
.Y(n_284)
);

BUFx10_ASAP7_75t_L g285 ( 
.A(n_173),
.Y(n_285)
);

NOR2xp67_ASAP7_75t_L g286 ( 
.A(n_147),
.B(n_153),
.Y(n_286)
);

BUFx5_ASAP7_75t_L g287 ( 
.A(n_257),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_231),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_221),
.Y(n_289)
);

BUFx6f_ASAP7_75t_L g290 ( 
.A(n_146),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_95),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_272),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_189),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_168),
.Y(n_294)
);

CKINVDCx16_ASAP7_75t_R g295 ( 
.A(n_256),
.Y(n_295)
);

BUFx3_ASAP7_75t_L g296 ( 
.A(n_37),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_206),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_180),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_142),
.Y(n_299)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_229),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_95),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_269),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_37),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_119),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_65),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_116),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_192),
.Y(n_307)
);

CKINVDCx16_ASAP7_75t_R g308 ( 
.A(n_181),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_190),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_225),
.Y(n_310)
);

BUFx3_ASAP7_75t_L g311 ( 
.A(n_239),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_170),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_204),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_110),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_167),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_96),
.Y(n_316)
);

INVx2_ASAP7_75t_SL g317 ( 
.A(n_59),
.Y(n_317)
);

CKINVDCx16_ASAP7_75t_R g318 ( 
.A(n_100),
.Y(n_318)
);

CKINVDCx16_ASAP7_75t_R g319 ( 
.A(n_222),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_237),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_223),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_163),
.Y(n_322)
);

BUFx6f_ASAP7_75t_L g323 ( 
.A(n_132),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_81),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_150),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_273),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_101),
.Y(n_327)
);

BUFx6f_ASAP7_75t_L g328 ( 
.A(n_151),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_91),
.Y(n_329)
);

CKINVDCx16_ASAP7_75t_R g330 ( 
.A(n_11),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_144),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_47),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_213),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_240),
.Y(n_334)
);

BUFx10_ASAP7_75t_L g335 ( 
.A(n_197),
.Y(n_335)
);

INVx1_ASAP7_75t_SL g336 ( 
.A(n_36),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_164),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_155),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_214),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_171),
.Y(n_340)
);

CKINVDCx20_ASAP7_75t_R g341 ( 
.A(n_210),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_3),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_19),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_98),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_28),
.Y(n_345)
);

BUFx3_ASAP7_75t_L g346 ( 
.A(n_143),
.Y(n_346)
);

HB1xp67_ASAP7_75t_L g347 ( 
.A(n_219),
.Y(n_347)
);

CKINVDCx20_ASAP7_75t_R g348 ( 
.A(n_62),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_165),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_182),
.B(n_130),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_254),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_227),
.Y(n_352)
);

INVx1_ASAP7_75t_SL g353 ( 
.A(n_152),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_3),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_183),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_34),
.Y(n_356)
);

CKINVDCx16_ASAP7_75t_R g357 ( 
.A(n_158),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_191),
.Y(n_358)
);

BUFx6f_ASAP7_75t_L g359 ( 
.A(n_255),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g360 ( 
.A(n_187),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_L g361 ( 
.A(n_251),
.B(n_265),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_228),
.Y(n_362)
);

BUFx8_ASAP7_75t_SL g363 ( 
.A(n_193),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_270),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_79),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_133),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_115),
.Y(n_367)
);

BUFx3_ASAP7_75t_L g368 ( 
.A(n_52),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_128),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_195),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_82),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_207),
.Y(n_372)
);

CKINVDCx20_ASAP7_75t_R g373 ( 
.A(n_162),
.Y(n_373)
);

INVxp67_ASAP7_75t_L g374 ( 
.A(n_220),
.Y(n_374)
);

BUFx6f_ASAP7_75t_L g375 ( 
.A(n_230),
.Y(n_375)
);

BUFx5_ASAP7_75t_L g376 ( 
.A(n_17),
.Y(n_376)
);

INVx2_ASAP7_75t_L g377 ( 
.A(n_57),
.Y(n_377)
);

BUFx6f_ASAP7_75t_L g378 ( 
.A(n_129),
.Y(n_378)
);

CKINVDCx20_ASAP7_75t_R g379 ( 
.A(n_241),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_217),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_198),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_8),
.Y(n_382)
);

CKINVDCx20_ASAP7_75t_R g383 ( 
.A(n_114),
.Y(n_383)
);

INVx2_ASAP7_75t_L g384 ( 
.A(n_188),
.Y(n_384)
);

CKINVDCx16_ASAP7_75t_R g385 ( 
.A(n_82),
.Y(n_385)
);

CKINVDCx20_ASAP7_75t_R g386 ( 
.A(n_69),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_57),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_7),
.Y(n_388)
);

INVxp67_ASAP7_75t_SL g389 ( 
.A(n_127),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_235),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_75),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_2),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_266),
.Y(n_393)
);

CKINVDCx20_ASAP7_75t_R g394 ( 
.A(n_56),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_140),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_154),
.Y(n_396)
);

INVx1_ASAP7_75t_SL g397 ( 
.A(n_61),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_24),
.Y(n_398)
);

CKINVDCx20_ASAP7_75t_R g399 ( 
.A(n_244),
.Y(n_399)
);

HB1xp67_ASAP7_75t_L g400 ( 
.A(n_141),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_58),
.Y(n_401)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_264),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_149),
.Y(n_403)
);

CKINVDCx14_ASAP7_75t_R g404 ( 
.A(n_92),
.Y(n_404)
);

XNOR2xp5_ASAP7_75t_L g405 ( 
.A(n_243),
.B(n_64),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_27),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_101),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_0),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_139),
.Y(n_409)
);

BUFx6f_ASAP7_75t_L g410 ( 
.A(n_166),
.Y(n_410)
);

BUFx2_ASAP7_75t_L g411 ( 
.A(n_85),
.Y(n_411)
);

BUFx10_ASAP7_75t_L g412 ( 
.A(n_205),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_61),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_196),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_16),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_263),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_145),
.Y(n_417)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_120),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_245),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_376),
.Y(n_420)
);

AND2x4_ASAP7_75t_L g421 ( 
.A(n_311),
.B(n_0),
.Y(n_421)
);

INVxp67_ASAP7_75t_L g422 ( 
.A(n_411),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_376),
.B(n_404),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_318),
.Y(n_424)
);

BUFx6f_ASAP7_75t_L g425 ( 
.A(n_280),
.Y(n_425)
);

INVx2_ASAP7_75t_L g426 ( 
.A(n_376),
.Y(n_426)
);

OA21x2_ASAP7_75t_L g427 ( 
.A1(n_279),
.A2(n_1),
.B(n_2),
.Y(n_427)
);

AND2x6_ASAP7_75t_L g428 ( 
.A(n_280),
.B(n_290),
.Y(n_428)
);

BUFx6f_ASAP7_75t_L g429 ( 
.A(n_290),
.Y(n_429)
);

OR2x2_ASAP7_75t_L g430 ( 
.A(n_317),
.B(n_4),
.Y(n_430)
);

AND2x2_ASAP7_75t_L g431 ( 
.A(n_296),
.B(n_368),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_376),
.Y(n_432)
);

AND2x2_ASAP7_75t_L g433 ( 
.A(n_330),
.B(n_385),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_376),
.Y(n_434)
);

AND2x4_ASAP7_75t_L g435 ( 
.A(n_346),
.B(n_5),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_275),
.Y(n_436)
);

NOR2x1_ASAP7_75t_L g437 ( 
.A(n_286),
.B(n_5),
.Y(n_437)
);

INVx4_ASAP7_75t_L g438 ( 
.A(n_290),
.Y(n_438)
);

BUFx6f_ASAP7_75t_L g439 ( 
.A(n_323),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_347),
.B(n_6),
.Y(n_440)
);

INVx2_ASAP7_75t_L g441 ( 
.A(n_287),
.Y(n_441)
);

HB1xp67_ASAP7_75t_L g442 ( 
.A(n_301),
.Y(n_442)
);

OA21x2_ASAP7_75t_L g443 ( 
.A1(n_281),
.A2(n_289),
.B(n_288),
.Y(n_443)
);

BUFx6f_ASAP7_75t_L g444 ( 
.A(n_323),
.Y(n_444)
);

BUFx6f_ASAP7_75t_L g445 ( 
.A(n_323),
.Y(n_445)
);

AND2x4_ASAP7_75t_L g446 ( 
.A(n_300),
.B(n_6),
.Y(n_446)
);

AND2x4_ASAP7_75t_L g447 ( 
.A(n_384),
.B(n_7),
.Y(n_447)
);

INVx3_ASAP7_75t_L g448 ( 
.A(n_377),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_276),
.Y(n_449)
);

AND2x6_ASAP7_75t_L g450 ( 
.A(n_328),
.B(n_109),
.Y(n_450)
);

BUFx12f_ASAP7_75t_L g451 ( 
.A(n_278),
.Y(n_451)
);

BUFx6f_ASAP7_75t_L g452 ( 
.A(n_328),
.Y(n_452)
);

BUFx6f_ASAP7_75t_L g453 ( 
.A(n_328),
.Y(n_453)
);

AOI22xp5_ASAP7_75t_L g454 ( 
.A1(n_291),
.A2(n_10),
.B1(n_8),
.B2(n_9),
.Y(n_454)
);

BUFx6f_ASAP7_75t_L g455 ( 
.A(n_359),
.Y(n_455)
);

INVx2_ASAP7_75t_L g456 ( 
.A(n_287),
.Y(n_456)
);

BUFx6f_ASAP7_75t_L g457 ( 
.A(n_359),
.Y(n_457)
);

INVx2_ASAP7_75t_L g458 ( 
.A(n_287),
.Y(n_458)
);

AND2x2_ASAP7_75t_SL g459 ( 
.A(n_295),
.B(n_10),
.Y(n_459)
);

BUFx6f_ASAP7_75t_L g460 ( 
.A(n_359),
.Y(n_460)
);

AND2x2_ASAP7_75t_L g461 ( 
.A(n_308),
.B(n_11),
.Y(n_461)
);

INVx3_ASAP7_75t_L g462 ( 
.A(n_278),
.Y(n_462)
);

OR2x2_ASAP7_75t_L g463 ( 
.A(n_324),
.B(n_12),
.Y(n_463)
);

INVx5_ASAP7_75t_L g464 ( 
.A(n_375),
.Y(n_464)
);

HB1xp67_ASAP7_75t_L g465 ( 
.A(n_342),
.Y(n_465)
);

AOI22xp5_ASAP7_75t_SL g466 ( 
.A1(n_348),
.A2(n_14),
.B1(n_12),
.B2(n_13),
.Y(n_466)
);

AND2x2_ASAP7_75t_L g467 ( 
.A(n_319),
.B(n_13),
.Y(n_467)
);

AND2x4_ASAP7_75t_L g468 ( 
.A(n_402),
.B(n_14),
.Y(n_468)
);

INVxp67_ASAP7_75t_L g469 ( 
.A(n_345),
.Y(n_469)
);

OAI21x1_ASAP7_75t_L g470 ( 
.A1(n_418),
.A2(n_112),
.B(n_111),
.Y(n_470)
);

INVx2_ASAP7_75t_SL g471 ( 
.A(n_285),
.Y(n_471)
);

BUFx3_ASAP7_75t_L g472 ( 
.A(n_285),
.Y(n_472)
);

INVx2_ASAP7_75t_L g473 ( 
.A(n_354),
.Y(n_473)
);

INVx3_ASAP7_75t_L g474 ( 
.A(n_335),
.Y(n_474)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_371),
.Y(n_475)
);

OAI22xp5_ASAP7_75t_SL g476 ( 
.A1(n_386),
.A2(n_18),
.B1(n_15),
.B2(n_17),
.Y(n_476)
);

INVx2_ASAP7_75t_L g477 ( 
.A(n_391),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_398),
.Y(n_478)
);

INVx2_ASAP7_75t_L g479 ( 
.A(n_401),
.Y(n_479)
);

AND2x6_ASAP7_75t_L g480 ( 
.A(n_378),
.B(n_113),
.Y(n_480)
);

BUFx6f_ASAP7_75t_L g481 ( 
.A(n_378),
.Y(n_481)
);

BUFx6f_ASAP7_75t_L g482 ( 
.A(n_378),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_407),
.Y(n_483)
);

INVx2_ASAP7_75t_L g484 ( 
.A(n_408),
.Y(n_484)
);

BUFx12f_ASAP7_75t_L g485 ( 
.A(n_335),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g486 ( 
.A(n_400),
.B(n_19),
.Y(n_486)
);

BUFx6f_ASAP7_75t_L g487 ( 
.A(n_410),
.Y(n_487)
);

HB1xp67_ASAP7_75t_L g488 ( 
.A(n_283),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_423),
.B(n_293),
.Y(n_489)
);

INVx2_ASAP7_75t_L g490 ( 
.A(n_426),
.Y(n_490)
);

AND2x2_ASAP7_75t_L g491 ( 
.A(n_431),
.B(n_357),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_SL g492 ( 
.A(n_459),
.B(n_412),
.Y(n_492)
);

NAND2xp33_ASAP7_75t_L g493 ( 
.A(n_461),
.B(n_410),
.Y(n_493)
);

INVx6_ASAP7_75t_L g494 ( 
.A(n_438),
.Y(n_494)
);

INVx8_ASAP7_75t_L g495 ( 
.A(n_464),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_425),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_420),
.Y(n_497)
);

OR2x2_ASAP7_75t_L g498 ( 
.A(n_488),
.B(n_336),
.Y(n_498)
);

INVx2_ASAP7_75t_L g499 ( 
.A(n_432),
.Y(n_499)
);

INVx2_ASAP7_75t_L g500 ( 
.A(n_434),
.Y(n_500)
);

INVx2_ASAP7_75t_L g501 ( 
.A(n_429),
.Y(n_501)
);

INVxp67_ASAP7_75t_SL g502 ( 
.A(n_423),
.Y(n_502)
);

INVx2_ASAP7_75t_L g503 ( 
.A(n_439),
.Y(n_503)
);

INVx2_ASAP7_75t_L g504 ( 
.A(n_439),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_444),
.Y(n_505)
);

BUFx6f_ASAP7_75t_L g506 ( 
.A(n_444),
.Y(n_506)
);

INVx3_ASAP7_75t_L g507 ( 
.A(n_444),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_445),
.Y(n_508)
);

INVx3_ASAP7_75t_L g509 ( 
.A(n_445),
.Y(n_509)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_445),
.Y(n_510)
);

INVx3_ASAP7_75t_L g511 ( 
.A(n_452),
.Y(n_511)
);

CKINVDCx6p67_ASAP7_75t_R g512 ( 
.A(n_451),
.Y(n_512)
);

OR2x2_ASAP7_75t_L g513 ( 
.A(n_488),
.B(n_397),
.Y(n_513)
);

INVx6_ASAP7_75t_L g514 ( 
.A(n_438),
.Y(n_514)
);

OR2x2_ASAP7_75t_L g515 ( 
.A(n_433),
.B(n_303),
.Y(n_515)
);

INVx2_ASAP7_75t_L g516 ( 
.A(n_453),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_SL g517 ( 
.A(n_459),
.B(n_412),
.Y(n_517)
);

INVx4_ASAP7_75t_L g518 ( 
.A(n_450),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_SL g519 ( 
.A(n_467),
.B(n_305),
.Y(n_519)
);

INVx3_ASAP7_75t_L g520 ( 
.A(n_455),
.Y(n_520)
);

BUFx2_ASAP7_75t_L g521 ( 
.A(n_424),
.Y(n_521)
);

NAND2xp33_ASAP7_75t_L g522 ( 
.A(n_440),
.B(n_316),
.Y(n_522)
);

AO22x2_ASAP7_75t_L g523 ( 
.A1(n_421),
.A2(n_282),
.B1(n_298),
.B2(n_294),
.Y(n_523)
);

AND2x2_ASAP7_75t_L g524 ( 
.A(n_473),
.B(n_353),
.Y(n_524)
);

OAI22xp33_ASAP7_75t_SL g525 ( 
.A1(n_440),
.A2(n_329),
.B1(n_332),
.B2(n_327),
.Y(n_525)
);

INVx2_ASAP7_75t_L g526 ( 
.A(n_457),
.Y(n_526)
);

CKINVDCx6p67_ASAP7_75t_R g527 ( 
.A(n_485),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_SL g528 ( 
.A(n_491),
.B(n_436),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_497),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_502),
.B(n_443),
.Y(n_530)
);

INVx8_ASAP7_75t_L g531 ( 
.A(n_491),
.Y(n_531)
);

AND2x6_ASAP7_75t_L g532 ( 
.A(n_489),
.B(n_421),
.Y(n_532)
);

NOR2x1p5_ASAP7_75t_L g533 ( 
.A(n_512),
.B(n_462),
.Y(n_533)
);

NOR2xp33_ASAP7_75t_L g534 ( 
.A(n_519),
.B(n_436),
.Y(n_534)
);

NOR2xp33_ASAP7_75t_L g535 ( 
.A(n_519),
.B(n_449),
.Y(n_535)
);

BUFx6f_ASAP7_75t_SL g536 ( 
.A(n_527),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_SL g537 ( 
.A(n_492),
.B(n_449),
.Y(n_537)
);

INVx2_ASAP7_75t_L g538 ( 
.A(n_501),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_493),
.B(n_443),
.Y(n_539)
);

NAND3xp33_ASAP7_75t_L g540 ( 
.A(n_492),
.B(n_486),
.C(n_422),
.Y(n_540)
);

HB1xp67_ASAP7_75t_L g541 ( 
.A(n_498),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_497),
.Y(n_542)
);

NAND2xp33_ASAP7_75t_L g543 ( 
.A(n_517),
.B(n_450),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_499),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_SL g545 ( 
.A(n_517),
.B(n_525),
.Y(n_545)
);

INVx2_ASAP7_75t_L g546 ( 
.A(n_503),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_500),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_490),
.Y(n_548)
);

AOI22xp33_ASAP7_75t_L g549 ( 
.A1(n_523),
.A2(n_447),
.B1(n_468),
.B2(n_446),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_L g550 ( 
.A(n_490),
.B(n_441),
.Y(n_550)
);

NOR2xp33_ASAP7_75t_L g551 ( 
.A(n_515),
.B(n_424),
.Y(n_551)
);

NOR2xp33_ASAP7_75t_L g552 ( 
.A(n_494),
.B(n_462),
.Y(n_552)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_503),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_SL g554 ( 
.A(n_524),
.B(n_474),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_504),
.Y(n_555)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_504),
.Y(n_556)
);

INVx2_ASAP7_75t_SL g557 ( 
.A(n_498),
.Y(n_557)
);

NAND2xp33_ASAP7_75t_L g558 ( 
.A(n_523),
.B(n_450),
.Y(n_558)
);

AND2x2_ASAP7_75t_L g559 ( 
.A(n_513),
.B(n_471),
.Y(n_559)
);

NOR2xp33_ASAP7_75t_L g560 ( 
.A(n_494),
.B(n_472),
.Y(n_560)
);

A2O1A1Ixp33_ASAP7_75t_L g561 ( 
.A1(n_522),
.A2(n_486),
.B(n_468),
.C(n_447),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_L g562 ( 
.A(n_510),
.B(n_456),
.Y(n_562)
);

INVx5_ASAP7_75t_L g563 ( 
.A(n_495),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_SL g564 ( 
.A(n_513),
.B(n_435),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_L g565 ( 
.A(n_516),
.B(n_457),
.Y(n_565)
);

INVxp67_ASAP7_75t_L g566 ( 
.A(n_521),
.Y(n_566)
);

NOR2xp33_ASAP7_75t_L g567 ( 
.A(n_494),
.B(n_422),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_L g568 ( 
.A(n_526),
.B(n_458),
.Y(n_568)
);

BUFx6f_ASAP7_75t_L g569 ( 
.A(n_506),
.Y(n_569)
);

OR2x6_ASAP7_75t_L g570 ( 
.A(n_523),
.B(n_476),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_507),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_L g572 ( 
.A(n_509),
.B(n_457),
.Y(n_572)
);

NOR2xp33_ASAP7_75t_L g573 ( 
.A(n_514),
.B(n_430),
.Y(n_573)
);

NOR2xp33_ASAP7_75t_L g574 ( 
.A(n_514),
.B(n_374),
.Y(n_574)
);

INVxp33_ASAP7_75t_L g575 ( 
.A(n_496),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_L g576 ( 
.A(n_509),
.B(n_460),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_SL g577 ( 
.A(n_518),
.B(n_437),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_L g578 ( 
.A(n_511),
.B(n_460),
.Y(n_578)
);

INVxp67_ASAP7_75t_L g579 ( 
.A(n_522),
.Y(n_579)
);

CKINVDCx5p33_ASAP7_75t_R g580 ( 
.A(n_512),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_520),
.Y(n_581)
);

OAI22xp5_ASAP7_75t_L g582 ( 
.A1(n_527),
.A2(n_454),
.B1(n_394),
.B2(n_463),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_562),
.Y(n_583)
);

AOI22xp5_ASAP7_75t_L g584 ( 
.A1(n_579),
.A2(n_535),
.B1(n_534),
.B2(n_545),
.Y(n_584)
);

O2A1O1Ixp33_ASAP7_75t_L g585 ( 
.A1(n_530),
.A2(n_469),
.B(n_442),
.C(n_465),
.Y(n_585)
);

INVx2_ASAP7_75t_L g586 ( 
.A(n_548),
.Y(n_586)
);

AO32x2_ASAP7_75t_L g587 ( 
.A1(n_582),
.A2(n_476),
.A3(n_427),
.B1(n_466),
.B2(n_470),
.Y(n_587)
);

AOI21xp5_ASAP7_75t_L g588 ( 
.A1(n_577),
.A2(n_350),
.B(n_389),
.Y(n_588)
);

OAI21xp5_ASAP7_75t_L g589 ( 
.A1(n_561),
.A2(n_427),
.B(n_302),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_562),
.Y(n_590)
);

O2A1O1Ixp33_ASAP7_75t_L g591 ( 
.A1(n_543),
.A2(n_564),
.B(n_558),
.C(n_554),
.Y(n_591)
);

INVx2_ASAP7_75t_L g592 ( 
.A(n_529),
.Y(n_592)
);

BUFx6f_ASAP7_75t_L g593 ( 
.A(n_569),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_SL g594 ( 
.A(n_559),
.B(n_292),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_568),
.Y(n_595)
);

AOI21xp33_ASAP7_75t_L g596 ( 
.A1(n_540),
.A2(n_405),
.B(n_466),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_L g597 ( 
.A(n_574),
.B(n_520),
.Y(n_597)
);

AO21x1_ASAP7_75t_L g598 ( 
.A1(n_537),
.A2(n_361),
.B(n_313),
.Y(n_598)
);

AO22x1_ASAP7_75t_L g599 ( 
.A1(n_551),
.A2(n_344),
.B1(n_356),
.B2(n_343),
.Y(n_599)
);

OAI22xp5_ASAP7_75t_L g600 ( 
.A1(n_549),
.A2(n_322),
.B1(n_331),
.B2(n_299),
.Y(n_600)
);

CKINVDCx5p33_ASAP7_75t_R g601 ( 
.A(n_536),
.Y(n_601)
);

INVx4_ASAP7_75t_L g602 ( 
.A(n_531),
.Y(n_602)
);

AO32x1_ASAP7_75t_L g603 ( 
.A1(n_555),
.A2(n_314),
.A3(n_326),
.B1(n_320),
.B2(n_312),
.Y(n_603)
);

AOI21x1_ASAP7_75t_L g604 ( 
.A1(n_568),
.A2(n_508),
.B(n_505),
.Y(n_604)
);

NOR2xp67_ASAP7_75t_L g605 ( 
.A(n_566),
.B(n_580),
.Y(n_605)
);

NOR2xp33_ASAP7_75t_L g606 ( 
.A(n_567),
.B(n_341),
.Y(n_606)
);

INVx3_ASAP7_75t_L g607 ( 
.A(n_538),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_SL g608 ( 
.A(n_552),
.B(n_360),
.Y(n_608)
);

CKINVDCx6p67_ASAP7_75t_R g609 ( 
.A(n_541),
.Y(n_609)
);

NOR2x1_ASAP7_75t_L g610 ( 
.A(n_533),
.B(n_373),
.Y(n_610)
);

INVx5_ASAP7_75t_L g611 ( 
.A(n_532),
.Y(n_611)
);

BUFx2_ASAP7_75t_L g612 ( 
.A(n_531),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_565),
.Y(n_613)
);

BUFx6f_ASAP7_75t_L g614 ( 
.A(n_569),
.Y(n_614)
);

AOI21xp5_ASAP7_75t_L g615 ( 
.A1(n_550),
.A2(n_544),
.B(n_542),
.Y(n_615)
);

AOI21xp5_ASAP7_75t_L g616 ( 
.A1(n_547),
.A2(n_340),
.B(n_337),
.Y(n_616)
);

OAI21xp5_ASAP7_75t_L g617 ( 
.A1(n_528),
.A2(n_351),
.B(n_349),
.Y(n_617)
);

NOR2xp33_ASAP7_75t_L g618 ( 
.A(n_560),
.B(n_379),
.Y(n_618)
);

AOI21xp5_ASAP7_75t_L g619 ( 
.A1(n_563),
.A2(n_358),
.B(n_352),
.Y(n_619)
);

AND2x2_ASAP7_75t_L g620 ( 
.A(n_575),
.B(n_465),
.Y(n_620)
);

AOI21xp5_ASAP7_75t_L g621 ( 
.A1(n_572),
.A2(n_578),
.B(n_576),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_L g622 ( 
.A(n_546),
.B(n_409),
.Y(n_622)
);

INVx2_ASAP7_75t_L g623 ( 
.A(n_553),
.Y(n_623)
);

NOR2xp33_ASAP7_75t_L g624 ( 
.A(n_571),
.B(n_383),
.Y(n_624)
);

OAI21xp5_ASAP7_75t_L g625 ( 
.A1(n_581),
.A2(n_416),
.B(n_414),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_L g626 ( 
.A(n_556),
.B(n_417),
.Y(n_626)
);

OR2x2_ASAP7_75t_L g627 ( 
.A(n_570),
.B(n_478),
.Y(n_627)
);

OAI21x1_ASAP7_75t_L g628 ( 
.A1(n_539),
.A2(n_477),
.B(n_475),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_573),
.B(n_480),
.Y(n_629)
);

AO21x1_ASAP7_75t_L g630 ( 
.A1(n_558),
.A2(n_483),
.B(n_479),
.Y(n_630)
);

INVx2_ASAP7_75t_L g631 ( 
.A(n_548),
.Y(n_631)
);

A2O1A1Ixp33_ASAP7_75t_L g632 ( 
.A1(n_561),
.A2(n_484),
.B(n_277),
.C(n_284),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_SL g633 ( 
.A(n_534),
.B(n_399),
.Y(n_633)
);

BUFx2_ASAP7_75t_L g634 ( 
.A(n_557),
.Y(n_634)
);

AOI21x1_ASAP7_75t_L g635 ( 
.A1(n_530),
.A2(n_428),
.B(n_506),
.Y(n_635)
);

INVx1_ASAP7_75t_SL g636 ( 
.A(n_559),
.Y(n_636)
);

NOR2xp33_ASAP7_75t_R g637 ( 
.A(n_580),
.B(n_274),
.Y(n_637)
);

INVx1_ASAP7_75t_SL g638 ( 
.A(n_559),
.Y(n_638)
);

NOR2xp33_ASAP7_75t_L g639 ( 
.A(n_534),
.B(n_365),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_562),
.Y(n_640)
);

INVxp67_ASAP7_75t_L g641 ( 
.A(n_559),
.Y(n_641)
);

BUFx12f_ASAP7_75t_L g642 ( 
.A(n_580),
.Y(n_642)
);

AOI21xp33_ASAP7_75t_L g643 ( 
.A1(n_534),
.A2(n_387),
.B(n_382),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_L g644 ( 
.A(n_573),
.B(n_297),
.Y(n_644)
);

AOI21x1_ASAP7_75t_L g645 ( 
.A1(n_530),
.A2(n_428),
.B(n_481),
.Y(n_645)
);

A2O1A1Ixp33_ASAP7_75t_L g646 ( 
.A1(n_561),
.A2(n_306),
.B(n_307),
.C(n_304),
.Y(n_646)
);

OR2x6_ASAP7_75t_L g647 ( 
.A(n_557),
.B(n_448),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_573),
.B(n_309),
.Y(n_648)
);

AOI22xp5_ASAP7_75t_L g649 ( 
.A1(n_579),
.A2(n_315),
.B1(n_321),
.B2(n_310),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_SL g650 ( 
.A(n_534),
.B(n_325),
.Y(n_650)
);

O2A1O1Ixp33_ASAP7_75t_SL g651 ( 
.A1(n_561),
.A2(n_428),
.B(n_363),
.C(n_392),
.Y(n_651)
);

A2O1A1Ixp33_ASAP7_75t_L g652 ( 
.A1(n_561),
.A2(n_334),
.B(n_338),
.C(n_333),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_L g653 ( 
.A(n_573),
.B(n_339),
.Y(n_653)
);

AOI21xp5_ASAP7_75t_L g654 ( 
.A1(n_530),
.A2(n_487),
.B(n_482),
.Y(n_654)
);

AOI21xp5_ASAP7_75t_L g655 ( 
.A1(n_530),
.A2(n_487),
.B(n_355),
.Y(n_655)
);

AOI21x1_ASAP7_75t_L g656 ( 
.A1(n_635),
.A2(n_645),
.B(n_629),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_586),
.Y(n_657)
);

AND2x2_ASAP7_75t_L g658 ( 
.A(n_636),
.B(n_388),
.Y(n_658)
);

AOI221x1_ASAP7_75t_L g659 ( 
.A1(n_632),
.A2(n_428),
.B1(n_364),
.B2(n_366),
.C(n_362),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_631),
.Y(n_660)
);

BUFx2_ASAP7_75t_L g661 ( 
.A(n_634),
.Y(n_661)
);

OAI21x1_ASAP7_75t_L g662 ( 
.A1(n_621),
.A2(n_615),
.B(n_604),
.Y(n_662)
);

OAI22xp5_ASAP7_75t_L g663 ( 
.A1(n_584),
.A2(n_369),
.B1(n_370),
.B2(n_367),
.Y(n_663)
);

BUFx6f_ASAP7_75t_L g664 ( 
.A(n_593),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_SL g665 ( 
.A(n_638),
.B(n_372),
.Y(n_665)
);

NOR2x1_ASAP7_75t_SL g666 ( 
.A(n_611),
.B(n_117),
.Y(n_666)
);

AO22x2_ASAP7_75t_L g667 ( 
.A1(n_600),
.A2(n_22),
.B1(n_20),
.B2(n_21),
.Y(n_667)
);

NAND2x1p5_ASAP7_75t_L g668 ( 
.A(n_602),
.B(n_118),
.Y(n_668)
);

INVx4_ASAP7_75t_L g669 ( 
.A(n_602),
.Y(n_669)
);

CKINVDCx6p67_ASAP7_75t_R g670 ( 
.A(n_642),
.Y(n_670)
);

INVxp67_ASAP7_75t_L g671 ( 
.A(n_620),
.Y(n_671)
);

AO21x1_ASAP7_75t_L g672 ( 
.A1(n_589),
.A2(n_20),
.B(n_21),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_606),
.B(n_380),
.Y(n_673)
);

AOI21xp33_ASAP7_75t_L g674 ( 
.A1(n_633),
.A2(n_618),
.B(n_641),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_583),
.B(n_381),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_590),
.B(n_390),
.Y(n_676)
);

INVx2_ASAP7_75t_SL g677 ( 
.A(n_647),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_L g678 ( 
.A(n_595),
.B(n_393),
.Y(n_678)
);

NOR2xp33_ASAP7_75t_L g679 ( 
.A(n_594),
.B(n_406),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_640),
.B(n_395),
.Y(n_680)
);

OR2x6_ASAP7_75t_L g681 ( 
.A(n_612),
.B(n_22),
.Y(n_681)
);

AOI21xp5_ASAP7_75t_SL g682 ( 
.A1(n_591),
.A2(n_614),
.B(n_593),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_644),
.B(n_396),
.Y(n_683)
);

AND2x4_ASAP7_75t_L g684 ( 
.A(n_627),
.B(n_592),
.Y(n_684)
);

NOR2x1_ASAP7_75t_SL g685 ( 
.A(n_611),
.B(n_121),
.Y(n_685)
);

BUFx2_ASAP7_75t_L g686 ( 
.A(n_609),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_SL g687 ( 
.A(n_648),
.B(n_403),
.Y(n_687)
);

AOI221x1_ASAP7_75t_L g688 ( 
.A1(n_646),
.A2(n_419),
.B1(n_125),
.B2(n_126),
.C(n_124),
.Y(n_688)
);

A2O1A1Ixp33_ASAP7_75t_L g689 ( 
.A1(n_643),
.A2(n_415),
.B(n_413),
.C(n_25),
.Y(n_689)
);

O2A1O1Ixp33_ASAP7_75t_L g690 ( 
.A1(n_585),
.A2(n_25),
.B(n_23),
.C(n_24),
.Y(n_690)
);

NOR2x1_ASAP7_75t_SL g691 ( 
.A(n_611),
.B(n_123),
.Y(n_691)
);

CKINVDCx5p33_ASAP7_75t_R g692 ( 
.A(n_637),
.Y(n_692)
);

INVx2_ASAP7_75t_L g693 ( 
.A(n_623),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_L g694 ( 
.A(n_653),
.B(n_23),
.Y(n_694)
);

A2O1A1Ixp33_ASAP7_75t_L g695 ( 
.A1(n_617),
.A2(n_30),
.B(n_28),
.C(n_29),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_L g696 ( 
.A(n_613),
.B(n_29),
.Y(n_696)
);

AND2x4_ASAP7_75t_L g697 ( 
.A(n_610),
.B(n_131),
.Y(n_697)
);

AO31x2_ASAP7_75t_L g698 ( 
.A1(n_630),
.A2(n_33),
.A3(n_31),
.B(n_32),
.Y(n_698)
);

AOI211x1_ASAP7_75t_L g699 ( 
.A1(n_598),
.A2(n_35),
.B(n_32),
.C(n_33),
.Y(n_699)
);

AO21x1_ASAP7_75t_L g700 ( 
.A1(n_588),
.A2(n_35),
.B(n_38),
.Y(n_700)
);

AOI21xp33_ASAP7_75t_L g701 ( 
.A1(n_650),
.A2(n_38),
.B(n_39),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_L g702 ( 
.A(n_624),
.B(n_40),
.Y(n_702)
);

OAI21xp5_ASAP7_75t_L g703 ( 
.A1(n_652),
.A2(n_135),
.B(n_134),
.Y(n_703)
);

AND2x2_ASAP7_75t_L g704 ( 
.A(n_608),
.B(n_40),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_L g705 ( 
.A(n_597),
.B(n_41),
.Y(n_705)
);

A2O1A1Ixp33_ASAP7_75t_L g706 ( 
.A1(n_596),
.A2(n_43),
.B(n_41),
.C(n_42),
.Y(n_706)
);

AND2x4_ASAP7_75t_L g707 ( 
.A(n_605),
.B(n_136),
.Y(n_707)
);

NAND3xp33_ASAP7_75t_L g708 ( 
.A(n_599),
.B(n_43),
.C(n_44),
.Y(n_708)
);

OAI21xp5_ASAP7_75t_L g709 ( 
.A1(n_655),
.A2(n_138),
.B(n_137),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_L g710 ( 
.A(n_654),
.B(n_45),
.Y(n_710)
);

AND2x4_ASAP7_75t_L g711 ( 
.A(n_607),
.B(n_148),
.Y(n_711)
);

AO31x2_ASAP7_75t_L g712 ( 
.A1(n_622),
.A2(n_48),
.A3(n_46),
.B(n_47),
.Y(n_712)
);

AOI211x1_ASAP7_75t_L g713 ( 
.A1(n_616),
.A2(n_51),
.B(n_49),
.C(n_50),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_L g714 ( 
.A(n_649),
.B(n_51),
.Y(n_714)
);

INVx2_ASAP7_75t_L g715 ( 
.A(n_626),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_625),
.B(n_52),
.Y(n_716)
);

NOR3xp33_ASAP7_75t_L g717 ( 
.A(n_601),
.B(n_53),
.C(n_54),
.Y(n_717)
);

OAI21xp5_ASAP7_75t_SL g718 ( 
.A1(n_587),
.A2(n_54),
.B(n_55),
.Y(n_718)
);

OAI22xp5_ASAP7_75t_L g719 ( 
.A1(n_619),
.A2(n_160),
.B1(n_161),
.B2(n_159),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_651),
.B(n_55),
.Y(n_720)
);

BUFx6f_ASAP7_75t_SL g721 ( 
.A(n_587),
.Y(n_721)
);

A2O1A1Ixp33_ASAP7_75t_L g722 ( 
.A1(n_603),
.A2(n_59),
.B(n_56),
.C(n_58),
.Y(n_722)
);

BUFx6f_ASAP7_75t_L g723 ( 
.A(n_603),
.Y(n_723)
);

OAI22xp5_ASAP7_75t_L g724 ( 
.A1(n_584),
.A2(n_174),
.B1(n_175),
.B2(n_169),
.Y(n_724)
);

AND2x4_ASAP7_75t_L g725 ( 
.A(n_602),
.B(n_176),
.Y(n_725)
);

OR2x2_ASAP7_75t_L g726 ( 
.A(n_636),
.B(n_60),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_L g727 ( 
.A(n_639),
.B(n_62),
.Y(n_727)
);

NAND3xp33_ASAP7_75t_L g728 ( 
.A(n_639),
.B(n_63),
.C(n_64),
.Y(n_728)
);

OAI22xp5_ASAP7_75t_L g729 ( 
.A1(n_584),
.A2(n_178),
.B1(n_179),
.B2(n_177),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_639),
.B(n_63),
.Y(n_730)
);

AOI21xp33_ASAP7_75t_L g731 ( 
.A1(n_639),
.A2(n_65),
.B(n_66),
.Y(n_731)
);

INVx3_ASAP7_75t_L g732 ( 
.A(n_609),
.Y(n_732)
);

OA22x2_ASAP7_75t_L g733 ( 
.A1(n_584),
.A2(n_66),
.B1(n_67),
.B2(n_68),
.Y(n_733)
);

NOR2xp33_ASAP7_75t_L g734 ( 
.A(n_606),
.B(n_67),
.Y(n_734)
);

OAI22xp5_ASAP7_75t_L g735 ( 
.A1(n_584),
.A2(n_208),
.B1(n_268),
.B2(n_267),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_L g736 ( 
.A(n_639),
.B(n_68),
.Y(n_736)
);

INVx3_ASAP7_75t_L g737 ( 
.A(n_609),
.Y(n_737)
);

NAND2x1p5_ASAP7_75t_L g738 ( 
.A(n_602),
.B(n_184),
.Y(n_738)
);

OAI21xp33_ASAP7_75t_L g739 ( 
.A1(n_639),
.A2(n_69),
.B(n_70),
.Y(n_739)
);

BUFx12f_ASAP7_75t_L g740 ( 
.A(n_642),
.Y(n_740)
);

NOR2x1_ASAP7_75t_SL g741 ( 
.A(n_611),
.B(n_186),
.Y(n_741)
);

AOI21xp33_ASAP7_75t_L g742 ( 
.A1(n_639),
.A2(n_70),
.B(n_71),
.Y(n_742)
);

AO31x2_ASAP7_75t_L g743 ( 
.A1(n_630),
.A2(n_72),
.A3(n_73),
.B(n_74),
.Y(n_743)
);

AO31x2_ASAP7_75t_L g744 ( 
.A1(n_630),
.A2(n_74),
.A3(n_75),
.B(n_76),
.Y(n_744)
);

AOI221x1_ASAP7_75t_L g745 ( 
.A1(n_632),
.A2(n_216),
.B1(n_262),
.B2(n_261),
.C(n_260),
.Y(n_745)
);

INVx5_ASAP7_75t_L g746 ( 
.A(n_593),
.Y(n_746)
);

INVx5_ASAP7_75t_L g747 ( 
.A(n_593),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_639),
.B(n_77),
.Y(n_748)
);

AO31x2_ASAP7_75t_L g749 ( 
.A1(n_630),
.A2(n_77),
.A3(n_78),
.B(n_79),
.Y(n_749)
);

NAND3xp33_ASAP7_75t_L g750 ( 
.A(n_639),
.B(n_78),
.C(n_80),
.Y(n_750)
);

BUFx3_ASAP7_75t_L g751 ( 
.A(n_661),
.Y(n_751)
);

NAND3xp33_ASAP7_75t_L g752 ( 
.A(n_734),
.B(n_80),
.C(n_81),
.Y(n_752)
);

BUFx12f_ASAP7_75t_L g753 ( 
.A(n_740),
.Y(n_753)
);

OAI21xp5_ASAP7_75t_L g754 ( 
.A1(n_727),
.A2(n_212),
.B(n_253),
.Y(n_754)
);

OAI21xp5_ASAP7_75t_L g755 ( 
.A1(n_730),
.A2(n_211),
.B(n_252),
.Y(n_755)
);

AOI22xp33_ASAP7_75t_L g756 ( 
.A1(n_721),
.A2(n_83),
.B1(n_84),
.B2(n_85),
.Y(n_756)
);

OA21x2_ASAP7_75t_L g757 ( 
.A1(n_688),
.A2(n_215),
.B(n_250),
.Y(n_757)
);

NAND3xp33_ASAP7_75t_L g758 ( 
.A(n_679),
.B(n_83),
.C(n_84),
.Y(n_758)
);

AND2x4_ASAP7_75t_L g759 ( 
.A(n_684),
.B(n_194),
.Y(n_759)
);

AO21x2_ASAP7_75t_L g760 ( 
.A1(n_703),
.A2(n_224),
.B(n_249),
.Y(n_760)
);

INVx1_ASAP7_75t_SL g761 ( 
.A(n_726),
.Y(n_761)
);

OAI21xp5_ASAP7_75t_L g762 ( 
.A1(n_736),
.A2(n_209),
.B(n_248),
.Y(n_762)
);

AOI222xp33_ASAP7_75t_L g763 ( 
.A1(n_671),
.A2(n_718),
.B1(n_739),
.B2(n_667),
.C1(n_702),
.C2(n_704),
.Y(n_763)
);

AO21x2_ASAP7_75t_L g764 ( 
.A1(n_682),
.A2(n_203),
.B(n_247),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_657),
.Y(n_765)
);

INVx1_ASAP7_75t_SL g766 ( 
.A(n_686),
.Y(n_766)
);

OR2x2_ASAP7_75t_L g767 ( 
.A(n_658),
.B(n_86),
.Y(n_767)
);

AO21x2_ASAP7_75t_L g768 ( 
.A1(n_709),
.A2(n_226),
.B(n_246),
.Y(n_768)
);

AOI22xp33_ASAP7_75t_L g769 ( 
.A1(n_748),
.A2(n_86),
.B1(n_87),
.B2(n_88),
.Y(n_769)
);

CKINVDCx5p33_ASAP7_75t_R g770 ( 
.A(n_692),
.Y(n_770)
);

OAI22xp33_ASAP7_75t_L g771 ( 
.A1(n_714),
.A2(n_87),
.B1(n_88),
.B2(n_89),
.Y(n_771)
);

OAI211xp5_ASAP7_75t_L g772 ( 
.A1(n_731),
.A2(n_89),
.B(n_90),
.C(n_91),
.Y(n_772)
);

AND3x2_ASAP7_75t_L g773 ( 
.A(n_717),
.B(n_92),
.C(n_93),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_L g774 ( 
.A(n_673),
.B(n_93),
.Y(n_774)
);

CKINVDCx20_ASAP7_75t_R g775 ( 
.A(n_670),
.Y(n_775)
);

BUFx2_ASAP7_75t_L g776 ( 
.A(n_681),
.Y(n_776)
);

HB1xp67_ASAP7_75t_L g777 ( 
.A(n_677),
.Y(n_777)
);

BUFx6f_ASAP7_75t_L g778 ( 
.A(n_664),
.Y(n_778)
);

BUFx10_ASAP7_75t_L g779 ( 
.A(n_707),
.Y(n_779)
);

BUFx3_ASAP7_75t_L g780 ( 
.A(n_732),
.Y(n_780)
);

OA21x2_ASAP7_75t_L g781 ( 
.A1(n_745),
.A2(n_201),
.B(n_242),
.Y(n_781)
);

BUFx6f_ASAP7_75t_L g782 ( 
.A(n_664),
.Y(n_782)
);

INVx2_ASAP7_75t_L g783 ( 
.A(n_660),
.Y(n_783)
);

AO31x2_ASAP7_75t_L g784 ( 
.A1(n_672),
.A2(n_94),
.A3(n_97),
.B(n_98),
.Y(n_784)
);

AO31x2_ASAP7_75t_L g785 ( 
.A1(n_722),
.A2(n_99),
.A3(n_100),
.B(n_102),
.Y(n_785)
);

CKINVDCx5p33_ASAP7_75t_R g786 ( 
.A(n_737),
.Y(n_786)
);

BUFx12f_ASAP7_75t_L g787 ( 
.A(n_681),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_715),
.Y(n_788)
);

OR2x6_ASAP7_75t_L g789 ( 
.A(n_725),
.B(n_99),
.Y(n_789)
);

NAND2x1p5_ASAP7_75t_L g790 ( 
.A(n_669),
.B(n_232),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_664),
.Y(n_791)
);

INVx5_ASAP7_75t_L g792 ( 
.A(n_746),
.Y(n_792)
);

NAND2x1p5_ASAP7_75t_L g793 ( 
.A(n_746),
.B(n_200),
.Y(n_793)
);

BUFx4_ASAP7_75t_SL g794 ( 
.A(n_708),
.Y(n_794)
);

INVx1_ASAP7_75t_SL g795 ( 
.A(n_696),
.Y(n_795)
);

AND2x4_ASAP7_75t_L g796 ( 
.A(n_707),
.B(n_199),
.Y(n_796)
);

AND2x2_ASAP7_75t_L g797 ( 
.A(n_675),
.B(n_103),
.Y(n_797)
);

AOI22xp5_ASAP7_75t_L g798 ( 
.A1(n_694),
.A2(n_233),
.B1(n_238),
.B2(n_236),
.Y(n_798)
);

BUFx2_ASAP7_75t_L g799 ( 
.A(n_711),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_L g800 ( 
.A(n_676),
.B(n_678),
.Y(n_800)
);

AND2x2_ASAP7_75t_L g801 ( 
.A(n_680),
.B(n_103),
.Y(n_801)
);

INVx2_ASAP7_75t_L g802 ( 
.A(n_747),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_L g803 ( 
.A(n_683),
.B(n_104),
.Y(n_803)
);

INVx2_ASAP7_75t_L g804 ( 
.A(n_747),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_L g805 ( 
.A(n_705),
.B(n_105),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_710),
.Y(n_806)
);

INVx2_ASAP7_75t_SL g807 ( 
.A(n_665),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_733),
.Y(n_808)
);

CKINVDCx20_ASAP7_75t_R g809 ( 
.A(n_687),
.Y(n_809)
);

CKINVDCx6p67_ASAP7_75t_R g810 ( 
.A(n_697),
.Y(n_810)
);

OR2x2_ASAP7_75t_L g811 ( 
.A(n_663),
.B(n_105),
.Y(n_811)
);

BUFx4f_ASAP7_75t_L g812 ( 
.A(n_668),
.Y(n_812)
);

AND2x2_ASAP7_75t_L g813 ( 
.A(n_689),
.B(n_106),
.Y(n_813)
);

CKINVDCx11_ASAP7_75t_R g814 ( 
.A(n_724),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_L g815 ( 
.A(n_716),
.B(n_107),
.Y(n_815)
);

NOR2xp67_ASAP7_75t_L g816 ( 
.A(n_728),
.B(n_234),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_700),
.Y(n_817)
);

AOI31xp67_ASAP7_75t_L g818 ( 
.A1(n_720),
.A2(n_258),
.A3(n_107),
.B(n_108),
.Y(n_818)
);

OR2x2_ASAP7_75t_L g819 ( 
.A(n_706),
.B(n_750),
.Y(n_819)
);

AOI222xp33_ASAP7_75t_L g820 ( 
.A1(n_667),
.A2(n_695),
.B1(n_735),
.B2(n_729),
.C1(n_719),
.C2(n_742),
.Y(n_820)
);

AOI22xp33_ASAP7_75t_SL g821 ( 
.A1(n_666),
.A2(n_741),
.B1(n_685),
.B2(n_691),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_698),
.Y(n_822)
);

INVx4_ASAP7_75t_L g823 ( 
.A(n_738),
.Y(n_823)
);

INVx1_ASAP7_75t_SL g824 ( 
.A(n_701),
.Y(n_824)
);

INVxp67_ASAP7_75t_SL g825 ( 
.A(n_690),
.Y(n_825)
);

AO31x2_ASAP7_75t_L g826 ( 
.A1(n_723),
.A2(n_713),
.A3(n_698),
.B(n_743),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_743),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_744),
.Y(n_828)
);

BUFx6f_ASAP7_75t_L g829 ( 
.A(n_744),
.Y(n_829)
);

INVx2_ASAP7_75t_L g830 ( 
.A(n_749),
.Y(n_830)
);

INVx1_ASAP7_75t_SL g831 ( 
.A(n_712),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_749),
.Y(n_832)
);

OAI21x1_ASAP7_75t_SL g833 ( 
.A1(n_672),
.A2(n_630),
.B(n_666),
.Y(n_833)
);

AO31x2_ASAP7_75t_L g834 ( 
.A1(n_672),
.A2(n_659),
.A3(n_688),
.B(n_722),
.Y(n_834)
);

OR2x6_ASAP7_75t_L g835 ( 
.A(n_661),
.B(n_740),
.Y(n_835)
);

AO21x1_ASAP7_75t_L g836 ( 
.A1(n_727),
.A2(n_736),
.B(n_730),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_693),
.Y(n_837)
);

INVx1_ASAP7_75t_SL g838 ( 
.A(n_661),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_L g839 ( 
.A(n_673),
.B(n_502),
.Y(n_839)
);

OR2x2_ASAP7_75t_L g840 ( 
.A(n_671),
.B(n_557),
.Y(n_840)
);

CKINVDCx5p33_ASAP7_75t_R g841 ( 
.A(n_692),
.Y(n_841)
);

NOR2xp33_ASAP7_75t_L g842 ( 
.A(n_674),
.B(n_606),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_657),
.Y(n_843)
);

BUFx12f_ASAP7_75t_L g844 ( 
.A(n_740),
.Y(n_844)
);

OAI21x1_ASAP7_75t_L g845 ( 
.A1(n_656),
.A2(n_628),
.B(n_662),
.Y(n_845)
);

AO22x2_ASAP7_75t_L g846 ( 
.A1(n_718),
.A2(n_699),
.B1(n_582),
.B2(n_713),
.Y(n_846)
);

OR2x2_ASAP7_75t_L g847 ( 
.A(n_838),
.B(n_761),
.Y(n_847)
);

AND2x2_ASAP7_75t_L g848 ( 
.A(n_795),
.B(n_842),
.Y(n_848)
);

INVx2_ASAP7_75t_SL g849 ( 
.A(n_751),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_788),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_788),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_L g852 ( 
.A(n_800),
.B(n_839),
.Y(n_852)
);

INVx2_ASAP7_75t_L g853 ( 
.A(n_765),
.Y(n_853)
);

INVx2_ASAP7_75t_L g854 ( 
.A(n_843),
.Y(n_854)
);

INVx1_ASAP7_75t_SL g855 ( 
.A(n_840),
.Y(n_855)
);

INVx2_ASAP7_75t_L g856 ( 
.A(n_783),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_837),
.Y(n_857)
);

AND2x4_ASAP7_75t_L g858 ( 
.A(n_799),
.B(n_759),
.Y(n_858)
);

BUFx2_ASAP7_75t_L g859 ( 
.A(n_776),
.Y(n_859)
);

BUFx2_ASAP7_75t_L g860 ( 
.A(n_777),
.Y(n_860)
);

CKINVDCx5p33_ASAP7_75t_R g861 ( 
.A(n_770),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_808),
.Y(n_862)
);

AO21x2_ASAP7_75t_L g863 ( 
.A1(n_845),
.A2(n_817),
.B(n_836),
.Y(n_863)
);

AND2x2_ASAP7_75t_L g864 ( 
.A(n_824),
.B(n_797),
.Y(n_864)
);

INVx2_ASAP7_75t_SL g865 ( 
.A(n_780),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_791),
.Y(n_866)
);

CKINVDCx20_ASAP7_75t_R g867 ( 
.A(n_775),
.Y(n_867)
);

INVx2_ASAP7_75t_L g868 ( 
.A(n_806),
.Y(n_868)
);

INVx1_ASAP7_75t_SL g869 ( 
.A(n_766),
.Y(n_869)
);

HB1xp67_ASAP7_75t_L g870 ( 
.A(n_792),
.Y(n_870)
);

CKINVDCx20_ASAP7_75t_R g871 ( 
.A(n_841),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_763),
.B(n_817),
.Y(n_872)
);

INVxp67_ASAP7_75t_L g873 ( 
.A(n_767),
.Y(n_873)
);

CKINVDCx5p33_ASAP7_75t_R g874 ( 
.A(n_753),
.Y(n_874)
);

AND2x2_ASAP7_75t_SL g875 ( 
.A(n_781),
.B(n_757),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_801),
.B(n_803),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_819),
.Y(n_877)
);

O2A1O1Ixp33_ASAP7_75t_L g878 ( 
.A1(n_825),
.A2(n_771),
.B(n_815),
.C(n_774),
.Y(n_878)
);

AND2x2_ASAP7_75t_L g879 ( 
.A(n_810),
.B(n_813),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_802),
.Y(n_880)
);

AO21x2_ASAP7_75t_L g881 ( 
.A1(n_833),
.A2(n_822),
.B(n_828),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_804),
.Y(n_882)
);

INVx2_ASAP7_75t_L g883 ( 
.A(n_830),
.Y(n_883)
);

INVx2_ASAP7_75t_L g884 ( 
.A(n_778),
.Y(n_884)
);

OAI22xp5_ASAP7_75t_L g885 ( 
.A1(n_756),
.A2(n_781),
.B1(n_757),
.B2(n_846),
.Y(n_885)
);

INVx3_ASAP7_75t_L g886 ( 
.A(n_778),
.Y(n_886)
);

AO21x2_ASAP7_75t_L g887 ( 
.A1(n_822),
.A2(n_828),
.B(n_827),
.Y(n_887)
);

INVx2_ASAP7_75t_L g888 ( 
.A(n_782),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_805),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_827),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_832),
.Y(n_891)
);

BUFx3_ASAP7_75t_L g892 ( 
.A(n_786),
.Y(n_892)
);

HB1xp67_ASAP7_75t_L g893 ( 
.A(n_789),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_832),
.Y(n_894)
);

INVx4_ASAP7_75t_L g895 ( 
.A(n_835),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_785),
.Y(n_896)
);

BUFx6f_ASAP7_75t_L g897 ( 
.A(n_779),
.Y(n_897)
);

CKINVDCx5p33_ASAP7_75t_R g898 ( 
.A(n_844),
.Y(n_898)
);

OAI22xp5_ASAP7_75t_L g899 ( 
.A1(n_846),
.A2(n_796),
.B1(n_811),
.B2(n_789),
.Y(n_899)
);

BUFx2_ASAP7_75t_L g900 ( 
.A(n_787),
.Y(n_900)
);

CKINVDCx6p67_ASAP7_75t_R g901 ( 
.A(n_779),
.Y(n_901)
);

INVx2_ASAP7_75t_SL g902 ( 
.A(n_812),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_831),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_SL g904 ( 
.A(n_820),
.B(n_755),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_784),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_L g906 ( 
.A(n_807),
.B(n_816),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_829),
.Y(n_907)
);

BUFx4f_ASAP7_75t_SL g908 ( 
.A(n_809),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_826),
.Y(n_909)
);

BUFx3_ASAP7_75t_L g910 ( 
.A(n_812),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_793),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_818),
.Y(n_912)
);

INVx2_ASAP7_75t_L g913 ( 
.A(n_823),
.Y(n_913)
);

HB1xp67_ASAP7_75t_L g914 ( 
.A(n_794),
.Y(n_914)
);

HB1xp67_ASAP7_75t_L g915 ( 
.A(n_834),
.Y(n_915)
);

INVx2_ASAP7_75t_L g916 ( 
.A(n_764),
.Y(n_916)
);

CKINVDCx20_ASAP7_75t_R g917 ( 
.A(n_814),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_758),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_772),
.Y(n_919)
);

AND2x2_ASAP7_75t_L g920 ( 
.A(n_848),
.B(n_769),
.Y(n_920)
);

BUFx2_ASAP7_75t_L g921 ( 
.A(n_847),
.Y(n_921)
);

BUFx2_ASAP7_75t_L g922 ( 
.A(n_859),
.Y(n_922)
);

INVxp67_ASAP7_75t_L g923 ( 
.A(n_860),
.Y(n_923)
);

INVxp67_ASAP7_75t_L g924 ( 
.A(n_855),
.Y(n_924)
);

AND2x2_ASAP7_75t_L g925 ( 
.A(n_864),
.B(n_752),
.Y(n_925)
);

HB1xp67_ASAP7_75t_L g926 ( 
.A(n_883),
.Y(n_926)
);

AND2x2_ASAP7_75t_L g927 ( 
.A(n_879),
.B(n_773),
.Y(n_927)
);

OR2x2_ASAP7_75t_L g928 ( 
.A(n_876),
.B(n_790),
.Y(n_928)
);

AND2x2_ASAP7_75t_L g929 ( 
.A(n_877),
.B(n_834),
.Y(n_929)
);

INVxp67_ASAP7_75t_L g930 ( 
.A(n_855),
.Y(n_930)
);

BUFx3_ASAP7_75t_L g931 ( 
.A(n_892),
.Y(n_931)
);

BUFx2_ASAP7_75t_L g932 ( 
.A(n_869),
.Y(n_932)
);

INVx1_ASAP7_75t_L g933 ( 
.A(n_850),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_L g934 ( 
.A(n_852),
.B(n_754),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_L g935 ( 
.A(n_889),
.B(n_762),
.Y(n_935)
);

OR2x2_ASAP7_75t_L g936 ( 
.A(n_876),
.B(n_768),
.Y(n_936)
);

AND2x2_ASAP7_75t_L g937 ( 
.A(n_873),
.B(n_798),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_851),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_853),
.Y(n_939)
);

AND2x2_ASAP7_75t_L g940 ( 
.A(n_873),
.B(n_760),
.Y(n_940)
);

BUFx6f_ASAP7_75t_L g941 ( 
.A(n_910),
.Y(n_941)
);

INVx1_ASAP7_75t_L g942 ( 
.A(n_854),
.Y(n_942)
);

AND2x2_ASAP7_75t_L g943 ( 
.A(n_868),
.B(n_821),
.Y(n_943)
);

INVx3_ASAP7_75t_L g944 ( 
.A(n_881),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_L g945 ( 
.A(n_872),
.B(n_919),
.Y(n_945)
);

AND2x2_ASAP7_75t_L g946 ( 
.A(n_872),
.B(n_862),
.Y(n_946)
);

INVx3_ASAP7_75t_L g947 ( 
.A(n_881),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_L g948 ( 
.A(n_918),
.B(n_858),
.Y(n_948)
);

BUFx3_ASAP7_75t_L g949 ( 
.A(n_892),
.Y(n_949)
);

OR2x2_ASAP7_75t_L g950 ( 
.A(n_869),
.B(n_856),
.Y(n_950)
);

INVx2_ASAP7_75t_L g951 ( 
.A(n_857),
.Y(n_951)
);

BUFx2_ASAP7_75t_L g952 ( 
.A(n_849),
.Y(n_952)
);

INVxp67_ASAP7_75t_SL g953 ( 
.A(n_903),
.Y(n_953)
);

INVx5_ASAP7_75t_SL g954 ( 
.A(n_901),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_L g955 ( 
.A(n_878),
.B(n_906),
.Y(n_955)
);

INVx1_ASAP7_75t_L g956 ( 
.A(n_890),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_891),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_L g958 ( 
.A(n_878),
.B(n_906),
.Y(n_958)
);

AND2x2_ASAP7_75t_L g959 ( 
.A(n_914),
.B(n_880),
.Y(n_959)
);

INVx2_ASAP7_75t_L g960 ( 
.A(n_887),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_894),
.Y(n_961)
);

INVx2_ASAP7_75t_L g962 ( 
.A(n_887),
.Y(n_962)
);

OR2x2_ASAP7_75t_L g963 ( 
.A(n_893),
.B(n_882),
.Y(n_963)
);

AND2x2_ASAP7_75t_L g964 ( 
.A(n_899),
.B(n_866),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_L g965 ( 
.A(n_893),
.B(n_904),
.Y(n_965)
);

AND2x2_ASAP7_75t_L g966 ( 
.A(n_914),
.B(n_884),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_L g967 ( 
.A(n_904),
.B(n_861),
.Y(n_967)
);

AND2x2_ASAP7_75t_L g968 ( 
.A(n_888),
.B(n_861),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_L g969 ( 
.A(n_910),
.B(n_908),
.Y(n_969)
);

AND2x4_ASAP7_75t_SL g970 ( 
.A(n_871),
.B(n_895),
.Y(n_970)
);

BUFx3_ASAP7_75t_L g971 ( 
.A(n_871),
.Y(n_971)
);

INVxp67_ASAP7_75t_L g972 ( 
.A(n_870),
.Y(n_972)
);

AND2x2_ASAP7_75t_L g973 ( 
.A(n_886),
.B(n_902),
.Y(n_973)
);

BUFx3_ASAP7_75t_L g974 ( 
.A(n_865),
.Y(n_974)
);

CKINVDCx5p33_ASAP7_75t_R g975 ( 
.A(n_867),
.Y(n_975)
);

BUFx2_ASAP7_75t_L g976 ( 
.A(n_908),
.Y(n_976)
);

INVx2_ASAP7_75t_SL g977 ( 
.A(n_897),
.Y(n_977)
);

OAI22xp5_ASAP7_75t_L g978 ( 
.A1(n_913),
.A2(n_917),
.B1(n_911),
.B2(n_885),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_909),
.Y(n_979)
);

AND2x2_ASAP7_75t_L g980 ( 
.A(n_929),
.B(n_896),
.Y(n_980)
);

INVxp67_ASAP7_75t_L g981 ( 
.A(n_932),
.Y(n_981)
);

INVx1_ASAP7_75t_L g982 ( 
.A(n_956),
.Y(n_982)
);

INVx1_ASAP7_75t_L g983 ( 
.A(n_957),
.Y(n_983)
);

BUFx2_ASAP7_75t_L g984 ( 
.A(n_921),
.Y(n_984)
);

AOI22xp5_ASAP7_75t_L g985 ( 
.A1(n_967),
.A2(n_917),
.B1(n_867),
.B2(n_900),
.Y(n_985)
);

AOI22xp5_ASAP7_75t_L g986 ( 
.A1(n_925),
.A2(n_874),
.B1(n_898),
.B2(n_885),
.Y(n_986)
);

INVxp67_ASAP7_75t_SL g987 ( 
.A(n_924),
.Y(n_987)
);

INVx1_ASAP7_75t_L g988 ( 
.A(n_961),
.Y(n_988)
);

INVx1_ASAP7_75t_L g989 ( 
.A(n_953),
.Y(n_989)
);

AND2x2_ASAP7_75t_L g990 ( 
.A(n_964),
.B(n_905),
.Y(n_990)
);

BUFx2_ASAP7_75t_L g991 ( 
.A(n_922),
.Y(n_991)
);

INVx1_ASAP7_75t_L g992 ( 
.A(n_979),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_933),
.Y(n_993)
);

HB1xp67_ASAP7_75t_L g994 ( 
.A(n_924),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_938),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_L g996 ( 
.A(n_945),
.B(n_870),
.Y(n_996)
);

HB1xp67_ASAP7_75t_L g997 ( 
.A(n_930),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_L g998 ( 
.A(n_955),
.B(n_915),
.Y(n_998)
);

OR2x2_ASAP7_75t_L g999 ( 
.A(n_965),
.B(n_915),
.Y(n_999)
);

OR2x2_ASAP7_75t_L g1000 ( 
.A(n_936),
.B(n_863),
.Y(n_1000)
);

OR2x2_ASAP7_75t_L g1001 ( 
.A(n_960),
.B(n_863),
.Y(n_1001)
);

NOR2xp33_ASAP7_75t_L g1002 ( 
.A(n_958),
.B(n_907),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_L g1003 ( 
.A(n_930),
.B(n_920),
.Y(n_1003)
);

INVxp67_ASAP7_75t_SL g1004 ( 
.A(n_926),
.Y(n_1004)
);

INVx1_ASAP7_75t_SL g1005 ( 
.A(n_968),
.Y(n_1005)
);

OR2x2_ASAP7_75t_L g1006 ( 
.A(n_950),
.B(n_912),
.Y(n_1006)
);

AND2x2_ASAP7_75t_L g1007 ( 
.A(n_946),
.B(n_875),
.Y(n_1007)
);

INVxp67_ASAP7_75t_L g1008 ( 
.A(n_952),
.Y(n_1008)
);

AND2x2_ASAP7_75t_L g1009 ( 
.A(n_940),
.B(n_875),
.Y(n_1009)
);

INVx1_ASAP7_75t_L g1010 ( 
.A(n_951),
.Y(n_1010)
);

INVx4_ASAP7_75t_R g1011 ( 
.A(n_971),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_SL g1012 ( 
.A(n_934),
.B(n_916),
.Y(n_1012)
);

INVx1_ASAP7_75t_SL g1013 ( 
.A(n_966),
.Y(n_1013)
);

NOR2xp33_ASAP7_75t_L g1014 ( 
.A(n_948),
.B(n_928),
.Y(n_1014)
);

OR2x6_ASAP7_75t_SL g1015 ( 
.A(n_978),
.B(n_898),
.Y(n_1015)
);

OR2x2_ASAP7_75t_L g1016 ( 
.A(n_1000),
.B(n_960),
.Y(n_1016)
);

INVxp67_ASAP7_75t_L g1017 ( 
.A(n_984),
.Y(n_1017)
);

INVxp67_ASAP7_75t_L g1018 ( 
.A(n_994),
.Y(n_1018)
);

INVx1_ASAP7_75t_L g1019 ( 
.A(n_992),
.Y(n_1019)
);

INVxp67_ASAP7_75t_SL g1020 ( 
.A(n_1004),
.Y(n_1020)
);

NAND2xp5_ASAP7_75t_L g1021 ( 
.A(n_1014),
.B(n_935),
.Y(n_1021)
);

INVx1_ASAP7_75t_L g1022 ( 
.A(n_989),
.Y(n_1022)
);

INVx2_ASAP7_75t_L g1023 ( 
.A(n_1010),
.Y(n_1023)
);

OR2x2_ASAP7_75t_L g1024 ( 
.A(n_1000),
.B(n_962),
.Y(n_1024)
);

NAND2xp5_ASAP7_75t_L g1025 ( 
.A(n_1014),
.B(n_939),
.Y(n_1025)
);

OR2x2_ASAP7_75t_L g1026 ( 
.A(n_999),
.B(n_944),
.Y(n_1026)
);

NAND2xp5_ASAP7_75t_SL g1027 ( 
.A(n_1002),
.B(n_943),
.Y(n_1027)
);

AND2x2_ASAP7_75t_L g1028 ( 
.A(n_1009),
.B(n_944),
.Y(n_1028)
);

AND2x2_ASAP7_75t_L g1029 ( 
.A(n_1009),
.B(n_944),
.Y(n_1029)
);

AND2x2_ASAP7_75t_L g1030 ( 
.A(n_1007),
.B(n_947),
.Y(n_1030)
);

AND2x2_ASAP7_75t_L g1031 ( 
.A(n_1007),
.B(n_980),
.Y(n_1031)
);

INVx1_ASAP7_75t_L g1032 ( 
.A(n_982),
.Y(n_1032)
);

HB1xp67_ASAP7_75t_L g1033 ( 
.A(n_997),
.Y(n_1033)
);

OR2x2_ASAP7_75t_L g1034 ( 
.A(n_1006),
.B(n_1001),
.Y(n_1034)
);

NAND2xp5_ASAP7_75t_L g1035 ( 
.A(n_987),
.B(n_942),
.Y(n_1035)
);

NOR2xp33_ASAP7_75t_L g1036 ( 
.A(n_1005),
.B(n_976),
.Y(n_1036)
);

INVxp67_ASAP7_75t_SL g1037 ( 
.A(n_1012),
.Y(n_1037)
);

INVx1_ASAP7_75t_L g1038 ( 
.A(n_983),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_988),
.Y(n_1039)
);

OR2x2_ASAP7_75t_L g1040 ( 
.A(n_1003),
.B(n_963),
.Y(n_1040)
);

INVx1_ASAP7_75t_L g1041 ( 
.A(n_993),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_995),
.Y(n_1042)
);

INVx2_ASAP7_75t_L g1043 ( 
.A(n_1019),
.Y(n_1043)
);

HB1xp67_ASAP7_75t_L g1044 ( 
.A(n_1016),
.Y(n_1044)
);

AND2x2_ASAP7_75t_L g1045 ( 
.A(n_1031),
.B(n_991),
.Y(n_1045)
);

OAI21xp33_ASAP7_75t_L g1046 ( 
.A1(n_1027),
.A2(n_986),
.B(n_1002),
.Y(n_1046)
);

OR2x2_ASAP7_75t_L g1047 ( 
.A(n_1034),
.B(n_1031),
.Y(n_1047)
);

AND2x2_ASAP7_75t_L g1048 ( 
.A(n_1030),
.B(n_1028),
.Y(n_1048)
);

CKINVDCx16_ASAP7_75t_R g1049 ( 
.A(n_1036),
.Y(n_1049)
);

AOI21xp33_ASAP7_75t_L g1050 ( 
.A1(n_1021),
.A2(n_998),
.B(n_996),
.Y(n_1050)
);

NOR2x1_ASAP7_75t_L g1051 ( 
.A(n_1025),
.B(n_1012),
.Y(n_1051)
);

OR2x2_ASAP7_75t_L g1052 ( 
.A(n_1026),
.B(n_1013),
.Y(n_1052)
);

INVx1_ASAP7_75t_L g1053 ( 
.A(n_1032),
.Y(n_1053)
);

INVx4_ASAP7_75t_L g1054 ( 
.A(n_1033),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_1038),
.Y(n_1055)
);

NAND2xp5_ASAP7_75t_L g1056 ( 
.A(n_1037),
.B(n_990),
.Y(n_1056)
);

OR2x2_ASAP7_75t_L g1057 ( 
.A(n_1024),
.B(n_981),
.Y(n_1057)
);

INVx2_ASAP7_75t_L g1058 ( 
.A(n_1023),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_1039),
.Y(n_1059)
);

INVx2_ASAP7_75t_L g1060 ( 
.A(n_1041),
.Y(n_1060)
);

INVx1_ASAP7_75t_L g1061 ( 
.A(n_1042),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_L g1062 ( 
.A(n_1044),
.B(n_1020),
.Y(n_1062)
);

INVx1_ASAP7_75t_L g1063 ( 
.A(n_1053),
.Y(n_1063)
);

NAND2xp5_ASAP7_75t_L g1064 ( 
.A(n_1050),
.B(n_1018),
.Y(n_1064)
);

INVx1_ASAP7_75t_L g1065 ( 
.A(n_1055),
.Y(n_1065)
);

INVx1_ASAP7_75t_L g1066 ( 
.A(n_1059),
.Y(n_1066)
);

INVx1_ASAP7_75t_L g1067 ( 
.A(n_1061),
.Y(n_1067)
);

INVx1_ASAP7_75t_L g1068 ( 
.A(n_1058),
.Y(n_1068)
);

AOI22xp33_ASAP7_75t_L g1069 ( 
.A1(n_1046),
.A2(n_1027),
.B1(n_927),
.B2(n_937),
.Y(n_1069)
);

AND2x2_ASAP7_75t_L g1070 ( 
.A(n_1048),
.B(n_1029),
.Y(n_1070)
);

NOR2xp67_ASAP7_75t_L g1071 ( 
.A(n_1054),
.B(n_1017),
.Y(n_1071)
);

INVx1_ASAP7_75t_L g1072 ( 
.A(n_1043),
.Y(n_1072)
);

INVx1_ASAP7_75t_L g1073 ( 
.A(n_1060),
.Y(n_1073)
);

INVx1_ASAP7_75t_L g1074 ( 
.A(n_1044),
.Y(n_1074)
);

OAI21xp33_ASAP7_75t_L g1075 ( 
.A1(n_1046),
.A2(n_1035),
.B(n_1029),
.Y(n_1075)
);

NAND2xp5_ASAP7_75t_L g1076 ( 
.A(n_1056),
.B(n_1022),
.Y(n_1076)
);

OAI22xp33_ASAP7_75t_L g1077 ( 
.A1(n_1049),
.A2(n_1015),
.B1(n_985),
.B2(n_1040),
.Y(n_1077)
);

OAI21xp5_ASAP7_75t_SL g1078 ( 
.A1(n_1069),
.A2(n_970),
.B(n_1050),
.Y(n_1078)
);

INVx1_ASAP7_75t_L g1079 ( 
.A(n_1063),
.Y(n_1079)
);

AOI22xp5_ASAP7_75t_L g1080 ( 
.A1(n_1075),
.A2(n_1051),
.B1(n_1056),
.B2(n_1054),
.Y(n_1080)
);

INVx1_ASAP7_75t_L g1081 ( 
.A(n_1065),
.Y(n_1081)
);

NAND2xp5_ASAP7_75t_L g1082 ( 
.A(n_1064),
.B(n_1045),
.Y(n_1082)
);

AOI21xp33_ASAP7_75t_SL g1083 ( 
.A1(n_1077),
.A2(n_975),
.B(n_874),
.Y(n_1083)
);

OAI221xp5_ASAP7_75t_L g1084 ( 
.A1(n_1071),
.A2(n_1076),
.B1(n_1062),
.B2(n_1057),
.C(n_1066),
.Y(n_1084)
);

INVx1_ASAP7_75t_SL g1085 ( 
.A(n_1062),
.Y(n_1085)
);

NAND2xp5_ASAP7_75t_L g1086 ( 
.A(n_1080),
.B(n_1085),
.Y(n_1086)
);

OAI21xp5_ASAP7_75t_L g1087 ( 
.A1(n_1083),
.A2(n_1076),
.B(n_1067),
.Y(n_1087)
);

O2A1O1Ixp33_ASAP7_75t_SL g1088 ( 
.A1(n_1084),
.A2(n_1074),
.B(n_1011),
.C(n_1008),
.Y(n_1088)
);

NOR3xp33_ASAP7_75t_SL g1089 ( 
.A(n_1078),
.B(n_975),
.C(n_969),
.Y(n_1089)
);

NAND2xp5_ASAP7_75t_L g1090 ( 
.A(n_1082),
.B(n_1070),
.Y(n_1090)
);

XNOR2xp5_ASAP7_75t_L g1091 ( 
.A(n_1089),
.B(n_970),
.Y(n_1091)
);

NAND2xp5_ASAP7_75t_SL g1092 ( 
.A(n_1087),
.B(n_1079),
.Y(n_1092)
);

AOI221xp5_ASAP7_75t_SL g1093 ( 
.A1(n_1086),
.A2(n_1081),
.B1(n_1073),
.B2(n_1072),
.C(n_923),
.Y(n_1093)
);

NAND2xp5_ASAP7_75t_SL g1094 ( 
.A(n_1090),
.B(n_1052),
.Y(n_1094)
);

INVx1_ASAP7_75t_L g1095 ( 
.A(n_1088),
.Y(n_1095)
);

OR2x2_ASAP7_75t_L g1096 ( 
.A(n_1086),
.B(n_1047),
.Y(n_1096)
);

NAND2xp5_ASAP7_75t_L g1097 ( 
.A(n_1093),
.B(n_1068),
.Y(n_1097)
);

OA211x2_ASAP7_75t_L g1098 ( 
.A1(n_1092),
.A2(n_923),
.B(n_972),
.C(n_954),
.Y(n_1098)
);

NOR2x1_ASAP7_75t_L g1099 ( 
.A(n_1095),
.B(n_971),
.Y(n_1099)
);

NOR3x1_ASAP7_75t_L g1100 ( 
.A(n_1097),
.B(n_1096),
.C(n_1094),
.Y(n_1100)
);

INVx1_ASAP7_75t_L g1101 ( 
.A(n_1099),
.Y(n_1101)
);

INVx1_ASAP7_75t_L g1102 ( 
.A(n_1101),
.Y(n_1102)
);

OAI22xp5_ASAP7_75t_L g1103 ( 
.A1(n_1102),
.A2(n_1098),
.B1(n_1091),
.B2(n_1100),
.Y(n_1103)
);

CKINVDCx20_ASAP7_75t_R g1104 ( 
.A(n_1103),
.Y(n_1104)
);

OAI21xp5_ASAP7_75t_L g1105 ( 
.A1(n_1104),
.A2(n_949),
.B(n_931),
.Y(n_1105)
);

OAI21xp5_ASAP7_75t_L g1106 ( 
.A1(n_1105),
.A2(n_974),
.B(n_959),
.Y(n_1106)
);

NAND2xp5_ASAP7_75t_L g1107 ( 
.A(n_1106),
.B(n_954),
.Y(n_1107)
);

OAI22xp33_ASAP7_75t_L g1108 ( 
.A1(n_1107),
.A2(n_941),
.B1(n_1015),
.B2(n_977),
.Y(n_1108)
);

NAND2xp5_ASAP7_75t_SL g1109 ( 
.A(n_1108),
.B(n_941),
.Y(n_1109)
);

AO21x2_ASAP7_75t_L g1110 ( 
.A1(n_1109),
.A2(n_973),
.B(n_972),
.Y(n_1110)
);


endmodule