module real_jpeg_31699_n_6 (n_5, n_4, n_0, n_1, n_2, n_3, n_6);

input n_5;
input n_4;
input n_0;
input n_1;
input n_2;
input n_3;

output n_6;

wire n_17;
wire n_8;
wire n_37;
wire n_21;
wire n_35;
wire n_38;
wire n_33;
wire n_29;
wire n_10;
wire n_31;
wire n_9;
wire n_12;
wire n_24;
wire n_34;
wire n_28;
wire n_23;
wire n_11;
wire n_14;
wire n_25;
wire n_7;
wire n_22;
wire n_18;
wire n_36;
wire n_40;
wire n_39;
wire n_26;
wire n_27;
wire n_20;
wire n_19;
wire n_32;
wire n_30;
wire n_16;
wire n_15;
wire n_13;

OR2x2_ASAP7_75t_L g17 ( 
.A(n_0),
.B(n_18),
.Y(n_17)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

BUFx2_ASAP7_75t_R g13 ( 
.A(n_1),
.Y(n_13)
);

NAND2x1p5_ASAP7_75t_L g23 ( 
.A(n_1),
.B(n_24),
.Y(n_23)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

INVx4_ASAP7_75t_L g12 ( 
.A(n_2),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g16 ( 
.A(n_2),
.B(n_9),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_SL g27 ( 
.A(n_2),
.B(n_22),
.Y(n_27)
);

INVx2_ASAP7_75t_L g9 ( 
.A(n_3),
.Y(n_9)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_3),
.B(n_12),
.Y(n_39)
);

AO21x1_ASAP7_75t_L g22 ( 
.A1(n_4),
.A2(n_23),
.B(n_25),
.Y(n_22)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

AND2x2_ASAP7_75t_L g25 ( 
.A(n_5),
.B(n_26),
.Y(n_25)
);

AOI221xp5_ASAP7_75t_L g6 ( 
.A1(n_7),
.A2(n_19),
.B1(n_28),
.B2(n_35),
.C(n_36),
.Y(n_6)
);

NAND2xp5_ASAP7_75t_SL g7 ( 
.A(n_8),
.B(n_17),
.Y(n_7)
);

AOI22xp5_ASAP7_75t_L g8 ( 
.A1(n_9),
.A2(n_10),
.B1(n_14),
.B2(n_15),
.Y(n_8)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_9),
.B(n_12),
.Y(n_40)
);

INVx1_ASAP7_75t_L g10 ( 
.A(n_11),
.Y(n_10)
);

OAI21xp5_ASAP7_75t_L g31 ( 
.A1(n_11),
.A2(n_12),
.B(n_13),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_SL g11 ( 
.A(n_12),
.B(n_13),
.Y(n_11)
);

NAND2xp67_ASAP7_75t_SL g20 ( 
.A(n_12),
.B(n_21),
.Y(n_20)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_13),
.Y(n_14)
);

AOI22xp5_ASAP7_75t_L g37 ( 
.A1(n_13),
.A2(n_14),
.B1(n_38),
.B2(n_40),
.Y(n_37)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_16),
.Y(n_15)
);

AND2x2_ASAP7_75t_L g33 ( 
.A(n_18),
.B(n_34),
.Y(n_33)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_19),
.Y(n_35)
);

NAND2x1_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_27),
.Y(n_19)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

OAI21xp5_ASAP7_75t_L g28 ( 
.A1(n_29),
.A2(n_30),
.B(n_32),
.Y(n_28)
);

INVx2_ASAP7_75t_R g34 ( 
.A(n_29),
.Y(n_34)
);

CKINVDCx16_ASAP7_75t_R g30 ( 
.A(n_31),
.Y(n_30)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_34),
.B(n_37),
.Y(n_36)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);


endmodule