module fake_jpeg_12404_n_611 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_611);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_611;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_19;
wire n_182;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_579;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_349;
wire n_21;
wire n_393;
wire n_288;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_442;
wire n_299;
wire n_300;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_599;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_10),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_14),
.B(n_6),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_5),
.Y(n_21)
);

CKINVDCx14_ASAP7_75t_R g22 ( 
.A(n_4),
.Y(n_22)
);

INVx6_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

BUFx8_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_15),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_13),
.Y(n_28)
);

INVx11_ASAP7_75t_SL g29 ( 
.A(n_10),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

BUFx4f_ASAP7_75t_L g35 ( 
.A(n_12),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_6),
.Y(n_36)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_4),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_10),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_11),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_11),
.Y(n_40)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_16),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_15),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_8),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_16),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_9),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_1),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_5),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_14),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_12),
.Y(n_49)
);

INVx2_ASAP7_75t_SL g50 ( 
.A(n_5),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_1),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_15),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_6),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_2),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_2),
.Y(n_55)
);

BUFx5_ASAP7_75t_L g56 ( 
.A(n_6),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_11),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_5),
.Y(n_58)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_37),
.Y(n_59)
);

INVx5_ASAP7_75t_L g176 ( 
.A(n_59),
.Y(n_176)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_60),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_18),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_61),
.Y(n_126)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_26),
.Y(n_62)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_62),
.Y(n_132)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_49),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g165 ( 
.A(n_63),
.Y(n_165)
);

AND2x2_ASAP7_75t_L g64 ( 
.A(n_20),
.B(n_8),
.Y(n_64)
);

AND2x2_ASAP7_75t_L g152 ( 
.A(n_64),
.B(n_51),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_18),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_65),
.Y(n_127)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_49),
.Y(n_66)
);

BUFx12f_ASAP7_75t_L g174 ( 
.A(n_66),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_20),
.B(n_9),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_67),
.B(n_58),
.Y(n_125)
);

BUFx12f_ASAP7_75t_L g68 ( 
.A(n_24),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g131 ( 
.A(n_68),
.Y(n_131)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_49),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g137 ( 
.A(n_69),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_18),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_70),
.Y(n_144)
);

INVx2_ASAP7_75t_SL g71 ( 
.A(n_31),
.Y(n_71)
);

BUFx3_ASAP7_75t_L g138 ( 
.A(n_71),
.Y(n_138)
);

BUFx8_ASAP7_75t_L g72 ( 
.A(n_29),
.Y(n_72)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_72),
.Y(n_128)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_24),
.Y(n_73)
);

INVx3_ASAP7_75t_L g160 ( 
.A(n_73),
.Y(n_160)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_40),
.Y(n_74)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_74),
.Y(n_133)
);

INVx6_ASAP7_75t_SL g75 ( 
.A(n_24),
.Y(n_75)
);

CKINVDCx5p33_ASAP7_75t_R g150 ( 
.A(n_75),
.Y(n_150)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_26),
.Y(n_76)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_76),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_35),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_77),
.B(n_83),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_33),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_78),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_33),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_79),
.Y(n_156)
);

INVx11_ASAP7_75t_L g80 ( 
.A(n_31),
.Y(n_80)
);

INVx11_ASAP7_75t_L g134 ( 
.A(n_80),
.Y(n_134)
);

BUFx5_ASAP7_75t_L g81 ( 
.A(n_37),
.Y(n_81)
);

BUFx5_ASAP7_75t_L g169 ( 
.A(n_81),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_32),
.B(n_50),
.C(n_57),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_82),
.B(n_47),
.C(n_53),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_35),
.Y(n_83)
);

BUFx3_ASAP7_75t_L g84 ( 
.A(n_49),
.Y(n_84)
);

BUFx3_ASAP7_75t_L g167 ( 
.A(n_84),
.Y(n_167)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_35),
.Y(n_85)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_85),
.Y(n_136)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_27),
.Y(n_86)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_86),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_33),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_87),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_36),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g180 ( 
.A(n_88),
.Y(n_180)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_35),
.Y(n_89)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_89),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_36),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g196 ( 
.A(n_90),
.Y(n_196)
);

BUFx5_ASAP7_75t_L g91 ( 
.A(n_56),
.Y(n_91)
);

INVx4_ASAP7_75t_L g124 ( 
.A(n_91),
.Y(n_124)
);

BUFx5_ASAP7_75t_L g92 ( 
.A(n_56),
.Y(n_92)
);

INVx4_ASAP7_75t_L g143 ( 
.A(n_92),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_36),
.Y(n_93)
);

INVx6_ASAP7_75t_L g145 ( 
.A(n_93),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_39),
.Y(n_94)
);

INVx6_ASAP7_75t_L g168 ( 
.A(n_94),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_17),
.B(n_9),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_95),
.B(n_13),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_39),
.Y(n_96)
);

INVx6_ASAP7_75t_L g182 ( 
.A(n_96),
.Y(n_182)
);

INVx11_ASAP7_75t_L g97 ( 
.A(n_24),
.Y(n_97)
);

CKINVDCx14_ASAP7_75t_R g187 ( 
.A(n_97),
.Y(n_187)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_27),
.Y(n_98)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_98),
.Y(n_186)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_41),
.Y(n_99)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_99),
.Y(n_163)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_30),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_100),
.B(n_104),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_39),
.Y(n_101)
);

INVx8_ASAP7_75t_L g140 ( 
.A(n_101),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_52),
.Y(n_102)
);

INVx8_ASAP7_75t_L g151 ( 
.A(n_102),
.Y(n_151)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_41),
.Y(n_103)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_103),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_41),
.Y(n_104)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_32),
.Y(n_105)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_105),
.Y(n_185)
);

BUFx3_ASAP7_75t_L g106 ( 
.A(n_19),
.Y(n_106)
);

INVx5_ASAP7_75t_L g172 ( 
.A(n_106),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_52),
.Y(n_107)
);

INVx8_ASAP7_75t_L g155 ( 
.A(n_107),
.Y(n_155)
);

INVx2_ASAP7_75t_SL g108 ( 
.A(n_19),
.Y(n_108)
);

HB1xp67_ASAP7_75t_L g142 ( 
.A(n_108),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_30),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_109),
.B(n_110),
.Y(n_164)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_38),
.Y(n_110)
);

BUFx16f_ASAP7_75t_L g111 ( 
.A(n_19),
.Y(n_111)
);

INVx4_ASAP7_75t_SL g188 ( 
.A(n_111),
.Y(n_188)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_19),
.Y(n_112)
);

INVx3_ASAP7_75t_L g162 ( 
.A(n_112),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_52),
.Y(n_113)
);

INVx8_ASAP7_75t_L g158 ( 
.A(n_113),
.Y(n_158)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_38),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_114),
.B(n_117),
.Y(n_173)
);

INVx11_ASAP7_75t_L g115 ( 
.A(n_50),
.Y(n_115)
);

INVx8_ASAP7_75t_L g166 ( 
.A(n_115),
.Y(n_166)
);

BUFx3_ASAP7_75t_L g116 ( 
.A(n_19),
.Y(n_116)
);

INVx5_ASAP7_75t_L g191 ( 
.A(n_116),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_42),
.Y(n_117)
);

BUFx3_ASAP7_75t_L g118 ( 
.A(n_55),
.Y(n_118)
);

INVx4_ASAP7_75t_L g170 ( 
.A(n_118),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_57),
.Y(n_119)
);

INVx8_ASAP7_75t_L g195 ( 
.A(n_119),
.Y(n_195)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_55),
.Y(n_120)
);

INVx3_ASAP7_75t_L g171 ( 
.A(n_120),
.Y(n_171)
);

BUFx5_ASAP7_75t_L g121 ( 
.A(n_57),
.Y(n_121)
);

INVx4_ASAP7_75t_L g193 ( 
.A(n_121),
.Y(n_193)
);

INVx4_ASAP7_75t_L g122 ( 
.A(n_55),
.Y(n_122)
);

INVx3_ASAP7_75t_L g199 ( 
.A(n_122),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_42),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_123),
.B(n_44),
.Y(n_178)
);

NAND3xp33_ASAP7_75t_L g251 ( 
.A(n_125),
.B(n_192),
.C(n_197),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_SL g139 ( 
.A(n_64),
.B(n_58),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g242 ( 
.A(n_139),
.B(n_146),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_82),
.A2(n_23),
.B1(n_50),
.B2(n_34),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_141),
.A2(n_157),
.B1(n_22),
.B2(n_54),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_SL g146 ( 
.A(n_68),
.B(n_17),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_149),
.B(n_154),
.Y(n_221)
);

AND2x2_ASAP7_75t_L g212 ( 
.A(n_152),
.B(n_153),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_60),
.B(n_45),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_61),
.A2(n_23),
.B1(n_45),
.B2(n_44),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g161 ( 
.A(n_75),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_161),
.B(n_178),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_111),
.B(n_21),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_179),
.B(n_181),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_99),
.B(n_28),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_111),
.B(n_21),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_183),
.B(n_189),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_115),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_68),
.B(n_25),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_190),
.B(n_198),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_103),
.B(n_28),
.Y(n_192)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_112),
.Y(n_194)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_194),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_108),
.B(n_25),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_63),
.B(n_53),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_66),
.B(n_48),
.Y(n_200)
);

AND2x2_ASAP7_75t_L g226 ( 
.A(n_200),
.B(n_72),
.Y(n_226)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_120),
.Y(n_201)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_201),
.Y(n_222)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_122),
.Y(n_202)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_202),
.Y(n_246)
);

AOI22xp33_ASAP7_75t_SL g204 ( 
.A1(n_150),
.A2(n_59),
.B1(n_34),
.B2(n_71),
.Y(n_204)
);

AOI22xp33_ASAP7_75t_SL g309 ( 
.A1(n_204),
.A2(n_208),
.B1(n_216),
.B2(n_243),
.Y(n_309)
);

INVx6_ASAP7_75t_L g205 ( 
.A(n_126),
.Y(n_205)
);

INVx6_ASAP7_75t_L g288 ( 
.A(n_205),
.Y(n_288)
);

INVx8_ASAP7_75t_L g206 ( 
.A(n_126),
.Y(n_206)
);

BUFx2_ASAP7_75t_L g324 ( 
.A(n_206),
.Y(n_324)
);

INVx3_ASAP7_75t_L g207 ( 
.A(n_166),
.Y(n_207)
);

INVx3_ASAP7_75t_L g306 ( 
.A(n_207),
.Y(n_306)
);

AOI22xp33_ASAP7_75t_SL g208 ( 
.A1(n_124),
.A2(n_34),
.B1(n_73),
.B2(n_80),
.Y(n_208)
);

CKINVDCx11_ASAP7_75t_R g209 ( 
.A(n_161),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_209),
.B(n_259),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_164),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_210),
.B(n_214),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_L g280 ( 
.A1(n_211),
.A2(n_213),
.B1(n_233),
.B2(n_269),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_152),
.A2(n_113),
.B1(n_119),
.B2(n_70),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_173),
.Y(n_214)
);

BUFx6f_ASAP7_75t_L g215 ( 
.A(n_127),
.Y(n_215)
);

BUFx6f_ASAP7_75t_L g289 ( 
.A(n_215),
.Y(n_289)
);

AOI22xp33_ASAP7_75t_SL g216 ( 
.A1(n_124),
.A2(n_97),
.B1(n_23),
.B2(n_118),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g217 ( 
.A1(n_132),
.A2(n_79),
.B1(n_78),
.B2(n_107),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_217),
.A2(n_224),
.B1(n_244),
.B2(n_255),
.Y(n_275)
);

INVx3_ASAP7_75t_L g218 ( 
.A(n_166),
.Y(n_218)
);

INVx1_ASAP7_75t_SL g297 ( 
.A(n_218),
.Y(n_297)
);

BUFx6f_ASAP7_75t_L g220 ( 
.A(n_127),
.Y(n_220)
);

BUFx6f_ASAP7_75t_L g295 ( 
.A(n_220),
.Y(n_295)
);

BUFx6f_ASAP7_75t_L g223 ( 
.A(n_144),
.Y(n_223)
);

BUFx6f_ASAP7_75t_L g300 ( 
.A(n_223),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_177),
.A2(n_65),
.B1(n_87),
.B2(n_88),
.Y(n_224)
);

INVx6_ASAP7_75t_L g225 ( 
.A(n_144),
.Y(n_225)
);

INVx6_ASAP7_75t_L g310 ( 
.A(n_225),
.Y(n_310)
);

XNOR2x1_ASAP7_75t_L g286 ( 
.A(n_226),
.B(n_252),
.Y(n_286)
);

BUFx6f_ASAP7_75t_L g227 ( 
.A(n_148),
.Y(n_227)
);

INVx6_ASAP7_75t_L g318 ( 
.A(n_227),
.Y(n_318)
);

INVx4_ASAP7_75t_L g228 ( 
.A(n_165),
.Y(n_228)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_228),
.Y(n_277)
);

INVx11_ASAP7_75t_L g229 ( 
.A(n_134),
.Y(n_229)
);

INVx11_ASAP7_75t_L g278 ( 
.A(n_229),
.Y(n_278)
);

CKINVDCx16_ASAP7_75t_R g230 ( 
.A(n_142),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g291 ( 
.A(n_230),
.B(n_258),
.Y(n_291)
);

BUFx6f_ASAP7_75t_L g231 ( 
.A(n_148),
.Y(n_231)
);

INVx8_ASAP7_75t_L g293 ( 
.A(n_231),
.Y(n_293)
);

BUFx6f_ASAP7_75t_L g232 ( 
.A(n_156),
.Y(n_232)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_232),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_184),
.A2(n_90),
.B1(n_93),
.B2(n_94),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_186),
.Y(n_234)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_234),
.Y(n_276)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_130),
.Y(n_235)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_235),
.Y(n_282)
);

INVx3_ASAP7_75t_L g236 ( 
.A(n_170),
.Y(n_236)
);

INVx1_ASAP7_75t_SL g313 ( 
.A(n_236),
.Y(n_313)
);

INVx6_ASAP7_75t_L g237 ( 
.A(n_156),
.Y(n_237)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_237),
.Y(n_284)
);

INVx5_ASAP7_75t_L g238 ( 
.A(n_193),
.Y(n_238)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_238),
.Y(n_287)
);

INVx11_ASAP7_75t_L g239 ( 
.A(n_134),
.Y(n_239)
);

BUFx24_ASAP7_75t_L g303 ( 
.A(n_239),
.Y(n_303)
);

BUFx6f_ASAP7_75t_L g240 ( 
.A(n_159),
.Y(n_240)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_240),
.Y(n_292)
);

OA22x2_ASAP7_75t_L g241 ( 
.A1(n_185),
.A2(n_96),
.B1(n_102),
.B2(n_101),
.Y(n_241)
);

OA22x2_ASAP7_75t_L g317 ( 
.A1(n_241),
.A2(n_191),
.B1(n_172),
.B2(n_167),
.Y(n_317)
);

AOI22xp33_ASAP7_75t_SL g243 ( 
.A1(n_143),
.A2(n_84),
.B1(n_69),
.B2(n_106),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_L g244 ( 
.A1(n_135),
.A2(n_51),
.B1(n_54),
.B2(n_22),
.Y(n_244)
);

BUFx3_ASAP7_75t_L g245 ( 
.A(n_131),
.Y(n_245)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_245),
.Y(n_298)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_142),
.Y(n_248)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_248),
.Y(n_290)
);

INVx6_ASAP7_75t_L g249 ( 
.A(n_159),
.Y(n_249)
);

INVx2_ASAP7_75t_L g327 ( 
.A(n_249),
.Y(n_327)
);

BUFx12f_ASAP7_75t_L g250 ( 
.A(n_131),
.Y(n_250)
);

INVxp67_ASAP7_75t_L g325 ( 
.A(n_250),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_143),
.A2(n_176),
.B1(n_199),
.B2(n_171),
.Y(n_252)
);

INVx6_ASAP7_75t_L g253 ( 
.A(n_180),
.Y(n_253)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_253),
.Y(n_319)
);

INVx3_ASAP7_75t_L g254 ( 
.A(n_138),
.Y(n_254)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_254),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_L g255 ( 
.A1(n_133),
.A2(n_43),
.B1(n_47),
.B2(n_48),
.Y(n_255)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_136),
.Y(n_256)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_256),
.Y(n_331)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_147),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_257),
.B(n_262),
.Y(n_304)
);

CKINVDCx16_ASAP7_75t_R g258 ( 
.A(n_188),
.Y(n_258)
);

BUFx3_ASAP7_75t_L g259 ( 
.A(n_165),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_L g260 ( 
.A1(n_145),
.A2(n_43),
.B1(n_46),
.B2(n_116),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_260),
.A2(n_187),
.B1(n_128),
.B2(n_195),
.Y(n_281)
);

BUFx3_ASAP7_75t_L g261 ( 
.A(n_165),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_261),
.B(n_265),
.Y(n_312)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_163),
.Y(n_262)
);

O2A1O1Ixp33_ASAP7_75t_L g264 ( 
.A1(n_187),
.A2(n_46),
.B(n_92),
.C(n_91),
.Y(n_264)
);

AOI22x1_ASAP7_75t_L g308 ( 
.A1(n_264),
.A2(n_72),
.B1(n_176),
.B2(n_160),
.Y(n_308)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_175),
.Y(n_265)
);

BUFx12f_ASAP7_75t_L g266 ( 
.A(n_137),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_266),
.B(n_267),
.Y(n_323)
);

AOI21xp33_ASAP7_75t_L g267 ( 
.A1(n_169),
.A2(n_81),
.B(n_12),
.Y(n_267)
);

BUFx5_ASAP7_75t_L g268 ( 
.A(n_188),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_SL g314 ( 
.A(n_268),
.B(n_270),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_145),
.A2(n_121),
.B1(n_11),
.B2(n_13),
.Y(n_269)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_129),
.Y(n_270)
);

INVx6_ASAP7_75t_L g272 ( 
.A(n_180),
.Y(n_272)
);

AOI22xp33_ASAP7_75t_SL g316 ( 
.A1(n_272),
.A2(n_273),
.B1(n_274),
.B2(n_167),
.Y(n_316)
);

INVx6_ASAP7_75t_L g273 ( 
.A(n_196),
.Y(n_273)
);

BUFx6f_ASAP7_75t_L g274 ( 
.A(n_196),
.Y(n_274)
);

AND2x2_ASAP7_75t_L g339 ( 
.A(n_281),
.B(n_301),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_247),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_285),
.B(n_294),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_203),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_212),
.A2(n_182),
.B1(n_168),
.B2(n_195),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_L g361 ( 
.A1(n_296),
.A2(n_305),
.B1(n_315),
.B2(n_320),
.Y(n_361)
);

OAI22xp5_ASAP7_75t_L g299 ( 
.A1(n_221),
.A2(n_168),
.B1(n_182),
.B2(n_151),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g364 ( 
.A1(n_299),
.A2(n_302),
.B1(n_322),
.B2(n_329),
.Y(n_364)
);

AND2x2_ASAP7_75t_SL g301 ( 
.A(n_263),
.B(n_138),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_216),
.A2(n_151),
.B1(n_155),
.B2(n_158),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_212),
.A2(n_140),
.B1(n_158),
.B2(n_155),
.Y(n_305)
);

XOR2xp5_ASAP7_75t_L g307 ( 
.A(n_271),
.B(n_162),
.Y(n_307)
);

XOR2xp5_ASAP7_75t_L g349 ( 
.A(n_307),
.B(n_208),
.Y(n_349)
);

CKINVDCx16_ASAP7_75t_R g345 ( 
.A(n_308),
.Y(n_345)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_241),
.A2(n_140),
.B1(n_170),
.B2(n_193),
.Y(n_315)
);

INVxp67_ASAP7_75t_L g350 ( 
.A(n_316),
.Y(n_350)
);

BUFx2_ASAP7_75t_L g352 ( 
.A(n_317),
.Y(n_352)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_241),
.A2(n_137),
.B1(n_7),
.B2(n_16),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_SL g321 ( 
.A1(n_226),
.A2(n_174),
.B1(n_7),
.B2(n_13),
.Y(n_321)
);

AOI21xp5_ASAP7_75t_SL g346 ( 
.A1(n_321),
.A2(n_328),
.B(n_243),
.Y(n_346)
);

OAI22xp5_ASAP7_75t_L g322 ( 
.A1(n_204),
.A2(n_174),
.B1(n_4),
.B2(n_3),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_246),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_326),
.B(n_236),
.Y(n_341)
);

AOI22xp5_ASAP7_75t_SL g328 ( 
.A1(n_242),
.A2(n_174),
.B1(n_3),
.B2(n_14),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_L g329 ( 
.A1(n_251),
.A2(n_3),
.B1(n_16),
.B2(n_2),
.Y(n_329)
);

AND2x2_ASAP7_75t_SL g332 ( 
.A(n_251),
.B(n_0),
.Y(n_332)
);

CKINVDCx14_ASAP7_75t_R g354 ( 
.A(n_332),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_SL g333 ( 
.A(n_279),
.B(n_222),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_SL g404 ( 
.A(n_333),
.B(n_347),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_307),
.B(n_219),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_335),
.B(n_342),
.Y(n_395)
);

BUFx3_ASAP7_75t_L g336 ( 
.A(n_298),
.Y(n_336)
);

BUFx3_ASAP7_75t_L g392 ( 
.A(n_336),
.Y(n_392)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_306),
.Y(n_337)
);

INVx1_ASAP7_75t_SL g406 ( 
.A(n_337),
.Y(n_406)
);

INVx8_ASAP7_75t_L g338 ( 
.A(n_289),
.Y(n_338)
);

INVx1_ASAP7_75t_SL g409 ( 
.A(n_338),
.Y(n_409)
);

AOI22xp5_ASAP7_75t_SL g340 ( 
.A1(n_302),
.A2(n_264),
.B1(n_218),
.B2(n_207),
.Y(n_340)
);

OAI21xp5_ASAP7_75t_SL g379 ( 
.A1(n_340),
.A2(n_346),
.B(n_350),
.Y(n_379)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_341),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_301),
.B(n_206),
.Y(n_342)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_306),
.Y(n_343)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_343),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_301),
.B(n_237),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_344),
.B(n_348),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_L g347 ( 
.A(n_282),
.B(n_238),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_323),
.B(n_205),
.Y(n_348)
);

XNOR2xp5_ASAP7_75t_L g385 ( 
.A(n_349),
.B(n_362),
.Y(n_385)
);

INVx2_ASAP7_75t_L g351 ( 
.A(n_284),
.Y(n_351)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_351),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_304),
.B(n_272),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_SL g411 ( 
.A(n_353),
.B(n_356),
.Y(n_411)
);

INVxp67_ASAP7_75t_L g355 ( 
.A(n_311),
.Y(n_355)
);

NAND2xp33_ASAP7_75t_SL g412 ( 
.A(n_355),
.B(n_277),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_332),
.B(n_273),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_276),
.B(n_228),
.Y(n_357)
);

CKINVDCx14_ASAP7_75t_R g389 ( 
.A(n_357),
.Y(n_389)
);

NOR2xp33_ASAP7_75t_L g358 ( 
.A(n_291),
.B(n_245),
.Y(n_358)
);

INVxp67_ASAP7_75t_L g377 ( 
.A(n_358),
.Y(n_377)
);

CKINVDCx20_ASAP7_75t_R g359 ( 
.A(n_312),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g387 ( 
.A(n_359),
.Y(n_387)
);

OAI21xp5_ASAP7_75t_L g360 ( 
.A1(n_332),
.A2(n_239),
.B(n_229),
.Y(n_360)
);

INVxp67_ASAP7_75t_L g388 ( 
.A(n_360),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_314),
.B(n_280),
.Y(n_362)
);

BUFx12f_ASAP7_75t_L g363 ( 
.A(n_303),
.Y(n_363)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_363),
.Y(n_390)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_290),
.Y(n_365)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_365),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_296),
.B(n_253),
.Y(n_366)
);

XNOR2xp5_ASAP7_75t_L g397 ( 
.A(n_366),
.B(n_372),
.Y(n_397)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_284),
.Y(n_367)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_367),
.Y(n_391)
);

NOR2xp33_ASAP7_75t_L g368 ( 
.A(n_330),
.B(n_261),
.Y(n_368)
);

INVxp67_ASAP7_75t_L g402 ( 
.A(n_368),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_SL g369 ( 
.A(n_305),
.B(n_331),
.Y(n_369)
);

NOR3xp33_ASAP7_75t_L g410 ( 
.A(n_369),
.B(n_371),
.C(n_374),
.Y(n_410)
);

INVx13_ASAP7_75t_L g370 ( 
.A(n_325),
.Y(n_370)
);

CKINVDCx20_ASAP7_75t_R g401 ( 
.A(n_370),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_SL g371 ( 
.A(n_275),
.B(n_249),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_275),
.B(n_225),
.Y(n_372)
);

INVx2_ASAP7_75t_L g373 ( 
.A(n_327),
.Y(n_373)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_373),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_SL g374 ( 
.A(n_313),
.B(n_227),
.Y(n_374)
);

INVx3_ASAP7_75t_L g375 ( 
.A(n_327),
.Y(n_375)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_375),
.Y(n_405)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_319),
.Y(n_376)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_376),
.Y(n_413)
);

AOI22xp5_ASAP7_75t_SL g378 ( 
.A1(n_339),
.A2(n_286),
.B1(n_309),
.B2(n_317),
.Y(n_378)
);

OAI21xp5_ASAP7_75t_SL g427 ( 
.A1(n_378),
.A2(n_381),
.B(n_412),
.Y(n_427)
);

INVxp67_ASAP7_75t_L g419 ( 
.A(n_379),
.Y(n_419)
);

OAI22xp5_ASAP7_75t_SL g380 ( 
.A1(n_362),
.A2(n_320),
.B1(n_315),
.B2(n_281),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_380),
.B(n_393),
.Y(n_418)
);

AOI22xp5_ASAP7_75t_SL g381 ( 
.A1(n_339),
.A2(n_286),
.B1(n_317),
.B2(n_308),
.Y(n_381)
);

MAJx2_ASAP7_75t_L g383 ( 
.A(n_335),
.B(n_297),
.C(n_328),
.Y(n_383)
);

MAJx2_ASAP7_75t_L g436 ( 
.A(n_383),
.B(n_361),
.C(n_370),
.Y(n_436)
);

OAI22xp5_ASAP7_75t_SL g393 ( 
.A1(n_372),
.A2(n_317),
.B1(n_321),
.B2(n_308),
.Y(n_393)
);

AND2x6_ASAP7_75t_L g396 ( 
.A(n_348),
.B(n_303),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_L g428 ( 
.A(n_396),
.B(n_356),
.Y(n_428)
);

AOI22xp33_ASAP7_75t_L g398 ( 
.A1(n_345),
.A2(n_324),
.B1(n_297),
.B2(n_293),
.Y(n_398)
);

OAI22xp5_ASAP7_75t_L g431 ( 
.A1(n_398),
.A2(n_350),
.B1(n_303),
.B2(n_337),
.Y(n_431)
);

MAJIxp5_ASAP7_75t_L g399 ( 
.A(n_349),
.B(n_325),
.C(n_313),
.Y(n_399)
);

MAJIxp5_ASAP7_75t_L g423 ( 
.A(n_399),
.B(n_355),
.C(n_342),
.Y(n_423)
);

OAI21xp5_ASAP7_75t_SL g403 ( 
.A1(n_339),
.A2(n_277),
.B(n_298),
.Y(n_403)
);

INVxp67_ASAP7_75t_L g420 ( 
.A(n_403),
.Y(n_420)
);

AO21x2_ASAP7_75t_L g407 ( 
.A1(n_366),
.A2(n_345),
.B(n_352),
.Y(n_407)
);

OAI22xp5_ASAP7_75t_L g430 ( 
.A1(n_407),
.A2(n_340),
.B1(n_364),
.B2(n_369),
.Y(n_430)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_353),
.Y(n_408)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_408),
.Y(n_415)
);

OAI21xp5_ASAP7_75t_L g416 ( 
.A1(n_388),
.A2(n_346),
.B(n_360),
.Y(n_416)
);

AOI21x1_ASAP7_75t_SL g470 ( 
.A1(n_416),
.A2(n_417),
.B(n_414),
.Y(n_470)
);

FAx1_ASAP7_75t_L g417 ( 
.A(n_393),
.B(n_352),
.CI(n_354),
.CON(n_417),
.SN(n_417)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_408),
.B(n_359),
.Y(n_421)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_421),
.Y(n_468)
);

OAI22x1_ASAP7_75t_SL g422 ( 
.A1(n_407),
.A2(n_364),
.B1(n_352),
.B2(n_371),
.Y(n_422)
);

AOI22xp5_ASAP7_75t_L g467 ( 
.A1(n_422),
.A2(n_430),
.B1(n_444),
.B2(n_390),
.Y(n_467)
);

MAJIxp5_ASAP7_75t_L g458 ( 
.A(n_423),
.B(n_436),
.C(n_439),
.Y(n_458)
);

INVxp67_ASAP7_75t_L g424 ( 
.A(n_399),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_424),
.B(n_434),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_397),
.B(n_344),
.Y(n_425)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_425),
.Y(n_479)
);

NOR2xp33_ASAP7_75t_SL g426 ( 
.A(n_387),
.B(n_377),
.Y(n_426)
);

NOR2xp33_ASAP7_75t_SL g466 ( 
.A(n_426),
.B(n_432),
.Y(n_466)
);

OAI22xp5_ASAP7_75t_L g482 ( 
.A1(n_428),
.A2(n_288),
.B1(n_310),
.B2(n_292),
.Y(n_482)
);

NOR2xp33_ASAP7_75t_L g429 ( 
.A(n_389),
.B(n_334),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_SL g454 ( 
.A(n_429),
.B(n_433),
.Y(n_454)
);

AOI22xp33_ASAP7_75t_L g462 ( 
.A1(n_431),
.A2(n_390),
.B1(n_409),
.B2(n_406),
.Y(n_462)
);

NOR2xp33_ASAP7_75t_SL g432 ( 
.A(n_377),
.B(n_365),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_SL g433 ( 
.A(n_404),
.B(n_376),
.Y(n_433)
);

CKINVDCx20_ASAP7_75t_R g434 ( 
.A(n_401),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_397),
.B(n_343),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_435),
.B(n_441),
.Y(n_471)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_386),
.Y(n_437)
);

INVx1_ASAP7_75t_SL g461 ( 
.A(n_437),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_SL g438 ( 
.A(n_402),
.B(n_336),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_SL g459 ( 
.A(n_438),
.B(n_448),
.Y(n_459)
);

XNOR2xp5_ASAP7_75t_L g439 ( 
.A(n_385),
.B(n_361),
.Y(n_439)
);

XNOR2xp5_ASAP7_75t_L g440 ( 
.A(n_385),
.B(n_375),
.Y(n_440)
);

MAJIxp5_ASAP7_75t_L g465 ( 
.A(n_440),
.B(n_445),
.C(n_447),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_411),
.B(n_373),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_384),
.B(n_367),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_442),
.B(n_443),
.Y(n_475)
);

CKINVDCx20_ASAP7_75t_R g443 ( 
.A(n_395),
.Y(n_443)
);

OAI22xp5_ASAP7_75t_L g444 ( 
.A1(n_407),
.A2(n_378),
.B1(n_381),
.B2(n_388),
.Y(n_444)
);

XNOR2xp5_ASAP7_75t_L g445 ( 
.A(n_395),
.B(n_351),
.Y(n_445)
);

CKINVDCx20_ASAP7_75t_R g446 ( 
.A(n_400),
.Y(n_446)
);

CKINVDCx20_ASAP7_75t_R g481 ( 
.A(n_446),
.Y(n_481)
);

MAJIxp5_ASAP7_75t_L g447 ( 
.A(n_400),
.B(n_287),
.C(n_324),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_SL g448 ( 
.A(n_402),
.B(n_287),
.Y(n_448)
);

NOR2xp33_ASAP7_75t_L g449 ( 
.A(n_413),
.B(n_409),
.Y(n_449)
);

INVxp33_ASAP7_75t_L g457 ( 
.A(n_449),
.Y(n_457)
);

MAJIxp5_ASAP7_75t_L g450 ( 
.A(n_403),
.B(n_370),
.C(n_292),
.Y(n_450)
);

MAJIxp5_ASAP7_75t_L g472 ( 
.A(n_450),
.B(n_440),
.C(n_424),
.Y(n_472)
);

OAI22xp5_ASAP7_75t_SL g451 ( 
.A1(n_418),
.A2(n_407),
.B1(n_379),
.B2(n_396),
.Y(n_451)
);

AOI22xp5_ASAP7_75t_L g496 ( 
.A1(n_451),
.A2(n_452),
.B1(n_460),
.B2(n_464),
.Y(n_496)
);

OAI22xp5_ASAP7_75t_SL g452 ( 
.A1(n_418),
.A2(n_407),
.B1(n_380),
.B2(n_410),
.Y(n_452)
);

INVxp67_ASAP7_75t_L g453 ( 
.A(n_450),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_453),
.B(n_469),
.Y(n_494)
);

NOR2xp33_ASAP7_75t_L g456 ( 
.A(n_426),
.B(n_392),
.Y(n_456)
);

NOR2xp33_ASAP7_75t_SL g491 ( 
.A(n_456),
.B(n_463),
.Y(n_491)
);

OAI22xp5_ASAP7_75t_SL g460 ( 
.A1(n_443),
.A2(n_419),
.B1(n_446),
.B2(n_415),
.Y(n_460)
);

OAI22xp5_ASAP7_75t_SL g488 ( 
.A1(n_462),
.A2(n_480),
.B1(n_420),
.B2(n_363),
.Y(n_488)
);

NOR2xp33_ASAP7_75t_L g463 ( 
.A(n_432),
.B(n_392),
.Y(n_463)
);

OAI22xp5_ASAP7_75t_SL g464 ( 
.A1(n_419),
.A2(n_383),
.B1(n_406),
.B2(n_414),
.Y(n_464)
);

OAI22xp5_ASAP7_75t_L g497 ( 
.A1(n_467),
.A2(n_473),
.B1(n_477),
.B2(n_422),
.Y(n_497)
);

INVxp67_ASAP7_75t_L g469 ( 
.A(n_447),
.Y(n_469)
);

OAI21xp5_ASAP7_75t_L g495 ( 
.A1(n_470),
.A2(n_427),
.B(n_417),
.Y(n_495)
);

MAJIxp5_ASAP7_75t_L g483 ( 
.A(n_472),
.B(n_436),
.C(n_442),
.Y(n_483)
);

AND2x6_ASAP7_75t_L g473 ( 
.A(n_417),
.B(n_278),
.Y(n_473)
);

NOR3xp33_ASAP7_75t_L g474 ( 
.A(n_421),
.B(n_405),
.C(n_394),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_SL g501 ( 
.A(n_474),
.B(n_363),
.Y(n_501)
);

XOR2xp5_ASAP7_75t_L g476 ( 
.A(n_439),
.B(n_405),
.Y(n_476)
);

XOR2xp5_ASAP7_75t_L g489 ( 
.A(n_476),
.B(n_478),
.Y(n_489)
);

AOI22xp5_ASAP7_75t_L g477 ( 
.A1(n_430),
.A2(n_394),
.B1(n_391),
.B2(n_382),
.Y(n_477)
);

XOR2xp5_ASAP7_75t_L g478 ( 
.A(n_423),
.B(n_391),
.Y(n_478)
);

OAI22xp5_ASAP7_75t_SL g480 ( 
.A1(n_415),
.A2(n_382),
.B1(n_338),
.B2(n_363),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_482),
.B(n_310),
.Y(n_503)
);

MAJIxp5_ASAP7_75t_L g520 ( 
.A(n_483),
.B(n_484),
.C(n_487),
.Y(n_520)
);

MAJIxp5_ASAP7_75t_L g484 ( 
.A(n_472),
.B(n_435),
.C(n_445),
.Y(n_484)
);

NAND2xp33_ASAP7_75t_SL g485 ( 
.A(n_455),
.B(n_416),
.Y(n_485)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_485),
.Y(n_517)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_466),
.Y(n_486)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_486),
.Y(n_518)
);

MAJIxp5_ASAP7_75t_L g487 ( 
.A(n_478),
.B(n_425),
.C(n_420),
.Y(n_487)
);

AND2x2_ASAP7_75t_L g534 ( 
.A(n_488),
.B(n_497),
.Y(n_534)
);

XNOR2xp5_ASAP7_75t_L g490 ( 
.A(n_458),
.B(n_444),
.Y(n_490)
);

XNOR2xp5_ASAP7_75t_L g512 ( 
.A(n_490),
.B(n_506),
.Y(n_512)
);

AOI21xp5_ASAP7_75t_SL g492 ( 
.A1(n_468),
.A2(n_427),
.B(n_417),
.Y(n_492)
);

OAI21xp5_ASAP7_75t_L g516 ( 
.A1(n_492),
.A2(n_495),
.B(n_470),
.Y(n_516)
);

NOR2xp33_ASAP7_75t_L g493 ( 
.A(n_466),
.B(n_434),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g531 ( 
.A(n_493),
.B(n_507),
.Y(n_531)
);

AND2x2_ASAP7_75t_L g498 ( 
.A(n_455),
.B(n_441),
.Y(n_498)
);

CKINVDCx14_ASAP7_75t_R g527 ( 
.A(n_498),
.Y(n_527)
);

MAJIxp5_ASAP7_75t_L g499 ( 
.A(n_458),
.B(n_437),
.C(n_283),
.Y(n_499)
);

MAJIxp5_ASAP7_75t_L g522 ( 
.A(n_499),
.B(n_502),
.C(n_504),
.Y(n_522)
);

BUFx3_ASAP7_75t_L g500 ( 
.A(n_467),
.Y(n_500)
);

INVx2_ASAP7_75t_L g524 ( 
.A(n_500),
.Y(n_524)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_501),
.Y(n_521)
);

MAJIxp5_ASAP7_75t_L g502 ( 
.A(n_465),
.B(n_283),
.C(n_278),
.Y(n_502)
);

OAI22xp5_ASAP7_75t_L g515 ( 
.A1(n_503),
.A2(n_461),
.B1(n_481),
.B2(n_453),
.Y(n_515)
);

MAJIxp5_ASAP7_75t_L g504 ( 
.A(n_465),
.B(n_289),
.C(n_300),
.Y(n_504)
);

MAJIxp5_ASAP7_75t_L g505 ( 
.A(n_476),
.B(n_295),
.C(n_300),
.Y(n_505)
);

MAJIxp5_ASAP7_75t_L g528 ( 
.A(n_505),
.B(n_508),
.C(n_480),
.Y(n_528)
);

XNOR2xp5_ASAP7_75t_L g506 ( 
.A(n_464),
.B(n_288),
.Y(n_506)
);

NOR2xp33_ASAP7_75t_L g507 ( 
.A(n_457),
.B(n_318),
.Y(n_507)
);

MAJIxp5_ASAP7_75t_L g508 ( 
.A(n_469),
.B(n_295),
.C(n_232),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_468),
.Y(n_509)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_509),
.Y(n_525)
);

AND2x2_ASAP7_75t_L g510 ( 
.A(n_451),
.B(n_293),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_510),
.B(n_452),
.Y(n_514)
);

BUFx3_ASAP7_75t_L g511 ( 
.A(n_500),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_L g538 ( 
.A(n_511),
.B(n_533),
.Y(n_538)
);

OAI22xp5_ASAP7_75t_SL g513 ( 
.A1(n_496),
.A2(n_481),
.B1(n_477),
.B2(n_475),
.Y(n_513)
);

AOI22xp5_ASAP7_75t_L g548 ( 
.A1(n_513),
.A2(n_510),
.B1(n_496),
.B2(n_506),
.Y(n_548)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_514),
.Y(n_539)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_515),
.Y(n_543)
);

OAI21xp5_ASAP7_75t_L g540 ( 
.A1(n_516),
.A2(n_492),
.B(n_495),
.Y(n_540)
);

XNOR2xp5_ASAP7_75t_L g519 ( 
.A(n_489),
.B(n_460),
.Y(n_519)
);

XNOR2xp5_ASAP7_75t_L g537 ( 
.A(n_519),
.B(n_528),
.Y(n_537)
);

XOR2xp5_ASAP7_75t_L g523 ( 
.A(n_490),
.B(n_471),
.Y(n_523)
);

XOR2xp5_ASAP7_75t_L g535 ( 
.A(n_523),
.B(n_526),
.Y(n_535)
);

XOR2xp5_ASAP7_75t_L g526 ( 
.A(n_489),
.B(n_471),
.Y(n_526)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_491),
.Y(n_529)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_529),
.Y(n_547)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_498),
.Y(n_530)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_530),
.Y(n_551)
);

XOR2xp5_ASAP7_75t_L g532 ( 
.A(n_484),
.B(n_479),
.Y(n_532)
);

XOR2xp5_ASAP7_75t_L g541 ( 
.A(n_532),
.B(n_487),
.Y(n_541)
);

NOR2xp33_ASAP7_75t_L g533 ( 
.A(n_494),
.B(n_454),
.Y(n_533)
);

MAJIxp5_ASAP7_75t_L g536 ( 
.A(n_522),
.B(n_499),
.C(n_504),
.Y(n_536)
);

NOR2xp33_ASAP7_75t_L g562 ( 
.A(n_536),
.B(n_545),
.Y(n_562)
);

OAI21xp5_ASAP7_75t_L g567 ( 
.A1(n_540),
.A2(n_552),
.B(n_259),
.Y(n_567)
);

XNOR2xp5_ASAP7_75t_L g569 ( 
.A(n_541),
.B(n_544),
.Y(n_569)
);

AO221x1_ASAP7_75t_L g542 ( 
.A1(n_518),
.A2(n_479),
.B1(n_459),
.B2(n_461),
.C(n_473),
.Y(n_542)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_542),
.Y(n_555)
);

XOR2xp5_ASAP7_75t_L g544 ( 
.A(n_512),
.B(n_519),
.Y(n_544)
);

FAx1_ASAP7_75t_SL g545 ( 
.A(n_516),
.B(n_475),
.CI(n_483),
.CON(n_545),
.SN(n_545)
);

MAJIxp5_ASAP7_75t_L g546 ( 
.A(n_522),
.B(n_502),
.C(n_505),
.Y(n_546)
);

OAI21xp5_ASAP7_75t_SL g558 ( 
.A1(n_546),
.A2(n_520),
.B(n_528),
.Y(n_558)
);

OAI22xp5_ASAP7_75t_SL g554 ( 
.A1(n_548),
.A2(n_550),
.B1(n_524),
.B2(n_511),
.Y(n_554)
);

NOR2xp33_ASAP7_75t_L g549 ( 
.A(n_532),
.B(n_508),
.Y(n_549)
);

CKINVDCx20_ASAP7_75t_R g563 ( 
.A(n_549),
.Y(n_563)
);

AOI22xp5_ASAP7_75t_L g550 ( 
.A1(n_534),
.A2(n_318),
.B1(n_231),
.B2(n_240),
.Y(n_550)
);

AOI21xp5_ASAP7_75t_L g552 ( 
.A1(n_517),
.A2(n_250),
.B(n_266),
.Y(n_552)
);

XOR2xp5_ASAP7_75t_L g553 ( 
.A(n_512),
.B(n_266),
.Y(n_553)
);

XOR2xp5_ASAP7_75t_L g556 ( 
.A(n_553),
.B(n_526),
.Y(n_556)
);

AOI22xp5_ASAP7_75t_L g572 ( 
.A1(n_554),
.A2(n_538),
.B1(n_553),
.B2(n_545),
.Y(n_572)
);

XOR2xp5_ASAP7_75t_L g575 ( 
.A(n_556),
.B(n_560),
.Y(n_575)
);

AOI21x1_ASAP7_75t_L g557 ( 
.A1(n_540),
.A2(n_521),
.B(n_534),
.Y(n_557)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_557),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_SL g580 ( 
.A(n_558),
.B(n_559),
.Y(n_580)
);

OAI21xp5_ASAP7_75t_SL g559 ( 
.A1(n_539),
.A2(n_520),
.B(n_527),
.Y(n_559)
);

XOR2xp5_ASAP7_75t_L g560 ( 
.A(n_544),
.B(n_523),
.Y(n_560)
);

XOR2xp5_ASAP7_75t_L g561 ( 
.A(n_535),
.B(n_534),
.Y(n_561)
);

NOR2xp33_ASAP7_75t_L g571 ( 
.A(n_561),
.B(n_564),
.Y(n_571)
);

XOR2xp5_ASAP7_75t_L g564 ( 
.A(n_535),
.B(n_514),
.Y(n_564)
);

AOI22xp5_ASAP7_75t_L g565 ( 
.A1(n_543),
.A2(n_513),
.B1(n_524),
.B2(n_525),
.Y(n_565)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_565),
.Y(n_581)
);

XOR2xp5_ASAP7_75t_L g566 ( 
.A(n_537),
.B(n_531),
.Y(n_566)
);

NOR2xp33_ASAP7_75t_L g576 ( 
.A(n_566),
.B(n_568),
.Y(n_576)
);

CKINVDCx16_ASAP7_75t_R g577 ( 
.A(n_567),
.Y(n_577)
);

AOI22xp5_ASAP7_75t_L g568 ( 
.A1(n_547),
.A2(n_274),
.B1(n_215),
.B2(n_220),
.Y(n_568)
);

OAI21xp5_ASAP7_75t_L g570 ( 
.A1(n_562),
.A2(n_551),
.B(n_545),
.Y(n_570)
);

AO21x1_ASAP7_75t_L g590 ( 
.A1(n_570),
.A2(n_573),
.B(n_567),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_L g583 ( 
.A(n_572),
.B(n_574),
.Y(n_583)
);

OAI21xp5_ASAP7_75t_L g573 ( 
.A1(n_555),
.A2(n_548),
.B(n_552),
.Y(n_573)
);

MAJIxp5_ASAP7_75t_L g574 ( 
.A(n_566),
.B(n_536),
.C(n_537),
.Y(n_574)
);

NOR2xp33_ASAP7_75t_L g579 ( 
.A(n_563),
.B(n_546),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g584 ( 
.A(n_579),
.B(n_569),
.Y(n_584)
);

NOR2xp33_ASAP7_75t_SL g582 ( 
.A(n_569),
.B(n_541),
.Y(n_582)
);

NOR2xp33_ASAP7_75t_L g587 ( 
.A(n_582),
.B(n_556),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_L g594 ( 
.A(n_584),
.B(n_585),
.Y(n_594)
);

MAJIxp5_ASAP7_75t_L g585 ( 
.A(n_574),
.B(n_560),
.C(n_561),
.Y(n_585)
);

INVxp67_ASAP7_75t_L g586 ( 
.A(n_580),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_L g598 ( 
.A(n_586),
.B(n_588),
.Y(n_598)
);

NOR2xp33_ASAP7_75t_SL g593 ( 
.A(n_587),
.B(n_592),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_L g588 ( 
.A(n_570),
.B(n_565),
.Y(n_588)
);

MAJIxp5_ASAP7_75t_L g589 ( 
.A(n_575),
.B(n_564),
.C(n_550),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_L g599 ( 
.A(n_589),
.B(n_591),
.Y(n_599)
);

XNOR2xp5_ASAP7_75t_L g596 ( 
.A(n_590),
.B(n_581),
.Y(n_596)
);

AOI22xp5_ASAP7_75t_L g591 ( 
.A1(n_578),
.A2(n_223),
.B1(n_250),
.B2(n_3),
.Y(n_591)
);

CKINVDCx20_ASAP7_75t_R g592 ( 
.A(n_572),
.Y(n_592)
);

AOI322xp5_ASAP7_75t_L g595 ( 
.A1(n_586),
.A2(n_578),
.A3(n_581),
.B1(n_577),
.B2(n_571),
.C1(n_576),
.C2(n_573),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_SL g601 ( 
.A(n_595),
.B(n_596),
.Y(n_601)
);

MAJIxp5_ASAP7_75t_L g597 ( 
.A(n_583),
.B(n_575),
.C(n_1),
.Y(n_597)
);

NOR2xp33_ASAP7_75t_L g603 ( 
.A(n_597),
.B(n_0),
.Y(n_603)
);

OAI21xp5_ASAP7_75t_SL g600 ( 
.A1(n_594),
.A2(n_585),
.B(n_590),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_L g605 ( 
.A(n_600),
.B(n_603),
.Y(n_605)
);

XOR2xp5_ASAP7_75t_L g602 ( 
.A(n_599),
.B(n_0),
.Y(n_602)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_602),
.Y(n_604)
);

A2O1A1Ixp33_ASAP7_75t_L g606 ( 
.A1(n_605),
.A2(n_598),
.B(n_601),
.C(n_593),
.Y(n_606)
);

NOR3xp33_ASAP7_75t_L g608 ( 
.A(n_606),
.B(n_607),
.C(n_0),
.Y(n_608)
);

AOI21xp5_ASAP7_75t_R g607 ( 
.A1(n_604),
.A2(n_595),
.B(n_1),
.Y(n_607)
);

BUFx24_ASAP7_75t_SL g609 ( 
.A(n_608),
.Y(n_609)
);

FAx1_ASAP7_75t_SL g610 ( 
.A(n_609),
.B(n_1),
.CI(n_2),
.CON(n_610),
.SN(n_610)
);

MAJx2_ASAP7_75t_L g611 ( 
.A(n_610),
.B(n_2),
.C(n_601),
.Y(n_611)
);


endmodule