module fake_jpeg_16363_n_380 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_380);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_380;

wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_4),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_2),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_7),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_1),
.B(n_5),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_3),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_2),
.Y(n_24)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_5),
.B(n_0),
.Y(n_31)
);

INVx1_ASAP7_75t_SL g32 ( 
.A(n_9),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_0),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_13),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_34),
.Y(n_37)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_37),
.Y(n_76)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_36),
.Y(n_38)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_38),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_14),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_39),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g40 ( 
.A(n_17),
.B(n_7),
.Y(n_40)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_40),
.B(n_24),
.Y(n_85)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_14),
.Y(n_41)
);

INVx5_ASAP7_75t_L g112 ( 
.A(n_41),
.Y(n_112)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_19),
.Y(n_42)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_42),
.Y(n_68)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_30),
.Y(n_43)
);

INVx8_ASAP7_75t_L g88 ( 
.A(n_43),
.Y(n_88)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_19),
.Y(n_44)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_44),
.Y(n_96)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_26),
.Y(n_45)
);

INVx11_ASAP7_75t_L g110 ( 
.A(n_45),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g46 ( 
.A1(n_26),
.A2(n_13),
.B1(n_1),
.B2(n_2),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_46),
.A2(n_33),
.B1(n_29),
.B2(n_28),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_14),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_47),
.Y(n_77)
);

OR2x2_ASAP7_75t_L g48 ( 
.A(n_16),
.B(n_7),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_48),
.B(n_57),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_14),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_49),
.Y(n_80)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_50),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_20),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_51),
.Y(n_86)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_30),
.Y(n_52)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_52),
.Y(n_83)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_30),
.Y(n_53)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_53),
.Y(n_90)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_26),
.Y(n_54)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_54),
.Y(n_97)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_34),
.Y(n_55)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_55),
.Y(n_95)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_30),
.Y(n_56)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_56),
.Y(n_100)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_36),
.Y(n_57)
);

INVx2_ASAP7_75t_SL g58 ( 
.A(n_30),
.Y(n_58)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_58),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_20),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_59),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_20),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_60),
.Y(n_102)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_20),
.Y(n_61)
);

BUFx2_ASAP7_75t_L g78 ( 
.A(n_61),
.Y(n_78)
);

BUFx5_ASAP7_75t_L g62 ( 
.A(n_30),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_62),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_17),
.B(n_7),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_63),
.B(n_64),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_31),
.B(n_8),
.Y(n_64)
);

BUFx4f_ASAP7_75t_L g65 ( 
.A(n_39),
.Y(n_65)
);

INVx5_ASAP7_75t_SL g123 ( 
.A(n_65),
.Y(n_123)
);

NAND3xp33_ASAP7_75t_L g66 ( 
.A(n_48),
.B(n_32),
.C(n_31),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_66),
.B(n_72),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_37),
.A2(n_26),
.B1(n_25),
.B2(n_19),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_69),
.A2(n_84),
.B1(n_111),
.B2(n_15),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_55),
.B(n_27),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_58),
.B(n_32),
.Y(n_73)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_73),
.Y(n_117)
);

BUFx3_ASAP7_75t_L g74 ( 
.A(n_41),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_74),
.B(n_92),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_50),
.B(n_27),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_75),
.B(n_79),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_46),
.B(n_16),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_45),
.A2(n_32),
.B1(n_25),
.B2(n_33),
.Y(n_81)
);

AOI21xp5_ASAP7_75t_L g141 ( 
.A1(n_81),
.A2(n_36),
.B(n_3),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_42),
.B(n_23),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_82),
.B(n_85),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_L g84 ( 
.A1(n_54),
.A2(n_25),
.B1(n_22),
.B2(n_23),
.Y(n_84)
);

INVx4_ASAP7_75t_SL g91 ( 
.A(n_62),
.Y(n_91)
);

INVx5_ASAP7_75t_SL g164 ( 
.A(n_91),
.Y(n_164)
);

INVx13_ASAP7_75t_L g92 ( 
.A(n_58),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_93),
.A2(n_99),
.B1(n_106),
.B2(n_6),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_56),
.B(n_24),
.Y(n_98)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_98),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_44),
.A2(n_28),
.B1(n_18),
.B2(n_33),
.Y(n_99)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_43),
.Y(n_103)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_103),
.Y(n_137)
);

OR2x2_ASAP7_75t_L g104 ( 
.A(n_38),
.B(n_29),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_104),
.B(n_96),
.Y(n_160)
);

NOR4xp25_ASAP7_75t_SL g105 ( 
.A(n_41),
.B(n_12),
.C(n_1),
.D(n_2),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g148 ( 
.A(n_105),
.B(n_13),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_52),
.A2(n_15),
.B1(n_29),
.B2(n_28),
.Y(n_106)
);

BUFx12f_ASAP7_75t_L g107 ( 
.A(n_61),
.Y(n_107)
);

INVx5_ASAP7_75t_L g140 ( 
.A(n_107),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_57),
.B(n_35),
.Y(n_108)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_108),
.Y(n_145)
);

BUFx12f_ASAP7_75t_L g109 ( 
.A(n_61),
.Y(n_109)
);

INVx5_ASAP7_75t_L g153 ( 
.A(n_109),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_L g111 ( 
.A1(n_53),
.A2(n_22),
.B1(n_21),
.B2(n_18),
.Y(n_111)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_60),
.Y(n_113)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_113),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_L g171 ( 
.A1(n_115),
.A2(n_141),
.B1(n_162),
.B2(n_143),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_110),
.A2(n_15),
.B1(n_21),
.B2(n_18),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_116),
.A2(n_133),
.B1(n_144),
.B2(n_162),
.Y(n_199)
);

BUFx2_ASAP7_75t_L g118 ( 
.A(n_83),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_118),
.Y(n_177)
);

O2A1O1Ixp33_ASAP7_75t_L g120 ( 
.A1(n_67),
.A2(n_35),
.B(n_21),
.C(n_49),
.Y(n_120)
);

CKINVDCx14_ASAP7_75t_R g207 ( 
.A(n_120),
.Y(n_207)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_71),
.Y(n_124)
);

INVx3_ASAP7_75t_L g206 ( 
.A(n_124),
.Y(n_206)
);

OAI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_97),
.A2(n_59),
.B1(n_51),
.B2(n_47),
.Y(n_125)
);

OAI22xp33_ASAP7_75t_SL g178 ( 
.A1(n_125),
.A2(n_126),
.B1(n_112),
.B2(n_86),
.Y(n_178)
);

OAI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_97),
.A2(n_22),
.B1(n_36),
.B2(n_4),
.Y(n_126)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_87),
.Y(n_127)
);

BUFx3_ASAP7_75t_L g173 ( 
.A(n_127),
.Y(n_173)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_100),
.Y(n_128)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_128),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_104),
.B(n_36),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_130),
.B(n_13),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_85),
.A2(n_66),
.B1(n_81),
.B2(n_84),
.Y(n_131)
);

OR2x2_ASAP7_75t_L g193 ( 
.A(n_131),
.B(n_156),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_70),
.B(n_10),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g185 ( 
.A(n_132),
.B(n_149),
.Y(n_185)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_110),
.A2(n_10),
.B1(n_3),
.B2(n_4),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_71),
.Y(n_134)
);

BUFx3_ASAP7_75t_L g210 ( 
.A(n_134),
.Y(n_210)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_77),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_135),
.Y(n_209)
);

BUFx3_ASAP7_75t_L g138 ( 
.A(n_114),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_138),
.B(n_142),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_SL g182 ( 
.A1(n_141),
.A2(n_148),
.B(n_159),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_76),
.Y(n_142)
);

OA22x2_ASAP7_75t_L g143 ( 
.A1(n_95),
.A2(n_22),
.B1(n_36),
.B2(n_0),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_143),
.A2(n_96),
.B1(n_112),
.B2(n_0),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_68),
.A2(n_9),
.B1(n_4),
.B2(n_6),
.Y(n_144)
);

CKINVDCx16_ASAP7_75t_R g146 ( 
.A(n_89),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_146),
.B(n_152),
.Y(n_166)
);

INVx3_ASAP7_75t_L g147 ( 
.A(n_90),
.Y(n_147)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_147),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_78),
.Y(n_149)
);

INVx4_ASAP7_75t_L g150 ( 
.A(n_88),
.Y(n_150)
);

INVxp67_ASAP7_75t_L g167 ( 
.A(n_150),
.Y(n_167)
);

INVx4_ASAP7_75t_L g151 ( 
.A(n_88),
.Y(n_151)
);

INVxp67_ASAP7_75t_L g184 ( 
.A(n_151),
.Y(n_184)
);

CKINVDCx14_ASAP7_75t_R g152 ( 
.A(n_111),
.Y(n_152)
);

CKINVDCx16_ASAP7_75t_R g154 ( 
.A(n_91),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_154),
.B(n_155),
.Y(n_189)
);

INVxp67_ASAP7_75t_L g155 ( 
.A(n_101),
.Y(n_155)
);

CKINVDCx16_ASAP7_75t_R g156 ( 
.A(n_65),
.Y(n_156)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_77),
.Y(n_157)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_157),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_78),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_SL g186 ( 
.A(n_158),
.B(n_74),
.Y(n_186)
);

AND2x2_ASAP7_75t_L g159 ( 
.A(n_92),
.B(n_6),
.Y(n_159)
);

AND2x2_ASAP7_75t_L g176 ( 
.A(n_160),
.B(n_6),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g161 ( 
.A(n_65),
.Y(n_161)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_161),
.Y(n_174)
);

HB1xp67_ASAP7_75t_L g163 ( 
.A(n_68),
.Y(n_163)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_163),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_80),
.Y(n_165)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_165),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_SL g214 ( 
.A1(n_169),
.A2(n_195),
.B(n_203),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_171),
.A2(n_180),
.B1(n_187),
.B2(n_190),
.Y(n_216)
);

OAI22xp33_ASAP7_75t_L g175 ( 
.A1(n_150),
.A2(n_80),
.B1(n_102),
.B2(n_94),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_175),
.A2(n_164),
.B1(n_165),
.B2(n_135),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_176),
.B(n_192),
.Y(n_247)
);

AOI22xp33_ASAP7_75t_L g238 ( 
.A1(n_178),
.A2(n_206),
.B1(n_177),
.B2(n_209),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_131),
.A2(n_86),
.B1(n_102),
.B2(n_94),
.Y(n_180)
);

AOI211xp5_ASAP7_75t_L g183 ( 
.A1(n_148),
.A2(n_109),
.B(n_107),
.C(n_114),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_183),
.A2(n_176),
.B1(n_195),
.B2(n_200),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_186),
.B(n_153),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_136),
.A2(n_107),
.B1(n_109),
.B2(n_11),
.Y(n_187)
);

FAx1_ASAP7_75t_SL g237 ( 
.A(n_188),
.B(n_192),
.CI(n_191),
.CON(n_237),
.SN(n_237)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_115),
.A2(n_8),
.B1(n_10),
.B2(n_11),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_130),
.B(n_122),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_191),
.B(n_194),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_117),
.B(n_11),
.C(n_12),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_148),
.B(n_159),
.Y(n_194)
);

AND2x2_ASAP7_75t_L g195 ( 
.A(n_143),
.B(n_139),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_159),
.B(n_120),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_196),
.B(n_200),
.Y(n_222)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_119),
.Y(n_197)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_197),
.Y(n_217)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_119),
.Y(n_198)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_198),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_143),
.B(n_129),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_147),
.Y(n_201)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_201),
.Y(n_230)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_128),
.Y(n_202)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_202),
.Y(n_233)
);

AOI21xp5_ASAP7_75t_L g203 ( 
.A1(n_155),
.A2(n_137),
.B(n_161),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_151),
.A2(n_157),
.B1(n_123),
.B2(n_145),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_204),
.A2(n_174),
.B1(n_170),
.B2(n_201),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_127),
.B(n_121),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_205),
.B(n_211),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_140),
.B(n_153),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_SL g270 ( 
.A(n_212),
.B(n_221),
.Y(n_270)
);

AOI21xp5_ASAP7_75t_L g213 ( 
.A1(n_182),
.A2(n_140),
.B(n_164),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_SL g266 ( 
.A1(n_213),
.A2(n_215),
.B(n_218),
.Y(n_266)
);

AND2x2_ASAP7_75t_SL g218 ( 
.A(n_196),
.B(n_123),
.Y(n_218)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_168),
.Y(n_219)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_219),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_185),
.B(n_118),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_208),
.B(n_138),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_224),
.B(n_225),
.Y(n_262)
);

CKINVDCx16_ASAP7_75t_R g225 ( 
.A(n_205),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_226),
.A2(n_235),
.B1(n_236),
.B2(n_181),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_211),
.B(n_188),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_228),
.B(n_231),
.Y(n_255)
);

AOI22xp33_ASAP7_75t_SL g229 ( 
.A1(n_207),
.A2(n_124),
.B1(n_134),
.B2(n_199),
.Y(n_229)
);

INVxp67_ASAP7_75t_L g259 ( 
.A(n_229),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_166),
.B(n_187),
.Y(n_231)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_168),
.Y(n_232)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_232),
.Y(n_253)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_202),
.Y(n_234)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_234),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_169),
.A2(n_194),
.B1(n_193),
.B2(n_180),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_237),
.B(n_242),
.Y(n_275)
);

CKINVDCx16_ASAP7_75t_R g282 ( 
.A(n_238),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_197),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_239),
.B(n_241),
.Y(n_269)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_198),
.Y(n_240)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_240),
.Y(n_261)
);

INVx1_ASAP7_75t_SL g241 ( 
.A(n_193),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_179),
.B(n_174),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_195),
.A2(n_182),
.B1(n_183),
.B2(n_190),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_L g256 ( 
.A1(n_243),
.A2(n_246),
.B1(n_251),
.B2(n_206),
.Y(n_256)
);

INVxp33_ASAP7_75t_L g244 ( 
.A(n_204),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_244),
.B(n_248),
.Y(n_274)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_172),
.Y(n_245)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_245),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_203),
.A2(n_170),
.B1(n_177),
.B2(n_184),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_SL g272 ( 
.A1(n_247),
.A2(n_218),
.B(n_220),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_179),
.B(n_189),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_176),
.B(n_167),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_249),
.B(n_243),
.Y(n_273)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_172),
.Y(n_250)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_250),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_167),
.A2(n_184),
.B1(n_209),
.B2(n_181),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_215),
.B(n_173),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_254),
.B(n_232),
.C(n_234),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_256),
.A2(n_282),
.B1(n_274),
.B2(n_259),
.Y(n_299)
);

INVx4_ASAP7_75t_L g258 ( 
.A(n_230),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_258),
.B(n_276),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_SL g300 ( 
.A1(n_260),
.A2(n_272),
.B(n_273),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_235),
.A2(n_241),
.B1(n_222),
.B2(n_216),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_263),
.A2(n_281),
.B1(n_283),
.B2(n_273),
.Y(n_296)
);

OAI21xp5_ASAP7_75t_L g264 ( 
.A1(n_213),
.A2(n_173),
.B(n_175),
.Y(n_264)
);

OAI21xp5_ASAP7_75t_L g311 ( 
.A1(n_264),
.A2(n_265),
.B(n_271),
.Y(n_311)
);

OAI21xp5_ASAP7_75t_L g265 ( 
.A1(n_222),
.A2(n_210),
.B(n_231),
.Y(n_265)
);

OAI21xp5_ASAP7_75t_L g271 ( 
.A1(n_227),
.A2(n_210),
.B(n_249),
.Y(n_271)
);

OAI32xp33_ASAP7_75t_L g276 ( 
.A1(n_220),
.A2(n_214),
.A3(n_228),
.B1(n_227),
.B2(n_216),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_248),
.B(n_242),
.Y(n_277)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_277),
.Y(n_293)
);

NAND2xp33_ASAP7_75t_SL g278 ( 
.A(n_218),
.B(n_214),
.Y(n_278)
);

AO21x1_ASAP7_75t_L g294 ( 
.A1(n_278),
.A2(n_266),
.B(n_284),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_221),
.B(n_225),
.Y(n_279)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_279),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_218),
.B(n_246),
.Y(n_280)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_280),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_226),
.A2(n_247),
.B1(n_237),
.B2(n_236),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_237),
.A2(n_212),
.B1(n_230),
.B2(n_239),
.Y(n_283)
);

OAI21xp5_ASAP7_75t_SL g284 ( 
.A1(n_251),
.A2(n_217),
.B(n_240),
.Y(n_284)
);

AOI21xp5_ASAP7_75t_SL g286 ( 
.A1(n_284),
.A2(n_223),
.B(n_233),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_283),
.B(n_217),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_285),
.B(n_289),
.C(n_292),
.Y(n_324)
);

OAI21xp5_ASAP7_75t_SL g313 ( 
.A1(n_286),
.A2(n_294),
.B(n_270),
.Y(n_313)
);

FAx1_ASAP7_75t_SL g287 ( 
.A(n_275),
.B(n_223),
.CI(n_233),
.CON(n_287),
.SN(n_287)
);

NOR2xp33_ASAP7_75t_SL g319 ( 
.A(n_287),
.B(n_290),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_252),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_288),
.B(n_296),
.Y(n_317)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_266),
.B(n_245),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_SL g290 ( 
.A(n_277),
.B(n_219),
.Y(n_290)
);

XOR2xp5_ASAP7_75t_L g327 ( 
.A(n_291),
.B(n_258),
.Y(n_327)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_254),
.B(n_250),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_280),
.A2(n_260),
.B1(n_263),
.B2(n_281),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_L g316 ( 
.A1(n_298),
.A2(n_299),
.B1(n_301),
.B2(n_309),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_282),
.A2(n_264),
.B1(n_276),
.B2(n_275),
.Y(n_301)
);

INVxp67_ASAP7_75t_L g302 ( 
.A(n_256),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_SL g321 ( 
.A(n_302),
.B(n_268),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_252),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_303),
.B(n_306),
.Y(n_332)
);

XNOR2xp5_ASAP7_75t_L g304 ( 
.A(n_272),
.B(n_271),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_304),
.B(n_305),
.C(n_307),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_255),
.B(n_278),
.C(n_265),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_253),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_255),
.B(n_279),
.C(n_262),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_262),
.B(n_269),
.C(n_270),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_308),
.B(n_305),
.C(n_292),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_SL g309 ( 
.A1(n_274),
.A2(n_269),
.B1(n_267),
.B2(n_261),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_261),
.A2(n_267),
.B1(n_258),
.B2(n_257),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g329 ( 
.A1(n_312),
.A2(n_310),
.B1(n_291),
.B2(n_289),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_SL g335 ( 
.A(n_313),
.B(n_333),
.Y(n_335)
);

INVxp67_ASAP7_75t_L g314 ( 
.A(n_312),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_314),
.B(n_318),
.Y(n_346)
);

OAI21xp5_ASAP7_75t_SL g315 ( 
.A1(n_286),
.A2(n_297),
.B(n_302),
.Y(n_315)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_315),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_293),
.Y(n_318)
);

AOI21xp5_ASAP7_75t_L g320 ( 
.A1(n_311),
.A2(n_253),
.B(n_257),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_SL g336 ( 
.A1(n_320),
.A2(n_329),
.B1(n_322),
.B2(n_321),
.Y(n_336)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_321),
.Y(n_339)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_309),
.Y(n_322)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_322),
.Y(n_348)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_295),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_323),
.B(n_331),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_326),
.B(n_327),
.C(n_324),
.Y(n_343)
);

NOR3xp33_ASAP7_75t_L g328 ( 
.A(n_308),
.B(n_268),
.C(n_307),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_328),
.B(n_287),
.Y(n_334)
);

XOR2xp5_ASAP7_75t_L g330 ( 
.A(n_304),
.B(n_300),
.Y(n_330)
);

XOR2xp5_ASAP7_75t_L g344 ( 
.A(n_330),
.B(n_324),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_287),
.B(n_285),
.Y(n_331)
);

OAI21xp5_ASAP7_75t_L g333 ( 
.A1(n_311),
.A2(n_294),
.B(n_300),
.Y(n_333)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_334),
.Y(n_353)
);

XNOR2xp5_ASAP7_75t_SL g357 ( 
.A(n_336),
.B(n_315),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_319),
.B(n_332),
.Y(n_337)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_337),
.Y(n_358)
);

XNOR2xp5_ASAP7_75t_L g340 ( 
.A(n_327),
.B(n_301),
.Y(n_340)
);

XOR2xp5_ASAP7_75t_L g351 ( 
.A(n_340),
.B(n_344),
.Y(n_351)
);

OAI22xp5_ASAP7_75t_SL g341 ( 
.A1(n_314),
.A2(n_299),
.B1(n_298),
.B2(n_296),
.Y(n_341)
);

AOI22xp5_ASAP7_75t_L g354 ( 
.A1(n_341),
.A2(n_349),
.B1(n_316),
.B2(n_331),
.Y(n_354)
);

BUFx24_ASAP7_75t_SL g342 ( 
.A(n_318),
.Y(n_342)
);

OAI21xp5_ASAP7_75t_L g361 ( 
.A1(n_342),
.A2(n_350),
.B(n_347),
.Y(n_361)
);

MAJIxp5_ASAP7_75t_L g355 ( 
.A(n_343),
.B(n_345),
.C(n_329),
.Y(n_355)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_326),
.B(n_325),
.C(n_330),
.Y(n_345)
);

HB1xp67_ASAP7_75t_L g349 ( 
.A(n_323),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_L g350 ( 
.A(n_319),
.B(n_317),
.Y(n_350)
);

XOR2xp5_ASAP7_75t_L g352 ( 
.A(n_344),
.B(n_325),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g362 ( 
.A(n_352),
.B(n_355),
.C(n_356),
.Y(n_362)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_354),
.Y(n_365)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_343),
.B(n_320),
.C(n_333),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_SL g367 ( 
.A(n_357),
.B(n_359),
.Y(n_367)
);

XOR2xp5_ASAP7_75t_L g359 ( 
.A(n_345),
.B(n_313),
.Y(n_359)
);

MAJIxp5_ASAP7_75t_L g360 ( 
.A(n_340),
.B(n_316),
.C(n_336),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_360),
.B(n_361),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_358),
.B(n_339),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_364),
.B(n_366),
.Y(n_371)
);

HB1xp67_ASAP7_75t_L g366 ( 
.A(n_360),
.Y(n_366)
);

AOI22xp5_ASAP7_75t_L g368 ( 
.A1(n_365),
.A2(n_346),
.B1(n_348),
.B2(n_338),
.Y(n_368)
);

OAI22xp5_ASAP7_75t_SL g373 ( 
.A1(n_368),
.A2(n_369),
.B1(n_335),
.B2(n_371),
.Y(n_373)
);

AOI22xp5_ASAP7_75t_L g369 ( 
.A1(n_367),
.A2(n_356),
.B1(n_357),
.B2(n_353),
.Y(n_369)
);

OAI22xp5_ASAP7_75t_SL g370 ( 
.A1(n_363),
.A2(n_335),
.B1(n_341),
.B2(n_355),
.Y(n_370)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_370),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_373),
.B(n_369),
.Y(n_374)
);

AOI21x1_ASAP7_75t_L g376 ( 
.A1(n_374),
.A2(n_375),
.B(n_373),
.Y(n_376)
);

AND2x2_ASAP7_75t_SL g375 ( 
.A(n_372),
.B(n_366),
.Y(n_375)
);

MAJIxp5_ASAP7_75t_L g377 ( 
.A(n_376),
.B(n_362),
.C(n_359),
.Y(n_377)
);

XOR2xp5_ASAP7_75t_L g378 ( 
.A(n_377),
.B(n_352),
.Y(n_378)
);

MAJIxp5_ASAP7_75t_L g379 ( 
.A(n_378),
.B(n_351),
.C(n_368),
.Y(n_379)
);

XNOR2xp5_ASAP7_75t_L g380 ( 
.A(n_379),
.B(n_351),
.Y(n_380)
);


endmodule