module fake_jpeg_8668_n_59 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_59);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_59;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_55;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_31;
wire n_25;
wire n_56;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;

CKINVDCx20_ASAP7_75t_R g8 ( 
.A(n_6),
.Y(n_8)
);

BUFx4f_ASAP7_75t_L g9 ( 
.A(n_2),
.Y(n_9)
);

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_2),
.Y(n_10)
);

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_5),
.Y(n_11)
);

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_3),
.Y(n_12)
);

INVx8_ASAP7_75t_L g13 ( 
.A(n_1),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_3),
.Y(n_14)
);

INVx2_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_5),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_SL g17 ( 
.A(n_10),
.B(n_0),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_17),
.B(n_21),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_10),
.B(n_0),
.Y(n_18)
);

CKINVDCx14_ASAP7_75t_R g27 ( 
.A(n_18),
.Y(n_27)
);

INVx4_ASAP7_75t_SL g19 ( 
.A(n_12),
.Y(n_19)
);

INVx11_ASAP7_75t_L g28 ( 
.A(n_19),
.Y(n_28)
);

INVx8_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

AOI22xp33_ASAP7_75t_SL g26 ( 
.A1(n_20),
.A2(n_22),
.B1(n_15),
.B2(n_13),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_SL g21 ( 
.A(n_11),
.B(n_0),
.Y(n_21)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

BUFx2_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_23),
.Y(n_25)
);

INVxp67_ASAP7_75t_L g35 ( 
.A(n_26),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_17),
.B(n_15),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_29),
.B(n_21),
.Y(n_33)
);

AOI22xp33_ASAP7_75t_SL g30 ( 
.A1(n_20),
.A2(n_13),
.B1(n_22),
.B2(n_19),
.Y(n_30)
);

AOI22xp33_ASAP7_75t_SL g36 ( 
.A1(n_30),
.A2(n_23),
.B1(n_1),
.B2(n_7),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_SL g31 ( 
.A1(n_20),
.A2(n_11),
.B1(n_16),
.B2(n_14),
.Y(n_31)
);

AOI22xp5_ASAP7_75t_L g34 ( 
.A1(n_31),
.A2(n_32),
.B1(n_12),
.B2(n_23),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_L g32 ( 
.A1(n_19),
.A2(n_14),
.B1(n_16),
.B2(n_8),
.Y(n_32)
);

XNOR2xp5_ASAP7_75t_L g43 ( 
.A(n_33),
.B(n_34),
.Y(n_43)
);

OAI21xp5_ASAP7_75t_L g45 ( 
.A1(n_36),
.A2(n_39),
.B(n_24),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_24),
.B(n_29),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_SL g46 ( 
.A(n_37),
.B(n_38),
.Y(n_46)
);

OR2x2_ASAP7_75t_L g38 ( 
.A(n_28),
.B(n_32),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g39 ( 
.A1(n_31),
.A2(n_1),
.B1(n_4),
.B2(n_7),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

HB1xp67_ASAP7_75t_L g44 ( 
.A(n_40),
.Y(n_44)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_34),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_41),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_38),
.Y(n_42)
);

OAI21xp5_ASAP7_75t_L g47 ( 
.A1(n_42),
.A2(n_45),
.B(n_35),
.Y(n_47)
);

XOR2xp5_ASAP7_75t_L g51 ( 
.A(n_47),
.B(n_48),
.Y(n_51)
);

XNOR2xp5_ASAP7_75t_L g48 ( 
.A(n_43),
.B(n_39),
.Y(n_48)
);

MAJIxp5_ASAP7_75t_L g50 ( 
.A(n_43),
.B(n_46),
.C(n_45),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_50),
.B(n_35),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_52),
.B(n_53),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_49),
.A2(n_27),
.B1(n_25),
.B2(n_44),
.Y(n_53)
);

NAND3xp33_ASAP7_75t_L g55 ( 
.A(n_51),
.B(n_50),
.C(n_27),
.Y(n_55)
);

MAJIxp5_ASAP7_75t_L g56 ( 
.A(n_55),
.B(n_51),
.C(n_54),
.Y(n_56)
);

NAND2x1_ASAP7_75t_L g57 ( 
.A(n_56),
.B(n_4),
.Y(n_57)
);

NAND3xp33_ASAP7_75t_L g58 ( 
.A(n_57),
.B(n_25),
.C(n_7),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_58),
.B(n_57),
.Y(n_59)
);


endmodule