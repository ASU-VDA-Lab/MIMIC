module real_aes_8358_n_104 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_104);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_104;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_766;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_571;
wire n_376;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_537;
wire n_320;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_774;
wire n_106;
wire n_559;
wire n_466;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_755;
wire n_656;
wire n_178;
wire n_409;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_449;
wire n_182;
wire n_363;
wire n_417;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_527;
wire n_434;
wire n_505;
wire n_502;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_733;
wire n_552;
wire n_402;
wire n_602;
wire n_617;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_768;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_756;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_481;
wire n_148;
wire n_498;
wire n_765;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_753;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_456;
wire n_156;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_762;
wire n_212;
wire n_210;
wire n_325;
wire n_575;
wire n_479;
wire n_338;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_729;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g499 ( .A1(n_0), .A2(n_181), .B(n_500), .C(n_503), .Y(n_499) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_1), .B(n_494), .Y(n_505) );
NAND3xp33_ASAP7_75t_SL g111 ( .A(n_2), .B(n_112), .C(n_113), .Y(n_111) );
INVx1_ASAP7_75t_L g451 ( .A(n_2), .Y(n_451) );
INVx1_ASAP7_75t_L g230 ( .A(n_3), .Y(n_230) );
OAI211xp5_ASAP7_75t_L g122 ( .A1(n_4), .A2(n_123), .B(n_453), .C(n_456), .Y(n_122) );
OAI211xp5_ASAP7_75t_L g453 ( .A1(n_4), .A2(n_125), .B(n_444), .C(n_454), .Y(n_453) );
NAND2xp5_ASAP7_75t_SL g528 ( .A(n_5), .B(n_169), .Y(n_528) );
AOI21xp5_ASAP7_75t_L g547 ( .A1(n_6), .A2(n_478), .B(n_548), .Y(n_547) );
OAI22xp5_ASAP7_75t_SL g440 ( .A1(n_7), .A2(n_11), .B1(n_441), .B2(n_442), .Y(n_440) );
CKINVDCx20_ASAP7_75t_R g441 ( .A(n_7), .Y(n_441) );
AO21x2_ASAP7_75t_L g556 ( .A1(n_8), .A2(n_186), .B(n_557), .Y(n_556) );
AOI22xp33_ASAP7_75t_L g180 ( .A1(n_9), .A2(n_39), .B1(n_142), .B2(n_154), .Y(n_180) );
NAND2xp5_ASAP7_75t_L g219 ( .A(n_10), .B(n_186), .Y(n_219) );
CKINVDCx20_ASAP7_75t_R g442 ( .A(n_11), .Y(n_442) );
AOI22xp5_ASAP7_75t_L g461 ( .A1(n_11), .A2(n_127), .B1(n_442), .B2(n_443), .Y(n_461) );
AND2x6_ASAP7_75t_L g157 ( .A(n_12), .B(n_158), .Y(n_157) );
A2O1A1Ixp33_ASAP7_75t_L g569 ( .A1(n_13), .A2(n_157), .B(n_481), .C(n_570), .Y(n_569) );
AOI22xp33_ASAP7_75t_L g104 ( .A1(n_14), .A2(n_105), .B1(n_116), .B2(n_773), .Y(n_104) );
NAND2xp5_ASAP7_75t_L g109 ( .A(n_15), .B(n_110), .Y(n_109) );
NOR2xp33_ASAP7_75t_L g452 ( .A(n_15), .B(n_40), .Y(n_452) );
INVx1_ASAP7_75t_L g138 ( .A(n_16), .Y(n_138) );
NAND2xp5_ASAP7_75t_L g145 ( .A(n_17), .B(n_146), .Y(n_145) );
INVx1_ASAP7_75t_L g224 ( .A(n_18), .Y(n_224) );
NAND2xp5_ASAP7_75t_SL g562 ( .A(n_19), .B(n_169), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g202 ( .A(n_20), .B(n_184), .Y(n_202) );
AO32x2_ASAP7_75t_L g178 ( .A1(n_21), .A2(n_179), .A3(n_183), .B1(n_185), .B2(n_186), .Y(n_178) );
OAI22xp5_ASAP7_75t_L g763 ( .A1(n_22), .A2(n_58), .B1(n_764), .B2(n_765), .Y(n_763) );
CKINVDCx20_ASAP7_75t_R g765 ( .A(n_22), .Y(n_765) );
NAND2xp5_ASAP7_75t_SL g152 ( .A(n_23), .B(n_142), .Y(n_152) );
NAND2xp5_ASAP7_75t_L g232 ( .A(n_24), .B(n_184), .Y(n_232) );
AOI22xp33_ASAP7_75t_L g182 ( .A1(n_25), .A2(n_56), .B1(n_142), .B2(n_154), .Y(n_182) );
AOI22xp33_ASAP7_75t_SL g195 ( .A1(n_26), .A2(n_83), .B1(n_142), .B2(n_146), .Y(n_195) );
NAND2xp5_ASAP7_75t_SL g172 ( .A(n_27), .B(n_142), .Y(n_172) );
A2O1A1Ixp33_ASAP7_75t_L g480 ( .A1(n_28), .A2(n_185), .B(n_481), .C(n_483), .Y(n_480) );
A2O1A1Ixp33_ASAP7_75t_L g559 ( .A1(n_29), .A2(n_185), .B(n_481), .C(n_560), .Y(n_559) );
BUFx6f_ASAP7_75t_L g150 ( .A(n_30), .Y(n_150) );
NAND2xp5_ASAP7_75t_L g244 ( .A(n_31), .B(n_134), .Y(n_244) );
AOI21xp5_ASAP7_75t_L g495 ( .A1(n_32), .A2(n_478), .B(n_496), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g176 ( .A(n_33), .B(n_134), .Y(n_176) );
INVx2_ASAP7_75t_L g144 ( .A(n_34), .Y(n_144) );
A2O1A1Ixp33_ASAP7_75t_L g511 ( .A1(n_35), .A2(n_512), .B(n_513), .C(n_517), .Y(n_511) );
NAND2xp5_ASAP7_75t_SL g239 ( .A(n_36), .B(n_142), .Y(n_239) );
NAND2xp5_ASAP7_75t_L g159 ( .A(n_37), .B(n_134), .Y(n_159) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_38), .B(n_149), .Y(n_561) );
INVx1_ASAP7_75t_L g110 ( .A(n_40), .Y(n_110) );
NAND2xp5_ASAP7_75t_L g476 ( .A(n_41), .B(n_477), .Y(n_476) );
CKINVDCx20_ASAP7_75t_R g574 ( .A(n_42), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g541 ( .A(n_43), .B(n_169), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g558 ( .A(n_44), .B(n_478), .Y(n_558) );
A2O1A1Ixp33_ASAP7_75t_L g538 ( .A1(n_45), .A2(n_512), .B(n_517), .C(n_539), .Y(n_538) );
AOI22xp5_ASAP7_75t_L g760 ( .A1(n_46), .A2(n_761), .B1(n_762), .B2(n_763), .Y(n_760) );
CKINVDCx20_ASAP7_75t_R g761 ( .A(n_46), .Y(n_761) );
NAND2xp5_ASAP7_75t_SL g212 ( .A(n_47), .B(n_142), .Y(n_212) );
INVx1_ASAP7_75t_L g501 ( .A(n_48), .Y(n_501) );
AOI22xp33_ASAP7_75t_L g193 ( .A1(n_49), .A2(n_93), .B1(n_154), .B2(n_194), .Y(n_193) );
INVx1_ASAP7_75t_L g540 ( .A(n_50), .Y(n_540) );
NAND2xp5_ASAP7_75t_SL g215 ( .A(n_51), .B(n_142), .Y(n_215) );
NAND2xp5_ASAP7_75t_L g226 ( .A(n_52), .B(n_142), .Y(n_226) );
NAND2xp5_ASAP7_75t_L g456 ( .A(n_53), .B(n_447), .Y(n_456) );
NAND2xp5_ASAP7_75t_L g537 ( .A(n_54), .B(n_478), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g216 ( .A(n_55), .B(n_217), .Y(n_216) );
AOI22xp33_ASAP7_75t_SL g206 ( .A1(n_57), .A2(n_62), .B1(n_142), .B2(n_146), .Y(n_206) );
CKINVDCx20_ASAP7_75t_R g764 ( .A(n_58), .Y(n_764) );
CKINVDCx20_ASAP7_75t_R g490 ( .A(n_59), .Y(n_490) );
NAND2xp5_ASAP7_75t_SL g141 ( .A(n_60), .B(n_142), .Y(n_141) );
NAND2xp5_ASAP7_75t_SL g243 ( .A(n_61), .B(n_142), .Y(n_243) );
INVx1_ASAP7_75t_L g158 ( .A(n_63), .Y(n_158) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_64), .B(n_478), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_65), .B(n_494), .Y(n_553) );
A2O1A1Ixp33_ASAP7_75t_L g550 ( .A1(n_66), .A2(n_217), .B(n_227), .C(n_551), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g231 ( .A(n_67), .B(n_142), .Y(n_231) );
INVx1_ASAP7_75t_L g137 ( .A(n_68), .Y(n_137) );
CKINVDCx20_ASAP7_75t_R g121 ( .A(n_69), .Y(n_121) );
NAND2xp5_ASAP7_75t_SL g515 ( .A(n_70), .B(n_169), .Y(n_515) );
AO32x2_ASAP7_75t_L g191 ( .A1(n_71), .A2(n_185), .A3(n_186), .B1(n_192), .B2(n_196), .Y(n_191) );
NAND2xp5_ASAP7_75t_L g571 ( .A(n_72), .B(n_170), .Y(n_571) );
INVx1_ASAP7_75t_L g242 ( .A(n_73), .Y(n_242) );
INVx1_ASAP7_75t_L g167 ( .A(n_74), .Y(n_167) );
CKINVDCx16_ASAP7_75t_R g497 ( .A(n_75), .Y(n_497) );
NAND2xp5_ASAP7_75t_L g484 ( .A(n_76), .B(n_485), .Y(n_484) );
NOR2xp33_ASAP7_75t_L g125 ( .A(n_77), .B(n_126), .Y(n_125) );
CKINVDCx20_ASAP7_75t_R g445 ( .A(n_77), .Y(n_445) );
A2O1A1Ixp33_ASAP7_75t_L g525 ( .A1(n_78), .A2(n_481), .B(n_517), .C(n_526), .Y(n_525) );
NAND2xp5_ASAP7_75t_SL g168 ( .A(n_79), .B(n_146), .Y(n_168) );
CKINVDCx16_ASAP7_75t_R g549 ( .A(n_80), .Y(n_549) );
INVx1_ASAP7_75t_L g115 ( .A(n_81), .Y(n_115) );
NAND2xp5_ASAP7_75t_SL g486 ( .A(n_82), .B(n_487), .Y(n_486) );
NAND2xp5_ASAP7_75t_L g153 ( .A(n_84), .B(n_154), .Y(n_153) );
CKINVDCx20_ASAP7_75t_R g519 ( .A(n_85), .Y(n_519) );
NAND2xp5_ASAP7_75t_SL g173 ( .A(n_86), .B(n_146), .Y(n_173) );
AOI222xp33_ASAP7_75t_L g458 ( .A1(n_87), .A2(n_459), .B1(n_759), .B2(n_760), .C1(n_766), .C2(n_768), .Y(n_458) );
INVx2_ASAP7_75t_L g135 ( .A(n_88), .Y(n_135) );
CKINVDCx20_ASAP7_75t_R g532 ( .A(n_89), .Y(n_532) );
NAND2xp5_ASAP7_75t_SL g572 ( .A(n_90), .B(n_156), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g213 ( .A(n_91), .B(n_146), .Y(n_213) );
INVx2_ASAP7_75t_L g112 ( .A(n_92), .Y(n_112) );
OR2x2_ASAP7_75t_L g448 ( .A(n_92), .B(n_449), .Y(n_448) );
OR2x2_ASAP7_75t_L g464 ( .A(n_92), .B(n_450), .Y(n_464) );
AOI22xp33_ASAP7_75t_L g205 ( .A1(n_94), .A2(n_103), .B1(n_146), .B2(n_147), .Y(n_205) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_95), .B(n_478), .Y(n_510) );
INVx1_ASAP7_75t_L g514 ( .A(n_96), .Y(n_514) );
INVxp67_ASAP7_75t_L g552 ( .A(n_97), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g240 ( .A(n_98), .B(n_146), .Y(n_240) );
NAND2xp5_ASAP7_75t_L g114 ( .A(n_99), .B(n_115), .Y(n_114) );
INVx1_ASAP7_75t_L g527 ( .A(n_100), .Y(n_527) );
INVx1_ASAP7_75t_L g567 ( .A(n_101), .Y(n_567) );
AND2x2_ASAP7_75t_L g542 ( .A(n_102), .B(n_134), .Y(n_542) );
INVx1_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
CKINVDCx12_ASAP7_75t_R g107 ( .A(n_108), .Y(n_107) );
INVx1_ASAP7_75t_SL g774 ( .A(n_108), .Y(n_774) );
OR2x2_ASAP7_75t_L g108 ( .A(n_109), .B(n_111), .Y(n_108) );
OR2x2_ASAP7_75t_L g758 ( .A(n_112), .B(n_450), .Y(n_758) );
NOR2x2_ASAP7_75t_L g770 ( .A(n_112), .B(n_449), .Y(n_770) );
INVx1_ASAP7_75t_SL g113 ( .A(n_114), .Y(n_113) );
OA21x2_ASAP7_75t_L g116 ( .A1(n_117), .A2(n_122), .B(n_457), .Y(n_116) );
BUFx2_ASAP7_75t_SL g117 ( .A(n_118), .Y(n_117) );
CKINVDCx20_ASAP7_75t_R g118 ( .A(n_119), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
INVx1_ASAP7_75t_SL g772 ( .A(n_120), .Y(n_772) );
INVx2_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
INVx1_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
NOR3xp33_ASAP7_75t_L g124 ( .A(n_125), .B(n_444), .C(n_447), .Y(n_124) );
INVx1_ASAP7_75t_L g446 ( .A(n_126), .Y(n_446) );
OAI22xp5_ASAP7_75t_SL g126 ( .A1(n_127), .A2(n_439), .B1(n_440), .B2(n_443), .Y(n_126) );
INVx1_ASAP7_75t_L g443 ( .A(n_127), .Y(n_443) );
OR2x2_ASAP7_75t_L g127 ( .A(n_128), .B(n_361), .Y(n_127) );
NAND5xp2_ASAP7_75t_L g128 ( .A(n_129), .B(n_280), .C(n_295), .D(n_321), .E(n_343), .Y(n_128) );
NOR2xp33_ASAP7_75t_SL g129 ( .A(n_130), .B(n_260), .Y(n_129) );
OAI221xp5_ASAP7_75t_L g130 ( .A1(n_131), .A2(n_197), .B1(n_233), .B2(n_249), .C(n_250), .Y(n_130) );
NOR2xp33_ASAP7_75t_SL g131 ( .A(n_132), .B(n_187), .Y(n_131) );
NAND2xp5_ASAP7_75t_L g309 ( .A(n_132), .B(n_310), .Y(n_309) );
INVx1_ASAP7_75t_SL g437 ( .A(n_132), .Y(n_437) );
AND2x2_ASAP7_75t_L g132 ( .A(n_133), .B(n_160), .Y(n_132) );
INVx1_ASAP7_75t_L g277 ( .A(n_133), .Y(n_277) );
AND2x2_ASAP7_75t_L g279 ( .A(n_133), .B(n_178), .Y(n_279) );
AND2x2_ASAP7_75t_L g289 ( .A(n_133), .B(n_177), .Y(n_289) );
HB1xp67_ASAP7_75t_L g307 ( .A(n_133), .Y(n_307) );
INVx1_ASAP7_75t_L g317 ( .A(n_133), .Y(n_317) );
OR2x2_ASAP7_75t_L g355 ( .A(n_133), .B(n_254), .Y(n_355) );
INVx2_ASAP7_75t_L g405 ( .A(n_133), .Y(n_405) );
NAND2xp5_ASAP7_75t_L g422 ( .A(n_133), .B(n_253), .Y(n_422) );
OA21x2_ASAP7_75t_L g133 ( .A1(n_134), .A2(n_139), .B(n_159), .Y(n_133) );
OA21x2_ASAP7_75t_L g163 ( .A1(n_134), .A2(n_164), .B(n_176), .Y(n_163) );
INVx2_ASAP7_75t_L g196 ( .A(n_134), .Y(n_196) );
INVx1_ASAP7_75t_L g491 ( .A(n_134), .Y(n_491) );
AOI21xp5_ASAP7_75t_L g509 ( .A1(n_134), .A2(n_510), .B(n_511), .Y(n_509) );
AOI21xp5_ASAP7_75t_L g536 ( .A1(n_134), .A2(n_537), .B(n_538), .Y(n_536) );
AND2x2_ASAP7_75t_SL g134 ( .A(n_135), .B(n_136), .Y(n_134) );
AND2x2_ASAP7_75t_L g184 ( .A(n_135), .B(n_136), .Y(n_184) );
NAND2xp5_ASAP7_75t_L g136 ( .A(n_137), .B(n_138), .Y(n_136) );
OAI21xp5_ASAP7_75t_L g139 ( .A1(n_140), .A2(n_151), .B(n_157), .Y(n_139) );
AOI21xp5_ASAP7_75t_L g140 ( .A1(n_141), .A2(n_145), .B(n_148), .Y(n_140) );
INVx3_ASAP7_75t_L g166 ( .A(n_142), .Y(n_166) );
HB1xp67_ASAP7_75t_L g529 ( .A(n_142), .Y(n_529) );
BUFx6f_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
INVx1_ASAP7_75t_L g154 ( .A(n_143), .Y(n_154) );
BUFx3_ASAP7_75t_L g194 ( .A(n_143), .Y(n_194) );
AND2x6_ASAP7_75t_L g481 ( .A(n_143), .B(n_482), .Y(n_481) );
INVx2_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
INVx1_ASAP7_75t_L g147 ( .A(n_144), .Y(n_147) );
INVx1_ASAP7_75t_L g218 ( .A(n_144), .Y(n_218) );
INVx2_ASAP7_75t_L g225 ( .A(n_146), .Y(n_225) );
INVx3_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
INVx1_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
INVx1_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
BUFx6f_ASAP7_75t_L g156 ( .A(n_150), .Y(n_156) );
INVx3_ASAP7_75t_L g170 ( .A(n_150), .Y(n_170) );
BUFx6f_ASAP7_75t_L g175 ( .A(n_150), .Y(n_175) );
AND2x2_ASAP7_75t_L g479 ( .A(n_150), .B(n_218), .Y(n_479) );
INVx1_ASAP7_75t_L g482 ( .A(n_150), .Y(n_482) );
AOI21xp5_ASAP7_75t_L g151 ( .A1(n_152), .A2(n_153), .B(n_155), .Y(n_151) );
O2A1O1Ixp5_ASAP7_75t_L g241 ( .A1(n_155), .A2(n_229), .B(n_242), .C(n_243), .Y(n_241) );
INVx2_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
OAI22xp5_ASAP7_75t_L g179 ( .A1(n_156), .A2(n_180), .B1(n_181), .B2(n_182), .Y(n_179) );
OAI22xp5_ASAP7_75t_SL g192 ( .A1(n_156), .A2(n_170), .B1(n_193), .B2(n_195), .Y(n_192) );
OAI22xp5_ASAP7_75t_L g204 ( .A1(n_156), .A2(n_181), .B1(n_205), .B2(n_206), .Y(n_204) );
INVx4_ASAP7_75t_L g502 ( .A(n_156), .Y(n_502) );
OAI21xp5_ASAP7_75t_L g164 ( .A1(n_157), .A2(n_165), .B(n_171), .Y(n_164) );
BUFx3_ASAP7_75t_L g185 ( .A(n_157), .Y(n_185) );
OAI21xp5_ASAP7_75t_L g210 ( .A1(n_157), .A2(n_211), .B(n_214), .Y(n_210) );
OAI21xp5_ASAP7_75t_L g222 ( .A1(n_157), .A2(n_223), .B(n_228), .Y(n_222) );
AND2x4_ASAP7_75t_L g478 ( .A(n_157), .B(n_479), .Y(n_478) );
INVx4_ASAP7_75t_SL g504 ( .A(n_157), .Y(n_504) );
NAND2x1p5_ASAP7_75t_L g568 ( .A(n_157), .B(n_479), .Y(n_568) );
NOR2xp67_ASAP7_75t_L g160 ( .A(n_161), .B(n_177), .Y(n_160) );
INVx1_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
HB1xp67_ASAP7_75t_L g271 ( .A(n_162), .Y(n_271) );
NAND2xp5_ASAP7_75t_L g287 ( .A(n_162), .B(n_288), .Y(n_287) );
AND2x2_ASAP7_75t_SL g337 ( .A(n_162), .B(n_277), .Y(n_337) );
INVx2_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
HB1xp67_ASAP7_75t_L g189 ( .A(n_163), .Y(n_189) );
INVx2_ASAP7_75t_L g254 ( .A(n_163), .Y(n_254) );
OR2x2_ASAP7_75t_L g316 ( .A(n_163), .B(n_317), .Y(n_316) );
O2A1O1Ixp5_ASAP7_75t_SL g165 ( .A1(n_166), .A2(n_167), .B(n_168), .C(n_169), .Y(n_165) );
INVx2_ASAP7_75t_L g181 ( .A(n_169), .Y(n_181) );
AOI21xp5_ASAP7_75t_L g211 ( .A1(n_169), .A2(n_212), .B(n_213), .Y(n_211) );
AOI21xp5_ASAP7_75t_L g238 ( .A1(n_169), .A2(n_239), .B(n_240), .Y(n_238) );
NOR2xp33_ASAP7_75t_L g551 ( .A(n_169), .B(n_552), .Y(n_551) );
INVx5_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
AOI21xp5_ASAP7_75t_L g171 ( .A1(n_172), .A2(n_173), .B(n_174), .Y(n_171) );
INVx1_ASAP7_75t_L g227 ( .A(n_174), .Y(n_227) );
INVx4_ASAP7_75t_L g174 ( .A(n_175), .Y(n_174) );
INVx2_ASAP7_75t_L g485 ( .A(n_175), .Y(n_485) );
AND2x2_ASAP7_75t_L g255 ( .A(n_177), .B(n_191), .Y(n_255) );
AND2x2_ASAP7_75t_L g272 ( .A(n_177), .B(n_252), .Y(n_272) );
INVx2_ASAP7_75t_L g177 ( .A(n_178), .Y(n_177) );
AND2x2_ASAP7_75t_L g190 ( .A(n_178), .B(n_191), .Y(n_190) );
BUFx2_ASAP7_75t_L g275 ( .A(n_178), .Y(n_275) );
AND2x2_ASAP7_75t_L g404 ( .A(n_178), .B(n_405), .Y(n_404) );
AOI21xp5_ASAP7_75t_L g214 ( .A1(n_181), .A2(n_215), .B(n_216), .Y(n_214) );
O2A1O1Ixp33_ASAP7_75t_L g228 ( .A1(n_181), .A2(n_229), .B(n_230), .C(n_231), .Y(n_228) );
INVx2_ASAP7_75t_L g221 ( .A(n_183), .Y(n_221) );
NOR2xp33_ASAP7_75t_L g573 ( .A(n_183), .B(n_574), .Y(n_573) );
INVx1_ASAP7_75t_L g183 ( .A(n_184), .Y(n_183) );
BUFx6f_ASAP7_75t_L g186 ( .A(n_184), .Y(n_186) );
NAND3xp33_ASAP7_75t_L g203 ( .A(n_185), .B(n_204), .C(n_207), .Y(n_203) );
OAI21xp5_ASAP7_75t_L g237 ( .A1(n_185), .A2(n_238), .B(n_241), .Y(n_237) );
INVx4_ASAP7_75t_L g207 ( .A(n_186), .Y(n_207) );
OA21x2_ASAP7_75t_L g209 ( .A1(n_186), .A2(n_210), .B(n_219), .Y(n_209) );
HB1xp67_ASAP7_75t_L g546 ( .A(n_186), .Y(n_546) );
AOI21xp5_ASAP7_75t_L g557 ( .A1(n_186), .A2(n_558), .B(n_559), .Y(n_557) );
INVx1_ASAP7_75t_L g249 ( .A(n_187), .Y(n_249) );
AND2x2_ASAP7_75t_L g187 ( .A(n_188), .B(n_190), .Y(n_187) );
AND2x2_ASAP7_75t_L g367 ( .A(n_188), .B(n_255), .Y(n_367) );
INVx1_ASAP7_75t_L g188 ( .A(n_189), .Y(n_188) );
AND2x2_ASAP7_75t_L g368 ( .A(n_189), .B(n_279), .Y(n_368) );
O2A1O1Ixp33_ASAP7_75t_L g335 ( .A1(n_190), .A2(n_336), .B(n_338), .C(n_340), .Y(n_335) );
NAND2xp5_ASAP7_75t_L g345 ( .A(n_190), .B(n_336), .Y(n_345) );
AOI221xp5_ASAP7_75t_L g408 ( .A1(n_190), .A2(n_266), .B1(n_409), .B2(n_410), .C(n_412), .Y(n_408) );
INVx1_ASAP7_75t_L g252 ( .A(n_191), .Y(n_252) );
INVx1_ASAP7_75t_L g288 ( .A(n_191), .Y(n_288) );
BUFx6f_ASAP7_75t_L g297 ( .A(n_191), .Y(n_297) );
INVx2_ASAP7_75t_L g503 ( .A(n_194), .Y(n_503) );
HB1xp67_ASAP7_75t_L g516 ( .A(n_194), .Y(n_516) );
INVx1_ASAP7_75t_L g488 ( .A(n_196), .Y(n_488) );
INVx1_ASAP7_75t_SL g197 ( .A(n_198), .Y(n_197) );
AND2x2_ASAP7_75t_L g198 ( .A(n_199), .B(n_208), .Y(n_198) );
AND2x2_ASAP7_75t_L g314 ( .A(n_199), .B(n_259), .Y(n_314) );
NAND2xp5_ASAP7_75t_L g333 ( .A(n_199), .B(n_334), .Y(n_333) );
INVx2_ASAP7_75t_L g199 ( .A(n_200), .Y(n_199) );
NOR2xp33_ASAP7_75t_L g282 ( .A(n_200), .B(n_283), .Y(n_282) );
OR2x2_ASAP7_75t_L g406 ( .A(n_200), .B(n_407), .Y(n_406) );
INVx1_ASAP7_75t_L g438 ( .A(n_200), .Y(n_438) );
INVx2_ASAP7_75t_L g200 ( .A(n_201), .Y(n_200) );
INVx3_ASAP7_75t_L g268 ( .A(n_201), .Y(n_268) );
AND2x2_ASAP7_75t_L g294 ( .A(n_201), .B(n_248), .Y(n_294) );
NOR2x1_ASAP7_75t_L g303 ( .A(n_201), .B(n_304), .Y(n_303) );
AND2x2_ASAP7_75t_L g310 ( .A(n_201), .B(n_311), .Y(n_310) );
AND2x4_ASAP7_75t_L g201 ( .A(n_202), .B(n_203), .Y(n_201) );
INVx1_ASAP7_75t_L g246 ( .A(n_202), .Y(n_246) );
AO21x1_ASAP7_75t_L g245 ( .A1(n_204), .A2(n_207), .B(n_246), .Y(n_245) );
INVx3_ASAP7_75t_L g494 ( .A(n_207), .Y(n_494) );
NOR2xp33_ASAP7_75t_L g518 ( .A(n_207), .B(n_519), .Y(n_518) );
AO21x2_ASAP7_75t_L g523 ( .A1(n_207), .A2(n_524), .B(n_531), .Y(n_523) );
NOR2xp33_ASAP7_75t_L g531 ( .A(n_207), .B(n_532), .Y(n_531) );
AO21x2_ASAP7_75t_L g565 ( .A1(n_207), .A2(n_566), .B(n_573), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g385 ( .A(n_208), .B(n_350), .Y(n_385) );
INVx1_ASAP7_75t_SL g389 ( .A(n_208), .Y(n_389) );
AND2x2_ASAP7_75t_L g208 ( .A(n_209), .B(n_220), .Y(n_208) );
INVx3_ASAP7_75t_L g248 ( .A(n_209), .Y(n_248) );
AND2x2_ASAP7_75t_L g259 ( .A(n_209), .B(n_236), .Y(n_259) );
AND2x2_ASAP7_75t_L g281 ( .A(n_209), .B(n_282), .Y(n_281) );
AND2x2_ASAP7_75t_L g326 ( .A(n_209), .B(n_320), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g407 ( .A(n_209), .B(n_258), .Y(n_407) );
INVx2_ASAP7_75t_L g229 ( .A(n_217), .Y(n_229) );
INVx1_ASAP7_75t_L g217 ( .A(n_218), .Y(n_217) );
AND2x2_ASAP7_75t_L g247 ( .A(n_220), .B(n_248), .Y(n_247) );
INVx2_ASAP7_75t_L g258 ( .A(n_220), .Y(n_258) );
NAND2xp5_ASAP7_75t_L g283 ( .A(n_220), .B(n_236), .Y(n_283) );
AND2x2_ASAP7_75t_L g319 ( .A(n_220), .B(n_320), .Y(n_319) );
OA21x2_ASAP7_75t_L g220 ( .A1(n_221), .A2(n_222), .B(n_232), .Y(n_220) );
OA21x2_ASAP7_75t_L g236 ( .A1(n_221), .A2(n_237), .B(n_244), .Y(n_236) );
O2A1O1Ixp33_ASAP7_75t_L g223 ( .A1(n_224), .A2(n_225), .B(n_226), .C(n_227), .Y(n_223) );
AOI21xp5_ASAP7_75t_L g560 ( .A1(n_225), .A2(n_561), .B(n_562), .Y(n_560) );
AOI21xp5_ASAP7_75t_L g570 ( .A1(n_225), .A2(n_571), .B(n_572), .Y(n_570) );
O2A1O1Ixp33_ASAP7_75t_L g526 ( .A1(n_227), .A2(n_527), .B(n_528), .C(n_529), .Y(n_526) );
AOI21xp5_ASAP7_75t_L g483 ( .A1(n_229), .A2(n_484), .B(n_486), .Y(n_483) );
INVx1_ASAP7_75t_L g233 ( .A(n_234), .Y(n_233) );
AND2x2_ASAP7_75t_L g234 ( .A(n_235), .B(n_247), .Y(n_234) );
INVx1_ASAP7_75t_L g299 ( .A(n_235), .Y(n_299) );
AND2x2_ASAP7_75t_L g341 ( .A(n_235), .B(n_342), .Y(n_341) );
NAND2xp5_ASAP7_75t_SL g347 ( .A(n_235), .B(n_262), .Y(n_347) );
AOI21xp5_ASAP7_75t_SL g421 ( .A1(n_235), .A2(n_253), .B(n_276), .Y(n_421) );
AND2x2_ASAP7_75t_L g235 ( .A(n_236), .B(n_245), .Y(n_235) );
OR2x2_ASAP7_75t_L g264 ( .A(n_236), .B(n_245), .Y(n_264) );
AND2x2_ASAP7_75t_L g311 ( .A(n_236), .B(n_248), .Y(n_311) );
INVx2_ASAP7_75t_L g320 ( .A(n_236), .Y(n_320) );
INVx1_ASAP7_75t_L g426 ( .A(n_236), .Y(n_426) );
AND2x2_ASAP7_75t_L g350 ( .A(n_245), .B(n_320), .Y(n_350) );
INVx1_ASAP7_75t_L g375 ( .A(n_245), .Y(n_375) );
AND2x2_ASAP7_75t_L g284 ( .A(n_247), .B(n_268), .Y(n_284) );
AND2x2_ASAP7_75t_L g296 ( .A(n_247), .B(n_297), .Y(n_296) );
INVx2_ASAP7_75t_SL g414 ( .A(n_247), .Y(n_414) );
INVx2_ASAP7_75t_L g304 ( .A(n_248), .Y(n_304) );
AND2x2_ASAP7_75t_L g342 ( .A(n_248), .B(n_258), .Y(n_342) );
NAND2xp5_ASAP7_75t_L g425 ( .A(n_248), .B(n_426), .Y(n_425) );
OAI21xp33_ASAP7_75t_L g250 ( .A1(n_251), .A2(n_255), .B(n_256), .Y(n_250) );
AND2x2_ASAP7_75t_L g357 ( .A(n_251), .B(n_358), .Y(n_357) );
INVx1_ASAP7_75t_L g411 ( .A(n_251), .Y(n_411) );
AND2x2_ASAP7_75t_L g251 ( .A(n_252), .B(n_253), .Y(n_251) );
INVx1_ASAP7_75t_L g331 ( .A(n_252), .Y(n_331) );
BUFx2_ASAP7_75t_L g430 ( .A(n_252), .Y(n_430) );
BUFx2_ASAP7_75t_L g301 ( .A(n_253), .Y(n_301) );
AND2x2_ASAP7_75t_L g403 ( .A(n_253), .B(n_404), .Y(n_403) );
INVx2_ASAP7_75t_L g253 ( .A(n_254), .Y(n_253) );
INVx1_ASAP7_75t_L g386 ( .A(n_254), .Y(n_386) );
AND2x4_ASAP7_75t_L g313 ( .A(n_255), .B(n_276), .Y(n_313) );
NAND2xp5_ASAP7_75t_SL g349 ( .A(n_255), .B(n_337), .Y(n_349) );
AOI32xp33_ASAP7_75t_L g273 ( .A1(n_256), .A2(n_274), .A3(n_276), .B1(n_278), .B2(n_279), .Y(n_273) );
AND2x2_ASAP7_75t_L g256 ( .A(n_257), .B(n_259), .Y(n_256) );
INVx3_ASAP7_75t_L g262 ( .A(n_257), .Y(n_262) );
OR2x2_ASAP7_75t_L g398 ( .A(n_257), .B(n_354), .Y(n_398) );
INVx2_ASAP7_75t_L g257 ( .A(n_258), .Y(n_257) );
AND2x2_ASAP7_75t_L g267 ( .A(n_258), .B(n_268), .Y(n_267) );
AND2x2_ASAP7_75t_L g374 ( .A(n_258), .B(n_375), .Y(n_374) );
AND2x2_ASAP7_75t_L g266 ( .A(n_259), .B(n_267), .Y(n_266) );
AND2x2_ASAP7_75t_L g278 ( .A(n_259), .B(n_268), .Y(n_278) );
INVx1_ASAP7_75t_L g399 ( .A(n_259), .Y(n_399) );
NAND2xp5_ASAP7_75t_L g432 ( .A(n_259), .B(n_374), .Y(n_432) );
A2O1A1Ixp33_ASAP7_75t_L g260 ( .A1(n_261), .A2(n_265), .B(n_269), .C(n_273), .Y(n_260) );
OAI322xp33_ASAP7_75t_L g369 ( .A1(n_261), .A2(n_306), .A3(n_370), .B1(n_372), .B2(n_376), .C1(n_377), .C2(n_381), .Y(n_369) );
NAND2xp5_ASAP7_75t_L g261 ( .A(n_262), .B(n_263), .Y(n_261) );
INVxp67_ASAP7_75t_L g334 ( .A(n_262), .Y(n_334) );
INVx1_ASAP7_75t_SL g263 ( .A(n_264), .Y(n_263) );
OR2x2_ASAP7_75t_L g388 ( .A(n_264), .B(n_389), .Y(n_388) );
NOR2xp33_ASAP7_75t_L g435 ( .A(n_264), .B(n_304), .Y(n_435) );
INVxp67_ASAP7_75t_L g265 ( .A(n_266), .Y(n_265) );
INVx1_ASAP7_75t_L g327 ( .A(n_267), .Y(n_327) );
OR2x2_ASAP7_75t_L g413 ( .A(n_268), .B(n_414), .Y(n_413) );
INVx1_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
AND2x2_ASAP7_75t_L g270 ( .A(n_271), .B(n_272), .Y(n_270) );
NAND2xp5_ASAP7_75t_L g329 ( .A(n_271), .B(n_330), .Y(n_329) );
AND2x2_ASAP7_75t_L g322 ( .A(n_272), .B(n_301), .Y(n_322) );
AND2x2_ASAP7_75t_L g393 ( .A(n_272), .B(n_306), .Y(n_393) );
NAND2xp5_ASAP7_75t_L g415 ( .A(n_272), .B(n_380), .Y(n_415) );
AOI221xp5_ASAP7_75t_L g280 ( .A1(n_274), .A2(n_281), .B1(n_284), .B2(n_285), .C(n_290), .Y(n_280) );
OR2x2_ASAP7_75t_L g291 ( .A(n_274), .B(n_287), .Y(n_291) );
AND2x2_ASAP7_75t_L g379 ( .A(n_274), .B(n_380), .Y(n_379) );
AOI32xp33_ASAP7_75t_L g418 ( .A1(n_274), .A2(n_304), .A3(n_419), .B1(n_420), .B2(n_423), .Y(n_418) );
INVx2_ASAP7_75t_L g274 ( .A(n_275), .Y(n_274) );
NAND3xp33_ASAP7_75t_L g352 ( .A(n_275), .B(n_311), .C(n_334), .Y(n_352) );
AND2x2_ASAP7_75t_L g378 ( .A(n_275), .B(n_371), .Y(n_378) );
INVxp67_ASAP7_75t_L g358 ( .A(n_276), .Y(n_358) );
BUFx3_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
NAND2xp5_ASAP7_75t_SL g387 ( .A(n_279), .B(n_331), .Y(n_387) );
INVx2_ASAP7_75t_L g397 ( .A(n_279), .Y(n_397) );
NOR2xp33_ASAP7_75t_L g410 ( .A(n_279), .B(n_411), .Y(n_410) );
INVx1_ASAP7_75t_L g366 ( .A(n_282), .Y(n_366) );
OR2x2_ASAP7_75t_L g292 ( .A(n_283), .B(n_293), .Y(n_292) );
NOR2xp33_ASAP7_75t_L g402 ( .A(n_285), .B(n_403), .Y(n_402) );
AND2x2_ASAP7_75t_L g285 ( .A(n_286), .B(n_289), .Y(n_285) );
INVx1_ASAP7_75t_SL g286 ( .A(n_287), .Y(n_286) );
HB1xp67_ASAP7_75t_L g371 ( .A(n_288), .Y(n_371) );
AND2x2_ASAP7_75t_L g330 ( .A(n_289), .B(n_331), .Y(n_330) );
INVx1_ASAP7_75t_L g376 ( .A(n_289), .Y(n_376) );
HB1xp67_ASAP7_75t_L g401 ( .A(n_289), .Y(n_401) );
NOR2xp33_ASAP7_75t_L g290 ( .A(n_291), .B(n_292), .Y(n_290) );
AOI21xp33_ASAP7_75t_SL g315 ( .A1(n_291), .A2(n_316), .B(n_318), .Y(n_315) );
INVx1_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
AND2x2_ASAP7_75t_L g409 ( .A(n_294), .B(n_319), .Y(n_409) );
AOI211xp5_ASAP7_75t_L g295 ( .A1(n_296), .A2(n_298), .B(n_308), .C(n_315), .Y(n_295) );
AND2x2_ASAP7_75t_L g339 ( .A(n_297), .B(n_307), .Y(n_339) );
INVx2_ASAP7_75t_L g354 ( .A(n_297), .Y(n_354) );
OR2x2_ASAP7_75t_L g392 ( .A(n_297), .B(n_355), .Y(n_392) );
NAND2xp5_ASAP7_75t_L g434 ( .A(n_297), .B(n_435), .Y(n_434) );
AOI211xp5_ASAP7_75t_SL g298 ( .A1(n_299), .A2(n_300), .B(n_302), .C(n_305), .Y(n_298) );
INVxp67_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g338 ( .A(n_301), .B(n_339), .Y(n_338) );
OAI211xp5_ASAP7_75t_L g420 ( .A1(n_302), .A2(n_397), .B(n_421), .C(n_422), .Y(n_420) );
INVx1_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
NAND2x1p5_ASAP7_75t_L g318 ( .A(n_303), .B(n_319), .Y(n_318) );
AND2x2_ASAP7_75t_L g360 ( .A(n_304), .B(n_350), .Y(n_360) );
INVx1_ASAP7_75t_L g365 ( .A(n_304), .Y(n_365) );
INVx1_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
INVx1_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
NAND2xp5_ASAP7_75t_SL g308 ( .A(n_309), .B(n_312), .Y(n_308) );
INVxp33_ASAP7_75t_L g416 ( .A(n_310), .Y(n_416) );
AND2x2_ASAP7_75t_L g395 ( .A(n_311), .B(n_374), .Y(n_395) );
NAND2xp5_ASAP7_75t_L g312 ( .A(n_313), .B(n_314), .Y(n_312) );
AOI21xp5_ASAP7_75t_L g377 ( .A1(n_316), .A2(n_378), .B(n_379), .Y(n_377) );
OAI322xp33_ASAP7_75t_L g396 ( .A1(n_318), .A2(n_397), .A3(n_398), .B1(n_399), .B2(n_400), .C1(n_402), .C2(n_406), .Y(n_396) );
AOI221xp5_ASAP7_75t_L g321 ( .A1(n_322), .A2(n_323), .B1(n_328), .B2(n_332), .C(n_335), .Y(n_321) );
INVx2_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
OR2x2_ASAP7_75t_L g324 ( .A(n_325), .B(n_327), .Y(n_324) );
INVx1_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
AND2x2_ASAP7_75t_L g373 ( .A(n_326), .B(n_374), .Y(n_373) );
INVx1_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
INVx1_ASAP7_75t_L g417 ( .A(n_330), .Y(n_417) );
INVxp67_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
NOR2xp33_ASAP7_75t_L g419 ( .A(n_333), .B(n_353), .Y(n_419) );
INVx2_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
INVx1_ASAP7_75t_SL g340 ( .A(n_341), .Y(n_340) );
AND2x2_ASAP7_75t_L g382 ( .A(n_342), .B(n_350), .Y(n_382) );
AOI221xp5_ASAP7_75t_L g343 ( .A1(n_344), .A2(n_346), .B1(n_348), .B2(n_350), .C(n_351), .Y(n_343) );
INVx1_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
AOI221xp5_ASAP7_75t_L g362 ( .A1(n_346), .A2(n_363), .B1(n_367), .B2(n_368), .C(n_369), .Y(n_362) );
INVx1_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
INVxp67_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
NAND2xp5_ASAP7_75t_L g364 ( .A(n_350), .B(n_365), .Y(n_364) );
OAI22xp5_ASAP7_75t_L g351 ( .A1(n_352), .A2(n_353), .B1(n_356), .B2(n_359), .Y(n_351) );
OR2x2_ASAP7_75t_L g353 ( .A(n_354), .B(n_355), .Y(n_353) );
INVx2_ASAP7_75t_SL g380 ( .A(n_355), .Y(n_380) );
INVxp67_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
INVx1_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
NAND5xp2_ASAP7_75t_L g361 ( .A(n_362), .B(n_383), .C(n_408), .D(n_418), .E(n_428), .Y(n_361) );
NAND2xp5_ASAP7_75t_SL g363 ( .A(n_364), .B(n_366), .Y(n_363) );
NOR4xp25_ASAP7_75t_L g436 ( .A(n_365), .B(n_371), .C(n_437), .D(n_438), .Y(n_436) );
AOI221xp5_ASAP7_75t_L g428 ( .A1(n_368), .A2(n_429), .B1(n_431), .B2(n_433), .C(n_436), .Y(n_428) );
INVx1_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
INVx1_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
INVx1_ASAP7_75t_L g427 ( .A(n_374), .Y(n_427) );
OAI322xp33_ASAP7_75t_L g384 ( .A1(n_378), .A2(n_385), .A3(n_386), .B1(n_387), .B2(n_388), .C1(n_390), .C2(n_394), .Y(n_384) );
INVx1_ASAP7_75t_SL g381 ( .A(n_382), .Y(n_381) );
NOR2xp33_ASAP7_75t_L g383 ( .A(n_384), .B(n_396), .Y(n_383) );
NOR2xp33_ASAP7_75t_L g390 ( .A(n_391), .B(n_393), .Y(n_390) );
INVx2_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
INVx1_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
INVx1_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
AND2x2_ASAP7_75t_L g429 ( .A(n_404), .B(n_430), .Y(n_429) );
OAI22xp33_ASAP7_75t_L g412 ( .A1(n_413), .A2(n_415), .B1(n_416), .B2(n_417), .Y(n_412) );
INVx1_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
OR2x2_ASAP7_75t_L g424 ( .A(n_425), .B(n_427), .Y(n_424) );
INVx1_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
INVxp67_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
INVx1_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
NOR2xp33_ASAP7_75t_L g444 ( .A(n_445), .B(n_446), .Y(n_444) );
INVx1_ASAP7_75t_SL g447 ( .A(n_448), .Y(n_447) );
INVx2_ASAP7_75t_L g455 ( .A(n_448), .Y(n_455) );
INVx2_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
AND2x2_ASAP7_75t_L g450 ( .A(n_451), .B(n_452), .Y(n_450) );
INVx1_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
NAND3xp33_ASAP7_75t_L g457 ( .A(n_456), .B(n_458), .C(n_771), .Y(n_457) );
OAI22x1_ASAP7_75t_SL g459 ( .A1(n_460), .A2(n_462), .B1(n_465), .B2(n_756), .Y(n_459) );
INVx1_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
OAI22xp5_ASAP7_75t_SL g766 ( .A1(n_461), .A2(n_466), .B1(n_756), .B2(n_767), .Y(n_766) );
INVx2_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
INVx2_ASAP7_75t_L g767 ( .A(n_463), .Y(n_767) );
INVx1_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
INVx2_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
AND2x2_ASAP7_75t_SL g466 ( .A(n_467), .B(n_711), .Y(n_466) );
NOR2xp33_ASAP7_75t_L g467 ( .A(n_468), .B(n_646), .Y(n_467) );
NAND4xp25_ASAP7_75t_SL g468 ( .A(n_469), .B(n_591), .C(n_615), .D(n_638), .Y(n_468) );
AOI221xp5_ASAP7_75t_L g469 ( .A1(n_470), .A2(n_533), .B1(n_563), .B2(n_575), .C(n_578), .Y(n_469) );
INVx1_ASAP7_75t_L g470 ( .A(n_471), .Y(n_470) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_472), .B(n_506), .Y(n_471) );
AOI22xp33_ASAP7_75t_L g581 ( .A1(n_472), .A2(n_492), .B1(n_534), .B2(n_582), .Y(n_581) );
NAND2xp5_ASAP7_75t_L g649 ( .A(n_472), .B(n_507), .Y(n_649) );
AND2x2_ASAP7_75t_L g668 ( .A(n_472), .B(n_669), .Y(n_668) );
NAND2xp5_ASAP7_75t_L g738 ( .A(n_472), .B(n_652), .Y(n_738) );
AND2x4_ASAP7_75t_L g472 ( .A(n_473), .B(n_492), .Y(n_472) );
AND2x2_ASAP7_75t_L g606 ( .A(n_473), .B(n_507), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g620 ( .A(n_473), .B(n_621), .Y(n_620) );
OR2x2_ASAP7_75t_L g629 ( .A(n_473), .B(n_630), .Y(n_629) );
AND2x2_ASAP7_75t_L g634 ( .A(n_473), .B(n_493), .Y(n_634) );
INVx2_ASAP7_75t_L g666 ( .A(n_473), .Y(n_666) );
HB1xp67_ASAP7_75t_L g710 ( .A(n_473), .Y(n_710) );
AND2x2_ASAP7_75t_L g727 ( .A(n_473), .B(n_604), .Y(n_727) );
INVx5_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
AND2x2_ASAP7_75t_L g645 ( .A(n_474), .B(n_604), .Y(n_645) );
AND2x4_ASAP7_75t_L g659 ( .A(n_474), .B(n_492), .Y(n_659) );
HB1xp67_ASAP7_75t_L g663 ( .A(n_474), .Y(n_663) );
AND2x2_ASAP7_75t_L g683 ( .A(n_474), .B(n_598), .Y(n_683) );
AND2x2_ASAP7_75t_L g733 ( .A(n_474), .B(n_508), .Y(n_733) );
AND2x2_ASAP7_75t_L g743 ( .A(n_474), .B(n_493), .Y(n_743) );
OR2x6_ASAP7_75t_L g474 ( .A(n_475), .B(n_489), .Y(n_474) );
AOI21xp5_ASAP7_75t_SL g475 ( .A1(n_476), .A2(n_480), .B(n_488), .Y(n_475) );
BUFx2_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
INVx5_ASAP7_75t_L g498 ( .A(n_481), .Y(n_498) );
INVx2_ASAP7_75t_L g487 ( .A(n_485), .Y(n_487) );
O2A1O1Ixp33_ASAP7_75t_L g513 ( .A1(n_487), .A2(n_514), .B(n_515), .C(n_516), .Y(n_513) );
O2A1O1Ixp33_ASAP7_75t_L g539 ( .A1(n_487), .A2(n_516), .B(n_540), .C(n_541), .Y(n_539) );
NOR2xp33_ASAP7_75t_L g489 ( .A(n_490), .B(n_491), .Y(n_489) );
AND2x2_ASAP7_75t_L g599 ( .A(n_492), .B(n_507), .Y(n_599) );
HB1xp67_ASAP7_75t_L g614 ( .A(n_492), .Y(n_614) );
NAND2xp5_ASAP7_75t_L g640 ( .A(n_492), .B(n_641), .Y(n_640) );
INVx1_ASAP7_75t_L g689 ( .A(n_492), .Y(n_689) );
INVx2_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
AND2x2_ASAP7_75t_L g577 ( .A(n_493), .B(n_522), .Y(n_577) );
AND2x2_ASAP7_75t_L g604 ( .A(n_493), .B(n_523), .Y(n_604) );
OA21x2_ASAP7_75t_L g493 ( .A1(n_494), .A2(n_495), .B(n_505), .Y(n_493) );
O2A1O1Ixp33_ASAP7_75t_SL g496 ( .A1(n_497), .A2(n_498), .B(n_499), .C(n_504), .Y(n_496) );
INVx2_ASAP7_75t_L g512 ( .A(n_498), .Y(n_512) );
O2A1O1Ixp33_ASAP7_75t_L g548 ( .A1(n_498), .A2(n_504), .B(n_549), .C(n_550), .Y(n_548) );
NOR2xp33_ASAP7_75t_L g500 ( .A(n_501), .B(n_502), .Y(n_500) );
INVx1_ASAP7_75t_L g517 ( .A(n_504), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g662 ( .A(n_506), .B(n_663), .Y(n_662) );
AND2x2_ASAP7_75t_L g506 ( .A(n_507), .B(n_520), .Y(n_506) );
OR2x2_ASAP7_75t_L g630 ( .A(n_507), .B(n_521), .Y(n_630) );
AND2x2_ASAP7_75t_L g667 ( .A(n_507), .B(n_577), .Y(n_667) );
NAND2xp5_ASAP7_75t_L g678 ( .A(n_507), .B(n_598), .Y(n_678) );
HB1xp67_ASAP7_75t_L g682 ( .A(n_507), .Y(n_682) );
NAND2xp5_ASAP7_75t_L g751 ( .A(n_507), .B(n_634), .Y(n_751) );
INVx5_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
BUFx2_ASAP7_75t_L g576 ( .A(n_508), .Y(n_576) );
AND2x2_ASAP7_75t_L g585 ( .A(n_508), .B(n_521), .Y(n_585) );
AND2x2_ASAP7_75t_L g701 ( .A(n_508), .B(n_596), .Y(n_701) );
NAND2xp5_ASAP7_75t_L g723 ( .A(n_508), .B(n_634), .Y(n_723) );
OR2x6_ASAP7_75t_L g508 ( .A(n_509), .B(n_518), .Y(n_508) );
INVx1_ASAP7_75t_L g520 ( .A(n_521), .Y(n_520) );
HB1xp67_ASAP7_75t_L g669 ( .A(n_521), .Y(n_669) );
INVx2_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
HB1xp67_ASAP7_75t_L g621 ( .A(n_522), .Y(n_621) );
INVx2_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
BUFx2_ASAP7_75t_L g598 ( .A(n_523), .Y(n_598) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_525), .B(n_530), .Y(n_524) );
NOR2xp33_ASAP7_75t_L g533 ( .A(n_534), .B(n_543), .Y(n_533) );
NOR2xp33_ASAP7_75t_L g730 ( .A(n_534), .B(n_611), .Y(n_730) );
HB1xp67_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
NOR2xp33_ASAP7_75t_L g563 ( .A(n_535), .B(n_564), .Y(n_563) );
AND2x2_ASAP7_75t_L g582 ( .A(n_535), .B(n_583), .Y(n_582) );
INVx5_ASAP7_75t_SL g590 ( .A(n_535), .Y(n_590) );
OR2x2_ASAP7_75t_L g613 ( .A(n_535), .B(n_583), .Y(n_613) );
OR2x2_ASAP7_75t_L g623 ( .A(n_535), .B(n_624), .Y(n_623) );
AND2x2_ASAP7_75t_L g686 ( .A(n_535), .B(n_545), .Y(n_686) );
AND2x2_ASAP7_75t_SL g724 ( .A(n_535), .B(n_544), .Y(n_724) );
NOR4xp25_ASAP7_75t_L g745 ( .A(n_535), .B(n_666), .C(n_746), .D(n_747), .Y(n_745) );
AND2x2_ASAP7_75t_L g755 ( .A(n_535), .B(n_587), .Y(n_755) );
OR2x6_ASAP7_75t_L g535 ( .A(n_536), .B(n_542), .Y(n_535) );
INVx2_ASAP7_75t_L g543 ( .A(n_544), .Y(n_543) );
AND2x2_ASAP7_75t_L g580 ( .A(n_544), .B(n_576), .Y(n_580) );
NAND2xp5_ASAP7_75t_L g749 ( .A(n_544), .B(n_582), .Y(n_749) );
AND2x2_ASAP7_75t_L g544 ( .A(n_545), .B(n_554), .Y(n_544) );
OR2x2_ASAP7_75t_L g589 ( .A(n_545), .B(n_590), .Y(n_589) );
INVx3_ASAP7_75t_L g596 ( .A(n_545), .Y(n_596) );
NAND2xp5_ASAP7_75t_L g608 ( .A(n_545), .B(n_565), .Y(n_608) );
INVxp67_ASAP7_75t_L g611 ( .A(n_545), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g624 ( .A(n_545), .B(n_583), .Y(n_624) );
NAND2xp5_ASAP7_75t_L g677 ( .A(n_545), .B(n_555), .Y(n_677) );
AND2x2_ASAP7_75t_L g692 ( .A(n_545), .B(n_587), .Y(n_692) );
OR2x2_ASAP7_75t_L g721 ( .A(n_545), .B(n_555), .Y(n_721) );
OA21x2_ASAP7_75t_L g545 ( .A1(n_546), .A2(n_547), .B(n_553), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g625 ( .A(n_554), .B(n_626), .Y(n_625) );
NOR2xp33_ASAP7_75t_L g729 ( .A(n_554), .B(n_590), .Y(n_729) );
OR2x2_ASAP7_75t_L g750 ( .A(n_554), .B(n_627), .Y(n_750) );
INVx1_ASAP7_75t_SL g554 ( .A(n_555), .Y(n_554) );
OR2x2_ASAP7_75t_L g564 ( .A(n_555), .B(n_565), .Y(n_564) );
AND2x2_ASAP7_75t_L g587 ( .A(n_555), .B(n_583), .Y(n_587) );
NAND2xp5_ASAP7_75t_SL g602 ( .A(n_555), .B(n_565), .Y(n_602) );
AND2x2_ASAP7_75t_L g672 ( .A(n_555), .B(n_596), .Y(n_672) );
AND2x2_ASAP7_75t_L g706 ( .A(n_555), .B(n_590), .Y(n_706) );
INVx2_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g609 ( .A(n_556), .B(n_590), .Y(n_609) );
AND2x2_ASAP7_75t_L g637 ( .A(n_556), .B(n_565), .Y(n_637) );
NAND2xp5_ASAP7_75t_L g644 ( .A(n_563), .B(n_645), .Y(n_644) );
AOI221xp5_ASAP7_75t_L g704 ( .A1(n_564), .A2(n_652), .B1(n_688), .B2(n_705), .C(n_707), .Y(n_704) );
INVx5_ASAP7_75t_SL g583 ( .A(n_565), .Y(n_583) );
OAI21xp5_ASAP7_75t_L g566 ( .A1(n_567), .A2(n_568), .B(n_569), .Y(n_566) );
AND2x2_ASAP7_75t_L g575 ( .A(n_576), .B(n_577), .Y(n_575) );
OAI33xp33_ASAP7_75t_L g603 ( .A1(n_576), .A2(n_604), .A3(n_605), .B1(n_607), .B2(n_610), .B3(n_614), .Y(n_603) );
OR2x2_ASAP7_75t_L g619 ( .A(n_576), .B(n_620), .Y(n_619) );
AOI322xp5_ASAP7_75t_L g728 ( .A1(n_576), .A2(n_645), .A3(n_652), .B1(n_729), .B2(n_730), .C1(n_731), .C2(n_734), .Y(n_728) );
NAND2xp5_ASAP7_75t_L g746 ( .A(n_576), .B(n_604), .Y(n_746) );
A2O1A1Ixp33_ASAP7_75t_SL g752 ( .A1(n_576), .A2(n_604), .B(n_753), .C(n_755), .Y(n_752) );
AOI221xp5_ASAP7_75t_L g591 ( .A1(n_577), .A2(n_592), .B1(n_597), .B2(n_600), .C(n_603), .Y(n_591) );
INVx1_ASAP7_75t_L g684 ( .A(n_577), .Y(n_684) );
NAND2xp5_ASAP7_75t_L g732 ( .A(n_577), .B(n_733), .Y(n_732) );
OAI22xp33_ASAP7_75t_L g578 ( .A1(n_579), .A2(n_581), .B1(n_584), .B2(n_586), .Y(n_578) );
INVx1_ASAP7_75t_SL g579 ( .A(n_580), .Y(n_579) );
AND2x2_ASAP7_75t_L g661 ( .A(n_582), .B(n_596), .Y(n_661) );
AND2x2_ASAP7_75t_L g719 ( .A(n_582), .B(n_720), .Y(n_719) );
OR2x2_ASAP7_75t_L g627 ( .A(n_583), .B(n_590), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g655 ( .A(n_583), .B(n_596), .Y(n_655) );
INVx1_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
NAND2xp5_ASAP7_75t_L g657 ( .A(n_585), .B(n_658), .Y(n_657) );
NAND2xp5_ASAP7_75t_L g717 ( .A(n_585), .B(n_663), .Y(n_717) );
OAI321xp33_ASAP7_75t_L g736 ( .A1(n_585), .A2(n_658), .A3(n_737), .B1(n_738), .B2(n_739), .C(n_740), .Y(n_736) );
INVx1_ASAP7_75t_L g703 ( .A(n_586), .Y(n_703) );
NAND2xp5_ASAP7_75t_L g586 ( .A(n_587), .B(n_588), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g593 ( .A(n_587), .B(n_594), .Y(n_593) );
AND2x2_ASAP7_75t_L g642 ( .A(n_587), .B(n_590), .Y(n_642) );
AOI321xp33_ASAP7_75t_L g700 ( .A1(n_587), .A2(n_604), .A3(n_701), .B1(n_702), .B2(n_703), .C(n_704), .Y(n_700) );
INVx1_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
OR2x2_ASAP7_75t_L g617 ( .A(n_589), .B(n_602), .Y(n_617) );
NAND2xp5_ASAP7_75t_L g595 ( .A(n_590), .B(n_596), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g671 ( .A(n_590), .B(n_672), .Y(n_671) );
NAND2xp5_ASAP7_75t_L g713 ( .A(n_590), .B(n_676), .Y(n_713) );
INVx1_ASAP7_75t_L g592 ( .A(n_593), .Y(n_592) );
AND2x4_ASAP7_75t_L g636 ( .A(n_594), .B(n_637), .Y(n_636) );
INVx2_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
OR2x2_ASAP7_75t_L g601 ( .A(n_595), .B(n_602), .Y(n_601) );
INVx1_ASAP7_75t_L g709 ( .A(n_596), .Y(n_709) );
AND2x2_ASAP7_75t_L g597 ( .A(n_598), .B(n_599), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g651 ( .A(n_599), .B(n_652), .Y(n_651) );
INVx2_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
INVx1_ASAP7_75t_L g632 ( .A(n_604), .Y(n_632) );
INVx1_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
NOR2xp33_ASAP7_75t_L g690 ( .A(n_606), .B(n_641), .Y(n_690) );
OR2x2_ASAP7_75t_L g607 ( .A(n_608), .B(n_609), .Y(n_607) );
OR2x2_ASAP7_75t_L g654 ( .A(n_609), .B(n_655), .Y(n_654) );
INVx1_ASAP7_75t_SL g699 ( .A(n_609), .Y(n_699) );
OAI22xp5_ASAP7_75t_L g656 ( .A1(n_610), .A2(n_657), .B1(n_660), .B2(n_662), .Y(n_656) );
NAND2xp5_ASAP7_75t_L g610 ( .A(n_611), .B(n_612), .Y(n_610) );
INVx1_ASAP7_75t_SL g612 ( .A(n_613), .Y(n_612) );
OR2x2_ASAP7_75t_L g754 ( .A(n_613), .B(n_677), .Y(n_754) );
AOI221xp5_ASAP7_75t_L g615 ( .A1(n_616), .A2(n_618), .B1(n_622), .B2(n_628), .C(n_631), .Y(n_615) );
INVx1_ASAP7_75t_SL g616 ( .A(n_617), .Y(n_616) );
INVx2_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
BUFx2_ASAP7_75t_L g652 ( .A(n_621), .Y(n_652) );
NAND2xp5_ASAP7_75t_L g622 ( .A(n_623), .B(n_625), .Y(n_622) );
INVx1_ASAP7_75t_SL g698 ( .A(n_624), .Y(n_698) );
NAND2xp5_ASAP7_75t_L g675 ( .A(n_626), .B(n_676), .Y(n_675) );
AOI21xp5_ASAP7_75t_L g693 ( .A1(n_626), .A2(n_694), .B(n_696), .Y(n_693) );
INVx2_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
OR2x2_ASAP7_75t_L g739 ( .A(n_627), .B(n_721), .Y(n_739) );
INVx1_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
INVx2_ASAP7_75t_SL g641 ( .A(n_630), .Y(n_641) );
AOI21xp33_ASAP7_75t_L g631 ( .A1(n_632), .A2(n_633), .B(n_635), .Y(n_631) );
INVx1_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
INVx2_ASAP7_75t_SL g635 ( .A(n_636), .Y(n_635) );
AND2x2_ASAP7_75t_L g685 ( .A(n_637), .B(n_686), .Y(n_685) );
INVxp67_ASAP7_75t_L g747 ( .A(n_637), .Y(n_747) );
AOI21xp5_ASAP7_75t_L g638 ( .A1(n_639), .A2(n_642), .B(n_643), .Y(n_638) );
INVx1_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
NAND2xp5_ASAP7_75t_L g695 ( .A(n_641), .B(n_659), .Y(n_695) );
INVxp67_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
INVx1_ASAP7_75t_L g716 ( .A(n_645), .Y(n_716) );
NAND5xp2_ASAP7_75t_L g646 ( .A(n_647), .B(n_664), .C(n_673), .D(n_693), .E(n_700), .Y(n_646) );
O2A1O1Ixp33_ASAP7_75t_L g647 ( .A1(n_648), .A2(n_650), .B(n_653), .C(n_656), .Y(n_647) );
INVx1_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
INVx1_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
INVx1_ASAP7_75t_L g688 ( .A(n_652), .Y(n_688) );
CKINVDCx16_ASAP7_75t_R g653 ( .A(n_654), .Y(n_653) );
INVx1_ASAP7_75t_SL g658 ( .A(n_659), .Y(n_658) );
NOR2xp33_ASAP7_75t_L g725 ( .A(n_660), .B(n_726), .Y(n_725) );
INVx1_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
INVx1_ASAP7_75t_L g702 ( .A(n_662), .Y(n_702) );
OAI21xp5_ASAP7_75t_SL g664 ( .A1(n_665), .A2(n_668), .B(n_670), .Y(n_664) );
AOI221xp5_ASAP7_75t_L g718 ( .A1(n_665), .A2(n_719), .B1(n_722), .B2(n_724), .C(n_725), .Y(n_718) );
AND2x2_ASAP7_75t_L g665 ( .A(n_666), .B(n_667), .Y(n_665) );
AOI321xp33_ASAP7_75t_L g673 ( .A1(n_666), .A2(n_674), .A3(n_678), .B1(n_679), .B2(n_685), .C(n_687), .Y(n_673) );
INVx1_ASAP7_75t_L g670 ( .A(n_671), .Y(n_670) );
INVx1_ASAP7_75t_L g674 ( .A(n_675), .Y(n_674) );
INVx1_ASAP7_75t_SL g676 ( .A(n_677), .Y(n_676) );
INVx1_ASAP7_75t_L g744 ( .A(n_678), .Y(n_744) );
NAND2xp5_ASAP7_75t_SL g679 ( .A(n_680), .B(n_684), .Y(n_679) );
INVx1_ASAP7_75t_L g680 ( .A(n_681), .Y(n_680) );
AND2x2_ASAP7_75t_L g696 ( .A(n_681), .B(n_697), .Y(n_696) );
AND2x2_ASAP7_75t_L g681 ( .A(n_682), .B(n_683), .Y(n_681) );
NOR2xp67_ASAP7_75t_SL g708 ( .A(n_682), .B(n_689), .Y(n_708) );
AOI321xp33_ASAP7_75t_SL g740 ( .A1(n_685), .A2(n_741), .A3(n_742), .B1(n_743), .B2(n_744), .C(n_745), .Y(n_740) );
O2A1O1Ixp33_ASAP7_75t_L g687 ( .A1(n_688), .A2(n_689), .B(n_690), .C(n_691), .Y(n_687) );
INVx1_ASAP7_75t_SL g691 ( .A(n_692), .Y(n_691) );
INVx1_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
AND2x2_ASAP7_75t_L g697 ( .A(n_698), .B(n_699), .Y(n_697) );
NAND2xp5_ASAP7_75t_L g735 ( .A(n_698), .B(n_706), .Y(n_735) );
INVx1_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
NAND3xp33_ASAP7_75t_L g707 ( .A(n_708), .B(n_709), .C(n_710), .Y(n_707) );
NOR3xp33_ASAP7_75t_L g711 ( .A(n_712), .B(n_736), .C(n_748), .Y(n_711) );
OAI211xp5_ASAP7_75t_SL g712 ( .A1(n_713), .A2(n_714), .B(n_718), .C(n_728), .Y(n_712) );
INVxp67_ASAP7_75t_L g714 ( .A(n_715), .Y(n_714) );
NAND2xp5_ASAP7_75t_SL g715 ( .A(n_716), .B(n_717), .Y(n_715) );
OAI221xp5_ASAP7_75t_L g748 ( .A1(n_717), .A2(n_749), .B1(n_750), .B2(n_751), .C(n_752), .Y(n_748) );
INVx1_ASAP7_75t_L g737 ( .A(n_719), .Y(n_737) );
INVx1_ASAP7_75t_SL g720 ( .A(n_721), .Y(n_720) );
INVx1_ASAP7_75t_L g722 ( .A(n_723), .Y(n_722) );
INVx1_ASAP7_75t_SL g726 ( .A(n_727), .Y(n_726) );
INVx1_ASAP7_75t_L g731 ( .A(n_732), .Y(n_731) );
INVx1_ASAP7_75t_L g734 ( .A(n_735), .Y(n_734) );
INVx1_ASAP7_75t_SL g741 ( .A(n_739), .Y(n_741) );
INVx1_ASAP7_75t_L g742 ( .A(n_743), .Y(n_742) );
CKINVDCx14_ASAP7_75t_R g753 ( .A(n_754), .Y(n_753) );
INVx2_ASAP7_75t_L g756 ( .A(n_757), .Y(n_756) );
INVx1_ASAP7_75t_L g757 ( .A(n_758), .Y(n_757) );
CKINVDCx20_ASAP7_75t_R g759 ( .A(n_760), .Y(n_759) );
INVx1_ASAP7_75t_L g762 ( .A(n_763), .Y(n_762) );
INVx1_ASAP7_75t_SL g768 ( .A(n_769), .Y(n_768) );
INVx3_ASAP7_75t_SL g769 ( .A(n_770), .Y(n_769) );
INVx1_ASAP7_75t_SL g771 ( .A(n_772), .Y(n_771) );
INVx1_ASAP7_75t_L g773 ( .A(n_774), .Y(n_773) );
endmodule