module fake_jpeg_4374_n_106 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_106);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_106;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_3),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_3),
.Y(n_12)
);

CKINVDCx14_ASAP7_75t_R g13 ( 
.A(n_3),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_L g14 ( 
.A(n_5),
.B(n_9),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_10),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

BUFx24_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_5),
.Y(n_21)
);

INVxp67_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

AND2x2_ASAP7_75t_L g24 ( 
.A(n_11),
.B(n_0),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_24),
.B(n_27),
.Y(n_34)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_17),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_25),
.B(n_31),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_20),
.Y(n_26)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_13),
.B(n_23),
.Y(n_27)
);

BUFx2_ASAP7_75t_L g28 ( 
.A(n_17),
.Y(n_28)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_20),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_29),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_17),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_30),
.B(n_31),
.Y(n_36)
);

INVx2_ASAP7_75t_SL g31 ( 
.A(n_17),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_32),
.B(n_12),
.Y(n_41)
);

INVxp67_ASAP7_75t_L g48 ( 
.A(n_33),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_24),
.B(n_16),
.Y(n_39)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_39),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_40),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g55 ( 
.A(n_41),
.B(n_21),
.Y(n_55)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_30),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_42),
.B(n_30),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g43 ( 
.A1(n_37),
.A2(n_15),
.B1(n_29),
.B2(n_26),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_43),
.A2(n_21),
.B1(n_11),
.B2(n_19),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_45),
.B(n_46),
.Y(n_64)
);

HB1xp67_ASAP7_75t_L g46 ( 
.A(n_42),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_41),
.B(n_24),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_47),
.B(n_19),
.Y(n_60)
);

AOI21xp5_ASAP7_75t_L g50 ( 
.A1(n_34),
.A2(n_27),
.B(n_22),
.Y(n_50)
);

AOI21xp5_ASAP7_75t_L g67 ( 
.A1(n_50),
.A2(n_51),
.B(n_14),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g51 ( 
.A(n_34),
.B(n_32),
.C(n_16),
.Y(n_51)
);

O2A1O1Ixp33_ASAP7_75t_L g52 ( 
.A1(n_37),
.A2(n_25),
.B(n_28),
.C(n_31),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_52),
.B(n_54),
.Y(n_65)
);

A2O1A1Ixp33_ASAP7_75t_L g53 ( 
.A1(n_36),
.A2(n_24),
.B(n_22),
.C(n_15),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_53),
.B(n_55),
.Y(n_57)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_35),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_50),
.A2(n_37),
.B1(n_26),
.B2(n_29),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_56),
.A2(n_61),
.B1(n_43),
.B2(n_52),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_55),
.B(n_32),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_58),
.B(n_59),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_55),
.B(n_23),
.Y(n_59)
);

XNOR2xp5_ASAP7_75t_SL g76 ( 
.A(n_60),
.B(n_62),
.Y(n_76)
);

NAND2x1_ASAP7_75t_L g62 ( 
.A(n_47),
.B(n_30),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_48),
.B(n_18),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_63),
.B(n_66),
.Y(n_69)
);

INVxp67_ASAP7_75t_L g66 ( 
.A(n_45),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g73 ( 
.A(n_67),
.B(n_62),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_68),
.A2(n_54),
.B1(n_38),
.B2(n_26),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_60),
.B(n_44),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_70),
.B(n_73),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_62),
.A2(n_44),
.B1(n_53),
.B2(n_51),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_72),
.B(n_74),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_64),
.B(n_49),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_67),
.B(n_61),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_75),
.B(n_77),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g77 ( 
.A(n_65),
.Y(n_77)
);

A2O1A1O1Ixp25_ASAP7_75t_L g79 ( 
.A1(n_76),
.A2(n_57),
.B(n_56),
.C(n_66),
.D(n_36),
.Y(n_79)
);

OAI21xp5_ASAP7_75t_SL g90 ( 
.A1(n_79),
.A2(n_80),
.B(n_0),
.Y(n_90)
);

AOI322xp5_ASAP7_75t_SL g80 ( 
.A1(n_72),
.A2(n_8),
.A3(n_1),
.B1(n_2),
.B2(n_4),
.C1(n_6),
.C2(n_7),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_71),
.B(n_68),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_81),
.B(n_83),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_76),
.B(n_52),
.Y(n_83)
);

AOI221xp5_ASAP7_75t_L g89 ( 
.A1(n_84),
.A2(n_29),
.B1(n_35),
.B2(n_25),
.C(n_49),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_81),
.A2(n_77),
.B1(n_69),
.B2(n_38),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_86),
.B(n_87),
.Y(n_93)
);

AOI21xp5_ASAP7_75t_L g87 ( 
.A1(n_83),
.A2(n_18),
.B(n_49),
.Y(n_87)
);

AO21x1_ASAP7_75t_L g95 ( 
.A1(n_89),
.A2(n_91),
.B(n_28),
.Y(n_95)
);

OAI322xp33_ASAP7_75t_L g92 ( 
.A1(n_90),
.A2(n_85),
.A3(n_82),
.B1(n_78),
.B2(n_6),
.C1(n_7),
.C2(n_0),
.Y(n_92)
);

HB1xp67_ASAP7_75t_L g91 ( 
.A(n_79),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_92),
.B(n_1),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_88),
.A2(n_35),
.B1(n_28),
.B2(n_40),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_94),
.B(n_95),
.Y(n_96)
);

MAJx2_ASAP7_75t_L g97 ( 
.A(n_95),
.B(n_87),
.C(n_86),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_97),
.B(n_93),
.C(n_96),
.Y(n_99)
);

AOI21xp33_ASAP7_75t_L g100 ( 
.A1(n_98),
.A2(n_95),
.B(n_6),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_99),
.B(n_100),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_98),
.B(n_94),
.Y(n_101)
);

AOI21xp5_ASAP7_75t_SL g102 ( 
.A1(n_101),
.A2(n_4),
.B(n_7),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_102),
.B(n_4),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_104),
.B(n_103),
.Y(n_105)
);

NAND2xp33_ASAP7_75t_SL g106 ( 
.A(n_105),
.B(n_40),
.Y(n_106)
);


endmodule