module fake_jpeg_17450_n_317 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_317);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_317;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx12_ASAP7_75t_L g16 ( 
.A(n_12),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_2),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_9),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_4),
.Y(n_21)
);

INVx13_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_0),
.Y(n_23)
);

INVx8_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

BUFx12_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

BUFx8_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_4),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_34),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_35),
.B(n_37),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_20),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_36),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_16),
.B(n_15),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_30),
.Y(n_39)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_20),
.Y(n_40)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_40),
.Y(n_44)
);

OR2x2_ASAP7_75t_L g41 ( 
.A(n_18),
.B(n_0),
.Y(n_41)
);

INVx1_ASAP7_75t_SL g58 ( 
.A(n_41),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_20),
.Y(n_42)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_42),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_16),
.B(n_25),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_43),
.B(n_31),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_39),
.A2(n_27),
.B1(n_24),
.B2(n_32),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_46),
.A2(n_31),
.B1(n_17),
.B2(n_34),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_L g47 ( 
.A1(n_37),
.A2(n_27),
.B1(n_24),
.B2(n_22),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_47),
.A2(n_49),
.B1(n_57),
.B2(n_59),
.Y(n_89)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_38),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_48),
.B(n_61),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_38),
.A2(n_27),
.B1(n_24),
.B2(n_22),
.Y(n_49)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_52),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_53),
.B(n_35),
.Y(n_73)
);

NAND2xp33_ASAP7_75t_SL g54 ( 
.A(n_41),
.B(n_30),
.Y(n_54)
);

XOR2xp5_ASAP7_75t_SL g68 ( 
.A(n_54),
.B(n_41),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_L g57 ( 
.A1(n_35),
.A2(n_24),
.B1(n_22),
.B2(n_21),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_43),
.A2(n_17),
.B1(n_33),
.B2(n_32),
.Y(n_59)
);

INVx5_ASAP7_75t_L g60 ( 
.A(n_36),
.Y(n_60)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_60),
.Y(n_66)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_42),
.Y(n_61)
);

INVx13_ASAP7_75t_L g62 ( 
.A(n_36),
.Y(n_62)
);

INVx8_ASAP7_75t_L g87 ( 
.A(n_62),
.Y(n_87)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_36),
.Y(n_63)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_63),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_58),
.A2(n_22),
.B1(n_32),
.B2(n_33),
.Y(n_64)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_64),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_58),
.A2(n_34),
.B1(n_33),
.B2(n_17),
.Y(n_67)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_67),
.Y(n_120)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_68),
.B(n_85),
.Y(n_98)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_52),
.Y(n_69)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_69),
.Y(n_106)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_55),
.Y(n_71)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_71),
.Y(n_118)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_62),
.Y(n_72)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_72),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_73),
.B(n_91),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_50),
.B(n_41),
.Y(n_74)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_74),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_75),
.A2(n_77),
.B1(n_23),
.B2(n_61),
.Y(n_105)
);

OR2x2_ASAP7_75t_L g76 ( 
.A(n_53),
.B(n_31),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_76),
.B(n_94),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_60),
.A2(n_21),
.B1(n_29),
.B2(n_19),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_50),
.B(n_21),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_78),
.B(n_81),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_55),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_79),
.B(n_82),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_49),
.B(n_30),
.C(n_40),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_80),
.B(n_26),
.C(n_30),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_59),
.B(n_19),
.Y(n_81)
);

BUFx24_ASAP7_75t_SL g82 ( 
.A(n_54),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_48),
.B(n_19),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_83),
.B(n_84),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_48),
.B(n_16),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_62),
.B(n_0),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_51),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_88),
.B(n_97),
.Y(n_117)
);

OA22x2_ASAP7_75t_SL g90 ( 
.A1(n_51),
.A2(n_42),
.B1(n_40),
.B2(n_45),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g115 ( 
.A(n_90),
.B(n_92),
.Y(n_115)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_63),
.Y(n_91)
);

OR2x2_ASAP7_75t_SL g92 ( 
.A(n_44),
.B(n_29),
.Y(n_92)
);

AOI21xp33_ASAP7_75t_L g93 ( 
.A1(n_44),
.A2(n_29),
.B(n_18),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_93),
.B(n_95),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_44),
.B(n_40),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_45),
.B(n_16),
.Y(n_95)
);

OA22x2_ASAP7_75t_L g96 ( 
.A1(n_56),
.A2(n_42),
.B1(n_26),
.B2(n_18),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_96),
.A2(n_23),
.B1(n_56),
.B2(n_2),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_56),
.Y(n_97)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_69),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_99),
.Y(n_127)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_87),
.Y(n_100)
);

INVx11_ASAP7_75t_L g135 ( 
.A(n_100),
.Y(n_135)
);

INVx1_ASAP7_75t_SL g102 ( 
.A(n_85),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_102),
.B(n_116),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g146 ( 
.A(n_105),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_L g107 ( 
.A(n_68),
.B(n_26),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_107),
.B(n_111),
.C(n_122),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_66),
.A2(n_61),
.B1(n_45),
.B2(n_23),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_110),
.A2(n_72),
.B1(n_87),
.B2(n_66),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g111 ( 
.A(n_74),
.B(n_26),
.Y(n_111)
);

AND2x6_ASAP7_75t_L g113 ( 
.A(n_73),
.B(n_89),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_113),
.Y(n_130)
);

INVx13_ASAP7_75t_L g116 ( 
.A(n_87),
.Y(n_116)
);

AOI21xp5_ASAP7_75t_L g141 ( 
.A1(n_121),
.A2(n_125),
.B(n_85),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_78),
.B(n_16),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_123),
.B(n_83),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_89),
.A2(n_20),
.B1(n_10),
.B2(n_15),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_76),
.B(n_30),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_126),
.B(n_76),
.Y(n_129)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_117),
.Y(n_128)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_128),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_129),
.B(n_136),
.Y(n_167)
);

NAND2x1_ASAP7_75t_SL g131 ( 
.A(n_114),
.B(n_64),
.Y(n_131)
);

OAI22x1_ASAP7_75t_L g162 ( 
.A1(n_131),
.A2(n_144),
.B1(n_90),
.B2(n_96),
.Y(n_162)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_99),
.Y(n_132)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_132),
.Y(n_160)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_118),
.Y(n_134)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_134),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_112),
.B(n_73),
.Y(n_136)
);

INVx13_ASAP7_75t_L g137 ( 
.A(n_116),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_137),
.B(n_148),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_138),
.B(n_149),
.Y(n_158)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_118),
.Y(n_139)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_139),
.Y(n_170)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_108),
.Y(n_140)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_140),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_141),
.A2(n_120),
.B1(n_115),
.B2(n_102),
.Y(n_163)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_108),
.Y(n_143)
);

CKINVDCx16_ASAP7_75t_R g173 ( 
.A(n_143),
.Y(n_173)
);

XOR2xp5_ASAP7_75t_L g145 ( 
.A(n_107),
.B(n_80),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_145),
.B(n_122),
.C(n_109),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_112),
.B(n_67),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_147),
.B(n_152),
.Y(n_178)
);

INVxp67_ASAP7_75t_L g148 ( 
.A(n_124),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_100),
.B(n_106),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_106),
.Y(n_150)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_150),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_L g151 ( 
.A1(n_114),
.A2(n_81),
.B(n_92),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_151),
.B(n_96),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_101),
.B(n_94),
.Y(n_152)
);

HB1xp67_ASAP7_75t_L g153 ( 
.A(n_119),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_153),
.Y(n_161)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_121),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_154),
.B(n_155),
.Y(n_175)
);

INVx5_ASAP7_75t_L g155 ( 
.A(n_113),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_125),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_156),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_126),
.B(n_65),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_157),
.B(n_96),
.Y(n_180)
);

OAI21xp33_ASAP7_75t_L g212 ( 
.A1(n_162),
.A2(n_127),
.B(n_140),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_163),
.A2(n_177),
.B1(n_185),
.B2(n_135),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_164),
.B(n_165),
.C(n_169),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_145),
.B(n_142),
.C(n_130),
.Y(n_165)
);

INVxp33_ASAP7_75t_L g168 ( 
.A(n_127),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_168),
.B(n_171),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_142),
.B(n_111),
.C(n_119),
.Y(n_169)
);

AOI32xp33_ASAP7_75t_L g171 ( 
.A1(n_155),
.A2(n_120),
.A3(n_98),
.B1(n_115),
.B2(n_103),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_130),
.B(n_98),
.C(n_70),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_174),
.B(n_183),
.C(n_189),
.Y(n_207)
);

AOI322xp5_ASAP7_75t_L g176 ( 
.A1(n_151),
.A2(n_98),
.A3(n_115),
.B1(n_104),
.B2(n_90),
.C1(n_28),
.C2(n_96),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_176),
.B(n_187),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_154),
.A2(n_90),
.B1(n_70),
.B2(n_91),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_180),
.B(n_152),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_182),
.B(n_150),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g183 ( 
.A(n_157),
.B(n_71),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_141),
.A2(n_146),
.B1(n_156),
.B2(n_147),
.Y(n_185)
);

AO22x1_ASAP7_75t_L g186 ( 
.A1(n_131),
.A2(n_86),
.B1(n_72),
.B2(n_97),
.Y(n_186)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_186),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_134),
.Y(n_187)
);

INVxp67_ASAP7_75t_L g188 ( 
.A(n_133),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_188),
.B(n_132),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_136),
.B(n_86),
.C(n_30),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_129),
.B(n_28),
.Y(n_190)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_190),
.Y(n_195)
);

AOI21xp5_ASAP7_75t_L g191 ( 
.A1(n_175),
.A2(n_146),
.B(n_131),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_191),
.A2(n_210),
.B1(n_212),
.B2(n_186),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_172),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_193),
.B(n_197),
.Y(n_226)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_194),
.Y(n_220)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_159),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_167),
.B(n_148),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_198),
.B(n_200),
.Y(n_227)
);

INVxp67_ASAP7_75t_L g200 ( 
.A(n_159),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_166),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_201),
.B(n_202),
.Y(n_228)
);

OR2x2_ASAP7_75t_L g203 ( 
.A(n_177),
.B(n_128),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_SL g219 ( 
.A(n_203),
.B(n_211),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_160),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g229 ( 
.A1(n_205),
.A2(n_206),
.B1(n_213),
.B2(n_216),
.Y(n_229)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_170),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_167),
.B(n_139),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_SL g232 ( 
.A(n_208),
.B(n_209),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_179),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_179),
.Y(n_213)
);

CKINVDCx16_ASAP7_75t_R g214 ( 
.A(n_184),
.Y(n_214)
);

INVx2_ASAP7_75t_SL g238 ( 
.A(n_214),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_161),
.B(n_137),
.Y(n_215)
);

INVxp67_ASAP7_75t_L g240 ( 
.A(n_215),
.Y(n_240)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_183),
.Y(n_216)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_168),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_217),
.A2(n_135),
.B1(n_143),
.B2(n_173),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_165),
.B(n_127),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_218),
.B(n_164),
.C(n_169),
.Y(n_222)
);

FAx1_ASAP7_75t_SL g221 ( 
.A(n_209),
.B(n_178),
.CI(n_174),
.CON(n_221),
.SN(n_221)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_221),
.B(n_216),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_222),
.B(n_223),
.C(n_225),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_196),
.B(n_189),
.C(n_163),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_192),
.A2(n_181),
.B1(n_180),
.B2(n_162),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_224),
.A2(n_231),
.B1(n_235),
.B2(n_237),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_196),
.B(n_182),
.C(n_178),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_218),
.B(n_190),
.C(n_185),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_230),
.B(n_233),
.C(n_241),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_207),
.B(n_158),
.C(n_186),
.Y(n_233)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_234),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_192),
.A2(n_188),
.B1(n_1),
.B2(n_2),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_191),
.A2(n_28),
.B1(n_1),
.B2(n_3),
.Y(n_236)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_236),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_199),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_L g239 ( 
.A1(n_213),
.A2(n_198),
.B1(n_193),
.B2(n_205),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_239),
.A2(n_195),
.B1(n_208),
.B2(n_201),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_207),
.B(n_26),
.C(n_25),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_242),
.B(n_251),
.Y(n_273)
);

BUFx24_ASAP7_75t_SL g243 ( 
.A(n_221),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_243),
.B(n_244),
.Y(n_264)
);

INVxp67_ASAP7_75t_L g244 ( 
.A(n_226),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_240),
.B(n_206),
.Y(n_247)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_247),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_238),
.B(n_203),
.Y(n_248)
);

CKINVDCx14_ASAP7_75t_R g265 ( 
.A(n_248),
.Y(n_265)
);

NOR2xp67_ASAP7_75t_L g250 ( 
.A(n_221),
.B(n_195),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_SL g263 ( 
.A(n_250),
.B(n_252),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_225),
.B(n_204),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_228),
.Y(n_252)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_253),
.Y(n_261)
);

AOI21xp5_ASAP7_75t_SL g254 ( 
.A1(n_220),
.A2(n_210),
.B(n_194),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_L g270 ( 
.A1(n_254),
.A2(n_257),
.B(n_240),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_222),
.B(n_197),
.C(n_200),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_256),
.B(n_223),
.C(n_233),
.Y(n_262)
);

NAND3xp33_ASAP7_75t_L g257 ( 
.A(n_227),
.B(n_217),
.C(n_4),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_SL g258 ( 
.A(n_232),
.B(n_26),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_258),
.B(n_260),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_SL g260 ( 
.A(n_232),
.B(n_230),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_262),
.B(n_275),
.C(n_255),
.Y(n_278)
);

INVx11_ASAP7_75t_L g266 ( 
.A(n_244),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_266),
.B(n_257),
.Y(n_279)
);

AOI21xp5_ASAP7_75t_L g268 ( 
.A1(n_245),
.A2(n_224),
.B(n_219),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_SL g283 ( 
.A1(n_268),
.A2(n_274),
.B(n_3),
.Y(n_283)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_254),
.Y(n_269)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_269),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_L g280 ( 
.A1(n_270),
.A2(n_258),
.B1(n_260),
.B2(n_6),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_L g271 ( 
.A1(n_259),
.A2(n_229),
.B(n_237),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_271),
.A2(n_269),
.B1(n_274),
.B2(n_261),
.Y(n_287)
);

AOI21xp5_ASAP7_75t_L g274 ( 
.A1(n_246),
.A2(n_235),
.B(n_236),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_255),
.B(n_241),
.C(n_238),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_262),
.B(n_249),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g291 ( 
.A(n_276),
.B(n_287),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_SL g292 ( 
.A(n_278),
.B(n_284),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_279),
.B(n_281),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_280),
.A2(n_261),
.B1(n_264),
.B2(n_272),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g281 ( 
.A(n_263),
.B(n_10),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_265),
.B(n_25),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_282),
.B(n_285),
.Y(n_293)
);

AOI21xp5_ASAP7_75t_L g295 ( 
.A1(n_283),
.A2(n_288),
.B(n_272),
.Y(n_295)
);

NOR2xp67_ASAP7_75t_L g284 ( 
.A(n_270),
.B(n_10),
.Y(n_284)
);

NOR3xp33_ASAP7_75t_SL g285 ( 
.A(n_268),
.B(n_9),
.C(n_5),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_267),
.B(n_25),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_286),
.B(n_266),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_273),
.B(n_25),
.Y(n_288)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_289),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_294),
.B(n_298),
.Y(n_305)
);

OAI21xp5_ASAP7_75t_L g304 ( 
.A1(n_295),
.A2(n_296),
.B(n_7),
.Y(n_304)
);

AOI21xp5_ASAP7_75t_SL g296 ( 
.A1(n_277),
.A2(n_271),
.B(n_273),
.Y(n_296)
);

AOI22xp33_ASAP7_75t_L g297 ( 
.A1(n_283),
.A2(n_275),
.B1(n_3),
.B2(n_7),
.Y(n_297)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_297),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_285),
.B(n_6),
.Y(n_298)
);

NOR2x1_ASAP7_75t_L g299 ( 
.A(n_296),
.B(n_287),
.Y(n_299)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_299),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_291),
.B(n_278),
.C(n_276),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_300),
.B(n_303),
.C(n_299),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_291),
.B(n_292),
.C(n_288),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_302),
.B(n_306),
.Y(n_311)
);

AOI322xp5_ASAP7_75t_L g310 ( 
.A1(n_304),
.A2(n_297),
.A3(n_12),
.B1(n_14),
.B2(n_11),
.C1(n_25),
.C2(n_16),
.Y(n_310)
);

OAI21xp5_ASAP7_75t_SL g306 ( 
.A1(n_293),
.A2(n_7),
.B(n_8),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_301),
.B(n_290),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_307),
.B(n_300),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_309),
.B(n_11),
.C(n_14),
.Y(n_314)
);

NAND3xp33_ASAP7_75t_L g312 ( 
.A(n_310),
.B(n_305),
.C(n_14),
.Y(n_312)
);

OAI311xp33_ASAP7_75t_L g315 ( 
.A1(n_312),
.A2(n_313),
.A3(n_314),
.B1(n_311),
.C1(n_308),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_315),
.B(n_309),
.Y(n_316)
);

XOR2xp5_ASAP7_75t_L g317 ( 
.A(n_316),
.B(n_11),
.Y(n_317)
);


endmodule