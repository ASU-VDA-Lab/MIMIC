module fake_netlist_1_8566_n_17 (n_3, n_1, n_2, n_0, n_17);
input n_3;
input n_1;
input n_2;
input n_0;
output n_17;
wire n_11;
wire n_13;
wire n_16;
wire n_12;
wire n_6;
wire n_4;
wire n_9;
wire n_5;
wire n_14;
wire n_8;
wire n_15;
wire n_10;
wire n_7;
INVx2_ASAP7_75t_L g4 ( .A(n_3), .Y(n_4) );
INVx1_ASAP7_75t_L g5 ( .A(n_2), .Y(n_5) );
AND2x6_ASAP7_75t_L g6 ( .A(n_0), .B(n_1), .Y(n_6) );
BUFx3_ASAP7_75t_L g7 ( .A(n_5), .Y(n_7) );
INVx1_ASAP7_75t_L g8 ( .A(n_4), .Y(n_8) );
BUFx8_ASAP7_75t_L g9 ( .A(n_8), .Y(n_9) );
AND2x2_ASAP7_75t_SL g10 ( .A(n_8), .B(n_6), .Y(n_10) );
NOR2xp33_ASAP7_75t_L g11 ( .A(n_10), .B(n_7), .Y(n_11) );
NAND2xp5_ASAP7_75t_L g12 ( .A(n_11), .B(n_9), .Y(n_12) );
INVx2_ASAP7_75t_L g13 ( .A(n_12), .Y(n_13) );
INVx1_ASAP7_75t_L g14 ( .A(n_13), .Y(n_14) );
BUFx2_ASAP7_75t_L g15 ( .A(n_14), .Y(n_15) );
INVx1_ASAP7_75t_L g16 ( .A(n_15), .Y(n_16) );
INVx1_ASAP7_75t_L g17 ( .A(n_16), .Y(n_17) );
endmodule