module fake_jpeg_19314_n_324 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_324);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_324;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_13;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_145;
wire n_18;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_12;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx4f_ASAP7_75t_L g12 ( 
.A(n_1),
.Y(n_12)
);

CKINVDCx14_ASAP7_75t_R g13 ( 
.A(n_2),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_L g14 ( 
.A(n_2),
.B(n_4),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_8),
.Y(n_15)
);

BUFx10_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_6),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_6),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_0),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_2),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_8),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_25),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_15),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_26),
.B(n_27),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_SL g27 ( 
.A(n_14),
.B(n_19),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_28),
.Y(n_45)
);

INVx2_ASAP7_75t_R g29 ( 
.A(n_13),
.Y(n_29)
);

INVx4_ASAP7_75t_SL g46 ( 
.A(n_29),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_14),
.B(n_6),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_30),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_17),
.Y(n_31)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_31),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_17),
.Y(n_32)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_32),
.Y(n_38)
);

AND2x2_ASAP7_75t_L g33 ( 
.A(n_16),
.B(n_0),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_33),
.B(n_34),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_15),
.Y(n_34)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_32),
.Y(n_37)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_33),
.B(n_12),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_39),
.B(n_33),
.Y(n_63)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_32),
.Y(n_41)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

OAI22xp33_ASAP7_75t_SL g43 ( 
.A1(n_29),
.A2(n_20),
.B1(n_23),
.B2(n_19),
.Y(n_43)
);

OAI22xp33_ASAP7_75t_L g53 ( 
.A1(n_43),
.A2(n_29),
.B1(n_34),
.B2(n_26),
.Y(n_53)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_45),
.Y(n_47)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_47),
.Y(n_85)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_44),
.Y(n_48)
);

INVx2_ASAP7_75t_SL g68 ( 
.A(n_48),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_36),
.B(n_33),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_49),
.B(n_50),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_40),
.B(n_27),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_45),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_51),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_53),
.A2(n_43),
.B1(n_46),
.B2(n_29),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g54 ( 
.A(n_40),
.B(n_27),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_54),
.B(n_55),
.Y(n_82)
);

INVx13_ASAP7_75t_L g55 ( 
.A(n_46),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_45),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_56),
.Y(n_83)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_35),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_57),
.Y(n_67)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_44),
.Y(n_58)
);

BUFx2_ASAP7_75t_L g77 ( 
.A(n_58),
.Y(n_77)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_35),
.Y(n_59)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_59),
.Y(n_73)
);

INVx3_ASAP7_75t_SL g60 ( 
.A(n_44),
.Y(n_60)
);

BUFx2_ASAP7_75t_L g86 ( 
.A(n_60),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_46),
.A2(n_29),
.B1(n_19),
.B2(n_21),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_62),
.A2(n_46),
.B1(n_25),
.B2(n_28),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g66 ( 
.A(n_63),
.B(n_36),
.C(n_39),
.Y(n_66)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_45),
.Y(n_64)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_64),
.Y(n_75)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_37),
.Y(n_65)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_65),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_66),
.B(n_72),
.Y(n_91)
);

CKINVDCx14_ASAP7_75t_R g103 ( 
.A(n_71),
.Y(n_103)
);

AOI21xp5_ASAP7_75t_SL g72 ( 
.A1(n_50),
.A2(n_40),
.B(n_49),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_63),
.A2(n_36),
.B1(n_39),
.B2(n_46),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_74),
.A2(n_80),
.B1(n_33),
.B2(n_28),
.Y(n_108)
);

XNOR2xp5_ASAP7_75t_L g78 ( 
.A(n_49),
.B(n_36),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_78),
.B(n_84),
.Y(n_92)
);

BUFx24_ASAP7_75t_SL g79 ( 
.A(n_54),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_79),
.Y(n_96)
);

MAJx2_ASAP7_75t_L g81 ( 
.A(n_62),
.B(n_39),
.C(n_42),
.Y(n_81)
);

AND2x6_ASAP7_75t_L g88 ( 
.A(n_81),
.B(n_55),
.Y(n_88)
);

XOR2xp5_ASAP7_75t_L g84 ( 
.A(n_47),
.B(n_42),
.Y(n_84)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_67),
.Y(n_87)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_87),
.Y(n_120)
);

XOR2x1_ASAP7_75t_L g114 ( 
.A(n_88),
.B(n_81),
.Y(n_114)
);

BUFx3_ASAP7_75t_L g89 ( 
.A(n_67),
.Y(n_89)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_89),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_68),
.A2(n_52),
.B1(n_61),
.B2(n_65),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_90),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_82),
.B(n_51),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_93),
.B(n_99),
.Y(n_113)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_70),
.Y(n_94)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_94),
.Y(n_112)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_70),
.Y(n_95)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_95),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_L g97 ( 
.A1(n_69),
.A2(n_83),
.B1(n_85),
.B2(n_71),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_97),
.A2(n_75),
.B1(n_44),
.B2(n_60),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_76),
.B(n_42),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_98),
.B(n_55),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_84),
.B(n_64),
.Y(n_99)
);

AND2x2_ASAP7_75t_SL g100 ( 
.A(n_76),
.B(n_56),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_100),
.B(n_101),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_69),
.B(n_26),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_68),
.A2(n_52),
.B1(n_61),
.B2(n_65),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_102),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_73),
.Y(n_104)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_104),
.Y(n_138)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_73),
.Y(n_105)
);

HB1xp67_ASAP7_75t_L g124 ( 
.A(n_105),
.Y(n_124)
);

INVx13_ASAP7_75t_L g106 ( 
.A(n_75),
.Y(n_106)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_106),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_85),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_107),
.B(n_86),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_108),
.A2(n_74),
.B1(n_72),
.B2(n_78),
.Y(n_115)
);

XOR2xp5_ASAP7_75t_L g109 ( 
.A(n_92),
.B(n_66),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_L g143 ( 
.A(n_109),
.B(n_119),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_110),
.B(n_129),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_114),
.A2(n_127),
.B1(n_87),
.B2(n_41),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_115),
.B(n_130),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_91),
.B(n_35),
.C(n_25),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_116),
.B(n_122),
.C(n_100),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_117),
.B(n_131),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g119 ( 
.A(n_92),
.B(n_30),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_103),
.A2(n_60),
.B1(n_44),
.B2(n_25),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_121),
.A2(n_134),
.B1(n_37),
.B2(n_41),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_91),
.B(n_35),
.C(n_32),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_L g127 ( 
.A1(n_88),
.A2(n_34),
.B(n_13),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_88),
.A2(n_60),
.B1(n_35),
.B2(n_41),
.Y(n_129)
);

BUFx24_ASAP7_75t_SL g130 ( 
.A(n_96),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_101),
.Y(n_131)
);

OAI32xp33_ASAP7_75t_L g132 ( 
.A1(n_98),
.A2(n_14),
.A3(n_48),
.B1(n_58),
.B2(n_52),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_132),
.B(n_133),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_108),
.A2(n_37),
.B1(n_41),
.B2(n_58),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_106),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_135),
.B(n_136),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_93),
.Y(n_136)
);

AOI21xp33_ASAP7_75t_SL g137 ( 
.A1(n_99),
.A2(n_77),
.B(n_68),
.Y(n_137)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_137),
.Y(n_142)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_133),
.Y(n_139)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_139),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_114),
.Y(n_144)
);

BUFx2_ASAP7_75t_L g202 ( 
.A(n_144),
.Y(n_202)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_112),
.Y(n_145)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_145),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_146),
.A2(n_37),
.B1(n_38),
.B2(n_31),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_147),
.B(n_159),
.C(n_169),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_113),
.B(n_125),
.Y(n_149)
);

CKINVDCx14_ASAP7_75t_R g176 ( 
.A(n_149),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_113),
.B(n_95),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_150),
.B(n_151),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_115),
.B(n_94),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_118),
.Y(n_152)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_152),
.Y(n_190)
);

INVxp67_ASAP7_75t_L g153 ( 
.A(n_129),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_153),
.B(n_155),
.Y(n_185)
);

AND2x6_ASAP7_75t_L g154 ( 
.A(n_127),
.B(n_100),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_154),
.B(n_162),
.Y(n_175)
);

INVxp67_ASAP7_75t_L g155 ( 
.A(n_116),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_124),
.Y(n_156)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_156),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_123),
.B(n_105),
.Y(n_157)
);

CKINVDCx16_ASAP7_75t_R g183 ( 
.A(n_157),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_109),
.B(n_100),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_158),
.B(n_160),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_122),
.B(n_107),
.C(n_104),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_123),
.B(n_120),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g178 ( 
.A(n_161),
.Y(n_178)
);

HB1xp67_ASAP7_75t_L g162 ( 
.A(n_125),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_119),
.B(n_96),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_165),
.B(n_166),
.Y(n_189)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_138),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_132),
.B(n_104),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_167),
.B(n_168),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_120),
.B(n_89),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_134),
.B(n_48),
.C(n_61),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_128),
.B(n_89),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_170),
.B(n_172),
.Y(n_194)
);

OAI22x1_ASAP7_75t_L g171 ( 
.A1(n_111),
.A2(n_106),
.B1(n_86),
.B2(n_77),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_SL g181 ( 
.A1(n_171),
.A2(n_173),
.B(n_126),
.Y(n_181)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_138),
.Y(n_172)
);

AND2x2_ASAP7_75t_L g173 ( 
.A(n_121),
.B(n_59),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_SL g177 ( 
.A(n_140),
.B(n_21),
.Y(n_177)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_177),
.Y(n_203)
);

NOR4xp25_ASAP7_75t_L g180 ( 
.A(n_154),
.B(n_126),
.C(n_111),
.D(n_24),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_180),
.B(n_22),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_SL g208 ( 
.A1(n_181),
.A2(n_182),
.B(n_184),
.Y(n_208)
);

AOI21xp5_ASAP7_75t_L g182 ( 
.A1(n_142),
.A2(n_9),
.B(n_11),
.Y(n_182)
);

AND2x2_ASAP7_75t_SL g184 ( 
.A(n_164),
.B(n_59),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_163),
.B(n_57),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_187),
.B(n_195),
.Y(n_209)
);

A2O1A1O1Ixp25_ASAP7_75t_L g188 ( 
.A1(n_144),
.A2(n_142),
.B(n_155),
.C(n_153),
.D(n_164),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_SL g219 ( 
.A1(n_188),
.A2(n_13),
.B(n_18),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_143),
.B(n_22),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_192),
.B(n_22),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_193),
.A2(n_169),
.B1(n_146),
.B2(n_173),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_159),
.B(n_57),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_141),
.A2(n_38),
.B1(n_20),
.B2(n_21),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_197),
.A2(n_173),
.B1(n_24),
.B2(n_23),
.Y(n_207)
);

A2O1A1Ixp33_ASAP7_75t_L g198 ( 
.A1(n_141),
.A2(n_24),
.B(n_15),
.C(n_18),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_198),
.B(n_23),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_156),
.B(n_148),
.Y(n_199)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_199),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_200),
.B(n_147),
.C(n_143),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_204),
.B(n_200),
.C(n_196),
.Y(n_229)
);

AOI21xp5_ASAP7_75t_L g205 ( 
.A1(n_175),
.A2(n_171),
.B(n_160),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_205),
.B(n_226),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_206),
.A2(n_212),
.B1(n_186),
.B2(n_190),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_207),
.A2(n_213),
.B1(n_214),
.B2(n_222),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_176),
.B(n_158),
.Y(n_210)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_210),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_211),
.B(n_182),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_191),
.A2(n_38),
.B1(n_20),
.B2(n_31),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_184),
.A2(n_38),
.B1(n_1),
.B2(n_0),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_184),
.A2(n_0),
.B1(n_1),
.B2(n_31),
.Y(n_214)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_215),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_216),
.B(n_218),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_187),
.B(n_12),
.Y(n_217)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_217),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_178),
.B(n_12),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_219),
.B(n_221),
.Y(n_239)
);

HB1xp67_ASAP7_75t_L g221 ( 
.A(n_188),
.Y(n_221)
);

AOI22xp33_ASAP7_75t_L g222 ( 
.A1(n_174),
.A2(n_18),
.B1(n_17),
.B2(n_2),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_185),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_223),
.A2(n_193),
.B1(n_179),
.B2(n_190),
.Y(n_234)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_194),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_224),
.B(n_225),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_178),
.B(n_12),
.Y(n_225)
);

BUFx2_ASAP7_75t_L g226 ( 
.A(n_197),
.Y(n_226)
);

AOI21xp5_ASAP7_75t_L g227 ( 
.A1(n_185),
.A2(n_181),
.B(n_180),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_227),
.B(n_202),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_229),
.B(n_233),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_204),
.B(n_195),
.C(n_196),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_230),
.B(n_238),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_227),
.B(n_192),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_234),
.A2(n_248),
.B1(n_212),
.B2(n_214),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_235),
.B(n_237),
.Y(n_257)
);

XNOR2x1_ASAP7_75t_L g237 ( 
.A(n_208),
.B(n_202),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_209),
.B(n_189),
.C(n_179),
.Y(n_238)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_240),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_241),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_206),
.A2(n_202),
.B1(n_201),
.B2(n_183),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_243),
.B(n_246),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_205),
.B(n_198),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_SL g247 ( 
.A(n_215),
.B(n_177),
.Y(n_247)
);

OA21x2_ASAP7_75t_SL g260 ( 
.A1(n_247),
.A2(n_211),
.B(n_223),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_220),
.A2(n_186),
.B1(n_201),
.B2(n_17),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_208),
.B(n_22),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_249),
.B(n_225),
.Y(n_256)
);

HB1xp67_ASAP7_75t_L g251 ( 
.A(n_238),
.Y(n_251)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_251),
.Y(n_271)
);

A2O1A1O1Ixp25_ASAP7_75t_L g255 ( 
.A1(n_237),
.A2(n_219),
.B(n_209),
.C(n_203),
.D(n_213),
.Y(n_255)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_255),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_256),
.B(n_258),
.Y(n_269)
);

AO21x1_ASAP7_75t_L g258 ( 
.A1(n_239),
.A2(n_216),
.B(n_217),
.Y(n_258)
);

OAI21xp5_ASAP7_75t_L g259 ( 
.A1(n_230),
.A2(n_218),
.B(n_226),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_259),
.A2(n_260),
.B1(n_242),
.B2(n_233),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_SL g261 ( 
.A(n_232),
.B(n_207),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_261),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_262),
.B(n_264),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_244),
.B(n_17),
.Y(n_264)
);

A2O1A1Ixp33_ASAP7_75t_SL g265 ( 
.A1(n_243),
.A2(n_249),
.B(n_245),
.C(n_246),
.Y(n_265)
);

OAI21xp5_ASAP7_75t_SL g279 ( 
.A1(n_265),
.A2(n_1),
.B(n_3),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_236),
.B(n_9),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_266),
.B(n_8),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_SL g282 ( 
.A(n_268),
.B(n_257),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_253),
.A2(n_228),
.B1(n_229),
.B2(n_231),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_272),
.B(n_5),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_252),
.A2(n_247),
.B1(n_235),
.B2(n_4),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_274),
.B(n_276),
.Y(n_281)
);

NOR2xp67_ASAP7_75t_SL g275 ( 
.A(n_251),
.B(n_9),
.Y(n_275)
);

OAI21xp5_ASAP7_75t_L g283 ( 
.A1(n_275),
.A2(n_255),
.B(n_265),
.Y(n_283)
);

AOI21xp5_ASAP7_75t_L g277 ( 
.A1(n_254),
.A2(n_8),
.B(n_3),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_277),
.B(n_278),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_265),
.A2(n_10),
.B1(n_3),
.B2(n_4),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_279),
.B(n_280),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_263),
.B(n_32),
.C(n_12),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g299 ( 
.A(n_282),
.B(n_288),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_283),
.B(n_286),
.Y(n_294)
);

OAI21xp5_ASAP7_75t_L g285 ( 
.A1(n_273),
.A2(n_265),
.B(n_250),
.Y(n_285)
);

AOI21xp5_ASAP7_75t_L g302 ( 
.A1(n_285),
.A2(n_290),
.B(n_5),
.Y(n_302)
);

INVxp67_ASAP7_75t_L g286 ( 
.A(n_272),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_SL g287 ( 
.A(n_270),
.B(n_257),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_287),
.B(n_291),
.Y(n_298)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_280),
.B(n_258),
.Y(n_288)
);

OAI21xp5_ASAP7_75t_SL g290 ( 
.A1(n_271),
.A2(n_32),
.B(n_7),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_SL g291 ( 
.A(n_269),
.B(n_5),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_SL g292 ( 
.A(n_269),
.B(n_268),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_292),
.B(n_278),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_293),
.A2(n_5),
.B1(n_10),
.B2(n_11),
.Y(n_303)
);

OAI21xp5_ASAP7_75t_L g295 ( 
.A1(n_286),
.A2(n_279),
.B(n_277),
.Y(n_295)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_295),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_296),
.B(n_297),
.Y(n_306)
);

AOI21xp5_ASAP7_75t_SL g297 ( 
.A1(n_289),
.A2(n_267),
.B(n_274),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_SL g300 ( 
.A1(n_281),
.A2(n_16),
.B(n_7),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_300),
.B(n_303),
.Y(n_311)
);

OA21x2_ASAP7_75t_SL g301 ( 
.A1(n_282),
.A2(n_284),
.B(n_7),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_301),
.B(n_16),
.C(n_10),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_L g307 ( 
.A(n_302),
.B(n_296),
.Y(n_307)
);

BUFx4f_ASAP7_75t_SL g304 ( 
.A(n_292),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_304),
.B(n_10),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_291),
.B(n_16),
.Y(n_305)
);

INVxp67_ASAP7_75t_L g313 ( 
.A(n_305),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_SL g317 ( 
.A(n_307),
.B(n_308),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_298),
.B(n_16),
.Y(n_308)
);

HB1xp67_ASAP7_75t_L g315 ( 
.A(n_309),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_312),
.B(n_305),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_306),
.B(n_299),
.C(n_294),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_314),
.B(n_316),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_317),
.B(n_304),
.Y(n_319)
);

AO21x2_ASAP7_75t_L g320 ( 
.A1(n_319),
.A2(n_315),
.B(n_310),
.Y(n_320)
);

XOR2xp5_ASAP7_75t_L g321 ( 
.A(n_320),
.B(n_318),
.Y(n_321)
);

AOI21xp5_ASAP7_75t_L g322 ( 
.A1(n_321),
.A2(n_311),
.B(n_313),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_L g323 ( 
.A1(n_322),
.A2(n_313),
.B1(n_16),
.B2(n_11),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_323),
.B(n_16),
.Y(n_324)
);


endmodule