module fake_jpeg_6418_n_77 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_77);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_77;

wire n_10;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_40;
wire n_71;
wire n_30;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_61;
wire n_45;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_11;
wire n_56;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_22;
wire n_35;
wire n_48;
wire n_46;
wire n_9;
wire n_36;
wire n_62;
wire n_43;
wire n_32;

INVx1_ASAP7_75t_L g9 ( 
.A(n_3),
.Y(n_9)
);

INVx1_ASAP7_75t_L g10 ( 
.A(n_7),
.Y(n_10)
);

BUFx4f_ASAP7_75t_L g11 ( 
.A(n_2),
.Y(n_11)
);

INVx6_ASAP7_75t_L g12 ( 
.A(n_6),
.Y(n_12)
);

BUFx16f_ASAP7_75t_L g13 ( 
.A(n_1),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_5),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_4),
.Y(n_15)
);

BUFx3_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

INVx3_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

INVx11_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_18),
.B(n_20),
.Y(n_24)
);

INVx5_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_19),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

AOI21xp33_ASAP7_75t_L g21 ( 
.A1(n_13),
.A2(n_15),
.B(n_14),
.Y(n_21)
);

AOI21xp5_ASAP7_75t_L g30 ( 
.A1(n_21),
.A2(n_23),
.B(n_16),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_22),
.Y(n_28)
);

OAI21xp5_ASAP7_75t_L g23 ( 
.A1(n_15),
.A2(n_14),
.B(n_9),
.Y(n_23)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_19),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_26),
.B(n_22),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_23),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_SL g36 ( 
.A(n_27),
.B(n_12),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_SL g29 ( 
.A1(n_18),
.A2(n_12),
.B1(n_17),
.B2(n_9),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_L g32 ( 
.A1(n_29),
.A2(n_12),
.B1(n_17),
.B2(n_10),
.Y(n_32)
);

XOR2xp5_ASAP7_75t_L g34 ( 
.A(n_30),
.B(n_19),
.Y(n_34)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_24),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_31),
.B(n_28),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g45 ( 
.A1(n_32),
.A2(n_17),
.B1(n_28),
.B2(n_25),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_27),
.B(n_21),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_SL g44 ( 
.A(n_33),
.B(n_35),
.Y(n_44)
);

AOI21xp5_ASAP7_75t_L g47 ( 
.A1(n_34),
.A2(n_11),
.B(n_22),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_30),
.B(n_10),
.Y(n_35)
);

OAI21xp5_ASAP7_75t_L g39 ( 
.A1(n_36),
.A2(n_24),
.B(n_11),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_37),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_25),
.B(n_16),
.Y(n_38)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_38),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_SL g49 ( 
.A(n_39),
.B(n_34),
.Y(n_49)
);

AOI21xp5_ASAP7_75t_L g41 ( 
.A1(n_33),
.A2(n_26),
.B(n_16),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_41),
.A2(n_45),
.B1(n_47),
.B2(n_18),
.Y(n_50)
);

CKINVDCx14_ASAP7_75t_R g54 ( 
.A(n_43),
.Y(n_54)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

INVx13_ASAP7_75t_L g55 ( 
.A(n_46),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_44),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_48),
.B(n_49),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_50),
.A2(n_53),
.B1(n_11),
.B2(n_5),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_41),
.B(n_0),
.Y(n_51)
);

OAI322xp33_ASAP7_75t_L g61 ( 
.A1(n_51),
.A2(n_7),
.A3(n_8),
.B1(n_3),
.B2(n_4),
.C1(n_1),
.C2(n_2),
.Y(n_61)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_45),
.Y(n_52)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_52),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_39),
.A2(n_11),
.B1(n_20),
.B2(n_6),
.Y(n_53)
);

MAJIxp5_ASAP7_75t_L g57 ( 
.A(n_49),
.B(n_42),
.C(n_40),
.Y(n_57)
);

XOR2xp5_ASAP7_75t_L g63 ( 
.A(n_57),
.B(n_60),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_52),
.A2(n_51),
.B1(n_48),
.B2(n_50),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_58),
.A2(n_59),
.B1(n_53),
.B2(n_54),
.Y(n_66)
);

NAND3xp33_ASAP7_75t_L g65 ( 
.A(n_61),
.B(n_8),
.C(n_2),
.Y(n_65)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_60),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_62),
.A2(n_64),
.B1(n_58),
.B2(n_56),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g69 ( 
.A(n_63),
.B(n_55),
.C(n_20),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_57),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_65),
.A2(n_66),
.B1(n_56),
.B2(n_59),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_67),
.B(n_68),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g70 ( 
.A(n_69),
.B(n_55),
.C(n_65),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_70),
.B(n_72),
.Y(n_74)
);

XOR2xp5_ASAP7_75t_L g72 ( 
.A(n_69),
.B(n_55),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_71),
.Y(n_73)
);

OAI21xp5_ASAP7_75t_L g75 ( 
.A1(n_73),
.A2(n_72),
.B(n_3),
.Y(n_75)
);

OAI21xp5_ASAP7_75t_L g76 ( 
.A1(n_75),
.A2(n_74),
.B(n_1),
.Y(n_76)
);

XNOR2xp5_ASAP7_75t_L g77 ( 
.A(n_76),
.B(n_4),
.Y(n_77)
);


endmodule