module real_jpeg_495_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_312;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_L g36 ( 
.A1(n_1),
.A2(n_31),
.B1(n_37),
.B2(n_38),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_1),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_1),
.A2(n_37),
.B1(n_43),
.B2(n_45),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_1),
.A2(n_37),
.B1(n_66),
.B2(n_68),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_1),
.A2(n_37),
.B1(n_59),
.B2(n_60),
.Y(n_317)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_3),
.A2(n_59),
.B1(n_60),
.B2(n_128),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_3),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_SL g178 ( 
.A1(n_3),
.A2(n_66),
.B1(n_68),
.B2(n_128),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_SL g203 ( 
.A1(n_3),
.A2(n_43),
.B1(n_45),
.B2(n_128),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_3),
.A2(n_31),
.B1(n_38),
.B2(n_128),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_4),
.A2(n_59),
.B1(n_60),
.B2(n_162),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_4),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_SL g194 ( 
.A1(n_4),
.A2(n_66),
.B1(n_68),
.B2(n_162),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g232 ( 
.A1(n_4),
.A2(n_43),
.B1(n_45),
.B2(n_162),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_L g265 ( 
.A1(n_4),
.A2(n_31),
.B1(n_38),
.B2(n_162),
.Y(n_265)
);

BUFx5_ASAP7_75t_L g82 ( 
.A(n_5),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g181 ( 
.A1(n_6),
.A2(n_59),
.B1(n_60),
.B2(n_182),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_6),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_SL g193 ( 
.A1(n_6),
.A2(n_66),
.B1(n_68),
.B2(n_182),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_6),
.A2(n_43),
.B1(n_45),
.B2(n_182),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_6),
.A2(n_31),
.B1(n_38),
.B2(n_182),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_L g51 ( 
.A1(n_7),
.A2(n_43),
.B1(n_45),
.B2(n_52),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_7),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_7),
.A2(n_52),
.B1(n_66),
.B2(n_68),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_7),
.A2(n_31),
.B1(n_38),
.B2(n_52),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g309 ( 
.A1(n_7),
.A2(n_52),
.B1(n_59),
.B2(n_60),
.Y(n_309)
);

BUFx8_ASAP7_75t_L g61 ( 
.A(n_8),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_9),
.A2(n_66),
.B1(n_68),
.B2(n_78),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_9),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_9),
.A2(n_59),
.B1(n_60),
.B2(n_78),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_L g120 ( 
.A1(n_9),
.A2(n_43),
.B1(n_45),
.B2(n_78),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_9),
.A2(n_31),
.B1(n_38),
.B2(n_78),
.Y(n_175)
);

BUFx16f_ASAP7_75t_L g48 ( 
.A(n_10),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_11),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_12),
.B(n_59),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_12),
.B(n_163),
.Y(n_197)
);

INVx1_ASAP7_75t_SL g208 ( 
.A(n_12),
.Y(n_208)
);

AOI21xp5_ASAP7_75t_L g219 ( 
.A1(n_12),
.A2(n_59),
.B(n_172),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_12),
.B(n_81),
.Y(n_233)
);

AOI21xp33_ASAP7_75t_L g240 ( 
.A1(n_12),
.A2(n_68),
.B(n_241),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_12),
.B(n_31),
.C(n_48),
.Y(n_249)
);

OAI22xp33_ASAP7_75t_SL g252 ( 
.A1(n_12),
.A2(n_43),
.B1(n_45),
.B2(n_208),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_12),
.B(n_34),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_12),
.B(n_53),
.Y(n_263)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_13),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g41 ( 
.A1(n_14),
.A2(n_42),
.B1(n_43),
.B2(n_45),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_14),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_14),
.A2(n_42),
.B1(n_66),
.B2(n_68),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_14),
.A2(n_42),
.B1(n_59),
.B2(n_60),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_14),
.A2(n_31),
.B1(n_38),
.B2(n_42),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_15),
.A2(n_59),
.B1(n_60),
.B2(n_70),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_15),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_15),
.A2(n_66),
.B1(n_68),
.B2(n_70),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_15),
.A2(n_43),
.B1(n_45),
.B2(n_70),
.Y(n_204)
);

OAI22xp33_ASAP7_75t_SL g212 ( 
.A1(n_15),
.A2(n_31),
.B1(n_38),
.B2(n_70),
.Y(n_212)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_16),
.A2(n_59),
.B1(n_60),
.B2(n_72),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_16),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_16),
.A2(n_66),
.B1(n_68),
.B2(n_72),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_16),
.A2(n_43),
.B1(n_45),
.B2(n_72),
.Y(n_154)
);

OAI22xp33_ASAP7_75t_L g199 ( 
.A1(n_16),
.A2(n_31),
.B1(n_38),
.B2(n_72),
.Y(n_199)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_17),
.Y(n_44)
);

XNOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_314),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

AOI21xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_301),
.B(n_313),
.Y(n_20)
);

AO21x1_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_142),
.B(n_298),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_129),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_SL g23 ( 
.A(n_24),
.B(n_102),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_24),
.B(n_102),
.Y(n_299)
);

XOR2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_73),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_25),
.B(n_88),
.C(n_100),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_54),
.B(n_55),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_26),
.A2(n_27),
.B1(n_105),
.B2(n_106),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_27),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_39),
.Y(n_27)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_28),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_28),
.A2(n_54),
.B1(n_55),
.B2(n_107),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_28),
.A2(n_39),
.B1(n_40),
.B2(n_54),
.Y(n_150)
);

AOI21xp5_ASAP7_75t_L g28 ( 
.A1(n_29),
.A2(n_33),
.B(n_35),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_29),
.A2(n_33),
.B1(n_116),
.B2(n_157),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_29),
.A2(n_33),
.B1(n_211),
.B2(n_213),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_29),
.A2(n_33),
.B1(n_269),
.B2(n_270),
.Y(n_268)
);

INVx1_ASAP7_75t_SL g29 ( 
.A(n_30),
.Y(n_29)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_30),
.A2(n_34),
.B1(n_36),
.B2(n_115),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_30),
.A2(n_34),
.B1(n_175),
.B2(n_176),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_30),
.A2(n_34),
.B1(n_175),
.B2(n_199),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_30),
.A2(n_34),
.B1(n_212),
.B2(n_235),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_30),
.A2(n_34),
.B1(n_208),
.B2(n_261),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_30),
.A2(n_34),
.B1(n_261),
.B2(n_265),
.Y(n_264)
);

AND2x2_ASAP7_75t_L g30 ( 
.A(n_31),
.B(n_33),
.Y(n_30)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_31),
.Y(n_38)
);

OA22x2_ASAP7_75t_L g50 ( 
.A1(n_31),
.A2(n_38),
.B1(n_48),
.B2(n_49),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_31),
.B(n_259),
.Y(n_258)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVxp67_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g40 ( 
.A1(n_41),
.A2(n_46),
.B1(n_51),
.B2(n_53),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_41),
.A2(n_46),
.B1(n_53),
.B2(n_119),
.Y(n_118)
);

INVx4_ASAP7_75t_SL g45 ( 
.A(n_43),
.Y(n_45)
);

OAI22xp33_ASAP7_75t_L g47 ( 
.A1(n_43),
.A2(n_45),
.B1(n_48),
.B2(n_49),
.Y(n_47)
);

AO22x2_ASAP7_75t_SL g81 ( 
.A1(n_43),
.A2(n_45),
.B1(n_82),
.B2(n_83),
.Y(n_81)
);

OAI32xp33_ASAP7_75t_L g206 ( 
.A1(n_43),
.A2(n_68),
.A3(n_82),
.B1(n_207),
.B2(n_209),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_43),
.B(n_249),
.Y(n_248)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g209 ( 
.A(n_45),
.B(n_83),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_46),
.A2(n_51),
.B1(n_53),
.B2(n_87),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_L g94 ( 
.A1(n_46),
.A2(n_53),
.B(n_87),
.Y(n_94)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_46),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_46),
.A2(n_53),
.B1(n_202),
.B2(n_204),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_46),
.A2(n_53),
.B1(n_204),
.B2(n_223),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_46),
.A2(n_53),
.B1(n_231),
.B2(n_232),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_46),
.A2(n_53),
.B1(n_231),
.B2(n_252),
.Y(n_251)
);

AND2x2_ASAP7_75t_L g46 ( 
.A(n_47),
.B(n_50),
.Y(n_46)
);

INVx11_ASAP7_75t_L g49 ( 
.A(n_48),
.Y(n_49)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_50),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_50),
.A2(n_120),
.B1(n_154),
.B2(n_155),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_50),
.A2(n_155),
.B1(n_203),
.B2(n_243),
.Y(n_242)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_55),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_56),
.A2(n_65),
.B1(n_69),
.B2(n_71),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_56),
.A2(n_65),
.B1(n_71),
.B2(n_91),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_56),
.A2(n_65),
.B1(n_69),
.B2(n_126),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_56),
.A2(n_65),
.B1(n_91),
.B2(n_139),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_56),
.A2(n_65),
.B1(n_181),
.B2(n_183),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_56),
.A2(n_65),
.B1(n_181),
.B2(n_219),
.Y(n_218)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_57),
.A2(n_127),
.B1(n_161),
.B2(n_163),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_57),
.A2(n_163),
.B1(n_308),
.B2(n_309),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_SL g316 ( 
.A1(n_57),
.A2(n_163),
.B1(n_309),
.B2(n_317),
.Y(n_316)
);

AND2x2_ASAP7_75t_L g57 ( 
.A(n_58),
.B(n_65),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_59),
.A2(n_60),
.B1(n_62),
.B2(n_64),
.Y(n_58)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

AOI32xp33_ASAP7_75t_L g171 ( 
.A1(n_60),
.A2(n_64),
.A3(n_68),
.B1(n_172),
.B2(n_173),
.Y(n_171)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx6_ASAP7_75t_SL g64 ( 
.A(n_62),
.Y(n_64)
);

OA22x2_ASAP7_75t_L g65 ( 
.A1(n_62),
.A2(n_64),
.B1(n_66),
.B2(n_68),
.Y(n_65)
);

NAND2xp33_ASAP7_75t_SL g173 ( 
.A(n_62),
.B(n_66),
.Y(n_173)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_65),
.Y(n_163)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_66),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_L g84 ( 
.A1(n_66),
.A2(n_68),
.B1(n_82),
.B2(n_83),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_66),
.B(n_208),
.Y(n_207)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_74),
.A2(n_88),
.B1(n_100),
.B2(n_101),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_74),
.Y(n_100)
);

OAI21xp33_ASAP7_75t_L g109 ( 
.A1(n_74),
.A2(n_75),
.B(n_86),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_75),
.B(n_86),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_L g75 ( 
.A1(n_76),
.A2(n_79),
.B1(n_81),
.B2(n_85),
.Y(n_75)
);

INVxp33_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_77),
.A2(n_80),
.B1(n_122),
.B2(n_124),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_79),
.A2(n_81),
.B1(n_85),
.B2(n_97),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_79),
.A2(n_81),
.B1(n_123),
.B2(n_159),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_SL g305 ( 
.A1(n_79),
.A2(n_81),
.B(n_306),
.Y(n_305)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_80),
.A2(n_98),
.B1(n_124),
.B2(n_137),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_80),
.A2(n_124),
.B1(n_178),
.B2(n_179),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_80),
.A2(n_124),
.B1(n_193),
.B2(n_194),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_80),
.A2(n_124),
.B1(n_178),
.B2(n_194),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_80),
.A2(n_124),
.B1(n_193),
.B2(n_240),
.Y(n_239)
);

OR2x2_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_84),
.Y(n_80)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_81),
.Y(n_124)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_82),
.Y(n_83)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_88),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_89),
.A2(n_90),
.B1(n_92),
.B2(n_93),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_89),
.A2(n_90),
.B1(n_132),
.B2(n_133),
.Y(n_131)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_90),
.B(n_94),
.C(n_96),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_90),
.B(n_133),
.C(n_140),
.Y(n_302)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_94),
.A2(n_95),
.B1(n_96),
.B2(n_99),
.Y(n_93)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_94),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_94),
.A2(n_99),
.B1(n_135),
.B2(n_136),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_94),
.B(n_136),
.C(n_138),
.Y(n_312)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_98),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_108),
.C(n_110),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_103),
.A2(n_104),
.B1(n_108),
.B2(n_109),
.Y(n_145)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

XNOR2xp5_ASAP7_75t_L g144 ( 
.A(n_110),
.B(n_145),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_111),
.B(n_121),
.C(n_125),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_111),
.A2(n_112),
.B1(n_148),
.B2(n_149),
.Y(n_147)
);

CKINVDCx16_ASAP7_75t_R g111 ( 
.A(n_112),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_117),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_113),
.A2(n_114),
.B1(n_117),
.B2(n_118),
.Y(n_184)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

XOR2xp5_ASAP7_75t_L g148 ( 
.A(n_121),
.B(n_125),
.Y(n_148)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_L g298 ( 
.A1(n_129),
.A2(n_299),
.B(n_300),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_SL g129 ( 
.A(n_130),
.B(n_141),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_130),
.B(n_141),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_140),
.Y(n_130)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_138),
.Y(n_133)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

CKINVDCx16_ASAP7_75t_R g306 ( 
.A(n_137),
.Y(n_306)
);

CKINVDCx16_ASAP7_75t_R g308 ( 
.A(n_139),
.Y(n_308)
);

AO21x1_ASAP7_75t_L g142 ( 
.A1(n_143),
.A2(n_164),
.B(n_297),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_144),
.B(n_146),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_144),
.B(n_146),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_150),
.C(n_151),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_147),
.B(n_150),
.Y(n_186)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_148),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_151),
.B(n_186),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_158),
.C(n_160),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_152),
.B(n_168),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_153),
.B(n_156),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_153),
.B(n_156),
.Y(n_288)
);

INVxp67_ASAP7_75t_L g223 ( 
.A(n_154),
.Y(n_223)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_157),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_158),
.B(n_160),
.Y(n_168)
);

CKINVDCx14_ASAP7_75t_R g179 ( 
.A(n_159),
.Y(n_179)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_161),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_L g164 ( 
.A1(n_165),
.A2(n_187),
.B(n_296),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_185),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_166),
.B(n_185),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_169),
.C(n_184),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_167),
.B(n_184),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_169),
.B(n_284),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_177),
.C(n_180),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_SL g286 ( 
.A(n_170),
.B(n_287),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_174),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_171),
.B(n_174),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_177),
.B(n_180),
.Y(n_287)
);

AOI31xp33_ASAP7_75t_L g187 ( 
.A1(n_188),
.A2(n_281),
.A3(n_290),
.B(n_293),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_L g188 ( 
.A1(n_189),
.A2(n_226),
.B(n_280),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_214),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_190),
.B(n_214),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_201),
.C(n_205),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g276 ( 
.A(n_191),
.B(n_277),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_195),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_192),
.B(n_196),
.C(n_200),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_196),
.A2(n_197),
.B1(n_198),
.B2(n_200),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_198),
.Y(n_200)
);

INVxp67_ASAP7_75t_L g213 ( 
.A(n_199),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_201),
.B(n_205),
.Y(n_277)
);

INVxp67_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_210),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_206),
.B(n_210),
.Y(n_237)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_207),
.Y(n_241)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

OR2x2_ASAP7_75t_L g290 ( 
.A(n_214),
.B(n_291),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_214),
.B(n_291),
.Y(n_294)
);

FAx1_ASAP7_75t_SL g214 ( 
.A(n_215),
.B(n_216),
.CI(n_217),
.CON(n_214),
.SN(n_214)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_220),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_218),
.B(n_221),
.C(n_225),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_221),
.A2(n_222),
.B1(n_224),
.B2(n_225),
.Y(n_220)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_221),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_222),
.Y(n_225)
);

AOI21xp5_ASAP7_75t_SL g226 ( 
.A1(n_227),
.A2(n_275),
.B(n_279),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_L g227 ( 
.A1(n_228),
.A2(n_244),
.B(n_274),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_236),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_229),
.B(n_236),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_233),
.C(n_234),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_230),
.B(n_233),
.Y(n_254)
);

INVxp67_ASAP7_75t_L g243 ( 
.A(n_232),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_234),
.B(n_254),
.Y(n_253)
);

INVxp67_ASAP7_75t_L g270 ( 
.A(n_235),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_238),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_237),
.B(n_239),
.C(n_242),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_242),
.Y(n_238)
);

AOI21xp5_ASAP7_75t_L g244 ( 
.A1(n_245),
.A2(n_255),
.B(n_273),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_253),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_246),
.B(n_253),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_250),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_247),
.A2(n_248),
.B1(n_250),
.B2(n_251),
.Y(n_271)
);

CKINVDCx16_ASAP7_75t_R g247 ( 
.A(n_248),
.Y(n_247)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

OAI21xp5_ASAP7_75t_L g255 ( 
.A1(n_256),
.A2(n_267),
.B(n_272),
.Y(n_255)
);

AOI21xp5_ASAP7_75t_L g256 ( 
.A1(n_257),
.A2(n_262),
.B(n_266),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_260),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_263),
.B(n_264),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_263),
.B(n_264),
.Y(n_266)
);

INVxp67_ASAP7_75t_L g269 ( 
.A(n_265),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_268),
.B(n_271),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_268),
.B(n_271),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_276),
.B(n_278),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_276),
.B(n_278),
.Y(n_279)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

OAI21xp5_ASAP7_75t_L g293 ( 
.A1(n_282),
.A2(n_294),
.B(n_295),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_SL g282 ( 
.A(n_283),
.B(n_285),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_283),
.B(n_285),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_286),
.B(n_288),
.C(n_289),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_286),
.B(n_292),
.Y(n_291)
);

XOR2xp5_ASAP7_75t_L g292 ( 
.A(n_288),
.B(n_289),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_SL g301 ( 
.A(n_302),
.B(n_303),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_302),
.B(n_303),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_304),
.B(n_312),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_305),
.A2(n_307),
.B1(n_310),
.B2(n_311),
.Y(n_304)
);

CKINVDCx16_ASAP7_75t_R g310 ( 
.A(n_305),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_307),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_307),
.B(n_310),
.C(n_312),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_315),
.B(n_319),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_316),
.B(n_318),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_316),
.Y(n_320)
);

CKINVDCx14_ASAP7_75t_R g321 ( 
.A(n_318),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_320),
.B(n_321),
.Y(n_319)
);


endmodule