module fake_jpeg_14267_n_49 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_49);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_49;

wire n_21;
wire n_33;
wire n_45;
wire n_23;
wire n_27;
wire n_22;
wire n_47;
wire n_40;
wire n_19;
wire n_20;
wire n_18;
wire n_35;
wire n_48;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_32;

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_16),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_12),
.Y(n_20)
);

INVx8_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

INVx5_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_17),
.Y(n_23)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_23),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_19),
.B(n_0),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_SL g33 ( 
.A(n_24),
.B(n_25),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_20),
.B(n_0),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_17),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_26),
.Y(n_28)
);

AOI21xp5_ASAP7_75t_L g27 ( 
.A1(n_22),
.A2(n_7),
.B(n_14),
.Y(n_27)
);

AOI22xp33_ASAP7_75t_SL g31 ( 
.A1(n_27),
.A2(n_21),
.B1(n_22),
.B2(n_18),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_23),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_SL g36 ( 
.A(n_29),
.B(n_31),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_26),
.B(n_21),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_32),
.B(n_26),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_34),
.B(n_35),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_32),
.Y(n_35)
);

OAI21xp5_ASAP7_75t_SL g37 ( 
.A1(n_33),
.A2(n_1),
.B(n_2),
.Y(n_37)
);

XOR2xp5_ASAP7_75t_L g42 ( 
.A(n_37),
.B(n_1),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_L g38 ( 
.A1(n_30),
.A2(n_18),
.B1(n_3),
.B2(n_4),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g39 ( 
.A1(n_38),
.A2(n_36),
.B1(n_30),
.B2(n_28),
.Y(n_39)
);

NAND2xp33_ASAP7_75t_R g45 ( 
.A(n_39),
.B(n_40),
.Y(n_45)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_38),
.Y(n_40)
);

MAJIxp5_ASAP7_75t_L g43 ( 
.A(n_42),
.B(n_3),
.C(n_4),
.Y(n_43)
);

MAJIxp5_ASAP7_75t_L g46 ( 
.A(n_43),
.B(n_44),
.C(n_42),
.Y(n_46)
);

OAI21x1_ASAP7_75t_L g44 ( 
.A1(n_41),
.A2(n_5),
.B(n_6),
.Y(n_44)
);

AOI21xp5_ASAP7_75t_L g47 ( 
.A1(n_46),
.A2(n_45),
.B(n_9),
.Y(n_47)
);

NAND4xp25_ASAP7_75t_L g48 ( 
.A(n_47),
.B(n_10),
.C(n_11),
.D(n_15),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_48),
.B(n_6),
.Y(n_49)
);


endmodule