module fake_jpeg_11445_n_188 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_51, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_52, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_188);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_51;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_52;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_188;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_76;
wire n_127;
wire n_154;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_91;
wire n_93;
wire n_54;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_9),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_32),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_24),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_47),
.Y(n_56)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_50),
.Y(n_57)
);

INVx1_ASAP7_75t_SL g58 ( 
.A(n_8),
.Y(n_58)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_43),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_27),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_5),
.Y(n_61)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_48),
.Y(n_62)
);

BUFx5_ASAP7_75t_L g63 ( 
.A(n_15),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_5),
.Y(n_64)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_0),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_31),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_14),
.Y(n_67)
);

INVx11_ASAP7_75t_L g68 ( 
.A(n_0),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_37),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_15),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_14),
.Y(n_71)
);

BUFx4f_ASAP7_75t_L g72 ( 
.A(n_2),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_9),
.Y(n_73)
);

BUFx12f_ASAP7_75t_L g74 ( 
.A(n_22),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_45),
.Y(n_75)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_44),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_29),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_1),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_51),
.Y(n_79)
);

INVx11_ASAP7_75t_SL g80 ( 
.A(n_52),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_13),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_64),
.B(n_1),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_82),
.B(n_67),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_68),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_83),
.B(n_75),
.Y(n_96)
);

BUFx3_ASAP7_75t_L g84 ( 
.A(n_74),
.Y(n_84)
);

BUFx12f_ASAP7_75t_L g100 ( 
.A(n_84),
.Y(n_100)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_74),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_85),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_77),
.Y(n_86)
);

INVx6_ASAP7_75t_L g92 ( 
.A(n_86),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_77),
.Y(n_87)
);

INVx6_ASAP7_75t_L g98 ( 
.A(n_87),
.Y(n_98)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_72),
.Y(n_88)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_88),
.Y(n_102)
);

INVx8_ASAP7_75t_L g89 ( 
.A(n_63),
.Y(n_89)
);

OR2x2_ASAP7_75t_L g97 ( 
.A(n_89),
.B(n_90),
.Y(n_97)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_72),
.Y(n_90)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_53),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_91),
.B(n_53),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_93),
.B(n_104),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_88),
.A2(n_65),
.B1(n_59),
.B2(n_62),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_95),
.A2(n_71),
.B1(n_76),
.B2(n_57),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_96),
.B(n_103),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_90),
.A2(n_58),
.B1(n_53),
.B2(n_65),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_99),
.A2(n_89),
.B1(n_85),
.B2(n_74),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_86),
.A2(n_71),
.B1(n_59),
.B2(n_87),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_101),
.A2(n_80),
.B1(n_99),
.B2(n_69),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_83),
.B(n_78),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_SL g104 ( 
.A1(n_91),
.A2(n_58),
.B(n_68),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_SL g105 ( 
.A(n_84),
.B(n_73),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_105),
.B(n_54),
.Y(n_110)
);

AND2x2_ASAP7_75t_L g115 ( 
.A(n_106),
.B(n_76),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_107),
.A2(n_120),
.B1(n_128),
.B2(n_28),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_97),
.Y(n_109)
);

HB1xp67_ASAP7_75t_L g139 ( 
.A(n_109),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_110),
.B(n_115),
.Y(n_133)
);

INVx6_ASAP7_75t_L g111 ( 
.A(n_92),
.Y(n_111)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_111),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_105),
.B(n_81),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_112),
.B(n_113),
.Y(n_132)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_94),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_92),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_116),
.B(n_118),
.Y(n_143)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_97),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_117),
.B(n_119),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_102),
.B(n_61),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_102),
.Y(n_119)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_98),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_121),
.B(n_122),
.Y(n_136)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_98),
.Y(n_122)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_94),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_123),
.B(n_124),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_104),
.B(n_70),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_95),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_125),
.B(n_127),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_126),
.A2(n_3),
.B1(n_4),
.B2(n_6),
.Y(n_138)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_100),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_100),
.A2(n_79),
.B1(n_56),
.B2(n_66),
.Y(n_128)
);

AND2x2_ASAP7_75t_L g129 ( 
.A(n_100),
.B(n_55),
.Y(n_129)
);

CKINVDCx16_ASAP7_75t_R g152 ( 
.A(n_129),
.Y(n_152)
);

NAND3xp33_ASAP7_75t_L g130 ( 
.A(n_109),
.B(n_25),
.C(n_49),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_130),
.B(n_144),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_117),
.B(n_60),
.C(n_80),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_SL g162 ( 
.A(n_131),
.B(n_134),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_108),
.B(n_21),
.C(n_42),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_114),
.B(n_2),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_137),
.B(n_13),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_138),
.A2(n_141),
.B1(n_145),
.B2(n_12),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_L g140 ( 
.A1(n_111),
.A2(n_3),
.B1(n_4),
.B2(n_6),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_140),
.A2(n_142),
.B1(n_23),
.B2(n_26),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_116),
.A2(n_7),
.B1(n_8),
.B2(n_10),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_129),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_113),
.A2(n_7),
.B1(n_10),
.B2(n_11),
.Y(n_145)
);

NOR3xp33_ASAP7_75t_SL g146 ( 
.A(n_115),
.B(n_11),
.C(n_12),
.Y(n_146)
);

NOR2xp67_ASAP7_75t_L g164 ( 
.A(n_146),
.B(n_30),
.Y(n_164)
);

A2O1A1O1Ixp25_ASAP7_75t_L g149 ( 
.A1(n_123),
.A2(n_33),
.B(n_41),
.C(n_16),
.D(n_17),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_149),
.B(n_46),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_129),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_151),
.B(n_152),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_153),
.B(n_154),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_155),
.B(n_156),
.Y(n_171)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_136),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_132),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_157),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_139),
.A2(n_150),
.B1(n_148),
.B2(n_142),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_158),
.A2(n_159),
.B1(n_164),
.B2(n_166),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_135),
.A2(n_18),
.B1(n_19),
.B2(n_20),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_160),
.A2(n_167),
.B1(n_168),
.B2(n_140),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_163),
.B(n_165),
.Y(n_174)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_147),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_131),
.B(n_34),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_143),
.A2(n_35),
.B1(n_36),
.B2(n_38),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_134),
.B(n_39),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_SL g173 ( 
.A(n_162),
.B(n_133),
.Y(n_173)
);

OAI322xp33_ASAP7_75t_L g176 ( 
.A1(n_173),
.A2(n_156),
.A3(n_162),
.B1(n_130),
.B2(n_161),
.C1(n_158),
.C2(n_146),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_175),
.B(n_153),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_L g180 ( 
.A1(n_176),
.A2(n_178),
.B(n_179),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_177),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_L g178 ( 
.A1(n_170),
.A2(n_159),
.B(n_149),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_170),
.B(n_167),
.Y(n_179)
);

AND2x2_ASAP7_75t_L g182 ( 
.A(n_180),
.B(n_172),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_182),
.Y(n_183)
);

AOI21xp5_ASAP7_75t_SL g184 ( 
.A1(n_183),
.A2(n_181),
.B(n_174),
.Y(n_184)
);

AOI21xp5_ASAP7_75t_L g185 ( 
.A1(n_184),
.A2(n_171),
.B(n_169),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_185),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_186),
.B(n_173),
.Y(n_187)
);

OR2x2_ASAP7_75t_L g188 ( 
.A(n_187),
.B(n_40),
.Y(n_188)
);


endmodule