module real_aes_13170_n_102 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_102);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_102;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_887;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_838;
wire n_485;
wire n_822;
wire n_846;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_207;
wire n_878;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_900;
wire n_328;
wire n_841;
wire n_318;
wire n_718;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_555;
wire n_421;
wire n_329;
wire n_766;
wire n_852;
wire n_132;
wire n_857;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_571;
wire n_376;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_894;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_865;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_884;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_886;
wire n_594;
wire n_856;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_889;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_870;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_883;
wire n_356;
wire n_478;
wire n_584;
wire n_896;
wire n_408;
wire n_553;
wire n_184;
wire n_578;
wire n_528;
wire n_372;
wire n_202;
wire n_892;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_875;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_559;
wire n_466;
wire n_636;
wire n_872;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_840;
wire n_570;
wire n_675;
wire n_530;
wire n_835;
wire n_104;
wire n_535;
wire n_732;
wire n_834;
wire n_882;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_781;
wire n_860;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_874;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_812;
wire n_817;
wire n_443;
wire n_565;
wire n_782;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_885;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_867;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_879;
wire n_331;
wire n_182;
wire n_417;
wire n_363;
wire n_449;
wire n_754;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_876;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_527;
wire n_505;
wire n_434;
wire n_502;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_552;
wire n_617;
wire n_402;
wire n_733;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_146;
wire n_880;
wire n_807;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_895;
wire n_832;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_869;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_898;
wire n_115;
wire n_604;
wire n_110;
wire n_734;
wire n_848;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_891;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_853;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_851;
wire n_133;
wire n_494;
wire n_711;
wire n_864;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_845;
wire n_850;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_893;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_847;
wire n_779;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_831;
wire n_290;
wire n_365;
wire n_653;
wire n_637;
wire n_526;
wire n_155;
wire n_899;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_866;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_858;
wire n_873;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_266;
wire n_183;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_861;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_839;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_863;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_888;
wire n_836;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_890;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_837;
wire n_871;
wire n_474;
wire n_829;
wire n_170;
wire n_375;
wire n_597;
wire n_640;
wire n_340;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_687;
wire n_729;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_601;
wire n_500;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_854;
wire n_403;
wire n_194;
wire n_137;
wire n_424;
wire n_225;
wire n_877;
wire n_802;
wire n_868;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_842;
wire n_259;
wire n_143;
wire n_849;
wire n_192;
wire n_475;
wire n_554;
wire n_897;
wire n_264;
wire n_855;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
wire n_862;
OA21x2_ASAP7_75t_L g128 ( .A1(n_0), .A2(n_52), .B(n_129), .Y(n_128) );
INVx1_ASAP7_75t_L g245 ( .A(n_0), .Y(n_245) );
OAI22xp5_ASAP7_75t_L g104 ( .A1(n_1), .A2(n_105), .B1(n_106), .B2(n_844), .Y(n_104) );
INVx1_ASAP7_75t_L g844 ( .A(n_1), .Y(n_844) );
NAND2xp5_ASAP7_75t_L g605 ( .A(n_2), .B(n_606), .Y(n_605) );
AND2x2_ASAP7_75t_L g164 ( .A(n_3), .B(n_150), .Y(n_164) );
OAI22xp5_ASAP7_75t_L g862 ( .A1(n_4), .A2(n_863), .B1(n_864), .B2(n_865), .Y(n_862) );
INVxp67_ASAP7_75t_L g863 ( .A(n_4), .Y(n_863) );
NAND2xp33_ASAP7_75t_L g620 ( .A(n_5), .B(n_147), .Y(n_620) );
AOI221xp5_ASAP7_75t_L g291 ( .A1(n_6), .A2(n_99), .B1(n_188), .B2(n_218), .C(n_241), .Y(n_291) );
NAND2xp5_ASAP7_75t_L g157 ( .A(n_7), .B(n_127), .Y(n_157) );
NAND2xp5_ASAP7_75t_L g639 ( .A(n_8), .B(n_578), .Y(n_639) );
NAND2xp5_ASAP7_75t_L g194 ( .A(n_9), .B(n_195), .Y(n_194) );
NAND2xp5_ASAP7_75t_L g132 ( .A(n_10), .B(n_133), .Y(n_132) );
CKINVDCx5p33_ASAP7_75t_R g571 ( .A(n_11), .Y(n_571) );
AOI22xp33_ASAP7_75t_L g102 ( .A1(n_12), .A2(n_103), .B1(n_885), .B2(n_898), .Y(n_102) );
BUFx3_ASAP7_75t_L g138 ( .A(n_13), .Y(n_138) );
INVx1_ASAP7_75t_L g144 ( .A(n_13), .Y(n_144) );
NAND2xp5_ASAP7_75t_L g171 ( .A(n_14), .B(n_172), .Y(n_171) );
A2O1A1Ixp33_ASAP7_75t_L g595 ( .A1(n_15), .A2(n_151), .B(n_532), .C(n_596), .Y(n_595) );
CKINVDCx5p33_ASAP7_75t_R g230 ( .A(n_16), .Y(n_230) );
BUFx10_ASAP7_75t_L g853 ( .A(n_17), .Y(n_853) );
CKINVDCx5p33_ASAP7_75t_R g556 ( .A(n_18), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g643 ( .A(n_19), .B(n_263), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g186 ( .A(n_20), .B(n_187), .Y(n_186) );
NAND2xp5_ASAP7_75t_L g227 ( .A(n_21), .B(n_223), .Y(n_227) );
OAI21xp33_ASAP7_75t_L g324 ( .A1(n_21), .A2(n_69), .B(n_325), .Y(n_324) );
NAND2xp5_ASAP7_75t_L g616 ( .A(n_22), .B(n_261), .Y(n_616) );
A2O1A1Ixp33_ASAP7_75t_L g586 ( .A1(n_23), .A2(n_587), .B(n_588), .C(n_590), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_24), .B(n_543), .Y(n_542) );
O2A1O1Ixp5_ASAP7_75t_L g292 ( .A1(n_25), .A2(n_152), .B(n_198), .C(n_293), .Y(n_292) );
AND2x2_ASAP7_75t_L g553 ( .A(n_26), .B(n_127), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g644 ( .A(n_27), .B(n_223), .Y(n_644) );
AOI22xp5_ASAP7_75t_L g865 ( .A1(n_28), .A2(n_32), .B1(n_109), .B2(n_866), .Y(n_865) );
CKINVDCx5p33_ASAP7_75t_R g866 ( .A(n_28), .Y(n_866) );
AOI22xp33_ASAP7_75t_L g580 ( .A1(n_29), .A2(n_80), .B1(n_195), .B2(n_211), .Y(n_580) );
INVx1_ASAP7_75t_L g156 ( .A(n_30), .Y(n_156) );
INVx1_ASAP7_75t_L g609 ( .A(n_31), .Y(n_609) );
INVx1_ASAP7_75t_L g109 ( .A(n_32), .Y(n_109) );
NOR2xp33_ASAP7_75t_L g233 ( .A(n_33), .B(n_148), .Y(n_233) );
NAND2xp5_ASAP7_75t_SL g638 ( .A(n_34), .B(n_211), .Y(n_638) );
NAND2xp5_ASAP7_75t_L g621 ( .A(n_35), .B(n_223), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g184 ( .A(n_36), .B(n_185), .Y(n_184) );
INVx1_ASAP7_75t_L g115 ( .A(n_37), .Y(n_115) );
AND3x2_ASAP7_75t_L g880 ( .A(n_37), .B(n_848), .C(n_850), .Y(n_880) );
NAND2xp5_ASAP7_75t_SL g541 ( .A(n_38), .B(n_188), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_39), .B(n_223), .Y(n_533) );
NAND2xp5_ASAP7_75t_SL g559 ( .A(n_40), .B(n_198), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g283 ( .A(n_41), .B(n_172), .Y(n_283) );
CKINVDCx5p33_ASAP7_75t_R g597 ( .A(n_42), .Y(n_597) );
AND2x4_ASAP7_75t_L g155 ( .A(n_43), .B(n_156), .Y(n_155) );
NAND2x1_ASAP7_75t_L g149 ( .A(n_44), .B(n_150), .Y(n_149) );
CKINVDCx5p33_ASAP7_75t_R g237 ( .A(n_45), .Y(n_237) );
AOI22x1_ASAP7_75t_L g106 ( .A1(n_46), .A2(n_107), .B1(n_842), .B2(n_843), .Y(n_106) );
INVx1_ASAP7_75t_L g843 ( .A(n_46), .Y(n_843) );
INVx1_ASAP7_75t_L g141 ( .A(n_47), .Y(n_141) );
CKINVDCx5p33_ASAP7_75t_R g255 ( .A(n_48), .Y(n_255) );
AND2x2_ASAP7_75t_L g162 ( .A(n_49), .B(n_163), .Y(n_162) );
NAND2xp5_ASAP7_75t_L g210 ( .A(n_50), .B(n_211), .Y(n_210) );
AOI22xp33_ASAP7_75t_L g577 ( .A1(n_51), .A2(n_94), .B1(n_211), .B2(n_578), .Y(n_577) );
INVx1_ASAP7_75t_L g246 ( .A(n_52), .Y(n_246) );
NAND2xp5_ASAP7_75t_L g265 ( .A(n_53), .B(n_127), .Y(n_265) );
INVx1_ASAP7_75t_L g129 ( .A(n_54), .Y(n_129) );
NAND2xp5_ASAP7_75t_SL g170 ( .A(n_55), .B(n_163), .Y(n_170) );
AND2x4_ASAP7_75t_L g890 ( .A(n_56), .B(n_891), .Y(n_890) );
NAND2xp5_ASAP7_75t_L g222 ( .A(n_57), .B(n_223), .Y(n_222) );
NAND2xp5_ASAP7_75t_L g146 ( .A(n_58), .B(n_147), .Y(n_146) );
NOR2xp67_ASAP7_75t_L g849 ( .A(n_59), .B(n_84), .Y(n_849) );
HB1xp67_ASAP7_75t_L g894 ( .A(n_59), .Y(n_894) );
NAND2xp5_ASAP7_75t_SL g280 ( .A(n_60), .B(n_211), .Y(n_280) );
AND2x2_ASAP7_75t_L g548 ( .A(n_61), .B(n_180), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g259 ( .A(n_62), .B(n_260), .Y(n_259) );
NAND2xp5_ASAP7_75t_L g560 ( .A(n_63), .B(n_543), .Y(n_560) );
INVx1_ASAP7_75t_L g891 ( .A(n_64), .Y(n_891) );
NAND2x1_ASAP7_75t_L g531 ( .A(n_65), .B(n_532), .Y(n_531) );
AND2x2_ASAP7_75t_L g168 ( .A(n_66), .B(n_127), .Y(n_168) );
NAND2xp5_ASAP7_75t_L g619 ( .A(n_67), .B(n_172), .Y(n_619) );
CKINVDCx5p33_ASAP7_75t_R g882 ( .A(n_68), .Y(n_882) );
CKINVDCx5p33_ASAP7_75t_R g297 ( .A(n_69), .Y(n_297) );
NAND2xp5_ASAP7_75t_SL g197 ( .A(n_70), .B(n_198), .Y(n_197) );
NAND2xp5_ASAP7_75t_L g279 ( .A(n_71), .B(n_195), .Y(n_279) );
NAND2xp5_ASAP7_75t_L g257 ( .A(n_72), .B(n_211), .Y(n_257) );
CKINVDCx5p33_ASAP7_75t_R g294 ( .A(n_73), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_74), .B(n_252), .Y(n_602) );
NAND2xp5_ASAP7_75t_SL g641 ( .A(n_75), .B(n_642), .Y(n_641) );
INVx2_ASAP7_75t_L g851 ( .A(n_76), .Y(n_851) );
HB1xp67_ASAP7_75t_L g897 ( .A(n_76), .Y(n_897) );
NAND2xp5_ASAP7_75t_SL g527 ( .A(n_77), .B(n_185), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g592 ( .A(n_78), .B(n_593), .Y(n_592) );
AOI21xp5_ASAP7_75t_SL g875 ( .A1(n_79), .A2(n_876), .B(n_881), .Y(n_875) );
NAND2xp5_ASAP7_75t_SL g216 ( .A(n_81), .B(n_217), .Y(n_216) );
NAND2xp5_ASAP7_75t_SL g547 ( .A(n_82), .B(n_188), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g285 ( .A(n_83), .B(n_223), .Y(n_285) );
HB1xp67_ASAP7_75t_L g896 ( .A(n_84), .Y(n_896) );
NAND2xp5_ASAP7_75t_L g179 ( .A(n_85), .B(n_180), .Y(n_179) );
NAND2xp5_ASAP7_75t_SL g282 ( .A(n_86), .B(n_163), .Y(n_282) );
CKINVDCx5p33_ASAP7_75t_R g530 ( .A(n_87), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g528 ( .A(n_88), .B(n_263), .Y(n_528) );
NAND2xp33_ASAP7_75t_SL g604 ( .A(n_89), .B(n_236), .Y(n_604) );
CKINVDCx5p33_ASAP7_75t_R g239 ( .A(n_90), .Y(n_239) );
NAND2xp5_ASAP7_75t_SL g601 ( .A(n_91), .B(n_163), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g219 ( .A(n_92), .B(n_187), .Y(n_219) );
NAND2xp5_ASAP7_75t_L g212 ( .A(n_93), .B(n_213), .Y(n_212) );
BUFx3_ASAP7_75t_L g134 ( .A(n_95), .Y(n_134) );
INVx1_ASAP7_75t_L g153 ( .A(n_95), .Y(n_153) );
INVx1_ASAP7_75t_L g192 ( .A(n_95), .Y(n_192) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_96), .B(n_238), .Y(n_546) );
CKINVDCx5p33_ASAP7_75t_R g589 ( .A(n_97), .Y(n_589) );
NAND2xp33_ASAP7_75t_L g617 ( .A(n_98), .B(n_142), .Y(n_617) );
NAND2xp5_ASAP7_75t_L g262 ( .A(n_100), .B(n_263), .Y(n_262) );
NAND2xp5_ASAP7_75t_SL g557 ( .A(n_101), .B(n_163), .Y(n_557) );
AO21x2_ASAP7_75t_L g103 ( .A1(n_104), .A2(n_845), .B(n_854), .Y(n_103) );
INVx1_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
INVx1_ASAP7_75t_L g842 ( .A(n_107), .Y(n_842) );
OA21x2_ASAP7_75t_L g107 ( .A1(n_108), .A2(n_116), .B(n_515), .Y(n_107) );
NAND2xp5_ASAP7_75t_L g108 ( .A(n_109), .B(n_110), .Y(n_108) );
NOR2xp33_ASAP7_75t_L g841 ( .A(n_109), .B(n_112), .Y(n_841) );
INVxp67_ASAP7_75t_SL g110 ( .A(n_111), .Y(n_110) );
BUFx8_ASAP7_75t_L g111 ( .A(n_112), .Y(n_111) );
AOI22xp5_ASAP7_75t_L g515 ( .A1(n_112), .A2(n_116), .B1(n_516), .B2(n_841), .Y(n_515) );
BUFx6f_ASAP7_75t_SL g112 ( .A(n_113), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_114), .Y(n_113) );
AND2x4_ASAP7_75t_L g887 ( .A(n_114), .B(n_888), .Y(n_887) );
BUFx2_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
NAND2xp5_ASAP7_75t_L g874 ( .A(n_115), .B(n_849), .Y(n_874) );
XNOR2xp5_ASAP7_75t_L g861 ( .A(n_116), .B(n_862), .Y(n_861) );
AND2x2_ASAP7_75t_L g116 ( .A(n_117), .B(n_450), .Y(n_116) );
NOR4xp25_ASAP7_75t_L g117 ( .A(n_118), .B(n_338), .C(n_391), .D(n_432), .Y(n_117) );
NAND2xp5_ASAP7_75t_L g118 ( .A(n_119), .B(n_312), .Y(n_118) );
AOI21xp5_ASAP7_75t_L g119 ( .A1(n_120), .A2(n_201), .B(n_266), .Y(n_119) );
AOI22xp5_ASAP7_75t_L g416 ( .A1(n_120), .A2(n_370), .B1(n_417), .B2(n_419), .Y(n_416) );
AND2x2_ASAP7_75t_L g120 ( .A(n_121), .B(n_158), .Y(n_120) );
HB1xp67_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
NAND2xp5_ASAP7_75t_L g445 ( .A(n_122), .B(n_160), .Y(n_445) );
INVx1_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
INVx2_ASAP7_75t_L g310 ( .A(n_123), .Y(n_310) );
AND2x2_ASAP7_75t_L g319 ( .A(n_123), .B(n_311), .Y(n_319) );
AND2x2_ASAP7_75t_L g345 ( .A(n_123), .B(n_272), .Y(n_345) );
NAND2xp5_ASAP7_75t_L g353 ( .A(n_123), .B(n_160), .Y(n_353) );
INVxp67_ASAP7_75t_L g361 ( .A(n_123), .Y(n_361) );
AND2x4_ASAP7_75t_SL g377 ( .A(n_123), .B(n_303), .Y(n_377) );
HB1xp67_ASAP7_75t_L g397 ( .A(n_123), .Y(n_397) );
INVx1_ASAP7_75t_L g413 ( .A(n_123), .Y(n_413) );
BUFx6f_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
OAI21x1_ASAP7_75t_L g124 ( .A1(n_125), .A2(n_130), .B(n_157), .Y(n_124) );
INVx1_ASAP7_75t_SL g125 ( .A(n_126), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
INVxp33_ASAP7_75t_L g175 ( .A(n_127), .Y(n_175) );
BUFx6f_ASAP7_75t_L g207 ( .A(n_127), .Y(n_207) );
INVx1_ASAP7_75t_L g298 ( .A(n_127), .Y(n_298) );
NOR2xp67_ASAP7_75t_SL g539 ( .A(n_127), .B(n_243), .Y(n_539) );
INVxp67_ASAP7_75t_SL g552 ( .A(n_127), .Y(n_552) );
BUFx6f_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
INVx1_ASAP7_75t_L g181 ( .A(n_128), .Y(n_181) );
BUFx2_ASAP7_75t_L g276 ( .A(n_128), .Y(n_276) );
INVxp33_ASAP7_75t_L g610 ( .A(n_128), .Y(n_610) );
INVx1_ASAP7_75t_L g247 ( .A(n_129), .Y(n_247) );
OAI21x1_ASAP7_75t_L g130 ( .A1(n_131), .A2(n_145), .B(n_154), .Y(n_130) );
OAI21xp5_ASAP7_75t_L g131 ( .A1(n_132), .A2(n_135), .B(n_139), .Y(n_131) );
INVx1_ASAP7_75t_L g590 ( .A(n_133), .Y(n_590) );
INVx2_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
NOR2xp33_ASAP7_75t_L g140 ( .A(n_134), .B(n_141), .Y(n_140) );
INVx1_ASAP7_75t_L g234 ( .A(n_134), .Y(n_234) );
INVx2_ASAP7_75t_L g284 ( .A(n_134), .Y(n_284) );
AOI211x1_ASAP7_75t_L g554 ( .A1(n_134), .A2(n_553), .B(n_555), .C(n_558), .Y(n_554) );
INVx1_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
INVx3_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
INVx3_ASAP7_75t_L g150 ( .A(n_137), .Y(n_150) );
INVx2_ASAP7_75t_L g172 ( .A(n_137), .Y(n_172) );
INVx2_ASAP7_75t_L g543 ( .A(n_137), .Y(n_543) );
INVx2_ASAP7_75t_L g578 ( .A(n_137), .Y(n_578) );
INVx2_ASAP7_75t_L g606 ( .A(n_137), .Y(n_606) );
BUFx6f_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
INVx2_ASAP7_75t_L g148 ( .A(n_138), .Y(n_148) );
BUFx6f_ASAP7_75t_L g196 ( .A(n_138), .Y(n_196) );
NAND2xp5_ASAP7_75t_L g139 ( .A(n_140), .B(n_142), .Y(n_139) );
INVx1_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
INVx2_ASAP7_75t_L g163 ( .A(n_143), .Y(n_163) );
INVx2_ASAP7_75t_L g198 ( .A(n_143), .Y(n_198) );
INVx2_ASAP7_75t_L g236 ( .A(n_143), .Y(n_236) );
BUFx6f_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
INVx2_ASAP7_75t_L g189 ( .A(n_144), .Y(n_189) );
AOI21x1_ASAP7_75t_L g145 ( .A1(n_146), .A2(n_149), .B(n_151), .Y(n_145) );
INVx1_ASAP7_75t_L g213 ( .A(n_147), .Y(n_213) );
INVx2_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
INVx1_ASAP7_75t_L g185 ( .A(n_148), .Y(n_185) );
INVx2_ASAP7_75t_L g211 ( .A(n_148), .Y(n_211) );
INVx2_ASAP7_75t_L g232 ( .A(n_148), .Y(n_232) );
AOI21xp5_ASAP7_75t_L g193 ( .A1(n_151), .A2(n_194), .B(n_197), .Y(n_193) );
INVx2_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
INVx2_ASAP7_75t_L g214 ( .A(n_152), .Y(n_214) );
INVx2_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
BUFx3_ASAP7_75t_L g166 ( .A(n_153), .Y(n_166) );
INVx1_ASAP7_75t_L g200 ( .A(n_154), .Y(n_200) );
OAI21xp5_ASAP7_75t_L g277 ( .A1(n_154), .A2(n_278), .B(n_281), .Y(n_277) );
AOI21xp5_ASAP7_75t_L g551 ( .A1(n_154), .A2(n_552), .B(n_553), .Y(n_551) );
AOI21xp5_ASAP7_75t_L g611 ( .A1(n_154), .A2(n_275), .B(n_608), .Y(n_611) );
OAI21x1_ASAP7_75t_L g614 ( .A1(n_154), .A2(n_615), .B(n_618), .Y(n_614) );
OAI21x1_ASAP7_75t_L g636 ( .A1(n_154), .A2(n_637), .B(n_640), .Y(n_636) );
BUFx6f_ASAP7_75t_SL g154 ( .A(n_155), .Y(n_154) );
INVx3_ASAP7_75t_L g177 ( .A(n_155), .Y(n_177) );
INVx2_ASAP7_75t_L g221 ( .A(n_155), .Y(n_221) );
INVx1_ASAP7_75t_L g243 ( .A(n_155), .Y(n_243) );
INVx1_ASAP7_75t_L g575 ( .A(n_155), .Y(n_575) );
INVx2_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
INVx2_ASAP7_75t_L g315 ( .A(n_159), .Y(n_315) );
INVxp67_ASAP7_75t_L g427 ( .A(n_159), .Y(n_427) );
OR2x2_ASAP7_75t_L g159 ( .A(n_160), .B(n_178), .Y(n_159) );
INVx2_ASAP7_75t_L g303 ( .A(n_160), .Y(n_303) );
AND2x2_ASAP7_75t_L g398 ( .A(n_160), .B(n_337), .Y(n_398) );
INVx1_ASAP7_75t_L g406 ( .A(n_160), .Y(n_406) );
AO21x2_ASAP7_75t_L g160 ( .A1(n_161), .A2(n_167), .B(n_174), .Y(n_160) );
OAI21xp5_ASAP7_75t_L g161 ( .A1(n_162), .A2(n_164), .B(n_165), .Y(n_161) );
INVx1_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
INVx2_ASAP7_75t_L g173 ( .A(n_166), .Y(n_173) );
O2A1O1Ixp5_ASAP7_75t_L g529 ( .A1(n_166), .A2(n_251), .B(n_530), .C(n_531), .Y(n_529) );
NAND3xp33_ASAP7_75t_L g579 ( .A(n_166), .B(n_328), .C(n_574), .Y(n_579) );
NOR2xp67_ASAP7_75t_L g167 ( .A(n_168), .B(n_169), .Y(n_167) );
AOI21xp33_ASAP7_75t_L g174 ( .A1(n_168), .A2(n_175), .B(n_176), .Y(n_174) );
AOI21xp5_ASAP7_75t_L g169 ( .A1(n_170), .A2(n_171), .B(n_173), .Y(n_169) );
AOI21xp5_ASAP7_75t_L g540 ( .A1(n_173), .A2(n_541), .B(n_542), .Y(n_540) );
INVx2_ASAP7_75t_L g176 ( .A(n_177), .Y(n_176) );
NOR3xp33_ASAP7_75t_L g290 ( .A(n_177), .B(n_291), .C(n_292), .Y(n_290) );
AND2x2_ASAP7_75t_L g302 ( .A(n_178), .B(n_303), .Y(n_302) );
INVx3_ASAP7_75t_L g337 ( .A(n_178), .Y(n_337) );
INVx1_ASAP7_75t_L g344 ( .A(n_178), .Y(n_344) );
AND2x2_ASAP7_75t_L g360 ( .A(n_178), .B(n_361), .Y(n_360) );
INVx1_ASAP7_75t_L g366 ( .A(n_178), .Y(n_366) );
HB1xp67_ASAP7_75t_L g394 ( .A(n_178), .Y(n_394) );
AND2x2_ASAP7_75t_L g453 ( .A(n_178), .B(n_369), .Y(n_453) );
AND2x4_ASAP7_75t_L g178 ( .A(n_179), .B(n_182), .Y(n_178) );
NOR2xp33_ASAP7_75t_L g199 ( .A(n_180), .B(n_200), .Y(n_199) );
BUFx6f_ASAP7_75t_L g223 ( .A(n_180), .Y(n_223) );
INVx2_ASAP7_75t_L g180 ( .A(n_181), .Y(n_180) );
OAI21xp5_ASAP7_75t_L g182 ( .A1(n_183), .A2(n_193), .B(n_199), .Y(n_182) );
AOI21xp5_ASAP7_75t_L g183 ( .A1(n_184), .A2(n_186), .B(n_190), .Y(n_183) );
INVx2_ASAP7_75t_L g187 ( .A(n_188), .Y(n_187) );
INVx1_ASAP7_75t_L g587 ( .A(n_188), .Y(n_587) );
NOR2xp33_ASAP7_75t_L g596 ( .A(n_188), .B(n_597), .Y(n_596) );
BUFx6f_ASAP7_75t_L g188 ( .A(n_189), .Y(n_188) );
INVx3_ASAP7_75t_L g218 ( .A(n_189), .Y(n_218) );
AOI21xp5_ASAP7_75t_L g215 ( .A1(n_190), .A2(n_216), .B(n_219), .Y(n_215) );
AOI21xp5_ASAP7_75t_L g258 ( .A1(n_190), .A2(n_259), .B(n_262), .Y(n_258) );
AOI21xp5_ASAP7_75t_L g278 ( .A1(n_190), .A2(n_279), .B(n_280), .Y(n_278) );
AOI21xp5_ASAP7_75t_L g526 ( .A1(n_190), .A2(n_527), .B(n_528), .Y(n_526) );
AOI21xp5_ASAP7_75t_L g558 ( .A1(n_190), .A2(n_559), .B(n_560), .Y(n_558) );
AO21x1_ASAP7_75t_L g600 ( .A1(n_190), .A2(n_601), .B(n_602), .Y(n_600) );
AOI21xp5_ASAP7_75t_L g640 ( .A1(n_190), .A2(n_641), .B(n_643), .Y(n_640) );
BUFx10_ASAP7_75t_L g190 ( .A(n_191), .Y(n_190) );
INVx1_ASAP7_75t_L g191 ( .A(n_192), .Y(n_191) );
BUFx3_ASAP7_75t_L g241 ( .A(n_192), .Y(n_241) );
INVx2_ASAP7_75t_L g195 ( .A(n_196), .Y(n_195) );
INVx2_ASAP7_75t_L g238 ( .A(n_196), .Y(n_238) );
INVx1_ASAP7_75t_L g252 ( .A(n_196), .Y(n_252) );
INVx2_ASAP7_75t_L g261 ( .A(n_196), .Y(n_261) );
NAND2xp5_ASAP7_75t_SL g293 ( .A(n_196), .B(n_294), .Y(n_293) );
AOI22xp33_ASAP7_75t_L g457 ( .A1(n_201), .A2(n_424), .B1(n_458), .B2(n_460), .Y(n_457) );
AND2x2_ASAP7_75t_L g201 ( .A(n_202), .B(n_224), .Y(n_201) );
OR2x2_ASAP7_75t_L g321 ( .A(n_202), .B(n_322), .Y(n_321) );
AND2x2_ASAP7_75t_L g456 ( .A(n_202), .B(n_415), .Y(n_456) );
INVx2_ASAP7_75t_L g202 ( .A(n_203), .Y(n_202) );
INVx1_ASAP7_75t_L g203 ( .A(n_204), .Y(n_203) );
AND2x2_ASAP7_75t_L g342 ( .A(n_204), .B(n_307), .Y(n_342) );
INVx1_ASAP7_75t_L g204 ( .A(n_205), .Y(n_204) );
AND2x2_ASAP7_75t_L g379 ( .A(n_205), .B(n_289), .Y(n_379) );
OAI21xp5_ASAP7_75t_L g205 ( .A1(n_206), .A2(n_208), .B(n_222), .Y(n_205) );
OAI21x1_ASAP7_75t_L g248 ( .A1(n_206), .A2(n_249), .B(n_265), .Y(n_248) );
OAI21x1_ASAP7_75t_L g300 ( .A1(n_206), .A2(n_208), .B(n_222), .Y(n_300) );
OAI21x1_ASAP7_75t_L g330 ( .A1(n_206), .A2(n_249), .B(n_265), .Y(n_330) );
OAI21x1_ASAP7_75t_L g524 ( .A1(n_206), .A2(n_525), .B(n_533), .Y(n_524) );
OAI21xp5_ASAP7_75t_L g635 ( .A1(n_206), .A2(n_636), .B(n_644), .Y(n_635) );
OAI21x1_ASAP7_75t_L g661 ( .A1(n_206), .A2(n_636), .B(n_644), .Y(n_661) );
BUFx6f_ASAP7_75t_L g206 ( .A(n_207), .Y(n_206) );
OAI21x1_ASAP7_75t_L g208 ( .A1(n_209), .A2(n_215), .B(n_220), .Y(n_208) );
AOI21xp5_ASAP7_75t_L g209 ( .A1(n_210), .A2(n_212), .B(n_214), .Y(n_209) );
INVx1_ASAP7_75t_L g576 ( .A(n_214), .Y(n_576) );
OAI21xp5_ASAP7_75t_L g555 ( .A1(n_217), .A2(n_556), .B(n_557), .Y(n_555) );
INVx2_ASAP7_75t_L g217 ( .A(n_218), .Y(n_217) );
INVx2_ASAP7_75t_L g532 ( .A(n_218), .Y(n_532) );
NOR2xp33_ASAP7_75t_L g588 ( .A(n_218), .B(n_589), .Y(n_588) );
INVx2_ASAP7_75t_L g642 ( .A(n_218), .Y(n_642) );
OAI21xp5_ASAP7_75t_L g525 ( .A1(n_220), .A2(n_526), .B(n_529), .Y(n_525) );
INVx1_ASAP7_75t_L g220 ( .A(n_221), .Y(n_220) );
INVx2_ASAP7_75t_SL g264 ( .A(n_221), .Y(n_264) );
AND2x4_ASAP7_75t_SL g304 ( .A(n_224), .B(n_305), .Y(n_304) );
NAND2x1p5_ASAP7_75t_L g461 ( .A(n_224), .B(n_462), .Y(n_461) );
AND2x2_ASAP7_75t_L g486 ( .A(n_224), .B(n_288), .Y(n_486) );
AND2x4_ASAP7_75t_L g224 ( .A(n_225), .B(n_248), .Y(n_224) );
INVx2_ASAP7_75t_L g225 ( .A(n_226), .Y(n_225) );
INVx2_ASAP7_75t_L g269 ( .A(n_226), .Y(n_269) );
AND2x2_ASAP7_75t_L g372 ( .A(n_226), .B(n_373), .Y(n_372) );
INVx1_ASAP7_75t_L g390 ( .A(n_226), .Y(n_390) );
AND2x2_ASAP7_75t_L g415 ( .A(n_226), .B(n_248), .Y(n_415) );
AND2x4_ASAP7_75t_L g226 ( .A(n_227), .B(n_228), .Y(n_226) );
NAND3xp33_ASAP7_75t_L g323 ( .A(n_228), .B(n_324), .C(n_326), .Y(n_323) );
NAND3xp33_ASAP7_75t_L g228 ( .A(n_229), .B(n_235), .C(n_242), .Y(n_228) );
A2O1A1Ixp33_ASAP7_75t_L g229 ( .A1(n_230), .A2(n_231), .B(n_233), .C(n_234), .Y(n_229) );
INVx2_ASAP7_75t_SL g231 ( .A(n_232), .Y(n_231) );
AOI21xp5_ASAP7_75t_L g545 ( .A1(n_234), .A2(n_546), .B(n_547), .Y(n_545) );
AOI21xp5_ASAP7_75t_L g615 ( .A1(n_234), .A2(n_616), .B(n_617), .Y(n_615) );
OAI221xp5_ASAP7_75t_L g235 ( .A1(n_236), .A2(n_237), .B1(n_238), .B2(n_239), .C(n_240), .Y(n_235) );
INVx2_ASAP7_75t_L g263 ( .A(n_236), .Y(n_263) );
INVx1_ASAP7_75t_L g240 ( .A(n_241), .Y(n_240) );
OAI22xp5_ASAP7_75t_L g250 ( .A1(n_241), .A2(n_251), .B1(n_253), .B2(n_257), .Y(n_250) );
INVx2_ASAP7_75t_SL g256 ( .A(n_241), .Y(n_256) );
NOR2xp33_ASAP7_75t_L g242 ( .A(n_243), .B(n_244), .Y(n_242) );
INVx2_ASAP7_75t_L g328 ( .A(n_244), .Y(n_328) );
AOI21x1_ASAP7_75t_L g244 ( .A1(n_245), .A2(n_246), .B(n_247), .Y(n_244) );
AO21x2_ASAP7_75t_L g295 ( .A1(n_245), .A2(n_246), .B(n_247), .Y(n_295) );
INVx1_ASAP7_75t_L g270 ( .A(n_248), .Y(n_270) );
OAI21x1_ASAP7_75t_L g249 ( .A1(n_250), .A2(n_258), .B(n_264), .Y(n_249) );
INVx2_ASAP7_75t_L g251 ( .A(n_252), .Y(n_251) );
NAND2xp5_ASAP7_75t_L g253 ( .A(n_254), .B(n_256), .Y(n_253) );
INVx2_ASAP7_75t_L g254 ( .A(n_255), .Y(n_254) );
INVx2_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
NAND2xp5_ASAP7_75t_L g591 ( .A(n_264), .B(n_295), .Y(n_591) );
AO32x1_ASAP7_75t_L g266 ( .A1(n_267), .A2(n_286), .A3(n_301), .B1(n_304), .B2(n_308), .Y(n_266) );
AOI32xp33_ASAP7_75t_L g479 ( .A1(n_267), .A2(n_419), .A3(n_480), .B1(n_481), .B2(n_482), .Y(n_479) );
AND2x2_ASAP7_75t_L g267 ( .A(n_268), .B(n_271), .Y(n_267) );
AND2x2_ASAP7_75t_L g341 ( .A(n_268), .B(n_342), .Y(n_341) );
AND2x2_ASAP7_75t_L g347 ( .A(n_268), .B(n_288), .Y(n_347) );
AND2x2_ASAP7_75t_L g399 ( .A(n_268), .B(n_379), .Y(n_399) );
AND2x4_ASAP7_75t_L g268 ( .A(n_269), .B(n_270), .Y(n_268) );
INVx1_ASAP7_75t_L g334 ( .A(n_269), .Y(n_334) );
INVx1_ASAP7_75t_L g388 ( .A(n_271), .Y(n_388) );
NAND2xp5_ASAP7_75t_L g426 ( .A(n_271), .B(n_427), .Y(n_426) );
AND2x2_ASAP7_75t_L g447 ( .A(n_271), .B(n_377), .Y(n_447) );
AND2x2_ASAP7_75t_L g508 ( .A(n_271), .B(n_398), .Y(n_508) );
INVx2_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
AND2x2_ASAP7_75t_L g314 ( .A(n_272), .B(n_310), .Y(n_314) );
INVx1_ASAP7_75t_L g272 ( .A(n_273), .Y(n_272) );
BUFx3_ASAP7_75t_L g311 ( .A(n_273), .Y(n_311) );
OAI21x1_ASAP7_75t_L g273 ( .A1(n_274), .A2(n_277), .B(n_285), .Y(n_273) );
INVx1_ASAP7_75t_L g274 ( .A(n_275), .Y(n_274) );
INVx1_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
BUFx3_ASAP7_75t_L g325 ( .A(n_276), .Y(n_325) );
AOI21xp5_ASAP7_75t_L g281 ( .A1(n_282), .A2(n_283), .B(n_284), .Y(n_281) );
AO21x1_ASAP7_75t_L g603 ( .A1(n_284), .A2(n_604), .B(n_605), .Y(n_603) );
AOI21xp5_ASAP7_75t_L g637 ( .A1(n_284), .A2(n_638), .B(n_639), .Y(n_637) );
NAND2xp5_ASAP7_75t_L g332 ( .A(n_286), .B(n_333), .Y(n_332) );
INVx2_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_287), .B(n_510), .Y(n_509) );
INVx1_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
NAND2xp5_ASAP7_75t_L g371 ( .A(n_288), .B(n_372), .Y(n_371) );
AND2x2_ASAP7_75t_L g501 ( .A(n_288), .B(n_431), .Y(n_501) );
AND2x2_ASAP7_75t_L g505 ( .A(n_288), .B(n_506), .Y(n_505) );
AND2x2_ASAP7_75t_L g288 ( .A(n_289), .B(n_299), .Y(n_288) );
INVx2_ASAP7_75t_L g307 ( .A(n_289), .Y(n_307) );
INVx1_ASAP7_75t_L g481 ( .A(n_289), .Y(n_481) );
AO21x2_ASAP7_75t_L g289 ( .A1(n_290), .A2(n_295), .B(n_296), .Y(n_289) );
NAND2xp33_ASAP7_75t_L g326 ( .A(n_290), .B(n_327), .Y(n_326) );
NOR2xp33_ASAP7_75t_L g570 ( .A(n_295), .B(n_571), .Y(n_570) );
INVx2_ASAP7_75t_L g593 ( .A(n_295), .Y(n_593) );
NOR2xp33_ASAP7_75t_R g296 ( .A(n_297), .B(n_298), .Y(n_296) );
INVx2_ASAP7_75t_L g306 ( .A(n_299), .Y(n_306) );
INVx2_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
INVxp67_ASAP7_75t_L g385 ( .A(n_300), .Y(n_385) );
NAND2x1p5_ASAP7_75t_L g466 ( .A(n_301), .B(n_467), .Y(n_466) );
BUFx3_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
NAND2xp5_ASAP7_75t_L g470 ( .A(n_302), .B(n_403), .Y(n_470) );
AND2x2_ASAP7_75t_L g503 ( .A(n_302), .B(n_388), .Y(n_503) );
BUFx2_ASAP7_75t_L g358 ( .A(n_303), .Y(n_358) );
NAND2xp5_ASAP7_75t_L g354 ( .A(n_304), .B(n_355), .Y(n_354) );
NAND2xp5_ASAP7_75t_L g429 ( .A(n_305), .B(n_430), .Y(n_429) );
AND2x4_ASAP7_75t_L g305 ( .A(n_306), .B(n_307), .Y(n_305) );
INVx2_ASAP7_75t_L g463 ( .A(n_306), .Y(n_463) );
AND2x2_ASAP7_75t_L g389 ( .A(n_307), .B(n_390), .Y(n_389) );
HB1xp67_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
AND2x2_ASAP7_75t_L g514 ( .A(n_309), .B(n_365), .Y(n_514) );
AND2x2_ASAP7_75t_L g309 ( .A(n_310), .B(n_311), .Y(n_309) );
INVx3_ASAP7_75t_L g369 ( .A(n_311), .Y(n_369) );
AND2x2_ASAP7_75t_L g424 ( .A(n_311), .B(n_406), .Y(n_424) );
OAI211xp5_ASAP7_75t_L g312 ( .A1(n_313), .A2(n_316), .B(n_320), .C(n_335), .Y(n_312) );
AND2x2_ASAP7_75t_L g313 ( .A(n_314), .B(n_315), .Y(n_313) );
AND2x2_ASAP7_75t_L g455 ( .A(n_314), .B(n_358), .Y(n_455) );
NAND2xp5_ASAP7_75t_L g484 ( .A(n_314), .B(n_404), .Y(n_484) );
HB1xp67_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
INVx2_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
BUFx2_ASAP7_75t_L g331 ( .A(n_318), .Y(n_331) );
INVx2_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
NAND2xp5_ASAP7_75t_L g477 ( .A(n_319), .B(n_394), .Y(n_477) );
HB1xp67_ASAP7_75t_L g492 ( .A(n_319), .Y(n_492) );
OAI21xp5_ASAP7_75t_L g320 ( .A1(n_321), .A2(n_331), .B(n_332), .Y(n_320) );
INVx1_ASAP7_75t_L g454 ( .A(n_321), .Y(n_454) );
INVx1_ASAP7_75t_L g513 ( .A(n_322), .Y(n_513) );
OR2x2_ASAP7_75t_L g322 ( .A(n_323), .B(n_329), .Y(n_322) );
OR2x2_ASAP7_75t_L g349 ( .A(n_323), .B(n_350), .Y(n_349) );
INVx1_ASAP7_75t_L g386 ( .A(n_323), .Y(n_386) );
INVx1_ASAP7_75t_L g421 ( .A(n_323), .Y(n_421) );
OAI21x1_ASAP7_75t_L g613 ( .A1(n_325), .A2(n_614), .B(n_621), .Y(n_613) );
HB1xp67_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
NAND3xp33_ASAP7_75t_L g573 ( .A(n_328), .B(n_574), .C(n_576), .Y(n_573) );
INVx2_ASAP7_75t_L g350 ( .A(n_329), .Y(n_350) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_329), .B(n_383), .Y(n_382) );
INVx1_ASAP7_75t_L g475 ( .A(n_329), .Y(n_475) );
BUFx3_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
INVx1_ASAP7_75t_L g373 ( .A(n_330), .Y(n_373) );
INVx1_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
AND2x2_ASAP7_75t_L g378 ( .A(n_334), .B(n_379), .Y(n_378) );
INVx1_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
OR2x2_ASAP7_75t_L g443 ( .A(n_336), .B(n_444), .Y(n_443) );
OAI21xp5_ASAP7_75t_SL g485 ( .A1(n_336), .A2(n_486), .B(n_487), .Y(n_485) );
O2A1O1Ixp33_ASAP7_75t_L g487 ( .A1(n_336), .A2(n_488), .B(n_491), .C(n_493), .Y(n_487) );
INVx1_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
OR2x2_ASAP7_75t_L g405 ( .A(n_337), .B(n_406), .Y(n_405) );
NAND4xp25_ASAP7_75t_L g338 ( .A(n_339), .B(n_354), .C(n_362), .D(n_380), .Y(n_338) );
AND2x2_ASAP7_75t_L g339 ( .A(n_340), .B(n_346), .Y(n_339) );
NAND2xp5_ASAP7_75t_L g340 ( .A(n_341), .B(n_343), .Y(n_340) );
AOI22xp33_ASAP7_75t_L g422 ( .A1(n_341), .A2(n_423), .B1(n_425), .B2(n_428), .Y(n_422) );
AND2x4_ASAP7_75t_L g439 ( .A(n_342), .B(n_440), .Y(n_439) );
AND2x2_ASAP7_75t_L g343 ( .A(n_344), .B(n_345), .Y(n_343) );
AND2x2_ASAP7_75t_L g351 ( .A(n_344), .B(n_352), .Y(n_351) );
AND2x2_ASAP7_75t_L g493 ( .A(n_344), .B(n_494), .Y(n_493) );
OAI21xp5_ASAP7_75t_L g346 ( .A1(n_347), .A2(n_348), .B(n_351), .Y(n_346) );
INVx1_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
AND2x4_ASAP7_75t_L g480 ( .A(n_352), .B(n_365), .Y(n_480) );
INVx1_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
INVx1_ASAP7_75t_L g435 ( .A(n_353), .Y(n_435) );
INVxp67_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
AND2x2_ASAP7_75t_L g356 ( .A(n_357), .B(n_359), .Y(n_356) );
AOI32xp33_ASAP7_75t_L g380 ( .A1(n_357), .A2(n_381), .A3(n_384), .B1(n_387), .B2(n_389), .Y(n_380) );
INVx1_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
INVx1_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
AND2x2_ASAP7_75t_L g497 ( .A(n_360), .B(n_369), .Y(n_497) );
AOI22xp33_ASAP7_75t_L g362 ( .A1(n_363), .A2(n_370), .B1(n_374), .B2(n_378), .Y(n_362) );
AND2x2_ASAP7_75t_L g363 ( .A(n_364), .B(n_367), .Y(n_363) );
INVx1_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
OR2x2_ASAP7_75t_L g375 ( .A(n_365), .B(n_376), .Y(n_375) );
INVx2_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
OR2x2_ASAP7_75t_L g412 ( .A(n_366), .B(n_413), .Y(n_412) );
INVx1_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
HB1xp67_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
INVx1_ASAP7_75t_L g383 ( .A(n_369), .Y(n_383) );
INVx1_ASAP7_75t_L g403 ( .A(n_369), .Y(n_403) );
AND2x2_ASAP7_75t_L g434 ( .A(n_369), .B(n_435), .Y(n_434) );
INVx1_ASAP7_75t_L g446 ( .A(n_369), .Y(n_446) );
OAI21xp5_ASAP7_75t_L g502 ( .A1(n_370), .A2(n_428), .B(n_503), .Y(n_502) );
INVx1_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
INVx1_ASAP7_75t_L g449 ( .A(n_372), .Y(n_449) );
BUFx3_ASAP7_75t_L g440 ( .A(n_373), .Y(n_440) );
INVx1_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
INVx1_ASAP7_75t_L g418 ( .A(n_376), .Y(n_418) );
INVx2_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
AND2x2_ASAP7_75t_L g387 ( .A(n_377), .B(n_388), .Y(n_387) );
AND2x2_ASAP7_75t_L g393 ( .A(n_377), .B(n_394), .Y(n_393) );
OAI21xp5_ASAP7_75t_L g504 ( .A1(n_378), .A2(n_480), .B(n_505), .Y(n_504) );
AND2x2_ASAP7_75t_L g414 ( .A(n_379), .B(n_415), .Y(n_414) );
INVx1_ASAP7_75t_L g472 ( .A(n_379), .Y(n_472) );
INVx1_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
INVx1_ASAP7_75t_L g409 ( .A(n_383), .Y(n_409) );
AND2x2_ASAP7_75t_L g384 ( .A(n_385), .B(n_386), .Y(n_384) );
INVx2_ASAP7_75t_L g420 ( .A(n_385), .Y(n_420) );
INVx2_ASAP7_75t_L g431 ( .A(n_390), .Y(n_431) );
NAND4xp25_ASAP7_75t_L g391 ( .A(n_392), .B(n_400), .C(n_416), .D(n_422), .Y(n_391) );
OAI21xp33_ASAP7_75t_L g392 ( .A1(n_393), .A2(n_395), .B(n_399), .Y(n_392) );
AND2x2_ASAP7_75t_L g395 ( .A(n_396), .B(n_398), .Y(n_395) );
INVxp67_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
NAND2xp5_ASAP7_75t_L g408 ( .A(n_398), .B(n_409), .Y(n_408) );
OAI31xp33_ASAP7_75t_L g400 ( .A1(n_401), .A2(n_407), .A3(n_410), .B(n_414), .Y(n_400) );
INVx1_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
NAND2xp5_ASAP7_75t_L g402 ( .A(n_403), .B(n_404), .Y(n_402) );
NOR2xp67_ASAP7_75t_L g459 ( .A(n_403), .B(n_405), .Y(n_459) );
INVx3_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
INVx1_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
INVx1_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
BUFx2_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
AND2x2_ASAP7_75t_L g423 ( .A(n_413), .B(n_424), .Y(n_423) );
BUFx2_ASAP7_75t_L g467 ( .A(n_413), .Y(n_467) );
INVx1_ASAP7_75t_L g494 ( .A(n_413), .Y(n_494) );
AND2x2_ASAP7_75t_L g489 ( .A(n_415), .B(n_490), .Y(n_489) );
HB1xp67_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
AND2x2_ASAP7_75t_L g419 ( .A(n_420), .B(n_421), .Y(n_419) );
AOI32xp33_ASAP7_75t_L g468 ( .A1(n_420), .A2(n_448), .A3(n_469), .B1(n_471), .B2(n_476), .Y(n_468) );
NAND2xp5_ASAP7_75t_L g473 ( .A(n_420), .B(n_474), .Y(n_473) );
INVx1_ASAP7_75t_L g511 ( .A(n_420), .Y(n_511) );
INVx2_ASAP7_75t_L g483 ( .A(n_423), .Y(n_483) );
INVx1_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
INVx1_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
INVx2_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
HB1xp67_ASAP7_75t_L g438 ( .A(n_431), .Y(n_438) );
OAI21xp5_ASAP7_75t_L g432 ( .A1(n_433), .A2(n_436), .B(n_441), .Y(n_432) );
INVxp67_ASAP7_75t_SL g433 ( .A(n_434), .Y(n_433) );
INVx1_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
AND2x2_ASAP7_75t_L g437 ( .A(n_438), .B(n_439), .Y(n_437) );
OAI21xp33_ASAP7_75t_SL g464 ( .A1(n_439), .A2(n_460), .B(n_465), .Y(n_464) );
INVx1_ASAP7_75t_L g500 ( .A(n_440), .Y(n_500) );
INVx2_ASAP7_75t_L g506 ( .A(n_440), .Y(n_506) );
OAI21xp5_ASAP7_75t_L g441 ( .A1(n_442), .A2(n_447), .B(n_448), .Y(n_441) );
INVx1_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
OR2x2_ASAP7_75t_L g444 ( .A(n_445), .B(n_446), .Y(n_444) );
INVx1_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
NOR3xp33_ASAP7_75t_L g450 ( .A(n_451), .B(n_478), .C(n_495), .Y(n_450) );
NAND4xp25_ASAP7_75t_SL g451 ( .A(n_452), .B(n_457), .C(n_464), .D(n_468), .Y(n_451) );
AOI22xp5_ASAP7_75t_L g452 ( .A1(n_453), .A2(n_454), .B1(n_455), .B2(n_456), .Y(n_452) );
BUFx2_ASAP7_75t_SL g458 ( .A(n_459), .Y(n_458) );
INVx1_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
INVx1_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
INVx2_ASAP7_75t_SL g465 ( .A(n_466), .Y(n_465) );
INVx1_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
NAND2xp33_ASAP7_75t_SL g471 ( .A(n_472), .B(n_473), .Y(n_471) );
INVx1_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
INVx1_ASAP7_75t_L g512 ( .A(n_475), .Y(n_512) );
INVx1_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
NAND2xp5_ASAP7_75t_L g478 ( .A(n_479), .B(n_485), .Y(n_478) );
INVx1_ASAP7_75t_L g490 ( .A(n_481), .Y(n_490) );
NAND2xp5_ASAP7_75t_L g482 ( .A(n_483), .B(n_484), .Y(n_482) );
INVx1_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
INVx1_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
NAND4xp25_ASAP7_75t_L g495 ( .A(n_496), .B(n_502), .C(n_504), .D(n_507), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_497), .B(n_498), .Y(n_496) );
INVx1_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
NAND2x1p5_ASAP7_75t_L g499 ( .A(n_500), .B(n_501), .Y(n_499) );
AOI22xp5_ASAP7_75t_L g507 ( .A1(n_508), .A2(n_509), .B1(n_513), .B2(n_514), .Y(n_507) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_511), .B(n_512), .Y(n_510) );
NAND4xp75_ASAP7_75t_L g516 ( .A(n_517), .B(n_706), .C(n_754), .D(n_807), .Y(n_516) );
OA211x2_ASAP7_75t_L g517 ( .A1(n_518), .A2(n_566), .B(n_622), .C(n_677), .Y(n_517) );
NOR2xp33_ASAP7_75t_SL g518 ( .A(n_519), .B(n_561), .Y(n_518) );
INVx2_ASAP7_75t_L g519 ( .A(n_520), .Y(n_519) );
AOI21xp5_ASAP7_75t_SL g767 ( .A1(n_520), .A2(n_768), .B(n_770), .Y(n_767) );
OR2x2_ASAP7_75t_L g520 ( .A(n_521), .B(n_534), .Y(n_520) );
AND2x2_ASAP7_75t_L g720 ( .A(n_521), .B(n_535), .Y(n_720) );
INVx1_ASAP7_75t_L g827 ( .A(n_521), .Y(n_827) );
OR2x2_ASAP7_75t_L g838 ( .A(n_521), .B(n_839), .Y(n_838) );
NAND2xp5_ASAP7_75t_L g840 ( .A(n_521), .B(n_673), .Y(n_840) );
INVx2_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
AND2x2_ASAP7_75t_L g733 ( .A(n_522), .B(n_634), .Y(n_733) );
INVx1_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
INVx2_ASAP7_75t_L g565 ( .A(n_523), .Y(n_565) );
INVx1_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
INVx1_ASAP7_75t_L g650 ( .A(n_524), .Y(n_650) );
INVx1_ASAP7_75t_L g712 ( .A(n_524), .Y(n_712) );
INVx1_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
AND2x4_ASAP7_75t_SL g535 ( .A(n_536), .B(n_549), .Y(n_535) );
AND2x2_ASAP7_75t_L g651 ( .A(n_536), .B(n_550), .Y(n_651) );
AND2x2_ASAP7_75t_L g673 ( .A(n_536), .B(n_635), .Y(n_673) );
OR2x2_ASAP7_75t_L g769 ( .A(n_536), .B(n_688), .Y(n_769) );
INVx2_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
AND2x4_ASAP7_75t_L g645 ( .A(n_537), .B(n_646), .Y(n_645) );
OR2x2_ASAP7_75t_L g660 ( .A(n_537), .B(n_661), .Y(n_660) );
INVx1_ASAP7_75t_L g667 ( .A(n_537), .Y(n_667) );
NAND2xp5_ASAP7_75t_L g689 ( .A(n_537), .B(n_650), .Y(n_689) );
AND2x2_ASAP7_75t_L g831 ( .A(n_537), .B(n_681), .Y(n_831) );
AND2x4_ASAP7_75t_L g537 ( .A(n_538), .B(n_544), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_539), .B(n_540), .Y(n_538) );
AOI21xp5_ASAP7_75t_L g544 ( .A1(n_539), .A2(n_545), .B(n_548), .Y(n_544) );
INVx2_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
INVx1_ASAP7_75t_L g564 ( .A(n_550), .Y(n_564) );
INVx1_ASAP7_75t_L g646 ( .A(n_550), .Y(n_646) );
HB1xp67_ASAP7_75t_L g658 ( .A(n_550), .Y(n_658) );
AND2x2_ASAP7_75t_L g668 ( .A(n_550), .B(n_635), .Y(n_668) );
BUFx2_ASAP7_75t_L g671 ( .A(n_550), .Y(n_671) );
INVx2_ASAP7_75t_L g688 ( .A(n_550), .Y(n_688) );
AND2x2_ASAP7_75t_L g830 ( .A(n_550), .B(n_565), .Y(n_830) );
OR2x6_ASAP7_75t_L g550 ( .A(n_551), .B(n_554), .Y(n_550) );
HB1xp67_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
INVx1_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
OR2x2_ASAP7_75t_L g563 ( .A(n_564), .B(n_565), .Y(n_563) );
AND2x2_ASAP7_75t_L g811 ( .A(n_564), .B(n_565), .Y(n_811) );
NAND2xp5_ASAP7_75t_L g566 ( .A(n_567), .B(n_581), .Y(n_566) );
AND2x2_ASAP7_75t_L g795 ( .A(n_567), .B(n_684), .Y(n_795) );
INVx2_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
AND2x2_ASAP7_75t_L g744 ( .A(n_568), .B(n_624), .Y(n_744) );
AND2x2_ASAP7_75t_L g789 ( .A(n_568), .B(n_598), .Y(n_789) );
INVx1_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
INVx1_ASAP7_75t_L g630 ( .A(n_569), .Y(n_630) );
INVxp67_ASAP7_75t_L g663 ( .A(n_569), .Y(n_663) );
INVx1_ASAP7_75t_L g693 ( .A(n_569), .Y(n_693) );
HB1xp67_ASAP7_75t_L g699 ( .A(n_569), .Y(n_699) );
AND2x2_ASAP7_75t_L g727 ( .A(n_569), .B(n_613), .Y(n_727) );
AND2x2_ASAP7_75t_L g774 ( .A(n_569), .B(n_626), .Y(n_774) );
AND2x2_ASAP7_75t_L g787 ( .A(n_569), .B(n_627), .Y(n_787) );
OR2x2_ASAP7_75t_L g569 ( .A(n_570), .B(n_572), .Y(n_569) );
OAI22xp5_ASAP7_75t_L g572 ( .A1(n_573), .A2(n_577), .B1(n_579), .B2(n_580), .Y(n_572) );
INVx1_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
INVx1_ASAP7_75t_L g779 ( .A(n_581), .Y(n_779) );
AND2x2_ASAP7_75t_L g581 ( .A(n_582), .B(n_598), .Y(n_581) );
INVx1_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
BUFx2_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
AND2x2_ASAP7_75t_L g684 ( .A(n_584), .B(n_629), .Y(n_684) );
INVx1_ASAP7_75t_L g697 ( .A(n_584), .Y(n_697) );
AND2x2_ASAP7_75t_L g730 ( .A(n_584), .B(n_688), .Y(n_730) );
HB1xp67_ASAP7_75t_L g765 ( .A(n_584), .Y(n_765) );
INVx1_ASAP7_75t_L g825 ( .A(n_584), .Y(n_825) );
NAND2x1p5_ASAP7_75t_L g584 ( .A(n_585), .B(n_594), .Y(n_584) );
NAND2x1p5_ASAP7_75t_L g626 ( .A(n_585), .B(n_594), .Y(n_626) );
OA21x2_ASAP7_75t_L g585 ( .A1(n_586), .A2(n_591), .B(n_592), .Y(n_585) );
AOI21xp5_ASAP7_75t_L g618 ( .A1(n_590), .A2(n_619), .B(n_620), .Y(n_618) );
OR2x2_ASAP7_75t_L g594 ( .A(n_591), .B(n_595), .Y(n_594) );
INVx3_ASAP7_75t_L g749 ( .A(n_598), .Y(n_749) );
AND2x2_ASAP7_75t_L g823 ( .A(n_598), .B(n_824), .Y(n_823) );
AND2x2_ASAP7_75t_L g598 ( .A(n_599), .B(n_612), .Y(n_598) );
INVx2_ASAP7_75t_L g629 ( .A(n_599), .Y(n_629) );
OR2x2_ASAP7_75t_L g657 ( .A(n_599), .B(n_626), .Y(n_657) );
AND2x2_ASAP7_75t_L g664 ( .A(n_599), .B(n_626), .Y(n_664) );
INVx1_ASAP7_75t_L g676 ( .A(n_599), .Y(n_676) );
AND2x2_ASAP7_75t_L g691 ( .A(n_599), .B(n_613), .Y(n_691) );
AND2x2_ASAP7_75t_L g696 ( .A(n_599), .B(n_697), .Y(n_696) );
AO31x2_ASAP7_75t_L g599 ( .A1(n_600), .A2(n_603), .A3(n_607), .B(n_611), .Y(n_599) );
INVx1_ASAP7_75t_L g607 ( .A(n_608), .Y(n_607) );
NOR2xp33_ASAP7_75t_L g608 ( .A(n_609), .B(n_610), .Y(n_608) );
INVx1_ASAP7_75t_L g612 ( .A(n_613), .Y(n_612) );
INVx1_ASAP7_75t_L g627 ( .A(n_613), .Y(n_627) );
INVx1_ASAP7_75t_L g655 ( .A(n_613), .Y(n_655) );
AND2x2_ASAP7_75t_L g702 ( .A(n_613), .B(n_625), .Y(n_702) );
AND2x2_ASAP7_75t_L g751 ( .A(n_613), .B(n_630), .Y(n_751) );
AOI211xp5_ASAP7_75t_L g622 ( .A1(n_623), .A2(n_631), .B(n_647), .C(n_652), .Y(n_622) );
AND2x2_ASAP7_75t_L g647 ( .A(n_623), .B(n_648), .Y(n_647) );
AND2x2_ASAP7_75t_L g623 ( .A(n_624), .B(n_628), .Y(n_623) );
AND2x2_ASAP7_75t_L g624 ( .A(n_625), .B(n_627), .Y(n_624) );
INVx2_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
AND2x2_ASAP7_75t_L g692 ( .A(n_626), .B(n_693), .Y(n_692) );
AND2x4_ASAP7_75t_L g701 ( .A(n_628), .B(n_702), .Y(n_701) );
AND2x2_ASAP7_75t_L g628 ( .A(n_629), .B(n_630), .Y(n_628) );
INVx1_ASAP7_75t_L g758 ( .A(n_629), .Y(n_758) );
INVx1_ASAP7_75t_L g631 ( .A(n_632), .Y(n_631) );
NAND2xp5_ASAP7_75t_SL g815 ( .A(n_632), .B(n_816), .Y(n_815) );
NAND2xp5_ASAP7_75t_L g632 ( .A(n_633), .B(n_645), .Y(n_632) );
NAND2xp5_ASAP7_75t_L g741 ( .A(n_633), .B(n_742), .Y(n_741) );
INVx1_ASAP7_75t_L g790 ( .A(n_633), .Y(n_790) );
INVx1_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
INVx1_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
AND2x2_ASAP7_75t_L g777 ( .A(n_645), .B(n_778), .Y(n_777) );
AOI22xp5_ASAP7_75t_L g834 ( .A1(n_645), .A2(n_821), .B1(n_835), .B2(n_837), .Y(n_834) );
AND2x2_ASAP7_75t_L g648 ( .A(n_649), .B(n_651), .Y(n_648) );
OR2x2_ASAP7_75t_L g659 ( .A(n_649), .B(n_660), .Y(n_659) );
AND2x2_ASAP7_75t_L g735 ( .A(n_649), .B(n_673), .Y(n_735) );
INVx1_ASAP7_75t_L g649 ( .A(n_650), .Y(n_649) );
AND2x2_ASAP7_75t_L g680 ( .A(n_650), .B(n_681), .Y(n_680) );
AND2x2_ASAP7_75t_L g704 ( .A(n_650), .B(n_705), .Y(n_704) );
HB1xp67_ASAP7_75t_L g778 ( .A(n_650), .Y(n_778) );
OAI322xp33_ASAP7_75t_L g652 ( .A1(n_653), .A2(n_656), .A3(n_659), .B1(n_662), .B2(n_665), .C1(n_669), .C2(n_674), .Y(n_652) );
INVx2_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
NOR2xp33_ASAP7_75t_L g718 ( .A(n_654), .B(n_719), .Y(n_718) );
BUFx3_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
NAND2xp5_ASAP7_75t_L g675 ( .A(n_655), .B(n_676), .Y(n_675) );
INVxp67_ASAP7_75t_SL g716 ( .A(n_655), .Y(n_716) );
OR2x2_ASAP7_75t_L g656 ( .A(n_657), .B(n_658), .Y(n_656) );
OR2x2_ASAP7_75t_L g836 ( .A(n_657), .B(n_726), .Y(n_836) );
NAND2xp5_ASAP7_75t_L g679 ( .A(n_658), .B(n_680), .Y(n_679) );
AO21x1_ASAP7_75t_L g763 ( .A1(n_659), .A2(n_736), .B(n_764), .Y(n_763) );
INVx4_ASAP7_75t_L g762 ( .A(n_660), .Y(n_762) );
INVx2_ASAP7_75t_L g681 ( .A(n_661), .Y(n_681) );
NAND2xp5_ASAP7_75t_L g662 ( .A(n_663), .B(n_664), .Y(n_662) );
NAND2xp5_ASAP7_75t_L g683 ( .A(n_663), .B(n_684), .Y(n_683) );
INVx2_ASAP7_75t_L g719 ( .A(n_664), .Y(n_719) );
NAND2x1_ASAP7_75t_L g665 ( .A(n_666), .B(n_668), .Y(n_665) );
INVx1_ASAP7_75t_L g710 ( .A(n_666), .Y(n_710) );
AND2x4_ASAP7_75t_SL g722 ( .A(n_666), .B(n_723), .Y(n_722) );
INVx4_ASAP7_75t_R g666 ( .A(n_667), .Y(n_666) );
NAND2xp5_ASAP7_75t_L g800 ( .A(n_667), .B(n_711), .Y(n_800) );
AND2x2_ASAP7_75t_L g806 ( .A(n_668), .B(n_778), .Y(n_806) );
OR2x2_ASAP7_75t_L g669 ( .A(n_670), .B(n_672), .Y(n_669) );
INVx1_ASAP7_75t_L g670 ( .A(n_671), .Y(n_670) );
NAND2xp5_ASAP7_75t_L g761 ( .A(n_671), .B(n_762), .Y(n_761) );
NAND2xp5_ASAP7_75t_L g802 ( .A(n_671), .B(n_733), .Y(n_802) );
INVx1_ASAP7_75t_L g833 ( .A(n_671), .Y(n_833) );
INVx1_ASAP7_75t_L g672 ( .A(n_673), .Y(n_672) );
HB1xp67_ASAP7_75t_L g753 ( .A(n_673), .Y(n_753) );
NAND2xp5_ASAP7_75t_L g832 ( .A(n_673), .B(n_833), .Y(n_832) );
BUFx3_ASAP7_75t_L g674 ( .A(n_675), .Y(n_674) );
NAND2xp5_ASAP7_75t_L g715 ( .A(n_676), .B(n_716), .Y(n_715) );
INVx1_ASAP7_75t_L g738 ( .A(n_676), .Y(n_738) );
AOI221xp5_ASAP7_75t_L g677 ( .A1(n_678), .A2(n_682), .B1(n_685), .B2(n_690), .C(n_694), .Y(n_677) );
INVx1_ASAP7_75t_L g678 ( .A(n_679), .Y(n_678) );
NAND2xp5_ASAP7_75t_L g801 ( .A(n_680), .B(n_687), .Y(n_801) );
NAND2xp5_ASAP7_75t_L g816 ( .A(n_680), .B(n_817), .Y(n_816) );
INVx1_ASAP7_75t_L g705 ( .A(n_681), .Y(n_705) );
OR2x2_ASAP7_75t_L g724 ( .A(n_681), .B(n_712), .Y(n_724) );
AOI22xp33_ASAP7_75t_SL g721 ( .A1(n_682), .A2(n_720), .B1(n_722), .B2(n_725), .Y(n_721) );
INVx1_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
AND2x4_ASAP7_75t_SL g821 ( .A(n_684), .B(n_787), .Y(n_821) );
INVx1_ASAP7_75t_L g685 ( .A(n_686), .Y(n_685) );
OR2x2_ASAP7_75t_L g686 ( .A(n_687), .B(n_689), .Y(n_686) );
NAND2xp5_ASAP7_75t_L g703 ( .A(n_687), .B(n_704), .Y(n_703) );
NAND2xp5_ASAP7_75t_L g783 ( .A(n_687), .B(n_784), .Y(n_783) );
NAND2xp5_ASAP7_75t_L g805 ( .A(n_687), .B(n_733), .Y(n_805) );
BUFx3_ASAP7_75t_L g687 ( .A(n_688), .Y(n_687) );
AND2x2_ASAP7_75t_L g793 ( .A(n_688), .B(n_705), .Y(n_793) );
INVx1_ASAP7_75t_L g742 ( .A(n_689), .Y(n_742) );
AND2x2_ASAP7_75t_L g690 ( .A(n_691), .B(n_692), .Y(n_690) );
AND2x2_ASAP7_75t_L g803 ( .A(n_691), .B(n_774), .Y(n_803) );
INVx2_ASAP7_75t_L g717 ( .A(n_692), .Y(n_717) );
INVx1_ASAP7_75t_L g731 ( .A(n_693), .Y(n_731) );
O2A1O1Ixp33_ASAP7_75t_L g694 ( .A1(n_695), .A2(n_698), .B(n_700), .C(n_703), .Y(n_694) );
AOI21xp33_ASAP7_75t_L g828 ( .A1(n_695), .A2(n_829), .B(n_832), .Y(n_828) );
INVx1_ASAP7_75t_L g695 ( .A(n_696), .Y(n_695) );
NAND2xp5_ASAP7_75t_L g750 ( .A(n_696), .B(n_751), .Y(n_750) );
OR2x2_ASAP7_75t_L g748 ( .A(n_698), .B(n_749), .Y(n_748) );
INVx1_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
INVx2_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
O2A1O1Ixp33_ASAP7_75t_L g822 ( .A1(n_701), .A2(n_823), .B(n_826), .C(n_828), .Y(n_822) );
NOR3x1_ASAP7_75t_SL g706 ( .A(n_707), .B(n_728), .C(n_745), .Y(n_706) );
NAND2xp5_ASAP7_75t_SL g707 ( .A(n_708), .B(n_721), .Y(n_707) );
AOI22xp5_ASAP7_75t_L g708 ( .A1(n_709), .A2(n_713), .B1(n_718), .B2(n_720), .Y(n_708) );
NOR2xp33_ASAP7_75t_L g709 ( .A(n_710), .B(n_711), .Y(n_709) );
BUFx2_ASAP7_75t_L g711 ( .A(n_712), .Y(n_711) );
INVx2_ASAP7_75t_L g713 ( .A(n_714), .Y(n_713) );
OR2x2_ASAP7_75t_L g714 ( .A(n_715), .B(n_717), .Y(n_714) );
INVx2_ASAP7_75t_L g775 ( .A(n_720), .Y(n_775) );
INVx1_ASAP7_75t_L g747 ( .A(n_722), .Y(n_747) );
INVx2_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
OR2x2_ASAP7_75t_L g768 ( .A(n_724), .B(n_769), .Y(n_768) );
INVx1_ASAP7_75t_L g784 ( .A(n_724), .Y(n_784) );
INVx1_ASAP7_75t_L g725 ( .A(n_726), .Y(n_725) );
INVx2_ASAP7_75t_L g726 ( .A(n_727), .Y(n_726) );
AND2x2_ASAP7_75t_L g737 ( .A(n_727), .B(n_738), .Y(n_737) );
OAI322xp33_ASAP7_75t_L g728 ( .A1(n_729), .A2(n_731), .A3(n_732), .B1(n_734), .B2(n_736), .C1(n_739), .C2(n_743), .Y(n_728) );
INVx1_ASAP7_75t_L g729 ( .A(n_730), .Y(n_729) );
AND2x2_ASAP7_75t_L g788 ( .A(n_730), .B(n_789), .Y(n_788) );
INVx2_ASAP7_75t_L g732 ( .A(n_733), .Y(n_732) );
NOR2xp33_ASAP7_75t_L g820 ( .A(n_733), .B(n_762), .Y(n_820) );
INVx2_ASAP7_75t_SL g734 ( .A(n_735), .Y(n_734) );
INVx2_ASAP7_75t_SL g736 ( .A(n_737), .Y(n_736) );
INVx1_ASAP7_75t_L g771 ( .A(n_738), .Y(n_771) );
INVx1_ASAP7_75t_L g739 ( .A(n_740), .Y(n_739) );
INVx1_ASAP7_75t_L g740 ( .A(n_741), .Y(n_740) );
AOI21xp33_ASAP7_75t_L g791 ( .A1(n_741), .A2(n_792), .B(n_794), .Y(n_791) );
INVx2_ASAP7_75t_L g743 ( .A(n_744), .Y(n_743) );
AND2x2_ASAP7_75t_L g757 ( .A(n_744), .B(n_758), .Y(n_757) );
HB1xp67_ASAP7_75t_L g745 ( .A(n_746), .Y(n_745) );
OAI22xp5_ASAP7_75t_L g746 ( .A1(n_747), .A2(n_748), .B1(n_750), .B2(n_752), .Y(n_746) );
INVx2_ASAP7_75t_L g814 ( .A(n_748), .Y(n_814) );
INVx1_ASAP7_75t_L g812 ( .A(n_750), .Y(n_812) );
NAND2xp5_ASAP7_75t_L g764 ( .A(n_751), .B(n_765), .Y(n_764) );
NAND2xp5_ASAP7_75t_L g770 ( .A(n_751), .B(n_771), .Y(n_770) );
AOI222xp33_ASAP7_75t_L g796 ( .A1(n_751), .A2(n_785), .B1(n_797), .B2(n_803), .C1(n_804), .C2(n_806), .Y(n_796) );
INVx1_ASAP7_75t_L g752 ( .A(n_753), .Y(n_752) );
NOR2x1_ASAP7_75t_L g754 ( .A(n_755), .B(n_780), .Y(n_754) );
OAI211xp5_ASAP7_75t_L g755 ( .A1(n_756), .A2(n_759), .B(n_763), .C(n_766), .Y(n_755) );
INVx1_ASAP7_75t_L g756 ( .A(n_757), .Y(n_756) );
INVx1_ASAP7_75t_L g786 ( .A(n_758), .Y(n_786) );
INVxp67_ASAP7_75t_SL g759 ( .A(n_760), .Y(n_759) );
INVx1_ASAP7_75t_L g760 ( .A(n_761), .Y(n_760) );
AND2x4_ASAP7_75t_L g826 ( .A(n_762), .B(n_827), .Y(n_826) );
NOR2xp67_ASAP7_75t_L g766 ( .A(n_767), .B(n_772), .Y(n_766) );
INVx2_ASAP7_75t_L g817 ( .A(n_769), .Y(n_817) );
OAI22xp5_ASAP7_75t_L g772 ( .A1(n_773), .A2(n_775), .B1(n_776), .B2(n_779), .Y(n_772) );
INVx1_ASAP7_75t_L g773 ( .A(n_774), .Y(n_773) );
INVx1_ASAP7_75t_L g776 ( .A(n_777), .Y(n_776) );
NAND2xp5_ASAP7_75t_L g780 ( .A(n_781), .B(n_796), .Y(n_780) );
AOI221xp5_ASAP7_75t_L g781 ( .A1(n_782), .A2(n_785), .B1(n_788), .B2(n_790), .C(n_791), .Y(n_781) );
INVx1_ASAP7_75t_L g782 ( .A(n_783), .Y(n_782) );
AND2x2_ASAP7_75t_L g785 ( .A(n_786), .B(n_787), .Y(n_785) );
INVx1_ASAP7_75t_L g792 ( .A(n_793), .Y(n_792) );
INVx2_ASAP7_75t_L g794 ( .A(n_795), .Y(n_794) );
NAND3xp33_ASAP7_75t_SL g797 ( .A(n_798), .B(n_801), .C(n_802), .Y(n_797) );
INVx1_ASAP7_75t_L g798 ( .A(n_799), .Y(n_798) );
INVx1_ASAP7_75t_L g799 ( .A(n_800), .Y(n_799) );
INVx1_ASAP7_75t_L g804 ( .A(n_805), .Y(n_804) );
OAI21xp5_ASAP7_75t_L g809 ( .A1(n_806), .A2(n_810), .B(n_812), .Y(n_809) );
NOR2x1_ASAP7_75t_L g807 ( .A(n_808), .B(n_818), .Y(n_807) );
NAND2xp5_ASAP7_75t_L g808 ( .A(n_809), .B(n_813), .Y(n_808) );
HB1xp67_ASAP7_75t_L g810 ( .A(n_811), .Y(n_810) );
NAND2xp5_ASAP7_75t_L g813 ( .A(n_814), .B(n_815), .Y(n_813) );
NAND3xp33_ASAP7_75t_SL g818 ( .A(n_819), .B(n_822), .C(n_834), .Y(n_818) );
NAND2xp5_ASAP7_75t_L g819 ( .A(n_820), .B(n_821), .Y(n_819) );
INVx2_ASAP7_75t_L g824 ( .A(n_825), .Y(n_824) );
NAND2xp5_ASAP7_75t_L g829 ( .A(n_830), .B(n_831), .Y(n_829) );
INVx2_ASAP7_75t_L g839 ( .A(n_831), .Y(n_839) );
INVx2_ASAP7_75t_L g835 ( .A(n_836), .Y(n_835) );
NAND2xp33_ASAP7_75t_SL g837 ( .A(n_838), .B(n_840), .Y(n_837) );
INVx6_ASAP7_75t_L g845 ( .A(n_846), .Y(n_845) );
OR2x6_ASAP7_75t_L g846 ( .A(n_847), .B(n_852), .Y(n_846) );
AND2x2_ASAP7_75t_L g847 ( .A(n_848), .B(n_850), .Y(n_847) );
HB1xp67_ASAP7_75t_L g848 ( .A(n_849), .Y(n_848) );
BUFx2_ASAP7_75t_L g850 ( .A(n_851), .Y(n_850) );
INVx1_ASAP7_75t_L g873 ( .A(n_851), .Y(n_873) );
INVx3_ASAP7_75t_L g852 ( .A(n_853), .Y(n_852) );
CKINVDCx11_ASAP7_75t_R g857 ( .A(n_853), .Y(n_857) );
NAND2xp5_ASAP7_75t_L g879 ( .A(n_853), .B(n_880), .Y(n_879) );
OAI21xp33_ASAP7_75t_L g854 ( .A1(n_855), .A2(n_858), .B(n_875), .Y(n_854) );
INVx4_ASAP7_75t_L g855 ( .A(n_856), .Y(n_855) );
BUFx6f_ASAP7_75t_L g856 ( .A(n_857), .Y(n_856) );
INVx1_ASAP7_75t_L g858 ( .A(n_859), .Y(n_858) );
INVx1_ASAP7_75t_L g859 ( .A(n_860), .Y(n_859) );
NAND2xp5_ASAP7_75t_L g860 ( .A(n_861), .B(n_867), .Y(n_860) );
INVx1_ASAP7_75t_L g864 ( .A(n_865), .Y(n_864) );
INVx1_ASAP7_75t_L g867 ( .A(n_868), .Y(n_867) );
CKINVDCx8_ASAP7_75t_R g868 ( .A(n_869), .Y(n_868) );
BUFx6f_ASAP7_75t_L g869 ( .A(n_870), .Y(n_869) );
BUFx3_ASAP7_75t_L g884 ( .A(n_870), .Y(n_884) );
BUFx3_ASAP7_75t_L g870 ( .A(n_871), .Y(n_870) );
INVx2_ASAP7_75t_L g871 ( .A(n_872), .Y(n_871) );
NOR2x1p5_ASAP7_75t_L g872 ( .A(n_873), .B(n_874), .Y(n_872) );
CKINVDCx5p33_ASAP7_75t_R g876 ( .A(n_877), .Y(n_876) );
BUFx6f_ASAP7_75t_L g877 ( .A(n_878), .Y(n_877) );
BUFx6f_ASAP7_75t_L g878 ( .A(n_879), .Y(n_878) );
NOR2x1p5_ASAP7_75t_L g881 ( .A(n_882), .B(n_883), .Y(n_881) );
BUFx3_ASAP7_75t_L g883 ( .A(n_884), .Y(n_883) );
BUFx6f_ASAP7_75t_L g885 ( .A(n_886), .Y(n_885) );
BUFx6f_ASAP7_75t_L g900 ( .A(n_886), .Y(n_900) );
AND3x4_ASAP7_75t_L g886 ( .A(n_887), .B(n_892), .C(n_897), .Y(n_886) );
INVx1_ASAP7_75t_L g888 ( .A(n_889), .Y(n_888) );
INVx1_ASAP7_75t_L g889 ( .A(n_890), .Y(n_889) );
INVx1_ASAP7_75t_L g892 ( .A(n_893), .Y(n_892) );
NAND2xp5_ASAP7_75t_L g893 ( .A(n_894), .B(n_895), .Y(n_893) );
INVx1_ASAP7_75t_L g895 ( .A(n_896), .Y(n_895) );
BUFx2_ASAP7_75t_L g898 ( .A(n_899), .Y(n_898) );
INVx5_ASAP7_75t_L g899 ( .A(n_900), .Y(n_899) );
endmodule