module fake_jpeg_29413_n_55 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_55);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_55;

wire n_21;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_23;
wire n_27;
wire n_22;
wire n_47;
wire n_51;
wire n_40;
wire n_19;
wire n_20;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_32;

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

INVx11_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

BUFx8_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

O2A1O1Ixp33_ASAP7_75t_SL g26 ( 
.A1(n_24),
.A2(n_18),
.B(n_17),
.C(n_16),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g32 ( 
.A1(n_26),
.A2(n_25),
.B1(n_22),
.B2(n_19),
.Y(n_32)
);

OAI32xp33_ASAP7_75t_L g27 ( 
.A1(n_20),
.A2(n_14),
.A3(n_13),
.B1(n_11),
.B2(n_4),
.Y(n_27)
);

A2O1A1Ixp33_ASAP7_75t_SL g36 ( 
.A1(n_27),
.A2(n_25),
.B(n_20),
.C(n_3),
.Y(n_36)
);

XNOR2xp5_ASAP7_75t_L g28 ( 
.A(n_21),
.B(n_0),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_SL g37 ( 
.A(n_28),
.B(n_30),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_L g29 ( 
.A1(n_22),
.A2(n_10),
.B1(n_2),
.B2(n_3),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_SL g35 ( 
.A1(n_29),
.A2(n_23),
.B1(n_20),
.B2(n_19),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_24),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_24),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_31),
.B(n_0),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g39 ( 
.A1(n_32),
.A2(n_23),
.B1(n_27),
.B2(n_28),
.Y(n_39)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_30),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_33),
.Y(n_40)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_26),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_34),
.B(n_38),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g42 ( 
.A1(n_35),
.A2(n_2),
.B1(n_6),
.B2(n_7),
.Y(n_42)
);

NAND3xp33_ASAP7_75t_L g45 ( 
.A(n_36),
.B(n_8),
.C(n_9),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g47 ( 
.A1(n_39),
.A2(n_42),
.B1(n_45),
.B2(n_35),
.Y(n_47)
);

MAJIxp5_ASAP7_75t_L g41 ( 
.A(n_37),
.B(n_10),
.C(n_4),
.Y(n_41)
);

MAJIxp5_ASAP7_75t_L g49 ( 
.A(n_41),
.B(n_36),
.C(n_9),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_33),
.B(n_7),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_44),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_47),
.A2(n_48),
.B1(n_36),
.B2(n_40),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g48 ( 
.A1(n_43),
.A2(n_32),
.B1(n_36),
.B2(n_8),
.Y(n_48)
);

MAJIxp5_ASAP7_75t_L g50 ( 
.A(n_49),
.B(n_41),
.C(n_42),
.Y(n_50)
);

MAJx2_ASAP7_75t_L g52 ( 
.A(n_50),
.B(n_51),
.C(n_49),
.Y(n_52)
);

BUFx24_ASAP7_75t_SL g53 ( 
.A(n_52),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_53),
.A2(n_50),
.B1(n_46),
.B2(n_40),
.Y(n_54)
);

INVxp67_ASAP7_75t_SL g55 ( 
.A(n_54),
.Y(n_55)
);


endmodule