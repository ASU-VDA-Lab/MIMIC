module real_jpeg_33782_n_20 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_639, n_7, n_18, n_3, n_5, n_4, n_1, n_19, n_16, n_15, n_13, n_20);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_639;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_19;
input n_16;
input n_15;
input n_13;

output n_20;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_598;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_630;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_541;
wire n_441;
wire n_557;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_553;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_574;
wire n_627;
wire n_595;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_203;
wire n_198;
wire n_500;
wire n_562;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_578;
wire n_456;
wire n_620;
wire n_259;
wire n_556;
wire n_507;
wire n_57;
wire n_157;
wire n_84;
wire n_560;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_565;
wire n_466;
wire n_623;
wire n_353;
wire n_453;
wire n_551;
wire n_230;
wire n_417;
wire n_428;
wire n_216;
wire n_128;
wire n_202;
wire n_605;
wire n_483;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_550;
wire n_233;
wire n_73;
wire n_621;
wire n_532;
wire n_516;
wire n_348;
wire n_473;
wire n_252;
wire n_601;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_288;
wire n_83;
wire n_525;
wire n_221;
wire n_393;
wire n_489;
wire n_611;
wire n_104;
wire n_153;
wire n_634;
wire n_443;
wire n_599;
wire n_337;
wire n_544;
wire n_131;
wire n_439;
wire n_607;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_561;
wire n_98;
wire n_469;
wire n_378;
wire n_200;
wire n_432;
wire n_465;
wire n_569;
wire n_335;
wire n_214;
wire n_113;
wire n_566;
wire n_543;
wire n_251;
wire n_459;
wire n_576;
wire n_139;
wire n_33;
wire n_631;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_577;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_564;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_262;
wire n_334;
wire n_383;
wire n_593;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_590;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_612;
wire n_110;
wire n_195;
wire n_592;
wire n_533;
wire n_289;
wire n_117;
wire n_614;
wire n_193;
wire n_411;
wire n_382;
wire n_278;
wire n_314;
wire n_103;
wire n_559;
wire n_232;
wire n_582;
wire n_615;
wire n_448;
wire n_212;
wire n_284;
wire n_579;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_583;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_589;
wire n_524;
wire n_25;
wire n_480;
wire n_542;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_632;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_633;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_215;
wire n_176;
wire n_323;
wire n_596;
wire n_312;
wire n_617;
wire n_325;
wire n_307;
wire n_316;
wire n_594;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_604;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_412;
wire n_120;
wire n_572;
wire n_155;
wire n_405;
wire n_586;
wire n_548;
wire n_319;
wire n_487;
wire n_93;
wire n_242;
wire n_493;
wire n_637;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_613;
wire n_265;
wire n_231;
wire n_44;
wire n_635;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_531;
wire n_285;
wire n_546;
wire n_112;
wire n_554;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_616;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_563;
wire n_558;
wire n_510;
wire n_396;
wire n_501;
wire n_600;
wire n_392;
wire n_575;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_584;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_622;
wire n_183;
wire n_248;
wire n_192;
wire n_624;
wire n_537;
wire n_318;
wire n_603;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_204;
wire n_158;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_628;
wire n_413;
wire n_585;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_581;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_534;
wire n_256;
wire n_520;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_545;
wire n_484;
wire n_587;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_343;
wire n_292;
wire n_486;
wire n_64;
wire n_608;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_400;
wire n_174;
wire n_388;
wire n_255;
wire n_299;
wire n_243;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_602;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_571;
wire n_610;
wire n_573;
wire n_379;
wire n_141;
wire n_555;
wire n_65;
wire n_188;
wire n_636;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_570;
wire n_28;
wire n_606;
wire n_245;
wire n_451;
wire n_626;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_597;
wire n_618;
wire n_609;
wire n_94;
wire n_547;
wire n_309;
wire n_294;
wire n_619;
wire n_116;
wire n_416;
wire n_513;
wire n_588;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_567;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_549;
wire n_70;
wire n_568;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_580;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_629;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_552;
wire n_408;
wire n_85;
wire n_591;
wire n_625;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

BUFx6f_ASAP7_75t_L g187 ( 
.A(n_0),
.Y(n_187)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_0),
.Y(n_191)
);

BUFx3_ASAP7_75t_L g348 ( 
.A(n_0),
.Y(n_348)
);

BUFx12f_ASAP7_75t_L g549 ( 
.A(n_0),
.Y(n_549)
);

AOI22xp5_ASAP7_75t_L g20 ( 
.A1(n_1),
.A2(n_16),
.B1(n_21),
.B2(n_24),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_2),
.Y(n_47)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_2),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_3),
.A2(n_117),
.B1(n_120),
.B2(n_121),
.Y(n_116)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_3),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_3),
.A2(n_120),
.B1(n_154),
.B2(n_204),
.Y(n_203)
);

AOI22xp33_ASAP7_75t_SL g234 ( 
.A1(n_3),
.A2(n_120),
.B1(n_235),
.B2(n_241),
.Y(n_234)
);

AOI22xp33_ASAP7_75t_L g255 ( 
.A1(n_3),
.A2(n_120),
.B1(n_256),
.B2(n_257),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_4),
.A2(n_296),
.B1(n_298),
.B2(n_299),
.Y(n_295)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_4),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_SL g352 ( 
.A1(n_4),
.A2(n_298),
.B1(n_353),
.B2(n_357),
.Y(n_352)
);

AOI22xp5_ASAP7_75t_L g505 ( 
.A1(n_4),
.A2(n_298),
.B1(n_506),
.B2(n_507),
.Y(n_505)
);

OAI22xp5_ASAP7_75t_L g591 ( 
.A1(n_4),
.A2(n_298),
.B1(n_592),
.B2(n_596),
.Y(n_591)
);

AO22x1_ASAP7_75t_L g148 ( 
.A1(n_5),
.A2(n_149),
.B1(n_152),
.B2(n_153),
.Y(n_148)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_5),
.Y(n_152)
);

AO22x1_ASAP7_75t_L g195 ( 
.A1(n_5),
.A2(n_152),
.B1(n_196),
.B2(n_199),
.Y(n_195)
);

AOI22xp33_ASAP7_75t_SL g224 ( 
.A1(n_5),
.A2(n_152),
.B1(n_225),
.B2(n_226),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_L g31 ( 
.A1(n_6),
.A2(n_32),
.B(n_36),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_6),
.B(n_37),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_6),
.A2(n_273),
.B1(n_277),
.B2(n_278),
.Y(n_272)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_6),
.Y(n_277)
);

AOI22xp33_ASAP7_75t_SL g309 ( 
.A1(n_6),
.A2(n_277),
.B1(n_310),
.B2(n_311),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_SL g440 ( 
.A1(n_6),
.A2(n_277),
.B1(n_441),
.B2(n_445),
.Y(n_440)
);

OAI22xp33_ASAP7_75t_SL g210 ( 
.A1(n_7),
.A2(n_73),
.B1(n_211),
.B2(n_214),
.Y(n_210)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_7),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_7),
.A2(n_214),
.B1(n_304),
.B2(n_308),
.Y(n_303)
);

AOI22xp33_ASAP7_75t_SL g411 ( 
.A1(n_7),
.A2(n_214),
.B1(n_412),
.B2(n_415),
.Y(n_411)
);

OAI22xp5_ASAP7_75t_SL g515 ( 
.A1(n_7),
.A2(n_214),
.B1(n_342),
.B2(n_516),
.Y(n_515)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_8),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_8),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g338 ( 
.A(n_8),
.Y(n_338)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_9),
.Y(n_81)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_9),
.Y(n_88)
);

INVx4_ASAP7_75t_L g142 ( 
.A(n_10),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_10),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g194 ( 
.A(n_10),
.Y(n_194)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_10),
.Y(n_511)
);

AOI22x1_ASAP7_75t_SL g287 ( 
.A1(n_11),
.A2(n_288),
.B1(n_291),
.B2(n_294),
.Y(n_287)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_11),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g419 ( 
.A1(n_11),
.A2(n_294),
.B1(n_420),
.B2(n_422),
.Y(n_419)
);

AOI22xp33_ASAP7_75t_L g521 ( 
.A1(n_11),
.A2(n_164),
.B1(n_294),
.B2(n_522),
.Y(n_521)
);

AOI22xp33_ASAP7_75t_SL g536 ( 
.A1(n_11),
.A2(n_294),
.B1(n_537),
.B2(n_539),
.Y(n_536)
);

INVx4_ASAP7_75t_L g130 ( 
.A(n_12),
.Y(n_130)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_12),
.Y(n_139)
);

INVx2_ASAP7_75t_L g496 ( 
.A(n_12),
.Y(n_496)
);

OAI21xp5_ASAP7_75t_L g63 ( 
.A1(n_13),
.A2(n_64),
.B(n_70),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_13),
.B(n_71),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_13),
.A2(n_98),
.B1(n_174),
.B2(n_175),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_13),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_13),
.A2(n_164),
.B1(n_174),
.B2(n_282),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_L g341 ( 
.A1(n_13),
.A2(n_174),
.B1(n_342),
.B2(n_343),
.Y(n_341)
);

AOI22xp33_ASAP7_75t_L g363 ( 
.A1(n_14),
.A2(n_317),
.B1(n_364),
.B2(n_365),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_14),
.Y(n_364)
);

AOI22xp33_ASAP7_75t_SL g427 ( 
.A1(n_14),
.A2(n_364),
.B1(n_428),
.B2(n_431),
.Y(n_427)
);

OAI22xp5_ASAP7_75t_SL g483 ( 
.A1(n_14),
.A2(n_364),
.B1(n_484),
.B2(n_487),
.Y(n_483)
);

AOI22xp5_ASAP7_75t_SL g530 ( 
.A1(n_14),
.A2(n_364),
.B1(n_531),
.B2(n_535),
.Y(n_530)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_15),
.A2(n_93),
.B1(n_97),
.B2(n_103),
.Y(n_92)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_15),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_15),
.A2(n_103),
.B1(n_164),
.B2(n_166),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_L g261 ( 
.A1(n_15),
.A2(n_103),
.B1(n_262),
.B2(n_264),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g23 ( 
.A(n_16),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_17),
.B(n_336),
.Y(n_335)
);

AOI21xp5_ASAP7_75t_L g407 ( 
.A1(n_17),
.A2(n_335),
.B(n_408),
.Y(n_407)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_17),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_SL g518 ( 
.A(n_17),
.B(n_78),
.Y(n_518)
);

OAI22xp33_ASAP7_75t_SL g547 ( 
.A1(n_17),
.A2(n_188),
.B1(n_530),
.B2(n_548),
.Y(n_547)
);

OAI32xp33_ASAP7_75t_L g567 ( 
.A1(n_17),
.A2(n_105),
.A3(n_568),
.B1(n_572),
.B2(n_576),
.Y(n_567)
);

AOI22xp33_ASAP7_75t_L g588 ( 
.A1(n_17),
.A2(n_97),
.B1(n_449),
.B2(n_589),
.Y(n_588)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_18),
.Y(n_84)
);

BUFx3_ASAP7_75t_L g91 ( 
.A(n_18),
.Y(n_91)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_18),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g414 ( 
.A(n_18),
.Y(n_414)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_19),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_19),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_19),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_19),
.Y(n_108)
);

BUFx4f_ASAP7_75t_SL g21 ( 
.A(n_22),
.Y(n_21)
);

BUFx12_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

XOR2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_245),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_243),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_216),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_27),
.B(n_216),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_158),
.C(n_178),
.Y(n_27)
);

XNOR2xp5_ASAP7_75t_L g634 ( 
.A(n_28),
.B(n_158),
.Y(n_634)
);

XNOR2xp5_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_75),
.Y(n_28)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_29),
.B(n_218),
.C(n_219),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_29),
.B(n_230),
.Y(n_229)
);

BUFx2_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

AOI22xp5_ASAP7_75t_L g30 ( 
.A1(n_31),
.A2(n_40),
.B1(n_61),
.B2(n_63),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_31),
.A2(n_40),
.B1(n_210),
.B2(n_215),
.Y(n_209)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_34),
.Y(n_297)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g213 ( 
.A(n_35),
.Y(n_213)
);

BUFx6f_ASAP7_75t_L g242 ( 
.A(n_35),
.Y(n_242)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_35),
.Y(n_290)
);

INVx2_ASAP7_75t_SL g37 ( 
.A(n_38),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_L g41 ( 
.A1(n_38),
.A2(n_42),
.B1(n_45),
.B2(n_48),
.Y(n_41)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_38),
.Y(n_366)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_39),
.Y(n_69)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_40),
.Y(n_231)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_40),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g361 ( 
.A1(n_40),
.A2(n_215),
.B1(n_362),
.B2(n_367),
.Y(n_361)
);

AOI22xp5_ASAP7_75t_SL g384 ( 
.A1(n_40),
.A2(n_61),
.B1(n_210),
.B2(n_385),
.Y(n_384)
);

AND2x2_ASAP7_75t_L g40 ( 
.A(n_41),
.B(n_50),
.Y(n_40)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx3_ASAP7_75t_L g240 ( 
.A(n_44),
.Y(n_240)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_47),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_47),
.Y(n_60)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_47),
.Y(n_329)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_50),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_51),
.A2(n_54),
.B1(n_57),
.B2(n_60),
.Y(n_50)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_51),
.Y(n_114)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_52),
.Y(n_177)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_53),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g356 ( 
.A(n_53),
.Y(n_356)
);

BUFx5_ASAP7_75t_L g430 ( 
.A(n_53),
.Y(n_430)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g324 ( 
.A(n_56),
.Y(n_324)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_59),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_59),
.Y(n_123)
);

INVx2_ASAP7_75t_L g333 ( 
.A(n_59),
.Y(n_333)
);

BUFx6f_ASAP7_75t_L g359 ( 
.A(n_59),
.Y(n_359)
);

BUFx6f_ASAP7_75t_L g435 ( 
.A(n_59),
.Y(n_435)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_61),
.Y(n_233)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_62),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_L g285 ( 
.A1(n_62),
.A2(n_286),
.B1(n_287),
.B2(n_295),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_SL g406 ( 
.A1(n_62),
.A2(n_231),
.B1(n_363),
.B2(n_407),
.Y(n_406)
);

NOR2x1_ASAP7_75t_R g448 ( 
.A(n_62),
.B(n_449),
.Y(n_448)
);

INVxp67_ASAP7_75t_L g232 ( 
.A(n_63),
.Y(n_232)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx2_ASAP7_75t_SL g66 ( 
.A(n_67),
.Y(n_66)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_69),
.Y(n_74)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx3_ASAP7_75t_SL g72 ( 
.A(n_73),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_74),
.Y(n_293)
);

XOR2xp5_ASAP7_75t_L g75 ( 
.A(n_76),
.B(n_124),
.Y(n_75)
);

HB1xp67_ASAP7_75t_L g219 ( 
.A(n_76),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_77),
.A2(n_92),
.B1(n_104),
.B2(n_115),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g223 ( 
.A1(n_77),
.A2(n_92),
.B1(n_104),
.B2(n_224),
.Y(n_223)
);

OAI22x1_ASAP7_75t_L g302 ( 
.A1(n_77),
.A2(n_104),
.B1(n_303),
.B2(n_309),
.Y(n_302)
);

OA22x2_ASAP7_75t_L g351 ( 
.A1(n_77),
.A2(n_104),
.B1(n_303),
.B2(n_352),
.Y(n_351)
);

OAI22xp5_ASAP7_75t_L g418 ( 
.A1(n_77),
.A2(n_104),
.B1(n_352),
.B2(n_419),
.Y(n_418)
);

OAI22xp5_ASAP7_75t_L g426 ( 
.A1(n_77),
.A2(n_104),
.B1(n_419),
.B2(n_427),
.Y(n_426)
);

OAI22xp5_ASAP7_75t_SL g587 ( 
.A1(n_77),
.A2(n_104),
.B1(n_427),
.B2(n_588),
.Y(n_587)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g171 ( 
.A1(n_78),
.A2(n_116),
.B1(n_172),
.B2(n_173),
.Y(n_171)
);

AOI22x1_ASAP7_75t_L g386 ( 
.A1(n_78),
.A2(n_172),
.B1(n_173),
.B2(n_387),
.Y(n_386)
);

BUFx2_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

AO21x2_ASAP7_75t_L g104 ( 
.A1(n_79),
.A2(n_105),
.B(n_111),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_80),
.A2(n_82),
.B1(n_85),
.B2(n_89),
.Y(n_79)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

BUFx3_ASAP7_75t_L g110 ( 
.A(n_81),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g487 ( 
.A(n_82),
.Y(n_487)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

BUFx3_ASAP7_75t_L g283 ( 
.A(n_83),
.Y(n_283)
);

INVx4_ASAP7_75t_L g482 ( 
.A(n_83),
.Y(n_482)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_84),
.Y(n_132)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_84),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g417 ( 
.A(n_84),
.Y(n_417)
);

BUFx6f_ASAP7_75t_L g523 ( 
.A(n_84),
.Y(n_523)
);

INVx2_ASAP7_75t_L g575 ( 
.A(n_84),
.Y(n_575)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_88),
.Y(n_113)
);

INVxp67_ASAP7_75t_SL g89 ( 
.A(n_90),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx2_ASAP7_75t_SL g151 ( 
.A(n_91),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_91),
.Y(n_165)
);

INVx2_ASAP7_75t_L g486 ( 
.A(n_91),
.Y(n_486)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx4_ASAP7_75t_L g312 ( 
.A(n_96),
.Y(n_312)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx8_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx2_ASAP7_75t_SL g172 ( 
.A(n_104),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_106),
.B(n_109),
.Y(n_105)
);

INVx5_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

BUFx2_ASAP7_75t_L g225 ( 
.A(n_107),
.Y(n_225)
);

INVx4_ASAP7_75t_L g319 ( 
.A(n_107),
.Y(n_319)
);

INVx8_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g228 ( 
.A(n_108),
.Y(n_228)
);

INVx5_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_112),
.B(n_114),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

BUFx2_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx4_ASAP7_75t_L g307 ( 
.A(n_119),
.Y(n_307)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx2_ASAP7_75t_SL g424 ( 
.A(n_123),
.Y(n_424)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_124),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_124),
.B(n_223),
.Y(n_222)
);

NAND2x1_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_148),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_147),
.Y(n_125)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_126),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_126),
.A2(n_147),
.B1(n_163),
.B2(n_203),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g271 ( 
.A1(n_126),
.A2(n_147),
.B1(n_272),
.B2(n_281),
.Y(n_271)
);

OAI22xp33_ASAP7_75t_SL g369 ( 
.A1(n_126),
.A2(n_147),
.B1(n_203),
.B2(n_281),
.Y(n_369)
);

OAI22xp5_ASAP7_75t_L g410 ( 
.A1(n_126),
.A2(n_147),
.B1(n_272),
.B2(n_411),
.Y(n_410)
);

OAI22xp5_ASAP7_75t_L g519 ( 
.A1(n_126),
.A2(n_147),
.B1(n_520),
.B2(n_521),
.Y(n_519)
);

OAI21xp5_ASAP7_75t_L g612 ( 
.A1(n_126),
.A2(n_613),
.B(n_614),
.Y(n_612)
);

AO21x2_ASAP7_75t_L g126 ( 
.A1(n_127),
.A2(n_133),
.B(n_140),
.Y(n_126)
);

NAND2xp33_ASAP7_75t_SL g127 ( 
.A(n_128),
.B(n_131),
.Y(n_127)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_130),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_130),
.Y(n_144)
);

INVx4_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g501 ( 
.A(n_133),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_137),
.Y(n_133)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_134),
.Y(n_207)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_135),
.Y(n_280)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

BUFx3_ASAP7_75t_L g157 ( 
.A(n_136),
.Y(n_157)
);

BUFx5_ASAP7_75t_L g595 ( 
.A(n_136),
.Y(n_595)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_140),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_141),
.A2(n_143),
.B1(n_144),
.B2(n_145),
.Y(n_140)
);

INVx4_ASAP7_75t_L g500 ( 
.A(n_141),
.Y(n_500)
);

BUFx2_ASAP7_75t_L g516 ( 
.A(n_141),
.Y(n_516)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_142),
.Y(n_198)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_142),
.Y(n_201)
);

BUFx6f_ASAP7_75t_L g266 ( 
.A(n_142),
.Y(n_266)
);

BUFx6f_ASAP7_75t_L g444 ( 
.A(n_142),
.Y(n_444)
);

INVx3_ASAP7_75t_L g542 ( 
.A(n_142),
.Y(n_542)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g344 ( 
.A(n_146),
.Y(n_344)
);

INVx1_ASAP7_75t_SL g161 ( 
.A(n_147),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_SL g545 ( 
.A(n_147),
.B(n_449),
.Y(n_545)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_148),
.A2(n_161),
.B1(n_162),
.B2(n_170),
.Y(n_160)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

INVx3_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVx2_ASAP7_75t_L g479 ( 
.A(n_156),
.Y(n_479)
);

INVx5_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_157),
.Y(n_276)
);

HB1xp67_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

OAI21xp33_ASAP7_75t_L g398 ( 
.A1(n_159),
.A2(n_160),
.B(n_171),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_171),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g476 ( 
.A1(n_161),
.A2(n_170),
.B1(n_477),
.B2(n_483),
.Y(n_476)
);

AOI22xp5_ASAP7_75t_SL g590 ( 
.A1(n_161),
.A2(n_170),
.B1(n_591),
.B2(n_601),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_L g614 ( 
.A(n_161),
.B(n_615),
.Y(n_614)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

INVx1_ASAP7_75t_SL g166 ( 
.A(n_167),
.Y(n_166)
);

BUFx2_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

INVx3_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_175),
.Y(n_589)
);

INVx3_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g633 ( 
.A(n_178),
.B(n_634),
.Y(n_633)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_179),
.A2(n_181),
.B1(n_208),
.B2(n_639),
.Y(n_178)
);

INVxp67_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g399 ( 
.A(n_180),
.B(n_400),
.Y(n_399)
);

AND2x2_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_202),
.Y(n_180)
);

HB1xp67_ASAP7_75t_L g380 ( 
.A(n_181),
.Y(n_380)
);

XOR2xp5_ASAP7_75t_L g400 ( 
.A(n_181),
.B(n_209),
.Y(n_400)
);

AND2x2_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_195),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_188),
.Y(n_182)
);

INVx3_ASAP7_75t_SL g183 ( 
.A(n_184),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_184),
.B(n_195),
.Y(n_371)
);

BUFx6f_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

INVx3_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

HB1xp67_ASAP7_75t_L g513 ( 
.A(n_187),
.Y(n_513)
);

BUFx6f_ASAP7_75t_L g544 ( 
.A(n_187),
.Y(n_544)
);

BUFx3_ASAP7_75t_L g583 ( 
.A(n_187),
.Y(n_583)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_188),
.A2(n_255),
.B1(n_261),
.B2(n_267),
.Y(n_254)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_188),
.Y(n_345)
);

OAI21xp5_ASAP7_75t_L g370 ( 
.A1(n_188),
.A2(n_261),
.B(n_371),
.Y(n_370)
);

OAI22xp5_ASAP7_75t_SL g529 ( 
.A1(n_188),
.A2(n_530),
.B1(n_536),
.B2(n_543),
.Y(n_529)
);

OR2x2_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_192),
.Y(n_188)
);

HB1xp67_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_191),
.Y(n_270)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_191),
.Y(n_439)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_193),
.Y(n_263)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_193),
.Y(n_506)
);

BUFx6f_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_194),
.Y(n_256)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_194),
.Y(n_260)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_194),
.Y(n_342)
);

INVx2_ASAP7_75t_L g447 ( 
.A(n_194),
.Y(n_447)
);

INVx5_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_200),
.Y(n_535)
);

INVx3_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

HB1xp67_ASAP7_75t_L g379 ( 
.A(n_202),
.Y(n_379)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

HB1xp67_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

INVx3_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_220),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_229),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

INVx3_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

INVx8_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

HB1xp67_ASAP7_75t_L g308 ( 
.A(n_228),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_231),
.A2(n_232),
.B1(n_233),
.B2(n_234),
.Y(n_230)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

BUFx4f_ASAP7_75t_SL g241 ( 
.A(n_242),
.Y(n_241)
);

INVx3_ASAP7_75t_SL g300 ( 
.A(n_242),
.Y(n_300)
);

BUFx12f_ASAP7_75t_L g318 ( 
.A(n_242),
.Y(n_318)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_SL g245 ( 
.A1(n_246),
.A2(n_632),
.B(n_636),
.Y(n_245)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_L g247 ( 
.A1(n_248),
.A2(n_469),
.B(n_627),
.Y(n_247)
);

NAND4xp25_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_388),
.C(n_403),
.D(n_462),
.Y(n_248)
);

A2O1A1O1Ixp25_ASAP7_75t_L g627 ( 
.A1(n_249),
.A2(n_388),
.B(n_628),
.C(n_630),
.D(n_631),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_372),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g630 ( 
.A(n_250),
.B(n_372),
.Y(n_630)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_314),
.C(n_368),
.Y(n_250)
);

HB1xp67_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

XNOR2x1_ASAP7_75t_L g468 ( 
.A(n_252),
.B(n_368),
.Y(n_468)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_284),
.Y(n_252)
);

HB1xp67_ASAP7_75t_L g374 ( 
.A(n_253),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_254),
.B(n_271),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g457 ( 
.A(n_254),
.B(n_271),
.Y(n_457)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_255),
.Y(n_346)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

INVx4_ASAP7_75t_L g534 ( 
.A(n_260),
.Y(n_534)
);

HB1xp67_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

BUFx2_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_266),
.Y(n_538)
);

INVx4_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_SL g555 ( 
.A1(n_268),
.A2(n_556),
.B1(n_557),
.B2(n_558),
.Y(n_555)
);

INVx4_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

INVx2_ASAP7_75t_SL g269 ( 
.A(n_270),
.Y(n_269)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

INVx2_ASAP7_75t_SL g275 ( 
.A(n_276),
.Y(n_275)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

INVx2_ASAP7_75t_SL g282 ( 
.A(n_283),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_L g284 ( 
.A1(n_285),
.A2(n_301),
.B1(n_302),
.B2(n_313),
.Y(n_284)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_285),
.Y(n_313)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_287),
.Y(n_367)
);

INVx2_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

INVx4_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

INVx3_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_295),
.Y(n_385)
);

BUFx3_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

HB1xp67_ASAP7_75t_L g376 ( 
.A(n_301),
.Y(n_376)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

INVx3_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

INVx2_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

INVx2_ASAP7_75t_L g310 ( 
.A(n_307),
.Y(n_310)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_309),
.Y(n_387)
);

INVx3_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);

HB1xp67_ASAP7_75t_L g375 ( 
.A(n_313),
.Y(n_375)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_314),
.Y(n_467)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_315),
.B(n_349),
.C(n_360),
.Y(n_314)
);

XOR2xp5_ASAP7_75t_L g453 ( 
.A(n_315),
.B(n_454),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_316),
.B(n_339),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_L g450 ( 
.A1(n_316),
.A2(n_339),
.B1(n_340),
.B2(n_451),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_316),
.Y(n_451)
);

OAI32xp33_ASAP7_75t_SL g316 ( 
.A1(n_317),
.A2(n_319),
.A3(n_320),
.B1(n_325),
.B2(n_334),
.Y(n_316)
);

INVx11_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

INVx1_ASAP7_75t_SL g320 ( 
.A(n_321),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

BUFx3_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

INVx5_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_326),
.B(n_330),
.Y(n_325)
);

INVx2_ASAP7_75t_SL g326 ( 
.A(n_327),
.Y(n_326)
);

BUFx2_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_331),
.Y(n_330)
);

BUFx2_ASAP7_75t_L g331 ( 
.A(n_332),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_335),
.Y(n_334)
);

INVx4_ASAP7_75t_SL g336 ( 
.A(n_337),
.Y(n_336)
);

BUFx6f_ASAP7_75t_L g337 ( 
.A(n_338),
.Y(n_337)
);

INVx1_ASAP7_75t_SL g339 ( 
.A(n_340),
.Y(n_339)
);

AOI22xp5_ASAP7_75t_L g340 ( 
.A1(n_341),
.A2(n_345),
.B1(n_346),
.B2(n_347),
.Y(n_340)
);

AOI22xp5_ASAP7_75t_L g437 ( 
.A1(n_341),
.A2(n_345),
.B1(n_438),
.B2(n_440),
.Y(n_437)
);

BUFx3_ASAP7_75t_L g343 ( 
.A(n_344),
.Y(n_343)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_344),
.Y(n_492)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_345),
.Y(n_504)
);

AOI22xp5_ASAP7_75t_L g580 ( 
.A1(n_345),
.A2(n_440),
.B1(n_515),
.B2(n_581),
.Y(n_580)
);

BUFx6f_ASAP7_75t_L g347 ( 
.A(n_348),
.Y(n_347)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_350),
.Y(n_349)
);

INVxp67_ASAP7_75t_L g350 ( 
.A(n_351),
.Y(n_350)
);

XOR2xp5_ASAP7_75t_L g454 ( 
.A(n_351),
.B(n_455),
.Y(n_454)
);

INVx2_ASAP7_75t_SL g353 ( 
.A(n_354),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_355),
.Y(n_354)
);

INVx2_ASAP7_75t_SL g355 ( 
.A(n_356),
.Y(n_355)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_356),
.Y(n_421)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_356),
.Y(n_571)
);

INVxp33_ASAP7_75t_L g357 ( 
.A(n_358),
.Y(n_357)
);

HB1xp67_ASAP7_75t_L g358 ( 
.A(n_359),
.Y(n_358)
);

HB1xp67_ASAP7_75t_L g360 ( 
.A(n_361),
.Y(n_360)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_361),
.Y(n_455)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_363),
.Y(n_362)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_365),
.Y(n_408)
);

INVx2_ASAP7_75t_SL g365 ( 
.A(n_366),
.Y(n_365)
);

XOR2x2_ASAP7_75t_L g368 ( 
.A(n_369),
.B(n_370),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_369),
.B(n_370),
.Y(n_382)
);

XNOR2xp5_ASAP7_75t_L g372 ( 
.A(n_373),
.B(n_377),
.Y(n_372)
);

MAJIxp5_ASAP7_75t_L g389 ( 
.A(n_373),
.B(n_390),
.C(n_391),
.Y(n_389)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_374),
.B(n_375),
.C(n_376),
.Y(n_373)
);

XNOR2xp5_ASAP7_75t_L g377 ( 
.A(n_378),
.B(n_381),
.Y(n_377)
);

INVxp33_ASAP7_75t_L g391 ( 
.A(n_378),
.Y(n_391)
);

XNOR2x2_ASAP7_75t_L g378 ( 
.A(n_379),
.B(n_380),
.Y(n_378)
);

HB1xp67_ASAP7_75t_L g390 ( 
.A(n_381),
.Y(n_390)
);

XOR2xp5_ASAP7_75t_L g381 ( 
.A(n_382),
.B(n_383),
.Y(n_381)
);

INVxp67_ASAP7_75t_SL g394 ( 
.A(n_382),
.Y(n_394)
);

XNOR2xp5_ASAP7_75t_L g383 ( 
.A(n_384),
.B(n_386),
.Y(n_383)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_384),
.Y(n_395)
);

INVxp33_ASAP7_75t_SL g396 ( 
.A(n_386),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_389),
.B(n_392),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_L g631 ( 
.A(n_389),
.B(n_392),
.Y(n_631)
);

XNOR2xp5_ASAP7_75t_L g392 ( 
.A(n_393),
.B(n_397),
.Y(n_392)
);

MAJIxp5_ASAP7_75t_L g635 ( 
.A(n_393),
.B(n_399),
.C(n_401),
.Y(n_635)
);

MAJIxp5_ASAP7_75t_L g393 ( 
.A(n_394),
.B(n_395),
.C(n_396),
.Y(n_393)
);

AOI22xp5_ASAP7_75t_L g397 ( 
.A1(n_398),
.A2(n_399),
.B1(n_401),
.B2(n_402),
.Y(n_397)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_398),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_399),
.Y(n_402)
);

OR2x2_ASAP7_75t_L g403 ( 
.A(n_404),
.B(n_452),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_404),
.B(n_452),
.Y(n_629)
);

MAJIxp5_ASAP7_75t_SL g404 ( 
.A(n_405),
.B(n_425),
.C(n_450),
.Y(n_404)
);

XNOR2xp5_ASAP7_75t_L g623 ( 
.A(n_405),
.B(n_624),
.Y(n_623)
);

XNOR2xp5_ASAP7_75t_L g405 ( 
.A(n_406),
.B(n_409),
.Y(n_405)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_406),
.Y(n_460)
);

XOR2xp5_ASAP7_75t_L g409 ( 
.A(n_410),
.B(n_418),
.Y(n_409)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_410),
.Y(n_461)
);

INVxp67_ASAP7_75t_SL g615 ( 
.A(n_411),
.Y(n_615)
);

INVx3_ASAP7_75t_L g412 ( 
.A(n_413),
.Y(n_412)
);

BUFx6f_ASAP7_75t_L g413 ( 
.A(n_414),
.Y(n_413)
);

BUFx6f_ASAP7_75t_L g579 ( 
.A(n_414),
.Y(n_579)
);

INVx2_ASAP7_75t_L g600 ( 
.A(n_414),
.Y(n_600)
);

INVx2_ASAP7_75t_SL g415 ( 
.A(n_416),
.Y(n_415)
);

INVx2_ASAP7_75t_SL g416 ( 
.A(n_417),
.Y(n_416)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_418),
.Y(n_459)
);

BUFx3_ASAP7_75t_L g420 ( 
.A(n_421),
.Y(n_420)
);

INVx2_ASAP7_75t_L g422 ( 
.A(n_423),
.Y(n_422)
);

INVx2_ASAP7_75t_L g423 ( 
.A(n_424),
.Y(n_423)
);

XNOR2xp5_ASAP7_75t_L g624 ( 
.A(n_425),
.B(n_450),
.Y(n_624)
);

MAJIxp5_ASAP7_75t_L g425 ( 
.A(n_426),
.B(n_436),
.C(n_448),
.Y(n_425)
);

XNOR2xp5_ASAP7_75t_SL g607 ( 
.A(n_426),
.B(n_608),
.Y(n_607)
);

INVx2_ASAP7_75t_L g428 ( 
.A(n_429),
.Y(n_428)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_430),
.Y(n_429)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_432),
.Y(n_431)
);

INVx2_ASAP7_75t_L g432 ( 
.A(n_433),
.Y(n_432)
);

INVx2_ASAP7_75t_L g433 ( 
.A(n_434),
.Y(n_433)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_435),
.Y(n_434)
);

OAI22xp5_ASAP7_75t_L g608 ( 
.A1(n_436),
.A2(n_437),
.B1(n_448),
.B2(n_609),
.Y(n_608)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_437),
.Y(n_436)
);

HB1xp67_ASAP7_75t_L g438 ( 
.A(n_439),
.Y(n_438)
);

INVx2_ASAP7_75t_L g441 ( 
.A(n_442),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_443),
.Y(n_442)
);

INVx4_ASAP7_75t_L g443 ( 
.A(n_444),
.Y(n_443)
);

INVx2_ASAP7_75t_L g445 ( 
.A(n_446),
.Y(n_445)
);

INVx4_ASAP7_75t_L g446 ( 
.A(n_447),
.Y(n_446)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_448),
.Y(n_609)
);

OAI21xp33_ASAP7_75t_SL g477 ( 
.A1(n_449),
.A2(n_478),
.B(n_480),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_449),
.B(n_481),
.Y(n_480)
);

NOR2xp33_ASAP7_75t_L g551 ( 
.A(n_449),
.B(n_543),
.Y(n_551)
);

NOR2xp33_ASAP7_75t_L g576 ( 
.A(n_449),
.B(n_577),
.Y(n_576)
);

XNOR2xp5_ASAP7_75t_L g452 ( 
.A(n_453),
.B(n_456),
.Y(n_452)
);

MAJIxp5_ASAP7_75t_L g463 ( 
.A(n_453),
.B(n_464),
.C(n_465),
.Y(n_463)
);

XNOR2xp5_ASAP7_75t_L g456 ( 
.A(n_457),
.B(n_458),
.Y(n_456)
);

HB1xp67_ASAP7_75t_L g464 ( 
.A(n_457),
.Y(n_464)
);

HB1xp67_ASAP7_75t_L g465 ( 
.A(n_458),
.Y(n_465)
);

MAJIxp5_ASAP7_75t_L g458 ( 
.A(n_459),
.B(n_460),
.C(n_461),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_463),
.B(n_466),
.Y(n_462)
);

MAJIxp5_ASAP7_75t_L g628 ( 
.A(n_463),
.B(n_466),
.C(n_629),
.Y(n_628)
);

XNOR2x1_ASAP7_75t_L g466 ( 
.A(n_467),
.B(n_468),
.Y(n_466)
);

AOI21x1_ASAP7_75t_L g469 ( 
.A1(n_470),
.A2(n_622),
.B(n_626),
.Y(n_469)
);

OAI21x1_ASAP7_75t_L g470 ( 
.A1(n_471),
.A2(n_605),
.B(n_621),
.Y(n_470)
);

AOI21x1_ASAP7_75t_L g471 ( 
.A1(n_472),
.A2(n_563),
.B(n_604),
.Y(n_471)
);

OAI21x1_ASAP7_75t_L g472 ( 
.A1(n_473),
.A2(n_526),
.B(n_562),
.Y(n_472)
);

AND2x2_ASAP7_75t_L g473 ( 
.A(n_474),
.B(n_502),
.Y(n_473)
);

OR2x2_ASAP7_75t_L g562 ( 
.A(n_474),
.B(n_502),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_SL g474 ( 
.A(n_475),
.B(n_488),
.Y(n_474)
);

AOI22xp5_ASAP7_75t_L g554 ( 
.A1(n_475),
.A2(n_476),
.B1(n_488),
.B2(n_489),
.Y(n_554)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_476),
.Y(n_475)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_479),
.Y(n_478)
);

INVxp67_ASAP7_75t_L g497 ( 
.A(n_480),
.Y(n_497)
);

INVx2_ASAP7_75t_L g481 ( 
.A(n_482),
.Y(n_481)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_483),
.Y(n_520)
);

BUFx2_ASAP7_75t_L g484 ( 
.A(n_485),
.Y(n_484)
);

INVx3_ASAP7_75t_SL g485 ( 
.A(n_486),
.Y(n_485)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_489),
.Y(n_488)
);

AOI22xp5_ASAP7_75t_L g489 ( 
.A1(n_490),
.A2(n_497),
.B1(n_498),
.B2(n_501),
.Y(n_489)
);

NAND2xp33_ASAP7_75t_SL g490 ( 
.A(n_491),
.B(n_493),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_492),
.Y(n_491)
);

BUFx2_ASAP7_75t_L g493 ( 
.A(n_494),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_495),
.Y(n_494)
);

BUFx6f_ASAP7_75t_L g495 ( 
.A(n_496),
.Y(n_495)
);

INVx3_ASAP7_75t_L g498 ( 
.A(n_499),
.Y(n_498)
);

INVx3_ASAP7_75t_L g499 ( 
.A(n_500),
.Y(n_499)
);

XNOR2xp5_ASAP7_75t_L g502 ( 
.A(n_503),
.B(n_517),
.Y(n_502)
);

MAJIxp5_ASAP7_75t_L g564 ( 
.A(n_503),
.B(n_519),
.C(n_524),
.Y(n_564)
);

OAI22xp5_ASAP7_75t_L g503 ( 
.A1(n_504),
.A2(n_505),
.B1(n_512),
.B2(n_514),
.Y(n_503)
);

INVxp67_ASAP7_75t_L g557 ( 
.A(n_504),
.Y(n_557)
);

INVxp67_ASAP7_75t_L g558 ( 
.A(n_505),
.Y(n_558)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_508),
.Y(n_507)
);

BUFx2_ASAP7_75t_L g508 ( 
.A(n_509),
.Y(n_508)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_510),
.Y(n_509)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_511),
.Y(n_510)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_513),
.Y(n_512)
);

INVxp67_ASAP7_75t_L g514 ( 
.A(n_515),
.Y(n_514)
);

OAI22xp5_ASAP7_75t_L g517 ( 
.A1(n_518),
.A2(n_519),
.B1(n_524),
.B2(n_525),
.Y(n_517)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_518),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_519),
.Y(n_525)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_521),
.Y(n_601)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_523),
.Y(n_522)
);

OAI31xp33_ASAP7_75t_L g526 ( 
.A1(n_527),
.A2(n_553),
.A3(n_559),
.B(n_561),
.Y(n_526)
);

NOR2xp33_ASAP7_75t_L g527 ( 
.A(n_528),
.B(n_546),
.Y(n_527)
);

NOR2xp33_ASAP7_75t_L g528 ( 
.A(n_529),
.B(n_545),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_SL g560 ( 
.A(n_529),
.B(n_545),
.Y(n_560)
);

INVx2_ASAP7_75t_L g531 ( 
.A(n_532),
.Y(n_531)
);

INVx2_ASAP7_75t_L g532 ( 
.A(n_533),
.Y(n_532)
);

INVx4_ASAP7_75t_L g533 ( 
.A(n_534),
.Y(n_533)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_535),
.Y(n_552)
);

INVxp67_ASAP7_75t_L g556 ( 
.A(n_536),
.Y(n_556)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_538),
.Y(n_537)
);

BUFx3_ASAP7_75t_L g539 ( 
.A(n_540),
.Y(n_539)
);

INVx2_ASAP7_75t_L g540 ( 
.A(n_541),
.Y(n_540)
);

INVx2_ASAP7_75t_L g541 ( 
.A(n_542),
.Y(n_541)
);

INVx8_ASAP7_75t_L g543 ( 
.A(n_544),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_SL g546 ( 
.A(n_547),
.B(n_550),
.Y(n_546)
);

INVx8_ASAP7_75t_L g548 ( 
.A(n_549),
.Y(n_548)
);

NOR2xp33_ASAP7_75t_SL g550 ( 
.A(n_551),
.B(n_552),
.Y(n_550)
);

NOR2xp33_ASAP7_75t_SL g553 ( 
.A(n_554),
.B(n_555),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g561 ( 
.A(n_554),
.B(n_555),
.Y(n_561)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_560),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_L g563 ( 
.A(n_564),
.B(n_565),
.Y(n_563)
);

NOR2xp67_ASAP7_75t_SL g604 ( 
.A(n_564),
.B(n_565),
.Y(n_604)
);

XNOR2xp5_ASAP7_75t_L g565 ( 
.A(n_566),
.B(n_586),
.Y(n_565)
);

MAJIxp5_ASAP7_75t_L g620 ( 
.A(n_566),
.B(n_590),
.C(n_603),
.Y(n_620)
);

AOI22xp5_ASAP7_75t_L g566 ( 
.A1(n_567),
.A2(n_580),
.B1(n_584),
.B2(n_585),
.Y(n_566)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_567),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_L g611 ( 
.A(n_567),
.B(n_585),
.Y(n_611)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_569),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_570),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_571),
.Y(n_570)
);

INVx2_ASAP7_75t_L g572 ( 
.A(n_573),
.Y(n_572)
);

INVx3_ASAP7_75t_L g573 ( 
.A(n_574),
.Y(n_573)
);

INVx3_ASAP7_75t_L g574 ( 
.A(n_575),
.Y(n_574)
);

INVx1_ASAP7_75t_SL g577 ( 
.A(n_578),
.Y(n_577)
);

BUFx6f_ASAP7_75t_L g578 ( 
.A(n_579),
.Y(n_578)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_580),
.Y(n_585)
);

INVx3_ASAP7_75t_L g581 ( 
.A(n_582),
.Y(n_581)
);

INVx3_ASAP7_75t_L g582 ( 
.A(n_583),
.Y(n_582)
);

AOI22xp5_ASAP7_75t_L g586 ( 
.A1(n_587),
.A2(n_590),
.B1(n_602),
.B2(n_603),
.Y(n_586)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_587),
.Y(n_603)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_590),
.Y(n_602)
);

INVxp67_ASAP7_75t_L g613 ( 
.A(n_591),
.Y(n_613)
);

INVx2_ASAP7_75t_L g592 ( 
.A(n_593),
.Y(n_592)
);

INVx2_ASAP7_75t_L g593 ( 
.A(n_594),
.Y(n_593)
);

INVx2_ASAP7_75t_L g594 ( 
.A(n_595),
.Y(n_594)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_597),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_598),
.Y(n_597)
);

INVx4_ASAP7_75t_L g598 ( 
.A(n_599),
.Y(n_598)
);

INVx4_ASAP7_75t_L g599 ( 
.A(n_600),
.Y(n_599)
);

NOR2xp67_ASAP7_75t_L g605 ( 
.A(n_606),
.B(n_620),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g621 ( 
.A(n_606),
.B(n_620),
.Y(n_621)
);

OAI22xp5_ASAP7_75t_L g606 ( 
.A1(n_607),
.A2(n_610),
.B1(n_618),
.B2(n_619),
.Y(n_606)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_607),
.Y(n_619)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_610),
.Y(n_618)
);

OAI22xp5_ASAP7_75t_L g610 ( 
.A1(n_611),
.A2(n_612),
.B1(n_616),
.B2(n_617),
.Y(n_610)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_611),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_612),
.Y(n_617)
);

MAJIxp5_ASAP7_75t_L g625 ( 
.A(n_612),
.B(n_616),
.C(n_619),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_SL g622 ( 
.A(n_623),
.B(n_625),
.Y(n_622)
);

NOR2xp67_ASAP7_75t_L g626 ( 
.A(n_623),
.B(n_625),
.Y(n_626)
);

NOR2xp33_ASAP7_75t_SL g632 ( 
.A(n_633),
.B(n_635),
.Y(n_632)
);

AND2x2_ASAP7_75t_L g637 ( 
.A(n_633),
.B(n_635),
.Y(n_637)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_637),
.Y(n_636)
);


endmodule