module real_jpeg_26298_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_247;
wire n_146;
wire n_249;
wire n_83;
wire n_78;
wire n_166;
wire n_286;
wire n_176;
wire n_215;
wire n_221;
wire n_288;
wire n_292;
wire n_194;
wire n_104;
wire n_153;
wire n_161;
wire n_207;
wire n_280;
wire n_64;
wire n_177;
wire n_291;
wire n_236;
wire n_47;
wire n_131;
wire n_271;
wire n_281;
wire n_163;
wire n_276;
wire n_22;
wire n_287;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_105;
wire n_40;
wire n_173;
wire n_243;
wire n_255;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_164;
wire n_48;
wire n_293;
wire n_200;
wire n_275;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_242;
wire n_141;
wire n_139;
wire n_33;
wire n_65;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_290;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_285;
wire n_172;
wire n_45;
wire n_211;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_262;
wire n_222;
wire n_118;
wire n_220;
wire n_294;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_198;
wire n_192;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_205;
wire n_258;
wire n_289;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_259;
wire n_103;
wire n_225;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_284;
wire n_277;
wire n_226;
wire n_185;
wire n_125;
wire n_240;
wire n_209;
wire n_55;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_97;
wire n_75;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_169;
wire n_88;
wire n_59;
wire n_279;
wire n_167;
wire n_128;
wire n_213;
wire n_295;
wire n_179;
wire n_202;
wire n_133;
wire n_216;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_181;
wire n_85;
wire n_283;
wire n_256;
wire n_101;
wire n_274;
wire n_182;
wire n_273;
wire n_96;
wire n_253;
wire n_269;
wire n_89;

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_0),
.Y(n_61)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_1),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_2),
.A2(n_67),
.B1(n_73),
.B2(n_122),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_2),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g159 ( 
.A1(n_2),
.A2(n_60),
.B1(n_63),
.B2(n_122),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_2),
.A2(n_42),
.B1(n_43),
.B2(n_122),
.Y(n_213)
);

AOI22xp33_ASAP7_75t_L g247 ( 
.A1(n_2),
.A2(n_29),
.B1(n_31),
.B2(n_122),
.Y(n_247)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

AOI21xp5_ASAP7_75t_L g163 ( 
.A1(n_4),
.A2(n_73),
.B(n_164),
.Y(n_163)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_4),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_4),
.B(n_59),
.Y(n_196)
);

OAI22xp33_ASAP7_75t_L g231 ( 
.A1(n_4),
.A2(n_42),
.B1(n_43),
.B2(n_166),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_4),
.B(n_29),
.C(n_47),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_4),
.B(n_82),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_4),
.A2(n_97),
.B1(n_256),
.B2(n_259),
.Y(n_258)
);

INVx8_ASAP7_75t_SL g62 ( 
.A(n_5),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_6),
.A2(n_71),
.B1(n_72),
.B2(n_75),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_6),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_6),
.A2(n_60),
.B1(n_63),
.B2(n_71),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_6),
.A2(n_42),
.B1(n_43),
.B2(n_71),
.Y(n_214)
);

AOI22xp33_ASAP7_75t_L g242 ( 
.A1(n_6),
.A2(n_29),
.B1(n_31),
.B2(n_71),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_7),
.A2(n_66),
.B1(n_67),
.B2(n_169),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_7),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_7),
.A2(n_60),
.B1(n_63),
.B2(n_169),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g232 ( 
.A1(n_7),
.A2(n_42),
.B1(n_43),
.B2(n_169),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_7),
.A2(n_29),
.B1(n_31),
.B2(n_169),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_8),
.A2(n_42),
.B1(n_43),
.B2(n_53),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_8),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_8),
.A2(n_29),
.B1(n_31),
.B2(n_53),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_8),
.A2(n_53),
.B1(n_60),
.B2(n_63),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_SL g41 ( 
.A1(n_9),
.A2(n_42),
.B1(n_43),
.B2(n_44),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_9),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_9),
.A2(n_44),
.B1(n_60),
.B2(n_63),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_9),
.A2(n_29),
.B1(n_31),
.B2(n_44),
.Y(n_185)
);

BUFx5_ASAP7_75t_L g83 ( 
.A(n_10),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g33 ( 
.A1(n_11),
.A2(n_29),
.B1(n_31),
.B2(n_34),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_11),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_11),
.A2(n_34),
.B1(n_60),
.B2(n_63),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_L g94 ( 
.A1(n_11),
.A2(n_34),
.B1(n_42),
.B2(n_43),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_L g140 ( 
.A1(n_11),
.A2(n_34),
.B1(n_67),
.B2(n_68),
.Y(n_140)
);

INVx13_ASAP7_75t_L g68 ( 
.A(n_12),
.Y(n_68)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_13),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_SL g28 ( 
.A1(n_14),
.A2(n_29),
.B1(n_30),
.B2(n_31),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_14),
.Y(n_30)
);

AOI22xp33_ASAP7_75t_L g78 ( 
.A1(n_14),
.A2(n_30),
.B1(n_67),
.B2(n_73),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_14),
.A2(n_30),
.B1(n_60),
.B2(n_63),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_14),
.A2(n_30),
.B1(n_42),
.B2(n_43),
.Y(n_131)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_15),
.Y(n_37)
);

INVx6_ASAP7_75t_L g110 ( 
.A(n_15),
.Y(n_110)
);

INVx3_ASAP7_75t_L g259 ( 
.A(n_15),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_149),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_147),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_123),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_19),
.B(n_123),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_90),
.C(n_101),
.Y(n_19)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_20),
.A2(n_21),
.B1(n_90),
.B2(n_294),
.Y(n_293)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_54),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_22),
.B(n_56),
.C(n_79),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_38),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_23),
.A2(n_24),
.B1(n_38),
.B2(n_39),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_24),
.Y(n_23)
);

AND2x2_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_32),
.Y(n_24)
);

OAI21xp5_ASAP7_75t_L g241 ( 
.A1(n_25),
.A2(n_97),
.B(n_242),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_28),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

BUFx2_ASAP7_75t_L g250 ( 
.A(n_27),
.Y(n_250)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_28),
.Y(n_100)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_29),
.Y(n_31)
);

AOI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_29),
.A2(n_31),
.B1(n_47),
.B2(n_49),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_31),
.B(n_36),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_SL g260 ( 
.A(n_31),
.B(n_261),
.Y(n_260)
);

OAI21xp5_ASAP7_75t_L g193 ( 
.A1(n_32),
.A2(n_185),
.B(n_194),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g32 ( 
.A(n_33),
.B(n_35),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_33),
.B(n_107),
.Y(n_106)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_35),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_35),
.A2(n_105),
.B1(n_109),
.B2(n_184),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_35),
.A2(n_246),
.B1(n_248),
.B2(n_249),
.Y(n_245)
);

INVx5_ASAP7_75t_L g194 ( 
.A(n_36),
.Y(n_194)
);

INVx5_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_37),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_39),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g39 ( 
.A1(n_40),
.A2(n_45),
.B1(n_51),
.B2(n_52),
.Y(n_39)
);

INVxp67_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

OAI21xp5_ASAP7_75t_L g111 ( 
.A1(n_41),
.A2(n_50),
.B(n_112),
.Y(n_111)
);

OAI22xp33_ASAP7_75t_L g46 ( 
.A1(n_42),
.A2(n_43),
.B1(n_47),
.B2(n_49),
.Y(n_46)
);

AO22x1_ASAP7_75t_L g82 ( 
.A1(n_42),
.A2(n_43),
.B1(n_83),
.B2(n_84),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_42),
.B(n_84),
.Y(n_209)
);

INVx2_ASAP7_75t_SL g42 ( 
.A(n_43),
.Y(n_42)
);

OAI32xp33_ASAP7_75t_L g207 ( 
.A1(n_43),
.A2(n_63),
.A3(n_83),
.B1(n_208),
.B2(n_209),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_43),
.B(n_234),
.Y(n_233)
);

AOI21xp5_ASAP7_75t_L g92 ( 
.A1(n_45),
.A2(n_52),
.B(n_93),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_45),
.B(n_113),
.Y(n_112)
);

AOI21xp5_ASAP7_75t_L g157 ( 
.A1(n_45),
.A2(n_93),
.B(n_131),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_45),
.A2(n_51),
.B1(n_213),
.B2(n_214),
.Y(n_212)
);

AOI21xp5_ASAP7_75t_L g224 ( 
.A1(n_45),
.A2(n_129),
.B(n_214),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_45),
.A2(n_51),
.B1(n_231),
.B2(n_232),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_45),
.A2(n_51),
.B1(n_213),
.B2(n_232),
.Y(n_239)
);

AND2x2_ASAP7_75t_L g45 ( 
.A(n_46),
.B(n_50),
.Y(n_45)
);

INVx13_ASAP7_75t_L g49 ( 
.A(n_47),
.Y(n_49)
);

BUFx24_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_50),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_50),
.B(n_94),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_50),
.B(n_130),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g254 ( 
.A(n_50),
.B(n_166),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_55),
.A2(n_56),
.B1(n_79),
.B2(n_80),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

AOI21xp5_ASAP7_75t_L g56 ( 
.A1(n_57),
.A2(n_70),
.B(n_77),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_57),
.A2(n_59),
.B1(n_70),
.B2(n_121),
.Y(n_120)
);

AOI21xp5_ASAP7_75t_L g137 ( 
.A1(n_57),
.A2(n_138),
.B(n_139),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_57),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_57),
.A2(n_59),
.B1(n_121),
.B2(n_168),
.Y(n_175)
);

AND2x2_ASAP7_75t_SL g57 ( 
.A(n_58),
.B(n_65),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_58),
.B(n_78),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_58),
.B(n_140),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_58),
.A2(n_162),
.B1(n_163),
.B2(n_167),
.Y(n_161)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_60),
.A2(n_62),
.B1(n_63),
.B2(n_64),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_60),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_L g88 ( 
.A1(n_60),
.A2(n_63),
.B1(n_83),
.B2(n_84),
.Y(n_88)
);

A2O1A1Ixp33_ASAP7_75t_L g180 ( 
.A1(n_60),
.A2(n_64),
.B(n_165),
.C(n_181),
.Y(n_180)
);

HAxp5_ASAP7_75t_SL g208 ( 
.A(n_60),
.B(n_166),
.CON(n_208),
.SN(n_208)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_62),
.Y(n_64)
);

OAI22xp33_ASAP7_75t_L g65 ( 
.A1(n_62),
.A2(n_64),
.B1(n_66),
.B2(n_69),
.Y(n_65)
);

NAND3xp33_ASAP7_75t_L g181 ( 
.A(n_62),
.B(n_63),
.C(n_76),
.Y(n_181)
);

INVx8_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx11_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_68),
.Y(n_69)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_68),
.Y(n_74)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_68),
.Y(n_76)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx8_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_76),
.B(n_166),
.Y(n_165)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_78),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_80),
.Y(n_79)
);

OAI21xp5_ASAP7_75t_L g80 ( 
.A1(n_81),
.A2(n_85),
.B(n_86),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_81),
.A2(n_85),
.B1(n_118),
.B2(n_133),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_81),
.A2(n_118),
.B1(n_159),
.B2(n_160),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_81),
.A2(n_118),
.B1(n_159),
.B2(n_198),
.Y(n_197)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_82),
.B(n_88),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_82),
.B(n_89),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_82),
.B(n_117),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_82),
.A2(n_87),
.B1(n_199),
.B2(n_208),
.Y(n_211)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_83),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_87),
.B(n_89),
.Y(n_86)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_87),
.Y(n_118)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_90),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_91),
.A2(n_92),
.B1(n_95),
.B2(n_96),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_92),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_92),
.B(n_95),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_94),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_95),
.A2(n_96),
.B1(n_137),
.B2(n_141),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_96),
.Y(n_95)
);

AOI21xp5_ASAP7_75t_L g96 ( 
.A1(n_97),
.A2(n_98),
.B(n_100),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_L g103 ( 
.A1(n_97),
.A2(n_104),
.B(n_106),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_L g210 ( 
.A1(n_97),
.A2(n_100),
.B(n_106),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_97),
.A2(n_98),
.B1(n_247),
.B2(n_256),
.Y(n_255)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_101),
.B(n_293),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_114),
.C(n_120),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_SL g284 ( 
.A(n_102),
.B(n_285),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_111),
.Y(n_102)
);

XOR2xp5_ASAP7_75t_L g154 ( 
.A(n_103),
.B(n_111),
.Y(n_154)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx5_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx8_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx5_ASAP7_75t_L g263 ( 
.A(n_110),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_112),
.B(n_128),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_114),
.A2(n_115),
.B1(n_120),
.B2(n_286),
.Y(n_285)
);

CKINVDCx14_ASAP7_75t_R g114 ( 
.A(n_115),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_L g115 ( 
.A1(n_116),
.A2(n_118),
.B(n_119),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

OAI21xp33_ASAP7_75t_L g177 ( 
.A1(n_118),
.A2(n_160),
.B(n_178),
.Y(n_177)
);

CKINVDCx14_ASAP7_75t_R g286 ( 
.A(n_120),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_124),
.A2(n_125),
.B1(n_145),
.B2(n_146),
.Y(n_123)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_126),
.A2(n_135),
.B1(n_143),
.B2(n_144),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_126),
.Y(n_143)
);

AOI21xp5_ASAP7_75t_L g126 ( 
.A1(n_127),
.A2(n_132),
.B(n_134),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_127),
.B(n_132),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_135),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_SL g135 ( 
.A(n_136),
.B(n_142),
.Y(n_135)
);

CKINVDCx16_ASAP7_75t_R g141 ( 
.A(n_137),
.Y(n_141)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_145),
.Y(n_146)
);

INVxp67_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_SL g149 ( 
.A1(n_150),
.A2(n_290),
.B(n_295),
.Y(n_149)
);

O2A1O1Ixp33_ASAP7_75t_SL g150 ( 
.A1(n_151),
.A2(n_200),
.B(n_278),
.C(n_289),
.Y(n_150)
);

AND2x2_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_186),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_152),
.B(n_186),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_172),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_154),
.A2(n_155),
.B1(n_170),
.B2(n_171),
.Y(n_153)
);

CKINVDCx16_ASAP7_75t_R g170 ( 
.A(n_154),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_154),
.B(n_171),
.C(n_172),
.Y(n_279)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_155),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_158),
.C(n_161),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_156),
.A2(n_157),
.B1(n_158),
.B2(n_189),
.Y(n_188)
);

CKINVDCx16_ASAP7_75t_R g156 ( 
.A(n_157),
.Y(n_156)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_158),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_SL g187 ( 
.A(n_161),
.B(n_188),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_165),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_166),
.B(n_262),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_168),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_173),
.B(n_179),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_174),
.A2(n_175),
.B1(n_176),
.B2(n_177),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_175),
.B(n_176),
.C(n_179),
.Y(n_287)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_182),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_180),
.A2(n_182),
.B1(n_183),
.B2(n_191),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_180),
.Y(n_191)
);

CKINVDCx16_ASAP7_75t_R g182 ( 
.A(n_183),
.Y(n_182)
);

INVxp67_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_190),
.C(n_192),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_187),
.B(n_276),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_190),
.B(n_192),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_195),
.C(n_197),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_193),
.A2(n_195),
.B1(n_196),
.B2(n_219),
.Y(n_218)
);

CKINVDCx14_ASAP7_75t_R g219 ( 
.A(n_193),
.Y(n_219)
);

CKINVDCx16_ASAP7_75t_R g195 ( 
.A(n_196),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_197),
.B(n_218),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_199),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_202),
.Y(n_200)
);

AOI21xp5_ASAP7_75t_L g202 ( 
.A1(n_203),
.A2(n_273),
.B(n_277),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_L g203 ( 
.A1(n_204),
.A2(n_226),
.B(n_272),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_215),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_205),
.B(n_215),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_211),
.C(n_212),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_206),
.B(n_270),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_SL g206 ( 
.A(n_207),
.B(n_210),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_207),
.B(n_210),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_211),
.B(n_212),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_216),
.A2(n_217),
.B1(n_220),
.B2(n_221),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_216),
.B(n_223),
.C(n_225),
.Y(n_274)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_222),
.A2(n_223),
.B1(n_224),
.B2(n_225),
.Y(n_221)
);

CKINVDCx16_ASAP7_75t_R g225 ( 
.A(n_222),
.Y(n_225)
);

CKINVDCx14_ASAP7_75t_R g223 ( 
.A(n_224),
.Y(n_223)
);

AOI21xp5_ASAP7_75t_L g226 ( 
.A1(n_227),
.A2(n_267),
.B(n_271),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_SL g227 ( 
.A1(n_228),
.A2(n_243),
.B(n_266),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_235),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_229),
.B(n_235),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_SL g229 ( 
.A(n_230),
.B(n_233),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_230),
.B(n_233),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_241),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_237),
.A2(n_238),
.B1(n_239),
.B2(n_240),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_237),
.B(n_240),
.C(n_241),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_238),
.Y(n_237)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_239),
.Y(n_240)
);

INVxp67_ASAP7_75t_L g248 ( 
.A(n_242),
.Y(n_248)
);

AOI21xp33_ASAP7_75t_L g243 ( 
.A1(n_244),
.A2(n_252),
.B(n_265),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_251),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_245),
.B(n_251),
.Y(n_265)
);

CKINVDCx14_ASAP7_75t_R g246 ( 
.A(n_247),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_250),
.Y(n_249)
);

OAI21xp5_ASAP7_75t_SL g252 ( 
.A1(n_253),
.A2(n_257),
.B(n_264),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_255),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_254),
.B(n_255),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g257 ( 
.A(n_258),
.B(n_260),
.Y(n_257)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_268),
.B(n_269),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_SL g271 ( 
.A(n_268),
.B(n_269),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_274),
.B(n_275),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_SL g277 ( 
.A(n_274),
.B(n_275),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_279),
.B(n_280),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_279),
.B(n_280),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_281),
.A2(n_282),
.B1(n_287),
.B2(n_288),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_283),
.B(n_284),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_283),
.B(n_284),
.C(n_288),
.Y(n_291)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_287),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_291),
.B(n_292),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_SL g295 ( 
.A(n_291),
.B(n_292),
.Y(n_295)
);


endmodule