module fake_jpeg_29795_n_115 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_115);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_115;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_43;
wire n_100;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_32),
.Y(n_37)
);

OR2x2_ASAP7_75t_L g38 ( 
.A(n_7),
.B(n_6),
.Y(n_38)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_6),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_10),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_4),
.Y(n_41)
);

BUFx12_ASAP7_75t_L g42 ( 
.A(n_35),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_5),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_13),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_27),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_17),
.Y(n_46)
);

INVx11_ASAP7_75t_L g47 ( 
.A(n_0),
.Y(n_47)
);

BUFx10_ASAP7_75t_L g48 ( 
.A(n_24),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_47),
.Y(n_49)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_49),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g50 ( 
.A(n_41),
.B(n_0),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_50),
.B(n_54),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_43),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_51),
.A2(n_43),
.B1(n_48),
.B2(n_44),
.Y(n_69)
);

BUFx4f_ASAP7_75t_SL g52 ( 
.A(n_48),
.Y(n_52)
);

INVx13_ASAP7_75t_L g63 ( 
.A(n_52),
.Y(n_63)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_53),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_SL g54 ( 
.A(n_38),
.B(n_1),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_38),
.B(n_2),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_55),
.B(n_3),
.Y(n_67)
);

BUFx10_ASAP7_75t_L g56 ( 
.A(n_48),
.Y(n_56)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_56),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g57 ( 
.A(n_54),
.B(n_37),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_57),
.B(n_67),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_50),
.B(n_45),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_59),
.B(n_66),
.Y(n_77)
);

AOI21xp33_ASAP7_75t_L g61 ( 
.A1(n_49),
.A2(n_44),
.B(n_40),
.Y(n_61)
);

OAI21xp5_ASAP7_75t_SL g78 ( 
.A1(n_61),
.A2(n_69),
.B(n_4),
.Y(n_78)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_53),
.B(n_39),
.Y(n_65)
);

AOI21xp5_ASAP7_75t_L g74 ( 
.A1(n_65),
.A2(n_56),
.B(n_42),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_52),
.B(n_45),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_52),
.B(n_40),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_68),
.B(n_12),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_65),
.A2(n_48),
.B1(n_56),
.B2(n_46),
.Y(n_70)
);

AOI21xp5_ASAP7_75t_L g88 ( 
.A1(n_70),
.A2(n_78),
.B(n_79),
.Y(n_88)
);

INVxp67_ASAP7_75t_L g71 ( 
.A(n_65),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_71),
.B(n_75),
.Y(n_89)
);

O2A1O1Ixp33_ASAP7_75t_L g72 ( 
.A1(n_66),
.A2(n_52),
.B(n_56),
.C(n_42),
.Y(n_72)
);

OAI21xp5_ASAP7_75t_L g90 ( 
.A1(n_72),
.A2(n_15),
.B(n_18),
.Y(n_90)
);

HB1xp67_ASAP7_75t_L g73 ( 
.A(n_64),
.Y(n_73)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_73),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_SL g92 ( 
.A1(n_74),
.A2(n_20),
.B(n_21),
.Y(n_92)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_62),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_62),
.A2(n_47),
.B1(n_42),
.B2(n_7),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_76),
.A2(n_81),
.B1(n_23),
.B2(n_25),
.Y(n_96)
);

AOI21xp5_ASAP7_75t_L g79 ( 
.A1(n_59),
.A2(n_5),
.B(n_8),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_63),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_80),
.B(n_83),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_60),
.A2(n_8),
.B1(n_9),
.B2(n_11),
.Y(n_81)
);

NOR2x1_ASAP7_75t_L g82 ( 
.A(n_58),
.B(n_9),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_82),
.B(n_14),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_85),
.B(n_91),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_77),
.B(n_63),
.C(n_16),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_87),
.B(n_95),
.C(n_29),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g102 ( 
.A(n_90),
.B(n_94),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_82),
.B(n_19),
.Y(n_91)
);

AOI21xp5_ASAP7_75t_L g101 ( 
.A1(n_92),
.A2(n_96),
.B(n_97),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_84),
.B(n_80),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_71),
.B(n_22),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_SL g97 ( 
.A1(n_76),
.A2(n_26),
.B(n_28),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_L g98 ( 
.A1(n_88),
.A2(n_72),
.B(n_30),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_98),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_90),
.A2(n_36),
.B1(n_31),
.B2(n_33),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_100),
.B(n_103),
.Y(n_105)
);

XOR2xp5_ASAP7_75t_L g104 ( 
.A(n_89),
.B(n_34),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_104),
.B(n_87),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_L g109 ( 
.A1(n_107),
.A2(n_108),
.B(n_102),
.Y(n_109)
);

AOI321xp33_ASAP7_75t_L g108 ( 
.A1(n_102),
.A2(n_86),
.A3(n_93),
.B1(n_96),
.B2(n_101),
.C(n_99),
.Y(n_108)
);

FAx1_ASAP7_75t_SL g111 ( 
.A(n_109),
.B(n_110),
.CI(n_104),
.CON(n_111),
.SN(n_111)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_105),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_L g112 ( 
.A1(n_111),
.A2(n_106),
.B(n_88),
.Y(n_112)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_112),
.Y(n_113)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_113),
.Y(n_114)
);

XOR2xp5_ASAP7_75t_L g115 ( 
.A(n_114),
.B(n_111),
.Y(n_115)
);


endmodule