module fake_jpeg_16441_n_76 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_76);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_76;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_23;
wire n_10;
wire n_69;
wire n_27;
wire n_64;
wire n_55;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_73;
wire n_19;
wire n_20;
wire n_18;
wire n_59;
wire n_35;
wire n_48;
wire n_68;
wire n_52;
wire n_71;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_65;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_72;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_74;
wire n_11;
wire n_62;
wire n_17;
wire n_25;
wire n_31;
wire n_56;
wire n_67;
wire n_75;
wire n_37;
wire n_43;
wire n_29;
wire n_50;
wire n_12;
wire n_32;
wire n_70;
wire n_15;
wire n_66;

INVx6_ASAP7_75t_SL g9 ( 
.A(n_5),
.Y(n_9)
);

CKINVDCx12_ASAP7_75t_R g10 ( 
.A(n_3),
.Y(n_10)
);

INVxp67_ASAP7_75t_L g11 ( 
.A(n_8),
.Y(n_11)
);

NOR2xp33_ASAP7_75t_L g12 ( 
.A(n_4),
.B(n_1),
.Y(n_12)
);

INVx11_ASAP7_75t_L g13 ( 
.A(n_2),
.Y(n_13)
);

INVx13_ASAP7_75t_L g14 ( 
.A(n_6),
.Y(n_14)
);

BUFx4f_ASAP7_75t_L g15 ( 
.A(n_4),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_2),
.Y(n_16)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

INVx8_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_20),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_SL g21 ( 
.A(n_18),
.B(n_12),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_21),
.B(n_22),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_15),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_17),
.Y(n_23)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_23),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_11),
.B(n_0),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_24),
.B(n_27),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_25),
.Y(n_35)
);

OR2x4_ASAP7_75t_L g26 ( 
.A(n_15),
.B(n_0),
.Y(n_26)
);

AOI21xp5_ASAP7_75t_L g30 ( 
.A1(n_26),
.A2(n_11),
.B(n_0),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_16),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_14),
.Y(n_28)
);

CKINVDCx16_ASAP7_75t_R g29 ( 
.A(n_28),
.Y(n_29)
);

OAI21xp5_ASAP7_75t_L g50 ( 
.A1(n_30),
.A2(n_31),
.B(n_38),
.Y(n_50)
);

OA22x2_ASAP7_75t_L g31 ( 
.A1(n_26),
.A2(n_19),
.B1(n_17),
.B2(n_14),
.Y(n_31)
);

AOI21xp5_ASAP7_75t_L g46 ( 
.A1(n_31),
.A2(n_34),
.B(n_37),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g32 ( 
.A1(n_23),
.A2(n_19),
.B1(n_13),
.B2(n_9),
.Y(n_32)
);

AOI22xp33_ASAP7_75t_SL g42 ( 
.A1(n_32),
.A2(n_40),
.B1(n_10),
.B2(n_27),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_22),
.B(n_1),
.Y(n_34)
);

MAJIxp5_ASAP7_75t_L g44 ( 
.A(n_34),
.B(n_37),
.C(n_30),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_25),
.B(n_6),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_L g40 ( 
.A1(n_20),
.A2(n_9),
.B1(n_8),
.B2(n_7),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_39),
.Y(n_41)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

INVxp67_ASAP7_75t_L g56 ( 
.A(n_42),
.Y(n_56)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_35),
.Y(n_43)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_43),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_44),
.B(n_46),
.Y(n_58)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_45),
.Y(n_51)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_33),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_47),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_36),
.B(n_29),
.Y(n_48)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_48),
.Y(n_52)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_31),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_49),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_54),
.B(n_46),
.Y(n_59)
);

MAJIxp5_ASAP7_75t_L g66 ( 
.A(n_59),
.B(n_60),
.C(n_61),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_52),
.B(n_44),
.Y(n_60)
);

XNOR2xp5_ASAP7_75t_L g61 ( 
.A(n_58),
.B(n_50),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_52),
.B(n_50),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_62),
.A2(n_56),
.B1(n_53),
.B2(n_51),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g63 ( 
.A(n_58),
.B(n_31),
.Y(n_63)
);

AOI21xp5_ASAP7_75t_L g65 ( 
.A1(n_63),
.A2(n_64),
.B(n_56),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_55),
.B(n_42),
.Y(n_64)
);

XNOR2xp5_ASAP7_75t_L g69 ( 
.A(n_65),
.B(n_67),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_61),
.Y(n_68)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_68),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_66),
.Y(n_71)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_71),
.B(n_68),
.Y(n_72)
);

AOI21xp5_ASAP7_75t_SL g74 ( 
.A1(n_72),
.A2(n_73),
.B(n_69),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_70),
.B(n_57),
.C(n_53),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_74),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_75),
.B(n_38),
.Y(n_76)
);


endmodule