module fake_jpeg_30511_n_443 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_443);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_443;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

INVx1_ASAP7_75t_SL g22 ( 
.A(n_6),
.Y(n_22)
);

INVx2_ASAP7_75t_SL g23 ( 
.A(n_11),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_1),
.B(n_3),
.Y(n_24)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

CKINVDCx14_ASAP7_75t_R g29 ( 
.A(n_18),
.Y(n_29)
);

BUFx4f_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

INVxp67_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

INVx5_ASAP7_75t_L g35 ( 
.A(n_18),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_12),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_13),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_1),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_4),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_17),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_0),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_5),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_14),
.Y(n_43)
);

BUFx24_ASAP7_75t_L g44 ( 
.A(n_14),
.Y(n_44)
);

BUFx4f_ASAP7_75t_SL g45 ( 
.A(n_44),
.Y(n_45)
);

INVxp67_ASAP7_75t_SL g108 ( 
.A(n_45),
.Y(n_108)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_25),
.Y(n_46)
);

INVx11_ASAP7_75t_L g95 ( 
.A(n_46),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_21),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_47),
.Y(n_91)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_19),
.Y(n_48)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_48),
.Y(n_98)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_33),
.Y(n_49)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_49),
.Y(n_93)
);

INVx11_ASAP7_75t_L g50 ( 
.A(n_44),
.Y(n_50)
);

INVx5_ASAP7_75t_L g113 ( 
.A(n_50),
.Y(n_113)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_44),
.Y(n_51)
);

BUFx5_ASAP7_75t_L g90 ( 
.A(n_51),
.Y(n_90)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_33),
.Y(n_52)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_52),
.Y(n_96)
);

HB1xp67_ASAP7_75t_L g53 ( 
.A(n_25),
.Y(n_53)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_53),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_36),
.B(n_37),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_54),
.B(n_58),
.Y(n_101)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_26),
.Y(n_55)
);

INVx5_ASAP7_75t_L g119 ( 
.A(n_55),
.Y(n_119)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_19),
.Y(n_56)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_56),
.Y(n_115)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_25),
.Y(n_57)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_57),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_24),
.B(n_9),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_20),
.Y(n_59)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_59),
.Y(n_107)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_34),
.Y(n_60)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_60),
.Y(n_103)
);

INVx11_ASAP7_75t_L g61 ( 
.A(n_44),
.Y(n_61)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_61),
.Y(n_110)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_31),
.Y(n_62)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_62),
.Y(n_136)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_34),
.Y(n_63)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_63),
.Y(n_92)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_26),
.Y(n_64)
);

INVx4_ASAP7_75t_L g116 ( 
.A(n_64),
.Y(n_116)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_34),
.Y(n_65)
);

INVx4_ASAP7_75t_L g134 ( 
.A(n_65),
.Y(n_134)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_21),
.Y(n_66)
);

INVx8_ASAP7_75t_L g100 ( 
.A(n_66),
.Y(n_100)
);

BUFx12f_ASAP7_75t_L g67 ( 
.A(n_21),
.Y(n_67)
);

BUFx4f_ASAP7_75t_SL g120 ( 
.A(n_67),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_24),
.B(n_9),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_68),
.B(n_79),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_42),
.Y(n_69)
);

INVx8_ASAP7_75t_L g104 ( 
.A(n_69),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_30),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_70),
.B(n_75),
.Y(n_137)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_20),
.Y(n_71)
);

INVx4_ASAP7_75t_SL g94 ( 
.A(n_71),
.Y(n_94)
);

BUFx10_ASAP7_75t_L g72 ( 
.A(n_30),
.Y(n_72)
);

INVx1_ASAP7_75t_SL g121 ( 
.A(n_72),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_42),
.Y(n_73)
);

INVx8_ASAP7_75t_L g131 ( 
.A(n_73),
.Y(n_131)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_34),
.Y(n_74)
);

HB1xp67_ASAP7_75t_L g124 ( 
.A(n_74),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_30),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_31),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_76),
.B(n_78),
.Y(n_105)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_42),
.Y(n_77)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_77),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_30),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_43),
.B(n_9),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_36),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_80),
.B(n_82),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_27),
.Y(n_81)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_81),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_37),
.B(n_10),
.Y(n_82)
);

INVx8_ASAP7_75t_L g83 ( 
.A(n_27),
.Y(n_83)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_83),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_40),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_84),
.B(n_86),
.Y(n_133)
);

INVx8_ASAP7_75t_L g85 ( 
.A(n_23),
.Y(n_85)
);

CKINVDCx16_ASAP7_75t_R g123 ( 
.A(n_85),
.Y(n_123)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_28),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_35),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_87),
.Y(n_112)
);

BUFx3_ASAP7_75t_L g88 ( 
.A(n_35),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_88),
.Y(n_106)
);

INVx6_ASAP7_75t_SL g89 ( 
.A(n_23),
.Y(n_89)
);

INVx4_ASAP7_75t_SL g111 ( 
.A(n_89),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_58),
.B(n_43),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_102),
.B(n_109),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_72),
.Y(n_109)
);

CKINVDCx5p33_ASAP7_75t_R g118 ( 
.A(n_45),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_118),
.B(n_128),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_49),
.B(n_22),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_122),
.B(n_125),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_52),
.B(n_22),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_57),
.B(n_22),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_126),
.B(n_135),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_72),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_77),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_130),
.B(n_51),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_59),
.B(n_23),
.Y(n_135)
);

INVx4_ASAP7_75t_L g138 ( 
.A(n_113),
.Y(n_138)
);

INVx1_ASAP7_75t_SL g192 ( 
.A(n_138),
.Y(n_192)
);

INVxp67_ASAP7_75t_L g139 ( 
.A(n_137),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_139),
.B(n_146),
.Y(n_178)
);

AND2x2_ASAP7_75t_L g140 ( 
.A(n_122),
.B(n_89),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_140),
.B(n_154),
.C(n_112),
.Y(n_199)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_93),
.Y(n_142)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_142),
.Y(n_189)
);

INVx3_ASAP7_75t_L g144 ( 
.A(n_113),
.Y(n_144)
);

INVx4_ASAP7_75t_L g182 ( 
.A(n_144),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_135),
.A2(n_47),
.B1(n_73),
.B2(n_69),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_145),
.A2(n_66),
.B1(n_132),
.B2(n_131),
.Y(n_190)
);

BUFx6f_ASAP7_75t_L g147 ( 
.A(n_91),
.Y(n_147)
);

INVx6_ASAP7_75t_L g186 ( 
.A(n_147),
.Y(n_186)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_93),
.Y(n_148)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_148),
.Y(n_193)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_97),
.Y(n_149)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_149),
.Y(n_180)
);

CKINVDCx16_ASAP7_75t_R g150 ( 
.A(n_98),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_150),
.B(n_160),
.Y(n_187)
);

INVx3_ASAP7_75t_L g151 ( 
.A(n_103),
.Y(n_151)
);

INVx4_ASAP7_75t_L g198 ( 
.A(n_151),
.Y(n_198)
);

HB1xp67_ASAP7_75t_L g152 ( 
.A(n_103),
.Y(n_152)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_152),
.Y(n_181)
);

INVx3_ASAP7_75t_L g153 ( 
.A(n_92),
.Y(n_153)
);

INVx3_ASAP7_75t_L g184 ( 
.A(n_153),
.Y(n_184)
);

AND2x2_ASAP7_75t_L g154 ( 
.A(n_125),
.B(n_85),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_91),
.Y(n_155)
);

INVx3_ASAP7_75t_L g195 ( 
.A(n_155),
.Y(n_195)
);

AOI22xp33_ASAP7_75t_SL g157 ( 
.A1(n_94),
.A2(n_29),
.B1(n_35),
.B2(n_55),
.Y(n_157)
);

CKINVDCx16_ASAP7_75t_R g191 ( 
.A(n_157),
.Y(n_191)
);

AOI22xp33_ASAP7_75t_SL g158 ( 
.A1(n_94),
.A2(n_29),
.B1(n_71),
.B2(n_64),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_158),
.A2(n_167),
.B1(n_123),
.B2(n_112),
.Y(n_196)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_96),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_159),
.Y(n_176)
);

INVx4_ASAP7_75t_L g160 ( 
.A(n_92),
.Y(n_160)
);

INVx4_ASAP7_75t_L g161 ( 
.A(n_134),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_161),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_129),
.B(n_133),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_162),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_SL g163 ( 
.A(n_101),
.B(n_40),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_SL g177 ( 
.A(n_163),
.B(n_168),
.Y(n_177)
);

INVx11_ASAP7_75t_L g164 ( 
.A(n_119),
.Y(n_164)
);

OA22x2_ASAP7_75t_L g185 ( 
.A1(n_164),
.A2(n_121),
.B1(n_110),
.B2(n_116),
.Y(n_185)
);

INVx5_ASAP7_75t_L g165 ( 
.A(n_90),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_165),
.B(n_166),
.Y(n_175)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_96),
.Y(n_166)
);

HB1xp67_ASAP7_75t_L g167 ( 
.A(n_134),
.Y(n_167)
);

OR2x2_ASAP7_75t_L g168 ( 
.A(n_117),
.B(n_51),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_105),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_SL g203 ( 
.A(n_170),
.B(n_171),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_117),
.B(n_38),
.Y(n_171)
);

INVx3_ASAP7_75t_L g172 ( 
.A(n_106),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_172),
.B(n_111),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_115),
.B(n_38),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_173),
.B(n_174),
.Y(n_179)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_97),
.Y(n_174)
);

A2O1A1Ixp33_ASAP7_75t_L g183 ( 
.A1(n_169),
.A2(n_126),
.B(n_136),
.C(n_99),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_183),
.B(n_199),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_185),
.A2(n_190),
.B1(n_110),
.B2(n_50),
.Y(n_206)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_188),
.Y(n_214)
);

INVxp67_ASAP7_75t_L g220 ( 
.A(n_196),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_140),
.A2(n_154),
.B1(n_145),
.B2(n_139),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_200),
.A2(n_202),
.B1(n_116),
.B2(n_45),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_169),
.B(n_107),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_201),
.B(n_156),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_140),
.A2(n_32),
.B1(n_132),
.B2(n_114),
.Y(n_202)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_189),
.Y(n_204)
);

BUFx2_ASAP7_75t_L g240 ( 
.A(n_204),
.Y(n_240)
);

AND2x6_ASAP7_75t_L g205 ( 
.A(n_200),
.B(n_168),
.Y(n_205)
);

AO21x1_ASAP7_75t_L g238 ( 
.A1(n_205),
.A2(n_211),
.B(n_177),
.Y(n_238)
);

AND2x2_ASAP7_75t_L g248 ( 
.A(n_206),
.B(n_185),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_201),
.A2(n_156),
.B1(n_154),
.B2(n_100),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_207),
.A2(n_227),
.B1(n_194),
.B2(n_192),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_208),
.B(n_209),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_179),
.B(n_143),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_175),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_210),
.B(n_217),
.Y(n_229)
);

AND2x6_ASAP7_75t_L g211 ( 
.A(n_183),
.B(n_141),
.Y(n_211)
);

INVx3_ASAP7_75t_L g212 ( 
.A(n_186),
.Y(n_212)
);

INVx3_ASAP7_75t_L g232 ( 
.A(n_212),
.Y(n_232)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_189),
.Y(n_213)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_213),
.Y(n_241)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_193),
.Y(n_215)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_215),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_203),
.B(n_170),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_180),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_218),
.B(n_219),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_203),
.B(n_163),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_197),
.B(n_172),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_221),
.B(n_224),
.Y(n_244)
);

INVx8_ASAP7_75t_L g222 ( 
.A(n_186),
.Y(n_222)
);

BUFx3_ASAP7_75t_L g233 ( 
.A(n_222),
.Y(n_233)
);

INVxp67_ASAP7_75t_L g237 ( 
.A(n_223),
.Y(n_237)
);

BUFx24_ASAP7_75t_SL g224 ( 
.A(n_197),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_180),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_225),
.B(n_226),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_175),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_199),
.A2(n_100),
.B1(n_107),
.B2(n_104),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_208),
.B(n_177),
.C(n_179),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_228),
.B(n_246),
.C(n_209),
.Y(n_255)
);

AND2x2_ASAP7_75t_SL g230 ( 
.A(n_214),
.B(n_188),
.Y(n_230)
);

INVx1_ASAP7_75t_SL g267 ( 
.A(n_230),
.Y(n_267)
);

AOI22xp33_ASAP7_75t_L g234 ( 
.A1(n_214),
.A2(n_191),
.B1(n_190),
.B2(n_196),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_234),
.A2(n_239),
.B1(n_248),
.B2(n_227),
.Y(n_253)
);

AOI22xp33_ASAP7_75t_SL g235 ( 
.A1(n_212),
.A2(n_191),
.B1(n_192),
.B2(n_182),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_235),
.A2(n_222),
.B1(n_195),
.B2(n_186),
.Y(n_259)
);

OR2x2_ASAP7_75t_L g263 ( 
.A(n_238),
.B(n_211),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_210),
.A2(n_202),
.B1(n_178),
.B2(n_104),
.Y(n_239)
);

AOI22xp33_ASAP7_75t_L g242 ( 
.A1(n_206),
.A2(n_185),
.B1(n_187),
.B2(n_155),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_242),
.B(n_222),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_SL g243 ( 
.A(n_219),
.B(n_194),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_SL g262 ( 
.A(n_243),
.B(n_176),
.Y(n_262)
);

OAI21xp5_ASAP7_75t_L g245 ( 
.A1(n_216),
.A2(n_181),
.B(n_185),
.Y(n_245)
);

OAI21xp5_ASAP7_75t_L g268 ( 
.A1(n_245),
.A2(n_251),
.B(n_120),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_216),
.B(n_181),
.C(n_149),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_250),
.B(n_142),
.Y(n_272)
);

OAI21xp5_ASAP7_75t_L g251 ( 
.A1(n_220),
.A2(n_223),
.B(n_226),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_249),
.Y(n_252)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_252),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_253),
.A2(n_274),
.B1(n_232),
.B2(n_233),
.Y(n_300)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_249),
.Y(n_254)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_254),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_255),
.B(n_264),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_246),
.B(n_207),
.C(n_205),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_256),
.B(n_266),
.C(n_269),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_L g282 ( 
.A1(n_257),
.A2(n_259),
.B1(n_237),
.B2(n_233),
.Y(n_282)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_229),
.Y(n_258)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_258),
.Y(n_294)
);

AOI21xp5_ASAP7_75t_L g260 ( 
.A1(n_245),
.A2(n_225),
.B(n_218),
.Y(n_260)
);

OAI21xp5_ASAP7_75t_SL g295 ( 
.A1(n_260),
.A2(n_261),
.B(n_271),
.Y(n_295)
);

AOI21xp5_ASAP7_75t_L g261 ( 
.A1(n_251),
.A2(n_182),
.B(n_217),
.Y(n_261)
);

CKINVDCx14_ASAP7_75t_R g305 ( 
.A(n_262),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_263),
.B(n_265),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_231),
.B(n_174),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_240),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_231),
.B(n_124),
.Y(n_266)
);

AOI21xp5_ASAP7_75t_L g288 ( 
.A1(n_268),
.A2(n_248),
.B(n_236),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_230),
.B(n_176),
.C(n_198),
.Y(n_269)
);

INVx13_ASAP7_75t_L g270 ( 
.A(n_232),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_270),
.B(n_275),
.Y(n_298)
);

AND2x6_ASAP7_75t_L g271 ( 
.A(n_238),
.B(n_118),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_272),
.B(n_247),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_243),
.B(n_198),
.Y(n_273)
);

CKINVDCx16_ASAP7_75t_R g280 ( 
.A(n_273),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_248),
.A2(n_195),
.B1(n_147),
.B2(n_204),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_240),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_230),
.B(n_114),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_276),
.B(n_277),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_230),
.B(n_184),
.C(n_159),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_229),
.Y(n_278)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_278),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_236),
.B(n_215),
.Y(n_279)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_279),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_260),
.A2(n_248),
.B1(n_239),
.B2(n_250),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_SL g310 ( 
.A1(n_281),
.A2(n_297),
.B1(n_274),
.B2(n_268),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g331 ( 
.A1(n_282),
.A2(n_300),
.B1(n_303),
.B2(n_288),
.Y(n_331)
);

HB1xp67_ASAP7_75t_L g286 ( 
.A(n_258),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_286),
.B(n_308),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_SL g287 ( 
.A(n_278),
.B(n_244),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g328 ( 
.A(n_287),
.B(n_296),
.Y(n_328)
);

NAND2x1_ASAP7_75t_SL g332 ( 
.A(n_288),
.B(n_138),
.Y(n_332)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_256),
.B(n_238),
.Y(n_289)
);

XOR2xp5_ASAP7_75t_L g327 ( 
.A(n_289),
.B(n_111),
.Y(n_327)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_290),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_279),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_292),
.B(n_241),
.Y(n_321)
);

CKINVDCx16_ASAP7_75t_R g296 ( 
.A(n_252),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_254),
.A2(n_234),
.B1(n_232),
.B2(n_247),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_253),
.A2(n_228),
.B1(n_244),
.B2(n_233),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_267),
.Y(n_304)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_304),
.Y(n_316)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_267),
.Y(n_306)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_306),
.Y(n_323)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_269),
.Y(n_307)
);

CKINVDCx16_ASAP7_75t_R g317 ( 
.A(n_307),
.Y(n_317)
);

CKINVDCx16_ASAP7_75t_R g308 ( 
.A(n_261),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_299),
.B(n_255),
.C(n_266),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_309),
.B(n_314),
.C(n_283),
.Y(n_340)
);

AOI22xp5_ASAP7_75t_L g345 ( 
.A1(n_310),
.A2(n_304),
.B1(n_302),
.B2(n_290),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_L g312 ( 
.A1(n_305),
.A2(n_263),
.B1(n_259),
.B2(n_272),
.Y(n_312)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_312),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_L g313 ( 
.A1(n_291),
.A2(n_271),
.B1(n_277),
.B2(n_241),
.Y(n_313)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_313),
.Y(n_356)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_299),
.B(n_276),
.C(n_264),
.Y(n_314)
);

INVx2_ASAP7_75t_SL g318 ( 
.A(n_298),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_318),
.B(n_319),
.Y(n_343)
);

HB1xp67_ASAP7_75t_L g319 ( 
.A(n_294),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_280),
.B(n_184),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_SL g348 ( 
.A(n_320),
.B(n_324),
.Y(n_348)
);

A2O1A1Ixp33_ASAP7_75t_L g350 ( 
.A1(n_321),
.A2(n_332),
.B(n_120),
.C(n_108),
.Y(n_350)
);

INVx4_ASAP7_75t_L g322 ( 
.A(n_295),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_322),
.B(n_295),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_303),
.B(n_294),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_SL g325 ( 
.A(n_301),
.B(n_13),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_L g334 ( 
.A1(n_325),
.A2(n_329),
.B1(n_292),
.B2(n_293),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_301),
.B(n_213),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_SL g354 ( 
.A(n_326),
.B(n_330),
.Y(n_354)
);

XNOR2xp5_ASAP7_75t_SL g338 ( 
.A(n_327),
.B(n_285),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_SL g329 ( 
.A(n_284),
.B(n_293),
.Y(n_329)
);

NOR2x1_ASAP7_75t_L g330 ( 
.A(n_281),
.B(n_270),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_SL g339 ( 
.A1(n_331),
.A2(n_333),
.B1(n_297),
.B2(n_284),
.Y(n_339)
);

AOI22xp5_ASAP7_75t_L g333 ( 
.A1(n_300),
.A2(n_240),
.B1(n_193),
.B2(n_131),
.Y(n_333)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_334),
.Y(n_360)
);

XNOR2xp5_ASAP7_75t_L g335 ( 
.A(n_314),
.B(n_283),
.Y(n_335)
);

XNOR2xp5_ASAP7_75t_L g368 ( 
.A(n_335),
.B(n_337),
.Y(n_368)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_336),
.Y(n_364)
);

XOR2xp5_ASAP7_75t_L g337 ( 
.A(n_327),
.B(n_289),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g372 ( 
.A(n_338),
.B(n_340),
.C(n_341),
.Y(n_372)
);

AOI22xp5_ASAP7_75t_L g359 ( 
.A1(n_339),
.A2(n_330),
.B1(n_353),
.B2(n_342),
.Y(n_359)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_309),
.B(n_307),
.C(n_285),
.Y(n_341)
);

XOR2xp5_ASAP7_75t_L g342 ( 
.A(n_331),
.B(n_306),
.Y(n_342)
);

MAJIxp5_ASAP7_75t_L g374 ( 
.A(n_342),
.B(n_347),
.C(n_353),
.Y(n_374)
);

OAI22xp5_ASAP7_75t_SL g369 ( 
.A1(n_345),
.A2(n_164),
.B1(n_95),
.B2(n_121),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_325),
.B(n_302),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_346),
.B(n_349),
.Y(n_370)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_317),
.B(n_166),
.C(n_148),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_322),
.B(n_151),
.Y(n_349)
);

CKINVDCx14_ASAP7_75t_R g373 ( 
.A(n_350),
.Y(n_373)
);

OAI22xp5_ASAP7_75t_L g351 ( 
.A1(n_328),
.A2(n_81),
.B1(n_39),
.B2(n_28),
.Y(n_351)
);

AOI322xp5_ASAP7_75t_L g358 ( 
.A1(n_351),
.A2(n_311),
.A3(n_318),
.B1(n_323),
.B2(n_165),
.C1(n_315),
.C2(n_119),
.Y(n_358)
);

OAI22xp5_ASAP7_75t_SL g352 ( 
.A1(n_333),
.A2(n_127),
.B1(n_144),
.B2(n_39),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_352),
.B(n_318),
.Y(n_363)
);

XOR2xp5_ASAP7_75t_L g353 ( 
.A(n_310),
.B(n_120),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_L g355 ( 
.A(n_316),
.B(n_161),
.C(n_160),
.Y(n_355)
);

MAJIxp5_ASAP7_75t_L g376 ( 
.A(n_355),
.B(n_357),
.C(n_63),
.Y(n_376)
);

MAJIxp5_ASAP7_75t_L g357 ( 
.A(n_316),
.B(n_153),
.C(n_127),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_SL g380 ( 
.A(n_358),
.B(n_375),
.Y(n_380)
);

OAI22xp5_ASAP7_75t_SL g379 ( 
.A1(n_359),
.A2(n_373),
.B1(n_374),
.B2(n_362),
.Y(n_379)
);

A2O1A1O1Ixp25_ASAP7_75t_L g361 ( 
.A1(n_344),
.A2(n_315),
.B(n_321),
.C(n_323),
.D(n_332),
.Y(n_361)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_361),
.Y(n_384)
);

OAI21xp5_ASAP7_75t_L g362 ( 
.A1(n_354),
.A2(n_329),
.B(n_332),
.Y(n_362)
);

AOI21xp5_ASAP7_75t_L g387 ( 
.A1(n_362),
.A2(n_16),
.B(n_11),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_L g386 ( 
.A(n_363),
.B(n_367),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_343),
.B(n_348),
.Y(n_365)
);

OAI21x1_ASAP7_75t_L g392 ( 
.A1(n_365),
.A2(n_377),
.B(n_16),
.Y(n_392)
);

AOI21xp5_ASAP7_75t_L g366 ( 
.A1(n_356),
.A2(n_10),
.B(n_17),
.Y(n_366)
);

OAI21xp5_ASAP7_75t_L g383 ( 
.A1(n_366),
.A2(n_370),
.B(n_364),
.Y(n_383)
);

INVx13_ASAP7_75t_L g367 ( 
.A(n_350),
.Y(n_367)
);

XOR2xp5_ASAP7_75t_L g390 ( 
.A(n_369),
.B(n_67),
.Y(n_390)
);

HB1xp67_ASAP7_75t_L g371 ( 
.A(n_335),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_L g391 ( 
.A(n_371),
.B(n_376),
.Y(n_391)
);

CKINVDCx20_ASAP7_75t_R g375 ( 
.A(n_345),
.Y(n_375)
);

A2O1A1O1Ixp25_ASAP7_75t_L g377 ( 
.A1(n_337),
.A2(n_41),
.B(n_17),
.C(n_8),
.D(n_18),
.Y(n_377)
);

AOI22xp5_ASAP7_75t_L g378 ( 
.A1(n_360),
.A2(n_338),
.B1(n_341),
.B2(n_355),
.Y(n_378)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_378),
.Y(n_394)
);

AOI22xp5_ASAP7_75t_L g397 ( 
.A1(n_379),
.A2(n_390),
.B1(n_369),
.B2(n_359),
.Y(n_397)
);

MAJIxp5_ASAP7_75t_L g381 ( 
.A(n_372),
.B(n_340),
.C(n_357),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_381),
.B(n_382),
.Y(n_395)
);

MAJIxp5_ASAP7_75t_L g382 ( 
.A(n_372),
.B(n_347),
.C(n_74),
.Y(n_382)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_383),
.Y(n_406)
);

MAJIxp5_ASAP7_75t_L g385 ( 
.A(n_368),
.B(n_65),
.C(n_60),
.Y(n_385)
);

MAJIxp5_ASAP7_75t_L g400 ( 
.A(n_385),
.B(n_393),
.C(n_41),
.Y(n_400)
);

OAI21x1_ASAP7_75t_L g396 ( 
.A1(n_387),
.A2(n_367),
.B(n_363),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_SL g388 ( 
.A(n_365),
.B(n_16),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_L g403 ( 
.A(n_388),
.B(n_389),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_SL g389 ( 
.A(n_366),
.B(n_374),
.Y(n_389)
);

HB1xp67_ASAP7_75t_L g401 ( 
.A(n_392),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_SL g393 ( 
.A(n_368),
.B(n_7),
.Y(n_393)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_396),
.Y(n_416)
);

XNOR2xp5_ASAP7_75t_L g409 ( 
.A(n_397),
.B(n_378),
.Y(n_409)
);

OAI21xp5_ASAP7_75t_SL g398 ( 
.A1(n_381),
.A2(n_376),
.B(n_361),
.Y(n_398)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_398),
.Y(n_418)
);

AND2x2_ASAP7_75t_L g399 ( 
.A(n_379),
.B(n_377),
.Y(n_399)
);

CKINVDCx14_ASAP7_75t_R g408 ( 
.A(n_399),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_SL g413 ( 
.A(n_400),
.B(n_405),
.Y(n_413)
);

HB1xp67_ASAP7_75t_L g402 ( 
.A(n_383),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_402),
.B(n_90),
.Y(n_417)
);

INVx13_ASAP7_75t_L g404 ( 
.A(n_386),
.Y(n_404)
);

NOR2xp33_ASAP7_75t_L g414 ( 
.A(n_404),
.B(n_13),
.Y(n_414)
);

MAJIxp5_ASAP7_75t_L g405 ( 
.A(n_380),
.B(n_88),
.C(n_87),
.Y(n_405)
);

INVxp67_ASAP7_75t_L g407 ( 
.A(n_399),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_407),
.B(n_411),
.Y(n_422)
);

XOR2xp5_ASAP7_75t_L g420 ( 
.A(n_409),
.B(n_417),
.Y(n_420)
);

MAJIxp5_ASAP7_75t_L g410 ( 
.A(n_395),
.B(n_391),
.C(n_382),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_SL g425 ( 
.A(n_410),
.B(n_412),
.Y(n_425)
);

OAI21xp5_ASAP7_75t_L g411 ( 
.A1(n_402),
.A2(n_384),
.B(n_385),
.Y(n_411)
);

OAI21xp5_ASAP7_75t_SL g412 ( 
.A1(n_406),
.A2(n_390),
.B(n_15),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_SL g426 ( 
.A(n_414),
.B(n_415),
.Y(n_426)
);

OAI22xp5_ASAP7_75t_SL g415 ( 
.A1(n_394),
.A2(n_95),
.B1(n_67),
.B2(n_83),
.Y(n_415)
);

XNOR2xp5_ASAP7_75t_L g419 ( 
.A(n_409),
.B(n_403),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_419),
.B(n_423),
.Y(n_433)
);

AOI322xp5_ASAP7_75t_L g421 ( 
.A1(n_407),
.A2(n_404),
.A3(n_401),
.B1(n_34),
.B2(n_11),
.C1(n_6),
.C2(n_7),
.Y(n_421)
);

OAI321xp33_ASAP7_75t_L g428 ( 
.A1(n_421),
.A2(n_408),
.A3(n_8),
.B1(n_15),
.B2(n_6),
.C(n_413),
.Y(n_428)
);

NOR2xp33_ASAP7_75t_L g423 ( 
.A(n_410),
.B(n_401),
.Y(n_423)
);

XNOR2xp5_ASAP7_75t_L g424 ( 
.A(n_411),
.B(n_7),
.Y(n_424)
);

XOR2xp5_ASAP7_75t_L g431 ( 
.A(n_424),
.B(n_0),
.Y(n_431)
);

MAJIxp5_ASAP7_75t_L g427 ( 
.A(n_418),
.B(n_46),
.C(n_61),
.Y(n_427)
);

NOR2xp33_ASAP7_75t_L g432 ( 
.A(n_427),
.B(n_0),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_428),
.B(n_431),
.Y(n_437)
);

AOI21xp5_ASAP7_75t_L g429 ( 
.A1(n_425),
.A2(n_416),
.B(n_8),
.Y(n_429)
);

OAI21xp5_ASAP7_75t_L g435 ( 
.A1(n_429),
.A2(n_430),
.B(n_4),
.Y(n_435)
);

AOI21x1_ASAP7_75t_L g430 ( 
.A1(n_422),
.A2(n_15),
.B(n_3),
.Y(n_430)
);

NOR2xp33_ASAP7_75t_L g436 ( 
.A(n_432),
.B(n_420),
.Y(n_436)
);

AOI322xp5_ASAP7_75t_L g434 ( 
.A1(n_433),
.A2(n_426),
.A3(n_420),
.B1(n_427),
.B2(n_4),
.C1(n_3),
.C2(n_5),
.Y(n_434)
);

NOR3xp33_ASAP7_75t_L g439 ( 
.A(n_434),
.B(n_5),
.C(n_437),
.Y(n_439)
);

MAJIxp5_ASAP7_75t_L g438 ( 
.A(n_435),
.B(n_436),
.C(n_4),
.Y(n_438)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_438),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_440),
.Y(n_441)
);

XOR2xp5_ASAP7_75t_L g442 ( 
.A(n_441),
.B(n_439),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_SL g443 ( 
.A(n_442),
.B(n_5),
.Y(n_443)
);


endmodule