module fake_jpeg_2708_n_638 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_638);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_638;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_182;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_620;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_417;
wire n_362;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_637;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_615;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_599;
wire n_239;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

INVx11_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

INVx8_ASAP7_75t_SL g24 ( 
.A(n_6),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_19),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

BUFx10_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_14),
.Y(n_32)
);

CKINVDCx16_ASAP7_75t_R g33 ( 
.A(n_3),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_3),
.Y(n_34)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_8),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_3),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_0),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_8),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_5),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_2),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_0),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_15),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_5),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_18),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_14),
.B(n_15),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_15),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_4),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_19),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_4),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_19),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_9),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_16),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_3),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_15),
.Y(n_56)
);

INVxp33_ASAP7_75t_L g57 ( 
.A(n_17),
.Y(n_57)
);

BUFx12_ASAP7_75t_L g58 ( 
.A(n_24),
.Y(n_58)
);

CKINVDCx6p67_ASAP7_75t_R g133 ( 
.A(n_58),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_50),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_59),
.B(n_82),
.Y(n_138)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_20),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g173 ( 
.A(n_60),
.Y(n_173)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_28),
.Y(n_61)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_61),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_50),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g180 ( 
.A(n_62),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_50),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g190 ( 
.A(n_63),
.Y(n_190)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_50),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g197 ( 
.A(n_64),
.Y(n_197)
);

HB1xp67_ASAP7_75t_L g65 ( 
.A(n_28),
.Y(n_65)
);

HB1xp67_ASAP7_75t_L g136 ( 
.A(n_65),
.Y(n_136)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_28),
.Y(n_66)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_66),
.Y(n_137)
);

BUFx5_ASAP7_75t_L g67 ( 
.A(n_24),
.Y(n_67)
);

INVx4_ASAP7_75t_L g132 ( 
.A(n_67),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_25),
.B(n_18),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_68),
.B(n_89),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_20),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g218 ( 
.A(n_69),
.Y(n_218)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_20),
.Y(n_70)
);

INVx6_ASAP7_75t_L g148 ( 
.A(n_70),
.Y(n_148)
);

BUFx12f_ASAP7_75t_L g71 ( 
.A(n_35),
.Y(n_71)
);

INVx5_ASAP7_75t_L g135 ( 
.A(n_71),
.Y(n_135)
);

BUFx12_ASAP7_75t_L g72 ( 
.A(n_57),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g188 ( 
.A(n_72),
.Y(n_188)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_53),
.Y(n_73)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_73),
.Y(n_143)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_53),
.Y(n_74)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_74),
.Y(n_146)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_21),
.Y(n_75)
);

BUFx2_ASAP7_75t_L g209 ( 
.A(n_75),
.Y(n_209)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_53),
.Y(n_76)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_76),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_20),
.Y(n_77)
);

INVx6_ASAP7_75t_L g150 ( 
.A(n_77),
.Y(n_150)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_21),
.Y(n_78)
);

INVx2_ASAP7_75t_SL g162 ( 
.A(n_78),
.Y(n_162)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_21),
.Y(n_79)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_79),
.Y(n_142)
);

INVx6_ASAP7_75t_SL g80 ( 
.A(n_29),
.Y(n_80)
);

INVx8_ASAP7_75t_L g178 ( 
.A(n_80),
.Y(n_178)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_26),
.Y(n_81)
);

INVx3_ASAP7_75t_L g152 ( 
.A(n_81),
.Y(n_152)
);

CKINVDCx14_ASAP7_75t_R g82 ( 
.A(n_47),
.Y(n_82)
);

INVx8_ASAP7_75t_L g83 ( 
.A(n_22),
.Y(n_83)
);

INVx5_ASAP7_75t_L g145 ( 
.A(n_83),
.Y(n_145)
);

BUFx5_ASAP7_75t_L g84 ( 
.A(n_34),
.Y(n_84)
);

INVx4_ASAP7_75t_L g140 ( 
.A(n_84),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_47),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_85),
.B(n_86),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_39),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_36),
.Y(n_87)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_87),
.Y(n_147)
);

INVx2_ASAP7_75t_SL g88 ( 
.A(n_22),
.Y(n_88)
);

INVx4_ASAP7_75t_L g144 ( 
.A(n_88),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_25),
.B(n_0),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_46),
.B(n_52),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_90),
.B(n_93),
.Y(n_174)
);

INVx5_ASAP7_75t_L g91 ( 
.A(n_26),
.Y(n_91)
);

INVx4_ASAP7_75t_L g158 ( 
.A(n_91),
.Y(n_158)
);

BUFx5_ASAP7_75t_L g92 ( 
.A(n_34),
.Y(n_92)
);

INVx4_ASAP7_75t_L g163 ( 
.A(n_92),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_46),
.B(n_1),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_39),
.Y(n_94)
);

INVx5_ASAP7_75t_L g165 ( 
.A(n_94),
.Y(n_165)
);

INVx11_ASAP7_75t_L g95 ( 
.A(n_22),
.Y(n_95)
);

INVx4_ASAP7_75t_L g175 ( 
.A(n_95),
.Y(n_175)
);

INVx3_ASAP7_75t_SL g96 ( 
.A(n_35),
.Y(n_96)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_96),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_52),
.B(n_1),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_97),
.B(n_98),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_32),
.B(n_17),
.Y(n_98)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_36),
.Y(n_99)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_99),
.Y(n_149)
);

INVx2_ASAP7_75t_R g100 ( 
.A(n_33),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_100),
.B(n_45),
.Y(n_155)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_36),
.Y(n_101)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_101),
.Y(n_186)
);

INVx8_ASAP7_75t_L g102 ( 
.A(n_22),
.Y(n_102)
);

INVx5_ASAP7_75t_L g210 ( 
.A(n_102),
.Y(n_210)
);

INVx5_ASAP7_75t_L g103 ( 
.A(n_26),
.Y(n_103)
);

INVx4_ASAP7_75t_L g181 ( 
.A(n_103),
.Y(n_181)
);

INVx13_ASAP7_75t_L g104 ( 
.A(n_33),
.Y(n_104)
);

INVx5_ASAP7_75t_L g211 ( 
.A(n_104),
.Y(n_211)
);

BUFx16f_ASAP7_75t_L g105 ( 
.A(n_29),
.Y(n_105)
);

INVx5_ASAP7_75t_L g214 ( 
.A(n_105),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_32),
.B(n_2),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_106),
.B(n_109),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_39),
.Y(n_107)
);

INVx5_ASAP7_75t_L g215 ( 
.A(n_107),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_56),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_108),
.B(n_111),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_42),
.B(n_2),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_42),
.B(n_2),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_110),
.B(n_5),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_39),
.Y(n_111)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_35),
.Y(n_112)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_112),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_55),
.Y(n_113)
);

INVx5_ASAP7_75t_L g224 ( 
.A(n_113),
.Y(n_224)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_38),
.Y(n_114)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_114),
.Y(n_169)
);

INVx5_ASAP7_75t_L g115 ( 
.A(n_49),
.Y(n_115)
);

INVx4_ASAP7_75t_L g194 ( 
.A(n_115),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_55),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_116),
.B(n_117),
.Y(n_172)
);

OR2x2_ASAP7_75t_L g117 ( 
.A(n_38),
.B(n_4),
.Y(n_117)
);

INVx8_ASAP7_75t_L g118 ( 
.A(n_22),
.Y(n_118)
);

INVx4_ASAP7_75t_L g204 ( 
.A(n_118),
.Y(n_204)
);

BUFx12f_ASAP7_75t_L g119 ( 
.A(n_38),
.Y(n_119)
);

INVx4_ASAP7_75t_L g220 ( 
.A(n_119),
.Y(n_220)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_55),
.Y(n_120)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_120),
.Y(n_177)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_27),
.Y(n_121)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_121),
.Y(n_199)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_49),
.Y(n_122)
);

INVx3_ASAP7_75t_L g157 ( 
.A(n_122),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_56),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_123),
.B(n_124),
.Y(n_212)
);

AND2x2_ASAP7_75t_L g124 ( 
.A(n_22),
.B(n_4),
.Y(n_124)
);

INVx8_ASAP7_75t_L g125 ( 
.A(n_55),
.Y(n_125)
);

INVx3_ASAP7_75t_L g183 ( 
.A(n_125),
.Y(n_183)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_27),
.Y(n_126)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_126),
.Y(n_203)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_49),
.Y(n_127)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_127),
.Y(n_179)
);

BUFx10_ASAP7_75t_L g128 ( 
.A(n_29),
.Y(n_128)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_128),
.Y(n_182)
);

BUFx3_ASAP7_75t_L g129 ( 
.A(n_56),
.Y(n_129)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_129),
.Y(n_195)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_56),
.Y(n_130)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_130),
.Y(n_196)
);

A2O1A1Ixp33_ASAP7_75t_L g151 ( 
.A1(n_100),
.A2(n_45),
.B(n_51),
.C(n_48),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_151),
.B(n_168),
.Y(n_248)
);

AOI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_80),
.A2(n_23),
.B1(n_31),
.B2(n_41),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g241 ( 
.A1(n_153),
.A2(n_154),
.B1(n_156),
.B2(n_159),
.Y(n_241)
);

AOI22xp33_ASAP7_75t_SL g154 ( 
.A1(n_88),
.A2(n_23),
.B1(n_31),
.B2(n_41),
.Y(n_154)
);

OR2x2_ASAP7_75t_L g277 ( 
.A(n_155),
.B(n_206),
.Y(n_277)
);

AOI22xp33_ASAP7_75t_SL g156 ( 
.A1(n_105),
.A2(n_31),
.B1(n_23),
.B2(n_54),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_L g159 ( 
.A1(n_130),
.A2(n_77),
.B1(n_107),
.B2(n_94),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_SL g161 ( 
.A(n_124),
.B(n_51),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_SL g244 ( 
.A(n_161),
.B(n_167),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_105),
.Y(n_167)
);

A2O1A1Ixp33_ASAP7_75t_L g168 ( 
.A1(n_117),
.A2(n_48),
.B(n_54),
.C(n_41),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_SL g170 ( 
.A1(n_95),
.A2(n_54),
.B1(n_44),
.B2(n_43),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g267 ( 
.A1(n_170),
.A2(n_185),
.B1(n_192),
.B2(n_200),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_60),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_SL g295 ( 
.A(n_171),
.B(n_189),
.Y(n_295)
);

OAI22xp33_ASAP7_75t_SL g184 ( 
.A1(n_62),
.A2(n_64),
.B1(n_63),
.B2(n_73),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_184),
.A2(n_208),
.B1(n_125),
.B2(n_83),
.Y(n_238)
);

AOI22xp33_ASAP7_75t_SL g185 ( 
.A1(n_78),
.A2(n_44),
.B1(n_43),
.B2(n_40),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_SL g189 ( 
.A(n_75),
.B(n_44),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_61),
.B(n_74),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g288 ( 
.A(n_191),
.B(n_193),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_69),
.A2(n_43),
.B1(n_40),
.B2(n_37),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_112),
.B(n_40),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_198),
.B(n_217),
.Y(n_250)
);

AOI22xp33_ASAP7_75t_L g200 ( 
.A1(n_70),
.A2(n_37),
.B1(n_30),
.B2(n_27),
.Y(n_200)
);

AOI22xp33_ASAP7_75t_SL g201 ( 
.A1(n_79),
.A2(n_37),
.B1(n_30),
.B2(n_29),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g286 ( 
.A1(n_201),
.A2(n_205),
.B1(n_216),
.B2(n_211),
.Y(n_286)
);

AND2x2_ASAP7_75t_SL g202 ( 
.A(n_114),
.B(n_30),
.Y(n_202)
);

AND2x2_ASAP7_75t_L g245 ( 
.A(n_202),
.B(n_11),
.Y(n_245)
);

AOI22xp33_ASAP7_75t_SL g205 ( 
.A1(n_81),
.A2(n_29),
.B1(n_34),
.B2(n_7),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_SL g206 ( 
.A(n_91),
.B(n_5),
.Y(n_206)
);

AND2x4_ASAP7_75t_L g207 ( 
.A(n_122),
.B(n_29),
.Y(n_207)
);

INVx1_ASAP7_75t_SL g230 ( 
.A(n_207),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_113),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_208)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_96),
.Y(n_213)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_213),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_L g216 ( 
.A1(n_120),
.A2(n_6),
.B1(n_7),
.B2(n_9),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_127),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_103),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_219),
.B(n_223),
.Y(n_276)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_71),
.Y(n_221)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_221),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_SL g222 ( 
.A(n_115),
.B(n_9),
.Y(n_222)
);

OR2x2_ASAP7_75t_L g280 ( 
.A(n_222),
.B(n_226),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_71),
.B(n_17),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_129),
.B(n_9),
.C(n_10),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_225),
.B(n_104),
.C(n_72),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_119),
.B(n_10),
.Y(n_226)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_119),
.Y(n_227)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_227),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_202),
.B(n_10),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_228),
.B(n_232),
.Y(n_322)
);

INVxp67_ASAP7_75t_L g229 ( 
.A(n_133),
.Y(n_229)
);

INVxp67_ASAP7_75t_L g314 ( 
.A(n_229),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_231),
.B(n_258),
.C(n_266),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_212),
.B(n_10),
.Y(n_232)
);

OR2x2_ASAP7_75t_SL g233 ( 
.A(n_151),
.B(n_72),
.Y(n_233)
);

CKINVDCx16_ASAP7_75t_R g325 ( 
.A(n_233),
.Y(n_325)
);

AND2x2_ASAP7_75t_SL g234 ( 
.A(n_137),
.B(n_128),
.Y(n_234)
);

INVx1_ASAP7_75t_SL g359 ( 
.A(n_234),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_136),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_SL g343 ( 
.A(n_235),
.B(n_246),
.Y(n_343)
);

INVx4_ASAP7_75t_L g236 ( 
.A(n_144),
.Y(n_236)
);

INVx3_ASAP7_75t_L g326 ( 
.A(n_236),
.Y(n_326)
);

CKINVDCx16_ASAP7_75t_R g237 ( 
.A(n_133),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g371 ( 
.A(n_237),
.B(n_229),
.Y(n_371)
);

AOI22xp5_ASAP7_75t_L g340 ( 
.A1(n_238),
.A2(n_265),
.B1(n_278),
.B2(n_282),
.Y(n_340)
);

BUFx4f_ASAP7_75t_SL g239 ( 
.A(n_133),
.Y(n_239)
);

CKINVDCx16_ASAP7_75t_R g358 ( 
.A(n_239),
.Y(n_358)
);

AOI22xp33_ASAP7_75t_SL g240 ( 
.A1(n_207),
.A2(n_118),
.B1(n_102),
.B2(n_92),
.Y(n_240)
);

INVxp67_ASAP7_75t_L g321 ( 
.A(n_240),
.Y(n_321)
);

AOI22xp33_ASAP7_75t_L g242 ( 
.A1(n_184),
.A2(n_128),
.B1(n_12),
.B2(n_13),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_L g319 ( 
.A1(n_242),
.A2(n_255),
.B1(n_291),
.B2(n_300),
.Y(n_319)
);

AOI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_207),
.A2(n_84),
.B1(n_58),
.B2(n_67),
.Y(n_243)
);

INVxp67_ASAP7_75t_L g330 ( 
.A(n_243),
.Y(n_330)
);

AOI21xp33_ASAP7_75t_L g346 ( 
.A1(n_245),
.A2(n_273),
.B(n_286),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_136),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_139),
.Y(n_247)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_247),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_168),
.B(n_11),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_249),
.B(n_251),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_176),
.B(n_11),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_144),
.Y(n_252)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_252),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_199),
.B(n_11),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_253),
.B(n_254),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_203),
.B(n_12),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_172),
.A2(n_58),
.B1(n_13),
.B2(n_16),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_196),
.Y(n_256)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_256),
.Y(n_323)
);

INVxp67_ASAP7_75t_L g257 ( 
.A(n_160),
.Y(n_257)
);

INVxp67_ASAP7_75t_L g338 ( 
.A(n_257),
.Y(n_338)
);

AND2x2_ASAP7_75t_L g258 ( 
.A(n_188),
.B(n_12),
.Y(n_258)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_147),
.Y(n_260)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_260),
.Y(n_329)
);

O2A1O1Ixp33_ASAP7_75t_SL g261 ( 
.A1(n_200),
.A2(n_16),
.B(n_17),
.C(n_159),
.Y(n_261)
);

AOI21xp5_ASAP7_75t_SL g334 ( 
.A1(n_261),
.A2(n_309),
.B(n_241),
.Y(n_334)
);

CKINVDCx16_ASAP7_75t_R g262 ( 
.A(n_209),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g363 ( 
.A(n_262),
.B(n_281),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_149),
.B(n_186),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_263),
.B(n_269),
.Y(n_348)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_164),
.Y(n_264)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_264),
.Y(n_331)
);

OAI22xp33_ASAP7_75t_SL g265 ( 
.A1(n_138),
.A2(n_16),
.B1(n_205),
.B2(n_201),
.Y(n_265)
);

AND2x2_ASAP7_75t_L g266 ( 
.A(n_188),
.B(n_146),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_134),
.B(n_143),
.Y(n_269)
);

AND2x2_ASAP7_75t_L g270 ( 
.A(n_162),
.B(n_169),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_270),
.B(n_298),
.C(n_311),
.Y(n_347)
);

INVx6_ASAP7_75t_L g271 ( 
.A(n_180),
.Y(n_271)
);

BUFx6f_ASAP7_75t_L g337 ( 
.A(n_271),
.Y(n_337)
);

AOI22xp33_ASAP7_75t_SL g273 ( 
.A1(n_140),
.A2(n_163),
.B1(n_162),
.B2(n_209),
.Y(n_273)
);

INVx3_ASAP7_75t_L g274 ( 
.A(n_178),
.Y(n_274)
);

INVx3_ASAP7_75t_L g354 ( 
.A(n_274),
.Y(n_354)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_177),
.Y(n_275)
);

INVx2_ASAP7_75t_L g342 ( 
.A(n_275),
.Y(n_342)
);

OAI22xp33_ASAP7_75t_L g278 ( 
.A1(n_185),
.A2(n_153),
.B1(n_154),
.B2(n_156),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_187),
.B(n_131),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_279),
.B(n_292),
.Y(n_357)
);

OR2x2_ASAP7_75t_L g281 ( 
.A(n_141),
.B(n_174),
.Y(n_281)
);

OAI22xp33_ASAP7_75t_SL g282 ( 
.A1(n_183),
.A2(n_170),
.B1(n_173),
.B2(n_152),
.Y(n_282)
);

BUFx3_ASAP7_75t_L g283 ( 
.A(n_214),
.Y(n_283)
);

BUFx6f_ASAP7_75t_L g352 ( 
.A(n_283),
.Y(n_352)
);

INVx8_ASAP7_75t_L g284 ( 
.A(n_218),
.Y(n_284)
);

INVx2_ASAP7_75t_L g362 ( 
.A(n_284),
.Y(n_362)
);

BUFx6f_ASAP7_75t_L g285 ( 
.A(n_180),
.Y(n_285)
);

INVx8_ASAP7_75t_L g345 ( 
.A(n_285),
.Y(n_345)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_165),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g366 ( 
.A(n_287),
.B(n_307),
.Y(n_366)
);

BUFx2_ASAP7_75t_SL g289 ( 
.A(n_179),
.Y(n_289)
);

INVx2_ASAP7_75t_L g368 ( 
.A(n_289),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_178),
.B(n_157),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_SL g351 ( 
.A(n_290),
.B(n_294),
.Y(n_351)
);

OAI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_173),
.A2(n_148),
.B1(n_150),
.B2(n_166),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_142),
.B(n_195),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_204),
.Y(n_293)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_293),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_220),
.B(n_181),
.Y(n_294)
);

FAx1_ASAP7_75t_SL g296 ( 
.A(n_140),
.B(n_163),
.CI(n_182),
.CON(n_296),
.SN(n_296)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_296),
.B(n_297),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_220),
.B(n_181),
.Y(n_297)
);

AND2x2_ASAP7_75t_L g298 ( 
.A(n_158),
.B(n_194),
.Y(n_298)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_158),
.Y(n_299)
);

INVx2_ASAP7_75t_SL g341 ( 
.A(n_299),
.Y(n_341)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_218),
.A2(n_190),
.B1(n_197),
.B2(n_224),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_194),
.B(n_135),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_301),
.B(n_310),
.Y(n_315)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_148),
.Y(n_302)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_302),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_150),
.B(n_197),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_303),
.B(n_300),
.Y(n_365)
);

BUFx12f_ASAP7_75t_L g304 ( 
.A(n_190),
.Y(n_304)
);

INVx13_ASAP7_75t_L g353 ( 
.A(n_304),
.Y(n_353)
);

INVx2_ASAP7_75t_L g305 ( 
.A(n_215),
.Y(n_305)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_305),
.Y(n_355)
);

INVx5_ASAP7_75t_L g306 ( 
.A(n_145),
.Y(n_306)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_306),
.Y(n_360)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_210),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_204),
.Y(n_308)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_308),
.Y(n_364)
);

O2A1O1Ixp33_ASAP7_75t_SL g309 ( 
.A1(n_132),
.A2(n_175),
.B(n_168),
.C(n_200),
.Y(n_309)
);

INVxp67_ASAP7_75t_L g310 ( 
.A(n_132),
.Y(n_310)
);

AND2x2_ASAP7_75t_L g311 ( 
.A(n_175),
.B(n_100),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_244),
.B(n_264),
.Y(n_317)
);

CKINVDCx14_ASAP7_75t_R g376 ( 
.A(n_317),
.Y(n_376)
);

OAI22xp5_ASAP7_75t_SL g318 ( 
.A1(n_238),
.A2(n_248),
.B1(n_288),
.B2(n_230),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_L g377 ( 
.A1(n_318),
.A2(n_332),
.B1(n_333),
.B2(n_361),
.Y(n_377)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_263),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_SL g386 ( 
.A(n_320),
.B(n_324),
.Y(n_386)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_270),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_276),
.B(n_295),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g375 ( 
.A(n_327),
.B(n_344),
.Y(n_375)
);

OAI22xp5_ASAP7_75t_SL g332 ( 
.A1(n_230),
.A2(n_228),
.B1(n_309),
.B2(n_245),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_SL g333 ( 
.A1(n_309),
.A2(n_245),
.B1(n_249),
.B2(n_280),
.Y(n_333)
);

AND2x2_ASAP7_75t_L g401 ( 
.A(n_334),
.B(n_371),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_281),
.B(n_250),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g349 ( 
.A(n_270),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_SL g412 ( 
.A(n_349),
.B(n_359),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_L g356 ( 
.A(n_277),
.B(n_260),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_L g391 ( 
.A(n_356),
.B(n_370),
.Y(n_391)
);

OAI22xp5_ASAP7_75t_SL g361 ( 
.A1(n_280),
.A2(n_233),
.B1(n_261),
.B2(n_267),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_365),
.B(n_369),
.Y(n_373)
);

OAI22xp5_ASAP7_75t_L g367 ( 
.A1(n_231),
.A2(n_254),
.B1(n_253),
.B2(n_303),
.Y(n_367)
);

AOI22xp5_ASAP7_75t_L g389 ( 
.A1(n_367),
.A2(n_266),
.B1(n_298),
.B2(n_293),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_251),
.B(n_269),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_L g370 ( 
.A(n_277),
.B(n_279),
.Y(n_370)
);

NOR2x1p5_ASAP7_75t_L g372 ( 
.A(n_325),
.B(n_296),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_372),
.B(n_383),
.Y(n_435)
);

OAI21xp5_ASAP7_75t_L g374 ( 
.A1(n_312),
.A2(n_311),
.B(n_255),
.Y(n_374)
);

OAI21xp5_ASAP7_75t_L g449 ( 
.A1(n_374),
.A2(n_378),
.B(n_381),
.Y(n_449)
);

OAI21xp5_ASAP7_75t_SL g378 ( 
.A1(n_330),
.A2(n_243),
.B(n_311),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_313),
.Y(n_379)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_379),
.Y(n_419)
);

OAI22xp5_ASAP7_75t_SL g380 ( 
.A1(n_340),
.A2(n_261),
.B1(n_278),
.B2(n_234),
.Y(n_380)
);

AOI22xp5_ASAP7_75t_L g427 ( 
.A1(n_380),
.A2(n_387),
.B1(n_390),
.B2(n_395),
.Y(n_427)
);

OAI21xp5_ASAP7_75t_L g381 ( 
.A1(n_334),
.A2(n_258),
.B(n_232),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_313),
.Y(n_382)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_382),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_336),
.B(n_292),
.Y(n_383)
);

AOI21xp5_ASAP7_75t_L g384 ( 
.A1(n_346),
.A2(n_296),
.B(n_274),
.Y(n_384)
);

INVxp67_ASAP7_75t_L g436 ( 
.A(n_384),
.Y(n_436)
);

AOI21xp5_ASAP7_75t_SL g385 ( 
.A1(n_330),
.A2(n_258),
.B(n_247),
.Y(n_385)
);

OAI21xp33_ASAP7_75t_L g446 ( 
.A1(n_385),
.A2(n_415),
.B(n_314),
.Y(n_446)
);

OAI22xp5_ASAP7_75t_SL g387 ( 
.A1(n_340),
.A2(n_234),
.B1(n_302),
.B2(n_271),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_SL g388 ( 
.A(n_357),
.B(n_256),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_SL g432 ( 
.A(n_388),
.B(n_322),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_389),
.B(n_393),
.Y(n_437)
);

AOI22xp5_ASAP7_75t_L g390 ( 
.A1(n_361),
.A2(n_291),
.B1(n_266),
.B2(n_275),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_L g392 ( 
.A(n_331),
.B(n_239),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_SL g424 ( 
.A(n_392),
.B(n_399),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_336),
.B(n_308),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_329),
.Y(n_394)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_394),
.Y(n_425)
);

AOI22xp5_ASAP7_75t_L g395 ( 
.A1(n_332),
.A2(n_298),
.B1(n_305),
.B2(n_284),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_329),
.Y(n_396)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_396),
.Y(n_433)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_323),
.Y(n_397)
);

INVx2_ASAP7_75t_SL g420 ( 
.A(n_397),
.Y(n_420)
);

AOI32xp33_ASAP7_75t_L g398 ( 
.A1(n_357),
.A2(n_236),
.A3(n_299),
.B1(n_252),
.B2(n_259),
.Y(n_398)
);

AOI322xp5_ASAP7_75t_L g448 ( 
.A1(n_398),
.A2(n_353),
.A3(n_352),
.B1(n_338),
.B2(n_337),
.C1(n_355),
.C2(n_350),
.Y(n_448)
);

NOR2xp33_ASAP7_75t_SL g399 ( 
.A(n_320),
.B(n_268),
.Y(n_399)
);

AOI22xp5_ASAP7_75t_L g400 ( 
.A1(n_318),
.A2(n_285),
.B1(n_259),
.B2(n_306),
.Y(n_400)
);

AOI22xp5_ASAP7_75t_L g434 ( 
.A1(n_400),
.A2(n_408),
.B1(n_417),
.B2(n_314),
.Y(n_434)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_323),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_SL g429 ( 
.A(n_402),
.B(n_409),
.Y(n_429)
);

MAJIxp5_ASAP7_75t_L g403 ( 
.A(n_328),
.B(n_257),
.C(n_268),
.Y(n_403)
);

MAJIxp5_ASAP7_75t_L g444 ( 
.A(n_403),
.B(n_406),
.C(n_316),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_348),
.B(n_239),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_404),
.B(n_407),
.Y(n_443)
);

HB1xp67_ASAP7_75t_L g405 ( 
.A(n_360),
.Y(n_405)
);

CKINVDCx20_ASAP7_75t_R g430 ( 
.A(n_405),
.Y(n_430)
);

MAJIxp5_ASAP7_75t_L g406 ( 
.A(n_328),
.B(n_367),
.C(n_348),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_369),
.B(n_272),
.Y(n_407)
);

AOI22xp5_ASAP7_75t_L g408 ( 
.A1(n_365),
.A2(n_272),
.B1(n_310),
.B2(n_283),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_L g409 ( 
.A(n_331),
.B(n_304),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_339),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_410),
.B(n_413),
.Y(n_452)
);

NOR2xp33_ASAP7_75t_SL g411 ( 
.A(n_335),
.B(n_304),
.Y(n_411)
);

OR2x2_ASAP7_75t_L g423 ( 
.A(n_411),
.B(n_412),
.Y(n_423)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_339),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_364),
.Y(n_414)
);

AOI22xp33_ASAP7_75t_SL g445 ( 
.A1(n_414),
.A2(n_416),
.B1(n_341),
.B2(n_360),
.Y(n_445)
);

AND2x2_ASAP7_75t_L g415 ( 
.A(n_359),
.B(n_304),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_364),
.Y(n_416)
);

OAI22xp5_ASAP7_75t_SL g417 ( 
.A1(n_335),
.A2(n_324),
.B1(n_349),
.B2(n_321),
.Y(n_417)
);

AO22x1_ASAP7_75t_SL g418 ( 
.A1(n_333),
.A2(n_319),
.B1(n_347),
.B2(n_316),
.Y(n_418)
);

AOI22xp33_ASAP7_75t_L g441 ( 
.A1(n_418),
.A2(n_322),
.B1(n_343),
.B2(n_315),
.Y(n_441)
);

CKINVDCx16_ASAP7_75t_R g422 ( 
.A(n_401),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_SL g465 ( 
.A(n_422),
.B(n_428),
.Y(n_465)
);

XOR2xp5_ASAP7_75t_L g426 ( 
.A(n_406),
.B(n_347),
.Y(n_426)
);

MAJIxp5_ASAP7_75t_L g471 ( 
.A(n_426),
.B(n_440),
.C(n_444),
.Y(n_471)
);

CKINVDCx16_ASAP7_75t_R g428 ( 
.A(n_401),
.Y(n_428)
);

CKINVDCx16_ASAP7_75t_R g431 ( 
.A(n_404),
.Y(n_431)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_431),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_432),
.B(n_445),
.Y(n_459)
);

OAI22xp5_ASAP7_75t_L g474 ( 
.A1(n_434),
.A2(n_438),
.B1(n_441),
.B2(n_442),
.Y(n_474)
);

AOI22xp5_ASAP7_75t_L g438 ( 
.A1(n_380),
.A2(n_319),
.B1(n_321),
.B2(n_351),
.Y(n_438)
);

OR2x2_ASAP7_75t_L g439 ( 
.A(n_386),
.B(n_351),
.Y(n_439)
);

OAI22xp33_ASAP7_75t_SL g468 ( 
.A1(n_439),
.A2(n_389),
.B1(n_372),
.B2(n_374),
.Y(n_468)
);

XNOR2xp5_ASAP7_75t_L g440 ( 
.A(n_383),
.B(n_403),
.Y(n_440)
);

AOI22xp5_ASAP7_75t_L g442 ( 
.A1(n_373),
.A2(n_366),
.B1(n_363),
.B2(n_354),
.Y(n_442)
);

OAI21xp5_ASAP7_75t_L g478 ( 
.A1(n_446),
.A2(n_448),
.B(n_451),
.Y(n_478)
);

MAJIxp5_ASAP7_75t_L g447 ( 
.A(n_377),
.B(n_354),
.C(n_355),
.Y(n_447)
);

MAJIxp5_ASAP7_75t_L g472 ( 
.A(n_447),
.B(n_454),
.C(n_455),
.Y(n_472)
);

BUFx3_ASAP7_75t_L g450 ( 
.A(n_395),
.Y(n_450)
);

NOR2xp33_ASAP7_75t_L g479 ( 
.A(n_450),
.B(n_456),
.Y(n_479)
);

AOI22xp5_ASAP7_75t_SL g451 ( 
.A1(n_401),
.A2(n_358),
.B1(n_362),
.B2(n_338),
.Y(n_451)
);

AOI22xp5_ASAP7_75t_L g453 ( 
.A1(n_373),
.A2(n_362),
.B1(n_337),
.B2(n_350),
.Y(n_453)
);

OAI22xp5_ASAP7_75t_L g490 ( 
.A1(n_453),
.A2(n_341),
.B1(n_337),
.B2(n_345),
.Y(n_490)
);

XNOR2xp5_ASAP7_75t_L g454 ( 
.A(n_393),
.B(n_342),
.Y(n_454)
);

MAJIxp5_ASAP7_75t_L g455 ( 
.A(n_377),
.B(n_326),
.C(n_342),
.Y(n_455)
);

CKINVDCx16_ASAP7_75t_R g456 ( 
.A(n_375),
.Y(n_456)
);

XOR2xp5_ASAP7_75t_L g457 ( 
.A(n_418),
.B(n_368),
.Y(n_457)
);

MAJIxp5_ASAP7_75t_L g473 ( 
.A(n_457),
.B(n_458),
.C(n_415),
.Y(n_473)
);

MAJIxp5_ASAP7_75t_L g458 ( 
.A(n_418),
.B(n_326),
.C(n_368),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_443),
.B(n_388),
.Y(n_460)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_460),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_443),
.B(n_407),
.Y(n_461)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_461),
.Y(n_516)
);

AOI22xp5_ASAP7_75t_L g462 ( 
.A1(n_438),
.A2(n_384),
.B1(n_417),
.B2(n_387),
.Y(n_462)
);

OAI22xp5_ASAP7_75t_L g528 ( 
.A1(n_462),
.A2(n_464),
.B1(n_480),
.B2(n_484),
.Y(n_528)
);

AOI22xp5_ASAP7_75t_L g464 ( 
.A1(n_427),
.A2(n_381),
.B1(n_390),
.B2(n_400),
.Y(n_464)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_452),
.Y(n_466)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_466),
.Y(n_502)
);

OAI32xp33_ASAP7_75t_L g467 ( 
.A1(n_437),
.A2(n_399),
.A3(n_391),
.B1(n_411),
.B2(n_372),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_467),
.B(n_475),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_SL g499 ( 
.A(n_468),
.B(n_492),
.Y(n_499)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_452),
.Y(n_469)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_469),
.Y(n_517)
);

CKINVDCx20_ASAP7_75t_R g470 ( 
.A(n_429),
.Y(n_470)
);

CKINVDCx5p33_ASAP7_75t_R g503 ( 
.A(n_470),
.Y(n_503)
);

HB1xp67_ASAP7_75t_L g523 ( 
.A(n_473),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_431),
.B(n_394),
.Y(n_475)
);

CKINVDCx20_ASAP7_75t_R g476 ( 
.A(n_439),
.Y(n_476)
);

INVxp67_ASAP7_75t_SL g506 ( 
.A(n_476),
.Y(n_506)
);

XOR2xp5_ASAP7_75t_L g477 ( 
.A(n_426),
.B(n_385),
.Y(n_477)
);

MAJIxp5_ASAP7_75t_L g496 ( 
.A(n_477),
.B(n_481),
.C(n_485),
.Y(n_496)
);

AOI22xp5_ASAP7_75t_L g480 ( 
.A1(n_427),
.A2(n_396),
.B1(n_382),
.B2(n_379),
.Y(n_480)
);

XOR2xp5_ASAP7_75t_L g481 ( 
.A(n_440),
.B(n_444),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_454),
.B(n_402),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g511 ( 
.A(n_482),
.B(n_486),
.Y(n_511)
);

XNOR2x1_ASAP7_75t_L g483 ( 
.A(n_457),
.B(n_415),
.Y(n_483)
);

XNOR2xp5_ASAP7_75t_SL g497 ( 
.A(n_483),
.B(n_435),
.Y(n_497)
);

AOI22xp5_ASAP7_75t_L g484 ( 
.A1(n_458),
.A2(n_408),
.B1(n_414),
.B2(n_413),
.Y(n_484)
);

MAJIxp5_ASAP7_75t_L g485 ( 
.A(n_449),
.B(n_378),
.C(n_397),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g486 ( 
.A(n_424),
.B(n_410),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_430),
.B(n_416),
.Y(n_487)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_487),
.Y(n_521)
);

XOR2xp5_ASAP7_75t_L g488 ( 
.A(n_449),
.B(n_398),
.Y(n_488)
);

MAJIxp5_ASAP7_75t_L g504 ( 
.A(n_488),
.B(n_493),
.C(n_494),
.Y(n_504)
);

NOR2xp33_ASAP7_75t_L g489 ( 
.A(n_442),
.B(n_376),
.Y(n_489)
);

CKINVDCx14_ASAP7_75t_R g501 ( 
.A(n_489),
.Y(n_501)
);

AOI22xp5_ASAP7_75t_L g509 ( 
.A1(n_490),
.A2(n_420),
.B1(n_419),
.B2(n_421),
.Y(n_509)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_420),
.Y(n_491)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_491),
.Y(n_527)
);

NOR2xp33_ASAP7_75t_L g492 ( 
.A(n_432),
.B(n_352),
.Y(n_492)
);

MAJIxp5_ASAP7_75t_L g493 ( 
.A(n_437),
.B(n_341),
.C(n_352),
.Y(n_493)
);

MAJIxp5_ASAP7_75t_L g494 ( 
.A(n_447),
.B(n_353),
.C(n_345),
.Y(n_494)
);

MAJIxp5_ASAP7_75t_L g495 ( 
.A(n_436),
.B(n_435),
.C(n_455),
.Y(n_495)
);

MAJIxp5_ASAP7_75t_L g508 ( 
.A(n_495),
.B(n_430),
.C(n_453),
.Y(n_508)
);

XNOR2x1_ASAP7_75t_L g539 ( 
.A(n_497),
.B(n_482),
.Y(n_539)
);

AOI21xp5_ASAP7_75t_L g498 ( 
.A1(n_488),
.A2(n_436),
.B(n_423),
.Y(n_498)
);

INVxp67_ASAP7_75t_L g556 ( 
.A(n_498),
.Y(n_556)
);

OAI22xp5_ASAP7_75t_SL g500 ( 
.A1(n_462),
.A2(n_434),
.B1(n_450),
.B2(n_423),
.Y(n_500)
);

AOI22xp5_ASAP7_75t_L g544 ( 
.A1(n_500),
.A2(n_512),
.B1(n_518),
.B2(n_478),
.Y(n_544)
);

XNOR2xp5_ASAP7_75t_L g507 ( 
.A(n_477),
.B(n_451),
.Y(n_507)
);

XOR2xp5_ASAP7_75t_L g551 ( 
.A(n_507),
.B(n_520),
.Y(n_551)
);

MAJIxp5_ASAP7_75t_L g530 ( 
.A(n_508),
.B(n_513),
.C(n_515),
.Y(n_530)
);

OAI22xp5_ASAP7_75t_L g537 ( 
.A1(n_509),
.A2(n_491),
.B1(n_490),
.B2(n_494),
.Y(n_537)
);

INVx4_ASAP7_75t_L g510 ( 
.A(n_479),
.Y(n_510)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_510),
.Y(n_536)
);

OAI22xp5_ASAP7_75t_SL g512 ( 
.A1(n_464),
.A2(n_420),
.B1(n_419),
.B2(n_421),
.Y(n_512)
);

MAJIxp5_ASAP7_75t_L g513 ( 
.A(n_471),
.B(n_425),
.C(n_433),
.Y(n_513)
);

MAJIxp5_ASAP7_75t_L g515 ( 
.A(n_471),
.B(n_425),
.C(n_433),
.Y(n_515)
);

OAI22xp5_ASAP7_75t_SL g518 ( 
.A1(n_466),
.A2(n_469),
.B1(n_480),
.B2(n_476),
.Y(n_518)
);

OAI21xp5_ASAP7_75t_SL g519 ( 
.A1(n_459),
.A2(n_478),
.B(n_474),
.Y(n_519)
);

INVxp67_ASAP7_75t_L g540 ( 
.A(n_519),
.Y(n_540)
);

XNOR2xp5_ASAP7_75t_L g520 ( 
.A(n_481),
.B(n_485),
.Y(n_520)
);

NOR2xp33_ASAP7_75t_L g522 ( 
.A(n_470),
.B(n_486),
.Y(n_522)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_522),
.Y(n_547)
);

NOR2xp33_ASAP7_75t_L g524 ( 
.A(n_495),
.B(n_463),
.Y(n_524)
);

NOR2xp33_ASAP7_75t_L g532 ( 
.A(n_524),
.B(n_529),
.Y(n_532)
);

XOR2xp5_ASAP7_75t_L g525 ( 
.A(n_465),
.B(n_483),
.Y(n_525)
);

MAJIxp5_ASAP7_75t_L g535 ( 
.A(n_525),
.B(n_526),
.C(n_472),
.Y(n_535)
);

XOR2xp5_ASAP7_75t_L g526 ( 
.A(n_467),
.B(n_472),
.Y(n_526)
);

NOR2xp33_ASAP7_75t_L g529 ( 
.A(n_463),
.B(n_493),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g531 ( 
.A(n_503),
.B(n_475),
.Y(n_531)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_531),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_503),
.B(n_487),
.Y(n_533)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_533),
.Y(n_572)
);

OA21x2_ASAP7_75t_L g534 ( 
.A1(n_505),
.A2(n_459),
.B(n_484),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g560 ( 
.A(n_534),
.B(n_541),
.Y(n_560)
);

XNOR2xp5_ASAP7_75t_SL g573 ( 
.A(n_535),
.B(n_539),
.Y(n_573)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_537),
.Y(n_576)
);

NOR2xp33_ASAP7_75t_L g538 ( 
.A(n_513),
.B(n_460),
.Y(n_538)
);

NOR2xp33_ASAP7_75t_L g575 ( 
.A(n_538),
.B(n_543),
.Y(n_575)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_518),
.Y(n_541)
);

XNOR2xp5_ASAP7_75t_SL g542 ( 
.A(n_520),
.B(n_473),
.Y(n_542)
);

XNOR2xp5_ASAP7_75t_L g558 ( 
.A(n_542),
.B(n_555),
.Y(n_558)
);

NOR2xp33_ASAP7_75t_L g543 ( 
.A(n_515),
.B(n_461),
.Y(n_543)
);

OAI22xp5_ASAP7_75t_L g559 ( 
.A1(n_544),
.A2(n_534),
.B1(n_550),
.B2(n_540),
.Y(n_559)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_506),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_L g562 ( 
.A(n_545),
.B(n_546),
.Y(n_562)
);

OAI22xp5_ASAP7_75t_L g546 ( 
.A1(n_501),
.A2(n_505),
.B1(n_510),
.B2(n_528),
.Y(n_546)
);

MAJIxp5_ASAP7_75t_L g548 ( 
.A(n_523),
.B(n_496),
.C(n_504),
.Y(n_548)
);

MAJIxp5_ASAP7_75t_L g563 ( 
.A(n_548),
.B(n_496),
.C(n_504),
.Y(n_563)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_527),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_L g568 ( 
.A(n_549),
.B(n_553),
.Y(n_568)
);

INVxp67_ASAP7_75t_L g550 ( 
.A(n_519),
.Y(n_550)
);

NAND2x1_ASAP7_75t_SL g561 ( 
.A(n_550),
.B(n_500),
.Y(n_561)
);

OR2x2_ASAP7_75t_L g552 ( 
.A(n_499),
.B(n_502),
.Y(n_552)
);

CKINVDCx20_ASAP7_75t_R g564 ( 
.A(n_552),
.Y(n_564)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_521),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_511),
.B(n_514),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_L g569 ( 
.A(n_554),
.B(n_514),
.Y(n_569)
);

XNOR2xp5_ASAP7_75t_SL g555 ( 
.A(n_526),
.B(n_497),
.Y(n_555)
);

AOI22xp5_ASAP7_75t_L g581 ( 
.A1(n_559),
.A2(n_574),
.B1(n_541),
.B2(n_572),
.Y(n_581)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_561),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_SL g590 ( 
.A(n_563),
.B(n_567),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_SL g565 ( 
.A(n_547),
.B(n_511),
.Y(n_565)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_565),
.Y(n_588)
);

INVx13_ASAP7_75t_L g566 ( 
.A(n_545),
.Y(n_566)
);

INVxp33_ASAP7_75t_L g579 ( 
.A(n_566),
.Y(n_579)
);

MAJIxp5_ASAP7_75t_L g567 ( 
.A(n_530),
.B(n_508),
.C(n_525),
.Y(n_567)
);

HB1xp67_ASAP7_75t_L g593 ( 
.A(n_569),
.Y(n_593)
);

MAJIxp5_ASAP7_75t_L g570 ( 
.A(n_530),
.B(n_548),
.C(n_542),
.Y(n_570)
);

MAJIxp5_ASAP7_75t_L g586 ( 
.A(n_570),
.B(n_571),
.C(n_578),
.Y(n_586)
);

MAJIxp5_ASAP7_75t_L g571 ( 
.A(n_535),
.B(n_498),
.C(n_507),
.Y(n_571)
);

OAI21xp5_ASAP7_75t_L g574 ( 
.A1(n_534),
.A2(n_556),
.B(n_540),
.Y(n_574)
);

OAI21xp5_ASAP7_75t_L g592 ( 
.A1(n_574),
.A2(n_509),
.B(n_549),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_L g577 ( 
.A(n_533),
.B(n_516),
.Y(n_577)
);

NOR2xp33_ASAP7_75t_L g585 ( 
.A(n_577),
.B(n_536),
.Y(n_585)
);

MAJIxp5_ASAP7_75t_L g578 ( 
.A(n_551),
.B(n_517),
.C(n_512),
.Y(n_578)
);

XNOR2xp5_ASAP7_75t_L g580 ( 
.A(n_570),
.B(n_544),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_L g597 ( 
.A(n_580),
.B(n_587),
.Y(n_597)
);

OAI22xp5_ASAP7_75t_SL g611 ( 
.A1(n_581),
.A2(n_582),
.B1(n_568),
.B2(n_566),
.Y(n_611)
);

AOI22xp5_ASAP7_75t_L g582 ( 
.A1(n_576),
.A2(n_531),
.B1(n_556),
.B2(n_553),
.Y(n_582)
);

OAI22xp5_ASAP7_75t_SL g583 ( 
.A1(n_576),
.A2(n_552),
.B1(n_516),
.B2(n_554),
.Y(n_583)
);

AOI22xp5_ASAP7_75t_L g606 ( 
.A1(n_583),
.A2(n_569),
.B1(n_562),
.B2(n_565),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_585),
.Y(n_607)
);

NOR2xp33_ASAP7_75t_L g587 ( 
.A(n_564),
.B(n_536),
.Y(n_587)
);

MAJIxp5_ASAP7_75t_L g589 ( 
.A(n_563),
.B(n_551),
.C(n_532),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_L g604 ( 
.A(n_589),
.B(n_594),
.Y(n_604)
);

XOR2xp5_ASAP7_75t_L g591 ( 
.A(n_578),
.B(n_555),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_SL g599 ( 
.A(n_591),
.B(n_595),
.Y(n_599)
);

OAI21xp5_ASAP7_75t_L g609 ( 
.A1(n_592),
.A2(n_561),
.B(n_568),
.Y(n_609)
);

NOR2xp33_ASAP7_75t_L g594 ( 
.A(n_564),
.B(n_539),
.Y(n_594)
);

MAJIxp5_ASAP7_75t_L g595 ( 
.A(n_567),
.B(n_571),
.C(n_573),
.Y(n_595)
);

OAI21xp5_ASAP7_75t_L g596 ( 
.A1(n_561),
.A2(n_572),
.B(n_557),
.Y(n_596)
);

OAI21x1_ASAP7_75t_SL g603 ( 
.A1(n_596),
.A2(n_577),
.B(n_560),
.Y(n_603)
);

NOR2xp33_ASAP7_75t_L g598 ( 
.A(n_590),
.B(n_588),
.Y(n_598)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_598),
.Y(n_615)
);

AND2x2_ASAP7_75t_L g600 ( 
.A(n_596),
.B(n_560),
.Y(n_600)
);

AOI22xp5_ASAP7_75t_L g616 ( 
.A1(n_600),
.A2(n_606),
.B1(n_611),
.B2(n_593),
.Y(n_616)
);

NOR2xp33_ASAP7_75t_L g601 ( 
.A(n_580),
.B(n_575),
.Y(n_601)
);

NOR2xp33_ASAP7_75t_L g613 ( 
.A(n_601),
.B(n_608),
.Y(n_613)
);

AOI21xp5_ASAP7_75t_L g602 ( 
.A1(n_582),
.A2(n_562),
.B(n_557),
.Y(n_602)
);

AOI21xp5_ASAP7_75t_L g614 ( 
.A1(n_602),
.A2(n_603),
.B(n_609),
.Y(n_614)
);

MAJIxp5_ASAP7_75t_L g605 ( 
.A(n_586),
.B(n_559),
.C(n_573),
.Y(n_605)
);

NOR2xp67_ASAP7_75t_SL g621 ( 
.A(n_605),
.B(n_610),
.Y(n_621)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_579),
.Y(n_608)
);

MAJIxp5_ASAP7_75t_L g610 ( 
.A(n_586),
.B(n_575),
.C(n_558),
.Y(n_610)
);

OAI22xp5_ASAP7_75t_SL g612 ( 
.A1(n_606),
.A2(n_581),
.B1(n_592),
.B2(n_584),
.Y(n_612)
);

OR2x2_ASAP7_75t_L g625 ( 
.A(n_612),
.B(n_617),
.Y(n_625)
);

XNOR2xp5_ASAP7_75t_L g626 ( 
.A(n_616),
.B(n_620),
.Y(n_626)
);

MAJIxp5_ASAP7_75t_L g617 ( 
.A(n_605),
.B(n_589),
.C(n_595),
.Y(n_617)
);

NOR2xp33_ASAP7_75t_L g618 ( 
.A(n_607),
.B(n_583),
.Y(n_618)
);

CKINVDCx20_ASAP7_75t_R g628 ( 
.A(n_618),
.Y(n_628)
);

OAI21xp5_ASAP7_75t_SL g619 ( 
.A1(n_602),
.A2(n_579),
.B(n_566),
.Y(n_619)
);

OAI21xp5_ASAP7_75t_SL g627 ( 
.A1(n_619),
.A2(n_609),
.B(n_600),
.Y(n_627)
);

NOR2xp33_ASAP7_75t_L g620 ( 
.A(n_604),
.B(n_591),
.Y(n_620)
);

AND2x2_ASAP7_75t_L g622 ( 
.A(n_617),
.B(n_610),
.Y(n_622)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_622),
.Y(n_630)
);

NOR2xp67_ASAP7_75t_L g623 ( 
.A(n_612),
.B(n_611),
.Y(n_623)
);

AOI21xp5_ASAP7_75t_L g629 ( 
.A1(n_623),
.A2(n_627),
.B(n_614),
.Y(n_629)
);

MAJIxp5_ASAP7_75t_L g624 ( 
.A(n_615),
.B(n_599),
.C(n_597),
.Y(n_624)
);

NOR2xp33_ASAP7_75t_SL g631 ( 
.A(n_624),
.B(n_613),
.Y(n_631)
);

MAJIxp5_ASAP7_75t_L g634 ( 
.A(n_629),
.B(n_625),
.C(n_628),
.Y(n_634)
);

NOR2xp33_ASAP7_75t_L g633 ( 
.A(n_631),
.B(n_632),
.Y(n_633)
);

NOR2xp33_ASAP7_75t_SL g632 ( 
.A(n_622),
.B(n_600),
.Y(n_632)
);

MAJIxp5_ASAP7_75t_L g635 ( 
.A(n_634),
.B(n_630),
.C(n_621),
.Y(n_635)
);

MAJIxp5_ASAP7_75t_L g636 ( 
.A(n_635),
.B(n_626),
.C(n_633),
.Y(n_636)
);

NOR2xp33_ASAP7_75t_L g637 ( 
.A(n_636),
.B(n_623),
.Y(n_637)
);

XNOR2xp5_ASAP7_75t_L g638 ( 
.A(n_637),
.B(n_614),
.Y(n_638)
);


endmodule