module fake_jpeg_19809_n_131 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_131);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_131;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_91;
wire n_93;
wire n_54;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

BUFx3_ASAP7_75t_L g43 ( 
.A(n_13),
.Y(n_43)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_21),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_12),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_6),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_30),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_16),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_41),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_42),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_2),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_3),
.Y(n_53)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_24),
.Y(n_54)
);

BUFx4f_ASAP7_75t_SL g55 ( 
.A(n_20),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_7),
.Y(n_56)
);

INVx1_ASAP7_75t_SL g57 ( 
.A(n_11),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_1),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_25),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_18),
.Y(n_60)
);

CKINVDCx14_ASAP7_75t_R g61 ( 
.A(n_15),
.Y(n_61)
);

INVx11_ASAP7_75t_SL g62 ( 
.A(n_40),
.Y(n_62)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_4),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_0),
.Y(n_64)
);

CKINVDCx14_ASAP7_75t_R g65 ( 
.A(n_36),
.Y(n_65)
);

CKINVDCx11_ASAP7_75t_R g66 ( 
.A(n_62),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_66),
.B(n_69),
.Y(n_73)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_46),
.Y(n_67)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_67),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_52),
.Y(n_68)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_68),
.Y(n_79)
);

INVx6_ASAP7_75t_SL g69 ( 
.A(n_52),
.Y(n_69)
);

NAND3xp33_ASAP7_75t_L g70 ( 
.A(n_65),
.B(n_0),
.C(n_1),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_70),
.B(n_71),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_51),
.B(n_2),
.Y(n_71)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_62),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_72),
.B(n_55),
.Y(n_77)
);

INVx13_ASAP7_75t_L g76 ( 
.A(n_66),
.Y(n_76)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_76),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_77),
.Y(n_87)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_68),
.Y(n_78)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_78),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_67),
.B(n_64),
.C(n_44),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_80),
.B(n_64),
.C(n_65),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_72),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_81),
.B(n_55),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_69),
.B(n_56),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_82),
.B(n_50),
.Y(n_91)
);

O2A1O1Ixp33_ASAP7_75t_L g83 ( 
.A1(n_66),
.A2(n_45),
.B(n_47),
.C(n_48),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_83),
.A2(n_61),
.B1(n_58),
.B2(n_49),
.Y(n_89)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_84),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_78),
.A2(n_79),
.B1(n_63),
.B2(n_57),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_85),
.A2(n_43),
.B1(n_53),
.B2(n_7),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_88),
.B(n_90),
.Y(n_104)
);

O2A1O1Ixp33_ASAP7_75t_L g108 ( 
.A1(n_89),
.A2(n_5),
.B(n_6),
.C(n_8),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_74),
.B(n_61),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_91),
.B(n_73),
.Y(n_97)
);

INVx1_ASAP7_75t_SL g92 ( 
.A(n_76),
.Y(n_92)
);

OR2x2_ASAP7_75t_L g110 ( 
.A(n_92),
.B(n_5),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_75),
.B(n_60),
.Y(n_93)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_93),
.Y(n_103)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_83),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_95),
.B(n_96),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_80),
.B(n_59),
.C(n_54),
.Y(n_96)
);

NOR3xp33_ASAP7_75t_SL g114 ( 
.A(n_97),
.B(n_19),
.C(n_22),
.Y(n_114)
);

CKINVDCx14_ASAP7_75t_R g99 ( 
.A(n_85),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_99),
.B(n_101),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_86),
.B(n_3),
.Y(n_101)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_94),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_102),
.A2(n_107),
.B1(n_100),
.B2(n_99),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_92),
.B(n_4),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_105),
.B(n_26),
.C(n_28),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_106),
.A2(n_109),
.B1(n_110),
.B2(n_8),
.Y(n_111)
);

HB1xp67_ASAP7_75t_L g107 ( 
.A(n_87),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_108),
.A2(n_10),
.B1(n_14),
.B2(n_17),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_87),
.A2(n_27),
.B1(n_37),
.B2(n_9),
.Y(n_109)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_111),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_L g119 ( 
.A1(n_112),
.A2(n_114),
.B(n_115),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_L g115 ( 
.A(n_104),
.B(n_23),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_116),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_118),
.B(n_98),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_L g123 ( 
.A1(n_121),
.A2(n_122),
.B(n_110),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_120),
.A2(n_113),
.B1(n_116),
.B2(n_107),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_123),
.B(n_122),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_SL g125 ( 
.A1(n_124),
.A2(n_103),
.B(n_114),
.Y(n_125)
);

AO21x1_ASAP7_75t_L g126 ( 
.A1(n_125),
.A2(n_119),
.B(n_117),
.Y(n_126)
);

OR2x2_ASAP7_75t_L g127 ( 
.A(n_126),
.B(n_29),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_SL g128 ( 
.A1(n_127),
.A2(n_39),
.B(n_32),
.Y(n_128)
);

OAI21x1_ASAP7_75t_L g129 ( 
.A1(n_128),
.A2(n_31),
.B(n_33),
.Y(n_129)
);

XOR2xp5_ASAP7_75t_L g130 ( 
.A(n_129),
.B(n_34),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_L g131 ( 
.A(n_130),
.B(n_35),
.Y(n_131)
);


endmodule