module fake_jpeg_7244_n_131 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_131);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_131;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_8),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_3),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_9),
.Y(n_13)
);

INVx13_ASAP7_75t_L g14 ( 
.A(n_3),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_9),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_10),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_0),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_7),
.Y(n_19)
);

CKINVDCx12_ASAP7_75t_R g20 ( 
.A(n_2),
.Y(n_20)
);

INVx11_ASAP7_75t_SL g21 ( 
.A(n_0),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_5),
.Y(n_22)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_23),
.Y(n_32)
);

INVx4_ASAP7_75t_SL g24 ( 
.A(n_14),
.Y(n_24)
);

AOI22xp33_ASAP7_75t_SL g41 ( 
.A1(n_24),
.A2(n_31),
.B1(n_12),
.B2(n_13),
.Y(n_41)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_25),
.B(n_27),
.Y(n_35)
);

INVx5_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_21),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_22),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_SL g33 ( 
.A(n_28),
.B(n_30),
.Y(n_33)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_21),
.Y(n_29)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_22),
.Y(n_30)
);

INVx5_ASAP7_75t_L g31 ( 
.A(n_20),
.Y(n_31)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_27),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_34),
.B(n_37),
.Y(n_49)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_27),
.Y(n_37)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_23),
.Y(n_38)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_38),
.Y(n_42)
);

AND2x2_ASAP7_75t_L g39 ( 
.A(n_25),
.B(n_0),
.Y(n_39)
);

AOI21xp5_ASAP7_75t_L g56 ( 
.A1(n_39),
.A2(n_12),
.B(n_17),
.Y(n_56)
);

CKINVDCx16_ASAP7_75t_R g52 ( 
.A(n_41),
.Y(n_52)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_35),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_43),
.B(n_45),
.Y(n_74)
);

OAI22xp33_ASAP7_75t_SL g44 ( 
.A1(n_41),
.A2(n_24),
.B1(n_26),
.B2(n_29),
.Y(n_44)
);

OAI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_44),
.A2(n_24),
.B1(n_29),
.B2(n_40),
.Y(n_67)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

AND2x6_ASAP7_75t_L g46 ( 
.A(n_39),
.B(n_5),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_46),
.A2(n_53),
.B1(n_55),
.B2(n_19),
.Y(n_79)
);

CKINVDCx12_ASAP7_75t_R g47 ( 
.A(n_33),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_47),
.B(n_48),
.Y(n_62)
);

INVx13_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_50),
.B(n_57),
.Y(n_76)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_33),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_51),
.B(n_30),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_34),
.A2(n_23),
.B1(n_25),
.B2(n_26),
.Y(n_53)
);

AND2x2_ASAP7_75t_L g54 ( 
.A(n_39),
.B(n_13),
.Y(n_54)
);

AOI21xp5_ASAP7_75t_L g70 ( 
.A1(n_54),
.A2(n_61),
.B(n_15),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_37),
.A2(n_29),
.B1(n_23),
.B2(n_13),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_SL g63 ( 
.A(n_56),
.B(n_60),
.Y(n_63)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_36),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_36),
.B(n_30),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_58),
.B(n_59),
.Y(n_77)
);

INVx13_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_40),
.Y(n_60)
);

MAJIxp5_ASAP7_75t_L g61 ( 
.A(n_39),
.B(n_24),
.C(n_31),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_51),
.B(n_28),
.Y(n_64)
);

OR2x2_ASAP7_75t_L g81 ( 
.A(n_64),
.B(n_47),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_65),
.B(n_73),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_54),
.B(n_32),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_66),
.B(n_69),
.Y(n_86)
);

O2A1O1Ixp33_ASAP7_75t_L g90 ( 
.A1(n_67),
.A2(n_60),
.B(n_59),
.C(n_57),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_52),
.A2(n_31),
.B1(n_12),
.B2(n_17),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_68),
.A2(n_55),
.B1(n_48),
.B2(n_32),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_54),
.B(n_28),
.Y(n_69)
);

OAI21xp5_ASAP7_75t_SL g85 ( 
.A1(n_70),
.A2(n_72),
.B(n_53),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_56),
.B(n_17),
.Y(n_71)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_71),
.Y(n_80)
);

AOI21xp5_ASAP7_75t_L g72 ( 
.A1(n_52),
.A2(n_32),
.B(n_40),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_49),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_43),
.B(n_15),
.Y(n_75)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_75),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_45),
.B(n_15),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_78),
.B(n_61),
.C(n_49),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_79),
.B(n_46),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_81),
.B(n_82),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_SL g101 ( 
.A1(n_85),
.A2(n_87),
.B(n_88),
.Y(n_101)
);

AOI21xp5_ASAP7_75t_SL g87 ( 
.A1(n_71),
.A2(n_69),
.B(n_66),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_89),
.A2(n_94),
.B1(n_80),
.B2(n_84),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_90),
.A2(n_74),
.B1(n_79),
.B2(n_63),
.Y(n_97)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_76),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_91),
.B(n_77),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_L g92 ( 
.A1(n_63),
.A2(n_18),
.B(n_19),
.Y(n_92)
);

A2O1A1O1Ixp25_ASAP7_75t_L g98 ( 
.A1(n_92),
.A2(n_74),
.B(n_62),
.C(n_78),
.D(n_75),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_73),
.B(n_42),
.C(n_50),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_93),
.B(n_94),
.C(n_16),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_70),
.B(n_42),
.C(n_19),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_96),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_97),
.A2(n_99),
.B1(n_80),
.B2(n_84),
.Y(n_107)
);

XNOR2xp5_ASAP7_75t_L g112 ( 
.A(n_98),
.B(n_100),
.Y(n_112)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_83),
.Y(n_99)
);

XOR2xp5_ASAP7_75t_L g102 ( 
.A(n_82),
.B(n_72),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_102),
.B(n_104),
.C(n_88),
.Y(n_113)
);

A2O1A1O1Ixp25_ASAP7_75t_L g103 ( 
.A1(n_92),
.A2(n_64),
.B(n_65),
.C(n_20),
.D(n_3),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_L g109 ( 
.A1(n_103),
.A2(n_105),
.B(n_86),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_L g104 ( 
.A(n_87),
.B(n_7),
.Y(n_104)
);

XOR2xp5_ASAP7_75t_L g106 ( 
.A(n_102),
.B(n_85),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_106),
.B(n_113),
.C(n_11),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_L g117 ( 
.A(n_107),
.B(n_108),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_101),
.A2(n_90),
.B1(n_98),
.B2(n_97),
.Y(n_108)
);

AOI321xp33_ASAP7_75t_L g116 ( 
.A1(n_109),
.A2(n_16),
.A3(n_11),
.B1(n_18),
.B2(n_4),
.C(n_5),
.Y(n_116)
);

AOI21xp5_ASAP7_75t_L g110 ( 
.A1(n_101),
.A2(n_86),
.B(n_93),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_110),
.B(n_7),
.Y(n_115)
);

AOI322xp5_ASAP7_75t_L g114 ( 
.A1(n_112),
.A2(n_95),
.A3(n_104),
.B1(n_105),
.B2(n_103),
.C1(n_81),
.C2(n_16),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_114),
.B(n_116),
.Y(n_120)
);

BUFx24_ASAP7_75t_SL g118 ( 
.A(n_111),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_118),
.B(n_119),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_117),
.A2(n_108),
.B1(n_113),
.B2(n_106),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_SL g124 ( 
.A1(n_121),
.A2(n_123),
.B(n_2),
.Y(n_124)
);

AOI21xp5_ASAP7_75t_L g123 ( 
.A1(n_115),
.A2(n_18),
.B(n_6),
.Y(n_123)
);

XNOR2xp5_ASAP7_75t_L g126 ( 
.A(n_124),
.B(n_125),
.Y(n_126)
);

AOI21xp5_ASAP7_75t_SL g125 ( 
.A1(n_120),
.A2(n_6),
.B(n_8),
.Y(n_125)
);

AOI322xp5_ASAP7_75t_L g127 ( 
.A1(n_124),
.A2(n_0),
.A3(n_1),
.B1(n_8),
.B2(n_10),
.C1(n_122),
.C2(n_120),
.Y(n_127)
);

AOI21xp5_ASAP7_75t_L g129 ( 
.A1(n_127),
.A2(n_10),
.B(n_1),
.Y(n_129)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_126),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_128),
.B(n_129),
.C(n_126),
.Y(n_130)
);

BUFx24_ASAP7_75t_SL g131 ( 
.A(n_130),
.Y(n_131)
);


endmodule