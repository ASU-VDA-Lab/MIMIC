module fake_netlist_5_1237_n_1911 (n_137, n_168, n_164, n_91, n_82, n_122, n_142, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_165, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_60, n_155, n_152, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_125, n_35, n_167, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_157, n_29, n_79, n_131, n_151, n_47, n_173, n_25, n_53, n_160, n_8, n_158, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_159, n_163, n_95, n_119, n_169, n_59, n_26, n_133, n_55, n_99, n_2, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_162, n_27, n_170, n_64, n_77, n_102, n_106, n_161, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_174, n_134, n_32, n_41, n_104, n_172, n_103, n_56, n_51, n_63, n_97, n_141, n_166, n_11, n_171, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_1911);

input n_137;
input n_168;
input n_164;
input n_91;
input n_82;
input n_122;
input n_142;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_165;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_60;
input n_155;
input n_152;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_125;
input n_35;
input n_167;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_157;
input n_29;
input n_79;
input n_131;
input n_151;
input n_47;
input n_173;
input n_25;
input n_53;
input n_160;
input n_8;
input n_158;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_159;
input n_163;
input n_95;
input n_119;
input n_169;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_162;
input n_27;
input n_170;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_174;
input n_134;
input n_32;
input n_41;
input n_104;
input n_172;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_166;
input n_11;
input n_171;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_1911;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1729;
wire n_1166;
wire n_1751;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1859;
wire n_1677;
wire n_1150;
wire n_226;
wire n_1780;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1738;
wire n_1021;
wire n_551;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1695;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_1789;
wire n_1666;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_1545;
wire n_864;
wire n_859;
wire n_951;
wire n_1264;
wire n_447;
wire n_247;
wire n_1494;
wire n_292;
wire n_625;
wire n_854;
wire n_1462;
wire n_1799;
wire n_1580;
wire n_674;
wire n_417;
wire n_1806;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_1869;
wire n_1607;
wire n_1563;
wire n_606;
wire n_275;
wire n_877;
wire n_1696;
wire n_755;
wire n_1118;
wire n_1686;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1860;
wire n_1359;
wire n_530;
wire n_1107;
wire n_1728;
wire n_556;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_1896;
wire n_929;
wire n_1124;
wire n_1818;
wire n_902;
wire n_1576;
wire n_191;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1705;
wire n_1257;
wire n_1182;
wire n_579;
wire n_1698;
wire n_1261;
wire n_938;
wire n_1098;
wire n_320;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_519;
wire n_406;
wire n_1016;
wire n_1243;
wire n_546;
wire n_1280;
wire n_1845;
wire n_281;
wire n_240;
wire n_291;
wire n_231;
wire n_257;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_317;
wire n_1236;
wire n_1633;
wire n_569;
wire n_1778;
wire n_227;
wire n_920;
wire n_1289;
wire n_1517;
wire n_335;
wire n_1669;
wire n_370;
wire n_976;
wire n_343;
wire n_1449;
wire n_308;
wire n_1566;
wire n_297;
wire n_1078;
wire n_1670;
wire n_775;
wire n_219;
wire n_600;
wire n_1484;
wire n_1374;
wire n_1328;
wire n_223;
wire n_264;
wire n_1877;
wire n_1831;
wire n_1598;
wire n_1723;
wire n_955;
wire n_1850;
wire n_339;
wire n_1146;
wire n_882;
wire n_183;
wire n_243;
wire n_1097;
wire n_1036;
wire n_1749;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_215;
wire n_350;
wire n_196;
wire n_798;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_290;
wire n_580;
wire n_1040;
wire n_1872;
wire n_1852;
wire n_578;
wire n_926;
wire n_344;
wire n_1218;
wire n_422;
wire n_475;
wire n_777;
wire n_1070;
wire n_1547;
wire n_1030;
wire n_1755;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1801;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_663;
wire n_845;
wire n_1862;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_1796;
wire n_680;
wire n_1473;
wire n_1587;
wire n_395;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_214;
wire n_1748;
wire n_1672;
wire n_675;
wire n_888;
wire n_1880;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1384;
wire n_1556;
wire n_184;
wire n_446;
wire n_1863;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_1706;
wire n_468;
wire n_213;
wire n_342;
wire n_464;
wire n_363;
wire n_1582;
wire n_197;
wire n_1069;
wire n_1784;
wire n_1075;
wire n_1836;
wire n_1450;
wire n_1322;
wire n_1471;
wire n_1750;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_1700;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1599;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_907;
wire n_1447;
wire n_1377;
wire n_190;
wire n_989;
wire n_1039;
wire n_228;
wire n_283;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_310;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_1667;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1248;
wire n_230;
wire n_1331;
wire n_953;
wire n_1014;
wire n_279;
wire n_1241;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_1819;
wire n_476;
wire n_1527;
wire n_534;
wire n_1882;
wire n_884;
wire n_345;
wire n_944;
wire n_1754;
wire n_1623;
wire n_1854;
wire n_1565;
wire n_1809;
wire n_1856;
wire n_182;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_857;
wire n_832;
wire n_207;
wire n_561;
wire n_1319;
wire n_1825;
wire n_1883;
wire n_1906;
wire n_1712;
wire n_1387;
wire n_1532;
wire n_1027;
wire n_971;
wire n_1156;
wire n_326;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1775;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_1709;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1538;
wire n_1838;
wire n_1199;
wire n_1847;
wire n_1779;
wire n_352;
wire n_1884;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_1841;
wire n_1660;
wire n_887;
wire n_1905;
wire n_300;
wire n_809;
wire n_870;
wire n_931;
wire n_599;
wire n_1711;
wire n_1662;
wire n_1891;
wire n_1481;
wire n_434;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1629;
wire n_1293;
wire n_965;
wire n_1876;
wire n_1743;
wire n_935;
wire n_1175;
wire n_817;
wire n_360;
wire n_1479;
wire n_1810;
wire n_1888;
wire n_759;
wire n_1892;
wire n_806;
wire n_1766;
wire n_1477;
wire n_324;
wire n_1635;
wire n_1571;
wire n_187;
wire n_1189;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_784;
wire n_1733;
wire n_1244;
wire n_431;
wire n_1194;
wire n_1815;
wire n_615;
wire n_851;
wire n_1759;
wire n_843;
wire n_1788;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_1679;
wire n_776;
wire n_1798;
wire n_1790;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1746;
wire n_1647;
wire n_1829;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_1674;
wire n_1833;
wire n_1830;
wire n_1710;
wire n_284;
wire n_1128;
wire n_1734;
wire n_744;
wire n_629;
wire n_590;
wire n_1308;
wire n_1767;
wire n_254;
wire n_1680;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_526;
wire n_293;
wire n_372;
wire n_677;
wire n_244;
wire n_1333;
wire n_1121;
wire n_314;
wire n_368;
wire n_433;
wire n_604;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_498;
wire n_1468;
wire n_1559;
wire n_1765;
wire n_1866;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_624;
wire n_252;
wire n_1380;
wire n_1744;
wire n_1617;
wire n_295;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_1837;
wire n_1839;
wire n_610;
wire n_1760;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_1832;
wire n_259;
wire n_448;
wire n_1851;
wire n_758;
wire n_999;
wire n_1656;
wire n_1158;
wire n_1509;
wire n_1874;
wire n_563;
wire n_1145;
wire n_878;
wire n_524;
wire n_394;
wire n_204;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_1871;
wire n_331;
wire n_906;
wire n_1163;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_1781;
wire n_658;
wire n_1740;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_1773;
wire n_592;
wire n_1169;
wire n_1596;
wire n_1692;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_1095;
wire n_1828;
wire n_1614;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_1431;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1640;
wire n_1732;
wire n_1009;
wire n_1148;
wire n_750;
wire n_742;
wire n_995;
wire n_454;
wire n_1609;
wire n_374;
wire n_185;
wire n_396;
wire n_1887;
wire n_1383;
wire n_1073;
wire n_255;
wire n_662;
wire n_459;
wire n_218;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1721;
wire n_1758;
wire n_1574;
wire n_473;
wire n_1309;
wire n_1878;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_1800;
wire n_1548;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_208;
wire n_743;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_1240;
wire n_1820;
wire n_829;
wire n_1612;
wire n_1416;
wire n_1724;
wire n_361;
wire n_1237;
wire n_700;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1785;
wire n_1568;
wire n_1006;
wire n_329;
wire n_274;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_1870;
wire n_309;
wire n_512;
wire n_1591;
wire n_322;
wire n_1682;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1349;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_1909;
wire n_224;
wire n_1562;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_239;
wire n_630;
wire n_1902;
wire n_504;
wire n_1823;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_1875;
wire n_1304;
wire n_1324;
wire n_987;
wire n_1846;
wire n_261;
wire n_1885;
wire n_1455;
wire n_767;
wire n_993;
wire n_1903;
wire n_1407;
wire n_1551;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_1805;
wire n_1816;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_1849;
wire n_729;
wire n_1131;
wire n_1084;
wire n_970;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_340;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_1645;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_1684;
wire n_233;
wire n_1717;
wire n_572;
wire n_366;
wire n_815;
wire n_1795;
wire n_1821;
wire n_327;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_1708;
wire n_426;
wire n_1438;
wire n_1082;
wire n_1840;
wire n_589;
wire n_716;
wire n_1630;
wire n_562;
wire n_1436;
wire n_1691;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_1776;
wire n_531;
wire n_1757;
wire n_890;
wire n_1897;
wire n_764;
wire n_1056;
wire n_1424;
wire n_960;
wire n_1893;
wire n_222;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_634;
wire n_199;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_1519;
wire n_256;
wire n_950;
wire n_1553;
wire n_1811;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1808;
wire n_1060;
wire n_1141;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_968;
wire n_912;
wire n_315;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_1699;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_1050;
wire n_841;
wire n_802;
wire n_1608;
wire n_983;
wire n_1844;
wire n_280;
wire n_1305;
wire n_873;
wire n_1826;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_1644;
wire n_690;
wire n_583;
wire n_302;
wire n_1343;
wire n_1203;
wire n_1631;
wire n_821;
wire n_1763;
wire n_1768;
wire n_321;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1719;
wire n_1288;
wire n_212;
wire n_385;
wire n_507;
wire n_1560;
wire n_1605;
wire n_330;
wire n_1228;
wire n_972;
wire n_692;
wire n_820;
wire n_1200;
wire n_1301;
wire n_1363;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_1688;
wire n_945;
wire n_492;
wire n_1504;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_286;
wire n_1643;
wire n_883;
wire n_470;
wire n_325;
wire n_449;
wire n_1594;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_856;
wire n_1793;
wire n_918;
wire n_942;
wire n_1804;
wire n_189;
wire n_1147;
wire n_1557;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_195;
wire n_356;
wire n_894;
wire n_1636;
wire n_1730;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1865;
wire n_1470;
wire n_1096;
wire n_234;
wire n_1575;
wire n_1697;
wire n_1735;
wire n_833;
wire n_1646;
wire n_225;
wire n_1307;
wire n_1881;
wire n_988;
wire n_814;
wire n_192;
wire n_1549;
wire n_1201;
wire n_1114;
wire n_655;
wire n_1616;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_1807;
wire n_387;
wire n_1149;
wire n_398;
wire n_1671;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_211;
wire n_1824;
wire n_1219;
wire n_1204;
wire n_178;
wire n_1814;
wire n_1035;
wire n_287;
wire n_555;
wire n_783;
wire n_1848;
wire n_1188;
wire n_1722;
wire n_661;
wire n_1802;
wire n_849;
wire n_584;
wire n_681;
wire n_336;
wire n_1638;
wire n_1786;
wire n_430;
wire n_510;
wire n_216;
wire n_311;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_1655;
wire n_445;
wire n_749;
wire n_1895;
wire n_1134;
wire n_1358;
wire n_717;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_249;
wire n_304;
wire n_1338;
wire n_577;
wire n_1522;
wire n_1687;
wire n_1637;
wire n_1419;
wire n_338;
wire n_1653;
wire n_693;
wire n_1506;
wire n_836;
wire n_990;
wire n_1886;
wire n_1389;
wire n_1894;
wire n_975;
wire n_1908;
wire n_1256;
wire n_1702;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_306;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_1843;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1164;
wire n_1659;
wire n_1834;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_1572;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1736;
wire n_1685;
wire n_601;
wire n_917;
wire n_1714;
wire n_966;
wire n_253;
wire n_1116;
wire n_1661;
wire n_1212;
wire n_1541;
wire n_206;
wire n_217;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_1731;
wire n_818;
wire n_861;
wire n_1713;
wire n_1183;
wire n_1658;
wire n_899;
wire n_1253;
wire n_210;
wire n_1737;
wire n_1904;
wire n_774;
wire n_1628;
wire n_1335;
wire n_1514;
wire n_1777;
wire n_1059;
wire n_1345;
wire n_176;
wire n_1133;
wire n_1771;
wire n_1899;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_707;
wire n_1168;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_1584;
wire n_665;
wire n_1726;
wire n_1835;
wire n_1440;
wire n_177;
wire n_421;
wire n_1853;
wire n_1356;
wire n_1787;
wire n_910;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1774;
wire n_1725;
wire n_205;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_179;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_1812;
wire n_735;
wire n_232;
wire n_1109;
wire n_895;
wire n_1310;
wire n_1803;
wire n_202;
wire n_427;
wire n_1399;
wire n_1543;
wire n_791;
wire n_732;
wire n_1533;
wire n_193;
wire n_808;
wire n_797;
wire n_1025;
wire n_500;
wire n_1067;
wire n_1720;
wire n_435;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1742;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_594;
wire n_200;
wire n_1291;
wire n_1297;
wire n_1753;
wire n_1782;
wire n_1155;
wire n_1418;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_985;
wire n_1855;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1703;
wire n_1352;
wire n_626;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_305;
wire n_676;
wire n_294;
wire n_318;
wire n_653;
wire n_642;
wire n_1602;
wire n_194;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_268;
wire n_664;
wire n_503;
wire n_235;
wire n_1372;
wire n_605;
wire n_1273;
wire n_1822;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_1783;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_1907;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_1898;
wire n_581;
wire n_382;
wire n_554;
wire n_1625;
wire n_898;
wire n_1762;
wire n_1013;
wire n_1452;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_1791;
wire n_198;
wire n_1890;
wire n_1747;
wire n_714;
wire n_1683;
wire n_1817;
wire n_909;
wire n_1530;
wire n_1497;
wire n_997;
wire n_932;
wire n_612;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_508;
wire n_506;
wire n_1320;
wire n_1663;
wire n_737;
wire n_1718;
wire n_986;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1715;
wire n_1281;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_1889;
wire n_209;
wire n_1792;
wire n_1564;
wire n_1868;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1376;
wire n_941;
wire n_981;
wire n_1569;
wire n_867;
wire n_186;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_518;
wire n_505;
wire n_1772;
wire n_282;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1861;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1901;
wire n_1900;
wire n_1620;
wire n_381;
wire n_220;
wire n_390;
wire n_1330;
wire n_1867;
wire n_481;
wire n_1675;
wire n_1727;
wire n_1554;
wire n_1745;
wire n_769;
wire n_1046;
wire n_271;
wire n_934;
wire n_1618;
wire n_826;
wire n_1813;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_428;
wire n_379;
wire n_1341;
wire n_570;
wire n_1641;
wire n_1361;
wire n_1707;
wire n_853;
wire n_377;
wire n_751;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_704;
wire n_787;
wire n_1770;
wire n_961;
wire n_1756;
wire n_771;
wire n_276;
wire n_1716;
wire n_1225;
wire n_1520;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_181;
wire n_1873;
wire n_1411;
wire n_221;
wire n_622;
wire n_1577;
wire n_1087;
wire n_386;
wire n_994;
wire n_1701;
wire n_848;
wire n_1550;
wire n_1498;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1857;
wire n_1344;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_1797;
wire n_432;
wire n_1769;
wire n_839;
wire n_1210;
wire n_1364;
wire n_328;
wire n_1250;
wire n_369;
wire n_1842;
wire n_871;
wire n_685;
wire n_598;
wire n_608;
wire n_928;
wire n_1367;
wire n_1460;
wire n_772;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_402;
wire n_413;
wire n_1086;
wire n_796;
wire n_1858;
wire n_1619;
wire n_236;
wire n_1502;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_903;
wire n_1525;
wire n_1752;
wire n_740;
wire n_203;
wire n_384;
wire n_1404;
wire n_1794;
wire n_1315;
wire n_277;
wire n_1061;
wire n_1910;
wire n_333;
wire n_1298;
wire n_1652;
wire n_462;
wire n_1193;
wire n_1676;
wire n_1255;
wire n_258;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_188;
wire n_844;
wire n_201;
wire n_471;
wire n_852;
wire n_1487;
wire n_1864;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_1673;
wire n_465;
wire n_1321;
wire n_362;
wire n_273;
wire n_585;
wire n_1739;
wire n_270;
wire n_616;
wire n_745;
wire n_1654;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_1761;
wire n_641;
wire n_730;
wire n_1325;
wire n_1595;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_180;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_229;
wire n_437;
wire n_1642;
wire n_403;
wire n_453;
wire n_1130;
wire n_720;
wire n_1526;
wire n_863;
wire n_805;
wire n_1604;
wire n_1275;
wire n_1764;
wire n_712;
wire n_246;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_269;
wire n_285;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1741;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_1621;
wire n_251;
wire n_566;
wire n_565;
wire n_1448;
wire n_1507;
wire n_1398;
wire n_1879;
wire n_597;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_651;
wire n_1340;
wire n_334;
wire n_811;
wire n_1558;
wire n_807;
wire n_835;
wire n_175;
wire n_666;
wire n_262;
wire n_1433;
wire n_1704;
wire n_1254;
wire n_1026;
wire n_1234;
wire n_319;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_242;
wire n_1681;
wire n_1018;
wire n_1693;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_1180;
wire n_1827;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;
wire n_278;

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_122),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_127),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_24),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_33),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_62),
.Y(n_179)
);

INVx1_ASAP7_75t_SL g180 ( 
.A(n_100),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_81),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_11),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_160),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_0),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_80),
.Y(n_185)
);

INVxp67_ASAP7_75t_L g186 ( 
.A(n_52),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_95),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_128),
.Y(n_188)
);

BUFx6f_ASAP7_75t_L g189 ( 
.A(n_102),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_153),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_32),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_35),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_159),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_38),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_74),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_104),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_162),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_163),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_133),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_129),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_107),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_111),
.Y(n_202)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_138),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_18),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_118),
.Y(n_205)
);

INVx1_ASAP7_75t_SL g206 ( 
.A(n_33),
.Y(n_206)
);

INVx2_ASAP7_75t_SL g207 ( 
.A(n_60),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_156),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_0),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_48),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_79),
.Y(n_211)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_55),
.Y(n_212)
);

INVxp33_ASAP7_75t_R g213 ( 
.A(n_51),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_50),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_77),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_125),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_126),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_10),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_113),
.Y(n_219)
);

BUFx2_ASAP7_75t_L g220 ( 
.A(n_73),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_88),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_78),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_52),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_112),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_168),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_99),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_124),
.Y(n_227)
);

BUFx10_ASAP7_75t_L g228 ( 
.A(n_101),
.Y(n_228)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_1),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_114),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_27),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_50),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_21),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_30),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_11),
.Y(n_235)
);

CKINVDCx16_ASAP7_75t_R g236 ( 
.A(n_167),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_161),
.Y(n_237)
);

INVx2_ASAP7_75t_SL g238 ( 
.A(n_132),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_26),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_83),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_39),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_13),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_32),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_48),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_62),
.Y(n_245)
);

INVx1_ASAP7_75t_SL g246 ( 
.A(n_47),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_123),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_71),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_12),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_20),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_143),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_94),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_157),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_154),
.Y(n_254)
);

INVx1_ASAP7_75t_SL g255 ( 
.A(n_27),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_28),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_8),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_3),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_58),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_65),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_93),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_150),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_17),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_119),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_61),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_31),
.Y(n_266)
);

BUFx2_ASAP7_75t_L g267 ( 
.A(n_56),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_142),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_134),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_19),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_103),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_19),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_170),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_31),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_35),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_173),
.Y(n_276)
);

BUFx10_ASAP7_75t_L g277 ( 
.A(n_85),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_68),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_110),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_169),
.Y(n_280)
);

INVx1_ASAP7_75t_SL g281 ( 
.A(n_64),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_10),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_57),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_69),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_130),
.Y(n_285)
);

BUFx6f_ASAP7_75t_L g286 ( 
.A(n_121),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_166),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_92),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_23),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_135),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_39),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_57),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_44),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_165),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_18),
.Y(n_295)
);

BUFx5_ASAP7_75t_L g296 ( 
.A(n_152),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_70),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_15),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_28),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_63),
.Y(n_300)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_155),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_59),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_146),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_43),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_151),
.Y(n_305)
);

INVx2_ASAP7_75t_L g306 ( 
.A(n_116),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_59),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_90),
.Y(n_308)
);

INVx1_ASAP7_75t_SL g309 ( 
.A(n_158),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_24),
.Y(n_310)
);

BUFx6f_ASAP7_75t_L g311 ( 
.A(n_97),
.Y(n_311)
);

INVxp67_ASAP7_75t_SL g312 ( 
.A(n_75),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_13),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_29),
.Y(n_314)
);

BUFx6f_ASAP7_75t_L g315 ( 
.A(n_61),
.Y(n_315)
);

INVx1_ASAP7_75t_SL g316 ( 
.A(n_30),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_55),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_41),
.Y(n_318)
);

BUFx10_ASAP7_75t_L g319 ( 
.A(n_46),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_60),
.Y(n_320)
);

CKINVDCx16_ASAP7_75t_R g321 ( 
.A(n_82),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_136),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_117),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_96),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_1),
.Y(n_325)
);

BUFx3_ASAP7_75t_L g326 ( 
.A(n_58),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_5),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_45),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_145),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_91),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_42),
.Y(n_331)
);

BUFx8_ASAP7_75t_SL g332 ( 
.A(n_140),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_21),
.Y(n_333)
);

INVx2_ASAP7_75t_L g334 ( 
.A(n_8),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_17),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_22),
.Y(n_336)
);

CKINVDCx16_ASAP7_75t_R g337 ( 
.A(n_22),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_87),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g339 ( 
.A(n_25),
.Y(n_339)
);

CKINVDCx16_ASAP7_75t_R g340 ( 
.A(n_20),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_105),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_5),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_42),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_148),
.Y(n_344)
);

BUFx3_ASAP7_75t_L g345 ( 
.A(n_46),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_36),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_98),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_29),
.Y(n_348)
);

INVxp33_ASAP7_75t_SL g349 ( 
.A(n_178),
.Y(n_349)
);

INVxp67_ASAP7_75t_L g350 ( 
.A(n_267),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_315),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_315),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_337),
.Y(n_353)
);

CKINVDCx16_ASAP7_75t_R g354 ( 
.A(n_340),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_326),
.Y(n_355)
);

CKINVDCx20_ASAP7_75t_R g356 ( 
.A(n_201),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_326),
.Y(n_357)
);

INVxp67_ASAP7_75t_SL g358 ( 
.A(n_220),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_345),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_345),
.Y(n_360)
);

INVxp33_ASAP7_75t_L g361 ( 
.A(n_177),
.Y(n_361)
);

INVxp33_ASAP7_75t_SL g362 ( 
.A(n_178),
.Y(n_362)
);

INVxp67_ASAP7_75t_SL g363 ( 
.A(n_315),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_315),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_315),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_212),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_212),
.Y(n_367)
);

INVxp67_ASAP7_75t_SL g368 ( 
.A(n_183),
.Y(n_368)
);

BUFx6f_ASAP7_75t_L g369 ( 
.A(n_189),
.Y(n_369)
);

CKINVDCx20_ASAP7_75t_R g370 ( 
.A(n_208),
.Y(n_370)
);

INVxp67_ASAP7_75t_L g371 ( 
.A(n_319),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_229),
.Y(n_372)
);

CKINVDCx16_ASAP7_75t_R g373 ( 
.A(n_236),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_229),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_334),
.Y(n_375)
);

CKINVDCx20_ASAP7_75t_R g376 ( 
.A(n_247),
.Y(n_376)
);

CKINVDCx20_ASAP7_75t_R g377 ( 
.A(n_248),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_334),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_239),
.Y(n_379)
);

CKINVDCx20_ASAP7_75t_R g380 ( 
.A(n_285),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_214),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_243),
.Y(n_382)
);

HB1xp67_ASAP7_75t_L g383 ( 
.A(n_179),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_218),
.Y(n_384)
);

HB1xp67_ASAP7_75t_L g385 ( 
.A(n_179),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_245),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_249),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_256),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_257),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_223),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_259),
.Y(n_391)
);

CKINVDCx20_ASAP7_75t_R g392 ( 
.A(n_324),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_270),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_274),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_231),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_282),
.Y(n_396)
);

CKINVDCx20_ASAP7_75t_R g397 ( 
.A(n_329),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_233),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_292),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_235),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_293),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_304),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_314),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_241),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_325),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_327),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_343),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_185),
.Y(n_408)
);

CKINVDCx20_ASAP7_75t_R g409 ( 
.A(n_332),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_187),
.Y(n_410)
);

HB1xp67_ASAP7_75t_L g411 ( 
.A(n_182),
.Y(n_411)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_296),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_242),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_195),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_197),
.Y(n_415)
);

CKINVDCx20_ASAP7_75t_R g416 ( 
.A(n_321),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_211),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_244),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_215),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_221),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_224),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_207),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_207),
.Y(n_423)
);

CKINVDCx14_ASAP7_75t_R g424 ( 
.A(n_319),
.Y(n_424)
);

CKINVDCx20_ASAP7_75t_R g425 ( 
.A(n_216),
.Y(n_425)
);

INVxp67_ASAP7_75t_L g426 ( 
.A(n_319),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_250),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_203),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_203),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_301),
.Y(n_430)
);

INVxp67_ASAP7_75t_L g431 ( 
.A(n_182),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_258),
.Y(n_432)
);

CKINVDCx20_ASAP7_75t_R g433 ( 
.A(n_217),
.Y(n_433)
);

CKINVDCx20_ASAP7_75t_R g434 ( 
.A(n_219),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_263),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_301),
.Y(n_436)
);

INVx1_ASAP7_75t_SL g437 ( 
.A(n_232),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_265),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_266),
.Y(n_439)
);

INVxp33_ASAP7_75t_SL g440 ( 
.A(n_184),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_351),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_351),
.Y(n_442)
);

AND2x2_ASAP7_75t_L g443 ( 
.A(n_368),
.B(n_238),
.Y(n_443)
);

AND2x2_ASAP7_75t_L g444 ( 
.A(n_363),
.B(n_238),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_409),
.Y(n_445)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_369),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_352),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_352),
.Y(n_448)
);

BUFx6f_ASAP7_75t_L g449 ( 
.A(n_369),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_364),
.Y(n_450)
);

HB1xp67_ASAP7_75t_L g451 ( 
.A(n_383),
.Y(n_451)
);

INVxp33_ASAP7_75t_SL g452 ( 
.A(n_353),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_364),
.Y(n_453)
);

OAI22xp5_ASAP7_75t_L g454 ( 
.A1(n_350),
.A2(n_234),
.B1(n_331),
.B2(n_333),
.Y(n_454)
);

BUFx6f_ASAP7_75t_L g455 ( 
.A(n_369),
.Y(n_455)
);

AND2x4_ASAP7_75t_L g456 ( 
.A(n_365),
.B(n_306),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_365),
.Y(n_457)
);

NAND2xp33_ASAP7_75t_L g458 ( 
.A(n_408),
.B(n_189),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_428),
.Y(n_459)
);

INVx3_ASAP7_75t_L g460 ( 
.A(n_369),
.Y(n_460)
);

BUFx6f_ASAP7_75t_L g461 ( 
.A(n_369),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_428),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_429),
.Y(n_463)
);

INVx2_ASAP7_75t_L g464 ( 
.A(n_412),
.Y(n_464)
);

AND2x2_ASAP7_75t_L g465 ( 
.A(n_410),
.B(n_306),
.Y(n_465)
);

NOR2xp33_ASAP7_75t_L g466 ( 
.A(n_358),
.B(n_349),
.Y(n_466)
);

INVx3_ASAP7_75t_L g467 ( 
.A(n_412),
.Y(n_467)
);

OAI22xp5_ASAP7_75t_L g468 ( 
.A1(n_416),
.A2(n_318),
.B1(n_339),
.B2(n_316),
.Y(n_468)
);

CKINVDCx5p33_ASAP7_75t_R g469 ( 
.A(n_425),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_429),
.Y(n_470)
);

INVx2_ASAP7_75t_L g471 ( 
.A(n_430),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_430),
.Y(n_472)
);

AND2x2_ASAP7_75t_L g473 ( 
.A(n_414),
.B(n_230),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_436),
.Y(n_474)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_436),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_379),
.Y(n_476)
);

BUFx3_ASAP7_75t_L g477 ( 
.A(n_415),
.Y(n_477)
);

BUFx2_ASAP7_75t_L g478 ( 
.A(n_353),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_379),
.Y(n_479)
);

BUFx6f_ASAP7_75t_L g480 ( 
.A(n_366),
.Y(n_480)
);

INVx2_ASAP7_75t_L g481 ( 
.A(n_366),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_367),
.Y(n_482)
);

BUFx2_ASAP7_75t_L g483 ( 
.A(n_381),
.Y(n_483)
);

OAI22xp5_ASAP7_75t_L g484 ( 
.A1(n_371),
.A2(n_206),
.B1(n_255),
.B2(n_246),
.Y(n_484)
);

AND2x2_ASAP7_75t_L g485 ( 
.A(n_417),
.B(n_237),
.Y(n_485)
);

INVx3_ASAP7_75t_L g486 ( 
.A(n_367),
.Y(n_486)
);

CKINVDCx5p33_ASAP7_75t_R g487 ( 
.A(n_433),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_372),
.Y(n_488)
);

INVx3_ASAP7_75t_L g489 ( 
.A(n_372),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_419),
.B(n_175),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_374),
.Y(n_491)
);

INVxp67_ASAP7_75t_L g492 ( 
.A(n_385),
.Y(n_492)
);

NAND2xp33_ASAP7_75t_SL g493 ( 
.A(n_361),
.B(n_184),
.Y(n_493)
);

INVx3_ASAP7_75t_L g494 ( 
.A(n_374),
.Y(n_494)
);

CKINVDCx20_ASAP7_75t_R g495 ( 
.A(n_356),
.Y(n_495)
);

INVx2_ASAP7_75t_L g496 ( 
.A(n_375),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_375),
.Y(n_497)
);

AND2x4_ASAP7_75t_L g498 ( 
.A(n_420),
.B(n_240),
.Y(n_498)
);

AND2x4_ASAP7_75t_L g499 ( 
.A(n_421),
.B(n_253),
.Y(n_499)
);

CKINVDCx20_ASAP7_75t_R g500 ( 
.A(n_370),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_378),
.Y(n_501)
);

AND2x6_ASAP7_75t_L g502 ( 
.A(n_378),
.B(n_189),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_382),
.Y(n_503)
);

INVx2_ASAP7_75t_L g504 ( 
.A(n_386),
.Y(n_504)
);

CKINVDCx20_ASAP7_75t_R g505 ( 
.A(n_376),
.Y(n_505)
);

INVx2_ASAP7_75t_L g506 ( 
.A(n_387),
.Y(n_506)
);

INVx2_ASAP7_75t_L g507 ( 
.A(n_388),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_389),
.Y(n_508)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_391),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_393),
.Y(n_510)
);

BUFx6f_ASAP7_75t_L g511 ( 
.A(n_394),
.Y(n_511)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_396),
.Y(n_512)
);

CKINVDCx5p33_ASAP7_75t_R g513 ( 
.A(n_434),
.Y(n_513)
);

AND2x4_ASAP7_75t_L g514 ( 
.A(n_355),
.B(n_254),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_399),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_401),
.Y(n_516)
);

INVx2_ASAP7_75t_L g517 ( 
.A(n_402),
.Y(n_517)
);

NOR2xp33_ASAP7_75t_L g518 ( 
.A(n_362),
.B(n_180),
.Y(n_518)
);

INVx3_ASAP7_75t_L g519 ( 
.A(n_403),
.Y(n_519)
);

NOR2xp33_ASAP7_75t_L g520 ( 
.A(n_518),
.B(n_373),
.Y(n_520)
);

AOI21x1_ASAP7_75t_L g521 ( 
.A1(n_456),
.A2(n_261),
.B(n_260),
.Y(n_521)
);

INVx2_ASAP7_75t_SL g522 ( 
.A(n_451),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_L g523 ( 
.A(n_444),
.B(n_381),
.Y(n_523)
);

INVxp67_ASAP7_75t_L g524 ( 
.A(n_518),
.Y(n_524)
);

BUFx3_ASAP7_75t_L g525 ( 
.A(n_477),
.Y(n_525)
);

INVxp67_ASAP7_75t_SL g526 ( 
.A(n_460),
.Y(n_526)
);

AOI22xp33_ASAP7_75t_SL g527 ( 
.A1(n_468),
.A2(n_424),
.B1(n_437),
.B2(n_354),
.Y(n_527)
);

INVx2_ASAP7_75t_L g528 ( 
.A(n_464),
.Y(n_528)
);

INVx2_ASAP7_75t_L g529 ( 
.A(n_464),
.Y(n_529)
);

INVx2_ASAP7_75t_L g530 ( 
.A(n_464),
.Y(n_530)
);

INVxp33_ASAP7_75t_SL g531 ( 
.A(n_469),
.Y(n_531)
);

NOR2xp33_ASAP7_75t_L g532 ( 
.A(n_466),
.B(n_440),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_444),
.B(n_384),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_519),
.Y(n_534)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_464),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_519),
.Y(n_536)
);

INVx2_ASAP7_75t_L g537 ( 
.A(n_441),
.Y(n_537)
);

INVx1_ASAP7_75t_SL g538 ( 
.A(n_495),
.Y(n_538)
);

INVx2_ASAP7_75t_SL g539 ( 
.A(n_451),
.Y(n_539)
);

INVx2_ASAP7_75t_L g540 ( 
.A(n_441),
.Y(n_540)
);

INVx4_ASAP7_75t_L g541 ( 
.A(n_467),
.Y(n_541)
);

NOR3xp33_ASAP7_75t_L g542 ( 
.A(n_454),
.B(n_431),
.C(n_426),
.Y(n_542)
);

INVx4_ASAP7_75t_L g543 ( 
.A(n_467),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_519),
.Y(n_544)
);

BUFx6f_ASAP7_75t_SL g545 ( 
.A(n_514),
.Y(n_545)
);

AND2x2_ASAP7_75t_L g546 ( 
.A(n_443),
.B(n_357),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_519),
.Y(n_547)
);

OR2x6_ASAP7_75t_L g548 ( 
.A(n_514),
.B(n_269),
.Y(n_548)
);

BUFx2_ASAP7_75t_L g549 ( 
.A(n_493),
.Y(n_549)
);

CKINVDCx5p33_ASAP7_75t_R g550 ( 
.A(n_487),
.Y(n_550)
);

BUFx6f_ASAP7_75t_L g551 ( 
.A(n_449),
.Y(n_551)
);

CKINVDCx20_ASAP7_75t_R g552 ( 
.A(n_495),
.Y(n_552)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_442),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_SL g554 ( 
.A(n_466),
.B(n_384),
.Y(n_554)
);

NAND3xp33_ASAP7_75t_L g555 ( 
.A(n_443),
.B(n_406),
.C(n_405),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_519),
.Y(n_556)
);

INVx2_ASAP7_75t_L g557 ( 
.A(n_442),
.Y(n_557)
);

INVx4_ASAP7_75t_L g558 ( 
.A(n_467),
.Y(n_558)
);

INVx2_ASAP7_75t_L g559 ( 
.A(n_447),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_SL g560 ( 
.A(n_493),
.B(n_390),
.Y(n_560)
);

INVx2_ASAP7_75t_L g561 ( 
.A(n_447),
.Y(n_561)
);

INVx3_ASAP7_75t_L g562 ( 
.A(n_449),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_SL g563 ( 
.A(n_492),
.B(n_390),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_448),
.Y(n_564)
);

CKINVDCx5p33_ASAP7_75t_R g565 ( 
.A(n_513),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_448),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_450),
.Y(n_567)
);

INVx2_ASAP7_75t_L g568 ( 
.A(n_450),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_453),
.Y(n_569)
);

AND2x2_ASAP7_75t_L g570 ( 
.A(n_443),
.B(n_359),
.Y(n_570)
);

INVx2_ASAP7_75t_L g571 ( 
.A(n_453),
.Y(n_571)
);

INVx3_ASAP7_75t_L g572 ( 
.A(n_449),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_457),
.Y(n_573)
);

INVxp33_ASAP7_75t_L g574 ( 
.A(n_454),
.Y(n_574)
);

INVx2_ASAP7_75t_L g575 ( 
.A(n_457),
.Y(n_575)
);

INVx3_ASAP7_75t_L g576 ( 
.A(n_449),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_456),
.Y(n_577)
);

INVx4_ASAP7_75t_L g578 ( 
.A(n_467),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_L g579 ( 
.A(n_444),
.B(n_395),
.Y(n_579)
);

INVx2_ASAP7_75t_L g580 ( 
.A(n_496),
.Y(n_580)
);

INVx3_ASAP7_75t_L g581 ( 
.A(n_449),
.Y(n_581)
);

INVx2_ASAP7_75t_L g582 ( 
.A(n_467),
.Y(n_582)
);

AND2x6_ASAP7_75t_L g583 ( 
.A(n_473),
.B(n_189),
.Y(n_583)
);

INVx3_ASAP7_75t_L g584 ( 
.A(n_449),
.Y(n_584)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_496),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_456),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_456),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_456),
.Y(n_588)
);

INVx2_ASAP7_75t_L g589 ( 
.A(n_496),
.Y(n_589)
);

INVx2_ASAP7_75t_L g590 ( 
.A(n_496),
.Y(n_590)
);

OR2x6_ASAP7_75t_L g591 ( 
.A(n_514),
.B(n_273),
.Y(n_591)
);

INVx2_ASAP7_75t_L g592 ( 
.A(n_497),
.Y(n_592)
);

INVx5_ASAP7_75t_L g593 ( 
.A(n_502),
.Y(n_593)
);

XNOR2xp5_ASAP7_75t_L g594 ( 
.A(n_468),
.B(n_377),
.Y(n_594)
);

AND2x2_ASAP7_75t_SL g595 ( 
.A(n_483),
.B(n_189),
.Y(n_595)
);

AND3x2_ASAP7_75t_L g596 ( 
.A(n_478),
.B(n_186),
.C(n_483),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_SL g597 ( 
.A(n_492),
.B(n_395),
.Y(n_597)
);

BUFx6f_ASAP7_75t_L g598 ( 
.A(n_449),
.Y(n_598)
);

INVx2_ASAP7_75t_L g599 ( 
.A(n_497),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_477),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_477),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_477),
.Y(n_602)
);

INVx2_ASAP7_75t_SL g603 ( 
.A(n_490),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_SL g604 ( 
.A(n_483),
.B(n_398),
.Y(n_604)
);

INVx2_ASAP7_75t_SL g605 ( 
.A(n_490),
.Y(n_605)
);

INVx2_ASAP7_75t_L g606 ( 
.A(n_497),
.Y(n_606)
);

CKINVDCx20_ASAP7_75t_R g607 ( 
.A(n_500),
.Y(n_607)
);

AO22x2_ASAP7_75t_L g608 ( 
.A1(n_484),
.A2(n_290),
.B1(n_308),
.B2(n_305),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_504),
.Y(n_609)
);

INVx2_ASAP7_75t_SL g610 ( 
.A(n_473),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_504),
.Y(n_611)
);

AOI21x1_ASAP7_75t_L g612 ( 
.A1(n_465),
.A2(n_294),
.B(n_287),
.Y(n_612)
);

BUFx6f_ASAP7_75t_L g613 ( 
.A(n_449),
.Y(n_613)
);

BUFx2_ASAP7_75t_L g614 ( 
.A(n_478),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_504),
.Y(n_615)
);

INVx3_ASAP7_75t_L g616 ( 
.A(n_455),
.Y(n_616)
);

CKINVDCx5p33_ASAP7_75t_R g617 ( 
.A(n_500),
.Y(n_617)
);

INVx2_ASAP7_75t_L g618 ( 
.A(n_497),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_504),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_506),
.Y(n_620)
);

CKINVDCx6p67_ASAP7_75t_R g621 ( 
.A(n_505),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_506),
.Y(n_622)
);

INVx4_ASAP7_75t_L g623 ( 
.A(n_455),
.Y(n_623)
);

BUFx6f_ASAP7_75t_L g624 ( 
.A(n_455),
.Y(n_624)
);

INVx2_ASAP7_75t_L g625 ( 
.A(n_480),
.Y(n_625)
);

BUFx2_ASAP7_75t_L g626 ( 
.A(n_478),
.Y(n_626)
);

INVx2_ASAP7_75t_L g627 ( 
.A(n_480),
.Y(n_627)
);

AOI22xp33_ASAP7_75t_L g628 ( 
.A1(n_514),
.A2(n_411),
.B1(n_407),
.B2(n_360),
.Y(n_628)
);

INVx3_ASAP7_75t_L g629 ( 
.A(n_455),
.Y(n_629)
);

INVx2_ASAP7_75t_SL g630 ( 
.A(n_473),
.Y(n_630)
);

INVx2_ASAP7_75t_L g631 ( 
.A(n_480),
.Y(n_631)
);

AND2x2_ASAP7_75t_L g632 ( 
.A(n_514),
.B(n_422),
.Y(n_632)
);

INVx2_ASAP7_75t_L g633 ( 
.A(n_480),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_L g634 ( 
.A(n_485),
.B(n_398),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_506),
.Y(n_635)
);

NOR2xp33_ASAP7_75t_L g636 ( 
.A(n_452),
.B(n_400),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_506),
.Y(n_637)
);

NOR2xp33_ASAP7_75t_L g638 ( 
.A(n_498),
.B(n_404),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_507),
.Y(n_639)
);

NOR2xp33_ASAP7_75t_L g640 ( 
.A(n_498),
.B(n_404),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_507),
.Y(n_641)
);

NOR2xp33_ASAP7_75t_L g642 ( 
.A(n_498),
.B(n_413),
.Y(n_642)
);

INVx3_ASAP7_75t_L g643 ( 
.A(n_455),
.Y(n_643)
);

INVx2_ASAP7_75t_L g644 ( 
.A(n_480),
.Y(n_644)
);

BUFx6f_ASAP7_75t_L g645 ( 
.A(n_455),
.Y(n_645)
);

AOI22xp33_ASAP7_75t_L g646 ( 
.A1(n_485),
.A2(n_286),
.B1(n_311),
.B2(n_323),
.Y(n_646)
);

NOR2xp33_ASAP7_75t_L g647 ( 
.A(n_498),
.B(n_413),
.Y(n_647)
);

CKINVDCx5p33_ASAP7_75t_R g648 ( 
.A(n_505),
.Y(n_648)
);

INVx2_ASAP7_75t_L g649 ( 
.A(n_480),
.Y(n_649)
);

INVx2_ASAP7_75t_L g650 ( 
.A(n_480),
.Y(n_650)
);

NOR2xp33_ASAP7_75t_L g651 ( 
.A(n_499),
.B(n_418),
.Y(n_651)
);

NOR2xp33_ASAP7_75t_L g652 ( 
.A(n_499),
.B(n_418),
.Y(n_652)
);

INVxp33_ASAP7_75t_SL g653 ( 
.A(n_445),
.Y(n_653)
);

NAND2xp33_ASAP7_75t_SL g654 ( 
.A(n_484),
.B(n_427),
.Y(n_654)
);

INVx3_ASAP7_75t_L g655 ( 
.A(n_455),
.Y(n_655)
);

BUFx6f_ASAP7_75t_SL g656 ( 
.A(n_499),
.Y(n_656)
);

AOI22xp5_ASAP7_75t_L g657 ( 
.A1(n_499),
.A2(n_317),
.B1(n_210),
.B2(n_209),
.Y(n_657)
);

INVx2_ASAP7_75t_L g658 ( 
.A(n_480),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_507),
.Y(n_659)
);

INVx2_ASAP7_75t_L g660 ( 
.A(n_471),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_507),
.Y(n_661)
);

INVx2_ASAP7_75t_L g662 ( 
.A(n_471),
.Y(n_662)
);

INVx5_ASAP7_75t_L g663 ( 
.A(n_502),
.Y(n_663)
);

CKINVDCx5p33_ASAP7_75t_R g664 ( 
.A(n_499),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_509),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_L g666 ( 
.A(n_485),
.B(n_427),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_SL g667 ( 
.A(n_503),
.B(n_432),
.Y(n_667)
);

AOI22xp33_ASAP7_75t_L g668 ( 
.A1(n_465),
.A2(n_311),
.B1(n_286),
.B2(n_300),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_509),
.Y(n_669)
);

AOI22xp33_ASAP7_75t_SL g670 ( 
.A1(n_465),
.A2(n_380),
.B1(n_392),
.B2(n_397),
.Y(n_670)
);

INVx2_ASAP7_75t_L g671 ( 
.A(n_471),
.Y(n_671)
);

INVx2_ASAP7_75t_L g672 ( 
.A(n_537),
.Y(n_672)
);

INVxp67_ASAP7_75t_L g673 ( 
.A(n_532),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_577),
.Y(n_674)
);

NOR2xp33_ASAP7_75t_L g675 ( 
.A(n_524),
.B(n_603),
.Y(n_675)
);

INVx2_ASAP7_75t_L g676 ( 
.A(n_537),
.Y(n_676)
);

AND2x2_ASAP7_75t_SL g677 ( 
.A(n_595),
.B(n_286),
.Y(n_677)
);

AND2x2_ASAP7_75t_L g678 ( 
.A(n_610),
.B(n_503),
.Y(n_678)
);

INVx4_ASAP7_75t_L g679 ( 
.A(n_541),
.Y(n_679)
);

NAND2xp33_ASAP7_75t_SL g680 ( 
.A(n_603),
.B(n_286),
.Y(n_680)
);

BUFx6f_ASAP7_75t_L g681 ( 
.A(n_525),
.Y(n_681)
);

NAND2xp33_ASAP7_75t_SL g682 ( 
.A(n_605),
.B(n_286),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_605),
.B(n_511),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_600),
.Y(n_684)
);

NOR2xp33_ASAP7_75t_L g685 ( 
.A(n_520),
.B(n_432),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_577),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_610),
.B(n_511),
.Y(n_687)
);

AND2x2_ASAP7_75t_L g688 ( 
.A(n_630),
.B(n_508),
.Y(n_688)
);

AO22x2_ASAP7_75t_L g689 ( 
.A1(n_554),
.A2(n_338),
.B1(n_297),
.B2(n_312),
.Y(n_689)
);

A2O1A1Ixp33_ASAP7_75t_L g690 ( 
.A1(n_630),
.A2(n_476),
.B(n_479),
.C(n_515),
.Y(n_690)
);

INVx2_ASAP7_75t_L g691 ( 
.A(n_540),
.Y(n_691)
);

O2A1O1Ixp33_ASAP7_75t_L g692 ( 
.A1(n_523),
.A2(n_476),
.B(n_479),
.C(n_515),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_L g693 ( 
.A(n_595),
.B(n_511),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_SL g694 ( 
.A(n_595),
.B(n_435),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_600),
.B(n_511),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_SL g696 ( 
.A(n_533),
.B(n_435),
.Y(n_696)
);

BUFx3_ASAP7_75t_L g697 ( 
.A(n_525),
.Y(n_697)
);

INVxp67_ASAP7_75t_L g698 ( 
.A(n_614),
.Y(n_698)
);

NOR3xp33_ASAP7_75t_L g699 ( 
.A(n_604),
.B(n_439),
.C(n_438),
.Y(n_699)
);

O2A1O1Ixp33_ASAP7_75t_L g700 ( 
.A1(n_579),
.A2(n_508),
.B(n_516),
.C(n_510),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_601),
.B(n_511),
.Y(n_701)
);

INVx4_ASAP7_75t_L g702 ( 
.A(n_541),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_L g703 ( 
.A(n_601),
.B(n_511),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_L g704 ( 
.A(n_602),
.B(n_511),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_SL g705 ( 
.A(n_634),
.B(n_438),
.Y(n_705)
);

INVx2_ASAP7_75t_L g706 ( 
.A(n_540),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_SL g707 ( 
.A(n_666),
.B(n_439),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_L g708 ( 
.A(n_602),
.B(n_486),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_586),
.B(n_486),
.Y(n_709)
);

INVx2_ASAP7_75t_L g710 ( 
.A(n_553),
.Y(n_710)
);

INVx2_ASAP7_75t_L g711 ( 
.A(n_553),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_SL g712 ( 
.A(n_664),
.B(n_175),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_587),
.Y(n_713)
);

NOR2xp33_ASAP7_75t_L g714 ( 
.A(n_563),
.B(n_597),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_L g715 ( 
.A(n_587),
.B(n_486),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_588),
.B(n_486),
.Y(n_716)
);

INVx2_ASAP7_75t_SL g717 ( 
.A(n_546),
.Y(n_717)
);

AOI221xp5_ASAP7_75t_L g718 ( 
.A1(n_574),
.A2(n_320),
.B1(n_191),
.B2(n_192),
.C(n_194),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_588),
.Y(n_719)
);

INVx2_ASAP7_75t_L g720 ( 
.A(n_557),
.Y(n_720)
);

INVx2_ASAP7_75t_SL g721 ( 
.A(n_546),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_564),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_L g723 ( 
.A(n_564),
.B(n_486),
.Y(n_723)
);

AOI22xp33_ASAP7_75t_L g724 ( 
.A1(n_632),
.A2(n_296),
.B1(n_311),
.B2(n_509),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_L g725 ( 
.A(n_566),
.B(n_489),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_L g726 ( 
.A(n_566),
.B(n_489),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_SL g727 ( 
.A(n_664),
.B(n_176),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_L g728 ( 
.A(n_567),
.B(n_573),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_SL g729 ( 
.A(n_638),
.B(n_176),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_SL g730 ( 
.A(n_640),
.B(n_181),
.Y(n_730)
);

NOR2xp33_ASAP7_75t_L g731 ( 
.A(n_636),
.B(n_213),
.Y(n_731)
);

AND2x2_ASAP7_75t_L g732 ( 
.A(n_570),
.B(n_632),
.Y(n_732)
);

AND2x4_ASAP7_75t_L g733 ( 
.A(n_525),
.B(n_510),
.Y(n_733)
);

INVx2_ASAP7_75t_L g734 ( 
.A(n_559),
.Y(n_734)
);

INVx2_ASAP7_75t_L g735 ( 
.A(n_559),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_L g736 ( 
.A(n_567),
.B(n_489),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_SL g737 ( 
.A(n_642),
.B(n_181),
.Y(n_737)
);

O2A1O1Ixp33_ASAP7_75t_L g738 ( 
.A1(n_570),
.A2(n_516),
.B(n_458),
.C(n_512),
.Y(n_738)
);

AOI22xp33_ASAP7_75t_L g739 ( 
.A1(n_573),
.A2(n_296),
.B1(n_311),
.B2(n_509),
.Y(n_739)
);

INVx2_ASAP7_75t_L g740 ( 
.A(n_561),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_561),
.Y(n_741)
);

INVx2_ASAP7_75t_L g742 ( 
.A(n_568),
.Y(n_742)
);

NOR2xp33_ASAP7_75t_L g743 ( 
.A(n_647),
.B(n_281),
.Y(n_743)
);

INVx2_ASAP7_75t_L g744 ( 
.A(n_568),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_SL g745 ( 
.A(n_651),
.B(n_188),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_L g746 ( 
.A(n_526),
.B(n_489),
.Y(n_746)
);

NAND3xp33_ASAP7_75t_L g747 ( 
.A(n_652),
.B(n_275),
.C(n_272),
.Y(n_747)
);

NAND2xp33_ASAP7_75t_L g748 ( 
.A(n_646),
.B(n_668),
.Y(n_748)
);

INVxp67_ASAP7_75t_L g749 ( 
.A(n_614),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_SL g750 ( 
.A(n_522),
.B(n_188),
.Y(n_750)
);

INVx2_ASAP7_75t_L g751 ( 
.A(n_569),
.Y(n_751)
);

OAI221xp5_ASAP7_75t_L g752 ( 
.A1(n_657),
.A2(n_309),
.B1(n_512),
.B2(n_517),
.C(n_463),
.Y(n_752)
);

NOR2xp33_ASAP7_75t_L g753 ( 
.A(n_549),
.B(n_190),
.Y(n_753)
);

NAND3xp33_ASAP7_75t_L g754 ( 
.A(n_628),
.B(n_289),
.C(n_283),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_SL g755 ( 
.A(n_539),
.B(n_190),
.Y(n_755)
);

NOR2xp67_ASAP7_75t_L g756 ( 
.A(n_555),
.B(n_512),
.Y(n_756)
);

NOR2xp33_ASAP7_75t_L g757 ( 
.A(n_667),
.B(n_193),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_569),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_571),
.Y(n_759)
);

NAND3x1_ASAP7_75t_L g760 ( 
.A(n_542),
.B(n_423),
.C(n_422),
.Y(n_760)
);

AOI22xp33_ASAP7_75t_L g761 ( 
.A1(n_548),
.A2(n_296),
.B1(n_517),
.B2(n_494),
.Y(n_761)
);

NOR2xp33_ASAP7_75t_L g762 ( 
.A(n_560),
.B(n_193),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_571),
.Y(n_763)
);

AOI22xp33_ASAP7_75t_L g764 ( 
.A1(n_548),
.A2(n_296),
.B1(n_517),
.B2(n_494),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_SL g765 ( 
.A(n_527),
.B(n_196),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_SL g766 ( 
.A(n_657),
.B(n_196),
.Y(n_766)
);

INVx3_ASAP7_75t_L g767 ( 
.A(n_541),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_575),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_L g769 ( 
.A(n_534),
.B(n_489),
.Y(n_769)
);

INVx2_ASAP7_75t_L g770 ( 
.A(n_575),
.Y(n_770)
);

HB1xp67_ASAP7_75t_L g771 ( 
.A(n_626),
.Y(n_771)
);

NAND3xp33_ASAP7_75t_L g772 ( 
.A(n_654),
.B(n_295),
.C(n_291),
.Y(n_772)
);

OAI22xp5_ASAP7_75t_L g773 ( 
.A1(n_656),
.A2(n_200),
.B1(n_322),
.B2(n_330),
.Y(n_773)
);

CKINVDCx5p33_ASAP7_75t_R g774 ( 
.A(n_550),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_609),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_534),
.B(n_494),
.Y(n_776)
);

INVxp67_ASAP7_75t_L g777 ( 
.A(n_626),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_L g778 ( 
.A(n_536),
.B(n_494),
.Y(n_778)
);

NOR2xp33_ASAP7_75t_L g779 ( 
.A(n_531),
.B(n_198),
.Y(n_779)
);

AND2x4_ASAP7_75t_L g780 ( 
.A(n_548),
.B(n_517),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_536),
.B(n_494),
.Y(n_781)
);

AND2x2_ASAP7_75t_L g782 ( 
.A(n_555),
.B(n_459),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_L g783 ( 
.A(n_544),
.B(n_547),
.Y(n_783)
);

NOR2xp33_ASAP7_75t_L g784 ( 
.A(n_653),
.B(n_198),
.Y(n_784)
);

INVx2_ASAP7_75t_L g785 ( 
.A(n_528),
.Y(n_785)
);

NOR2xp33_ASAP7_75t_L g786 ( 
.A(n_596),
.B(n_199),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_L g787 ( 
.A(n_544),
.B(n_460),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_L g788 ( 
.A(n_547),
.B(n_460),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_SL g789 ( 
.A(n_670),
.B(n_199),
.Y(n_789)
);

AOI21xp5_ASAP7_75t_L g790 ( 
.A1(n_541),
.A2(n_455),
.B(n_461),
.Y(n_790)
);

INVx2_ASAP7_75t_L g791 ( 
.A(n_528),
.Y(n_791)
);

AOI22xp33_ASAP7_75t_L g792 ( 
.A1(n_548),
.A2(n_296),
.B1(n_502),
.B2(n_471),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_L g793 ( 
.A(n_556),
.B(n_460),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_609),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_L g795 ( 
.A(n_556),
.B(n_460),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_L g796 ( 
.A(n_543),
.B(n_558),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_543),
.B(n_462),
.Y(n_797)
);

INVx2_ASAP7_75t_L g798 ( 
.A(n_529),
.Y(n_798)
);

NOR3xp33_ASAP7_75t_L g799 ( 
.A(n_538),
.B(n_423),
.C(n_348),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_SL g800 ( 
.A(n_543),
.B(n_200),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_611),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_SL g802 ( 
.A(n_543),
.B(n_202),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_L g803 ( 
.A(n_558),
.B(n_462),
.Y(n_803)
);

OAI22x1_ASAP7_75t_SL g804 ( 
.A1(n_617),
.A2(n_210),
.B1(n_209),
.B2(n_302),
.Y(n_804)
);

AND2x2_ASAP7_75t_L g805 ( 
.A(n_608),
.B(n_463),
.Y(n_805)
);

OR2x2_ASAP7_75t_L g806 ( 
.A(n_594),
.B(n_191),
.Y(n_806)
);

AND2x2_ASAP7_75t_L g807 ( 
.A(n_608),
.B(n_470),
.Y(n_807)
);

NOR3xp33_ASAP7_75t_L g808 ( 
.A(n_617),
.B(n_299),
.C(n_298),
.Y(n_808)
);

INVx2_ASAP7_75t_SL g809 ( 
.A(n_548),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_558),
.B(n_470),
.Y(n_810)
);

INVx2_ASAP7_75t_L g811 ( 
.A(n_529),
.Y(n_811)
);

NOR2xp33_ASAP7_75t_L g812 ( 
.A(n_558),
.B(n_202),
.Y(n_812)
);

BUFx2_ASAP7_75t_L g813 ( 
.A(n_552),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_611),
.Y(n_814)
);

INVx2_ASAP7_75t_L g815 ( 
.A(n_530),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_SL g816 ( 
.A(n_578),
.B(n_205),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_615),
.Y(n_817)
);

BUFx6f_ASAP7_75t_L g818 ( 
.A(n_551),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_L g819 ( 
.A(n_578),
.B(n_472),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_L g820 ( 
.A(n_578),
.B(n_474),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_SL g821 ( 
.A(n_550),
.B(n_205),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_SL g822 ( 
.A(n_565),
.B(n_303),
.Y(n_822)
);

BUFx6f_ASAP7_75t_L g823 ( 
.A(n_551),
.Y(n_823)
);

AND2x2_ASAP7_75t_L g824 ( 
.A(n_608),
.B(n_474),
.Y(n_824)
);

BUFx8_ASAP7_75t_L g825 ( 
.A(n_545),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_615),
.Y(n_826)
);

INVx2_ASAP7_75t_L g827 ( 
.A(n_530),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_619),
.Y(n_828)
);

NOR2xp33_ASAP7_75t_L g829 ( 
.A(n_565),
.B(n_303),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_SL g830 ( 
.A(n_594),
.B(n_322),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_562),
.B(n_446),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_L g832 ( 
.A(n_562),
.B(n_446),
.Y(n_832)
);

INVx2_ASAP7_75t_L g833 ( 
.A(n_535),
.Y(n_833)
);

INVx2_ASAP7_75t_L g834 ( 
.A(n_535),
.Y(n_834)
);

INVx2_ASAP7_75t_SL g835 ( 
.A(n_591),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_619),
.Y(n_836)
);

INVx2_ASAP7_75t_SL g837 ( 
.A(n_591),
.Y(n_837)
);

CKINVDCx5p33_ASAP7_75t_R g838 ( 
.A(n_774),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_L g839 ( 
.A(n_743),
.B(n_675),
.Y(n_839)
);

BUFx6f_ASAP7_75t_L g840 ( 
.A(n_681),
.Y(n_840)
);

INVx2_ASAP7_75t_L g841 ( 
.A(n_672),
.Y(n_841)
);

INVx2_ASAP7_75t_L g842 ( 
.A(n_672),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_SL g843 ( 
.A(n_677),
.B(n_593),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_L g844 ( 
.A(n_677),
.B(n_591),
.Y(n_844)
);

BUFx6f_ASAP7_75t_L g845 ( 
.A(n_681),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_SL g846 ( 
.A(n_767),
.B(n_679),
.Y(n_846)
);

INVx3_ASAP7_75t_L g847 ( 
.A(n_681),
.Y(n_847)
);

NOR2xp33_ASAP7_75t_L g848 ( 
.A(n_673),
.B(n_591),
.Y(n_848)
);

INVx2_ASAP7_75t_L g849 ( 
.A(n_676),
.Y(n_849)
);

AND2x4_ASAP7_75t_L g850 ( 
.A(n_717),
.B(n_591),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_SL g851 ( 
.A(n_767),
.B(n_593),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_674),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_674),
.Y(n_853)
);

OR2x6_ASAP7_75t_L g854 ( 
.A(n_813),
.B(n_608),
.Y(n_854)
);

INVx2_ASAP7_75t_SL g855 ( 
.A(n_771),
.Y(n_855)
);

INVx5_ASAP7_75t_L g856 ( 
.A(n_767),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_732),
.B(n_620),
.Y(n_857)
);

NOR2xp33_ASAP7_75t_L g858 ( 
.A(n_685),
.B(n_656),
.Y(n_858)
);

INVx2_ASAP7_75t_L g859 ( 
.A(n_676),
.Y(n_859)
);

AND2x6_ASAP7_75t_SL g860 ( 
.A(n_731),
.B(n_621),
.Y(n_860)
);

AOI22xp33_ASAP7_75t_L g861 ( 
.A1(n_689),
.A2(n_748),
.B1(n_732),
.B2(n_686),
.Y(n_861)
);

AND2x6_ASAP7_75t_SL g862 ( 
.A(n_829),
.B(n_607),
.Y(n_862)
);

CKINVDCx5p33_ASAP7_75t_R g863 ( 
.A(n_813),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_686),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_678),
.B(n_620),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_L g866 ( 
.A(n_678),
.B(n_622),
.Y(n_866)
);

NOR2xp67_ASAP7_75t_L g867 ( 
.A(n_747),
.B(n_648),
.Y(n_867)
);

BUFx6f_ASAP7_75t_L g868 ( 
.A(n_681),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_L g869 ( 
.A(n_688),
.B(n_622),
.Y(n_869)
);

BUFx3_ASAP7_75t_L g870 ( 
.A(n_825),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_713),
.Y(n_871)
);

INVxp67_ASAP7_75t_L g872 ( 
.A(n_750),
.Y(n_872)
);

OR2x2_ASAP7_75t_L g873 ( 
.A(n_806),
.B(n_648),
.Y(n_873)
);

AND2x4_ASAP7_75t_L g874 ( 
.A(n_717),
.B(n_482),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_L g875 ( 
.A(n_688),
.B(n_635),
.Y(n_875)
);

INVx3_ASAP7_75t_L g876 ( 
.A(n_681),
.Y(n_876)
);

NOR2xp33_ASAP7_75t_L g877 ( 
.A(n_698),
.B(n_656),
.Y(n_877)
);

NOR2xp33_ASAP7_75t_L g878 ( 
.A(n_749),
.B(n_545),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_719),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_SL g880 ( 
.A(n_679),
.B(n_593),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_759),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_L g882 ( 
.A(n_722),
.B(n_721),
.Y(n_882)
);

INVx2_ASAP7_75t_SL g883 ( 
.A(n_805),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_L g884 ( 
.A(n_721),
.B(n_635),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_L g885 ( 
.A(n_782),
.B(n_637),
.Y(n_885)
);

INVx1_ASAP7_75t_SL g886 ( 
.A(n_806),
.Y(n_886)
);

CKINVDCx5p33_ASAP7_75t_R g887 ( 
.A(n_825),
.Y(n_887)
);

INVxp67_ASAP7_75t_L g888 ( 
.A(n_755),
.Y(n_888)
);

AOI22xp5_ASAP7_75t_L g889 ( 
.A1(n_714),
.A2(n_545),
.B1(n_583),
.B2(n_665),
.Y(n_889)
);

BUFx2_ASAP7_75t_L g890 ( 
.A(n_777),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_SL g891 ( 
.A(n_679),
.B(n_593),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_L g892 ( 
.A(n_782),
.B(n_637),
.Y(n_892)
);

CKINVDCx5p33_ASAP7_75t_R g893 ( 
.A(n_825),
.Y(n_893)
);

INVx2_ASAP7_75t_L g894 ( 
.A(n_691),
.Y(n_894)
);

CKINVDCx20_ASAP7_75t_R g895 ( 
.A(n_830),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_L g896 ( 
.A(n_728),
.B(n_639),
.Y(n_896)
);

AND2x2_ASAP7_75t_L g897 ( 
.A(n_753),
.B(n_779),
.Y(n_897)
);

OAI22xp5_ASAP7_75t_SL g898 ( 
.A1(n_752),
.A2(n_784),
.B1(n_757),
.B2(n_786),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_SL g899 ( 
.A(n_702),
.B(n_593),
.Y(n_899)
);

CKINVDCx5p33_ASAP7_75t_R g900 ( 
.A(n_696),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_763),
.Y(n_901)
);

INVx2_ASAP7_75t_L g902 ( 
.A(n_706),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_SL g903 ( 
.A(n_702),
.B(n_593),
.Y(n_903)
);

INVx2_ASAP7_75t_L g904 ( 
.A(n_706),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_768),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_768),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_L g907 ( 
.A(n_733),
.B(n_756),
.Y(n_907)
);

INVx2_ASAP7_75t_L g908 ( 
.A(n_710),
.Y(n_908)
);

AOI22xp33_ASAP7_75t_L g909 ( 
.A1(n_689),
.A2(n_583),
.B1(n_669),
.B2(n_665),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_710),
.Y(n_910)
);

NOR2x2_ASAP7_75t_L g911 ( 
.A(n_766),
.B(n_228),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_SL g912 ( 
.A(n_702),
.B(n_663),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_L g913 ( 
.A(n_733),
.B(n_639),
.Y(n_913)
);

NOR2xp67_ASAP7_75t_L g914 ( 
.A(n_772),
.B(n_612),
.Y(n_914)
);

BUFx3_ASAP7_75t_L g915 ( 
.A(n_733),
.Y(n_915)
);

NAND3xp33_ASAP7_75t_SL g916 ( 
.A(n_718),
.B(n_194),
.C(n_192),
.Y(n_916)
);

AOI22xp33_ASAP7_75t_L g917 ( 
.A1(n_689),
.A2(n_583),
.B1(n_669),
.B2(n_641),
.Y(n_917)
);

INVx5_ASAP7_75t_L g918 ( 
.A(n_818),
.Y(n_918)
);

AOI22xp5_ASAP7_75t_L g919 ( 
.A1(n_694),
.A2(n_583),
.B1(n_661),
.B2(n_659),
.Y(n_919)
);

AND2x6_ASAP7_75t_SL g920 ( 
.A(n_762),
.B(n_488),
.Y(n_920)
);

AO22x1_ASAP7_75t_L g921 ( 
.A1(n_699),
.A2(n_328),
.B1(n_204),
.B2(n_302),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_SL g922 ( 
.A(n_780),
.B(n_663),
.Y(n_922)
);

NOR2xp33_ASAP7_75t_L g923 ( 
.A(n_705),
.B(n_641),
.Y(n_923)
);

CKINVDCx5p33_ASAP7_75t_R g924 ( 
.A(n_707),
.Y(n_924)
);

AND2x4_ASAP7_75t_L g925 ( 
.A(n_697),
.B(n_488),
.Y(n_925)
);

INVx4_ASAP7_75t_L g926 ( 
.A(n_697),
.Y(n_926)
);

NOR3xp33_ASAP7_75t_SL g927 ( 
.A(n_765),
.B(n_789),
.C(n_307),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_711),
.Y(n_928)
);

INVx2_ASAP7_75t_L g929 ( 
.A(n_711),
.Y(n_929)
);

INVx2_ASAP7_75t_L g930 ( 
.A(n_720),
.Y(n_930)
);

NAND2x1p5_ASAP7_75t_L g931 ( 
.A(n_780),
.B(n_663),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_L g932 ( 
.A(n_683),
.B(n_659),
.Y(n_932)
);

NOR2xp33_ASAP7_75t_L g933 ( 
.A(n_821),
.B(n_661),
.Y(n_933)
);

INVx2_ASAP7_75t_L g934 ( 
.A(n_720),
.Y(n_934)
);

AOI22xp5_ASAP7_75t_L g935 ( 
.A1(n_780),
.A2(n_583),
.B1(n_582),
.B2(n_633),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_L g936 ( 
.A(n_812),
.B(n_562),
.Y(n_936)
);

AOI21xp5_ASAP7_75t_L g937 ( 
.A1(n_796),
.A2(n_623),
.B(n_598),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_734),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_L g939 ( 
.A(n_690),
.B(n_572),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_L g940 ( 
.A(n_690),
.B(n_572),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_734),
.Y(n_941)
);

CKINVDCx20_ASAP7_75t_R g942 ( 
.A(n_822),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_735),
.Y(n_943)
);

NAND2x1p5_ASAP7_75t_L g944 ( 
.A(n_809),
.B(n_663),
.Y(n_944)
);

HB1xp67_ASAP7_75t_L g945 ( 
.A(n_805),
.Y(n_945)
);

NOR2x1p5_ASAP7_75t_L g946 ( 
.A(n_754),
.B(n_204),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_L g947 ( 
.A(n_684),
.B(n_572),
.Y(n_947)
);

INVx3_ASAP7_75t_L g948 ( 
.A(n_740),
.Y(n_948)
);

CKINVDCx20_ASAP7_75t_R g949 ( 
.A(n_729),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_L g950 ( 
.A(n_748),
.B(n_572),
.Y(n_950)
);

INVx3_ASAP7_75t_L g951 ( 
.A(n_740),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_742),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_SL g953 ( 
.A(n_693),
.B(n_663),
.Y(n_953)
);

BUFx3_ASAP7_75t_L g954 ( 
.A(n_809),
.Y(n_954)
);

AO22x1_ASAP7_75t_L g955 ( 
.A1(n_808),
.A2(n_799),
.B1(n_824),
.B2(n_807),
.Y(n_955)
);

NOR2x1p5_ASAP7_75t_L g956 ( 
.A(n_807),
.B(n_307),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_742),
.Y(n_957)
);

INVx3_ASAP7_75t_L g958 ( 
.A(n_744),
.Y(n_958)
);

AOI22xp5_ASAP7_75t_L g959 ( 
.A1(n_835),
.A2(n_583),
.B1(n_582),
.B2(n_625),
.Y(n_959)
);

BUFx12f_ASAP7_75t_L g960 ( 
.A(n_824),
.Y(n_960)
);

AO22x1_ASAP7_75t_L g961 ( 
.A1(n_835),
.A2(n_320),
.B1(n_310),
.B2(n_313),
.Y(n_961)
);

INVx2_ASAP7_75t_L g962 ( 
.A(n_744),
.Y(n_962)
);

BUFx2_ASAP7_75t_L g963 ( 
.A(n_760),
.Y(n_963)
);

INVx1_ASAP7_75t_L g964 ( 
.A(n_751),
.Y(n_964)
);

INVx1_ASAP7_75t_L g965 ( 
.A(n_751),
.Y(n_965)
);

AOI22xp33_ASAP7_75t_SL g966 ( 
.A1(n_689),
.A2(n_583),
.B1(n_228),
.B2(n_277),
.Y(n_966)
);

NOR2xp33_ASAP7_75t_L g967 ( 
.A(n_730),
.B(n_612),
.Y(n_967)
);

BUFx3_ASAP7_75t_L g968 ( 
.A(n_837),
.Y(n_968)
);

AND2x4_ASAP7_75t_L g969 ( 
.A(n_837),
.B(n_491),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_SL g970 ( 
.A(n_818),
.B(n_663),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_SL g971 ( 
.A(n_818),
.B(n_576),
.Y(n_971)
);

BUFx3_ASAP7_75t_L g972 ( 
.A(n_741),
.Y(n_972)
);

CKINVDCx5p33_ASAP7_75t_R g973 ( 
.A(n_804),
.Y(n_973)
);

CKINVDCx5p33_ASAP7_75t_R g974 ( 
.A(n_773),
.Y(n_974)
);

AOI22xp33_ASAP7_75t_L g975 ( 
.A1(n_770),
.A2(n_296),
.B1(n_662),
.B2(n_660),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_770),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_L g977 ( 
.A(n_758),
.B(n_576),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_L g978 ( 
.A(n_687),
.B(n_576),
.Y(n_978)
);

NAND2xp5_ASAP7_75t_L g979 ( 
.A(n_692),
.B(n_576),
.Y(n_979)
);

INVx2_ASAP7_75t_L g980 ( 
.A(n_785),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_SL g981 ( 
.A(n_818),
.B(n_581),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_SL g982 ( 
.A(n_818),
.B(n_581),
.Y(n_982)
);

NAND2x1p5_ASAP7_75t_L g983 ( 
.A(n_823),
.B(n_623),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_SL g984 ( 
.A(n_823),
.B(n_581),
.Y(n_984)
);

OR2x2_ASAP7_75t_SL g985 ( 
.A(n_760),
.B(n_228),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_SL g986 ( 
.A(n_823),
.B(n_581),
.Y(n_986)
);

HB1xp67_ASAP7_75t_L g987 ( 
.A(n_775),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_SL g988 ( 
.A(n_823),
.B(n_584),
.Y(n_988)
);

BUFx6f_ASAP7_75t_L g989 ( 
.A(n_823),
.Y(n_989)
);

INVx2_ASAP7_75t_L g990 ( 
.A(n_785),
.Y(n_990)
);

INVx2_ASAP7_75t_L g991 ( 
.A(n_791),
.Y(n_991)
);

OAI22xp5_ASAP7_75t_L g992 ( 
.A1(n_797),
.A2(n_330),
.B1(n_347),
.B2(n_341),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_SL g993 ( 
.A(n_709),
.B(n_584),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_L g994 ( 
.A(n_803),
.B(n_584),
.Y(n_994)
);

HB1xp67_ASAP7_75t_L g995 ( 
.A(n_794),
.Y(n_995)
);

BUFx6f_ASAP7_75t_L g996 ( 
.A(n_783),
.Y(n_996)
);

NOR2x2_ASAP7_75t_L g997 ( 
.A(n_737),
.B(n_277),
.Y(n_997)
);

AND2x4_ASAP7_75t_L g998 ( 
.A(n_712),
.B(n_491),
.Y(n_998)
);

NOR2xp33_ASAP7_75t_L g999 ( 
.A(n_745),
.B(n_623),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_SL g1000 ( 
.A(n_715),
.B(n_584),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_L g1001 ( 
.A(n_810),
.B(n_616),
.Y(n_1001)
);

INVx1_ASAP7_75t_L g1002 ( 
.A(n_794),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_L g1003 ( 
.A(n_819),
.B(n_616),
.Y(n_1003)
);

BUFx3_ASAP7_75t_L g1004 ( 
.A(n_801),
.Y(n_1004)
);

INVx1_ASAP7_75t_L g1005 ( 
.A(n_801),
.Y(n_1005)
);

HB1xp67_ASAP7_75t_L g1006 ( 
.A(n_814),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_814),
.Y(n_1007)
);

AND2x4_ASAP7_75t_L g1008 ( 
.A(n_727),
.B(n_501),
.Y(n_1008)
);

AOI22xp5_ASAP7_75t_L g1009 ( 
.A1(n_800),
.A2(n_582),
.B1(n_658),
.B2(n_625),
.Y(n_1009)
);

AOI22xp5_ASAP7_75t_L g1010 ( 
.A1(n_802),
.A2(n_644),
.B1(n_658),
.B2(n_631),
.Y(n_1010)
);

AND2x4_ASAP7_75t_L g1011 ( 
.A(n_817),
.B(n_501),
.Y(n_1011)
);

AOI22xp5_ASAP7_75t_L g1012 ( 
.A1(n_816),
.A2(n_627),
.B1(n_631),
.B2(n_650),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_L g1013 ( 
.A(n_820),
.B(n_616),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_L g1014 ( 
.A(n_700),
.B(n_616),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_L g1015 ( 
.A(n_817),
.B(n_629),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_L g1016 ( 
.A(n_826),
.B(n_629),
.Y(n_1016)
);

INVx1_ASAP7_75t_L g1017 ( 
.A(n_826),
.Y(n_1017)
);

INVx1_ASAP7_75t_L g1018 ( 
.A(n_836),
.Y(n_1018)
);

INVx1_ASAP7_75t_L g1019 ( 
.A(n_836),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_SL g1020 ( 
.A(n_716),
.B(n_629),
.Y(n_1020)
);

AOI22xp5_ASAP7_75t_L g1021 ( 
.A1(n_828),
.A2(n_627),
.B1(n_633),
.B2(n_650),
.Y(n_1021)
);

INVxp67_ASAP7_75t_L g1022 ( 
.A(n_890),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_L g1023 ( 
.A(n_839),
.B(n_746),
.Y(n_1023)
);

OR2x2_ASAP7_75t_L g1024 ( 
.A(n_886),
.B(n_723),
.Y(n_1024)
);

BUFx2_ASAP7_75t_L g1025 ( 
.A(n_863),
.Y(n_1025)
);

NAND2xp33_ASAP7_75t_L g1026 ( 
.A(n_856),
.B(n_725),
.Y(n_1026)
);

AOI21xp5_ASAP7_75t_L g1027 ( 
.A1(n_856),
.A2(n_790),
.B(n_623),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_L g1028 ( 
.A(n_885),
.B(n_726),
.Y(n_1028)
);

NOR2xp33_ASAP7_75t_L g1029 ( 
.A(n_898),
.B(n_736),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_L g1030 ( 
.A(n_892),
.B(n_791),
.Y(n_1030)
);

NOR2xp33_ASAP7_75t_L g1031 ( 
.A(n_872),
.B(n_769),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_SL g1032 ( 
.A(n_858),
.B(n_761),
.Y(n_1032)
);

NOR3xp33_ASAP7_75t_SL g1033 ( 
.A(n_974),
.B(n_313),
.C(n_310),
.Y(n_1033)
);

INVx1_ASAP7_75t_L g1034 ( 
.A(n_987),
.Y(n_1034)
);

BUFx3_ASAP7_75t_L g1035 ( 
.A(n_855),
.Y(n_1035)
);

INVx1_ASAP7_75t_L g1036 ( 
.A(n_987),
.Y(n_1036)
);

NAND2xp5_ASAP7_75t_SL g1037 ( 
.A(n_858),
.B(n_764),
.Y(n_1037)
);

INVx1_ASAP7_75t_L g1038 ( 
.A(n_995),
.Y(n_1038)
);

AOI21xp5_ASAP7_75t_L g1039 ( 
.A1(n_856),
.A2(n_701),
.B(n_695),
.Y(n_1039)
);

NOR2xp33_ASAP7_75t_SL g1040 ( 
.A(n_838),
.B(n_277),
.Y(n_1040)
);

OAI22xp5_ASAP7_75t_L g1041 ( 
.A1(n_861),
.A2(n_724),
.B1(n_739),
.B2(n_738),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_SL g1042 ( 
.A(n_848),
.B(n_680),
.Y(n_1042)
);

BUFx2_ASAP7_75t_SL g1043 ( 
.A(n_870),
.Y(n_1043)
);

NOR3xp33_ASAP7_75t_SL g1044 ( 
.A(n_973),
.B(n_328),
.C(n_317),
.Y(n_1044)
);

INVx3_ASAP7_75t_L g1045 ( 
.A(n_840),
.Y(n_1045)
);

OAI22xp5_ASAP7_75t_L g1046 ( 
.A1(n_861),
.A2(n_708),
.B1(n_792),
.B2(n_778),
.Y(n_1046)
);

AOI21xp5_ASAP7_75t_L g1047 ( 
.A1(n_846),
.A2(n_704),
.B(n_703),
.Y(n_1047)
);

HB1xp67_ASAP7_75t_L g1048 ( 
.A(n_945),
.Y(n_1048)
);

INVx2_ASAP7_75t_L g1049 ( 
.A(n_948),
.Y(n_1049)
);

INVx1_ASAP7_75t_SL g1050 ( 
.A(n_873),
.Y(n_1050)
);

O2A1O1Ixp33_ASAP7_75t_L g1051 ( 
.A1(n_916),
.A2(n_888),
.B(n_848),
.C(n_992),
.Y(n_1051)
);

NAND3xp33_ASAP7_75t_SL g1052 ( 
.A(n_900),
.B(n_335),
.C(n_336),
.Y(n_1052)
);

A2O1A1Ixp33_ASAP7_75t_SL g1053 ( 
.A1(n_967),
.A2(n_999),
.B(n_923),
.C(n_878),
.Y(n_1053)
);

AOI21xp5_ASAP7_75t_L g1054 ( 
.A1(n_846),
.A2(n_918),
.B(n_936),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_L g1055 ( 
.A(n_857),
.B(n_798),
.Y(n_1055)
);

O2A1O1Ixp33_ASAP7_75t_L g1056 ( 
.A1(n_882),
.A2(n_781),
.B(n_776),
.C(n_787),
.Y(n_1056)
);

INVx2_ASAP7_75t_L g1057 ( 
.A(n_948),
.Y(n_1057)
);

O2A1O1Ixp33_ASAP7_75t_L g1058 ( 
.A1(n_883),
.A2(n_788),
.B(n_793),
.C(n_795),
.Y(n_1058)
);

INVx2_ASAP7_75t_L g1059 ( 
.A(n_951),
.Y(n_1059)
);

INVx1_ASAP7_75t_L g1060 ( 
.A(n_995),
.Y(n_1060)
);

INVx3_ASAP7_75t_L g1061 ( 
.A(n_840),
.Y(n_1061)
);

OAI22xp5_ASAP7_75t_L g1062 ( 
.A1(n_909),
.A2(n_834),
.B1(n_833),
.B2(n_798),
.Y(n_1062)
);

NOR2x1_ASAP7_75t_L g1063 ( 
.A(n_926),
.B(n_811),
.Y(n_1063)
);

AOI22xp5_ASAP7_75t_L g1064 ( 
.A1(n_949),
.A2(n_895),
.B1(n_924),
.B2(n_956),
.Y(n_1064)
);

OA21x2_ASAP7_75t_L g1065 ( 
.A1(n_939),
.A2(n_831),
.B(n_832),
.Y(n_1065)
);

BUFx10_ASAP7_75t_L g1066 ( 
.A(n_860),
.Y(n_1066)
);

OR2x2_ASAP7_75t_L g1067 ( 
.A(n_945),
.B(n_811),
.Y(n_1067)
);

O2A1O1Ixp33_ASAP7_75t_L g1068 ( 
.A1(n_1006),
.A2(n_834),
.B(n_833),
.C(n_827),
.Y(n_1068)
);

CKINVDCx10_ASAP7_75t_R g1069 ( 
.A(n_854),
.Y(n_1069)
);

INVx1_ASAP7_75t_L g1070 ( 
.A(n_1006),
.Y(n_1070)
);

AND2x2_ASAP7_75t_L g1071 ( 
.A(n_874),
.B(n_335),
.Y(n_1071)
);

NOR2xp33_ASAP7_75t_SL g1072 ( 
.A(n_915),
.B(n_341),
.Y(n_1072)
);

OR2x6_ASAP7_75t_L g1073 ( 
.A(n_960),
.B(n_815),
.Y(n_1073)
);

BUFx6f_ASAP7_75t_L g1074 ( 
.A(n_989),
.Y(n_1074)
);

A2O1A1Ixp33_ASAP7_75t_L g1075 ( 
.A1(n_933),
.A2(n_682),
.B(n_815),
.C(n_827),
.Y(n_1075)
);

A2O1A1Ixp33_ASAP7_75t_SL g1076 ( 
.A1(n_967),
.A2(n_644),
.B(n_649),
.C(n_629),
.Y(n_1076)
);

AOI21xp5_ASAP7_75t_L g1077 ( 
.A1(n_918),
.A2(n_613),
.B(n_598),
.Y(n_1077)
);

AOI21xp5_ASAP7_75t_L g1078 ( 
.A1(n_918),
.A2(n_613),
.B(n_598),
.Y(n_1078)
);

O2A1O1Ixp33_ASAP7_75t_L g1079 ( 
.A1(n_923),
.A2(n_671),
.B(n_662),
.C(n_660),
.Y(n_1079)
);

O2A1O1Ixp33_ASAP7_75t_L g1080 ( 
.A1(n_933),
.A2(n_671),
.B(n_589),
.C(n_585),
.Y(n_1080)
);

OAI22xp5_ASAP7_75t_L g1081 ( 
.A1(n_909),
.A2(n_336),
.B1(n_342),
.B2(n_346),
.Y(n_1081)
);

AOI21xp5_ASAP7_75t_L g1082 ( 
.A1(n_918),
.A2(n_598),
.B(n_551),
.Y(n_1082)
);

INVx1_ASAP7_75t_SL g1083 ( 
.A(n_963),
.Y(n_1083)
);

NAND2xp5_ASAP7_75t_L g1084 ( 
.A(n_865),
.B(n_655),
.Y(n_1084)
);

NAND2xp5_ASAP7_75t_L g1085 ( 
.A(n_871),
.B(n_643),
.Y(n_1085)
);

AOI21xp5_ASAP7_75t_L g1086 ( 
.A1(n_937),
.A2(n_983),
.B(n_907),
.Y(n_1086)
);

NAND2xp5_ASAP7_75t_SL g1087 ( 
.A(n_915),
.B(n_344),
.Y(n_1087)
);

AOI21xp5_ASAP7_75t_L g1088 ( 
.A1(n_983),
.A2(n_851),
.B(n_994),
.Y(n_1088)
);

BUFx6f_ASAP7_75t_L g1089 ( 
.A(n_989),
.Y(n_1089)
);

OAI22xp5_ASAP7_75t_SL g1090 ( 
.A1(n_942),
.A2(n_342),
.B1(n_346),
.B2(n_347),
.Y(n_1090)
);

INVx1_ASAP7_75t_L g1091 ( 
.A(n_852),
.Y(n_1091)
);

INVxp67_ASAP7_75t_L g1092 ( 
.A(n_946),
.Y(n_1092)
);

NAND2xp5_ASAP7_75t_SL g1093 ( 
.A(n_850),
.B(n_344),
.Y(n_1093)
);

INVx2_ASAP7_75t_L g1094 ( 
.A(n_951),
.Y(n_1094)
);

INVx1_ASAP7_75t_L g1095 ( 
.A(n_853),
.Y(n_1095)
);

BUFx6f_ASAP7_75t_L g1096 ( 
.A(n_989),
.Y(n_1096)
);

AND2x2_ASAP7_75t_L g1097 ( 
.A(n_874),
.B(n_481),
.Y(n_1097)
);

NOR2xp67_ASAP7_75t_SL g1098 ( 
.A(n_989),
.B(n_222),
.Y(n_1098)
);

OAI22xp5_ASAP7_75t_L g1099 ( 
.A1(n_917),
.A2(n_521),
.B1(n_599),
.B2(n_606),
.Y(n_1099)
);

BUFx3_ASAP7_75t_L g1100 ( 
.A(n_870),
.Y(n_1100)
);

AOI22xp33_ASAP7_75t_L g1101 ( 
.A1(n_966),
.A2(n_288),
.B1(n_226),
.B2(n_227),
.Y(n_1101)
);

BUFx6f_ASAP7_75t_L g1102 ( 
.A(n_840),
.Y(n_1102)
);

A2O1A1Ixp33_ASAP7_75t_L g1103 ( 
.A1(n_999),
.A2(n_649),
.B(n_655),
.C(n_643),
.Y(n_1103)
);

INVx1_ASAP7_75t_L g1104 ( 
.A(n_864),
.Y(n_1104)
);

OR2x6_ASAP7_75t_SL g1105 ( 
.A(n_887),
.B(n_893),
.Y(n_1105)
);

NAND2xp5_ASAP7_75t_SL g1106 ( 
.A(n_996),
.B(n_225),
.Y(n_1106)
);

NOR2xp33_ASAP7_75t_L g1107 ( 
.A(n_920),
.B(n_643),
.Y(n_1107)
);

AOI21xp5_ASAP7_75t_L g1108 ( 
.A1(n_851),
.A2(n_598),
.B(n_645),
.Y(n_1108)
);

NAND2xp5_ASAP7_75t_L g1109 ( 
.A(n_866),
.B(n_655),
.Y(n_1109)
);

INVx4_ASAP7_75t_L g1110 ( 
.A(n_840),
.Y(n_1110)
);

INVx2_ASAP7_75t_SL g1111 ( 
.A(n_925),
.Y(n_1111)
);

AND2x2_ASAP7_75t_L g1112 ( 
.A(n_998),
.B(n_1008),
.Y(n_1112)
);

AOI21xp5_ASAP7_75t_L g1113 ( 
.A1(n_1001),
.A2(n_645),
.B(n_624),
.Y(n_1113)
);

AND2x2_ASAP7_75t_L g1114 ( 
.A(n_998),
.B(n_481),
.Y(n_1114)
);

AND2x2_ASAP7_75t_SL g1115 ( 
.A(n_917),
.B(n_481),
.Y(n_1115)
);

INVx4_ASAP7_75t_L g1116 ( 
.A(n_845),
.Y(n_1116)
);

O2A1O1Ixp33_ASAP7_75t_L g1117 ( 
.A1(n_879),
.A2(n_590),
.B(n_585),
.C(n_618),
.Y(n_1117)
);

OR2x6_ASAP7_75t_L g1118 ( 
.A(n_854),
.B(n_551),
.Y(n_1118)
);

CKINVDCx14_ASAP7_75t_R g1119 ( 
.A(n_854),
.Y(n_1119)
);

NOR2xp33_ASAP7_75t_L g1120 ( 
.A(n_955),
.B(n_643),
.Y(n_1120)
);

HB1xp67_ASAP7_75t_L g1121 ( 
.A(n_925),
.Y(n_1121)
);

BUFx3_ASAP7_75t_L g1122 ( 
.A(n_954),
.Y(n_1122)
);

AOI22x1_ASAP7_75t_L g1123 ( 
.A1(n_929),
.A2(n_962),
.B1(n_1005),
.B2(n_1002),
.Y(n_1123)
);

AOI21xp5_ASAP7_75t_L g1124 ( 
.A1(n_1003),
.A2(n_645),
.B(n_624),
.Y(n_1124)
);

NAND2xp5_ASAP7_75t_L g1125 ( 
.A(n_869),
.B(n_655),
.Y(n_1125)
);

AOI21xp5_ASAP7_75t_L g1126 ( 
.A1(n_1013),
.A2(n_645),
.B(n_624),
.Y(n_1126)
);

INVx5_ASAP7_75t_L g1127 ( 
.A(n_845),
.Y(n_1127)
);

BUFx3_ASAP7_75t_L g1128 ( 
.A(n_954),
.Y(n_1128)
);

NAND2xp5_ASAP7_75t_L g1129 ( 
.A(n_875),
.B(n_580),
.Y(n_1129)
);

AOI33xp33_ASAP7_75t_L g1130 ( 
.A1(n_1008),
.A2(n_1011),
.A3(n_1019),
.B1(n_1018),
.B2(n_1017),
.B3(n_1007),
.Y(n_1130)
);

INVx1_ASAP7_75t_L g1131 ( 
.A(n_881),
.Y(n_1131)
);

A2O1A1Ixp33_ASAP7_75t_L g1132 ( 
.A1(n_927),
.A2(n_580),
.B(n_589),
.C(n_618),
.Y(n_1132)
);

AOI22xp5_ASAP7_75t_L g1133 ( 
.A1(n_867),
.A2(n_927),
.B1(n_844),
.B2(n_878),
.Y(n_1133)
);

INVxp67_ASAP7_75t_L g1134 ( 
.A(n_877),
.Y(n_1134)
);

AOI21xp5_ASAP7_75t_L g1135 ( 
.A1(n_896),
.A2(n_645),
.B(n_624),
.Y(n_1135)
);

AOI21xp5_ASAP7_75t_L g1136 ( 
.A1(n_978),
.A2(n_624),
.B(n_613),
.Y(n_1136)
);

INVx4_ASAP7_75t_L g1137 ( 
.A(n_845),
.Y(n_1137)
);

NOR2xp33_ASAP7_75t_L g1138 ( 
.A(n_877),
.B(n_251),
.Y(n_1138)
);

NOR2x1_ASAP7_75t_L g1139 ( 
.A(n_926),
.B(n_590),
.Y(n_1139)
);

AOI21xp5_ASAP7_75t_L g1140 ( 
.A1(n_953),
.A2(n_613),
.B(n_461),
.Y(n_1140)
);

INVx2_ASAP7_75t_L g1141 ( 
.A(n_958),
.Y(n_1141)
);

AOI21xp5_ASAP7_75t_L g1142 ( 
.A1(n_953),
.A2(n_613),
.B(n_461),
.Y(n_1142)
);

INVx2_ASAP7_75t_SL g1143 ( 
.A(n_968),
.Y(n_1143)
);

NAND2xp5_ASAP7_75t_L g1144 ( 
.A(n_1011),
.B(n_592),
.Y(n_1144)
);

AOI21xp5_ASAP7_75t_L g1145 ( 
.A1(n_880),
.A2(n_899),
.B(n_891),
.Y(n_1145)
);

INVx2_ASAP7_75t_SL g1146 ( 
.A(n_968),
.Y(n_1146)
);

INVx5_ASAP7_75t_L g1147 ( 
.A(n_845),
.Y(n_1147)
);

INVx1_ASAP7_75t_L g1148 ( 
.A(n_901),
.Y(n_1148)
);

AOI21xp5_ASAP7_75t_L g1149 ( 
.A1(n_880),
.A2(n_899),
.B(n_891),
.Y(n_1149)
);

BUFx3_ASAP7_75t_L g1150 ( 
.A(n_969),
.Y(n_1150)
);

NAND2xp5_ASAP7_75t_L g1151 ( 
.A(n_1004),
.B(n_592),
.Y(n_1151)
);

NAND2xp5_ASAP7_75t_L g1152 ( 
.A(n_1004),
.B(n_599),
.Y(n_1152)
);

AO22x1_ASAP7_75t_L g1153 ( 
.A1(n_972),
.A2(n_252),
.B1(n_262),
.B2(n_264),
.Y(n_1153)
);

INVx2_ASAP7_75t_L g1154 ( 
.A(n_958),
.Y(n_1154)
);

O2A1O1Ixp5_ASAP7_75t_L g1155 ( 
.A1(n_1014),
.A2(n_521),
.B(n_606),
.C(n_475),
.Y(n_1155)
);

INVx2_ASAP7_75t_L g1156 ( 
.A(n_929),
.Y(n_1156)
);

AOI21xp5_ASAP7_75t_L g1157 ( 
.A1(n_903),
.A2(n_461),
.B(n_446),
.Y(n_1157)
);

NAND2xp5_ASAP7_75t_L g1158 ( 
.A(n_905),
.B(n_475),
.Y(n_1158)
);

NAND2xp5_ASAP7_75t_L g1159 ( 
.A(n_906),
.B(n_475),
.Y(n_1159)
);

AOI21xp5_ASAP7_75t_L g1160 ( 
.A1(n_903),
.A2(n_461),
.B(n_446),
.Y(n_1160)
);

NAND2xp5_ASAP7_75t_L g1161 ( 
.A(n_884),
.B(n_475),
.Y(n_1161)
);

INVx2_ASAP7_75t_L g1162 ( 
.A(n_962),
.Y(n_1162)
);

INVx2_ASAP7_75t_L g1163 ( 
.A(n_980),
.Y(n_1163)
);

BUFx2_ASAP7_75t_L g1164 ( 
.A(n_985),
.Y(n_1164)
);

INVx2_ASAP7_75t_L g1165 ( 
.A(n_990),
.Y(n_1165)
);

AOI21xp5_ASAP7_75t_L g1166 ( 
.A1(n_912),
.A2(n_461),
.B(n_268),
.Y(n_1166)
);

AO32x1_ASAP7_75t_L g1167 ( 
.A1(n_910),
.A2(n_2),
.A3(n_3),
.B1(n_4),
.B2(n_6),
.Y(n_1167)
);

INVx1_ASAP7_75t_L g1168 ( 
.A(n_928),
.Y(n_1168)
);

AOI21xp5_ASAP7_75t_L g1169 ( 
.A1(n_912),
.A2(n_932),
.B(n_913),
.Y(n_1169)
);

CKINVDCx5p33_ASAP7_75t_R g1170 ( 
.A(n_862),
.Y(n_1170)
);

BUFx4f_ASAP7_75t_SL g1171 ( 
.A(n_868),
.Y(n_1171)
);

INVx2_ASAP7_75t_SL g1172 ( 
.A(n_972),
.Y(n_1172)
);

OAI22xp5_ASAP7_75t_SL g1173 ( 
.A1(n_911),
.A2(n_271),
.B1(n_276),
.B2(n_278),
.Y(n_1173)
);

O2A1O1Ixp33_ASAP7_75t_SL g1174 ( 
.A1(n_843),
.A2(n_67),
.B(n_66),
.C(n_72),
.Y(n_1174)
);

OAI21xp5_ASAP7_75t_L g1175 ( 
.A1(n_1169),
.A2(n_950),
.B(n_914),
.Y(n_1175)
);

NAND4xp25_ASAP7_75t_SL g1176 ( 
.A(n_1101),
.B(n_997),
.C(n_921),
.D(n_889),
.Y(n_1176)
);

INVx3_ASAP7_75t_L g1177 ( 
.A(n_1110),
.Y(n_1177)
);

OAI21x1_ASAP7_75t_L g1178 ( 
.A1(n_1086),
.A2(n_940),
.B(n_1020),
.Y(n_1178)
);

NAND2xp5_ASAP7_75t_L g1179 ( 
.A(n_1023),
.B(n_961),
.Y(n_1179)
);

AOI221x1_ASAP7_75t_L g1180 ( 
.A1(n_1029),
.A2(n_979),
.B1(n_938),
.B2(n_952),
.C(n_964),
.Y(n_1180)
);

AOI21x1_ASAP7_75t_L g1181 ( 
.A1(n_1042),
.A2(n_1020),
.B(n_993),
.Y(n_1181)
);

OAI22xp5_ASAP7_75t_L g1182 ( 
.A1(n_1115),
.A2(n_843),
.B1(n_935),
.B2(n_868),
.Y(n_1182)
);

INVx1_ASAP7_75t_L g1183 ( 
.A(n_1091),
.Y(n_1183)
);

INVx1_ASAP7_75t_L g1184 ( 
.A(n_1095),
.Y(n_1184)
);

OAI21xp5_ASAP7_75t_L g1185 ( 
.A1(n_1075),
.A2(n_993),
.B(n_1000),
.Y(n_1185)
);

NAND2x1_ASAP7_75t_L g1186 ( 
.A(n_1110),
.B(n_868),
.Y(n_1186)
);

AO21x2_ASAP7_75t_L g1187 ( 
.A1(n_1076),
.A2(n_919),
.B(n_1000),
.Y(n_1187)
);

NOR2xp33_ASAP7_75t_L g1188 ( 
.A(n_1050),
.B(n_841),
.Y(n_1188)
);

AND2x2_ASAP7_75t_L g1189 ( 
.A(n_1112),
.B(n_842),
.Y(n_1189)
);

INVx2_ASAP7_75t_SL g1190 ( 
.A(n_1035),
.Y(n_1190)
);

OR2x6_ASAP7_75t_L g1191 ( 
.A(n_1043),
.B(n_868),
.Y(n_1191)
);

OA21x2_ASAP7_75t_L g1192 ( 
.A1(n_1155),
.A2(n_1016),
.B(n_1015),
.Y(n_1192)
);

OAI21x1_ASAP7_75t_L g1193 ( 
.A1(n_1123),
.A2(n_977),
.B(n_947),
.Y(n_1193)
);

A2O1A1Ixp33_ASAP7_75t_L g1194 ( 
.A1(n_1051),
.A2(n_959),
.B(n_976),
.C(n_941),
.Y(n_1194)
);

O2A1O1Ixp33_ASAP7_75t_L g1195 ( 
.A1(n_1053),
.A2(n_922),
.B(n_957),
.C(n_943),
.Y(n_1195)
);

INVx2_ASAP7_75t_L g1196 ( 
.A(n_1156),
.Y(n_1196)
);

AOI22xp33_ASAP7_75t_L g1197 ( 
.A1(n_1164),
.A2(n_922),
.B1(n_965),
.B2(n_849),
.Y(n_1197)
);

INVx1_ASAP7_75t_L g1198 ( 
.A(n_1104),
.Y(n_1198)
);

NAND2xp5_ASAP7_75t_L g1199 ( 
.A(n_1023),
.B(n_859),
.Y(n_1199)
);

AOI21xp5_ASAP7_75t_L g1200 ( 
.A1(n_1026),
.A2(n_986),
.B(n_971),
.Y(n_1200)
);

OR2x6_ASAP7_75t_L g1201 ( 
.A(n_1118),
.B(n_931),
.Y(n_1201)
);

INVx2_ASAP7_75t_L g1202 ( 
.A(n_1162),
.Y(n_1202)
);

OAI22xp5_ASAP7_75t_L g1203 ( 
.A1(n_1041),
.A2(n_975),
.B1(n_876),
.B2(n_847),
.Y(n_1203)
);

NAND2xp5_ASAP7_75t_L g1204 ( 
.A(n_1028),
.B(n_894),
.Y(n_1204)
);

NAND2xp5_ASAP7_75t_L g1205 ( 
.A(n_1031),
.B(n_902),
.Y(n_1205)
);

OAI21xp5_ASAP7_75t_L g1206 ( 
.A1(n_1103),
.A2(n_1012),
.B(n_1010),
.Y(n_1206)
);

INVx1_ASAP7_75t_L g1207 ( 
.A(n_1131),
.Y(n_1207)
);

AND2x4_ASAP7_75t_L g1208 ( 
.A(n_1150),
.B(n_847),
.Y(n_1208)
);

AOI21xp5_ASAP7_75t_L g1209 ( 
.A1(n_1088),
.A2(n_984),
.B(n_981),
.Y(n_1209)
);

AOI211x1_ASAP7_75t_L g1210 ( 
.A1(n_1034),
.A2(n_981),
.B(n_982),
.C(n_984),
.Y(n_1210)
);

AOI21x1_ASAP7_75t_L g1211 ( 
.A1(n_1054),
.A2(n_982),
.B(n_988),
.Y(n_1211)
);

A2O1A1Ixp33_ASAP7_75t_L g1212 ( 
.A1(n_1130),
.A2(n_1037),
.B(n_1032),
.C(n_1138),
.Y(n_1212)
);

NAND2xp5_ASAP7_75t_L g1213 ( 
.A(n_1114),
.B(n_904),
.Y(n_1213)
);

AOI21xp5_ASAP7_75t_L g1214 ( 
.A1(n_1027),
.A2(n_988),
.B(n_876),
.Y(n_1214)
);

OAI21x1_ASAP7_75t_SL g1215 ( 
.A1(n_1145),
.A2(n_1021),
.B(n_908),
.Y(n_1215)
);

AOI221xp5_ASAP7_75t_SL g1216 ( 
.A1(n_1081),
.A2(n_934),
.B1(n_930),
.B2(n_975),
.C(n_991),
.Y(n_1216)
);

HB1xp67_ASAP7_75t_L g1217 ( 
.A(n_1022),
.Y(n_1217)
);

NAND2x1p5_ASAP7_75t_L g1218 ( 
.A(n_1127),
.B(n_970),
.Y(n_1218)
);

AOI21x1_ASAP7_75t_SL g1219 ( 
.A1(n_1055),
.A2(n_1009),
.B(n_944),
.Y(n_1219)
);

NAND2xp5_ASAP7_75t_L g1220 ( 
.A(n_1097),
.B(n_944),
.Y(n_1220)
);

BUFx4f_ASAP7_75t_L g1221 ( 
.A(n_1073),
.Y(n_1221)
);

INVx2_ASAP7_75t_L g1222 ( 
.A(n_1067),
.Y(n_1222)
);

AOI21xp5_ASAP7_75t_SL g1223 ( 
.A1(n_1041),
.A2(n_461),
.B(n_279),
.Y(n_1223)
);

BUFx10_ASAP7_75t_L g1224 ( 
.A(n_1107),
.Y(n_1224)
);

INVx5_ASAP7_75t_L g1225 ( 
.A(n_1074),
.Y(n_1225)
);

NAND2xp5_ASAP7_75t_L g1226 ( 
.A(n_1024),
.B(n_284),
.Y(n_1226)
);

A2O1A1Ixp33_ASAP7_75t_L g1227 ( 
.A1(n_1120),
.A2(n_280),
.B(n_4),
.C(n_6),
.Y(n_1227)
);

AOI21x1_ASAP7_75t_L g1228 ( 
.A1(n_1047),
.A2(n_502),
.B(n_174),
.Y(n_1228)
);

NAND2xp5_ASAP7_75t_L g1229 ( 
.A(n_1030),
.B(n_2),
.Y(n_1229)
);

O2A1O1Ixp33_ASAP7_75t_L g1230 ( 
.A1(n_1134),
.A2(n_7),
.B(n_9),
.C(n_12),
.Y(n_1230)
);

AOI21xp5_ASAP7_75t_L g1231 ( 
.A1(n_1149),
.A2(n_1030),
.B(n_1135),
.Y(n_1231)
);

NAND2xp5_ASAP7_75t_L g1232 ( 
.A(n_1055),
.B(n_1148),
.Y(n_1232)
);

INVx1_ASAP7_75t_L g1233 ( 
.A(n_1168),
.Y(n_1233)
);

OAI21x1_ASAP7_75t_L g1234 ( 
.A1(n_1136),
.A2(n_131),
.B(n_172),
.Y(n_1234)
);

OAI21x1_ASAP7_75t_L g1235 ( 
.A1(n_1113),
.A2(n_1126),
.B(n_1124),
.Y(n_1235)
);

OR2x2_ASAP7_75t_L g1236 ( 
.A(n_1050),
.B(n_7),
.Y(n_1236)
);

OAI21xp5_ASAP7_75t_SL g1237 ( 
.A1(n_1052),
.A2(n_9),
.B(n_14),
.Y(n_1237)
);

BUFx3_ASAP7_75t_L g1238 ( 
.A(n_1100),
.Y(n_1238)
);

AOI21xp5_ASAP7_75t_L g1239 ( 
.A1(n_1039),
.A2(n_120),
.B(n_171),
.Y(n_1239)
);

AOI221x1_ASAP7_75t_L g1240 ( 
.A1(n_1132),
.A2(n_14),
.B1(n_15),
.B2(n_16),
.C(n_23),
.Y(n_1240)
);

AOI21xp5_ASAP7_75t_L g1241 ( 
.A1(n_1129),
.A2(n_1109),
.B(n_1084),
.Y(n_1241)
);

NAND3xp33_ASAP7_75t_L g1242 ( 
.A(n_1040),
.B(n_16),
.C(n_25),
.Y(n_1242)
);

NAND2xp5_ASAP7_75t_L g1243 ( 
.A(n_1129),
.B(n_26),
.Y(n_1243)
);

OAI21x1_ASAP7_75t_L g1244 ( 
.A1(n_1140),
.A2(n_76),
.B(n_164),
.Y(n_1244)
);

OAI21x1_ASAP7_75t_L g1245 ( 
.A1(n_1142),
.A2(n_115),
.B(n_149),
.Y(n_1245)
);

INVx3_ASAP7_75t_L g1246 ( 
.A(n_1116),
.Y(n_1246)
);

O2A1O1Ixp33_ASAP7_75t_L g1247 ( 
.A1(n_1092),
.A2(n_34),
.B(n_36),
.C(n_37),
.Y(n_1247)
);

OAI21x1_ASAP7_75t_L g1248 ( 
.A1(n_1157),
.A2(n_109),
.B(n_147),
.Y(n_1248)
);

NAND2xp5_ASAP7_75t_SL g1249 ( 
.A(n_1083),
.B(n_34),
.Y(n_1249)
);

OAI21x1_ASAP7_75t_L g1250 ( 
.A1(n_1160),
.A2(n_108),
.B(n_144),
.Y(n_1250)
);

BUFx2_ASAP7_75t_R g1251 ( 
.A(n_1105),
.Y(n_1251)
);

AOI21xp5_ASAP7_75t_L g1252 ( 
.A1(n_1084),
.A2(n_106),
.B(n_141),
.Y(n_1252)
);

AO21x1_ASAP7_75t_L g1253 ( 
.A1(n_1046),
.A2(n_37),
.B(n_38),
.Y(n_1253)
);

BUFx2_ASAP7_75t_L g1254 ( 
.A(n_1025),
.Y(n_1254)
);

AO31x2_ASAP7_75t_L g1255 ( 
.A1(n_1099),
.A2(n_502),
.A3(n_41),
.B(n_43),
.Y(n_1255)
);

OAI21x1_ASAP7_75t_L g1256 ( 
.A1(n_1108),
.A2(n_139),
.B(n_137),
.Y(n_1256)
);

AOI21xp5_ASAP7_75t_L g1257 ( 
.A1(n_1109),
.A2(n_89),
.B(n_86),
.Y(n_1257)
);

NAND3xp33_ASAP7_75t_L g1258 ( 
.A(n_1040),
.B(n_40),
.C(n_44),
.Y(n_1258)
);

NAND3x1_ASAP7_75t_L g1259 ( 
.A(n_1064),
.B(n_40),
.C(n_45),
.Y(n_1259)
);

BUFx6f_ASAP7_75t_L g1260 ( 
.A(n_1074),
.Y(n_1260)
);

NAND2xp5_ASAP7_75t_L g1261 ( 
.A(n_1036),
.B(n_47),
.Y(n_1261)
);

A2O1A1Ixp33_ASAP7_75t_L g1262 ( 
.A1(n_1058),
.A2(n_49),
.B(n_51),
.C(n_53),
.Y(n_1262)
);

INVx1_ASAP7_75t_L g1263 ( 
.A(n_1038),
.Y(n_1263)
);

INVx1_ASAP7_75t_L g1264 ( 
.A(n_1060),
.Y(n_1264)
);

AOI21xp5_ASAP7_75t_L g1265 ( 
.A1(n_1125),
.A2(n_84),
.B(n_502),
.Y(n_1265)
);

O2A1O1Ixp33_ASAP7_75t_SL g1266 ( 
.A1(n_1106),
.A2(n_49),
.B(n_53),
.C(n_54),
.Y(n_1266)
);

OAI21x1_ASAP7_75t_L g1267 ( 
.A1(n_1099),
.A2(n_502),
.B(n_54),
.Y(n_1267)
);

BUFx10_ASAP7_75t_L g1268 ( 
.A(n_1170),
.Y(n_1268)
);

OA21x2_ASAP7_75t_L g1269 ( 
.A1(n_1161),
.A2(n_502),
.B(n_56),
.Y(n_1269)
);

AOI21xp5_ASAP7_75t_L g1270 ( 
.A1(n_1125),
.A2(n_502),
.B(n_1161),
.Y(n_1270)
);

AOI21xp5_ASAP7_75t_L g1271 ( 
.A1(n_1046),
.A2(n_1056),
.B(n_1077),
.Y(n_1271)
);

O2A1O1Ixp5_ASAP7_75t_L g1272 ( 
.A1(n_1098),
.A2(n_1087),
.B(n_1093),
.C(n_1153),
.Y(n_1272)
);

O2A1O1Ixp33_ASAP7_75t_L g1273 ( 
.A1(n_1081),
.A2(n_1083),
.B(n_1048),
.C(n_1121),
.Y(n_1273)
);

CKINVDCx16_ASAP7_75t_R g1274 ( 
.A(n_1066),
.Y(n_1274)
);

HB1xp67_ASAP7_75t_L g1275 ( 
.A(n_1070),
.Y(n_1275)
);

INVx1_ASAP7_75t_L g1276 ( 
.A(n_1163),
.Y(n_1276)
);

OAI21x1_ASAP7_75t_L g1277 ( 
.A1(n_1158),
.A2(n_1159),
.B(n_1062),
.Y(n_1277)
);

OAI21x1_ASAP7_75t_L g1278 ( 
.A1(n_1158),
.A2(n_1159),
.B(n_1062),
.Y(n_1278)
);

INVx1_ASAP7_75t_L g1279 ( 
.A(n_1165),
.Y(n_1279)
);

AND2x4_ASAP7_75t_L g1280 ( 
.A(n_1073),
.B(n_1111),
.Y(n_1280)
);

OAI22xp5_ASAP7_75t_L g1281 ( 
.A1(n_1118),
.A2(n_1119),
.B1(n_1172),
.B2(n_1127),
.Y(n_1281)
);

AO31x2_ASAP7_75t_L g1282 ( 
.A1(n_1151),
.A2(n_1152),
.A3(n_1166),
.B(n_1085),
.Y(n_1282)
);

OAI21x1_ASAP7_75t_L g1283 ( 
.A1(n_1079),
.A2(n_1078),
.B(n_1082),
.Y(n_1283)
);

AOI21xp5_ASAP7_75t_L g1284 ( 
.A1(n_1127),
.A2(n_1147),
.B(n_1068),
.Y(n_1284)
);

NAND2xp5_ASAP7_75t_L g1285 ( 
.A(n_1071),
.B(n_1146),
.Y(n_1285)
);

NAND2xp5_ASAP7_75t_L g1286 ( 
.A(n_1151),
.B(n_1152),
.Y(n_1286)
);

AND2x4_ASAP7_75t_L g1287 ( 
.A(n_1073),
.B(n_1122),
.Y(n_1287)
);

OAI21x1_ASAP7_75t_L g1288 ( 
.A1(n_1080),
.A2(n_1117),
.B(n_1065),
.Y(n_1288)
);

OAI21x1_ASAP7_75t_L g1289 ( 
.A1(n_1065),
.A2(n_1139),
.B(n_1063),
.Y(n_1289)
);

NAND2xp5_ASAP7_75t_SL g1290 ( 
.A(n_1072),
.B(n_1128),
.Y(n_1290)
);

AND2x2_ASAP7_75t_L g1291 ( 
.A(n_1033),
.B(n_1044),
.Y(n_1291)
);

O2A1O1Ixp33_ASAP7_75t_SL g1292 ( 
.A1(n_1144),
.A2(n_1143),
.B(n_1049),
.C(n_1057),
.Y(n_1292)
);

INVx2_ASAP7_75t_L g1293 ( 
.A(n_1059),
.Y(n_1293)
);

AO31x2_ASAP7_75t_L g1294 ( 
.A1(n_1094),
.A2(n_1154),
.A3(n_1141),
.B(n_1116),
.Y(n_1294)
);

BUFx4f_ASAP7_75t_SL g1295 ( 
.A(n_1066),
.Y(n_1295)
);

O2A1O1Ixp5_ASAP7_75t_L g1296 ( 
.A1(n_1045),
.A2(n_1061),
.B(n_1137),
.C(n_1174),
.Y(n_1296)
);

NAND2xp5_ASAP7_75t_L g1297 ( 
.A(n_1045),
.B(n_1061),
.Y(n_1297)
);

INVx1_ASAP7_75t_L g1298 ( 
.A(n_1074),
.Y(n_1298)
);

AOI21xp5_ASAP7_75t_L g1299 ( 
.A1(n_1127),
.A2(n_1147),
.B(n_1072),
.Y(n_1299)
);

OAI21x1_ASAP7_75t_L g1300 ( 
.A1(n_1137),
.A2(n_1171),
.B(n_1102),
.Y(n_1300)
);

OR2x6_ASAP7_75t_L g1301 ( 
.A(n_1089),
.B(n_1096),
.Y(n_1301)
);

AOI21xp5_ASAP7_75t_L g1302 ( 
.A1(n_1089),
.A2(n_1096),
.B(n_1102),
.Y(n_1302)
);

BUFx4f_ASAP7_75t_SL g1303 ( 
.A(n_1102),
.Y(n_1303)
);

OAI21x1_ASAP7_75t_SL g1304 ( 
.A1(n_1167),
.A2(n_1069),
.B(n_1173),
.Y(n_1304)
);

INVxp67_ASAP7_75t_SL g1305 ( 
.A(n_1090),
.Y(n_1305)
);

AND2x4_ASAP7_75t_L g1306 ( 
.A(n_1112),
.B(n_1150),
.Y(n_1306)
);

A2O1A1Ixp33_ASAP7_75t_L g1307 ( 
.A1(n_1029),
.A2(n_743),
.B(n_839),
.C(n_897),
.Y(n_1307)
);

INVx1_ASAP7_75t_L g1308 ( 
.A(n_1091),
.Y(n_1308)
);

AOI221x1_ASAP7_75t_L g1309 ( 
.A1(n_1029),
.A2(n_689),
.B1(n_898),
.B2(n_839),
.C(n_685),
.Y(n_1309)
);

AOI21xp5_ASAP7_75t_L g1310 ( 
.A1(n_1026),
.A2(n_856),
.B(n_767),
.Y(n_1310)
);

OAI21x1_ASAP7_75t_L g1311 ( 
.A1(n_1086),
.A2(n_1123),
.B(n_1145),
.Y(n_1311)
);

A2O1A1Ixp33_ASAP7_75t_L g1312 ( 
.A1(n_1029),
.A2(n_743),
.B(n_839),
.C(n_897),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_1091),
.Y(n_1313)
);

OAI21xp5_ASAP7_75t_L g1314 ( 
.A1(n_1169),
.A2(n_1075),
.B(n_1103),
.Y(n_1314)
);

OAI21xp5_ASAP7_75t_L g1315 ( 
.A1(n_1169),
.A2(n_1075),
.B(n_1103),
.Y(n_1315)
);

AOI21xp5_ASAP7_75t_L g1316 ( 
.A1(n_1026),
.A2(n_856),
.B(n_767),
.Y(n_1316)
);

BUFx6f_ASAP7_75t_L g1317 ( 
.A(n_1074),
.Y(n_1317)
);

NAND2xp5_ASAP7_75t_L g1318 ( 
.A(n_1023),
.B(n_839),
.Y(n_1318)
);

AOI21x1_ASAP7_75t_L g1319 ( 
.A1(n_1042),
.A2(n_1086),
.B(n_1054),
.Y(n_1319)
);

AO31x2_ASAP7_75t_L g1320 ( 
.A1(n_1103),
.A2(n_1075),
.A3(n_1132),
.B(n_967),
.Y(n_1320)
);

AND2x2_ASAP7_75t_L g1321 ( 
.A(n_1112),
.B(n_1071),
.Y(n_1321)
);

OAI21x1_ASAP7_75t_L g1322 ( 
.A1(n_1086),
.A2(n_1123),
.B(n_1145),
.Y(n_1322)
);

CKINVDCx5p33_ASAP7_75t_R g1323 ( 
.A(n_1025),
.Y(n_1323)
);

INVx1_ASAP7_75t_L g1324 ( 
.A(n_1091),
.Y(n_1324)
);

OR2x6_ASAP7_75t_L g1325 ( 
.A(n_1043),
.B(n_1118),
.Y(n_1325)
);

OR2x2_ASAP7_75t_L g1326 ( 
.A(n_1050),
.B(n_886),
.Y(n_1326)
);

INVx2_ASAP7_75t_L g1327 ( 
.A(n_1156),
.Y(n_1327)
);

OAI22xp5_ASAP7_75t_L g1328 ( 
.A1(n_1115),
.A2(n_677),
.B1(n_839),
.B2(n_595),
.Y(n_1328)
);

AOI21xp5_ASAP7_75t_L g1329 ( 
.A1(n_1026),
.A2(n_856),
.B(n_767),
.Y(n_1329)
);

BUFx2_ASAP7_75t_L g1330 ( 
.A(n_1035),
.Y(n_1330)
);

HB1xp67_ASAP7_75t_L g1331 ( 
.A(n_1326),
.Y(n_1331)
);

INVx1_ASAP7_75t_SL g1332 ( 
.A(n_1254),
.Y(n_1332)
);

NAND2x1p5_ASAP7_75t_L g1333 ( 
.A(n_1225),
.B(n_1221),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_1183),
.Y(n_1334)
);

BUFx3_ASAP7_75t_L g1335 ( 
.A(n_1330),
.Y(n_1335)
);

BUFx2_ASAP7_75t_L g1336 ( 
.A(n_1323),
.Y(n_1336)
);

AOI21xp5_ASAP7_75t_L g1337 ( 
.A1(n_1329),
.A2(n_1175),
.B(n_1231),
.Y(n_1337)
);

INVx4_ASAP7_75t_L g1338 ( 
.A(n_1225),
.Y(n_1338)
);

OAI21x1_ASAP7_75t_L g1339 ( 
.A1(n_1311),
.A2(n_1322),
.B(n_1219),
.Y(n_1339)
);

BUFx12f_ASAP7_75t_L g1340 ( 
.A(n_1224),
.Y(n_1340)
);

OAI21x1_ASAP7_75t_L g1341 ( 
.A1(n_1319),
.A2(n_1235),
.B(n_1283),
.Y(n_1341)
);

INVx3_ASAP7_75t_L g1342 ( 
.A(n_1201),
.Y(n_1342)
);

CKINVDCx6p67_ASAP7_75t_R g1343 ( 
.A(n_1238),
.Y(n_1343)
);

INVx4_ASAP7_75t_SL g1344 ( 
.A(n_1255),
.Y(n_1344)
);

INVx1_ASAP7_75t_L g1345 ( 
.A(n_1184),
.Y(n_1345)
);

INVx1_ASAP7_75t_L g1346 ( 
.A(n_1198),
.Y(n_1346)
);

A2O1A1Ixp33_ASAP7_75t_L g1347 ( 
.A1(n_1312),
.A2(n_1328),
.B(n_1212),
.C(n_1258),
.Y(n_1347)
);

OAI21x1_ASAP7_75t_L g1348 ( 
.A1(n_1228),
.A2(n_1178),
.B(n_1193),
.Y(n_1348)
);

OAI21x1_ASAP7_75t_L g1349 ( 
.A1(n_1214),
.A2(n_1288),
.B(n_1209),
.Y(n_1349)
);

A2O1A1Ixp33_ASAP7_75t_L g1350 ( 
.A1(n_1328),
.A2(n_1242),
.B(n_1258),
.C(n_1237),
.Y(n_1350)
);

AOI222xp33_ASAP7_75t_L g1351 ( 
.A1(n_1237),
.A2(n_1305),
.B1(n_1242),
.B2(n_1249),
.C1(n_1321),
.C2(n_1291),
.Y(n_1351)
);

INVx2_ASAP7_75t_SL g1352 ( 
.A(n_1190),
.Y(n_1352)
);

AND2x4_ASAP7_75t_L g1353 ( 
.A(n_1201),
.B(n_1208),
.Y(n_1353)
);

OAI221xp5_ASAP7_75t_L g1354 ( 
.A1(n_1227),
.A2(n_1262),
.B1(n_1285),
.B2(n_1247),
.C(n_1230),
.Y(n_1354)
);

NAND2xp5_ASAP7_75t_L g1355 ( 
.A(n_1222),
.B(n_1189),
.Y(n_1355)
);

INVx1_ASAP7_75t_L g1356 ( 
.A(n_1207),
.Y(n_1356)
);

OAI21x1_ASAP7_75t_L g1357 ( 
.A1(n_1270),
.A2(n_1315),
.B(n_1314),
.Y(n_1357)
);

NAND2x1p5_ASAP7_75t_L g1358 ( 
.A(n_1225),
.B(n_1221),
.Y(n_1358)
);

NAND2xp5_ASAP7_75t_L g1359 ( 
.A(n_1205),
.B(n_1179),
.Y(n_1359)
);

OAI21x1_ASAP7_75t_L g1360 ( 
.A1(n_1315),
.A2(n_1211),
.B(n_1234),
.Y(n_1360)
);

AND2x2_ASAP7_75t_L g1361 ( 
.A(n_1306),
.B(n_1188),
.Y(n_1361)
);

INVx1_ASAP7_75t_L g1362 ( 
.A(n_1308),
.Y(n_1362)
);

NAND2x1p5_ASAP7_75t_L g1363 ( 
.A(n_1299),
.B(n_1177),
.Y(n_1363)
);

HB1xp67_ASAP7_75t_L g1364 ( 
.A(n_1217),
.Y(n_1364)
);

A2O1A1Ixp33_ASAP7_75t_L g1365 ( 
.A1(n_1175),
.A2(n_1267),
.B(n_1273),
.C(n_1206),
.Y(n_1365)
);

INVx1_ASAP7_75t_L g1366 ( 
.A(n_1313),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_1324),
.Y(n_1367)
);

NAND2x1_ASAP7_75t_L g1368 ( 
.A(n_1215),
.B(n_1191),
.Y(n_1368)
);

AOI22xp33_ASAP7_75t_L g1369 ( 
.A1(n_1253),
.A2(n_1176),
.B1(n_1304),
.B2(n_1229),
.Y(n_1369)
);

NAND2x1p5_ASAP7_75t_L g1370 ( 
.A(n_1177),
.B(n_1246),
.Y(n_1370)
);

OAI21x1_ASAP7_75t_L g1371 ( 
.A1(n_1289),
.A2(n_1278),
.B(n_1277),
.Y(n_1371)
);

AOI22xp33_ASAP7_75t_L g1372 ( 
.A1(n_1229),
.A2(n_1243),
.B1(n_1236),
.B2(n_1261),
.Y(n_1372)
);

INVx1_ASAP7_75t_L g1373 ( 
.A(n_1233),
.Y(n_1373)
);

NAND2xp5_ASAP7_75t_L g1374 ( 
.A(n_1232),
.B(n_1213),
.Y(n_1374)
);

OAI21x1_ASAP7_75t_L g1375 ( 
.A1(n_1248),
.A2(n_1250),
.B(n_1256),
.Y(n_1375)
);

BUFx2_ASAP7_75t_L g1376 ( 
.A(n_1306),
.Y(n_1376)
);

OAI21x1_ASAP7_75t_L g1377 ( 
.A1(n_1181),
.A2(n_1245),
.B(n_1244),
.Y(n_1377)
);

INVx3_ASAP7_75t_L g1378 ( 
.A(n_1201),
.Y(n_1378)
);

OAI21x1_ASAP7_75t_L g1379 ( 
.A1(n_1241),
.A2(n_1185),
.B(n_1200),
.Y(n_1379)
);

INVx2_ASAP7_75t_L g1380 ( 
.A(n_1202),
.Y(n_1380)
);

NOR2x1_ASAP7_75t_SL g1381 ( 
.A(n_1191),
.B(n_1325),
.Y(n_1381)
);

AOI21xp5_ASAP7_75t_L g1382 ( 
.A1(n_1206),
.A2(n_1223),
.B(n_1204),
.Y(n_1382)
);

INVx2_ASAP7_75t_L g1383 ( 
.A(n_1327),
.Y(n_1383)
);

OAI22xp5_ASAP7_75t_L g1384 ( 
.A1(n_1197),
.A2(n_1232),
.B1(n_1325),
.B2(n_1226),
.Y(n_1384)
);

NAND2x1p5_ASAP7_75t_L g1385 ( 
.A(n_1246),
.B(n_1186),
.Y(n_1385)
);

OAI21x1_ASAP7_75t_L g1386 ( 
.A1(n_1296),
.A2(n_1195),
.B(n_1284),
.Y(n_1386)
);

BUFx6f_ASAP7_75t_L g1387 ( 
.A(n_1260),
.Y(n_1387)
);

INVx1_ASAP7_75t_L g1388 ( 
.A(n_1263),
.Y(n_1388)
);

INVx2_ASAP7_75t_L g1389 ( 
.A(n_1276),
.Y(n_1389)
);

OAI21xp5_ASAP7_75t_L g1390 ( 
.A1(n_1309),
.A2(n_1272),
.B(n_1194),
.Y(n_1390)
);

INVx1_ASAP7_75t_L g1391 ( 
.A(n_1264),
.Y(n_1391)
);

OAI21x1_ASAP7_75t_L g1392 ( 
.A1(n_1239),
.A2(n_1192),
.B(n_1203),
.Y(n_1392)
);

NAND2x1p5_ASAP7_75t_L g1393 ( 
.A(n_1300),
.B(n_1287),
.Y(n_1393)
);

NAND2xp5_ASAP7_75t_L g1394 ( 
.A(n_1199),
.B(n_1243),
.Y(n_1394)
);

NAND2x1p5_ASAP7_75t_L g1395 ( 
.A(n_1287),
.B(n_1290),
.Y(n_1395)
);

NOR2xp33_ASAP7_75t_L g1396 ( 
.A(n_1275),
.B(n_1220),
.Y(n_1396)
);

BUFx2_ASAP7_75t_L g1397 ( 
.A(n_1303),
.Y(n_1397)
);

AOI21xp5_ASAP7_75t_L g1398 ( 
.A1(n_1204),
.A2(n_1182),
.B(n_1286),
.Y(n_1398)
);

AOI21xp5_ASAP7_75t_L g1399 ( 
.A1(n_1182),
.A2(n_1286),
.B(n_1203),
.Y(n_1399)
);

INVx2_ASAP7_75t_L g1400 ( 
.A(n_1279),
.Y(n_1400)
);

NAND2x1p5_ASAP7_75t_L g1401 ( 
.A(n_1280),
.B(n_1208),
.Y(n_1401)
);

INVx2_ASAP7_75t_SL g1402 ( 
.A(n_1224),
.Y(n_1402)
);

OAI21x1_ASAP7_75t_L g1403 ( 
.A1(n_1192),
.A2(n_1265),
.B(n_1257),
.Y(n_1403)
);

INVx1_ASAP7_75t_L g1404 ( 
.A(n_1293),
.Y(n_1404)
);

INVx1_ASAP7_75t_L g1405 ( 
.A(n_1294),
.Y(n_1405)
);

INVx2_ASAP7_75t_SL g1406 ( 
.A(n_1280),
.Y(n_1406)
);

AO21x2_ASAP7_75t_L g1407 ( 
.A1(n_1187),
.A2(n_1292),
.B(n_1252),
.Y(n_1407)
);

INVx2_ASAP7_75t_L g1408 ( 
.A(n_1294),
.Y(n_1408)
);

AOI22xp33_ASAP7_75t_L g1409 ( 
.A1(n_1325),
.A2(n_1259),
.B1(n_1281),
.B2(n_1268),
.Y(n_1409)
);

O2A1O1Ixp33_ASAP7_75t_L g1410 ( 
.A1(n_1266),
.A2(n_1281),
.B(n_1297),
.C(n_1191),
.Y(n_1410)
);

AOI22xp33_ASAP7_75t_L g1411 ( 
.A1(n_1268),
.A2(n_1187),
.B1(n_1269),
.B2(n_1240),
.Y(n_1411)
);

CKINVDCx11_ASAP7_75t_R g1412 ( 
.A(n_1274),
.Y(n_1412)
);

OAI21x1_ASAP7_75t_L g1413 ( 
.A1(n_1269),
.A2(n_1218),
.B(n_1302),
.Y(n_1413)
);

NOR2xp33_ASAP7_75t_L g1414 ( 
.A(n_1297),
.B(n_1298),
.Y(n_1414)
);

INVx1_ASAP7_75t_L g1415 ( 
.A(n_1294),
.Y(n_1415)
);

INVx2_ASAP7_75t_L g1416 ( 
.A(n_1320),
.Y(n_1416)
);

OAI21x1_ASAP7_75t_L g1417 ( 
.A1(n_1218),
.A2(n_1320),
.B(n_1210),
.Y(n_1417)
);

INVx3_ASAP7_75t_L g1418 ( 
.A(n_1260),
.Y(n_1418)
);

INVx2_ASAP7_75t_SL g1419 ( 
.A(n_1260),
.Y(n_1419)
);

NOR2xp67_ASAP7_75t_L g1420 ( 
.A(n_1317),
.B(n_1251),
.Y(n_1420)
);

AOI22xp33_ASAP7_75t_L g1421 ( 
.A1(n_1295),
.A2(n_1317),
.B1(n_1301),
.B2(n_1216),
.Y(n_1421)
);

AOI22xp33_ASAP7_75t_L g1422 ( 
.A1(n_1317),
.A2(n_1301),
.B1(n_1216),
.B2(n_1320),
.Y(n_1422)
);

OR2x2_ASAP7_75t_L g1423 ( 
.A(n_1282),
.B(n_1222),
.Y(n_1423)
);

OAI21x1_ASAP7_75t_L g1424 ( 
.A1(n_1282),
.A2(n_1322),
.B(n_1311),
.Y(n_1424)
);

OAI21x1_ASAP7_75t_L g1425 ( 
.A1(n_1282),
.A2(n_1322),
.B(n_1311),
.Y(n_1425)
);

INVx2_ASAP7_75t_SL g1426 ( 
.A(n_1238),
.Y(n_1426)
);

INVx1_ASAP7_75t_L g1427 ( 
.A(n_1183),
.Y(n_1427)
);

OAI22xp5_ASAP7_75t_L g1428 ( 
.A1(n_1307),
.A2(n_1312),
.B1(n_839),
.B2(n_1318),
.Y(n_1428)
);

AND2x2_ASAP7_75t_L g1429 ( 
.A(n_1321),
.B(n_1112),
.Y(n_1429)
);

BUFx8_ASAP7_75t_L g1430 ( 
.A(n_1330),
.Y(n_1430)
);

AO21x2_ASAP7_75t_L g1431 ( 
.A1(n_1271),
.A2(n_1175),
.B(n_1314),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_1183),
.Y(n_1432)
);

INVx2_ASAP7_75t_L g1433 ( 
.A(n_1196),
.Y(n_1433)
);

AOI22xp33_ASAP7_75t_L g1434 ( 
.A1(n_1253),
.A2(n_898),
.B1(n_839),
.B2(n_1242),
.Y(n_1434)
);

INVx4_ASAP7_75t_SL g1435 ( 
.A(n_1255),
.Y(n_1435)
);

INVx1_ASAP7_75t_L g1436 ( 
.A(n_1183),
.Y(n_1436)
);

NAND2xp5_ASAP7_75t_SL g1437 ( 
.A(n_1307),
.B(n_1312),
.Y(n_1437)
);

A2O1A1Ixp33_ASAP7_75t_L g1438 ( 
.A1(n_1307),
.A2(n_1312),
.B(n_839),
.C(n_1328),
.Y(n_1438)
);

AOI22xp33_ASAP7_75t_L g1439 ( 
.A1(n_1253),
.A2(n_898),
.B1(n_839),
.B2(n_1242),
.Y(n_1439)
);

INVx2_ASAP7_75t_SL g1440 ( 
.A(n_1238),
.Y(n_1440)
);

INVx1_ASAP7_75t_L g1441 ( 
.A(n_1183),
.Y(n_1441)
);

AOI22xp33_ASAP7_75t_L g1442 ( 
.A1(n_1253),
.A2(n_898),
.B1(n_839),
.B2(n_1242),
.Y(n_1442)
);

BUFx2_ASAP7_75t_L g1443 ( 
.A(n_1330),
.Y(n_1443)
);

AO21x2_ASAP7_75t_L g1444 ( 
.A1(n_1271),
.A2(n_1175),
.B(n_1314),
.Y(n_1444)
);

OAI21x1_ASAP7_75t_L g1445 ( 
.A1(n_1311),
.A2(n_1322),
.B(n_1219),
.Y(n_1445)
);

AND2x2_ASAP7_75t_L g1446 ( 
.A(n_1321),
.B(n_1112),
.Y(n_1446)
);

AND2x2_ASAP7_75t_L g1447 ( 
.A(n_1321),
.B(n_1112),
.Y(n_1447)
);

INVx2_ASAP7_75t_L g1448 ( 
.A(n_1196),
.Y(n_1448)
);

INVx2_ASAP7_75t_L g1449 ( 
.A(n_1196),
.Y(n_1449)
);

OAI22xp33_ASAP7_75t_L g1450 ( 
.A1(n_1242),
.A2(n_839),
.B1(n_1258),
.B2(n_1309),
.Y(n_1450)
);

AO31x2_ASAP7_75t_L g1451 ( 
.A1(n_1309),
.A2(n_1180),
.A3(n_1271),
.B(n_1240),
.Y(n_1451)
);

OAI21xp5_ASAP7_75t_L g1452 ( 
.A1(n_1307),
.A2(n_1312),
.B(n_897),
.Y(n_1452)
);

OAI21x1_ASAP7_75t_L g1453 ( 
.A1(n_1311),
.A2(n_1322),
.B(n_1219),
.Y(n_1453)
);

AOI22xp33_ASAP7_75t_L g1454 ( 
.A1(n_1253),
.A2(n_898),
.B1(n_839),
.B2(n_1242),
.Y(n_1454)
);

AND2x2_ASAP7_75t_L g1455 ( 
.A(n_1321),
.B(n_1112),
.Y(n_1455)
);

INVxp67_ASAP7_75t_L g1456 ( 
.A(n_1326),
.Y(n_1456)
);

OR2x2_ASAP7_75t_L g1457 ( 
.A(n_1222),
.B(n_1326),
.Y(n_1457)
);

INVx1_ASAP7_75t_L g1458 ( 
.A(n_1183),
.Y(n_1458)
);

CKINVDCx16_ASAP7_75t_R g1459 ( 
.A(n_1274),
.Y(n_1459)
);

INVx1_ASAP7_75t_L g1460 ( 
.A(n_1183),
.Y(n_1460)
);

BUFx3_ASAP7_75t_L g1461 ( 
.A(n_1330),
.Y(n_1461)
);

AOI22xp33_ASAP7_75t_L g1462 ( 
.A1(n_1253),
.A2(n_898),
.B1(n_839),
.B2(n_1242),
.Y(n_1462)
);

OAI21x1_ASAP7_75t_L g1463 ( 
.A1(n_1311),
.A2(n_1322),
.B(n_1219),
.Y(n_1463)
);

AND2x4_ASAP7_75t_L g1464 ( 
.A(n_1201),
.B(n_1208),
.Y(n_1464)
);

OAI21x1_ASAP7_75t_L g1465 ( 
.A1(n_1311),
.A2(n_1322),
.B(n_1219),
.Y(n_1465)
);

INVx1_ASAP7_75t_L g1466 ( 
.A(n_1183),
.Y(n_1466)
);

NAND2xp5_ASAP7_75t_L g1467 ( 
.A(n_1318),
.B(n_1307),
.Y(n_1467)
);

BUFx3_ASAP7_75t_L g1468 ( 
.A(n_1330),
.Y(n_1468)
);

CKINVDCx20_ASAP7_75t_R g1469 ( 
.A(n_1295),
.Y(n_1469)
);

OR2x6_ASAP7_75t_L g1470 ( 
.A(n_1299),
.B(n_1325),
.Y(n_1470)
);

A2O1A1Ixp33_ASAP7_75t_L g1471 ( 
.A1(n_1452),
.A2(n_1347),
.B(n_1350),
.C(n_1454),
.Y(n_1471)
);

A2O1A1Ixp33_ASAP7_75t_L g1472 ( 
.A1(n_1347),
.A2(n_1350),
.B(n_1434),
.C(n_1439),
.Y(n_1472)
);

AOI21xp5_ASAP7_75t_SL g1473 ( 
.A1(n_1428),
.A2(n_1438),
.B(n_1467),
.Y(n_1473)
);

O2A1O1Ixp33_ASAP7_75t_L g1474 ( 
.A1(n_1450),
.A2(n_1437),
.B(n_1438),
.C(n_1354),
.Y(n_1474)
);

AND2x2_ASAP7_75t_L g1475 ( 
.A(n_1429),
.B(n_1446),
.Y(n_1475)
);

AND2x2_ASAP7_75t_L g1476 ( 
.A(n_1447),
.B(n_1455),
.Y(n_1476)
);

AND2x2_ASAP7_75t_L g1477 ( 
.A(n_1361),
.B(n_1396),
.Y(n_1477)
);

NAND2xp5_ASAP7_75t_L g1478 ( 
.A(n_1394),
.B(n_1398),
.Y(n_1478)
);

AND2x4_ASAP7_75t_L g1479 ( 
.A(n_1342),
.B(n_1378),
.Y(n_1479)
);

OAI22xp5_ASAP7_75t_L g1480 ( 
.A1(n_1434),
.A2(n_1439),
.B1(n_1442),
.B2(n_1462),
.Y(n_1480)
);

OAI22xp5_ASAP7_75t_L g1481 ( 
.A1(n_1442),
.A2(n_1454),
.B1(n_1462),
.B2(n_1409),
.Y(n_1481)
);

NAND2xp5_ASAP7_75t_L g1482 ( 
.A(n_1374),
.B(n_1359),
.Y(n_1482)
);

AND2x2_ASAP7_75t_L g1483 ( 
.A(n_1396),
.B(n_1376),
.Y(n_1483)
);

HB1xp67_ASAP7_75t_L g1484 ( 
.A(n_1331),
.Y(n_1484)
);

AND2x2_ASAP7_75t_L g1485 ( 
.A(n_1457),
.B(n_1355),
.Y(n_1485)
);

OAI22xp5_ASAP7_75t_L g1486 ( 
.A1(n_1409),
.A2(n_1372),
.B1(n_1369),
.B2(n_1395),
.Y(n_1486)
);

OR2x6_ASAP7_75t_L g1487 ( 
.A(n_1470),
.B(n_1368),
.Y(n_1487)
);

INVx2_ASAP7_75t_SL g1488 ( 
.A(n_1430),
.Y(n_1488)
);

OA21x2_ASAP7_75t_L g1489 ( 
.A1(n_1386),
.A2(n_1425),
.B(n_1424),
.Y(n_1489)
);

HB1xp67_ASAP7_75t_L g1490 ( 
.A(n_1364),
.Y(n_1490)
);

INVx1_ASAP7_75t_L g1491 ( 
.A(n_1334),
.Y(n_1491)
);

OAI22xp5_ASAP7_75t_L g1492 ( 
.A1(n_1372),
.A2(n_1369),
.B1(n_1395),
.B2(n_1332),
.Y(n_1492)
);

AND2x2_ASAP7_75t_L g1493 ( 
.A(n_1456),
.B(n_1406),
.Y(n_1493)
);

NAND2xp5_ASAP7_75t_L g1494 ( 
.A(n_1399),
.B(n_1450),
.Y(n_1494)
);

INVx2_ASAP7_75t_L g1495 ( 
.A(n_1380),
.Y(n_1495)
);

OA21x2_ASAP7_75t_L g1496 ( 
.A1(n_1386),
.A2(n_1425),
.B(n_1424),
.Y(n_1496)
);

O2A1O1Ixp33_ASAP7_75t_L g1497 ( 
.A1(n_1437),
.A2(n_1390),
.B(n_1365),
.C(n_1384),
.Y(n_1497)
);

NAND2xp5_ASAP7_75t_L g1498 ( 
.A(n_1382),
.B(n_1423),
.Y(n_1498)
);

A2O1A1Ixp33_ASAP7_75t_L g1499 ( 
.A1(n_1410),
.A2(n_1411),
.B(n_1357),
.C(n_1379),
.Y(n_1499)
);

INVx3_ASAP7_75t_L g1500 ( 
.A(n_1353),
.Y(n_1500)
);

NAND2xp5_ASAP7_75t_L g1501 ( 
.A(n_1414),
.B(n_1431),
.Y(n_1501)
);

NAND2xp5_ASAP7_75t_L g1502 ( 
.A(n_1414),
.B(n_1444),
.Y(n_1502)
);

AND2x4_ASAP7_75t_L g1503 ( 
.A(n_1342),
.B(n_1378),
.Y(n_1503)
);

BUFx4f_ASAP7_75t_SL g1504 ( 
.A(n_1469),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_1345),
.Y(n_1505)
);

HB1xp67_ASAP7_75t_L g1506 ( 
.A(n_1388),
.Y(n_1506)
);

OA21x2_ASAP7_75t_L g1507 ( 
.A1(n_1392),
.A2(n_1360),
.B(n_1371),
.Y(n_1507)
);

NAND2xp5_ASAP7_75t_L g1508 ( 
.A(n_1451),
.B(n_1346),
.Y(n_1508)
);

OA21x2_ASAP7_75t_L g1509 ( 
.A1(n_1392),
.A2(n_1360),
.B(n_1371),
.Y(n_1509)
);

AND2x2_ASAP7_75t_L g1510 ( 
.A(n_1464),
.B(n_1401),
.Y(n_1510)
);

OAI22xp5_ASAP7_75t_L g1511 ( 
.A1(n_1421),
.A2(n_1420),
.B1(n_1443),
.B2(n_1468),
.Y(n_1511)
);

AND2x4_ASAP7_75t_L g1512 ( 
.A(n_1381),
.B(n_1470),
.Y(n_1512)
);

OR2x2_ASAP7_75t_L g1513 ( 
.A(n_1389),
.B(n_1400),
.Y(n_1513)
);

AND2x4_ASAP7_75t_L g1514 ( 
.A(n_1470),
.B(n_1335),
.Y(n_1514)
);

O2A1O1Ixp33_ASAP7_75t_L g1515 ( 
.A1(n_1351),
.A2(n_1402),
.B(n_1352),
.C(n_1391),
.Y(n_1515)
);

A2O1A1Ixp33_ASAP7_75t_L g1516 ( 
.A1(n_1411),
.A2(n_1421),
.B(n_1403),
.C(n_1460),
.Y(n_1516)
);

OAI22xp5_ASAP7_75t_L g1517 ( 
.A1(n_1461),
.A2(n_1468),
.B1(n_1333),
.B2(n_1358),
.Y(n_1517)
);

AND2x2_ASAP7_75t_L g1518 ( 
.A(n_1401),
.B(n_1383),
.Y(n_1518)
);

OR2x2_ASAP7_75t_L g1519 ( 
.A(n_1389),
.B(n_1400),
.Y(n_1519)
);

NAND2xp5_ASAP7_75t_L g1520 ( 
.A(n_1451),
.B(n_1356),
.Y(n_1520)
);

OAI22xp5_ASAP7_75t_L g1521 ( 
.A1(n_1333),
.A2(n_1358),
.B1(n_1393),
.B2(n_1336),
.Y(n_1521)
);

AOI21xp5_ASAP7_75t_L g1522 ( 
.A1(n_1349),
.A2(n_1341),
.B(n_1403),
.Y(n_1522)
);

AOI21xp5_ASAP7_75t_L g1523 ( 
.A1(n_1407),
.A2(n_1375),
.B(n_1363),
.Y(n_1523)
);

OAI22xp5_ASAP7_75t_L g1524 ( 
.A1(n_1393),
.A2(n_1422),
.B1(n_1466),
.B2(n_1441),
.Y(n_1524)
);

OAI22xp5_ASAP7_75t_L g1525 ( 
.A1(n_1422),
.A2(n_1366),
.B1(n_1436),
.B2(n_1373),
.Y(n_1525)
);

NAND2xp5_ASAP7_75t_L g1526 ( 
.A(n_1451),
.B(n_1458),
.Y(n_1526)
);

AOI21xp5_ASAP7_75t_L g1527 ( 
.A1(n_1348),
.A2(n_1453),
.B(n_1339),
.Y(n_1527)
);

O2A1O1Ixp5_ASAP7_75t_L g1528 ( 
.A1(n_1416),
.A2(n_1405),
.B(n_1415),
.C(n_1408),
.Y(n_1528)
);

OR2x2_ASAP7_75t_L g1529 ( 
.A(n_1362),
.B(n_1427),
.Y(n_1529)
);

AOI21xp5_ASAP7_75t_L g1530 ( 
.A1(n_1348),
.A2(n_1445),
.B(n_1465),
.Y(n_1530)
);

BUFx6f_ASAP7_75t_L g1531 ( 
.A(n_1387),
.Y(n_1531)
);

OR2x2_ASAP7_75t_L g1532 ( 
.A(n_1367),
.B(n_1432),
.Y(n_1532)
);

OAI22x1_ASAP7_75t_L g1533 ( 
.A1(n_1370),
.A2(n_1404),
.B1(n_1440),
.B2(n_1426),
.Y(n_1533)
);

BUFx2_ASAP7_75t_L g1534 ( 
.A(n_1430),
.Y(n_1534)
);

O2A1O1Ixp33_ASAP7_75t_L g1535 ( 
.A1(n_1433),
.A2(n_1449),
.B(n_1448),
.C(n_1397),
.Y(n_1535)
);

A2O1A1Ixp33_ASAP7_75t_L g1536 ( 
.A1(n_1417),
.A2(n_1413),
.B(n_1377),
.C(n_1463),
.Y(n_1536)
);

AOI221x1_ASAP7_75t_SL g1537 ( 
.A1(n_1433),
.A2(n_1449),
.B1(n_1448),
.B2(n_1412),
.C(n_1459),
.Y(n_1537)
);

AND2x2_ASAP7_75t_L g1538 ( 
.A(n_1418),
.B(n_1387),
.Y(n_1538)
);

AOI21xp5_ASAP7_75t_SL g1539 ( 
.A1(n_1338),
.A2(n_1370),
.B(n_1385),
.Y(n_1539)
);

NOR2xp67_ASAP7_75t_L g1540 ( 
.A(n_1340),
.B(n_1419),
.Y(n_1540)
);

O2A1O1Ixp33_ASAP7_75t_L g1541 ( 
.A1(n_1385),
.A2(n_1469),
.B(n_1344),
.C(n_1435),
.Y(n_1541)
);

AND2x2_ASAP7_75t_L g1542 ( 
.A(n_1387),
.B(n_1343),
.Y(n_1542)
);

OAI22xp5_ASAP7_75t_L g1543 ( 
.A1(n_1340),
.A2(n_1338),
.B1(n_1387),
.B2(n_1430),
.Y(n_1543)
);

OAI22xp5_ASAP7_75t_L g1544 ( 
.A1(n_1338),
.A2(n_1344),
.B1(n_1435),
.B2(n_1413),
.Y(n_1544)
);

INVxp67_ASAP7_75t_L g1545 ( 
.A(n_1364),
.Y(n_1545)
);

OR2x2_ASAP7_75t_L g1546 ( 
.A(n_1331),
.B(n_1457),
.Y(n_1546)
);

AND2x2_ASAP7_75t_L g1547 ( 
.A(n_1429),
.B(n_1446),
.Y(n_1547)
);

AND2x2_ASAP7_75t_L g1548 ( 
.A(n_1429),
.B(n_1446),
.Y(n_1548)
);

O2A1O1Ixp5_ASAP7_75t_L g1549 ( 
.A1(n_1437),
.A2(n_1390),
.B(n_1452),
.C(n_1312),
.Y(n_1549)
);

NAND2xp5_ASAP7_75t_L g1550 ( 
.A(n_1394),
.B(n_1398),
.Y(n_1550)
);

NAND2xp5_ASAP7_75t_L g1551 ( 
.A(n_1394),
.B(n_1398),
.Y(n_1551)
);

HB1xp67_ASAP7_75t_L g1552 ( 
.A(n_1331),
.Y(n_1552)
);

OA21x2_ASAP7_75t_L g1553 ( 
.A1(n_1386),
.A2(n_1180),
.B(n_1424),
.Y(n_1553)
);

OAI22xp5_ASAP7_75t_L g1554 ( 
.A1(n_1434),
.A2(n_1307),
.B1(n_1312),
.B2(n_839),
.Y(n_1554)
);

AOI21xp5_ASAP7_75t_L g1555 ( 
.A1(n_1337),
.A2(n_1316),
.B(n_1310),
.Y(n_1555)
);

NOR2xp67_ASAP7_75t_L g1556 ( 
.A(n_1402),
.B(n_1340),
.Y(n_1556)
);

NAND2xp5_ASAP7_75t_L g1557 ( 
.A(n_1394),
.B(n_1398),
.Y(n_1557)
);

OAI22xp5_ASAP7_75t_L g1558 ( 
.A1(n_1434),
.A2(n_1307),
.B1(n_1312),
.B2(n_839),
.Y(n_1558)
);

OAI22xp5_ASAP7_75t_L g1559 ( 
.A1(n_1434),
.A2(n_1307),
.B1(n_1312),
.B2(n_839),
.Y(n_1559)
);

OA22x2_ASAP7_75t_L g1560 ( 
.A1(n_1452),
.A2(n_1237),
.B1(n_1309),
.B2(n_1133),
.Y(n_1560)
);

AND2x2_ASAP7_75t_L g1561 ( 
.A(n_1429),
.B(n_1446),
.Y(n_1561)
);

A2O1A1Ixp33_ASAP7_75t_L g1562 ( 
.A1(n_1452),
.A2(n_1307),
.B(n_1312),
.C(n_897),
.Y(n_1562)
);

OAI22xp5_ASAP7_75t_L g1563 ( 
.A1(n_1434),
.A2(n_1307),
.B1(n_1312),
.B2(n_839),
.Y(n_1563)
);

NAND2xp5_ASAP7_75t_L g1564 ( 
.A(n_1394),
.B(n_1398),
.Y(n_1564)
);

INVxp67_ASAP7_75t_L g1565 ( 
.A(n_1364),
.Y(n_1565)
);

AND2x2_ASAP7_75t_L g1566 ( 
.A(n_1429),
.B(n_1446),
.Y(n_1566)
);

OA21x2_ASAP7_75t_L g1567 ( 
.A1(n_1386),
.A2(n_1180),
.B(n_1424),
.Y(n_1567)
);

AOI21xp5_ASAP7_75t_L g1568 ( 
.A1(n_1337),
.A2(n_1316),
.B(n_1310),
.Y(n_1568)
);

INVx1_ASAP7_75t_L g1569 ( 
.A(n_1508),
.Y(n_1569)
);

BUFx2_ASAP7_75t_L g1570 ( 
.A(n_1512),
.Y(n_1570)
);

OAI21x1_ASAP7_75t_L g1571 ( 
.A1(n_1522),
.A2(n_1530),
.B(n_1527),
.Y(n_1571)
);

AND2x4_ASAP7_75t_L g1572 ( 
.A(n_1512),
.B(n_1487),
.Y(n_1572)
);

AND2x2_ASAP7_75t_L g1573 ( 
.A(n_1501),
.B(n_1502),
.Y(n_1573)
);

INVx1_ASAP7_75t_L g1574 ( 
.A(n_1508),
.Y(n_1574)
);

AND2x2_ASAP7_75t_L g1575 ( 
.A(n_1501),
.B(n_1502),
.Y(n_1575)
);

OR2x2_ASAP7_75t_L g1576 ( 
.A(n_1498),
.B(n_1520),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_1520),
.Y(n_1577)
);

NOR2xp33_ASAP7_75t_L g1578 ( 
.A(n_1485),
.B(n_1482),
.Y(n_1578)
);

OR2x6_ASAP7_75t_L g1579 ( 
.A(n_1487),
.B(n_1555),
.Y(n_1579)
);

BUFx2_ASAP7_75t_L g1580 ( 
.A(n_1514),
.Y(n_1580)
);

NAND2xp5_ASAP7_75t_L g1581 ( 
.A(n_1478),
.B(n_1550),
.Y(n_1581)
);

AND2x4_ASAP7_75t_L g1582 ( 
.A(n_1536),
.B(n_1499),
.Y(n_1582)
);

INVx1_ASAP7_75t_L g1583 ( 
.A(n_1526),
.Y(n_1583)
);

NAND2xp5_ASAP7_75t_L g1584 ( 
.A(n_1478),
.B(n_1550),
.Y(n_1584)
);

HB1xp67_ASAP7_75t_L g1585 ( 
.A(n_1506),
.Y(n_1585)
);

BUFx2_ASAP7_75t_SL g1586 ( 
.A(n_1556),
.Y(n_1586)
);

INVx1_ASAP7_75t_L g1587 ( 
.A(n_1526),
.Y(n_1587)
);

OR2x2_ASAP7_75t_L g1588 ( 
.A(n_1498),
.B(n_1494),
.Y(n_1588)
);

INVx1_ASAP7_75t_L g1589 ( 
.A(n_1528),
.Y(n_1589)
);

HB1xp67_ASAP7_75t_L g1590 ( 
.A(n_1484),
.Y(n_1590)
);

AND2x4_ASAP7_75t_L g1591 ( 
.A(n_1479),
.B(n_1503),
.Y(n_1591)
);

NAND2xp5_ASAP7_75t_L g1592 ( 
.A(n_1551),
.B(n_1557),
.Y(n_1592)
);

INVxp67_ASAP7_75t_SL g1593 ( 
.A(n_1551),
.Y(n_1593)
);

OR2x2_ASAP7_75t_L g1594 ( 
.A(n_1494),
.B(n_1557),
.Y(n_1594)
);

AOI21xp5_ASAP7_75t_SL g1595 ( 
.A1(n_1562),
.A2(n_1471),
.B(n_1472),
.Y(n_1595)
);

HB1xp67_ASAP7_75t_L g1596 ( 
.A(n_1552),
.Y(n_1596)
);

INVx1_ASAP7_75t_L g1597 ( 
.A(n_1491),
.Y(n_1597)
);

NOR2x1_ASAP7_75t_L g1598 ( 
.A(n_1473),
.B(n_1564),
.Y(n_1598)
);

AND2x2_ASAP7_75t_L g1599 ( 
.A(n_1553),
.B(n_1567),
.Y(n_1599)
);

INVx1_ASAP7_75t_L g1600 ( 
.A(n_1505),
.Y(n_1600)
);

AOI21xp5_ASAP7_75t_SL g1601 ( 
.A1(n_1474),
.A2(n_1554),
.B(n_1558),
.Y(n_1601)
);

OR2x2_ASAP7_75t_L g1602 ( 
.A(n_1564),
.B(n_1546),
.Y(n_1602)
);

INVx1_ASAP7_75t_SL g1603 ( 
.A(n_1483),
.Y(n_1603)
);

INVx2_ASAP7_75t_L g1604 ( 
.A(n_1489),
.Y(n_1604)
);

AND2x4_ASAP7_75t_L g1605 ( 
.A(n_1523),
.B(n_1500),
.Y(n_1605)
);

OA21x2_ASAP7_75t_L g1606 ( 
.A1(n_1516),
.A2(n_1568),
.B(n_1555),
.Y(n_1606)
);

INVx2_ASAP7_75t_L g1607 ( 
.A(n_1489),
.Y(n_1607)
);

INVx3_ASAP7_75t_L g1608 ( 
.A(n_1507),
.Y(n_1608)
);

AND2x2_ASAP7_75t_L g1609 ( 
.A(n_1496),
.B(n_1507),
.Y(n_1609)
);

INVx1_ASAP7_75t_L g1610 ( 
.A(n_1513),
.Y(n_1610)
);

AOI21xp5_ASAP7_75t_L g1611 ( 
.A1(n_1559),
.A2(n_1563),
.B(n_1549),
.Y(n_1611)
);

AO21x2_ASAP7_75t_L g1612 ( 
.A1(n_1544),
.A2(n_1497),
.B(n_1480),
.Y(n_1612)
);

INVx2_ASAP7_75t_L g1613 ( 
.A(n_1509),
.Y(n_1613)
);

AND2x2_ASAP7_75t_L g1614 ( 
.A(n_1477),
.B(n_1495),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_1519),
.Y(n_1615)
);

INVx1_ASAP7_75t_SL g1616 ( 
.A(n_1490),
.Y(n_1616)
);

OAI21xp5_ASAP7_75t_L g1617 ( 
.A1(n_1497),
.A2(n_1481),
.B(n_1560),
.Y(n_1617)
);

AOI21xp5_ASAP7_75t_L g1618 ( 
.A1(n_1482),
.A2(n_1535),
.B(n_1560),
.Y(n_1618)
);

NAND2xp5_ASAP7_75t_L g1619 ( 
.A(n_1525),
.B(n_1532),
.Y(n_1619)
);

INVx1_ASAP7_75t_L g1620 ( 
.A(n_1529),
.Y(n_1620)
);

INVx2_ASAP7_75t_SL g1621 ( 
.A(n_1533),
.Y(n_1621)
);

HB1xp67_ASAP7_75t_L g1622 ( 
.A(n_1524),
.Y(n_1622)
);

OR2x6_ASAP7_75t_L g1623 ( 
.A(n_1541),
.B(n_1539),
.Y(n_1623)
);

INVx2_ASAP7_75t_L g1624 ( 
.A(n_1613),
.Y(n_1624)
);

INVx1_ASAP7_75t_L g1625 ( 
.A(n_1597),
.Y(n_1625)
);

INVx1_ASAP7_75t_L g1626 ( 
.A(n_1597),
.Y(n_1626)
);

INVx1_ASAP7_75t_L g1627 ( 
.A(n_1600),
.Y(n_1627)
);

NAND2xp5_ASAP7_75t_L g1628 ( 
.A(n_1573),
.B(n_1545),
.Y(n_1628)
);

INVx1_ASAP7_75t_L g1629 ( 
.A(n_1600),
.Y(n_1629)
);

NAND2x1p5_ASAP7_75t_L g1630 ( 
.A(n_1598),
.B(n_1518),
.Y(n_1630)
);

AND2x2_ASAP7_75t_L g1631 ( 
.A(n_1575),
.B(n_1566),
.Y(n_1631)
);

NAND2xp5_ASAP7_75t_L g1632 ( 
.A(n_1575),
.B(n_1565),
.Y(n_1632)
);

BUFx2_ASAP7_75t_L g1633 ( 
.A(n_1605),
.Y(n_1633)
);

BUFx2_ASAP7_75t_L g1634 ( 
.A(n_1605),
.Y(n_1634)
);

AND2x2_ASAP7_75t_L g1635 ( 
.A(n_1575),
.B(n_1561),
.Y(n_1635)
);

INVxp67_ASAP7_75t_L g1636 ( 
.A(n_1593),
.Y(n_1636)
);

INVx3_ASAP7_75t_L g1637 ( 
.A(n_1608),
.Y(n_1637)
);

INVxp67_ASAP7_75t_L g1638 ( 
.A(n_1593),
.Y(n_1638)
);

AND2x2_ASAP7_75t_L g1639 ( 
.A(n_1599),
.B(n_1548),
.Y(n_1639)
);

NOR2xp33_ASAP7_75t_L g1640 ( 
.A(n_1601),
.B(n_1492),
.Y(n_1640)
);

AOI22xp33_ASAP7_75t_L g1641 ( 
.A1(n_1617),
.A2(n_1486),
.B1(n_1475),
.B2(n_1476),
.Y(n_1641)
);

AOI22xp33_ASAP7_75t_L g1642 ( 
.A1(n_1617),
.A2(n_1547),
.B1(n_1511),
.B2(n_1493),
.Y(n_1642)
);

INVxp67_ASAP7_75t_SL g1643 ( 
.A(n_1589),
.Y(n_1643)
);

INVx5_ASAP7_75t_SL g1644 ( 
.A(n_1623),
.Y(n_1644)
);

AND2x4_ASAP7_75t_SL g1645 ( 
.A(n_1623),
.B(n_1579),
.Y(n_1645)
);

OAI22xp5_ASAP7_75t_L g1646 ( 
.A1(n_1595),
.A2(n_1515),
.B1(n_1534),
.B2(n_1488),
.Y(n_1646)
);

INVxp67_ASAP7_75t_SL g1647 ( 
.A(n_1589),
.Y(n_1647)
);

AND2x2_ASAP7_75t_L g1648 ( 
.A(n_1609),
.B(n_1510),
.Y(n_1648)
);

AOI22xp5_ASAP7_75t_L g1649 ( 
.A1(n_1611),
.A2(n_1521),
.B1(n_1517),
.B2(n_1543),
.Y(n_1649)
);

NOR2xp33_ASAP7_75t_L g1650 ( 
.A(n_1594),
.B(n_1538),
.Y(n_1650)
);

AND2x2_ASAP7_75t_L g1651 ( 
.A(n_1609),
.B(n_1541),
.Y(n_1651)
);

HB1xp67_ASAP7_75t_L g1652 ( 
.A(n_1585),
.Y(n_1652)
);

INVx4_ASAP7_75t_L g1653 ( 
.A(n_1623),
.Y(n_1653)
);

OR2x2_ASAP7_75t_L g1654 ( 
.A(n_1576),
.B(n_1531),
.Y(n_1654)
);

INVx1_ASAP7_75t_L g1655 ( 
.A(n_1625),
.Y(n_1655)
);

OR2x2_ASAP7_75t_L g1656 ( 
.A(n_1628),
.B(n_1602),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1625),
.Y(n_1657)
);

AOI22xp5_ASAP7_75t_L g1658 ( 
.A1(n_1640),
.A2(n_1611),
.B1(n_1598),
.B2(n_1612),
.Y(n_1658)
);

INVx1_ASAP7_75t_L g1659 ( 
.A(n_1626),
.Y(n_1659)
);

INVx2_ASAP7_75t_L g1660 ( 
.A(n_1624),
.Y(n_1660)
);

OAI221xp5_ASAP7_75t_L g1661 ( 
.A1(n_1640),
.A2(n_1537),
.B1(n_1592),
.B2(n_1584),
.C(n_1581),
.Y(n_1661)
);

OAI31xp33_ASAP7_75t_L g1662 ( 
.A1(n_1646),
.A2(n_1641),
.A3(n_1642),
.B(n_1622),
.Y(n_1662)
);

INVxp67_ASAP7_75t_L g1663 ( 
.A(n_1628),
.Y(n_1663)
);

AOI222xp33_ASAP7_75t_L g1664 ( 
.A1(n_1641),
.A2(n_1622),
.B1(n_1581),
.B2(n_1592),
.C1(n_1584),
.C2(n_1619),
.Y(n_1664)
);

OAI21x1_ASAP7_75t_L g1665 ( 
.A1(n_1637),
.A2(n_1571),
.B(n_1608),
.Y(n_1665)
);

OAI221xp5_ASAP7_75t_L g1666 ( 
.A1(n_1642),
.A2(n_1618),
.B1(n_1594),
.B2(n_1602),
.C(n_1621),
.Y(n_1666)
);

AND2x2_ASAP7_75t_L g1667 ( 
.A(n_1639),
.B(n_1570),
.Y(n_1667)
);

AND2x2_ASAP7_75t_L g1668 ( 
.A(n_1639),
.B(n_1570),
.Y(n_1668)
);

OAI221xp5_ASAP7_75t_L g1669 ( 
.A1(n_1649),
.A2(n_1646),
.B1(n_1630),
.B2(n_1618),
.C(n_1621),
.Y(n_1669)
);

AND2x2_ASAP7_75t_L g1670 ( 
.A(n_1648),
.B(n_1580),
.Y(n_1670)
);

AOI221xp5_ASAP7_75t_L g1671 ( 
.A1(n_1636),
.A2(n_1616),
.B1(n_1590),
.B2(n_1596),
.C(n_1578),
.Y(n_1671)
);

NOR2xp33_ASAP7_75t_L g1672 ( 
.A(n_1632),
.B(n_1616),
.Y(n_1672)
);

AOI22xp33_ASAP7_75t_L g1673 ( 
.A1(n_1649),
.A2(n_1612),
.B1(n_1606),
.B2(n_1588),
.Y(n_1673)
);

AND2x2_ASAP7_75t_L g1674 ( 
.A(n_1648),
.B(n_1580),
.Y(n_1674)
);

OAI211xp5_ASAP7_75t_SL g1675 ( 
.A1(n_1636),
.A2(n_1588),
.B(n_1619),
.C(n_1621),
.Y(n_1675)
);

AOI21xp5_ASAP7_75t_L g1676 ( 
.A1(n_1645),
.A2(n_1623),
.B(n_1612),
.Y(n_1676)
);

OAI33xp33_ASAP7_75t_L g1677 ( 
.A1(n_1632),
.A2(n_1577),
.A3(n_1569),
.B1(n_1587),
.B2(n_1583),
.B3(n_1574),
.Y(n_1677)
);

AND2x2_ASAP7_75t_L g1678 ( 
.A(n_1639),
.B(n_1603),
.Y(n_1678)
);

NAND2xp33_ASAP7_75t_R g1679 ( 
.A(n_1651),
.B(n_1623),
.Y(n_1679)
);

OAI31xp33_ASAP7_75t_SL g1680 ( 
.A1(n_1651),
.A2(n_1582),
.A3(n_1572),
.B(n_1591),
.Y(n_1680)
);

NOR2xp33_ASAP7_75t_L g1681 ( 
.A(n_1631),
.B(n_1590),
.Y(n_1681)
);

INVx4_ASAP7_75t_L g1682 ( 
.A(n_1653),
.Y(n_1682)
);

OA21x2_ASAP7_75t_L g1683 ( 
.A1(n_1624),
.A2(n_1604),
.B(n_1607),
.Y(n_1683)
);

OAI221xp5_ASAP7_75t_L g1684 ( 
.A1(n_1630),
.A2(n_1623),
.B1(n_1579),
.B2(n_1596),
.C(n_1586),
.Y(n_1684)
);

AOI22xp33_ASAP7_75t_L g1685 ( 
.A1(n_1650),
.A2(n_1612),
.B1(n_1606),
.B2(n_1582),
.Y(n_1685)
);

INVx1_ASAP7_75t_L g1686 ( 
.A(n_1627),
.Y(n_1686)
);

NAND3xp33_ASAP7_75t_L g1687 ( 
.A(n_1638),
.B(n_1606),
.C(n_1582),
.Y(n_1687)
);

INVxp67_ASAP7_75t_L g1688 ( 
.A(n_1650),
.Y(n_1688)
);

AOI221xp5_ASAP7_75t_L g1689 ( 
.A1(n_1638),
.A2(n_1582),
.B1(n_1620),
.B2(n_1585),
.C(n_1610),
.Y(n_1689)
);

INVx1_ASAP7_75t_L g1690 ( 
.A(n_1629),
.Y(n_1690)
);

AOI222xp33_ASAP7_75t_L g1691 ( 
.A1(n_1631),
.A2(n_1582),
.B1(n_1504),
.B2(n_1614),
.C1(n_1620),
.C2(n_1615),
.Y(n_1691)
);

AO21x2_ASAP7_75t_L g1692 ( 
.A1(n_1643),
.A2(n_1607),
.B(n_1604),
.Y(n_1692)
);

AND2x2_ASAP7_75t_SL g1693 ( 
.A(n_1645),
.B(n_1606),
.Y(n_1693)
);

BUFx3_ASAP7_75t_L g1694 ( 
.A(n_1654),
.Y(n_1694)
);

OR2x6_ASAP7_75t_L g1695 ( 
.A(n_1653),
.B(n_1579),
.Y(n_1695)
);

AND2x4_ASAP7_75t_SL g1696 ( 
.A(n_1653),
.B(n_1572),
.Y(n_1696)
);

INVx1_ASAP7_75t_L g1697 ( 
.A(n_1655),
.Y(n_1697)
);

NOR2xp33_ASAP7_75t_L g1698 ( 
.A(n_1688),
.B(n_1631),
.Y(n_1698)
);

AND2x2_ASAP7_75t_L g1699 ( 
.A(n_1667),
.B(n_1633),
.Y(n_1699)
);

HB1xp67_ASAP7_75t_L g1700 ( 
.A(n_1692),
.Y(n_1700)
);

INVx2_ASAP7_75t_L g1701 ( 
.A(n_1683),
.Y(n_1701)
);

INVx1_ASAP7_75t_L g1702 ( 
.A(n_1657),
.Y(n_1702)
);

BUFx3_ASAP7_75t_L g1703 ( 
.A(n_1692),
.Y(n_1703)
);

INVx4_ASAP7_75t_L g1704 ( 
.A(n_1682),
.Y(n_1704)
);

INVx2_ASAP7_75t_L g1705 ( 
.A(n_1660),
.Y(n_1705)
);

OR2x6_ASAP7_75t_L g1706 ( 
.A(n_1695),
.B(n_1653),
.Y(n_1706)
);

NOR2xp33_ASAP7_75t_L g1707 ( 
.A(n_1661),
.B(n_1635),
.Y(n_1707)
);

INVx2_ASAP7_75t_L g1708 ( 
.A(n_1665),
.Y(n_1708)
);

BUFx3_ASAP7_75t_L g1709 ( 
.A(n_1682),
.Y(n_1709)
);

INVx2_ASAP7_75t_SL g1710 ( 
.A(n_1696),
.Y(n_1710)
);

INVx2_ASAP7_75t_SL g1711 ( 
.A(n_1696),
.Y(n_1711)
);

INVx2_ASAP7_75t_L g1712 ( 
.A(n_1659),
.Y(n_1712)
);

NAND3xp33_ASAP7_75t_SL g1713 ( 
.A(n_1662),
.B(n_1630),
.C(n_1651),
.Y(n_1713)
);

INVx1_ASAP7_75t_L g1714 ( 
.A(n_1686),
.Y(n_1714)
);

NAND2xp5_ASAP7_75t_SL g1715 ( 
.A(n_1658),
.B(n_1630),
.Y(n_1715)
);

INVx1_ASAP7_75t_L g1716 ( 
.A(n_1690),
.Y(n_1716)
);

NOR2x1p5_ASAP7_75t_L g1717 ( 
.A(n_1687),
.B(n_1643),
.Y(n_1717)
);

INVx2_ASAP7_75t_L g1718 ( 
.A(n_1694),
.Y(n_1718)
);

INVx2_ASAP7_75t_L g1719 ( 
.A(n_1694),
.Y(n_1719)
);

BUFx6f_ASAP7_75t_L g1720 ( 
.A(n_1693),
.Y(n_1720)
);

INVx1_ASAP7_75t_L g1721 ( 
.A(n_1668),
.Y(n_1721)
);

INVx2_ASAP7_75t_L g1722 ( 
.A(n_1693),
.Y(n_1722)
);

INVx1_ASAP7_75t_L g1723 ( 
.A(n_1656),
.Y(n_1723)
);

INVx2_ASAP7_75t_L g1724 ( 
.A(n_1682),
.Y(n_1724)
);

BUFx2_ASAP7_75t_L g1725 ( 
.A(n_1695),
.Y(n_1725)
);

INVx1_ASAP7_75t_L g1726 ( 
.A(n_1697),
.Y(n_1726)
);

OR2x2_ASAP7_75t_L g1727 ( 
.A(n_1723),
.B(n_1647),
.Y(n_1727)
);

INVx1_ASAP7_75t_L g1728 ( 
.A(n_1697),
.Y(n_1728)
);

NAND4xp25_ASAP7_75t_L g1729 ( 
.A(n_1713),
.B(n_1673),
.C(n_1669),
.D(n_1685),
.Y(n_1729)
);

AOI221xp5_ASAP7_75t_L g1730 ( 
.A1(n_1713),
.A2(n_1666),
.B1(n_1673),
.B2(n_1671),
.C(n_1675),
.Y(n_1730)
);

INVx1_ASAP7_75t_L g1731 ( 
.A(n_1697),
.Y(n_1731)
);

INVx1_ASAP7_75t_L g1732 ( 
.A(n_1702),
.Y(n_1732)
);

NAND2xp5_ASAP7_75t_L g1733 ( 
.A(n_1707),
.B(n_1672),
.Y(n_1733)
);

NOR2xp33_ASAP7_75t_L g1734 ( 
.A(n_1707),
.B(n_1663),
.Y(n_1734)
);

HB1xp67_ASAP7_75t_L g1735 ( 
.A(n_1718),
.Y(n_1735)
);

AND2x2_ASAP7_75t_L g1736 ( 
.A(n_1725),
.B(n_1680),
.Y(n_1736)
);

INVx1_ASAP7_75t_L g1737 ( 
.A(n_1702),
.Y(n_1737)
);

INVx1_ASAP7_75t_L g1738 ( 
.A(n_1702),
.Y(n_1738)
);

AND2x2_ASAP7_75t_L g1739 ( 
.A(n_1725),
.B(n_1678),
.Y(n_1739)
);

INVx1_ASAP7_75t_L g1740 ( 
.A(n_1714),
.Y(n_1740)
);

OR2x2_ASAP7_75t_L g1741 ( 
.A(n_1723),
.B(n_1647),
.Y(n_1741)
);

INVx1_ASAP7_75t_L g1742 ( 
.A(n_1714),
.Y(n_1742)
);

INVx2_ASAP7_75t_L g1743 ( 
.A(n_1703),
.Y(n_1743)
);

OAI221xp5_ASAP7_75t_L g1744 ( 
.A1(n_1715),
.A2(n_1685),
.B1(n_1684),
.B2(n_1664),
.C(n_1679),
.Y(n_1744)
);

NAND2xp5_ASAP7_75t_L g1745 ( 
.A(n_1698),
.B(n_1672),
.Y(n_1745)
);

AND2x4_ASAP7_75t_L g1746 ( 
.A(n_1709),
.B(n_1634),
.Y(n_1746)
);

INVx1_ASAP7_75t_L g1747 ( 
.A(n_1714),
.Y(n_1747)
);

INVx2_ASAP7_75t_L g1748 ( 
.A(n_1703),
.Y(n_1748)
);

AND2x2_ASAP7_75t_L g1749 ( 
.A(n_1725),
.B(n_1678),
.Y(n_1749)
);

AND2x2_ASAP7_75t_L g1750 ( 
.A(n_1710),
.B(n_1670),
.Y(n_1750)
);

OR2x2_ASAP7_75t_L g1751 ( 
.A(n_1723),
.B(n_1652),
.Y(n_1751)
);

INVx2_ASAP7_75t_L g1752 ( 
.A(n_1703),
.Y(n_1752)
);

NAND2xp5_ASAP7_75t_L g1753 ( 
.A(n_1698),
.B(n_1681),
.Y(n_1753)
);

OR2x6_ASAP7_75t_L g1754 ( 
.A(n_1704),
.B(n_1676),
.Y(n_1754)
);

INVx1_ASAP7_75t_L g1755 ( 
.A(n_1716),
.Y(n_1755)
);

INVx1_ASAP7_75t_L g1756 ( 
.A(n_1716),
.Y(n_1756)
);

AOI22xp33_ASAP7_75t_L g1757 ( 
.A1(n_1715),
.A2(n_1579),
.B1(n_1645),
.B2(n_1644),
.Y(n_1757)
);

NAND2x1_ASAP7_75t_L g1758 ( 
.A(n_1710),
.B(n_1711),
.Y(n_1758)
);

INVx2_ASAP7_75t_L g1759 ( 
.A(n_1703),
.Y(n_1759)
);

AND2x4_ASAP7_75t_L g1760 ( 
.A(n_1709),
.B(n_1634),
.Y(n_1760)
);

OR2x2_ASAP7_75t_L g1761 ( 
.A(n_1721),
.B(n_1652),
.Y(n_1761)
);

INVx2_ASAP7_75t_L g1762 ( 
.A(n_1705),
.Y(n_1762)
);

NOR3xp33_ASAP7_75t_L g1763 ( 
.A(n_1704),
.B(n_1677),
.C(n_1689),
.Y(n_1763)
);

AND2x2_ASAP7_75t_L g1764 ( 
.A(n_1710),
.B(n_1674),
.Y(n_1764)
);

INVx2_ASAP7_75t_L g1765 ( 
.A(n_1705),
.Y(n_1765)
);

NAND2xp5_ASAP7_75t_L g1766 ( 
.A(n_1718),
.B(n_1681),
.Y(n_1766)
);

INVx2_ASAP7_75t_L g1767 ( 
.A(n_1705),
.Y(n_1767)
);

NAND2xp5_ASAP7_75t_L g1768 ( 
.A(n_1718),
.B(n_1635),
.Y(n_1768)
);

OR2x2_ASAP7_75t_L g1769 ( 
.A(n_1751),
.B(n_1718),
.Y(n_1769)
);

INVx1_ASAP7_75t_L g1770 ( 
.A(n_1726),
.Y(n_1770)
);

OR2x2_ASAP7_75t_L g1771 ( 
.A(n_1751),
.B(n_1719),
.Y(n_1771)
);

INVx1_ASAP7_75t_L g1772 ( 
.A(n_1726),
.Y(n_1772)
);

OR2x2_ASAP7_75t_L g1773 ( 
.A(n_1727),
.B(n_1741),
.Y(n_1773)
);

INVx2_ASAP7_75t_L g1774 ( 
.A(n_1743),
.Y(n_1774)
);

AND2x2_ASAP7_75t_L g1775 ( 
.A(n_1736),
.B(n_1719),
.Y(n_1775)
);

INVx1_ASAP7_75t_L g1776 ( 
.A(n_1728),
.Y(n_1776)
);

OR2x2_ASAP7_75t_L g1777 ( 
.A(n_1727),
.B(n_1719),
.Y(n_1777)
);

OR2x2_ASAP7_75t_L g1778 ( 
.A(n_1741),
.B(n_1719),
.Y(n_1778)
);

AND2x2_ASAP7_75t_L g1779 ( 
.A(n_1736),
.B(n_1711),
.Y(n_1779)
);

NAND2xp5_ASAP7_75t_L g1780 ( 
.A(n_1734),
.B(n_1721),
.Y(n_1780)
);

NAND2xp5_ASAP7_75t_L g1781 ( 
.A(n_1733),
.B(n_1721),
.Y(n_1781)
);

INVx1_ASAP7_75t_SL g1782 ( 
.A(n_1758),
.Y(n_1782)
);

NAND2xp5_ASAP7_75t_L g1783 ( 
.A(n_1763),
.B(n_1717),
.Y(n_1783)
);

INVx1_ASAP7_75t_L g1784 ( 
.A(n_1728),
.Y(n_1784)
);

AOI22xp33_ASAP7_75t_L g1785 ( 
.A1(n_1729),
.A2(n_1744),
.B1(n_1730),
.B2(n_1717),
.Y(n_1785)
);

INVx1_ASAP7_75t_L g1786 ( 
.A(n_1731),
.Y(n_1786)
);

INVx2_ASAP7_75t_L g1787 ( 
.A(n_1743),
.Y(n_1787)
);

AND2x2_ASAP7_75t_L g1788 ( 
.A(n_1739),
.B(n_1749),
.Y(n_1788)
);

INVx3_ASAP7_75t_L g1789 ( 
.A(n_1758),
.Y(n_1789)
);

AND2x4_ASAP7_75t_L g1790 ( 
.A(n_1739),
.B(n_1704),
.Y(n_1790)
);

NAND2xp5_ASAP7_75t_L g1791 ( 
.A(n_1745),
.B(n_1717),
.Y(n_1791)
);

AND2x2_ASAP7_75t_L g1792 ( 
.A(n_1749),
.B(n_1750),
.Y(n_1792)
);

INVx4_ASAP7_75t_L g1793 ( 
.A(n_1748),
.Y(n_1793)
);

NAND2xp5_ASAP7_75t_SL g1794 ( 
.A(n_1757),
.B(n_1720),
.Y(n_1794)
);

OAI32xp33_ASAP7_75t_L g1795 ( 
.A1(n_1766),
.A2(n_1700),
.A3(n_1679),
.B1(n_1722),
.B2(n_1709),
.Y(n_1795)
);

NAND2x1_ASAP7_75t_L g1796 ( 
.A(n_1754),
.B(n_1711),
.Y(n_1796)
);

AND2x2_ASAP7_75t_L g1797 ( 
.A(n_1750),
.B(n_1724),
.Y(n_1797)
);

OR2x6_ASAP7_75t_L g1798 ( 
.A(n_1754),
.B(n_1586),
.Y(n_1798)
);

INVx2_ASAP7_75t_SL g1799 ( 
.A(n_1764),
.Y(n_1799)
);

OR2x2_ASAP7_75t_L g1800 ( 
.A(n_1768),
.B(n_1712),
.Y(n_1800)
);

INVxp67_ASAP7_75t_L g1801 ( 
.A(n_1735),
.Y(n_1801)
);

NAND2xp5_ASAP7_75t_L g1802 ( 
.A(n_1753),
.B(n_1635),
.Y(n_1802)
);

NAND2xp5_ASAP7_75t_L g1803 ( 
.A(n_1764),
.B(n_1699),
.Y(n_1803)
);

INVx2_ASAP7_75t_L g1804 ( 
.A(n_1748),
.Y(n_1804)
);

NAND2xp5_ASAP7_75t_L g1805 ( 
.A(n_1785),
.B(n_1755),
.Y(n_1805)
);

INVxp67_ASAP7_75t_L g1806 ( 
.A(n_1779),
.Y(n_1806)
);

OAI21xp5_ASAP7_75t_L g1807 ( 
.A1(n_1783),
.A2(n_1759),
.B(n_1752),
.Y(n_1807)
);

NAND3xp33_ASAP7_75t_L g1808 ( 
.A(n_1801),
.B(n_1759),
.C(n_1752),
.Y(n_1808)
);

INVx2_ASAP7_75t_L g1809 ( 
.A(n_1792),
.Y(n_1809)
);

INVx1_ASAP7_75t_L g1810 ( 
.A(n_1770),
.Y(n_1810)
);

AND2x2_ASAP7_75t_L g1811 ( 
.A(n_1788),
.B(n_1746),
.Y(n_1811)
);

INVx2_ASAP7_75t_L g1812 ( 
.A(n_1792),
.Y(n_1812)
);

AND2x4_ASAP7_75t_L g1813 ( 
.A(n_1789),
.B(n_1731),
.Y(n_1813)
);

OAI22xp5_ASAP7_75t_L g1814 ( 
.A1(n_1791),
.A2(n_1720),
.B1(n_1644),
.B2(n_1754),
.Y(n_1814)
);

HB1xp67_ASAP7_75t_L g1815 ( 
.A(n_1788),
.Y(n_1815)
);

INVx1_ASAP7_75t_L g1816 ( 
.A(n_1772),
.Y(n_1816)
);

NAND2xp5_ASAP7_75t_L g1817 ( 
.A(n_1775),
.B(n_1724),
.Y(n_1817)
);

INVx1_ASAP7_75t_L g1818 ( 
.A(n_1776),
.Y(n_1818)
);

AND2x2_ASAP7_75t_L g1819 ( 
.A(n_1779),
.B(n_1746),
.Y(n_1819)
);

AND2x2_ASAP7_75t_L g1820 ( 
.A(n_1775),
.B(n_1746),
.Y(n_1820)
);

AND2x2_ASAP7_75t_L g1821 ( 
.A(n_1799),
.B(n_1760),
.Y(n_1821)
);

INVx1_ASAP7_75t_L g1822 ( 
.A(n_1784),
.Y(n_1822)
);

INVxp67_ASAP7_75t_L g1823 ( 
.A(n_1799),
.Y(n_1823)
);

OR2x6_ASAP7_75t_L g1824 ( 
.A(n_1796),
.B(n_1754),
.Y(n_1824)
);

HB1xp67_ASAP7_75t_L g1825 ( 
.A(n_1789),
.Y(n_1825)
);

AO21x2_ASAP7_75t_L g1826 ( 
.A1(n_1774),
.A2(n_1700),
.B(n_1738),
.Y(n_1826)
);

AND2x2_ASAP7_75t_L g1827 ( 
.A(n_1782),
.B(n_1760),
.Y(n_1827)
);

NOR2xp33_ASAP7_75t_L g1828 ( 
.A(n_1780),
.B(n_1724),
.Y(n_1828)
);

INVx1_ASAP7_75t_L g1829 ( 
.A(n_1786),
.Y(n_1829)
);

INVx1_ASAP7_75t_L g1830 ( 
.A(n_1773),
.Y(n_1830)
);

AND2x2_ASAP7_75t_L g1831 ( 
.A(n_1797),
.B(n_1760),
.Y(n_1831)
);

INVx1_ASAP7_75t_L g1832 ( 
.A(n_1815),
.Y(n_1832)
);

INVx2_ASAP7_75t_L g1833 ( 
.A(n_1825),
.Y(n_1833)
);

OAI21xp33_ASAP7_75t_L g1834 ( 
.A1(n_1805),
.A2(n_1794),
.B(n_1795),
.Y(n_1834)
);

AOI22xp33_ASAP7_75t_L g1835 ( 
.A1(n_1805),
.A2(n_1790),
.B1(n_1781),
.B2(n_1789),
.Y(n_1835)
);

AOI21xp5_ASAP7_75t_L g1836 ( 
.A1(n_1807),
.A2(n_1795),
.B(n_1796),
.Y(n_1836)
);

NOR2xp33_ASAP7_75t_L g1837 ( 
.A(n_1806),
.B(n_1790),
.Y(n_1837)
);

NAND2xp5_ASAP7_75t_L g1838 ( 
.A(n_1823),
.B(n_1797),
.Y(n_1838)
);

AND2x2_ASAP7_75t_L g1839 ( 
.A(n_1819),
.B(n_1790),
.Y(n_1839)
);

NAND2xp5_ASAP7_75t_L g1840 ( 
.A(n_1830),
.B(n_1803),
.Y(n_1840)
);

INVx1_ASAP7_75t_L g1841 ( 
.A(n_1809),
.Y(n_1841)
);

INVx1_ASAP7_75t_L g1842 ( 
.A(n_1809),
.Y(n_1842)
);

INVx2_ASAP7_75t_L g1843 ( 
.A(n_1820),
.Y(n_1843)
);

AOI211xp5_ASAP7_75t_SL g1844 ( 
.A1(n_1814),
.A2(n_1804),
.B(n_1774),
.C(n_1787),
.Y(n_1844)
);

AOI21xp33_ASAP7_75t_L g1845 ( 
.A1(n_1807),
.A2(n_1798),
.B(n_1771),
.Y(n_1845)
);

AOI21xp5_ASAP7_75t_L g1846 ( 
.A1(n_1808),
.A2(n_1798),
.B(n_1771),
.Y(n_1846)
);

INVx1_ASAP7_75t_L g1847 ( 
.A(n_1809),
.Y(n_1847)
);

INVx1_ASAP7_75t_L g1848 ( 
.A(n_1812),
.Y(n_1848)
);

AOI221xp5_ASAP7_75t_L g1849 ( 
.A1(n_1808),
.A2(n_1793),
.B1(n_1804),
.B2(n_1787),
.C(n_1773),
.Y(n_1849)
);

AOI221xp5_ASAP7_75t_L g1850 ( 
.A1(n_1828),
.A2(n_1793),
.B1(n_1769),
.B2(n_1778),
.C(n_1777),
.Y(n_1850)
);

AND2x2_ASAP7_75t_L g1851 ( 
.A(n_1819),
.B(n_1793),
.Y(n_1851)
);

NAND2xp5_ASAP7_75t_L g1852 ( 
.A(n_1830),
.B(n_1802),
.Y(n_1852)
);

AOI322xp5_ASAP7_75t_L g1853 ( 
.A1(n_1812),
.A2(n_1722),
.A3(n_1720),
.B1(n_1742),
.B2(n_1737),
.C1(n_1738),
.C2(n_1747),
.Y(n_1853)
);

NAND2xp5_ASAP7_75t_L g1854 ( 
.A(n_1843),
.B(n_1812),
.Y(n_1854)
);

NAND2xp5_ASAP7_75t_L g1855 ( 
.A(n_1843),
.B(n_1820),
.Y(n_1855)
);

NOR2xp33_ASAP7_75t_L g1856 ( 
.A(n_1832),
.B(n_1827),
.Y(n_1856)
);

OR2x6_ASAP7_75t_L g1857 ( 
.A(n_1833),
.B(n_1824),
.Y(n_1857)
);

NOR2xp33_ASAP7_75t_L g1858 ( 
.A(n_1834),
.B(n_1827),
.Y(n_1858)
);

INVx1_ASAP7_75t_L g1859 ( 
.A(n_1841),
.Y(n_1859)
);

NOR2x1p5_ASAP7_75t_L g1860 ( 
.A(n_1838),
.B(n_1817),
.Y(n_1860)
);

NOR2x1_ASAP7_75t_L g1861 ( 
.A(n_1833),
.B(n_1824),
.Y(n_1861)
);

AOI22xp33_ASAP7_75t_SL g1862 ( 
.A1(n_1836),
.A2(n_1811),
.B1(n_1814),
.B2(n_1831),
.Y(n_1862)
);

NOR2xp33_ASAP7_75t_SL g1863 ( 
.A(n_1851),
.B(n_1821),
.Y(n_1863)
);

NAND2xp5_ASAP7_75t_L g1864 ( 
.A(n_1835),
.B(n_1811),
.Y(n_1864)
);

OAI22xp5_ASAP7_75t_L g1865 ( 
.A1(n_1835),
.A2(n_1824),
.B1(n_1720),
.B2(n_1831),
.Y(n_1865)
);

AOI221xp5_ASAP7_75t_L g1866 ( 
.A1(n_1858),
.A2(n_1849),
.B1(n_1850),
.B2(n_1845),
.C(n_1837),
.Y(n_1866)
);

NAND2xp5_ASAP7_75t_SL g1867 ( 
.A(n_1863),
.B(n_1851),
.Y(n_1867)
);

OA22x2_ASAP7_75t_L g1868 ( 
.A1(n_1857),
.A2(n_1839),
.B1(n_1848),
.B2(n_1847),
.Y(n_1868)
);

AOI21xp5_ASAP7_75t_L g1869 ( 
.A1(n_1861),
.A2(n_1846),
.B(n_1844),
.Y(n_1869)
);

NOR4xp25_ASAP7_75t_L g1870 ( 
.A(n_1859),
.B(n_1842),
.C(n_1837),
.D(n_1840),
.Y(n_1870)
);

OAI221xp5_ASAP7_75t_L g1871 ( 
.A1(n_1862),
.A2(n_1852),
.B1(n_1853),
.B2(n_1824),
.C(n_1798),
.Y(n_1871)
);

AOI22xp33_ASAP7_75t_L g1872 ( 
.A1(n_1856),
.A2(n_1824),
.B1(n_1821),
.B2(n_1798),
.Y(n_1872)
);

NAND3xp33_ASAP7_75t_L g1873 ( 
.A(n_1865),
.B(n_1816),
.C(n_1810),
.Y(n_1873)
);

AOI21xp5_ASAP7_75t_L g1874 ( 
.A1(n_1864),
.A2(n_1813),
.B(n_1810),
.Y(n_1874)
);

AOI222xp33_ASAP7_75t_L g1875 ( 
.A1(n_1860),
.A2(n_1829),
.B1(n_1822),
.B2(n_1818),
.C1(n_1816),
.C2(n_1813),
.Y(n_1875)
);

OAI21xp33_ASAP7_75t_SL g1876 ( 
.A1(n_1869),
.A2(n_1857),
.B(n_1854),
.Y(n_1876)
);

INVx1_ASAP7_75t_L g1877 ( 
.A(n_1868),
.Y(n_1877)
);

OAI22xp33_ASAP7_75t_L g1878 ( 
.A1(n_1871),
.A2(n_1855),
.B1(n_1720),
.B2(n_1769),
.Y(n_1878)
);

AOI21xp5_ASAP7_75t_L g1879 ( 
.A1(n_1867),
.A2(n_1822),
.B(n_1818),
.Y(n_1879)
);

AOI211xp5_ASAP7_75t_SL g1880 ( 
.A1(n_1866),
.A2(n_1829),
.B(n_1813),
.C(n_1777),
.Y(n_1880)
);

AOI21xp5_ASAP7_75t_L g1881 ( 
.A1(n_1874),
.A2(n_1813),
.B(n_1826),
.Y(n_1881)
);

NOR2xp67_ASAP7_75t_L g1882 ( 
.A(n_1879),
.B(n_1873),
.Y(n_1882)
);

NAND2xp5_ASAP7_75t_L g1883 ( 
.A(n_1880),
.B(n_1870),
.Y(n_1883)
);

INVx1_ASAP7_75t_L g1884 ( 
.A(n_1877),
.Y(n_1884)
);

NOR2x1_ASAP7_75t_L g1885 ( 
.A(n_1881),
.B(n_1826),
.Y(n_1885)
);

NAND2xp5_ASAP7_75t_L g1886 ( 
.A(n_1876),
.B(n_1875),
.Y(n_1886)
);

NOR2xp33_ASAP7_75t_L g1887 ( 
.A(n_1878),
.B(n_1872),
.Y(n_1887)
);

OR3x2_ASAP7_75t_L g1888 ( 
.A(n_1877),
.B(n_1778),
.C(n_1800),
.Y(n_1888)
);

A2O1A1Ixp33_ASAP7_75t_L g1889 ( 
.A1(n_1882),
.A2(n_1883),
.B(n_1885),
.C(n_1886),
.Y(n_1889)
);

NOR2xp33_ASAP7_75t_R g1890 ( 
.A(n_1884),
.B(n_1709),
.Y(n_1890)
);

INVx1_ASAP7_75t_L g1891 ( 
.A(n_1888),
.Y(n_1891)
);

CKINVDCx5p33_ASAP7_75t_R g1892 ( 
.A(n_1887),
.Y(n_1892)
);

NOR2xp67_ASAP7_75t_L g1893 ( 
.A(n_1882),
.B(n_1732),
.Y(n_1893)
);

AOI211xp5_ASAP7_75t_L g1894 ( 
.A1(n_1883),
.A2(n_1540),
.B(n_1720),
.C(n_1800),
.Y(n_1894)
);

AND2x2_ASAP7_75t_SL g1895 ( 
.A(n_1891),
.B(n_1542),
.Y(n_1895)
);

NOR2x1_ASAP7_75t_L g1896 ( 
.A(n_1893),
.B(n_1826),
.Y(n_1896)
);

NAND3x1_ASAP7_75t_L g1897 ( 
.A(n_1892),
.B(n_1732),
.C(n_1737),
.Y(n_1897)
);

BUFx6f_ASAP7_75t_L g1898 ( 
.A(n_1895),
.Y(n_1898)
);

AOI322xp5_ASAP7_75t_L g1899 ( 
.A1(n_1898),
.A2(n_1889),
.A3(n_1896),
.B1(n_1890),
.B2(n_1894),
.C1(n_1897),
.C2(n_1722),
.Y(n_1899)
);

OAI21xp5_ASAP7_75t_L g1900 ( 
.A1(n_1899),
.A2(n_1898),
.B(n_1724),
.Y(n_1900)
);

XNOR2xp5_ASAP7_75t_L g1901 ( 
.A(n_1899),
.B(n_1898),
.Y(n_1901)
);

NAND4xp25_ASAP7_75t_L g1902 ( 
.A(n_1900),
.B(n_1898),
.C(n_1704),
.D(n_1691),
.Y(n_1902)
);

NOR4xp25_ASAP7_75t_L g1903 ( 
.A(n_1901),
.B(n_1740),
.C(n_1742),
.D(n_1747),
.Y(n_1903)
);

AOI22xp5_ASAP7_75t_L g1904 ( 
.A1(n_1902),
.A2(n_1903),
.B1(n_1826),
.B2(n_1756),
.Y(n_1904)
);

AOI22xp5_ASAP7_75t_L g1905 ( 
.A1(n_1902),
.A2(n_1756),
.B1(n_1740),
.B2(n_1704),
.Y(n_1905)
);

AOI222xp33_ASAP7_75t_SL g1906 ( 
.A1(n_1905),
.A2(n_1904),
.B1(n_1722),
.B2(n_1767),
.C1(n_1765),
.C2(n_1762),
.Y(n_1906)
);

XNOR2x1_ASAP7_75t_L g1907 ( 
.A(n_1906),
.B(n_1706),
.Y(n_1907)
);

AOI22xp5_ASAP7_75t_L g1908 ( 
.A1(n_1907),
.A2(n_1767),
.B1(n_1765),
.B2(n_1762),
.Y(n_1908)
);

XNOR2xp5_ASAP7_75t_L g1909 ( 
.A(n_1908),
.B(n_1706),
.Y(n_1909)
);

AOI221xp5_ASAP7_75t_L g1910 ( 
.A1(n_1909),
.A2(n_1704),
.B1(n_1708),
.B2(n_1720),
.C(n_1701),
.Y(n_1910)
);

AOI211xp5_ASAP7_75t_L g1911 ( 
.A1(n_1910),
.A2(n_1708),
.B(n_1720),
.C(n_1761),
.Y(n_1911)
);


endmodule