module real_jpeg_26861_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_201;
wire n_114;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_83;
wire n_78;
wire n_249;
wire n_166;
wire n_176;
wire n_221;
wire n_300;
wire n_215;
wire n_286;
wire n_288;
wire n_292;
wire n_194;
wire n_153;
wire n_104;
wire n_161;
wire n_207;
wire n_301;
wire n_280;
wire n_64;
wire n_177;
wire n_291;
wire n_236;
wire n_47;
wire n_131;
wire n_281;
wire n_271;
wire n_163;
wire n_276;
wire n_22;
wire n_287;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_299;
wire n_173;
wire n_255;
wire n_115;
wire n_243;
wire n_98;
wire n_27;
wire n_56;
wire n_200;
wire n_48;
wire n_164;
wire n_293;
wire n_184;
wire n_275;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_290;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_285;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_262;
wire n_222;
wire n_118;
wire n_220;
wire n_294;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_298;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_296;
wire n_134;
wire n_270;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_198;
wire n_192;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_110;
wire n_61;
wire n_205;
wire n_195;
wire n_258;
wire n_289;
wire n_117;
wire n_193;
wire n_99;
wire n_261;
wire n_86;
wire n_150;
wire n_41;
wire n_70;
wire n_74;
wire n_32;
wire n_20;
wire n_80;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_103;
wire n_259;
wire n_225;
wire n_232;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_284;
wire n_226;
wire n_277;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_297;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_279;
wire n_59;
wire n_169;
wire n_167;
wire n_128;
wire n_295;
wire n_179;
wire n_202;
wire n_213;
wire n_133;
wire n_216;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_283;
wire n_181;
wire n_101;
wire n_256;
wire n_274;
wire n_182;
wire n_253;
wire n_96;
wire n_269;
wire n_273;
wire n_89;

AOI22xp33_ASAP7_75t_SL g39 ( 
.A1(n_0),
.A2(n_29),
.B1(n_30),
.B2(n_40),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_0),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_0),
.A2(n_32),
.B1(n_33),
.B2(n_40),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_0),
.A2(n_40),
.B1(n_47),
.B2(n_48),
.Y(n_136)
);

INVx11_ASAP7_75t_L g88 ( 
.A(n_1),
.Y(n_88)
);

INVx5_ASAP7_75t_L g89 ( 
.A(n_1),
.Y(n_89)
);

HB1xp67_ASAP7_75t_L g140 ( 
.A(n_1),
.Y(n_140)
);

AOI21xp5_ASAP7_75t_L g182 ( 
.A1(n_1),
.A2(n_110),
.B(n_170),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g37 ( 
.A1(n_2),
.A2(n_29),
.B1(n_30),
.B2(n_38),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_2),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_2),
.A2(n_38),
.B1(n_75),
.B2(n_76),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_2),
.A2(n_32),
.B1(n_33),
.B2(n_38),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_2),
.A2(n_38),
.B1(n_47),
.B2(n_48),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_3),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_3),
.B(n_29),
.Y(n_193)
);

AOI21xp33_ASAP7_75t_L g197 ( 
.A1(n_3),
.A2(n_29),
.B(n_193),
.Y(n_197)
);

AOI22xp33_ASAP7_75t_SL g217 ( 
.A1(n_3),
.A2(n_32),
.B1(n_33),
.B2(n_151),
.Y(n_217)
);

AOI21xp5_ASAP7_75t_L g220 ( 
.A1(n_3),
.A2(n_11),
.B(n_47),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_3),
.B(n_117),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_L g243 ( 
.A1(n_3),
.A2(n_87),
.B1(n_88),
.B2(n_241),
.Y(n_243)
);

BUFx12_ASAP7_75t_L g73 ( 
.A(n_4),
.Y(n_73)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

INVx13_ASAP7_75t_L g75 ( 
.A(n_6),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_7),
.A2(n_75),
.B1(n_76),
.B2(n_123),
.Y(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_7),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_7),
.A2(n_29),
.B1(n_30),
.B2(n_123),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_SL g201 ( 
.A1(n_7),
.A2(n_32),
.B1(n_33),
.B2(n_123),
.Y(n_201)
);

AOI22xp33_ASAP7_75t_SL g228 ( 
.A1(n_7),
.A2(n_47),
.B1(n_48),
.B2(n_123),
.Y(n_228)
);

OAI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_8),
.A2(n_32),
.B1(n_33),
.B2(n_56),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_8),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_L g68 ( 
.A1(n_8),
.A2(n_29),
.B1(n_30),
.B2(n_56),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_L g81 ( 
.A1(n_8),
.A2(n_56),
.B1(n_75),
.B2(n_76),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_L g111 ( 
.A1(n_8),
.A2(n_47),
.B1(n_48),
.B2(n_56),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g43 ( 
.A1(n_9),
.A2(n_32),
.B1(n_33),
.B2(n_44),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_9),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_9),
.A2(n_44),
.B1(n_47),
.B2(n_48),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_9),
.A2(n_44),
.B1(n_75),
.B2(n_76),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_9),
.A2(n_29),
.B1(n_30),
.B2(n_44),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_10),
.A2(n_29),
.B1(n_30),
.B2(n_147),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_10),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_10),
.A2(n_75),
.B1(n_76),
.B2(n_147),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_SL g200 ( 
.A1(n_10),
.A2(n_32),
.B1(n_33),
.B2(n_147),
.Y(n_200)
);

AOI22xp33_ASAP7_75t_SL g233 ( 
.A1(n_10),
.A2(n_47),
.B1(n_48),
.B2(n_147),
.Y(n_233)
);

INVx11_ASAP7_75t_L g49 ( 
.A(n_11),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_12),
.A2(n_75),
.B1(n_76),
.B2(n_153),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_12),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_SL g179 ( 
.A1(n_12),
.A2(n_29),
.B1(n_30),
.B2(n_153),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_12),
.A2(n_32),
.B1(n_33),
.B2(n_153),
.Y(n_218)
);

AOI22xp33_ASAP7_75t_SL g241 ( 
.A1(n_12),
.A2(n_47),
.B1(n_48),
.B2(n_153),
.Y(n_241)
);

BUFx24_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_L g31 ( 
.A1(n_14),
.A2(n_32),
.B1(n_33),
.B2(n_35),
.Y(n_31)
);

INVx11_ASAP7_75t_SL g48 ( 
.A(n_15),
.Y(n_48)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_127),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_125),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_99),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_19),
.B(n_99),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g19 ( 
.A1(n_20),
.A2(n_21),
.B1(n_84),
.B2(n_85),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_23),
.B1(n_57),
.B2(n_58),
.Y(n_21)
);

CKINVDCx16_ASAP7_75t_R g22 ( 
.A(n_23),
.Y(n_22)
);

AOI21xp5_ASAP7_75t_L g104 ( 
.A1(n_23),
.A2(n_24),
.B(n_41),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_41),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_SL g24 ( 
.A1(n_25),
.A2(n_31),
.B1(n_36),
.B2(n_39),
.Y(n_24)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_25),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_25),
.B(n_68),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_25),
.A2(n_31),
.B1(n_146),
.B2(n_148),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_25),
.A2(n_31),
.B1(n_146),
.B2(n_179),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_25),
.A2(n_31),
.B1(n_179),
.B2(n_197),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_31),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_L g26 ( 
.A1(n_27),
.A2(n_28),
.B1(n_29),
.B2(n_30),
.Y(n_26)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_27),
.Y(n_35)
);

NAND2xp33_ASAP7_75t_SL g194 ( 
.A(n_27),
.B(n_33),
.Y(n_194)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_29),
.A2(n_30),
.B1(n_72),
.B2(n_73),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_29),
.B(n_72),
.Y(n_167)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_30),
.A2(n_79),
.B1(n_150),
.B2(n_167),
.Y(n_166)
);

AOI32xp33_ASAP7_75t_L g192 ( 
.A1(n_30),
.A2(n_32),
.A3(n_35),
.B1(n_193),
.B2(n_194),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_31),
.B(n_68),
.Y(n_67)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_31),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_31),
.B(n_164),
.Y(n_163)
);

OAI22xp33_ASAP7_75t_L g54 ( 
.A1(n_32),
.A2(n_33),
.B1(n_49),
.B2(n_50),
.Y(n_54)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

A2O1A1Ixp33_ASAP7_75t_L g219 ( 
.A1(n_33),
.A2(n_49),
.B(n_151),
.C(n_220),
.Y(n_219)
);

BUFx10_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_37),
.Y(n_36)
);

AOI21xp5_ASAP7_75t_L g116 ( 
.A1(n_37),
.A2(n_117),
.B(n_118),
.Y(n_116)
);

CKINVDCx16_ASAP7_75t_R g66 ( 
.A(n_39),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_42),
.B(n_51),
.Y(n_41)
);

OAI21xp5_ASAP7_75t_SL g210 ( 
.A1(n_42),
.A2(n_53),
.B(n_201),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_43),
.B(n_45),
.Y(n_42)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_43),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_45),
.B(n_55),
.Y(n_95)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_46),
.B(n_54),
.Y(n_53)
);

AOI21xp5_ASAP7_75t_L g61 ( 
.A1(n_46),
.A2(n_53),
.B(n_62),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_46),
.A2(n_53),
.B1(n_94),
.B2(n_115),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_L g134 ( 
.A1(n_46),
.A2(n_51),
.B(n_115),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_46),
.A2(n_53),
.B1(n_200),
.B2(n_201),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_46),
.A2(n_53),
.B1(n_217),
.B2(n_218),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_46),
.A2(n_53),
.B1(n_200),
.B2(n_218),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_SL g239 ( 
.A(n_46),
.B(n_151),
.Y(n_239)
);

OA22x2_ASAP7_75t_L g46 ( 
.A1(n_47),
.A2(n_48),
.B1(n_49),
.B2(n_50),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_47),
.B(n_88),
.Y(n_87)
);

INVx5_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g244 ( 
.A(n_48),
.B(n_245),
.Y(n_244)
);

INVx11_ASAP7_75t_L g50 ( 
.A(n_49),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_52),
.B(n_55),
.Y(n_51)
);

INVxp67_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

OAI21xp5_ASAP7_75t_SL g93 ( 
.A1(n_53),
.A2(n_94),
.B(n_95),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_SL g143 ( 
.A1(n_53),
.A2(n_62),
.B(n_95),
.Y(n_143)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_59),
.A2(n_69),
.B1(n_82),
.B2(n_83),
.Y(n_58)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_59),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_60),
.A2(n_61),
.B1(n_63),
.B2(n_64),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_61),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_64),
.Y(n_63)
);

AOI21xp5_ASAP7_75t_L g64 ( 
.A1(n_65),
.A2(n_66),
.B(n_67),
.Y(n_64)
);

AOI21xp5_ASAP7_75t_L g161 ( 
.A1(n_65),
.A2(n_162),
.B(n_163),
.Y(n_161)
);

AOI21xp5_ASAP7_75t_L g278 ( 
.A1(n_65),
.A2(n_67),
.B(n_279),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_69),
.Y(n_83)
);

OAI21xp5_ASAP7_75t_L g69 ( 
.A1(n_70),
.A2(n_74),
.B(n_77),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_70),
.B(n_81),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_70),
.A2(n_121),
.B1(n_158),
.B2(n_159),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_70),
.B(n_151),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_70),
.A2(n_121),
.B1(n_122),
.B2(n_159),
.Y(n_276)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

O2A1O1Ixp33_ASAP7_75t_L g78 ( 
.A1(n_71),
.A2(n_72),
.B(n_76),
.C(n_79),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_71),
.B(n_97),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_71),
.A2(n_78),
.B1(n_150),
.B2(n_152),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_72),
.B(n_76),
.Y(n_79)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx11_ASAP7_75t_L g76 ( 
.A(n_75),
.Y(n_76)
);

HAxp5_ASAP7_75t_SL g150 ( 
.A(n_76),
.B(n_151),
.CON(n_150),
.SN(n_150)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_78),
.B(n_80),
.Y(n_77)
);

AOI21xp5_ASAP7_75t_L g96 ( 
.A1(n_78),
.A2(n_97),
.B(n_98),
.Y(n_96)
);

CKINVDCx14_ASAP7_75t_R g121 ( 
.A(n_78),
.Y(n_121)
);

CKINVDCx16_ASAP7_75t_R g80 ( 
.A(n_81),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_85),
.Y(n_84)
);

AOI21xp5_ASAP7_75t_L g85 ( 
.A1(n_86),
.A2(n_92),
.B(n_96),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_86),
.B(n_93),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_86),
.A2(n_96),
.B1(n_102),
.B2(n_103),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_86),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g292 ( 
.A1(n_86),
.A2(n_93),
.B1(n_103),
.B2(n_293),
.Y(n_292)
);

AOI21xp5_ASAP7_75t_L g86 ( 
.A1(n_87),
.A2(n_89),
.B(n_90),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_87),
.B(n_111),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_L g135 ( 
.A1(n_87),
.A2(n_136),
.B(n_137),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_87),
.A2(n_89),
.B1(n_136),
.B2(n_169),
.Y(n_168)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_87),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_L g227 ( 
.A1(n_87),
.A2(n_112),
.B(n_228),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_87),
.A2(n_89),
.B1(n_233),
.B2(n_241),
.Y(n_240)
);

INVx11_ASAP7_75t_L g113 ( 
.A(n_88),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_88),
.B(n_151),
.Y(n_245)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_91),
.B(n_113),
.Y(n_112)
);

AOI21xp5_ASAP7_75t_L g190 ( 
.A1(n_91),
.A2(n_138),
.B(n_191),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g100 ( 
.A(n_92),
.B(n_101),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_93),
.Y(n_293)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_96),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_104),
.C(n_105),
.Y(n_99)
);

XOR2xp5_ASAP7_75t_L g300 ( 
.A(n_100),
.B(n_104),
.Y(n_300)
);

AOI22xp33_ASAP7_75t_SL g298 ( 
.A1(n_105),
.A2(n_106),
.B1(n_299),
.B2(n_300),
.Y(n_298)
);

CKINVDCx14_ASAP7_75t_R g105 ( 
.A(n_106),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_107),
.B(n_116),
.C(n_119),
.Y(n_106)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_107),
.B(n_289),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_114),
.Y(n_107)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_108),
.B(n_114),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_112),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_111),
.B(n_139),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_113),
.A2(n_191),
.B1(n_232),
.B2(n_234),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_116),
.A2(n_119),
.B1(n_120),
.B2(n_290),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_116),
.Y(n_290)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_SL g120 ( 
.A1(n_121),
.A2(n_122),
.B(n_124),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

AOI21xp5_ASAP7_75t_L g127 ( 
.A1(n_128),
.A2(n_296),
.B(n_301),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_SL g128 ( 
.A1(n_129),
.A2(n_283),
.B(n_295),
.Y(n_128)
);

O2A1O1Ixp33_ASAP7_75t_SL g129 ( 
.A1(n_130),
.A2(n_183),
.B(n_264),
.C(n_282),
.Y(n_129)
);

AND2x2_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_171),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_131),
.B(n_171),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_154),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_141),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_133),
.B(n_141),
.C(n_154),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_135),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_134),
.B(n_135),
.Y(n_273)
);

CKINVDCx16_ASAP7_75t_R g137 ( 
.A(n_138),
.Y(n_137)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_144),
.C(n_149),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_142),
.A2(n_143),
.B1(n_144),
.B2(n_145),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_143),
.Y(n_142)
);

CKINVDCx16_ASAP7_75t_R g144 ( 
.A(n_145),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g162 ( 
.A(n_148),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_SL g173 ( 
.A(n_149),
.B(n_174),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_152),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_SL g154 ( 
.A(n_155),
.B(n_165),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_156),
.A2(n_157),
.B1(n_160),
.B2(n_161),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_156),
.B(n_161),
.C(n_165),
.Y(n_280)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_161),
.Y(n_160)
);

CKINVDCx14_ASAP7_75t_R g279 ( 
.A(n_164),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_168),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g176 ( 
.A(n_166),
.B(n_168),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_175),
.C(n_177),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_172),
.A2(n_173),
.B1(n_259),
.B2(n_261),
.Y(n_258)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g259 ( 
.A1(n_175),
.A2(n_176),
.B1(n_177),
.B2(n_260),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_176),
.Y(n_175)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_177),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_180),
.C(n_181),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_SL g204 ( 
.A(n_178),
.B(n_205),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_180),
.A2(n_181),
.B1(n_182),
.B2(n_206),
.Y(n_205)
);

CKINVDCx14_ASAP7_75t_R g206 ( 
.A(n_180),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_182),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_SL g183 ( 
.A(n_184),
.B(n_263),
.Y(n_183)
);

AOI21xp5_ASAP7_75t_L g184 ( 
.A1(n_185),
.A2(n_256),
.B(n_262),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_L g185 ( 
.A1(n_186),
.A2(n_211),
.B(n_255),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_202),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g255 ( 
.A(n_187),
.B(n_202),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_188),
.B(n_195),
.C(n_198),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_188),
.A2(n_189),
.B1(n_252),
.B2(n_253),
.Y(n_251)
);

CKINVDCx16_ASAP7_75t_R g188 ( 
.A(n_189),
.Y(n_188)
);

XOR2xp5_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_192),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_190),
.B(n_192),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_L g253 ( 
.A1(n_195),
.A2(n_196),
.B1(n_198),
.B2(n_199),
.Y(n_253)
);

CKINVDCx16_ASAP7_75t_R g195 ( 
.A(n_196),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_199),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_203),
.A2(n_204),
.B1(n_207),
.B2(n_208),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_203),
.B(n_209),
.C(n_210),
.Y(n_257)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

CKINVDCx14_ASAP7_75t_R g207 ( 
.A(n_208),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_210),
.Y(n_208)
);

AOI21xp5_ASAP7_75t_L g211 ( 
.A1(n_212),
.A2(n_249),
.B(n_254),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_L g212 ( 
.A1(n_213),
.A2(n_229),
.B(n_248),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_221),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_214),
.B(n_221),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_SL g214 ( 
.A(n_215),
.B(n_219),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_215),
.A2(n_216),
.B1(n_219),
.B2(n_236),
.Y(n_235)
);

CKINVDCx16_ASAP7_75t_R g215 ( 
.A(n_216),
.Y(n_215)
);

CKINVDCx16_ASAP7_75t_R g236 ( 
.A(n_219),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_227),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_223),
.A2(n_224),
.B1(n_225),
.B2(n_226),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_223),
.B(n_226),
.C(n_227),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_224),
.Y(n_223)
);

CKINVDCx16_ASAP7_75t_R g225 ( 
.A(n_226),
.Y(n_225)
);

INVxp67_ASAP7_75t_L g234 ( 
.A(n_228),
.Y(n_234)
);

AOI21xp5_ASAP7_75t_L g229 ( 
.A1(n_230),
.A2(n_237),
.B(n_247),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_235),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_SL g247 ( 
.A(n_231),
.B(n_235),
.Y(n_247)
);

INVxp67_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

OAI21xp5_ASAP7_75t_SL g237 ( 
.A1(n_238),
.A2(n_242),
.B(n_246),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_240),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_239),
.B(n_240),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_243),
.B(n_244),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_251),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_SL g254 ( 
.A(n_250),
.B(n_251),
.Y(n_254)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_257),
.B(n_258),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_SL g262 ( 
.A(n_257),
.B(n_258),
.Y(n_262)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_259),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_266),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_SL g282 ( 
.A(n_265),
.B(n_266),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_267),
.A2(n_268),
.B1(n_280),
.B2(n_281),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_L g268 ( 
.A1(n_269),
.A2(n_270),
.B1(n_271),
.B2(n_272),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_269),
.B(n_272),
.C(n_281),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_270),
.Y(n_269)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_273),
.B(n_274),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_273),
.B(n_275),
.C(n_278),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_275),
.A2(n_276),
.B1(n_277),
.B2(n_278),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

CKINVDCx16_ASAP7_75t_R g277 ( 
.A(n_278),
.Y(n_277)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_280),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_284),
.B(n_285),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_SL g295 ( 
.A(n_284),
.B(n_285),
.Y(n_295)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_286),
.B(n_294),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_287),
.A2(n_288),
.B1(n_291),
.B2(n_292),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_287),
.B(n_292),
.C(n_294),
.Y(n_297)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_297),
.B(n_298),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_SL g301 ( 
.A(n_297),
.B(n_298),
.Y(n_301)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);


endmodule