module fake_jpeg_28174_n_169 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_169);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_169;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_9),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_8),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_10),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_4),
.Y(n_18)
);

INVx4_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_10),
.Y(n_23)
);

BUFx6f_ASAP7_75t_SL g24 ( 
.A(n_5),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_14),
.Y(n_26)
);

BUFx10_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_28),
.Y(n_31)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_31),
.Y(n_44)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_28),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_32),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_28),
.B(n_0),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_33),
.B(n_36),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_28),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_34),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_28),
.Y(n_35)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_24),
.Y(n_36)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_24),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_37),
.B(n_39),
.Y(n_51)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_27),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_38),
.B(n_40),
.Y(n_55)
);

CKINVDCx16_ASAP7_75t_R g39 ( 
.A(n_27),
.Y(n_39)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_27),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_SL g42 ( 
.A1(n_37),
.A2(n_19),
.B1(n_18),
.B2(n_26),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_42),
.A2(n_15),
.B1(n_23),
.B2(n_16),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g43 ( 
.A(n_33),
.B(n_18),
.Y(n_43)
);

OR2x2_ASAP7_75t_L g59 ( 
.A(n_43),
.B(n_23),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_39),
.B(n_21),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_45),
.B(n_54),
.Y(n_67)
);

OAI22xp33_ASAP7_75t_L g46 ( 
.A1(n_32),
.A2(n_19),
.B1(n_29),
.B2(n_27),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_46),
.A2(n_53),
.B1(n_25),
.B2(n_26),
.Y(n_68)
);

BUFx2_ASAP7_75t_L g49 ( 
.A(n_31),
.Y(n_49)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_49),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_34),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_50),
.B(n_52),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_32),
.B(n_17),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_36),
.A2(n_19),
.B1(n_20),
.B2(n_21),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_34),
.B(n_20),
.Y(n_54)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_57),
.B(n_58),
.Y(n_78)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g83 ( 
.A(n_59),
.B(n_64),
.Y(n_83)
);

AOI32xp33_ASAP7_75t_L g60 ( 
.A1(n_47),
.A2(n_40),
.A3(n_38),
.B1(n_27),
.B2(n_34),
.Y(n_60)
);

XNOR2xp5_ASAP7_75t_L g76 ( 
.A(n_60),
.B(n_68),
.Y(n_76)
);

OAI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_53),
.A2(n_40),
.B1(n_38),
.B2(n_17),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_61),
.A2(n_68),
.B1(n_70),
.B2(n_45),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_49),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_49),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_65),
.B(n_66),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_47),
.B(n_16),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_54),
.B(n_29),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_69),
.B(n_48),
.Y(n_77)
);

HB1xp67_ASAP7_75t_L g71 ( 
.A(n_41),
.Y(n_71)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_71),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_50),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_72),
.B(n_74),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_48),
.Y(n_73)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_73),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g74 ( 
.A(n_55),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_55),
.B(n_34),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_75),
.B(n_35),
.C(n_56),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_76),
.B(n_94),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_77),
.B(n_80),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_74),
.B(n_67),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_81),
.A2(n_75),
.B1(n_44),
.B2(n_22),
.Y(n_100)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_63),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_85),
.B(n_88),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_67),
.B(n_43),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_86),
.B(n_93),
.Y(n_104)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_60),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_69),
.A2(n_44),
.B1(n_51),
.B2(n_31),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_89),
.A2(n_81),
.B1(n_88),
.B2(n_93),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_72),
.B(n_15),
.Y(n_90)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_90),
.Y(n_106)
);

INVx8_ASAP7_75t_L g91 ( 
.A(n_57),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_91),
.A2(n_58),
.B1(n_44),
.B2(n_65),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_59),
.B(n_25),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_92),
.B(n_30),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_75),
.B(n_51),
.Y(n_93)
);

INVxp33_ASAP7_75t_L g96 ( 
.A(n_78),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_96),
.B(n_97),
.Y(n_114)
);

CKINVDCx16_ASAP7_75t_R g97 ( 
.A(n_87),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_98),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_100),
.B(n_107),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g115 ( 
.A(n_101),
.B(n_30),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_L g102 ( 
.A(n_80),
.B(n_62),
.Y(n_102)
);

XOR2xp5_ASAP7_75t_L g116 ( 
.A(n_102),
.B(n_84),
.Y(n_116)
);

INVx1_ASAP7_75t_SL g103 ( 
.A(n_79),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_103),
.B(n_105),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_76),
.A2(n_77),
.B1(n_94),
.B2(n_86),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_89),
.B(n_64),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_108),
.B(n_95),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_82),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_109),
.B(n_91),
.Y(n_121)
);

AOI221xp5_ASAP7_75t_L g112 ( 
.A1(n_107),
.A2(n_83),
.B1(n_85),
.B2(n_84),
.C(n_30),
.Y(n_112)
);

A2O1A1O1Ixp25_ASAP7_75t_L g133 ( 
.A1(n_112),
.A2(n_22),
.B(n_29),
.C(n_56),
.D(n_79),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_115),
.B(n_122),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_116),
.B(n_119),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_L g118 ( 
.A1(n_110),
.A2(n_83),
.B(n_62),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g136 ( 
.A(n_118),
.Y(n_136)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_95),
.Y(n_119)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_120),
.Y(n_127)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_121),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_106),
.B(n_13),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_102),
.B(n_91),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_123),
.B(n_124),
.Y(n_135)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_103),
.Y(n_124)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_108),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_125),
.A2(n_110),
.B1(n_104),
.B2(n_96),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_113),
.A2(n_105),
.B1(n_100),
.B2(n_99),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_126),
.A2(n_111),
.B1(n_22),
.B2(n_2),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_128),
.A2(n_133),
.B1(n_111),
.B2(n_124),
.Y(n_140)
);

NOR2x1_ASAP7_75t_L g129 ( 
.A(n_125),
.B(n_104),
.Y(n_129)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_129),
.Y(n_138)
);

MAJx2_ASAP7_75t_L g131 ( 
.A(n_116),
.B(n_110),
.C(n_35),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_131),
.B(n_132),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_123),
.B(n_56),
.C(n_73),
.Y(n_132)
);

AOI321xp33_ASAP7_75t_L g139 ( 
.A1(n_127),
.A2(n_118),
.A3(n_119),
.B1(n_117),
.B2(n_114),
.C(n_113),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g150 ( 
.A(n_139),
.B(n_130),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_140),
.B(n_142),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g141 ( 
.A(n_137),
.B(n_120),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_141),
.B(n_144),
.C(n_132),
.Y(n_147)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_135),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_143),
.B(n_1),
.Y(n_152)
);

XOR2xp5_ASAP7_75t_L g144 ( 
.A(n_131),
.B(n_0),
.Y(n_144)
);

XNOR2x1_ASAP7_75t_L g146 ( 
.A(n_128),
.B(n_0),
.Y(n_146)
);

AOI21xp5_ASAP7_75t_L g149 ( 
.A1(n_146),
.A2(n_1),
.B(n_2),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_SL g155 ( 
.A(n_147),
.B(n_145),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_138),
.A2(n_126),
.B1(n_129),
.B2(n_136),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_148),
.B(n_152),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_L g154 ( 
.A1(n_149),
.A2(n_134),
.B(n_136),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_SL g158 ( 
.A(n_150),
.B(n_153),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_146),
.Y(n_153)
);

AO21x1_ASAP7_75t_L g160 ( 
.A1(n_154),
.A2(n_151),
.B(n_133),
.Y(n_160)
);

AOI31xp33_ASAP7_75t_L g162 ( 
.A1(n_155),
.A2(n_1),
.A3(n_3),
.B(n_4),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_147),
.B(n_144),
.C(n_141),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_156),
.B(n_148),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_159),
.B(n_162),
.C(n_157),
.Y(n_163)
);

AOI21xp5_ASAP7_75t_SL g165 ( 
.A1(n_160),
.A2(n_161),
.B(n_5),
.Y(n_165)
);

A2O1A1Ixp33_ASAP7_75t_SL g161 ( 
.A1(n_158),
.A2(n_157),
.B(n_2),
.C(n_3),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_SL g166 ( 
.A1(n_163),
.A2(n_164),
.B(n_5),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_SL g164 ( 
.A(n_159),
.B(n_4),
.Y(n_164)
);

AOI21xp5_ASAP7_75t_SL g167 ( 
.A1(n_165),
.A2(n_6),
.B(n_7),
.Y(n_167)
);

O2A1O1Ixp33_ASAP7_75t_L g168 ( 
.A1(n_166),
.A2(n_167),
.B(n_6),
.C(n_7),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_168),
.B(n_6),
.Y(n_169)
);


endmodule