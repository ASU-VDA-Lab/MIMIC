module fake_jpeg_8468_n_62 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_62);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_62;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_23;
wire n_10;
wire n_27;
wire n_55;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_59;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_56;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_15;

INVx1_ASAP7_75t_L g9 ( 
.A(n_6),
.Y(n_9)
);

INVx2_ASAP7_75t_L g10 ( 
.A(n_0),
.Y(n_10)
);

INVx4_ASAP7_75t_L g11 ( 
.A(n_6),
.Y(n_11)
);

BUFx3_ASAP7_75t_L g12 ( 
.A(n_8),
.Y(n_12)
);

BUFx5_ASAP7_75t_L g13 ( 
.A(n_8),
.Y(n_13)
);

BUFx12f_ASAP7_75t_L g14 ( 
.A(n_7),
.Y(n_14)
);

INVx2_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_4),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_17),
.B(n_9),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_SL g24 ( 
.A(n_18),
.B(n_23),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

INVx1_ASAP7_75t_SL g26 ( 
.A(n_19),
.Y(n_26)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_20),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_21),
.Y(n_27)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_22),
.B(n_15),
.Y(n_29)
);

OR2x2_ASAP7_75t_SL g23 ( 
.A(n_17),
.B(n_0),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_SL g25 ( 
.A(n_22),
.B(n_10),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_SL g30 ( 
.A(n_25),
.B(n_15),
.Y(n_30)
);

OAI21xp5_ASAP7_75t_SL g31 ( 
.A1(n_29),
.A2(n_23),
.B(n_10),
.Y(n_31)
);

OAI21xp5_ASAP7_75t_L g41 ( 
.A1(n_30),
.A2(n_35),
.B(n_12),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g44 ( 
.A(n_31),
.B(n_16),
.Y(n_44)
);

AND2x2_ASAP7_75t_SL g32 ( 
.A(n_29),
.B(n_19),
.Y(n_32)
);

MAJIxp5_ASAP7_75t_L g43 ( 
.A(n_32),
.B(n_16),
.C(n_2),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_26),
.Y(n_33)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_33),
.Y(n_39)
);

O2A1O1Ixp33_ASAP7_75t_L g34 ( 
.A1(n_24),
.A2(n_21),
.B(n_20),
.C(n_11),
.Y(n_34)
);

AOI22xp5_ASAP7_75t_SL g38 ( 
.A1(n_34),
.A2(n_27),
.B1(n_26),
.B2(n_14),
.Y(n_38)
);

AOI21xp5_ASAP7_75t_L g35 ( 
.A1(n_28),
.A2(n_11),
.B(n_12),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_27),
.B(n_14),
.Y(n_36)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_36),
.Y(n_42)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_37),
.B(n_14),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_38),
.A2(n_44),
.B1(n_39),
.B2(n_2),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_40),
.B(n_1),
.Y(n_47)
);

XNOR2xp5_ASAP7_75t_L g48 ( 
.A(n_41),
.B(n_7),
.Y(n_48)
);

MAJIxp5_ASAP7_75t_L g45 ( 
.A(n_43),
.B(n_32),
.C(n_34),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_45),
.B(n_46),
.Y(n_51)
);

MAJIxp5_ASAP7_75t_L g46 ( 
.A(n_42),
.B(n_32),
.C(n_33),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_47),
.B(n_49),
.Y(n_52)
);

OAI21x1_ASAP7_75t_L g54 ( 
.A1(n_48),
.A2(n_50),
.B(n_1),
.Y(n_54)
);

MAJIxp5_ASAP7_75t_L g49 ( 
.A(n_43),
.B(n_1),
.C(n_2),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_47),
.B(n_38),
.Y(n_53)
);

XNOR2xp5_ASAP7_75t_L g55 ( 
.A(n_53),
.B(n_54),
.Y(n_55)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_51),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_56),
.B(n_57),
.Y(n_58)
);

AOI221xp5_ASAP7_75t_L g57 ( 
.A1(n_52),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.C(n_6),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g59 ( 
.A(n_55),
.B(n_57),
.C(n_4),
.Y(n_59)
);

HB1xp67_ASAP7_75t_L g60 ( 
.A(n_59),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_60),
.A2(n_58),
.B1(n_3),
.B2(n_5),
.Y(n_61)
);

XNOR2xp5_ASAP7_75t_L g62 ( 
.A(n_61),
.B(n_3),
.Y(n_62)
);


endmodule