module fake_jpeg_11483_n_387 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_387);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_387;

wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_19;
wire n_182;
wire n_385;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx8_ASAP7_75t_L g15 ( 
.A(n_9),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_6),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_1),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

INVxp67_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

INVx1_ASAP7_75t_SL g23 ( 
.A(n_9),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_7),
.B(n_5),
.Y(n_24)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_2),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_8),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_12),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_11),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_4),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_3),
.Y(n_39)
);

BUFx10_ASAP7_75t_L g40 ( 
.A(n_6),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_2),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_4),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_24),
.B(n_14),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_43),
.B(n_51),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_18),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_44),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_18),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_45),
.Y(n_119)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

INVx5_ASAP7_75t_L g120 ( 
.A(n_46),
.Y(n_120)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_22),
.Y(n_47)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_47),
.Y(n_86)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_22),
.Y(n_48)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_48),
.Y(n_116)
);

INVx6_ASAP7_75t_SL g49 ( 
.A(n_40),
.Y(n_49)
);

CKINVDCx6p67_ASAP7_75t_R g112 ( 
.A(n_49),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_18),
.Y(n_50)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_50),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_31),
.B(n_14),
.Y(n_51)
);

INVx6_ASAP7_75t_SL g52 ( 
.A(n_40),
.Y(n_52)
);

CKINVDCx14_ASAP7_75t_R g88 ( 
.A(n_52),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_15),
.Y(n_53)
);

INVx8_ASAP7_75t_L g130 ( 
.A(n_53),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_31),
.B(n_13),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_54),
.B(n_80),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_40),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_55),
.B(n_56),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_40),
.Y(n_56)
);

INVx11_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

CKINVDCx16_ASAP7_75t_R g103 ( 
.A(n_57),
.Y(n_103)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_25),
.Y(n_58)
);

INVx2_ASAP7_75t_SL g89 ( 
.A(n_58),
.Y(n_89)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_15),
.Y(n_59)
);

INVx5_ASAP7_75t_L g123 ( 
.A(n_59),
.Y(n_123)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_25),
.Y(n_60)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_60),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_35),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_61),
.B(n_72),
.Y(n_98)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_36),
.Y(n_62)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_62),
.Y(n_115)
);

INVx11_ASAP7_75t_L g63 ( 
.A(n_15),
.Y(n_63)
);

CKINVDCx14_ASAP7_75t_R g133 ( 
.A(n_63),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_30),
.Y(n_64)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_64),
.Y(n_127)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_26),
.Y(n_65)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_65),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_30),
.Y(n_66)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_66),
.Y(n_90)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_26),
.Y(n_67)
);

HB1xp67_ASAP7_75t_L g94 ( 
.A(n_67),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_30),
.Y(n_68)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_68),
.Y(n_111)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_26),
.Y(n_69)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_69),
.Y(n_118)
);

BUFx12f_ASAP7_75t_L g70 ( 
.A(n_16),
.Y(n_70)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_70),
.Y(n_124)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_32),
.Y(n_71)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_71),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g72 ( 
.A(n_16),
.B(n_12),
.Y(n_72)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_32),
.Y(n_73)
);

HB1xp67_ASAP7_75t_L g106 ( 
.A(n_73),
.Y(n_106)
);

BUFx12f_ASAP7_75t_L g74 ( 
.A(n_17),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_74),
.B(n_77),
.Y(n_102)
);

INVx6_ASAP7_75t_SL g75 ( 
.A(n_20),
.Y(n_75)
);

NAND2xp33_ASAP7_75t_SL g107 ( 
.A(n_75),
.B(n_76),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_26),
.Y(n_76)
);

CKINVDCx16_ASAP7_75t_R g77 ( 
.A(n_33),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_33),
.Y(n_78)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_78),
.B(n_79),
.Y(n_93)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_33),
.Y(n_79)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_33),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_35),
.B(n_12),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_81),
.B(n_11),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_39),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_82),
.B(n_83),
.Y(n_109)
);

INVx5_ASAP7_75t_L g83 ( 
.A(n_39),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_47),
.A2(n_73),
.B1(n_71),
.B2(n_48),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_85),
.A2(n_105),
.B1(n_122),
.B2(n_74),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_82),
.B(n_37),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_87),
.B(n_92),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_59),
.A2(n_23),
.B1(n_37),
.B2(n_27),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g165 ( 
.A1(n_91),
.A2(n_101),
.B1(n_117),
.B2(n_125),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_83),
.B(n_23),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_64),
.A2(n_68),
.B1(n_66),
.B2(n_44),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_95),
.A2(n_99),
.B1(n_108),
.B2(n_113),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_L g99 ( 
.A1(n_45),
.A2(n_42),
.B1(n_41),
.B2(n_38),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_46),
.A2(n_19),
.B1(n_21),
.B2(n_27),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_50),
.A2(n_42),
.B1(n_41),
.B2(n_38),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_53),
.A2(n_34),
.B1(n_28),
.B2(n_17),
.Y(n_108)
);

NAND3xp33_ASAP7_75t_L g150 ( 
.A(n_110),
.B(n_5),
.C(n_6),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_L g113 ( 
.A1(n_58),
.A2(n_34),
.B1(n_28),
.B2(n_29),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_60),
.A2(n_29),
.B1(n_21),
.B2(n_19),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_114),
.B(n_132),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_49),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_117)
);

OAI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_63),
.A2(n_11),
.B1(n_2),
.B2(n_3),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_52),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_70),
.B(n_1),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_126),
.B(n_131),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_70),
.B(n_4),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_67),
.A2(n_5),
.B1(n_6),
.B2(n_8),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_104),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g184 ( 
.A(n_134),
.Y(n_184)
);

INVx6_ASAP7_75t_L g135 ( 
.A(n_104),
.Y(n_135)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_135),
.Y(n_202)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_100),
.Y(n_137)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_137),
.Y(n_214)
);

CKINVDCx16_ASAP7_75t_R g138 ( 
.A(n_102),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_138),
.B(n_150),
.Y(n_182)
);

AND2x4_ASAP7_75t_L g139 ( 
.A(n_92),
.B(n_75),
.Y(n_139)
);

CKINVDCx16_ASAP7_75t_R g194 ( 
.A(n_139),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_140),
.A2(n_165),
.B1(n_179),
.B2(n_153),
.Y(n_222)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_97),
.Y(n_141)
);

INVx2_ASAP7_75t_SL g192 ( 
.A(n_141),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_98),
.B(n_74),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_SL g210 ( 
.A(n_142),
.B(n_147),
.Y(n_210)
);

INVx13_ASAP7_75t_L g143 ( 
.A(n_112),
.Y(n_143)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_143),
.Y(n_183)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_106),
.Y(n_145)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_145),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_121),
.B(n_80),
.Y(n_147)
);

CKINVDCx6p67_ASAP7_75t_R g148 ( 
.A(n_112),
.Y(n_148)
);

INVx13_ASAP7_75t_L g198 ( 
.A(n_148),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_129),
.B(n_79),
.Y(n_149)
);

INVxp67_ASAP7_75t_L g193 ( 
.A(n_149),
.Y(n_193)
);

INVx5_ASAP7_75t_L g151 ( 
.A(n_130),
.Y(n_151)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_151),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_112),
.B(n_65),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_152),
.B(n_154),
.Y(n_200)
);

INVx8_ASAP7_75t_L g153 ( 
.A(n_119),
.Y(n_153)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_153),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_SL g154 ( 
.A(n_126),
.B(n_62),
.Y(n_154)
);

INVx4_ASAP7_75t_L g156 ( 
.A(n_128),
.Y(n_156)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_156),
.Y(n_201)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_118),
.Y(n_157)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_157),
.Y(n_203)
);

INVxp67_ASAP7_75t_L g158 ( 
.A(n_94),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_158),
.B(n_164),
.Y(n_207)
);

AOI21xp33_ASAP7_75t_L g159 ( 
.A1(n_131),
.A2(n_57),
.B(n_62),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_R g188 ( 
.A(n_159),
.B(n_93),
.Y(n_188)
);

BUFx6f_ASAP7_75t_L g160 ( 
.A(n_119),
.Y(n_160)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_160),
.Y(n_204)
);

INVx6_ASAP7_75t_L g161 ( 
.A(n_84),
.Y(n_161)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_161),
.Y(n_205)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_84),
.Y(n_162)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_162),
.Y(n_206)
);

BUFx4f_ASAP7_75t_SL g163 ( 
.A(n_112),
.Y(n_163)
);

INVx13_ASAP7_75t_L g208 ( 
.A(n_163),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_88),
.B(n_76),
.Y(n_164)
);

INVx11_ASAP7_75t_L g166 ( 
.A(n_133),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_166),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_SL g167 ( 
.A(n_124),
.B(n_78),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_167),
.B(n_169),
.Y(n_219)
);

INVx4_ASAP7_75t_L g168 ( 
.A(n_128),
.Y(n_168)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_168),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_124),
.B(n_69),
.Y(n_169)
);

INVx2_ASAP7_75t_SL g170 ( 
.A(n_118),
.Y(n_170)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_170),
.Y(n_220)
);

AND2x4_ASAP7_75t_L g171 ( 
.A(n_87),
.B(n_9),
.Y(n_171)
);

AND2x2_ASAP7_75t_L g215 ( 
.A(n_171),
.B(n_176),
.Y(n_215)
);

INVx6_ASAP7_75t_L g172 ( 
.A(n_127),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_SL g209 ( 
.A1(n_172),
.A2(n_175),
.B1(n_177),
.B2(n_178),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_86),
.B(n_10),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_173),
.B(n_181),
.Y(n_186)
);

INVx13_ASAP7_75t_L g174 ( 
.A(n_107),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_174),
.Y(n_211)
);

INVx6_ASAP7_75t_L g175 ( 
.A(n_127),
.Y(n_175)
);

BUFx3_ASAP7_75t_L g176 ( 
.A(n_115),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_SL g177 ( 
.A1(n_105),
.A2(n_10),
.B1(n_107),
.B2(n_130),
.Y(n_177)
);

BUFx3_ASAP7_75t_L g178 ( 
.A(n_115),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_SL g179 ( 
.A1(n_120),
.A2(n_10),
.B1(n_123),
.B2(n_96),
.Y(n_179)
);

AOI21xp5_ASAP7_75t_L g199 ( 
.A1(n_179),
.A2(n_120),
.B(n_89),
.Y(n_199)
);

INVx5_ASAP7_75t_L g180 ( 
.A(n_123),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_180),
.A2(n_89),
.B1(n_93),
.B2(n_96),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_86),
.B(n_10),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_L g187 ( 
.A1(n_139),
.A2(n_109),
.B(n_89),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_SL g232 ( 
.A1(n_187),
.A2(n_188),
.B(n_199),
.Y(n_232)
);

OAI21xp5_ASAP7_75t_SL g189 ( 
.A1(n_174),
.A2(n_114),
.B(n_132),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_189),
.B(n_134),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_146),
.A2(n_90),
.B1(n_111),
.B2(n_116),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_195),
.A2(n_222),
.B1(n_158),
.B2(n_135),
.Y(n_235)
);

FAx1_ASAP7_75t_SL g196 ( 
.A(n_136),
.B(n_85),
.CI(n_116),
.CON(n_196),
.SN(n_196)
);

NOR2xp33_ASAP7_75t_SL g231 ( 
.A(n_196),
.B(n_163),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_144),
.B(n_90),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_212),
.B(n_213),
.Y(n_230)
);

A2O1A1Ixp33_ASAP7_75t_L g213 ( 
.A1(n_139),
.A2(n_93),
.B(n_111),
.C(n_103),
.Y(n_213)
);

CKINVDCx16_ASAP7_75t_R g227 ( 
.A(n_216),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_155),
.A2(n_171),
.B1(n_139),
.B2(n_177),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_217),
.A2(n_165),
.B1(n_171),
.B2(n_151),
.Y(n_226)
);

AND2x6_ASAP7_75t_L g221 ( 
.A(n_166),
.B(n_171),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_221),
.B(n_148),
.Y(n_223)
);

INVxp67_ASAP7_75t_L g275 ( 
.A(n_223),
.Y(n_275)
);

INVx5_ASAP7_75t_L g224 ( 
.A(n_183),
.Y(n_224)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_224),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_210),
.B(n_148),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_225),
.B(n_231),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_226),
.A2(n_215),
.B1(n_213),
.B2(n_221),
.Y(n_262)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_220),
.Y(n_228)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_228),
.Y(n_260)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_220),
.Y(n_229)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_229),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_212),
.B(n_170),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_233),
.B(n_236),
.Y(n_269)
);

INVx3_ASAP7_75t_SL g234 ( 
.A(n_183),
.Y(n_234)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_234),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_L g272 ( 
.A1(n_235),
.A2(n_243),
.B1(n_255),
.B2(n_256),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_211),
.B(n_168),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_203),
.Y(n_237)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_237),
.Y(n_266)
);

INVx3_ASAP7_75t_L g238 ( 
.A(n_202),
.Y(n_238)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_238),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_211),
.B(n_156),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_239),
.B(n_245),
.Y(n_271)
);

CKINVDCx14_ASAP7_75t_R g240 ( 
.A(n_208),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_240),
.B(n_241),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_SL g241 ( 
.A(n_193),
.B(n_163),
.Y(n_241)
);

AOI22x1_ASAP7_75t_SL g242 ( 
.A1(n_188),
.A2(n_178),
.B1(n_176),
.B2(n_143),
.Y(n_242)
);

OAI21xp5_ASAP7_75t_SL g280 ( 
.A1(n_242),
.A2(n_253),
.B(n_254),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_222),
.A2(n_161),
.B1(n_172),
.B2(n_175),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_210),
.B(n_180),
.Y(n_244)
);

INVxp67_ASAP7_75t_L g282 ( 
.A(n_244),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_215),
.B(n_162),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_246),
.B(n_216),
.Y(n_274)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_205),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_247),
.Y(n_264)
);

OAI21xp5_ASAP7_75t_SL g248 ( 
.A1(n_194),
.A2(n_160),
.B(n_217),
.Y(n_248)
);

AOI21xp5_ASAP7_75t_L g257 ( 
.A1(n_248),
.A2(n_199),
.B(n_187),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_219),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_249),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_207),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_250),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_SL g251 ( 
.A(n_193),
.B(n_200),
.Y(n_251)
);

OAI21xp5_ASAP7_75t_L g268 ( 
.A1(n_251),
.A2(n_192),
.B(n_185),
.Y(n_268)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_203),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_252),
.Y(n_276)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_190),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_190),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_SL g255 ( 
.A(n_192),
.B(n_186),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_195),
.A2(n_189),
.B1(n_215),
.B2(n_194),
.Y(n_256)
);

AOI21xp5_ASAP7_75t_L g292 ( 
.A1(n_257),
.A2(n_277),
.B(n_280),
.Y(n_292)
);

OAI22x1_ASAP7_75t_L g304 ( 
.A1(n_262),
.A2(n_253),
.B1(n_254),
.B2(n_247),
.Y(n_304)
);

OAI32xp33_ASAP7_75t_L g267 ( 
.A1(n_230),
.A2(n_196),
.A3(n_186),
.B1(n_182),
.B2(n_205),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_267),
.B(n_283),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_268),
.B(n_191),
.Y(n_306)
);

A2O1A1Ixp33_ASAP7_75t_SL g270 ( 
.A1(n_232),
.A2(n_209),
.B(n_208),
.C(n_196),
.Y(n_270)
);

AO22x1_ASAP7_75t_L g300 ( 
.A1(n_270),
.A2(n_234),
.B1(n_241),
.B2(n_224),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_274),
.B(n_233),
.C(n_249),
.Y(n_301)
);

AOI21xp5_ASAP7_75t_L g277 ( 
.A1(n_232),
.A2(n_185),
.B(n_201),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_256),
.A2(n_192),
.B1(n_206),
.B2(n_204),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_281),
.A2(n_285),
.B1(n_252),
.B2(n_237),
.Y(n_297)
);

OA21x2_ASAP7_75t_L g283 ( 
.A1(n_236),
.A2(n_218),
.B(n_201),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_226),
.A2(n_227),
.B1(n_231),
.B2(n_230),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_284),
.A2(n_238),
.B1(n_202),
.B2(n_214),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_L g285 ( 
.A1(n_235),
.A2(n_206),
.B1(n_197),
.B2(n_204),
.Y(n_285)
);

OA22x2_ASAP7_75t_L g286 ( 
.A1(n_243),
.A2(n_191),
.B1(n_197),
.B2(n_218),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_286),
.B(n_239),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_261),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_287),
.B(n_291),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_L g288 ( 
.A1(n_262),
.A2(n_227),
.B1(n_242),
.B2(n_246),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_288),
.A2(n_296),
.B1(n_302),
.B2(n_307),
.Y(n_316)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_260),
.Y(n_289)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_289),
.Y(n_311)
);

INVx1_ASAP7_75t_SL g291 ( 
.A(n_265),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_292),
.B(n_295),
.Y(n_319)
);

CKINVDCx14_ASAP7_75t_R g293 ( 
.A(n_259),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_293),
.B(n_308),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_273),
.B(n_251),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_SL g321 ( 
.A(n_294),
.B(n_304),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_271),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_L g296 ( 
.A1(n_257),
.A2(n_284),
.B1(n_273),
.B2(n_275),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_L g312 ( 
.A1(n_297),
.A2(n_299),
.B1(n_303),
.B2(n_269),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_298),
.B(n_305),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_272),
.A2(n_248),
.B1(n_250),
.B2(n_245),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_SL g330 ( 
.A(n_300),
.B(n_306),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_301),
.B(n_270),
.C(n_263),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_L g302 ( 
.A1(n_275),
.A2(n_234),
.B1(n_229),
.B2(n_228),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_281),
.A2(n_274),
.B1(n_282),
.B2(n_271),
.Y(n_303)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_260),
.Y(n_305)
);

INVx8_ASAP7_75t_L g308 ( 
.A(n_258),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_269),
.B(n_214),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_309),
.B(n_276),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_279),
.B(n_184),
.Y(n_310)
);

OAI322xp33_ASAP7_75t_L g325 ( 
.A1(n_310),
.A2(n_265),
.A3(n_198),
.B1(n_278),
.B2(n_270),
.C1(n_266),
.C2(n_283),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_L g341 ( 
.A1(n_312),
.A2(n_302),
.B1(n_304),
.B2(n_305),
.Y(n_341)
);

AOI322xp5_ASAP7_75t_L g314 ( 
.A1(n_296),
.A2(n_282),
.A3(n_280),
.B1(n_267),
.B2(n_270),
.C1(n_276),
.C2(n_277),
.Y(n_314)
);

AO21x1_ASAP7_75t_L g336 ( 
.A1(n_314),
.A2(n_321),
.B(n_320),
.Y(n_336)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_301),
.B(n_268),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_315),
.B(n_324),
.C(n_327),
.Y(n_338)
);

XNOR2xp5_ASAP7_75t_L g337 ( 
.A(n_318),
.B(n_328),
.Y(n_337)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_322),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_287),
.B(n_258),
.Y(n_323)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_323),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_303),
.B(n_270),
.C(n_263),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_SL g335 ( 
.A1(n_325),
.A2(n_329),
.B1(n_291),
.B2(n_307),
.Y(n_335)
);

AOI22xp5_ASAP7_75t_L g326 ( 
.A1(n_288),
.A2(n_283),
.B1(n_266),
.B2(n_264),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_L g331 ( 
.A1(n_326),
.A2(n_297),
.B1(n_298),
.B2(n_306),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_299),
.B(n_264),
.C(n_278),
.Y(n_327)
);

XOR2xp5_ASAP7_75t_L g328 ( 
.A(n_290),
.B(n_286),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_290),
.B(n_286),
.C(n_184),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_L g359 ( 
.A1(n_331),
.A2(n_311),
.B1(n_308),
.B2(n_286),
.Y(n_359)
);

OAI22xp5_ASAP7_75t_L g334 ( 
.A1(n_316),
.A2(n_295),
.B1(n_310),
.B2(n_309),
.Y(n_334)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_334),
.Y(n_348)
);

OAI22xp5_ASAP7_75t_SL g350 ( 
.A1(n_335),
.A2(n_336),
.B1(n_341),
.B2(n_316),
.Y(n_350)
);

CKINVDCx20_ASAP7_75t_R g339 ( 
.A(n_313),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g356 ( 
.A(n_339),
.B(n_342),
.Y(n_356)
);

XOR2xp5_ASAP7_75t_SL g340 ( 
.A(n_315),
.B(n_292),
.Y(n_340)
);

XOR2xp5_ASAP7_75t_L g351 ( 
.A(n_340),
.B(n_318),
.Y(n_351)
);

BUFx12_ASAP7_75t_L g342 ( 
.A(n_319),
.Y(n_342)
);

AND2x2_ASAP7_75t_L g343 ( 
.A(n_313),
.B(n_308),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_343),
.B(n_346),
.Y(n_349)
);

BUFx12_ASAP7_75t_L g344 ( 
.A(n_319),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_344),
.B(n_328),
.Y(n_357)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_320),
.Y(n_345)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_345),
.Y(n_353)
);

OAI21xp5_ASAP7_75t_L g346 ( 
.A1(n_330),
.A2(n_300),
.B(n_289),
.Y(n_346)
);

OAI21xp5_ASAP7_75t_SL g347 ( 
.A1(n_335),
.A2(n_300),
.B(n_324),
.Y(n_347)
);

OR2x2_ASAP7_75t_L g360 ( 
.A(n_347),
.B(n_354),
.Y(n_360)
);

AOI22xp5_ASAP7_75t_L g364 ( 
.A1(n_350),
.A2(n_346),
.B1(n_332),
.B2(n_345),
.Y(n_364)
);

AOI21xp5_ASAP7_75t_L g367 ( 
.A1(n_351),
.A2(n_338),
.B(n_352),
.Y(n_367)
);

XOR2xp5_ASAP7_75t_L g352 ( 
.A(n_337),
.B(n_327),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_L g366 ( 
.A(n_352),
.B(n_338),
.Y(n_366)
);

OAI21xp5_ASAP7_75t_SL g354 ( 
.A1(n_342),
.A2(n_329),
.B(n_326),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_343),
.B(n_322),
.Y(n_355)
);

OAI21x1_ASAP7_75t_SL g365 ( 
.A1(n_355),
.A2(n_343),
.B(n_344),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_357),
.B(n_358),
.Y(n_362)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_333),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_359),
.B(n_341),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_SL g361 ( 
.A(n_356),
.B(n_317),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_SL g373 ( 
.A(n_361),
.B(n_364),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_363),
.B(n_366),
.Y(n_370)
);

AOI21xp5_ASAP7_75t_L g369 ( 
.A1(n_365),
.A2(n_367),
.B(n_368),
.Y(n_369)
);

OAI21xp5_ASAP7_75t_L g368 ( 
.A1(n_349),
.A2(n_342),
.B(n_344),
.Y(n_368)
);

OAI21xp5_ASAP7_75t_SL g371 ( 
.A1(n_360),
.A2(n_349),
.B(n_355),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_371),
.B(n_372),
.Y(n_379)
);

OAI21xp5_ASAP7_75t_L g372 ( 
.A1(n_360),
.A2(n_347),
.B(n_354),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_L g374 ( 
.A(n_362),
.B(n_348),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_L g376 ( 
.A(n_374),
.B(n_375),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_L g375 ( 
.A(n_364),
.B(n_350),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_L g377 ( 
.A(n_370),
.B(n_359),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_377),
.B(n_378),
.Y(n_382)
);

XOR2xp5_ASAP7_75t_L g378 ( 
.A(n_369),
.B(n_337),
.Y(n_378)
);

AOI22xp5_ASAP7_75t_L g380 ( 
.A1(n_379),
.A2(n_372),
.B1(n_353),
.B2(n_368),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_380),
.B(n_381),
.Y(n_384)
);

OAI22xp5_ASAP7_75t_L g381 ( 
.A1(n_376),
.A2(n_373),
.B1(n_336),
.B2(n_378),
.Y(n_381)
);

NAND3xp33_ASAP7_75t_L g383 ( 
.A(n_382),
.B(n_340),
.C(n_351),
.Y(n_383)
);

OAI21x1_ASAP7_75t_L g385 ( 
.A1(n_383),
.A2(n_380),
.B(n_198),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_385),
.B(n_384),
.Y(n_386)
);

XNOR2x2_ASAP7_75t_SL g387 ( 
.A(n_386),
.B(n_184),
.Y(n_387)
);


endmodule