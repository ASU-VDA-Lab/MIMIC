module fake_aes_839_n_666 (n_53, n_67, n_45, n_20, n_2, n_38, n_44, n_64, n_54, n_62, n_36, n_47, n_37, n_69, n_34, n_5, n_23, n_8, n_28, n_31, n_22, n_46, n_48, n_58, n_57, n_11, n_25, n_16, n_26, n_13, n_30, n_33, n_50, n_52, n_49, n_59, n_73, n_3, n_18, n_60, n_66, n_32, n_0, n_41, n_1, n_35, n_55, n_65, n_12, n_9, n_70, n_17, n_63, n_14, n_10, n_15, n_56, n_71, n_42, n_24, n_19, n_61, n_21, n_6, n_4, n_74, n_72, n_51, n_29, n_43, n_7, n_68, n_40, n_27, n_39, n_666);
input n_53;
input n_67;
input n_45;
input n_20;
input n_2;
input n_38;
input n_44;
input n_64;
input n_54;
input n_62;
input n_36;
input n_47;
input n_37;
input n_69;
input n_34;
input n_5;
input n_23;
input n_8;
input n_28;
input n_31;
input n_22;
input n_46;
input n_48;
input n_58;
input n_57;
input n_11;
input n_25;
input n_16;
input n_26;
input n_13;
input n_30;
input n_33;
input n_50;
input n_52;
input n_49;
input n_59;
input n_73;
input n_3;
input n_18;
input n_60;
input n_66;
input n_32;
input n_0;
input n_41;
input n_1;
input n_35;
input n_55;
input n_65;
input n_12;
input n_9;
input n_70;
input n_17;
input n_63;
input n_14;
input n_10;
input n_15;
input n_56;
input n_71;
input n_42;
input n_24;
input n_19;
input n_61;
input n_21;
input n_6;
input n_4;
input n_74;
input n_72;
input n_51;
input n_29;
input n_43;
input n_7;
input n_68;
input n_40;
input n_27;
input n_39;
output n_666;
wire n_117;
wire n_663;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_383;
wire n_288;
wire n_661;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_642;
wire n_586;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_647;
wire n_367;
wire n_644;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_108;
wire n_91;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_307;
wire n_191;
wire n_634;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_77;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_90;
wire n_357;
wire n_653;
wire n_260;
wire n_78;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_75;
wire n_376;
wire n_639;
wire n_552;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_76;
wire n_520;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_487;
wire n_451;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_84;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_109;
wire n_132;
wire n_406;
wire n_395;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g75 ( .A(n_24), .Y(n_75) );
NOR2xp33_ASAP7_75t_L g76 ( .A(n_41), .B(n_46), .Y(n_76) );
CKINVDCx5p33_ASAP7_75t_R g77 ( .A(n_55), .Y(n_77) );
INVx1_ASAP7_75t_L g78 ( .A(n_39), .Y(n_78) );
INVx1_ASAP7_75t_L g79 ( .A(n_49), .Y(n_79) );
INVx1_ASAP7_75t_L g80 ( .A(n_56), .Y(n_80) );
INVx1_ASAP7_75t_L g81 ( .A(n_70), .Y(n_81) );
CKINVDCx20_ASAP7_75t_R g82 ( .A(n_69), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_47), .Y(n_83) );
INVx1_ASAP7_75t_L g84 ( .A(n_35), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_12), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_54), .Y(n_86) );
CKINVDCx5p33_ASAP7_75t_R g87 ( .A(n_25), .Y(n_87) );
BUFx2_ASAP7_75t_SL g88 ( .A(n_38), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_29), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_21), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_10), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_51), .Y(n_92) );
CKINVDCx14_ASAP7_75t_R g93 ( .A(n_73), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_71), .Y(n_94) );
INVx2_ASAP7_75t_L g95 ( .A(n_31), .Y(n_95) );
INVx2_ASAP7_75t_L g96 ( .A(n_12), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_1), .Y(n_97) );
CKINVDCx16_ASAP7_75t_R g98 ( .A(n_44), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_45), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_63), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_62), .Y(n_101) );
INVxp33_ASAP7_75t_SL g102 ( .A(n_60), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_68), .Y(n_103) );
INVx1_ASAP7_75t_SL g104 ( .A(n_11), .Y(n_104) );
CKINVDCx20_ASAP7_75t_R g105 ( .A(n_40), .Y(n_105) );
CKINVDCx20_ASAP7_75t_R g106 ( .A(n_48), .Y(n_106) );
CKINVDCx5p33_ASAP7_75t_R g107 ( .A(n_27), .Y(n_107) );
CKINVDCx5p33_ASAP7_75t_R g108 ( .A(n_8), .Y(n_108) );
CKINVDCx20_ASAP7_75t_R g109 ( .A(n_42), .Y(n_109) );
CKINVDCx5p33_ASAP7_75t_R g110 ( .A(n_66), .Y(n_110) );
INVxp33_ASAP7_75t_L g111 ( .A(n_22), .Y(n_111) );
INVx2_ASAP7_75t_L g112 ( .A(n_7), .Y(n_112) );
INVxp67_ASAP7_75t_SL g113 ( .A(n_11), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_6), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_15), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_72), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_6), .Y(n_117) );
INVxp67_ASAP7_75t_L g118 ( .A(n_50), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_5), .Y(n_119) );
CKINVDCx16_ASAP7_75t_R g120 ( .A(n_67), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_0), .Y(n_121) );
NAND2xp5_ASAP7_75t_L g122 ( .A(n_108), .B(n_0), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_84), .Y(n_123) );
INVx2_ASAP7_75t_L g124 ( .A(n_95), .Y(n_124) );
NAND2xp5_ASAP7_75t_L g125 ( .A(n_108), .B(n_1), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_84), .Y(n_126) );
NAND2xp5_ASAP7_75t_SL g127 ( .A(n_95), .B(n_2), .Y(n_127) );
AND2x4_ASAP7_75t_L g128 ( .A(n_96), .B(n_112), .Y(n_128) );
INVx1_ASAP7_75t_L g129 ( .A(n_86), .Y(n_129) );
INVx1_ASAP7_75t_L g130 ( .A(n_86), .Y(n_130) );
INVx1_ASAP7_75t_L g131 ( .A(n_89), .Y(n_131) );
INVx1_ASAP7_75t_L g132 ( .A(n_89), .Y(n_132) );
INVx2_ASAP7_75t_L g133 ( .A(n_75), .Y(n_133) );
BUFx2_ASAP7_75t_L g134 ( .A(n_98), .Y(n_134) );
NAND2xp5_ASAP7_75t_L g135 ( .A(n_91), .B(n_2), .Y(n_135) );
HB1xp67_ASAP7_75t_L g136 ( .A(n_85), .Y(n_136) );
INVx1_ASAP7_75t_L g137 ( .A(n_96), .Y(n_137) );
AND2x4_ASAP7_75t_L g138 ( .A(n_112), .B(n_3), .Y(n_138) );
AND2x4_ASAP7_75t_L g139 ( .A(n_85), .B(n_3), .Y(n_139) );
INVx2_ASAP7_75t_L g140 ( .A(n_78), .Y(n_140) );
NAND2xp5_ASAP7_75t_L g141 ( .A(n_97), .B(n_4), .Y(n_141) );
NAND2xp5_ASAP7_75t_L g142 ( .A(n_114), .B(n_4), .Y(n_142) );
OA21x2_ASAP7_75t_L g143 ( .A1(n_79), .A2(n_30), .B(n_65), .Y(n_143) );
OR2x6_ASAP7_75t_L g144 ( .A(n_88), .B(n_5), .Y(n_144) );
INVx3_ASAP7_75t_L g145 ( .A(n_80), .Y(n_145) );
BUFx2_ASAP7_75t_L g146 ( .A(n_120), .Y(n_146) );
HB1xp67_ASAP7_75t_L g147 ( .A(n_115), .Y(n_147) );
BUFx2_ASAP7_75t_L g148 ( .A(n_93), .Y(n_148) );
INVx2_ASAP7_75t_L g149 ( .A(n_81), .Y(n_149) );
INVx1_ASAP7_75t_L g150 ( .A(n_83), .Y(n_150) );
INVx1_ASAP7_75t_L g151 ( .A(n_90), .Y(n_151) );
BUFx6f_ASAP7_75t_L g152 ( .A(n_92), .Y(n_152) );
NAND3xp33_ASAP7_75t_L g153 ( .A(n_117), .B(n_28), .C(n_64), .Y(n_153) );
AND2x4_ASAP7_75t_L g154 ( .A(n_121), .B(n_7), .Y(n_154) );
NAND2xp5_ASAP7_75t_L g155 ( .A(n_119), .B(n_8), .Y(n_155) );
INVx1_ASAP7_75t_L g156 ( .A(n_94), .Y(n_156) );
INVx2_ASAP7_75t_L g157 ( .A(n_99), .Y(n_157) );
INVx2_ASAP7_75t_L g158 ( .A(n_100), .Y(n_158) );
INVx3_ASAP7_75t_L g159 ( .A(n_101), .Y(n_159) );
INVx2_ASAP7_75t_L g160 ( .A(n_103), .Y(n_160) );
INVx2_ASAP7_75t_L g161 ( .A(n_116), .Y(n_161) );
INVx1_ASAP7_75t_L g162 ( .A(n_88), .Y(n_162) );
NAND2x1p5_ASAP7_75t_L g163 ( .A(n_139), .B(n_104), .Y(n_163) );
BUFx6f_ASAP7_75t_L g164 ( .A(n_143), .Y(n_164) );
INVx2_ASAP7_75t_L g165 ( .A(n_152), .Y(n_165) );
INVx2_ASAP7_75t_L g166 ( .A(n_152), .Y(n_166) );
INVxp67_ASAP7_75t_L g167 ( .A(n_134), .Y(n_167) );
INVx2_ASAP7_75t_L g168 ( .A(n_152), .Y(n_168) );
INVx1_ASAP7_75t_L g169 ( .A(n_162), .Y(n_169) );
AND2x6_ASAP7_75t_L g170 ( .A(n_139), .B(n_76), .Y(n_170) );
NAND2x1p5_ASAP7_75t_L g171 ( .A(n_139), .B(n_102), .Y(n_171) );
INVx1_ASAP7_75t_L g172 ( .A(n_152), .Y(n_172) );
AND2x4_ASAP7_75t_L g173 ( .A(n_162), .B(n_128), .Y(n_173) );
BUFx2_ASAP7_75t_L g174 ( .A(n_148), .Y(n_174) );
NAND2xp5_ASAP7_75t_SL g175 ( .A(n_148), .B(n_77), .Y(n_175) );
BUFx3_ASAP7_75t_L g176 ( .A(n_128), .Y(n_176) );
INVx2_ASAP7_75t_L g177 ( .A(n_152), .Y(n_177) );
AND2x6_ASAP7_75t_L g178 ( .A(n_139), .B(n_102), .Y(n_178) );
INVx2_ASAP7_75t_L g179 ( .A(n_152), .Y(n_179) );
INVx2_ASAP7_75t_L g180 ( .A(n_124), .Y(n_180) );
INVx4_ASAP7_75t_L g181 ( .A(n_144), .Y(n_181) );
INVx2_ASAP7_75t_L g182 ( .A(n_124), .Y(n_182) );
OAI221xp5_ASAP7_75t_L g183 ( .A1(n_147), .A2(n_113), .B1(n_118), .B2(n_107), .C(n_110), .Y(n_183) );
INVx3_ASAP7_75t_L g184 ( .A(n_138), .Y(n_184) );
INVx1_ASAP7_75t_L g185 ( .A(n_124), .Y(n_185) );
CKINVDCx20_ASAP7_75t_R g186 ( .A(n_134), .Y(n_186) );
INVx2_ASAP7_75t_L g187 ( .A(n_137), .Y(n_187) );
INVx1_ASAP7_75t_L g188 ( .A(n_138), .Y(n_188) );
AND2x2_ASAP7_75t_L g189 ( .A(n_146), .B(n_111), .Y(n_189) );
INVx1_ASAP7_75t_L g190 ( .A(n_138), .Y(n_190) );
BUFx6f_ASAP7_75t_L g191 ( .A(n_143), .Y(n_191) );
INVx2_ASAP7_75t_L g192 ( .A(n_137), .Y(n_192) );
INVx1_ASAP7_75t_L g193 ( .A(n_138), .Y(n_193) );
AND2x2_ASAP7_75t_L g194 ( .A(n_146), .B(n_110), .Y(n_194) );
NAND2x1p5_ASAP7_75t_L g195 ( .A(n_154), .B(n_107), .Y(n_195) );
AND2x2_ASAP7_75t_L g196 ( .A(n_136), .B(n_87), .Y(n_196) );
AND2x4_ASAP7_75t_L g197 ( .A(n_128), .B(n_87), .Y(n_197) );
INVx1_ASAP7_75t_L g198 ( .A(n_123), .Y(n_198) );
INVxp67_ASAP7_75t_L g199 ( .A(n_122), .Y(n_199) );
NAND2xp5_ASAP7_75t_L g200 ( .A(n_150), .B(n_77), .Y(n_200) );
OAI22xp33_ASAP7_75t_L g201 ( .A1(n_144), .A2(n_109), .B1(n_106), .B2(n_105), .Y(n_201) );
AND2x4_ASAP7_75t_L g202 ( .A(n_128), .B(n_109), .Y(n_202) );
INVx1_ASAP7_75t_L g203 ( .A(n_123), .Y(n_203) );
BUFx6f_ASAP7_75t_L g204 ( .A(n_143), .Y(n_204) );
INVx1_ASAP7_75t_L g205 ( .A(n_126), .Y(n_205) );
NAND2xp5_ASAP7_75t_SL g206 ( .A(n_126), .B(n_106), .Y(n_206) );
AND3x1_ASAP7_75t_L g207 ( .A(n_125), .B(n_105), .C(n_82), .Y(n_207) );
INVx3_ASAP7_75t_L g208 ( .A(n_154), .Y(n_208) );
AO22x2_ASAP7_75t_L g209 ( .A1(n_154), .A2(n_82), .B1(n_10), .B2(n_13), .Y(n_209) );
INVx3_ASAP7_75t_L g210 ( .A(n_154), .Y(n_210) );
BUFx6f_ASAP7_75t_L g211 ( .A(n_143), .Y(n_211) );
INVx1_ASAP7_75t_L g212 ( .A(n_129), .Y(n_212) );
INVx4_ASAP7_75t_L g213 ( .A(n_144), .Y(n_213) );
INVx1_ASAP7_75t_L g214 ( .A(n_129), .Y(n_214) );
INVx5_ASAP7_75t_L g215 ( .A(n_144), .Y(n_215) );
INVx2_ASAP7_75t_L g216 ( .A(n_145), .Y(n_216) );
INVx1_ASAP7_75t_L g217 ( .A(n_130), .Y(n_217) );
INVx1_ASAP7_75t_L g218 ( .A(n_130), .Y(n_218) );
INVx1_ASAP7_75t_L g219 ( .A(n_131), .Y(n_219) );
INVxp67_ASAP7_75t_L g220 ( .A(n_144), .Y(n_220) );
BUFx6f_ASAP7_75t_L g221 ( .A(n_157), .Y(n_221) );
INVx2_ASAP7_75t_L g222 ( .A(n_145), .Y(n_222) );
BUFx2_ASAP7_75t_L g223 ( .A(n_181), .Y(n_223) );
NAND2xp5_ASAP7_75t_L g224 ( .A(n_199), .B(n_131), .Y(n_224) );
INVx2_ASAP7_75t_L g225 ( .A(n_221), .Y(n_225) );
BUFx6f_ASAP7_75t_L g226 ( .A(n_164), .Y(n_226) );
INVx1_ASAP7_75t_L g227 ( .A(n_216), .Y(n_227) );
BUFx6f_ASAP7_75t_L g228 ( .A(n_164), .Y(n_228) );
INVx5_ASAP7_75t_L g229 ( .A(n_215), .Y(n_229) );
INVx2_ASAP7_75t_L g230 ( .A(n_221), .Y(n_230) );
BUFx2_ASAP7_75t_L g231 ( .A(n_181), .Y(n_231) );
AND2x2_ASAP7_75t_L g232 ( .A(n_196), .B(n_156), .Y(n_232) );
AND2x2_ASAP7_75t_L g233 ( .A(n_196), .B(n_156), .Y(n_233) );
INVx2_ASAP7_75t_L g234 ( .A(n_221), .Y(n_234) );
NOR2xp33_ASAP7_75t_L g235 ( .A(n_175), .B(n_150), .Y(n_235) );
NAND2xp5_ASAP7_75t_L g236 ( .A(n_200), .B(n_132), .Y(n_236) );
AND2x4_ASAP7_75t_L g237 ( .A(n_181), .B(n_151), .Y(n_237) );
INVx1_ASAP7_75t_L g238 ( .A(n_216), .Y(n_238) );
INVx2_ASAP7_75t_L g239 ( .A(n_221), .Y(n_239) );
BUFx6f_ASAP7_75t_L g240 ( .A(n_164), .Y(n_240) );
INVx2_ASAP7_75t_L g241 ( .A(n_221), .Y(n_241) );
INVx1_ASAP7_75t_L g242 ( .A(n_222), .Y(n_242) );
BUFx6f_ASAP7_75t_SL g243 ( .A(n_213), .Y(n_243) );
INVx2_ASAP7_75t_SL g244 ( .A(n_215), .Y(n_244) );
CKINVDCx5p33_ASAP7_75t_R g245 ( .A(n_186), .Y(n_245) );
HB1xp67_ASAP7_75t_L g246 ( .A(n_174), .Y(n_246) );
AOI22xp33_ASAP7_75t_L g247 ( .A1(n_213), .A2(n_151), .B1(n_159), .B2(n_145), .Y(n_247) );
OR2x2_ASAP7_75t_L g248 ( .A(n_167), .B(n_155), .Y(n_248) );
NAND2xp5_ASAP7_75t_L g249 ( .A(n_197), .B(n_132), .Y(n_249) );
AOI22xp5_ASAP7_75t_L g250 ( .A1(n_213), .A2(n_145), .B1(n_159), .B2(n_135), .Y(n_250) );
INVx1_ASAP7_75t_L g251 ( .A(n_222), .Y(n_251) );
INVx1_ASAP7_75t_L g252 ( .A(n_185), .Y(n_252) );
NAND2xp5_ASAP7_75t_SL g253 ( .A(n_215), .B(n_141), .Y(n_253) );
INVx1_ASAP7_75t_L g254 ( .A(n_185), .Y(n_254) );
NAND2xp5_ASAP7_75t_L g255 ( .A(n_197), .B(n_159), .Y(n_255) );
BUFx3_ASAP7_75t_L g256 ( .A(n_176), .Y(n_256) );
HB1xp67_ASAP7_75t_L g257 ( .A(n_174), .Y(n_257) );
INVx2_ASAP7_75t_L g258 ( .A(n_165), .Y(n_258) );
INVx2_ASAP7_75t_SL g259 ( .A(n_215), .Y(n_259) );
AND2x6_ASAP7_75t_L g260 ( .A(n_208), .B(n_159), .Y(n_260) );
AND3x2_ASAP7_75t_SL g261 ( .A(n_209), .B(n_158), .C(n_149), .Y(n_261) );
AND2x4_ASAP7_75t_L g262 ( .A(n_215), .B(n_149), .Y(n_262) );
BUFx6f_ASAP7_75t_L g263 ( .A(n_164), .Y(n_263) );
NAND2xp5_ASAP7_75t_L g264 ( .A(n_197), .B(n_158), .Y(n_264) );
INVx2_ASAP7_75t_L g265 ( .A(n_165), .Y(n_265) );
NAND2xp5_ASAP7_75t_L g266 ( .A(n_169), .B(n_133), .Y(n_266) );
AND2x2_ASAP7_75t_L g267 ( .A(n_194), .B(n_140), .Y(n_267) );
INVx3_ASAP7_75t_L g268 ( .A(n_184), .Y(n_268) );
INVx1_ASAP7_75t_L g269 ( .A(n_198), .Y(n_269) );
INVx1_ASAP7_75t_L g270 ( .A(n_198), .Y(n_270) );
INVx2_ASAP7_75t_SL g271 ( .A(n_163), .Y(n_271) );
INVx2_ASAP7_75t_L g272 ( .A(n_166), .Y(n_272) );
INVx1_ASAP7_75t_L g273 ( .A(n_203), .Y(n_273) );
BUFx3_ASAP7_75t_L g274 ( .A(n_176), .Y(n_274) );
NAND2xp5_ASAP7_75t_L g275 ( .A(n_173), .B(n_133), .Y(n_275) );
AOI22xp33_ASAP7_75t_L g276 ( .A1(n_178), .A2(n_140), .B1(n_160), .B2(n_157), .Y(n_276) );
NAND2xp5_ASAP7_75t_SL g277 ( .A(n_195), .B(n_142), .Y(n_277) );
INVx2_ASAP7_75t_L g278 ( .A(n_166), .Y(n_278) );
AOI22xp5_ASAP7_75t_L g279 ( .A1(n_209), .A2(n_161), .B1(n_160), .B2(n_157), .Y(n_279) );
NAND2xp5_ASAP7_75t_L g280 ( .A(n_173), .B(n_161), .Y(n_280) );
AND2x2_ASAP7_75t_L g281 ( .A(n_194), .B(n_161), .Y(n_281) );
INVx1_ASAP7_75t_L g282 ( .A(n_203), .Y(n_282) );
OAI21x1_ASAP7_75t_L g283 ( .A1(n_208), .A2(n_160), .B(n_153), .Y(n_283) );
INVx2_ASAP7_75t_L g284 ( .A(n_168), .Y(n_284) );
INVx2_ASAP7_75t_SL g285 ( .A(n_163), .Y(n_285) );
INVx2_ASAP7_75t_L g286 ( .A(n_269), .Y(n_286) );
AND2x2_ASAP7_75t_L g287 ( .A(n_232), .B(n_202), .Y(n_287) );
BUFx6f_ASAP7_75t_L g288 ( .A(n_226), .Y(n_288) );
OR2x2_ASAP7_75t_L g289 ( .A(n_248), .B(n_201), .Y(n_289) );
BUFx6f_ASAP7_75t_L g290 ( .A(n_226), .Y(n_290) );
AND2x4_ASAP7_75t_L g291 ( .A(n_285), .B(n_220), .Y(n_291) );
NAND2xp5_ASAP7_75t_SL g292 ( .A(n_223), .B(n_195), .Y(n_292) );
AOI222xp33_ASAP7_75t_L g293 ( .A1(n_245), .A2(n_202), .B1(n_189), .B2(n_186), .C1(n_206), .C2(n_183), .Y(n_293) );
OAI21x1_ASAP7_75t_SL g294 ( .A1(n_279), .A2(n_193), .B(n_188), .Y(n_294) );
INVx2_ASAP7_75t_L g295 ( .A(n_269), .Y(n_295) );
AOI21xp5_ASAP7_75t_L g296 ( .A1(n_270), .A2(n_193), .B(n_188), .Y(n_296) );
AND2x4_ASAP7_75t_L g297 ( .A(n_271), .B(n_173), .Y(n_297) );
INVx3_ASAP7_75t_L g298 ( .A(n_229), .Y(n_298) );
INVx1_ASAP7_75t_L g299 ( .A(n_252), .Y(n_299) );
NOR2x1_ASAP7_75t_L g300 ( .A(n_277), .B(n_237), .Y(n_300) );
INVx4_ASAP7_75t_L g301 ( .A(n_229), .Y(n_301) );
INVx1_ASAP7_75t_L g302 ( .A(n_252), .Y(n_302) );
INVx1_ASAP7_75t_SL g303 ( .A(n_246), .Y(n_303) );
INVx2_ASAP7_75t_L g304 ( .A(n_270), .Y(n_304) );
OR2x2_ASAP7_75t_L g305 ( .A(n_248), .B(n_202), .Y(n_305) );
AND2x2_ASAP7_75t_L g306 ( .A(n_232), .B(n_209), .Y(n_306) );
BUFx6f_ASAP7_75t_L g307 ( .A(n_226), .Y(n_307) );
HB1xp67_ASAP7_75t_L g308 ( .A(n_257), .Y(n_308) );
BUFx6f_ASAP7_75t_L g309 ( .A(n_226), .Y(n_309) );
BUFx12f_ASAP7_75t_L g310 ( .A(n_245), .Y(n_310) );
AND2x6_ASAP7_75t_L g311 ( .A(n_237), .B(n_208), .Y(n_311) );
INVx2_ASAP7_75t_L g312 ( .A(n_273), .Y(n_312) );
INVxp67_ASAP7_75t_SL g313 ( .A(n_279), .Y(n_313) );
INVx2_ASAP7_75t_L g314 ( .A(n_273), .Y(n_314) );
BUFx12f_ASAP7_75t_L g315 ( .A(n_271), .Y(n_315) );
BUFx2_ASAP7_75t_L g316 ( .A(n_260), .Y(n_316) );
INVx1_ASAP7_75t_L g317 ( .A(n_254), .Y(n_317) );
AO32x2_ASAP7_75t_L g318 ( .A1(n_261), .A2(n_209), .A3(n_164), .B1(n_211), .B2(n_204), .Y(n_318) );
AOI21xp33_ASAP7_75t_L g319 ( .A1(n_285), .A2(n_189), .B(n_190), .Y(n_319) );
INVx3_ASAP7_75t_L g320 ( .A(n_229), .Y(n_320) );
INVx4_ASAP7_75t_L g321 ( .A(n_229), .Y(n_321) );
AND2x4_ASAP7_75t_L g322 ( .A(n_237), .B(n_223), .Y(n_322) );
AOI21xp33_ASAP7_75t_L g323 ( .A1(n_231), .A2(n_171), .B(n_163), .Y(n_323) );
INVx1_ASAP7_75t_L g324 ( .A(n_254), .Y(n_324) );
INVx2_ASAP7_75t_L g325 ( .A(n_282), .Y(n_325) );
NOR2xp33_ASAP7_75t_L g326 ( .A(n_224), .B(n_171), .Y(n_326) );
INVx2_ASAP7_75t_SL g327 ( .A(n_237), .Y(n_327) );
CKINVDCx8_ASAP7_75t_R g328 ( .A(n_229), .Y(n_328) );
INVx2_ASAP7_75t_L g329 ( .A(n_282), .Y(n_329) );
INVx2_ASAP7_75t_L g330 ( .A(n_227), .Y(n_330) );
HB1xp67_ASAP7_75t_L g331 ( .A(n_233), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_268), .Y(n_332) );
INVx2_ASAP7_75t_L g333 ( .A(n_227), .Y(n_333) );
CKINVDCx11_ASAP7_75t_R g334 ( .A(n_310), .Y(n_334) );
OAI22xp5_ASAP7_75t_L g335 ( .A1(n_313), .A2(n_171), .B1(n_195), .B2(n_250), .Y(n_335) );
HB1xp67_ASAP7_75t_L g336 ( .A(n_303), .Y(n_336) );
HB1xp67_ASAP7_75t_L g337 ( .A(n_303), .Y(n_337) );
INVx2_ASAP7_75t_L g338 ( .A(n_286), .Y(n_338) );
AND2x4_ASAP7_75t_L g339 ( .A(n_322), .B(n_229), .Y(n_339) );
BUFx2_ASAP7_75t_L g340 ( .A(n_308), .Y(n_340) );
BUFx3_ASAP7_75t_L g341 ( .A(n_328), .Y(n_341) );
OAI22xp5_ASAP7_75t_L g342 ( .A1(n_306), .A2(n_250), .B1(n_249), .B2(n_276), .Y(n_342) );
OAI221xp5_ASAP7_75t_L g343 ( .A1(n_293), .A2(n_235), .B1(n_207), .B2(n_233), .C(n_267), .Y(n_343) );
INVx8_ASAP7_75t_L g344 ( .A(n_315), .Y(n_344) );
OAI21xp5_ASAP7_75t_L g345 ( .A1(n_296), .A2(n_283), .B(n_236), .Y(n_345) );
CKINVDCx11_ASAP7_75t_R g346 ( .A(n_310), .Y(n_346) );
NAND2x1p5_ASAP7_75t_L g347 ( .A(n_322), .B(n_231), .Y(n_347) );
AOI22xp33_ASAP7_75t_SL g348 ( .A1(n_306), .A2(n_261), .B1(n_243), .B2(n_281), .Y(n_348) );
AND2x4_ASAP7_75t_L g349 ( .A(n_322), .B(n_281), .Y(n_349) );
AOI22xp33_ASAP7_75t_L g350 ( .A1(n_287), .A2(n_178), .B1(n_267), .B2(n_210), .Y(n_350) );
NAND2xp5_ASAP7_75t_L g351 ( .A(n_326), .B(n_264), .Y(n_351) );
AOI22xp33_ASAP7_75t_L g352 ( .A1(n_287), .A2(n_178), .B1(n_210), .B2(n_184), .Y(n_352) );
AOI22xp5_ASAP7_75t_L g353 ( .A1(n_322), .A2(n_178), .B1(n_243), .B2(n_260), .Y(n_353) );
AOI22xp33_ASAP7_75t_SL g354 ( .A1(n_289), .A2(n_261), .B1(n_243), .B2(n_178), .Y(n_354) );
OAI22xp5_ASAP7_75t_L g355 ( .A1(n_305), .A2(n_280), .B1(n_275), .B2(n_255), .Y(n_355) );
OAI22xp5_ASAP7_75t_L g356 ( .A1(n_305), .A2(n_247), .B1(n_210), .B2(n_184), .Y(n_356) );
INVx2_ASAP7_75t_SL g357 ( .A(n_315), .Y(n_357) );
CKINVDCx16_ASAP7_75t_R g358 ( .A(n_289), .Y(n_358) );
A2O1A1Ixp33_ASAP7_75t_L g359 ( .A1(n_286), .A2(n_266), .B(n_205), .C(n_218), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_331), .Y(n_360) );
OAI21x1_ASAP7_75t_L g361 ( .A1(n_295), .A2(n_283), .B(n_230), .Y(n_361) );
NOR2xp33_ASAP7_75t_L g362 ( .A(n_319), .B(n_274), .Y(n_362) );
OAI22xp33_ASAP7_75t_L g363 ( .A1(n_327), .A2(n_274), .B1(n_268), .B2(n_256), .Y(n_363) );
AOI22xp5_ASAP7_75t_L g364 ( .A1(n_358), .A2(n_311), .B1(n_178), .B2(n_291), .Y(n_364) );
AO22x1_ASAP7_75t_L g365 ( .A1(n_335), .A2(n_318), .B1(n_311), .B2(n_299), .Y(n_365) );
OAI222xp33_ASAP7_75t_L g366 ( .A1(n_348), .A2(n_292), .B1(n_299), .B2(n_317), .C1(n_302), .C2(n_324), .Y(n_366) );
INVx1_ASAP7_75t_L g367 ( .A(n_360), .Y(n_367) );
NAND2xp5_ASAP7_75t_L g368 ( .A(n_349), .B(n_302), .Y(n_368) );
NAND2xp5_ASAP7_75t_L g369 ( .A(n_349), .B(n_317), .Y(n_369) );
AOI22xp33_ASAP7_75t_L g370 ( .A1(n_343), .A2(n_178), .B1(n_294), .B2(n_311), .Y(n_370) );
AOI22xp33_ASAP7_75t_SL g371 ( .A1(n_336), .A2(n_294), .B1(n_311), .B2(n_316), .Y(n_371) );
AND2x2_ASAP7_75t_L g372 ( .A(n_349), .B(n_330), .Y(n_372) );
AOI22xp33_ASAP7_75t_SL g373 ( .A1(n_337), .A2(n_311), .B1(n_316), .B2(n_291), .Y(n_373) );
AOI22xp33_ASAP7_75t_L g374 ( .A1(n_354), .A2(n_311), .B1(n_323), .B2(n_170), .Y(n_374) );
AOI22xp33_ASAP7_75t_L g375 ( .A1(n_362), .A2(n_311), .B1(n_170), .B2(n_300), .Y(n_375) );
INVx1_ASAP7_75t_L g376 ( .A(n_338), .Y(n_376) );
O2A1O1Ixp5_ASAP7_75t_L g377 ( .A1(n_345), .A2(n_314), .B(n_295), .C(n_304), .Y(n_377) );
BUFx4f_ASAP7_75t_L g378 ( .A(n_347), .Y(n_378) );
BUFx3_ASAP7_75t_L g379 ( .A(n_344), .Y(n_379) );
NAND2xp5_ASAP7_75t_L g380 ( .A(n_351), .B(n_324), .Y(n_380) );
OAI22xp33_ASAP7_75t_L g381 ( .A1(n_340), .A2(n_344), .B1(n_353), .B2(n_347), .Y(n_381) );
AND2x2_ASAP7_75t_L g382 ( .A(n_338), .B(n_330), .Y(n_382) );
AOI22xp5_ASAP7_75t_L g383 ( .A1(n_355), .A2(n_291), .B1(n_327), .B2(n_297), .Y(n_383) );
INVx2_ASAP7_75t_L g384 ( .A(n_361), .Y(n_384) );
OAI221xp5_ASAP7_75t_L g385 ( .A1(n_350), .A2(n_300), .B1(n_312), .B2(n_329), .C(n_304), .Y(n_385) );
AOI22xp5_ASAP7_75t_L g386 ( .A1(n_362), .A2(n_291), .B1(n_297), .B2(n_260), .Y(n_386) );
INVx1_ASAP7_75t_L g387 ( .A(n_359), .Y(n_387) );
AND2x4_ASAP7_75t_L g388 ( .A(n_339), .B(n_301), .Y(n_388) );
OAI221xp5_ASAP7_75t_L g389 ( .A1(n_350), .A2(n_329), .B1(n_325), .B2(n_314), .C(n_312), .Y(n_389) );
OAI221xp5_ASAP7_75t_L g390 ( .A1(n_352), .A2(n_325), .B1(n_332), .B2(n_127), .C(n_256), .Y(n_390) );
INVx5_ASAP7_75t_L g391 ( .A(n_379), .Y(n_391) );
AOI22xp33_ASAP7_75t_L g392 ( .A1(n_370), .A2(n_342), .B1(n_170), .B2(n_352), .Y(n_392) );
INVx1_ASAP7_75t_L g393 ( .A(n_367), .Y(n_393) );
AOI22xp5_ASAP7_75t_L g394 ( .A1(n_364), .A2(n_356), .B1(n_344), .B2(n_357), .Y(n_394) );
AND2x4_ASAP7_75t_L g395 ( .A(n_388), .B(n_339), .Y(n_395) );
AOI33xp33_ASAP7_75t_L g396 ( .A1(n_381), .A2(n_192), .A3(n_187), .B1(n_212), .B2(n_217), .B3(n_205), .Y(n_396) );
INVx2_ASAP7_75t_SL g397 ( .A(n_378), .Y(n_397) );
AOI221xp5_ASAP7_75t_SL g398 ( .A1(n_366), .A2(n_359), .B1(n_192), .B2(n_187), .C(n_217), .Y(n_398) );
AND2x2_ASAP7_75t_L g399 ( .A(n_382), .B(n_318), .Y(n_399) );
NAND3xp33_ASAP7_75t_L g400 ( .A(n_387), .B(n_182), .C(n_180), .Y(n_400) );
NAND2xp5_ASAP7_75t_L g401 ( .A(n_380), .B(n_339), .Y(n_401) );
OR2x6_ASAP7_75t_L g402 ( .A(n_379), .B(n_341), .Y(n_402) );
NOR2x1_ASAP7_75t_SL g403 ( .A(n_378), .B(n_341), .Y(n_403) );
AOI21xp5_ASAP7_75t_L g404 ( .A1(n_365), .A2(n_309), .B(n_307), .Y(n_404) );
OAI21xp33_ASAP7_75t_L g405 ( .A1(n_387), .A2(n_180), .B(n_182), .Y(n_405) );
INVx1_ASAP7_75t_L g406 ( .A(n_376), .Y(n_406) );
AND2x2_ASAP7_75t_L g407 ( .A(n_372), .B(n_318), .Y(n_407) );
OR2x2_ASAP7_75t_L g408 ( .A(n_368), .B(n_333), .Y(n_408) );
AO21x2_ASAP7_75t_L g409 ( .A1(n_384), .A2(n_363), .B(n_318), .Y(n_409) );
AOI22xp33_ASAP7_75t_L g410 ( .A1(n_378), .A2(n_170), .B1(n_333), .B2(n_297), .Y(n_410) );
OR2x2_ASAP7_75t_L g411 ( .A(n_369), .B(n_297), .Y(n_411) );
AND2x2_ASAP7_75t_L g412 ( .A(n_372), .B(n_382), .Y(n_412) );
AOI21xp5_ASAP7_75t_L g413 ( .A1(n_365), .A2(n_307), .B(n_290), .Y(n_413) );
AOI222xp33_ASAP7_75t_L g414 ( .A1(n_374), .A2(n_346), .B1(n_334), .B2(n_170), .C1(n_214), .C2(n_218), .Y(n_414) );
AOI22xp33_ASAP7_75t_L g415 ( .A1(n_383), .A2(n_170), .B1(n_332), .B2(n_274), .Y(n_415) );
AND2x4_ASAP7_75t_L g416 ( .A(n_388), .B(n_301), .Y(n_416) );
AO21x2_ASAP7_75t_L g417 ( .A1(n_384), .A2(n_318), .B(n_253), .Y(n_417) );
AOI222xp33_ASAP7_75t_L g418 ( .A1(n_385), .A2(n_170), .B1(n_214), .B2(n_219), .C1(n_260), .C2(n_251), .Y(n_418) );
INVx1_ASAP7_75t_L g419 ( .A(n_376), .Y(n_419) );
AOI22xp33_ASAP7_75t_L g420 ( .A1(n_371), .A2(n_211), .B1(n_204), .B2(n_191), .Y(n_420) );
AOI222xp33_ASAP7_75t_L g421 ( .A1(n_389), .A2(n_219), .B1(n_260), .B2(n_251), .C1(n_238), .C2(n_242), .Y(n_421) );
INVx2_ASAP7_75t_L g422 ( .A(n_377), .Y(n_422) );
NAND3xp33_ASAP7_75t_L g423 ( .A(n_375), .B(n_172), .C(n_211), .Y(n_423) );
OAI211xp5_ASAP7_75t_L g424 ( .A1(n_373), .A2(n_328), .B(n_321), .C(n_301), .Y(n_424) );
AND2x2_ASAP7_75t_L g425 ( .A(n_388), .B(n_9), .Y(n_425) );
INVx2_ASAP7_75t_SL g426 ( .A(n_391), .Y(n_426) );
INVx2_ASAP7_75t_SL g427 ( .A(n_391), .Y(n_427) );
AOI22xp33_ASAP7_75t_L g428 ( .A1(n_392), .A2(n_390), .B1(n_386), .B2(n_211), .Y(n_428) );
INVx2_ASAP7_75t_L g429 ( .A(n_406), .Y(n_429) );
OAI31xp33_ASAP7_75t_L g430 ( .A1(n_397), .A2(n_262), .A3(n_320), .B(n_298), .Y(n_430) );
INVx1_ASAP7_75t_L g431 ( .A(n_393), .Y(n_431) );
NAND2xp5_ASAP7_75t_L g432 ( .A(n_412), .B(n_9), .Y(n_432) );
INVx2_ASAP7_75t_L g433 ( .A(n_419), .Y(n_433) );
INVx1_ASAP7_75t_L g434 ( .A(n_408), .Y(n_434) );
NOR2xp33_ASAP7_75t_L g435 ( .A(n_401), .B(n_13), .Y(n_435) );
NOR2xp67_ASAP7_75t_L g436 ( .A(n_391), .B(n_14), .Y(n_436) );
HB1xp67_ASAP7_75t_L g437 ( .A(n_409), .Y(n_437) );
AOI22xp5_ASAP7_75t_L g438 ( .A1(n_414), .A2(n_260), .B1(n_262), .B2(n_301), .Y(n_438) );
INVxp67_ASAP7_75t_SL g439 ( .A(n_399), .Y(n_439) );
OAI22xp5_ASAP7_75t_L g440 ( .A1(n_410), .A2(n_392), .B1(n_415), .B2(n_394), .Y(n_440) );
OAI33xp33_ASAP7_75t_L g441 ( .A1(n_411), .A2(n_172), .A3(n_15), .B1(n_16), .B2(n_17), .B3(n_14), .Y(n_441) );
INVx1_ASAP7_75t_L g442 ( .A(n_425), .Y(n_442) );
INVxp67_ASAP7_75t_SL g443 ( .A(n_399), .Y(n_443) );
INVx1_ASAP7_75t_L g444 ( .A(n_396), .Y(n_444) );
NAND2xp5_ASAP7_75t_L g445 ( .A(n_396), .B(n_16), .Y(n_445) );
INVx1_ASAP7_75t_L g446 ( .A(n_391), .Y(n_446) );
BUFx6f_ASAP7_75t_L g447 ( .A(n_416), .Y(n_447) );
INVx1_ASAP7_75t_L g448 ( .A(n_397), .Y(n_448) );
AND2x2_ASAP7_75t_L g449 ( .A(n_395), .B(n_17), .Y(n_449) );
AND2x4_ASAP7_75t_L g450 ( .A(n_416), .B(n_321), .Y(n_450) );
NAND3xp33_ASAP7_75t_L g451 ( .A(n_398), .B(n_168), .C(n_177), .Y(n_451) );
INVx1_ASAP7_75t_L g452 ( .A(n_407), .Y(n_452) );
BUFx3_ASAP7_75t_L g453 ( .A(n_402), .Y(n_453) );
HB1xp67_ASAP7_75t_L g454 ( .A(n_409), .Y(n_454) );
INVx1_ASAP7_75t_L g455 ( .A(n_395), .Y(n_455) );
AOI33xp33_ASAP7_75t_L g456 ( .A1(n_410), .A2(n_177), .A3(n_179), .B1(n_238), .B2(n_242), .B3(n_262), .Y(n_456) );
INVx2_ASAP7_75t_L g457 ( .A(n_422), .Y(n_457) );
OR2x2_ASAP7_75t_SL g458 ( .A(n_403), .B(n_402), .Y(n_458) );
INVx5_ASAP7_75t_L g459 ( .A(n_402), .Y(n_459) );
NAND2xp5_ASAP7_75t_L g460 ( .A(n_416), .B(n_191), .Y(n_460) );
OR2x2_ASAP7_75t_L g461 ( .A(n_395), .B(n_417), .Y(n_461) );
INVx1_ASAP7_75t_L g462 ( .A(n_400), .Y(n_462) );
OAI33xp33_ASAP7_75t_L g463 ( .A1(n_422), .A2(n_179), .A3(n_241), .B1(n_239), .B2(n_234), .B3(n_230), .Y(n_463) );
HB1xp67_ASAP7_75t_L g464 ( .A(n_417), .Y(n_464) );
INVx1_ASAP7_75t_SL g465 ( .A(n_404), .Y(n_465) );
AOI22xp33_ASAP7_75t_L g466 ( .A1(n_421), .A2(n_191), .B1(n_204), .B2(n_211), .Y(n_466) );
OAI321xp33_ASAP7_75t_L g467 ( .A1(n_420), .A2(n_191), .A3(n_204), .B1(n_225), .B2(n_234), .C(n_239), .Y(n_467) );
AND2x2_ASAP7_75t_L g468 ( .A(n_415), .B(n_321), .Y(n_468) );
OAI22xp5_ASAP7_75t_L g469 ( .A1(n_420), .A2(n_321), .B1(n_320), .B2(n_298), .Y(n_469) );
INVx3_ASAP7_75t_L g470 ( .A(n_424), .Y(n_470) );
INVx1_ASAP7_75t_L g471 ( .A(n_405), .Y(n_471) );
AND2x4_ASAP7_75t_L g472 ( .A(n_413), .B(n_320), .Y(n_472) );
INVx1_ASAP7_75t_L g473 ( .A(n_423), .Y(n_473) );
OR2x2_ASAP7_75t_L g474 ( .A(n_418), .B(n_298), .Y(n_474) );
INVx1_ASAP7_75t_L g475 ( .A(n_393), .Y(n_475) );
OR2x2_ASAP7_75t_L g476 ( .A(n_439), .B(n_204), .Y(n_476) );
INVx5_ASAP7_75t_L g477 ( .A(n_459), .Y(n_477) );
AND2x2_ASAP7_75t_L g478 ( .A(n_439), .B(n_443), .Y(n_478) );
INVx2_ASAP7_75t_L g479 ( .A(n_457), .Y(n_479) );
NOR2xp33_ASAP7_75t_L g480 ( .A(n_442), .B(n_18), .Y(n_480) );
AND2x4_ASAP7_75t_SL g481 ( .A(n_447), .B(n_309), .Y(n_481) );
NAND2xp5_ASAP7_75t_L g482 ( .A(n_434), .B(n_191), .Y(n_482) );
AND2x2_ASAP7_75t_L g483 ( .A(n_443), .B(n_19), .Y(n_483) );
NAND2xp5_ASAP7_75t_L g484 ( .A(n_431), .B(n_268), .Y(n_484) );
INVx2_ASAP7_75t_L g485 ( .A(n_457), .Y(n_485) );
AND2x2_ASAP7_75t_L g486 ( .A(n_452), .B(n_20), .Y(n_486) );
INVx1_ASAP7_75t_L g487 ( .A(n_475), .Y(n_487) );
OAI33xp33_ASAP7_75t_L g488 ( .A1(n_432), .A2(n_241), .A3(n_225), .B1(n_32), .B2(n_33), .B3(n_34), .Y(n_488) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_429), .B(n_260), .Y(n_489) );
AND2x2_ASAP7_75t_L g490 ( .A(n_429), .B(n_23), .Y(n_490) );
AND2x2_ASAP7_75t_L g491 ( .A(n_433), .B(n_26), .Y(n_491) );
INVxp67_ASAP7_75t_L g492 ( .A(n_426), .Y(n_492) );
NOR2xp33_ASAP7_75t_L g493 ( .A(n_435), .B(n_36), .Y(n_493) );
INVx1_ASAP7_75t_L g494 ( .A(n_433), .Y(n_494) );
AND2x2_ASAP7_75t_L g495 ( .A(n_461), .B(n_37), .Y(n_495) );
INVx2_ASAP7_75t_L g496 ( .A(n_464), .Y(n_496) );
INVx1_ASAP7_75t_SL g497 ( .A(n_427), .Y(n_497) );
INVx1_ASAP7_75t_L g498 ( .A(n_446), .Y(n_498) );
INVx3_ASAP7_75t_SL g499 ( .A(n_458), .Y(n_499) );
INVx2_ASAP7_75t_L g500 ( .A(n_464), .Y(n_500) );
HB1xp67_ASAP7_75t_L g501 ( .A(n_447), .Y(n_501) );
OR2x2_ASAP7_75t_L g502 ( .A(n_437), .B(n_43), .Y(n_502) );
OAI222xp33_ASAP7_75t_L g503 ( .A1(n_459), .A2(n_262), .B1(n_244), .B2(n_259), .C1(n_58), .C2(n_59), .Y(n_503) );
INVx1_ASAP7_75t_L g504 ( .A(n_448), .Y(n_504) );
INVx1_ASAP7_75t_L g505 ( .A(n_455), .Y(n_505) );
INVx1_ASAP7_75t_L g506 ( .A(n_453), .Y(n_506) );
AND2x2_ASAP7_75t_L g507 ( .A(n_437), .B(n_52), .Y(n_507) );
INVx1_ASAP7_75t_L g508 ( .A(n_453), .Y(n_508) );
INVx1_ASAP7_75t_L g509 ( .A(n_454), .Y(n_509) );
NOR3xp33_ASAP7_75t_SL g510 ( .A(n_441), .B(n_53), .C(n_57), .Y(n_510) );
INVx1_ASAP7_75t_L g511 ( .A(n_454), .Y(n_511) );
INVx1_ASAP7_75t_L g512 ( .A(n_444), .Y(n_512) );
OR2x2_ASAP7_75t_L g513 ( .A(n_447), .B(n_61), .Y(n_513) );
INVx1_ASAP7_75t_L g514 ( .A(n_472), .Y(n_514) );
AND2x2_ASAP7_75t_L g515 ( .A(n_472), .B(n_74), .Y(n_515) );
OR2x2_ASAP7_75t_L g516 ( .A(n_445), .B(n_226), .Y(n_516) );
AND2x2_ASAP7_75t_L g517 ( .A(n_465), .B(n_228), .Y(n_517) );
AND2x2_ASAP7_75t_L g518 ( .A(n_460), .B(n_449), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_435), .B(n_228), .Y(n_519) );
INVx1_ASAP7_75t_L g520 ( .A(n_436), .Y(n_520) );
AND2x2_ASAP7_75t_L g521 ( .A(n_468), .B(n_228), .Y(n_521) );
AND2x2_ASAP7_75t_L g522 ( .A(n_473), .B(n_228), .Y(n_522) );
INVx1_ASAP7_75t_L g523 ( .A(n_471), .Y(n_523) );
OR2x2_ASAP7_75t_L g524 ( .A(n_470), .B(n_228), .Y(n_524) );
INVx2_ASAP7_75t_L g525 ( .A(n_462), .Y(n_525) );
AND2x2_ASAP7_75t_L g526 ( .A(n_470), .B(n_240), .Y(n_526) );
OR2x2_ASAP7_75t_L g527 ( .A(n_440), .B(n_240), .Y(n_527) );
INVx1_ASAP7_75t_L g528 ( .A(n_459), .Y(n_528) );
NAND3xp33_ASAP7_75t_L g529 ( .A(n_456), .B(n_240), .C(n_263), .Y(n_529) );
INVx2_ASAP7_75t_L g530 ( .A(n_459), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_450), .B(n_240), .Y(n_531) );
NAND3xp33_ASAP7_75t_L g532 ( .A(n_456), .B(n_240), .C(n_263), .Y(n_532) );
AND2x4_ASAP7_75t_L g533 ( .A(n_514), .B(n_450), .Y(n_533) );
INVx1_ASAP7_75t_L g534 ( .A(n_487), .Y(n_534) );
AND2x2_ASAP7_75t_L g535 ( .A(n_518), .B(n_474), .Y(n_535) );
OAI21xp33_ASAP7_75t_L g536 ( .A1(n_512), .A2(n_428), .B(n_466), .Y(n_536) );
NOR2xp33_ASAP7_75t_L g537 ( .A(n_520), .B(n_463), .Y(n_537) );
INVxp67_ASAP7_75t_SL g538 ( .A(n_496), .Y(n_538) );
OAI22xp5_ASAP7_75t_L g539 ( .A1(n_499), .A2(n_466), .B1(n_428), .B2(n_438), .Y(n_539) );
INVx1_ASAP7_75t_L g540 ( .A(n_498), .Y(n_540) );
INVx1_ASAP7_75t_SL g541 ( .A(n_497), .Y(n_541) );
AND2x2_ASAP7_75t_L g542 ( .A(n_478), .B(n_451), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_478), .B(n_504), .Y(n_543) );
NOR2xp33_ASAP7_75t_L g544 ( .A(n_492), .B(n_469), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_505), .B(n_518), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_494), .B(n_430), .Y(n_546) );
INVx2_ASAP7_75t_L g547 ( .A(n_494), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_523), .B(n_263), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g549 ( .A(n_523), .B(n_263), .Y(n_549) );
OR2x2_ASAP7_75t_L g550 ( .A(n_509), .B(n_309), .Y(n_550) );
BUFx2_ASAP7_75t_L g551 ( .A(n_499), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g552 ( .A(n_511), .B(n_263), .Y(n_552) );
AND2x2_ASAP7_75t_L g553 ( .A(n_501), .B(n_309), .Y(n_553) );
INVxp67_ASAP7_75t_L g554 ( .A(n_525), .Y(n_554) );
OAI211xp5_ASAP7_75t_L g555 ( .A1(n_493), .A2(n_244), .B(n_259), .C(n_467), .Y(n_555) );
NAND2x1_ASAP7_75t_L g556 ( .A(n_528), .B(n_307), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g557 ( .A(n_506), .B(n_307), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g558 ( .A(n_508), .B(n_307), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g559 ( .A(n_525), .B(n_288), .Y(n_559) );
OAI21xp33_ASAP7_75t_L g560 ( .A1(n_510), .A2(n_258), .B(n_265), .Y(n_560) );
OAI31xp33_ASAP7_75t_L g561 ( .A1(n_503), .A2(n_258), .A3(n_265), .B(n_272), .Y(n_561) );
INVxp67_ASAP7_75t_L g562 ( .A(n_496), .Y(n_562) );
AND2x2_ASAP7_75t_L g563 ( .A(n_479), .B(n_290), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g564 ( .A(n_485), .B(n_288), .Y(n_564) );
INVx1_ASAP7_75t_L g565 ( .A(n_485), .Y(n_565) );
AND2x2_ASAP7_75t_L g566 ( .A(n_495), .B(n_288), .Y(n_566) );
OR2x2_ASAP7_75t_L g567 ( .A(n_500), .B(n_290), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g568 ( .A(n_507), .B(n_290), .Y(n_568) );
NOR2xp33_ASAP7_75t_L g569 ( .A(n_480), .B(n_290), .Y(n_569) );
OR2x2_ASAP7_75t_L g570 ( .A(n_500), .B(n_272), .Y(n_570) );
INVx2_ASAP7_75t_SL g571 ( .A(n_477), .Y(n_571) );
INVxp67_ASAP7_75t_L g572 ( .A(n_483), .Y(n_572) );
INVx1_ASAP7_75t_L g573 ( .A(n_502), .Y(n_573) );
NOR2x1_ASAP7_75t_L g574 ( .A(n_529), .B(n_278), .Y(n_574) );
OR2x2_ASAP7_75t_L g575 ( .A(n_476), .B(n_278), .Y(n_575) );
AND2x2_ASAP7_75t_L g576 ( .A(n_495), .B(n_507), .Y(n_576) );
AND2x2_ASAP7_75t_L g577 ( .A(n_483), .B(n_284), .Y(n_577) );
AND2x2_ASAP7_75t_L g578 ( .A(n_521), .B(n_284), .Y(n_578) );
OR2x2_ASAP7_75t_L g579 ( .A(n_476), .B(n_502), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g580 ( .A(n_482), .B(n_528), .Y(n_580) );
AND2x2_ASAP7_75t_L g581 ( .A(n_545), .B(n_521), .Y(n_581) );
INVxp67_ASAP7_75t_SL g582 ( .A(n_538), .Y(n_582) );
INVx1_ASAP7_75t_L g583 ( .A(n_540), .Y(n_583) );
INVx1_ASAP7_75t_L g584 ( .A(n_547), .Y(n_584) );
INVxp67_ASAP7_75t_L g585 ( .A(n_551), .Y(n_585) );
NAND2xp5_ASAP7_75t_L g586 ( .A(n_543), .B(n_530), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g587 ( .A(n_537), .B(n_530), .Y(n_587) );
INVx1_ASAP7_75t_L g588 ( .A(n_547), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g589 ( .A(n_537), .B(n_486), .Y(n_589) );
AND2x2_ASAP7_75t_L g590 ( .A(n_533), .B(n_517), .Y(n_590) );
AOI21xp33_ASAP7_75t_L g591 ( .A1(n_544), .A2(n_515), .B(n_486), .Y(n_591) );
INVx2_ASAP7_75t_L g592 ( .A(n_565), .Y(n_592) );
NOR3xp33_ASAP7_75t_L g593 ( .A(n_539), .B(n_560), .C(n_555), .Y(n_593) );
INVx1_ASAP7_75t_L g594 ( .A(n_534), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g595 ( .A(n_535), .B(n_515), .Y(n_595) );
NAND2xp33_ASAP7_75t_L g596 ( .A(n_571), .B(n_477), .Y(n_596) );
INVx1_ASAP7_75t_L g597 ( .A(n_580), .Y(n_597) );
AOI211x1_ASAP7_75t_L g598 ( .A1(n_536), .A2(n_532), .B(n_519), .C(n_484), .Y(n_598) );
INVx1_ASAP7_75t_L g599 ( .A(n_554), .Y(n_599) );
OAI221xp5_ASAP7_75t_L g600 ( .A1(n_544), .A2(n_541), .B1(n_572), .B2(n_546), .C(n_561), .Y(n_600) );
INVxp67_ASAP7_75t_L g601 ( .A(n_533), .Y(n_601) );
OAI222xp33_ASAP7_75t_L g602 ( .A1(n_572), .A2(n_477), .B1(n_513), .B2(n_491), .C1(n_490), .C2(n_527), .Y(n_602) );
HB1xp67_ASAP7_75t_L g603 ( .A(n_562), .Y(n_603) );
OR2x2_ASAP7_75t_L g604 ( .A(n_562), .B(n_527), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g605 ( .A(n_573), .B(n_516), .Y(n_605) );
INVx1_ASAP7_75t_SL g606 ( .A(n_571), .Y(n_606) );
INVx2_ASAP7_75t_SL g607 ( .A(n_556), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g608 ( .A(n_542), .B(n_516), .Y(n_608) );
INVx1_ASAP7_75t_SL g609 ( .A(n_533), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g610 ( .A(n_542), .B(n_490), .Y(n_610) );
INVx1_ASAP7_75t_L g611 ( .A(n_538), .Y(n_611) );
INVx1_ASAP7_75t_L g612 ( .A(n_579), .Y(n_612) );
AOI211x1_ASAP7_75t_L g613 ( .A1(n_576), .A2(n_491), .B(n_489), .C(n_526), .Y(n_613) );
HB1xp67_ASAP7_75t_L g614 ( .A(n_570), .Y(n_614) );
OAI22xp5_ASAP7_75t_L g615 ( .A1(n_574), .A2(n_477), .B1(n_513), .B2(n_531), .Y(n_615) );
INVxp67_ASAP7_75t_SL g616 ( .A(n_575), .Y(n_616) );
INVx1_ASAP7_75t_L g617 ( .A(n_578), .Y(n_617) );
INVx2_ASAP7_75t_L g618 ( .A(n_567), .Y(n_618) );
AOI21xp5_ASAP7_75t_L g619 ( .A1(n_568), .A2(n_488), .B(n_477), .Y(n_619) );
INVx1_ASAP7_75t_L g620 ( .A(n_578), .Y(n_620) );
NAND2xp5_ASAP7_75t_SL g621 ( .A(n_566), .B(n_550), .Y(n_621) );
XNOR2x1_ASAP7_75t_L g622 ( .A(n_577), .B(n_524), .Y(n_622) );
INVx1_ASAP7_75t_L g623 ( .A(n_548), .Y(n_623) );
AOI21xp33_ASAP7_75t_L g624 ( .A1(n_557), .A2(n_524), .B(n_526), .Y(n_624) );
O2A1O1Ixp33_ASAP7_75t_L g625 ( .A1(n_558), .A2(n_481), .B(n_522), .C(n_552), .Y(n_625) );
INVx1_ASAP7_75t_L g626 ( .A(n_549), .Y(n_626) );
INVx1_ASAP7_75t_SL g627 ( .A(n_553), .Y(n_627) );
INVx1_ASAP7_75t_L g628 ( .A(n_559), .Y(n_628) );
XOR2x2_ASAP7_75t_L g629 ( .A(n_569), .B(n_481), .Y(n_629) );
INVx1_ASAP7_75t_L g630 ( .A(n_564), .Y(n_630) );
O2A1O1Ixp33_ASAP7_75t_L g631 ( .A1(n_569), .A2(n_537), .B(n_512), .C(n_520), .Y(n_631) );
OAI21xp5_ASAP7_75t_L g632 ( .A1(n_563), .A2(n_537), .B(n_551), .Y(n_632) );
AOI221xp5_ASAP7_75t_L g633 ( .A1(n_537), .A2(n_512), .B1(n_534), .B2(n_545), .C(n_540), .Y(n_633) );
OAI21xp5_ASAP7_75t_L g634 ( .A1(n_593), .A2(n_585), .B(n_631), .Y(n_634) );
INVx1_ASAP7_75t_L g635 ( .A(n_587), .Y(n_635) );
NAND2xp5_ASAP7_75t_L g636 ( .A(n_633), .B(n_616), .Y(n_636) );
AOI21xp5_ASAP7_75t_L g637 ( .A1(n_596), .A2(n_607), .B(n_600), .Y(n_637) );
XNOR2xp5_ASAP7_75t_L g638 ( .A(n_622), .B(n_629), .Y(n_638) );
INVx2_ASAP7_75t_L g639 ( .A(n_611), .Y(n_639) );
AOI322xp5_ASAP7_75t_L g640 ( .A1(n_589), .A2(n_612), .A3(n_581), .B1(n_609), .B2(n_601), .C1(n_616), .C2(n_582), .Y(n_640) );
XNOR2xp5_ASAP7_75t_L g641 ( .A(n_581), .B(n_614), .Y(n_641) );
INVx1_ASAP7_75t_L g642 ( .A(n_603), .Y(n_642) );
NAND3xp33_ASAP7_75t_SL g643 ( .A(n_632), .B(n_606), .C(n_619), .Y(n_643) );
OAI21xp5_ASAP7_75t_L g644 ( .A1(n_596), .A2(n_607), .B(n_591), .Y(n_644) );
OAI21xp33_ASAP7_75t_L g645 ( .A1(n_597), .A2(n_586), .B(n_608), .Y(n_645) );
INVx1_ASAP7_75t_L g646 ( .A(n_599), .Y(n_646) );
NAND4xp25_ASAP7_75t_L g647 ( .A(n_637), .B(n_598), .C(n_613), .D(n_625), .Y(n_647) );
NAND3xp33_ASAP7_75t_L g648 ( .A(n_637), .B(n_611), .C(n_583), .Y(n_648) );
NOR3xp33_ASAP7_75t_SL g649 ( .A(n_643), .B(n_602), .C(n_615), .Y(n_649) );
AOI21xp33_ASAP7_75t_L g650 ( .A1(n_634), .A2(n_605), .B(n_594), .Y(n_650) );
OAI211xp5_ASAP7_75t_SL g651 ( .A1(n_640), .A2(n_621), .B(n_595), .C(n_610), .Y(n_651) );
NOR3xp33_ASAP7_75t_L g652 ( .A(n_643), .B(n_626), .C(n_623), .Y(n_652) );
NAND3xp33_ASAP7_75t_SL g653 ( .A(n_644), .B(n_627), .C(n_604), .Y(n_653) );
AOI22xp5_ASAP7_75t_L g654 ( .A1(n_647), .A2(n_638), .B1(n_636), .B2(n_635), .Y(n_654) );
AOI211xp5_ASAP7_75t_L g655 ( .A1(n_650), .A2(n_642), .B(n_645), .C(n_641), .Y(n_655) );
NAND2x1p5_ASAP7_75t_L g656 ( .A(n_648), .B(n_621), .Y(n_656) );
NAND4xp25_ASAP7_75t_L g657 ( .A(n_651), .B(n_646), .C(n_624), .D(n_604), .Y(n_657) );
AOI22xp5_ASAP7_75t_L g658 ( .A1(n_654), .A2(n_653), .B1(n_652), .B2(n_649), .Y(n_658) );
XNOR2xp5_ASAP7_75t_L g659 ( .A(n_655), .B(n_590), .Y(n_659) );
INVx1_ASAP7_75t_L g660 ( .A(n_657), .Y(n_660) );
INVx1_ASAP7_75t_L g661 ( .A(n_660), .Y(n_661) );
AOI21xp5_ASAP7_75t_L g662 ( .A1(n_658), .A2(n_656), .B(n_639), .Y(n_662) );
INVx1_ASAP7_75t_L g663 ( .A(n_661), .Y(n_663) );
OAI22x1_ASAP7_75t_L g664 ( .A1(n_663), .A2(n_659), .B1(n_662), .B2(n_618), .Y(n_664) );
AOI22xp33_ASAP7_75t_L g665 ( .A1(n_664), .A2(n_628), .B1(n_630), .B2(n_620), .Y(n_665) );
AOI221xp5_ASAP7_75t_L g666 ( .A1(n_665), .A2(n_617), .B1(n_588), .B2(n_584), .C(n_592), .Y(n_666) );
endmodule