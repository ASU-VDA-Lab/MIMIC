module fake_jpeg_27254_n_64 (n_13, n_21, n_1, n_10, n_23, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_64);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_64;

wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_27;
wire n_55;
wire n_51;
wire n_47;
wire n_40;
wire n_59;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_62;
wire n_31;
wire n_25;
wire n_56;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_32;

INVx1_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_SL g25 ( 
.A(n_9),
.B(n_17),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_19),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_10),
.Y(n_28)
);

BUFx4f_ASAP7_75t_L g29 ( 
.A(n_22),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_2),
.B(n_15),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_26),
.B(n_0),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_31),
.B(n_32),
.Y(n_42)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_29),
.Y(n_32)
);

CKINVDCx14_ASAP7_75t_R g33 ( 
.A(n_30),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_33),
.B(n_36),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_26),
.B(n_0),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_34),
.B(n_35),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_24),
.B(n_1),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_29),
.B(n_1),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_29),
.B(n_2),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_37),
.B(n_3),
.Y(n_49)
);

BUFx2_ASAP7_75t_L g38 ( 
.A(n_27),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_38),
.Y(n_39)
);

AOI22x1_ASAP7_75t_SL g40 ( 
.A1(n_36),
.A2(n_27),
.B1(n_14),
.B2(n_23),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_40),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g41 ( 
.A1(n_32),
.A2(n_28),
.B1(n_25),
.B2(n_24),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_41),
.A2(n_45),
.B1(n_5),
.B2(n_6),
.Y(n_55)
);

XNOR2xp5_ASAP7_75t_L g43 ( 
.A(n_37),
.B(n_38),
.Y(n_43)
);

XNOR2xp5_ASAP7_75t_SL g57 ( 
.A(n_43),
.B(n_7),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g45 ( 
.A1(n_36),
.A2(n_11),
.B1(n_20),
.B2(n_18),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_35),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_46),
.Y(n_52)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_38),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_48),
.B(n_49),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_50),
.A2(n_53),
.B1(n_54),
.B2(n_55),
.Y(n_58)
);

MAJIxp5_ASAP7_75t_L g51 ( 
.A(n_43),
.B(n_21),
.C(n_16),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_51),
.A2(n_57),
.B1(n_40),
.B2(n_41),
.Y(n_59)
);

MAJIxp5_ASAP7_75t_L g53 ( 
.A(n_47),
.B(n_13),
.C(n_12),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_44),
.B(n_4),
.Y(n_54)
);

INVxp67_ASAP7_75t_L g60 ( 
.A(n_59),
.Y(n_60)
);

AOI221x1_ASAP7_75t_L g61 ( 
.A1(n_60),
.A2(n_59),
.B1(n_57),
.B2(n_58),
.C(n_51),
.Y(n_61)
);

AOI21xp5_ASAP7_75t_L g62 ( 
.A1(n_61),
.A2(n_42),
.B(n_56),
.Y(n_62)
);

AO21x1_ASAP7_75t_L g63 ( 
.A1(n_62),
.A2(n_52),
.B(n_39),
.Y(n_63)
);

XOR2xp5_ASAP7_75t_L g64 ( 
.A(n_63),
.B(n_8),
.Y(n_64)
);


endmodule