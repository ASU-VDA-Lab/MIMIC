module fake_jpeg_22009_n_54 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_54);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_54;

wire n_13;
wire n_21;
wire n_53;
wire n_33;
wire n_45;
wire n_23;
wire n_10;
wire n_27;
wire n_47;
wire n_22;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_44;
wire n_38;
wire n_26;
wire n_28;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_31;
wire n_25;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;

CKINVDCx20_ASAP7_75t_R g8 ( 
.A(n_2),
.Y(n_8)
);

INVx8_ASAP7_75t_L g9 ( 
.A(n_1),
.Y(n_9)
);

CKINVDCx16_ASAP7_75t_R g10 ( 
.A(n_1),
.Y(n_10)
);

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_4),
.Y(n_11)
);

INVx2_ASAP7_75t_L g12 ( 
.A(n_4),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_3),
.Y(n_13)
);

BUFx12f_ASAP7_75t_L g14 ( 
.A(n_7),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

NAND3xp33_ASAP7_75t_L g16 ( 
.A(n_15),
.B(n_0),
.C(n_2),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_SL g23 ( 
.A(n_16),
.B(n_15),
.Y(n_23)
);

INVx6_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_17),
.Y(n_22)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_18),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_19),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

OR2x2_ASAP7_75t_L g27 ( 
.A(n_20),
.B(n_21),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

CKINVDCx14_ASAP7_75t_R g30 ( 
.A(n_23),
.Y(n_30)
);

NOR2x1_ASAP7_75t_L g24 ( 
.A(n_20),
.B(n_8),
.Y(n_24)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_24),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_24),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_29),
.B(n_31),
.Y(n_40)
);

INVxp67_ASAP7_75t_L g31 ( 
.A(n_27),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_22),
.Y(n_32)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_32),
.Y(n_41)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_22),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_33),
.B(n_34),
.Y(n_39)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_26),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_L g35 ( 
.A1(n_25),
.A2(n_12),
.B1(n_9),
.B2(n_18),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_L g37 ( 
.A1(n_35),
.A2(n_25),
.B1(n_13),
.B2(n_11),
.Y(n_37)
);

INVxp67_ASAP7_75t_L g36 ( 
.A(n_32),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_SL g43 ( 
.A(n_36),
.B(n_37),
.Y(n_43)
);

MAJIxp5_ASAP7_75t_L g38 ( 
.A(n_31),
.B(n_27),
.C(n_10),
.Y(n_38)
);

XNOR2xp5_ASAP7_75t_L g45 ( 
.A(n_38),
.B(n_30),
.Y(n_45)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_39),
.Y(n_42)
);

MAJIxp5_ASAP7_75t_L g47 ( 
.A(n_42),
.B(n_44),
.C(n_45),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_40),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_43),
.A2(n_28),
.B1(n_36),
.B2(n_41),
.Y(n_46)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_46),
.Y(n_49)
);

MAJIxp5_ASAP7_75t_L g48 ( 
.A(n_47),
.B(n_45),
.C(n_3),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g50 ( 
.A(n_48),
.B(n_6),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_50),
.B(n_0),
.Y(n_51)
);

OAI21x1_ASAP7_75t_SL g52 ( 
.A1(n_51),
.A2(n_5),
.B(n_6),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_52),
.B(n_49),
.Y(n_53)
);

BUFx24_ASAP7_75t_SL g54 ( 
.A(n_53),
.Y(n_54)
);


endmodule