module real_aes_10737_n_12 (n_4, n_0, n_3, n_5, n_2, n_7, n_8, n_6, n_9, n_1, n_10, n_11, n_12);
input n_4;
input n_0;
input n_3;
input n_5;
input n_2;
input n_7;
input n_8;
input n_6;
input n_9;
input n_1;
input n_10;
input n_11;
output n_12;
wire n_17;
wire n_22;
wire n_13;
wire n_24;
wire n_19;
wire n_25;
wire n_14;
wire n_16;
wire n_15;
wire n_23;
wire n_20;
wire n_18;
wire n_26;
wire n_21;
NOR2xp33_ASAP7_75t_R g21 ( .A(n_0), .B(n_5), .Y(n_21) );
NOR3xp33_ASAP7_75t_SL g19 ( .A(n_1), .B(n_7), .C(n_20), .Y(n_19) );
NAND2xp33_ASAP7_75t_R g20 ( .A(n_2), .B(n_21), .Y(n_20) );
CKINVDCx5p33_ASAP7_75t_R g22 ( .A(n_3), .Y(n_22) );
NOR4xp25_ASAP7_75t_SL g17 ( .A(n_4), .B(n_18), .C(n_22), .D(n_23), .Y(n_17) );
NAND2xp33_ASAP7_75t_SL g14 ( .A(n_6), .B(n_15), .Y(n_14) );
NAND2xp33_ASAP7_75t_R g26 ( .A(n_6), .B(n_10), .Y(n_26) );
AOI22xp33_ASAP7_75t_L g12 ( .A1(n_8), .A2(n_11), .B1(n_13), .B2(n_24), .Y(n_12) );
CKINVDCx5p33_ASAP7_75t_R g23 ( .A(n_9), .Y(n_23) );
CKINVDCx5p33_ASAP7_75t_R g15 ( .A(n_10), .Y(n_15) );
NOR2xp33_ASAP7_75t_R g13 ( .A(n_14), .B(n_16), .Y(n_13) );
NOR2xp33_ASAP7_75t_R g25 ( .A(n_16), .B(n_26), .Y(n_25) );
CKINVDCx5p33_ASAP7_75t_R g16 ( .A(n_17), .Y(n_16) );
CKINVDCx5p33_ASAP7_75t_R g18 ( .A(n_19), .Y(n_18) );
HB1xp67_ASAP7_75t_L g24 ( .A(n_25), .Y(n_24) );
endmodule