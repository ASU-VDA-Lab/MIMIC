module fake_jpeg_30011_n_258 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_258);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_258;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_182;
wire n_19;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx3_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_15),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_7),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_16),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_11),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_10),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_0),
.B(n_3),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_24),
.Y(n_35)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

BUFx12_ASAP7_75t_L g37 ( 
.A(n_17),
.Y(n_37)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_33),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_38),
.B(n_27),
.Y(n_44)
);

BUFx10_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_24),
.Y(n_40)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_40),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_33),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_41),
.B(n_27),
.Y(n_48)
);

INVx13_ASAP7_75t_L g42 ( 
.A(n_19),
.Y(n_42)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_42),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_18),
.Y(n_43)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_43),
.Y(n_56)
);

OR2x2_ASAP7_75t_L g75 ( 
.A(n_44),
.B(n_52),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g45 ( 
.A1(n_38),
.A2(n_25),
.B1(n_26),
.B2(n_34),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_L g71 ( 
.A1(n_45),
.A2(n_57),
.B1(n_61),
.B2(n_21),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_48),
.B(n_44),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_35),
.A2(n_19),
.B1(n_17),
.B2(n_34),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_51),
.A2(n_28),
.B1(n_43),
.B2(n_36),
.Y(n_70)
);

NAND2x1_ASAP7_75t_L g52 ( 
.A(n_35),
.B(n_40),
.Y(n_52)
);

HB1xp67_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_53),
.Y(n_69)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_54),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_38),
.A2(n_25),
.B1(n_26),
.B2(n_34),
.Y(n_57)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_42),
.Y(n_59)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_59),
.Y(n_72)
);

NAND2xp33_ASAP7_75t_SL g60 ( 
.A(n_39),
.B(n_17),
.Y(n_60)
);

NAND3xp33_ASAP7_75t_SL g96 ( 
.A(n_60),
.B(n_39),
.C(n_42),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_41),
.A2(n_26),
.B1(n_21),
.B2(n_23),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_37),
.B(n_30),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_62),
.B(n_20),
.Y(n_74)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_47),
.Y(n_64)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_64),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_65),
.B(n_74),
.Y(n_98)
);

INVx5_ASAP7_75t_L g66 ( 
.A(n_46),
.Y(n_66)
);

INVx4_ASAP7_75t_L g115 ( 
.A(n_66),
.Y(n_115)
);

OAI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_61),
.A2(n_43),
.B1(n_36),
.B2(n_23),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_67),
.A2(n_22),
.B1(n_37),
.B2(n_2),
.Y(n_109)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_47),
.Y(n_68)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_68),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_70),
.A2(n_71),
.B1(n_89),
.B2(n_93),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_49),
.B(n_39),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_73),
.B(n_80),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_52),
.B(n_30),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g119 ( 
.A(n_76),
.B(n_77),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_46),
.B(n_20),
.Y(n_77)
);

BUFx12_ASAP7_75t_L g78 ( 
.A(n_58),
.Y(n_78)
);

INVx13_ASAP7_75t_L g123 ( 
.A(n_78),
.Y(n_123)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_54),
.Y(n_79)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_79),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_49),
.B(n_39),
.Y(n_80)
);

INVx2_ASAP7_75t_SL g81 ( 
.A(n_59),
.Y(n_81)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_81),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_52),
.B(n_29),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_82),
.B(n_87),
.Y(n_104)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_56),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_83),
.Y(n_113)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_58),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_84),
.Y(n_99)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_56),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g122 ( 
.A(n_85),
.B(n_92),
.Y(n_122)
);

BUFx2_ASAP7_75t_L g86 ( 
.A(n_55),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_86),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_45),
.B(n_29),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_57),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_88),
.B(n_91),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_L g89 ( 
.A1(n_55),
.A2(n_43),
.B1(n_21),
.B2(n_23),
.Y(n_89)
);

BUFx3_ASAP7_75t_L g90 ( 
.A(n_55),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_90),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_50),
.B(n_32),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_50),
.B(n_32),
.Y(n_92)
);

INVx2_ASAP7_75t_SL g93 ( 
.A(n_50),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_93),
.B(n_94),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_60),
.B(n_12),
.Y(n_94)
);

INVx1_ASAP7_75t_SL g95 ( 
.A(n_46),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_L g103 ( 
.A1(n_95),
.A2(n_97),
.B1(n_28),
.B2(n_39),
.Y(n_103)
);

A2O1A1Ixp33_ASAP7_75t_SL g114 ( 
.A1(n_96),
.A2(n_0),
.B(n_4),
.C(n_5),
.Y(n_114)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_47),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_75),
.B(n_28),
.C(n_31),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_L g143 ( 
.A(n_101),
.B(n_106),
.Y(n_143)
);

A2O1A1Ixp33_ASAP7_75t_L g102 ( 
.A1(n_75),
.A2(n_31),
.B(n_22),
.C(n_12),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_102),
.B(n_124),
.Y(n_146)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_103),
.Y(n_130)
);

XOR2xp5_ASAP7_75t_L g106 ( 
.A(n_73),
.B(n_42),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g147 ( 
.A(n_109),
.B(n_111),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_110),
.A2(n_112),
.B1(n_93),
.B2(n_95),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_63),
.A2(n_37),
.B1(n_1),
.B2(n_2),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_80),
.A2(n_37),
.B1(n_2),
.B2(n_3),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_SL g139 ( 
.A1(n_114),
.A2(n_84),
.B(n_4),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_69),
.B(n_16),
.C(n_15),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_122),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_125),
.B(n_129),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_126),
.B(n_128),
.Y(n_163)
);

AOI21xp5_ASAP7_75t_L g127 ( 
.A1(n_105),
.A2(n_81),
.B(n_63),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g154 ( 
.A(n_127),
.Y(n_154)
);

AO22x2_ASAP7_75t_L g128 ( 
.A1(n_110),
.A2(n_68),
.B1(n_97),
.B2(n_64),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_98),
.B(n_72),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_107),
.B(n_72),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_131),
.B(n_134),
.Y(n_161)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_120),
.Y(n_132)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_132),
.Y(n_152)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_118),
.Y(n_133)
);

HB1xp67_ASAP7_75t_L g170 ( 
.A(n_133),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_119),
.B(n_81),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_122),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_135),
.B(n_139),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_106),
.A2(n_85),
.B1(n_83),
.B2(n_86),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_136),
.A2(n_137),
.B1(n_127),
.B2(n_143),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_104),
.A2(n_112),
.B1(n_122),
.B2(n_100),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_121),
.Y(n_138)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_138),
.Y(n_153)
);

INVx8_ASAP7_75t_L g140 ( 
.A(n_115),
.Y(n_140)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_140),
.Y(n_156)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_121),
.Y(n_141)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_141),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_100),
.B(n_66),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_142),
.B(n_144),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_105),
.B(n_90),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_101),
.B(n_78),
.Y(n_145)
);

CKINVDCx16_ASAP7_75t_R g174 ( 
.A(n_145),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_108),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_148),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_116),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_149),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_L g150 ( 
.A1(n_114),
.A2(n_78),
.B(n_4),
.Y(n_150)
);

OR2x2_ASAP7_75t_L g160 ( 
.A(n_150),
.B(n_114),
.Y(n_160)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_113),
.Y(n_151)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_151),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_159),
.B(n_143),
.Y(n_182)
);

INVxp67_ASAP7_75t_L g195 ( 
.A(n_160),
.Y(n_195)
);

OA21x2_ASAP7_75t_L g162 ( 
.A1(n_142),
.A2(n_114),
.B(n_109),
.Y(n_162)
);

AND2x2_ASAP7_75t_L g183 ( 
.A(n_162),
.B(n_137),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_144),
.Y(n_164)
);

OR2x2_ASAP7_75t_L g189 ( 
.A(n_164),
.B(n_133),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_147),
.A2(n_117),
.B1(n_102),
.B2(n_99),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_166),
.B(n_168),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_147),
.A2(n_99),
.B1(n_113),
.B2(n_111),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_147),
.A2(n_126),
.B1(n_130),
.B2(n_128),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_169),
.B(n_173),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_L g172 ( 
.A1(n_130),
.A2(n_115),
.B1(n_123),
.B2(n_7),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_L g181 ( 
.A1(n_172),
.A2(n_150),
.B1(n_140),
.B2(n_151),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_128),
.A2(n_0),
.B1(n_6),
.B2(n_8),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_128),
.A2(n_6),
.B1(n_9),
.B2(n_13),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_175),
.A2(n_6),
.B1(n_9),
.B2(n_14),
.Y(n_193)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_165),
.Y(n_178)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_178),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_161),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_SL g200 ( 
.A(n_180),
.B(n_188),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_181),
.A2(n_182),
.B1(n_193),
.B2(n_196),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_SL g209 ( 
.A1(n_183),
.A2(n_154),
.B(n_163),
.Y(n_209)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_165),
.Y(n_184)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_184),
.Y(n_202)
);

A2O1A1O1Ixp25_ASAP7_75t_L g185 ( 
.A1(n_167),
.A2(n_146),
.B(n_139),
.C(n_141),
.D(n_132),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_185),
.B(n_157),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_159),
.B(n_136),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_186),
.B(n_163),
.Y(n_199)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_167),
.B(n_158),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_187),
.B(n_154),
.C(n_160),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_155),
.Y(n_188)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_189),
.Y(n_204)
);

BUFx2_ASAP7_75t_L g190 ( 
.A(n_156),
.Y(n_190)
);

CKINVDCx14_ASAP7_75t_R g207 ( 
.A(n_190),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_176),
.Y(n_191)
);

CKINVDCx14_ASAP7_75t_R g208 ( 
.A(n_191),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_SL g192 ( 
.A(n_174),
.B(n_124),
.Y(n_192)
);

CKINVDCx16_ASAP7_75t_R g210 ( 
.A(n_192),
.Y(n_210)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_170),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_194),
.B(n_156),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_152),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_199),
.B(n_205),
.Y(n_222)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_201),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_179),
.A2(n_175),
.B1(n_166),
.B2(n_173),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_203),
.A2(n_190),
.B1(n_177),
.B2(n_153),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_189),
.B(n_164),
.Y(n_206)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_206),
.Y(n_221)
);

A2O1A1Ixp33_ASAP7_75t_SL g216 ( 
.A1(n_209),
.A2(n_195),
.B(n_162),
.C(n_183),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_211),
.B(n_212),
.Y(n_213)
);

XOR2x2_ASAP7_75t_L g212 ( 
.A(n_187),
.B(n_162),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_212),
.B(n_186),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_SL g229 ( 
.A(n_215),
.B(n_205),
.Y(n_229)
);

A2O1A1Ixp33_ASAP7_75t_SL g234 ( 
.A1(n_216),
.A2(n_171),
.B(n_152),
.C(n_123),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_211),
.B(n_183),
.C(n_195),
.Y(n_217)
);

AND2x2_ASAP7_75t_L g233 ( 
.A(n_217),
.B(n_153),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_L g218 ( 
.A1(n_210),
.A2(n_179),
.B1(n_193),
.B2(n_177),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_218),
.A2(n_204),
.B1(n_197),
.B2(n_202),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_208),
.B(n_200),
.Y(n_219)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_219),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_199),
.B(n_194),
.Y(n_220)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_220),
.Y(n_235)
);

OAI21xp5_ASAP7_75t_SL g223 ( 
.A1(n_206),
.A2(n_204),
.B(n_198),
.Y(n_223)
);

CKINVDCx14_ASAP7_75t_R g231 ( 
.A(n_223),
.Y(n_231)
);

INVx13_ASAP7_75t_L g224 ( 
.A(n_207),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_224),
.B(n_201),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_225),
.A2(n_169),
.B1(n_168),
.B2(n_197),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_227),
.B(n_232),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_228),
.A2(n_214),
.B1(n_215),
.B2(n_216),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_229),
.B(n_233),
.C(n_213),
.Y(n_236)
);

OA22x2_ASAP7_75t_L g230 ( 
.A1(n_221),
.A2(n_209),
.B1(n_185),
.B2(n_202),
.Y(n_230)
);

CKINVDCx16_ASAP7_75t_R g240 ( 
.A(n_230),
.Y(n_240)
);

INVxp67_ASAP7_75t_L g237 ( 
.A(n_234),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_236),
.B(n_235),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_231),
.B(n_222),
.C(n_213),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_238),
.B(n_241),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_239),
.A2(n_234),
.B1(n_216),
.B2(n_230),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_231),
.B(n_222),
.C(n_217),
.Y(n_241)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_242),
.Y(n_243)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_243),
.Y(n_248)
);

AOI21xp5_ASAP7_75t_L g251 ( 
.A1(n_244),
.A2(n_247),
.B(n_246),
.Y(n_251)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_246),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_240),
.B(n_226),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_L g249 ( 
.A1(n_245),
.A2(n_237),
.B(n_232),
.Y(n_249)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_249),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_251),
.B(n_244),
.Y(n_254)
);

NOR2xp67_ASAP7_75t_L g252 ( 
.A(n_248),
.B(n_250),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_252),
.B(n_254),
.C(n_237),
.Y(n_255)
);

AO21x1_ASAP7_75t_L g256 ( 
.A1(n_255),
.A2(n_253),
.B(n_234),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_256),
.B(n_216),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_257),
.B(n_224),
.Y(n_258)
);


endmodule