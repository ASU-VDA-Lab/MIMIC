module fake_jpeg_30378_n_61 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_61);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_61;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_23;
wire n_10;
wire n_27;
wire n_55;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_59;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_44;
wire n_26;
wire n_38;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_31;
wire n_25;
wire n_56;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;

BUFx6f_ASAP7_75t_L g8 ( 
.A(n_3),
.Y(n_8)
);

INVx1_ASAP7_75t_L g9 ( 
.A(n_4),
.Y(n_9)
);

BUFx3_ASAP7_75t_L g10 ( 
.A(n_2),
.Y(n_10)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_0),
.Y(n_11)
);

BUFx5_ASAP7_75t_L g12 ( 
.A(n_3),
.Y(n_12)
);

BUFx10_ASAP7_75t_L g13 ( 
.A(n_1),
.Y(n_13)
);

INVx2_ASAP7_75t_L g14 ( 
.A(n_5),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_2),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_7),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_17),
.B(n_6),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_18),
.B(n_20),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_19),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_17),
.B(n_6),
.Y(n_20)
);

OR2x2_ASAP7_75t_L g21 ( 
.A(n_16),
.B(n_0),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_21),
.B(n_23),
.Y(n_26)
);

BUFx10_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

OR2x2_ASAP7_75t_L g31 ( 
.A(n_22),
.B(n_12),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_13),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_14),
.B(n_0),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_24),
.B(n_14),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_SL g38 ( 
.A(n_27),
.B(n_28),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_21),
.B(n_9),
.Y(n_28)
);

OAI21xp5_ASAP7_75t_SL g29 ( 
.A1(n_24),
.A2(n_9),
.B(n_11),
.Y(n_29)
);

CKINVDCx16_ASAP7_75t_R g39 ( 
.A(n_29),
.Y(n_39)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_31),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_L g33 ( 
.A1(n_27),
.A2(n_23),
.B1(n_8),
.B2(n_15),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_L g41 ( 
.A1(n_33),
.A2(n_35),
.B1(n_12),
.B2(n_10),
.Y(n_41)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_30),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_34),
.B(n_37),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_L g35 ( 
.A1(n_29),
.A2(n_19),
.B1(n_11),
.B2(n_15),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_26),
.B(n_31),
.Y(n_36)
);

XNOR2xp5_ASAP7_75t_L g44 ( 
.A(n_36),
.B(n_22),
.Y(n_44)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_30),
.Y(n_37)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

NAND3xp33_ASAP7_75t_L g42 ( 
.A(n_40),
.B(n_25),
.C(n_2),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_L g48 ( 
.A1(n_41),
.A2(n_43),
.B1(n_32),
.B2(n_33),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_42),
.Y(n_51)
);

HB1xp67_ASAP7_75t_SL g43 ( 
.A(n_39),
.Y(n_43)
);

XNOR2xp5_ASAP7_75t_L g49 ( 
.A(n_44),
.B(n_38),
.Y(n_49)
);

AND2x6_ASAP7_75t_L g46 ( 
.A(n_36),
.B(n_22),
.Y(n_46)
);

MAJIxp5_ASAP7_75t_L g47 ( 
.A(n_46),
.B(n_40),
.C(n_32),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_47),
.B(n_50),
.Y(n_53)
);

OAI21xp5_ASAP7_75t_L g54 ( 
.A1(n_48),
.A2(n_19),
.B(n_10),
.Y(n_54)
);

MAJIxp5_ASAP7_75t_L g52 ( 
.A(n_49),
.B(n_46),
.C(n_42),
.Y(n_52)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_45),
.Y(n_50)
);

XOR2xp5_ASAP7_75t_L g56 ( 
.A(n_52),
.B(n_54),
.Y(n_56)
);

OAI322xp33_ASAP7_75t_L g55 ( 
.A1(n_53),
.A2(n_51),
.A3(n_49),
.B1(n_47),
.B2(n_13),
.C1(n_7),
.C2(n_37),
.Y(n_55)
);

MAJIxp5_ASAP7_75t_L g57 ( 
.A(n_55),
.B(n_34),
.C(n_3),
.Y(n_57)
);

OAI21xp5_ASAP7_75t_L g59 ( 
.A1(n_57),
.A2(n_58),
.B(n_1),
.Y(n_59)
);

MAJIxp5_ASAP7_75t_L g58 ( 
.A(n_56),
.B(n_22),
.C(n_13),
.Y(n_58)
);

OAI21xp5_ASAP7_75t_SL g60 ( 
.A1(n_59),
.A2(n_1),
.B(n_4),
.Y(n_60)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_60),
.B(n_4),
.Y(n_61)
);


endmodule