module fake_jpeg_8864_n_298 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_298);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_298;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_155;
wire n_207;
wire n_277;
wire n_31;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_21;
wire n_57;
wire n_187;
wire n_234;
wire n_288;
wire n_272;
wire n_284;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_247;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_145;
wire n_241;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_273;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_270;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_265;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

INVx1_ASAP7_75t_L g17 ( 
.A(n_14),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_14),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

INVx6_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_10),
.Y(n_26)
);

CKINVDCx16_ASAP7_75t_R g27 ( 
.A(n_9),
.Y(n_27)
);

BUFx24_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_1),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_15),
.B(n_8),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_16),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_3),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_10),
.Y(n_35)
);

INVx2_ASAP7_75t_SL g36 ( 
.A(n_24),
.Y(n_36)
);

NAND2x2_ASAP7_75t_L g47 ( 
.A(n_36),
.B(n_28),
.Y(n_47)
);

INVx5_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_37),
.Y(n_61)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_24),
.Y(n_38)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_38),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_22),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_39),
.B(n_35),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_19),
.B(n_0),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_40),
.B(n_45),
.Y(n_52)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_32),
.Y(n_41)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_41),
.Y(n_63)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

AND2x2_ASAP7_75t_L g51 ( 
.A(n_42),
.B(n_43),
.Y(n_51)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_28),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_19),
.B(n_0),
.Y(n_44)
);

OR2x2_ASAP7_75t_L g46 ( 
.A(n_44),
.B(n_24),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_21),
.B(n_0),
.Y(n_45)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_46),
.B(n_72),
.Y(n_91)
);

INVx1_ASAP7_75t_SL g90 ( 
.A(n_47),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_44),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_48),
.B(n_49),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_41),
.B(n_42),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_39),
.Y(n_50)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_50),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_L g53 ( 
.A1(n_40),
.A2(n_22),
.B1(n_21),
.B2(n_45),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_L g78 ( 
.A1(n_53),
.A2(n_64),
.B1(n_65),
.B2(n_23),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_54),
.Y(n_73)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_55),
.Y(n_74)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_56),
.B(n_57),
.Y(n_83)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_44),
.Y(n_58)
);

AOI21xp33_ASAP7_75t_L g87 ( 
.A1(n_58),
.A2(n_51),
.B(n_69),
.Y(n_87)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_37),
.Y(n_59)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_59),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_41),
.B(n_26),
.Y(n_60)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_60),
.Y(n_93)
);

BUFx12_ASAP7_75t_L g62 ( 
.A(n_38),
.Y(n_62)
);

CKINVDCx14_ASAP7_75t_R g75 ( 
.A(n_62),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_L g64 ( 
.A1(n_40),
.A2(n_22),
.B1(n_33),
.B2(n_18),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_40),
.A2(n_45),
.B1(n_42),
.B2(n_41),
.Y(n_65)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_36),
.Y(n_66)
);

INVx5_ASAP7_75t_L g89 ( 
.A(n_66),
.Y(n_89)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_37),
.Y(n_67)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_67),
.Y(n_80)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_37),
.Y(n_68)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_68),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_45),
.B(n_23),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_69),
.B(n_71),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_42),
.B(n_26),
.Y(n_71)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_47),
.Y(n_77)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_77),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_78),
.B(n_86),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_48),
.A2(n_58),
.B1(n_63),
.B2(n_27),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_79),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_L g81 ( 
.A1(n_63),
.A2(n_36),
.B1(n_33),
.B2(n_18),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_81),
.A2(n_29),
.B1(n_17),
.B2(n_30),
.Y(n_98)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_62),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g111 ( 
.A(n_87),
.B(n_43),
.Y(n_111)
);

AND2x6_ASAP7_75t_L g88 ( 
.A(n_51),
.B(n_16),
.Y(n_88)
);

AND2x6_ASAP7_75t_L g109 ( 
.A(n_88),
.B(n_11),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_50),
.Y(n_94)
);

INVx6_ASAP7_75t_L g118 ( 
.A(n_94),
.Y(n_118)
);

BUFx12_ASAP7_75t_L g95 ( 
.A(n_47),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_95),
.B(n_47),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_90),
.B(n_52),
.C(n_65),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_97),
.B(n_100),
.C(n_43),
.Y(n_123)
);

CKINVDCx16_ASAP7_75t_R g147 ( 
.A(n_98),
.Y(n_147)
);

INVx1_ASAP7_75t_SL g99 ( 
.A(n_74),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_99),
.B(n_102),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_90),
.B(n_52),
.C(n_92),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_76),
.B(n_51),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_101),
.B(n_103),
.Y(n_142)
);

INVx13_ASAP7_75t_L g102 ( 
.A(n_75),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_91),
.B(n_46),
.Y(n_103)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_83),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_104),
.B(n_113),
.Y(n_129)
);

BUFx24_ASAP7_75t_L g105 ( 
.A(n_80),
.Y(n_105)
);

BUFx3_ASAP7_75t_L g140 ( 
.A(n_105),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_77),
.A2(n_56),
.B1(n_70),
.B2(n_47),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_106),
.A2(n_61),
.B1(n_37),
.B2(n_43),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_91),
.B(n_54),
.Y(n_107)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_107),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_109),
.A2(n_17),
.B1(n_61),
.B2(n_27),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_L g126 ( 
.A1(n_111),
.A2(n_85),
.B(n_29),
.Y(n_126)
);

AOI21xp5_ASAP7_75t_L g146 ( 
.A1(n_112),
.A2(n_28),
.B(n_36),
.Y(n_146)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_91),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_93),
.B(n_62),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_114),
.B(n_115),
.Y(n_132)
);

INVx13_ASAP7_75t_L g115 ( 
.A(n_86),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_92),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_116),
.B(n_117),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_74),
.B(n_57),
.Y(n_117)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_89),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_119),
.B(n_121),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_88),
.B(n_68),
.Y(n_120)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_120),
.Y(n_127)
);

INVx13_ASAP7_75t_L g121 ( 
.A(n_80),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_123),
.B(n_25),
.C(n_35),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_125),
.A2(n_128),
.B1(n_135),
.B2(n_143),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_L g150 ( 
.A1(n_126),
.A2(n_144),
.B(n_108),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_96),
.A2(n_95),
.B1(n_59),
.B2(n_67),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_101),
.B(n_95),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g167 ( 
.A(n_130),
.B(n_16),
.Y(n_167)
);

INVx4_ASAP7_75t_L g131 ( 
.A(n_99),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_131),
.B(n_134),
.Y(n_153)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_107),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_133),
.B(n_116),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_120),
.A2(n_73),
.B1(n_84),
.B2(n_70),
.Y(n_135)
);

INVxp33_ASAP7_75t_L g137 ( 
.A(n_119),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_137),
.B(n_141),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_110),
.A2(n_84),
.B1(n_73),
.B2(n_82),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_L g161 ( 
.A1(n_138),
.A2(n_148),
.B(n_28),
.Y(n_161)
);

INVxp33_ASAP7_75t_L g141 ( 
.A(n_121),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_113),
.A2(n_55),
.B1(n_36),
.B2(n_66),
.Y(n_143)
);

AND2x2_ASAP7_75t_SL g144 ( 
.A(n_103),
.B(n_111),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_L g145 ( 
.A1(n_110),
.A2(n_89),
.B1(n_82),
.B2(n_36),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_145),
.A2(n_115),
.B1(n_94),
.B2(n_105),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_SL g160 ( 
.A1(n_146),
.A2(n_108),
.B(n_106),
.Y(n_160)
);

AND2x2_ASAP7_75t_L g148 ( 
.A(n_97),
.B(n_0),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_150),
.B(n_169),
.Y(n_203)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_139),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_151),
.B(n_154),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_SL g152 ( 
.A(n_144),
.B(n_111),
.Y(n_152)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_152),
.B(n_148),
.Y(n_193)
);

CKINVDCx16_ASAP7_75t_R g154 ( 
.A(n_139),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_L g155 ( 
.A(n_123),
.B(n_100),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_155),
.B(n_168),
.C(n_174),
.Y(n_178)
);

CKINVDCx16_ASAP7_75t_R g156 ( 
.A(n_136),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_156),
.B(n_164),
.Y(n_180)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_157),
.Y(n_184)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_136),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_158),
.B(n_162),
.Y(n_182)
);

XOR2x2_ASAP7_75t_SL g201 ( 
.A(n_160),
.B(n_146),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_161),
.A2(n_163),
.B1(n_165),
.B2(n_166),
.Y(n_198)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_124),
.Y(n_162)
);

AOI21xp5_ASAP7_75t_L g163 ( 
.A1(n_127),
.A2(n_109),
.B(n_104),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_124),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_147),
.A2(n_102),
.B1(n_98),
.B2(n_118),
.Y(n_165)
);

AOI21xp5_ASAP7_75t_L g166 ( 
.A1(n_127),
.A2(n_130),
.B(n_133),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_167),
.B(n_170),
.Y(n_199)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_144),
.B(n_102),
.Y(n_168)
);

AOI21xp5_ASAP7_75t_L g169 ( 
.A1(n_122),
.A2(n_105),
.B(n_118),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_145),
.Y(n_170)
);

CKINVDCx16_ASAP7_75t_R g171 ( 
.A(n_132),
.Y(n_171)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_171),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_172),
.Y(n_190)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_143),
.Y(n_173)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_173),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_144),
.B(n_25),
.Y(n_174)
);

OR2x2_ASAP7_75t_L g175 ( 
.A(n_129),
.B(n_30),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_175),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_SL g176 ( 
.A(n_142),
.B(n_12),
.Y(n_176)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_176),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_177),
.B(n_160),
.C(n_161),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_159),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_SL g206 ( 
.A(n_183),
.B(n_156),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_185),
.B(n_186),
.C(n_188),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_155),
.B(n_122),
.C(n_142),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_152),
.B(n_126),
.C(n_148),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_173),
.A2(n_134),
.B1(n_147),
.B2(n_135),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_192),
.A2(n_202),
.B1(n_171),
.B2(n_131),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_193),
.B(n_158),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_153),
.A2(n_170),
.B1(n_125),
.B2(n_166),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_194),
.A2(n_149),
.B1(n_165),
.B2(n_164),
.Y(n_207)
);

BUFx6f_ASAP7_75t_L g195 ( 
.A(n_151),
.Y(n_195)
);

BUFx6f_ASAP7_75t_L g226 ( 
.A(n_195),
.Y(n_226)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_169),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_196),
.B(n_197),
.Y(n_223)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_172),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_168),
.B(n_129),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_200),
.B(n_177),
.C(n_174),
.Y(n_208)
);

AO21x1_ASAP7_75t_L g221 ( 
.A1(n_201),
.A2(n_181),
.B(n_198),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_149),
.A2(n_128),
.B1(n_138),
.B2(n_132),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_SL g205 ( 
.A(n_203),
.B(n_150),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_SL g244 ( 
.A(n_205),
.B(n_215),
.Y(n_244)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_206),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_207),
.A2(n_225),
.B1(n_190),
.B2(n_184),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_208),
.B(n_213),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_178),
.B(n_163),
.C(n_148),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_209),
.B(n_214),
.C(n_219),
.Y(n_238)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_182),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_210),
.B(n_211),
.Y(n_237)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_182),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_180),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_SL g228 ( 
.A1(n_212),
.A2(n_217),
.B(n_218),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_178),
.B(n_162),
.Y(n_214)
);

FAx1_ASAP7_75t_SL g215 ( 
.A(n_201),
.B(n_167),
.CI(n_176),
.CON(n_215),
.SN(n_215)
);

OAI21xp5_ASAP7_75t_L g229 ( 
.A1(n_216),
.A2(n_185),
.B(n_189),
.Y(n_229)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_191),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_199),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_186),
.B(n_140),
.C(n_131),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_203),
.B(n_200),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_220),
.B(n_193),
.Y(n_239)
);

NAND3xp33_ASAP7_75t_L g234 ( 
.A(n_221),
.B(n_215),
.C(n_184),
.Y(n_234)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_194),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_SL g241 ( 
.A1(n_222),
.A2(n_189),
.B(n_179),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_202),
.A2(n_175),
.B1(n_140),
.B2(n_105),
.Y(n_224)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_224),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_190),
.A2(n_175),
.B1(n_35),
.B2(n_34),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_227),
.B(n_236),
.Y(n_255)
);

AOI21xp5_ASAP7_75t_L g248 ( 
.A1(n_229),
.A2(n_241),
.B(n_195),
.Y(n_248)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_223),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_232),
.B(n_235),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_216),
.A2(n_192),
.B1(n_205),
.B2(n_224),
.Y(n_233)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_233),
.Y(n_253)
);

OAI21xp5_ASAP7_75t_L g254 ( 
.A1(n_234),
.A2(n_25),
.B(n_2),
.Y(n_254)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_226),
.Y(n_235)
);

BUFx12_ASAP7_75t_L g236 ( 
.A(n_226),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_239),
.B(n_245),
.Y(n_247)
);

BUFx2_ASAP7_75t_L g240 ( 
.A(n_221),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_240),
.B(n_243),
.Y(n_256)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_219),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_214),
.B(n_188),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_231),
.A2(n_209),
.B1(n_204),
.B2(n_208),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_246),
.B(n_250),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_248),
.B(n_244),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_238),
.B(n_204),
.C(n_220),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_249),
.B(n_251),
.C(n_34),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_229),
.A2(n_213),
.B1(n_215),
.B2(n_187),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_238),
.B(n_242),
.C(n_239),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_245),
.B(n_242),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_252),
.B(n_244),
.C(n_228),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_254),
.Y(n_265)
);

OA21x2_ASAP7_75t_L g258 ( 
.A1(n_240),
.A2(n_140),
.B(n_35),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_258),
.B(n_259),
.Y(n_268)
);

AOI21xp5_ASAP7_75t_L g259 ( 
.A1(n_237),
.A2(n_1),
.B(n_2),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_257),
.B(n_230),
.Y(n_260)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_260),
.Y(n_279)
);

AND2x2_ASAP7_75t_L g261 ( 
.A(n_253),
.B(n_234),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_261),
.B(n_263),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_262),
.B(n_246),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_SL g263 ( 
.A(n_259),
.B(n_236),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_266),
.B(n_252),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_251),
.B(n_236),
.C(n_4),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_267),
.B(n_270),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_269),
.B(n_248),
.C(n_256),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_256),
.B(n_11),
.Y(n_270)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_273),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_L g274 ( 
.A1(n_264),
.A2(n_249),
.B(n_255),
.Y(n_274)
);

AOI21xp5_ASAP7_75t_SL g282 ( 
.A1(n_274),
.A2(n_261),
.B(n_271),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_SL g284 ( 
.A(n_275),
.B(n_276),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_268),
.A2(n_250),
.B1(n_258),
.B2(n_254),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_SL g281 ( 
.A(n_277),
.B(n_247),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_269),
.B(n_247),
.C(n_258),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_SL g286 ( 
.A(n_278),
.B(n_34),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_SL g288 ( 
.A(n_281),
.B(n_12),
.Y(n_288)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_282),
.Y(n_291)
);

OAI21x1_ASAP7_75t_L g283 ( 
.A1(n_278),
.A2(n_265),
.B(n_268),
.Y(n_283)
);

AOI332xp33_ASAP7_75t_L g289 ( 
.A1(n_283),
.A2(n_285),
.A3(n_9),
.B1(n_5),
.B2(n_6),
.B3(n_7),
.C1(n_8),
.C2(n_15),
.Y(n_289)
);

AOI21x1_ASAP7_75t_L g285 ( 
.A1(n_273),
.A2(n_11),
.B(n_5),
.Y(n_285)
);

AOI322xp5_ASAP7_75t_L g287 ( 
.A1(n_286),
.A2(n_279),
.A3(n_272),
.B1(n_275),
.B2(n_7),
.C1(n_8),
.C2(n_9),
.Y(n_287)
);

AOI322xp5_ASAP7_75t_L g293 ( 
.A1(n_287),
.A2(n_290),
.A3(n_1),
.B1(n_6),
.B2(n_20),
.C1(n_31),
.C2(n_291),
.Y(n_293)
);

AOI221xp5_ASAP7_75t_L g292 ( 
.A1(n_288),
.A2(n_5),
.B1(n_6),
.B2(n_13),
.C(n_280),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_L g294 ( 
.A1(n_289),
.A2(n_20),
.B1(n_31),
.B2(n_179),
.Y(n_294)
);

AOI322xp5_ASAP7_75t_L g290 ( 
.A1(n_284),
.A2(n_34),
.A3(n_31),
.B1(n_20),
.B2(n_7),
.C1(n_13),
.C2(n_15),
.Y(n_290)
);

INVxp67_ASAP7_75t_L g296 ( 
.A(n_292),
.Y(n_296)
);

AND2x2_ASAP7_75t_L g295 ( 
.A(n_293),
.B(n_294),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_295),
.B(n_20),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_297),
.B(n_296),
.Y(n_298)
);


endmodule