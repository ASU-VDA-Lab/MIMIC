module real_aes_4642_n_7 (n_4, n_0, n_3, n_5, n_2, n_6, n_1, n_7);
input n_4;
input n_0;
input n_3;
input n_5;
input n_2;
input n_6;
input n_1;
output n_7;
wire n_13;
wire n_15;
wire n_8;
wire n_9;
wire n_12;
wire n_14;
wire n_10;
wire n_11;
A2O1A1Ixp33_ASAP7_75t_SL g7 ( .A1(n_0), .A2(n_8), .B(n_11), .C(n_14), .Y(n_7) );
NOR2xp33_ASAP7_75t_L g8 ( .A(n_1), .B(n_9), .Y(n_8) );
INVx1_ASAP7_75t_L g12 ( .A(n_2), .Y(n_12) );
AND2x2_ASAP7_75t_L g14 ( .A(n_3), .B(n_15), .Y(n_14) );
O2A1O1Ixp33_ASAP7_75t_L g11 ( .A1(n_4), .A2(n_8), .B(n_12), .C(n_13), .Y(n_11) );
NAND2xp5_ASAP7_75t_L g13 ( .A(n_4), .B(n_12), .Y(n_13) );
BUFx3_ASAP7_75t_L g10 ( .A(n_5), .Y(n_10) );
INVx1_ASAP7_75t_L g15 ( .A(n_6), .Y(n_15) );
CKINVDCx20_ASAP7_75t_R g9 ( .A(n_10), .Y(n_9) );
endmodule