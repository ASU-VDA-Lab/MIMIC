module fake_jpeg_8532_n_333 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_333);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_333;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx8_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_12),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_10),
.B(n_7),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

INVxp67_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_4),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

INVx11_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_37),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_23),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_39),
.B(n_41),
.Y(n_57)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_16),
.Y(n_40)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_40),
.Y(n_59)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_26),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_24),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_42),
.B(n_45),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g43 ( 
.A(n_29),
.B(n_8),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_43),
.B(n_44),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_24),
.B(n_0),
.Y(n_44)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_17),
.Y(n_45)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_16),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_46),
.Y(n_71)
);

BUFx16f_ASAP7_75t_L g47 ( 
.A(n_37),
.Y(n_47)
);

INVx3_ASAP7_75t_SL g109 ( 
.A(n_47),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_L g48 ( 
.A1(n_42),
.A2(n_25),
.B1(n_44),
.B2(n_27),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_48),
.A2(n_19),
.B1(n_22),
.B2(n_28),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_44),
.B(n_25),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_49),
.B(n_50),
.Y(n_76)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_42),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

CKINVDCx16_ASAP7_75t_R g102 ( 
.A(n_51),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_43),
.B(n_21),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_53),
.B(n_56),
.Y(n_95)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_55),
.Y(n_93)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_36),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_37),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_58),
.B(n_63),
.Y(n_94)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_36),
.Y(n_60)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_60),
.B(n_62),
.Y(n_107)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_36),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_37),
.Y(n_63)
);

INVx6_ASAP7_75t_SL g64 ( 
.A(n_40),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_64),
.B(n_65),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_43),
.B(n_21),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_36),
.B(n_19),
.Y(n_66)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_66),
.Y(n_75)
);

CKINVDCx14_ASAP7_75t_R g67 ( 
.A(n_38),
.Y(n_67)
);

OR2x2_ASAP7_75t_L g88 ( 
.A(n_67),
.B(n_46),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_38),
.B(n_18),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_69),
.B(n_40),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_37),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_72),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g73 ( 
.A(n_64),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_73),
.B(n_77),
.Y(n_126)
);

OAI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_74),
.A2(n_81),
.B1(n_86),
.B2(n_88),
.Y(n_121)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_66),
.Y(n_77)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_57),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_79),
.B(n_82),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_49),
.A2(n_39),
.B1(n_27),
.B2(n_35),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_L g83 ( 
.A1(n_53),
.A2(n_39),
.B1(n_40),
.B2(n_22),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_83),
.A2(n_90),
.B1(n_96),
.B2(n_18),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_68),
.A2(n_31),
.B1(n_39),
.B2(n_28),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_84),
.Y(n_123)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_57),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_85),
.B(n_87),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_65),
.A2(n_35),
.B1(n_33),
.B2(n_34),
.Y(n_86)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_54),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_70),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_89),
.B(n_71),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_69),
.A2(n_34),
.B1(n_33),
.B2(n_30),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_59),
.A2(n_46),
.B1(n_30),
.B2(n_45),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_91),
.Y(n_130)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_54),
.Y(n_92)
);

CKINVDCx16_ASAP7_75t_R g119 ( 
.A(n_92),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_L g96 ( 
.A1(n_50),
.A2(n_46),
.B1(n_41),
.B2(n_45),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_70),
.A2(n_45),
.B1(n_41),
.B2(n_31),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_97),
.A2(n_103),
.B1(n_52),
.B2(n_62),
.Y(n_117)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_47),
.Y(n_98)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_98),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_51),
.Y(n_99)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_99),
.Y(n_116)
);

INVx5_ASAP7_75t_L g100 ( 
.A(n_47),
.Y(n_100)
);

INVx5_ASAP7_75t_L g131 ( 
.A(n_100),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_59),
.B(n_20),
.Y(n_101)
);

CKINVDCx16_ASAP7_75t_R g124 ( 
.A(n_101),
.Y(n_124)
);

OAI22xp33_ASAP7_75t_L g103 ( 
.A1(n_52),
.A2(n_38),
.B1(n_23),
.B2(n_32),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_47),
.Y(n_104)
);

CKINVDCx16_ASAP7_75t_R g134 ( 
.A(n_104),
.Y(n_134)
);

NAND2x1p5_ASAP7_75t_L g105 ( 
.A(n_68),
.B(n_16),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g138 ( 
.A(n_105),
.B(n_0),
.Y(n_138)
);

BUFx2_ASAP7_75t_L g106 ( 
.A(n_71),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_106),
.Y(n_111)
);

O2A1O1Ixp33_ASAP7_75t_L g108 ( 
.A1(n_58),
.A2(n_38),
.B(n_16),
.C(n_20),
.Y(n_108)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_108),
.Y(n_136)
);

BUFx3_ASAP7_75t_L g110 ( 
.A(n_55),
.Y(n_110)
);

INVx2_ASAP7_75t_SL g122 ( 
.A(n_110),
.Y(n_122)
);

XOR2xp5_ASAP7_75t_L g113 ( 
.A(n_76),
.B(n_18),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_113),
.B(n_128),
.C(n_140),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_106),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_115),
.B(n_120),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_117),
.A2(n_118),
.B1(n_135),
.B2(n_108),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_76),
.A2(n_60),
.B1(n_56),
.B2(n_63),
.Y(n_118)
);

INVx8_ASAP7_75t_L g125 ( 
.A(n_109),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_125),
.A2(n_100),
.B1(n_109),
.B2(n_93),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_84),
.A2(n_71),
.B1(n_17),
.B2(n_32),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_127),
.A2(n_73),
.B1(n_77),
.B2(n_75),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_L g128 ( 
.A(n_105),
.B(n_95),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g169 ( 
.A(n_129),
.B(n_0),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_95),
.B(n_72),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_132),
.B(n_139),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_89),
.A2(n_32),
.B1(n_20),
.B2(n_18),
.Y(n_135)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_107),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_137),
.B(n_103),
.Y(n_158)
);

AOI21xp5_ASAP7_75t_L g152 ( 
.A1(n_138),
.A2(n_107),
.B(n_80),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_105),
.B(n_72),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_94),
.B(n_55),
.C(n_51),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_129),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_141),
.B(n_142),
.Y(n_176)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_133),
.Y(n_142)
);

BUFx3_ASAP7_75t_L g144 ( 
.A(n_122),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_144),
.B(n_146),
.Y(n_181)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_132),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_122),
.B(n_85),
.Y(n_147)
);

CKINVDCx16_ASAP7_75t_R g202 ( 
.A(n_147),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_148),
.A2(n_153),
.B1(n_163),
.B2(n_125),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_128),
.B(n_79),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_149),
.B(n_155),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_118),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_150),
.B(n_154),
.Y(n_190)
);

OA21x2_ASAP7_75t_L g151 ( 
.A1(n_136),
.A2(n_107),
.B(n_75),
.Y(n_151)
);

OA21x2_ASAP7_75t_L g175 ( 
.A1(n_151),
.A2(n_135),
.B(n_112),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_L g200 ( 
.A1(n_152),
.A2(n_161),
.B(n_164),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_123),
.A2(n_97),
.B1(n_87),
.B2(n_92),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_122),
.B(n_93),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_113),
.B(n_88),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_156),
.B(n_131),
.Y(n_191)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_116),
.Y(n_157)
);

HB1xp67_ASAP7_75t_L g207 ( 
.A(n_157),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_SL g185 ( 
.A(n_158),
.B(n_173),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_139),
.B(n_98),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_159),
.B(n_162),
.Y(n_188)
);

INVxp67_ASAP7_75t_L g196 ( 
.A(n_160),
.Y(n_196)
);

AND2x2_ASAP7_75t_L g161 ( 
.A(n_137),
.B(n_109),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_138),
.B(n_104),
.Y(n_162)
);

O2A1O1Ixp33_ASAP7_75t_L g163 ( 
.A1(n_136),
.A2(n_106),
.B(n_32),
.C(n_51),
.Y(n_163)
);

AND2x2_ASAP7_75t_L g164 ( 
.A(n_140),
.B(n_0),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_123),
.A2(n_130),
.B1(n_117),
.B2(n_114),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_165),
.A2(n_171),
.B1(n_131),
.B2(n_115),
.Y(n_179)
);

OAI32xp33_ASAP7_75t_L g167 ( 
.A1(n_120),
.A2(n_102),
.A3(n_20),
.B1(n_12),
.B2(n_15),
.Y(n_167)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_167),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_138),
.B(n_61),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_168),
.B(n_169),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_127),
.B(n_61),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_170),
.B(n_134),
.C(n_111),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_130),
.A2(n_61),
.B1(n_78),
.B2(n_11),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_121),
.B(n_1),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_172),
.B(n_151),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_SL g173 ( 
.A(n_126),
.B(n_10),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_124),
.B(n_99),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_SL g186 ( 
.A(n_174),
.B(n_141),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_SL g232 ( 
.A1(n_175),
.A2(n_179),
.B(n_164),
.Y(n_232)
);

AND2x6_ASAP7_75t_L g177 ( 
.A(n_166),
.B(n_124),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_177),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_178),
.A2(n_191),
.B1(n_201),
.B2(n_198),
.Y(n_235)
);

AND2x2_ASAP7_75t_SL g183 ( 
.A(n_159),
.B(n_112),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_L g234 ( 
.A1(n_183),
.A2(n_157),
.B(n_2),
.Y(n_234)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_163),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_184),
.B(n_186),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_166),
.B(n_134),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_187),
.B(n_193),
.C(n_197),
.Y(n_214)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_145),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_189),
.B(n_192),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_169),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_SL g194 ( 
.A(n_152),
.B(n_13),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_194),
.B(n_198),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_149),
.B(n_111),
.C(n_119),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_142),
.B(n_116),
.Y(n_199)
);

CKINVDCx16_ASAP7_75t_R g209 ( 
.A(n_199),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_143),
.A2(n_78),
.B1(n_110),
.B2(n_99),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_146),
.B(n_1),
.Y(n_203)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_203),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_144),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_204),
.B(n_205),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_150),
.B(n_9),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_145),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_206),
.B(n_173),
.Y(n_217)
);

O2A1O1Ixp33_ASAP7_75t_SL g208 ( 
.A1(n_184),
.A2(n_172),
.B(n_151),
.C(n_168),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_SL g241 ( 
.A1(n_208),
.A2(n_225),
.B(n_226),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_180),
.A2(n_165),
.B1(n_167),
.B2(n_156),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_210),
.A2(n_221),
.B1(n_185),
.B2(n_78),
.Y(n_257)
);

AOI21xp5_ASAP7_75t_L g213 ( 
.A1(n_196),
.A2(n_161),
.B(n_162),
.Y(n_213)
);

A2O1A1Ixp33_ASAP7_75t_SL g258 ( 
.A1(n_213),
.A2(n_219),
.B(n_235),
.C(n_1),
.Y(n_258)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_207),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_215),
.B(n_220),
.Y(n_249)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_217),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_182),
.B(n_155),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_218),
.B(n_222),
.C(n_200),
.Y(n_248)
);

OA21x2_ASAP7_75t_L g219 ( 
.A1(n_180),
.A2(n_175),
.B(n_183),
.Y(n_219)
);

INVx5_ASAP7_75t_L g220 ( 
.A(n_204),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_196),
.A2(n_175),
.B1(n_202),
.B2(n_179),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_187),
.B(n_170),
.C(n_161),
.Y(n_222)
);

INVxp67_ASAP7_75t_L g223 ( 
.A(n_201),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_223),
.B(n_229),
.Y(n_243)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_181),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_176),
.Y(n_226)
);

NOR3xp33_ASAP7_75t_L g227 ( 
.A(n_194),
.B(n_164),
.C(n_171),
.Y(n_227)
);

NAND3xp33_ASAP7_75t_L g251 ( 
.A(n_227),
.B(n_188),
.C(n_195),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_186),
.B(n_11),
.Y(n_228)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_228),
.Y(n_238)
);

INVxp67_ASAP7_75t_L g229 ( 
.A(n_190),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_183),
.Y(n_230)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_230),
.Y(n_240)
);

CKINVDCx16_ASAP7_75t_R g255 ( 
.A(n_232),
.Y(n_255)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_234),
.Y(n_250)
);

AND2x2_ASAP7_75t_L g236 ( 
.A(n_230),
.B(n_193),
.Y(n_236)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_236),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_223),
.A2(n_206),
.B1(n_189),
.B2(n_177),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_239),
.A2(n_246),
.B1(n_224),
.B2(n_229),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_SL g242 ( 
.A(n_226),
.B(n_192),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_242),
.B(n_259),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_214),
.B(n_182),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_244),
.B(n_248),
.C(n_253),
.Y(n_264)
);

AND2x2_ASAP7_75t_L g245 ( 
.A(n_231),
.B(n_183),
.Y(n_245)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_245),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_216),
.A2(n_175),
.B1(n_202),
.B2(n_178),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_216),
.A2(n_210),
.B1(n_221),
.B2(n_219),
.Y(n_247)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_247),
.Y(n_263)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_251),
.Y(n_267)
);

CKINVDCx11_ASAP7_75t_R g252 ( 
.A(n_220),
.Y(n_252)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_252),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_214),
.B(n_197),
.C(n_200),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_222),
.B(n_188),
.C(n_195),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_254),
.B(n_256),
.C(n_224),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_218),
.B(n_203),
.C(n_185),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_L g265 ( 
.A1(n_257),
.A2(n_258),
.B1(n_234),
.B2(n_213),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_211),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_249),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_260),
.B(n_269),
.Y(n_279)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_265),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_266),
.B(n_268),
.C(n_278),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_244),
.B(n_253),
.C(n_248),
.Y(n_268)
);

INVxp67_ASAP7_75t_L g269 ( 
.A(n_243),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_245),
.B(n_233),
.Y(n_270)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_270),
.Y(n_287)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_245),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_271),
.B(n_274),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_241),
.B(n_212),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_254),
.B(n_232),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g292 ( 
.A(n_275),
.B(n_258),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_276),
.A2(n_277),
.B1(n_261),
.B2(n_262),
.Y(n_289)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_246),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_239),
.B(n_212),
.C(n_225),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_264),
.B(n_256),
.C(n_255),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_282),
.B(n_283),
.C(n_284),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_264),
.B(n_240),
.C(n_247),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_268),
.B(n_250),
.C(n_236),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_L g285 ( 
.A1(n_274),
.A2(n_257),
.B1(n_237),
.B2(n_258),
.Y(n_285)
);

INVxp67_ASAP7_75t_L g294 ( 
.A(n_285),
.Y(n_294)
);

INVx4_ASAP7_75t_L g286 ( 
.A(n_269),
.Y(n_286)
);

INVxp67_ASAP7_75t_L g299 ( 
.A(n_286),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_263),
.A2(n_258),
.B1(n_236),
.B2(n_219),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_288),
.A2(n_289),
.B1(n_281),
.B2(n_291),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_275),
.B(n_208),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_290),
.B(n_292),
.C(n_293),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_266),
.B(n_208),
.Y(n_293)
);

A2O1A1O1Ixp25_ASAP7_75t_L g295 ( 
.A1(n_292),
.A2(n_262),
.B(n_271),
.C(n_270),
.D(n_261),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_295),
.B(n_304),
.Y(n_312)
);

XOR2xp5_ASAP7_75t_L g314 ( 
.A(n_298),
.B(n_303),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_280),
.B(n_278),
.C(n_276),
.Y(n_300)
);

OAI21xp5_ASAP7_75t_L g310 ( 
.A1(n_300),
.A2(n_5),
.B(n_3),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_L g301 ( 
.A1(n_288),
.A2(n_272),
.B1(n_267),
.B2(n_209),
.Y(n_301)
);

INVxp67_ASAP7_75t_L g316 ( 
.A(n_301),
.Y(n_316)
);

OAI221xp5_ASAP7_75t_L g302 ( 
.A1(n_279),
.A2(n_238),
.B1(n_273),
.B2(n_215),
.C(n_13),
.Y(n_302)
);

NOR2xp67_ASAP7_75t_L g313 ( 
.A(n_302),
.B(n_4),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_280),
.B(n_15),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_283),
.A2(n_6),
.B1(n_14),
.B2(n_3),
.Y(n_304)
);

AO21x1_ASAP7_75t_SL g305 ( 
.A1(n_287),
.A2(n_284),
.B(n_286),
.Y(n_305)
);

NOR2x1_ASAP7_75t_R g315 ( 
.A(n_305),
.B(n_4),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_282),
.B(n_14),
.C(n_2),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_306),
.B(n_1),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_307),
.B(n_311),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_299),
.B(n_14),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_SL g321 ( 
.A(n_308),
.B(n_309),
.Y(n_321)
);

NOR2x1_ASAP7_75t_L g309 ( 
.A(n_305),
.B(n_2),
.Y(n_309)
);

XOR2xp5_ASAP7_75t_L g317 ( 
.A(n_310),
.B(n_296),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_299),
.B(n_4),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_313),
.B(n_294),
.Y(n_322)
);

AOI21xp5_ASAP7_75t_SL g319 ( 
.A1(n_315),
.A2(n_5),
.B(n_295),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_317),
.B(n_320),
.C(n_322),
.Y(n_325)
);

INVxp67_ASAP7_75t_L g324 ( 
.A(n_319),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_SL g320 ( 
.A(n_312),
.B(n_300),
.Y(n_320)
);

XOR2xp5_ASAP7_75t_L g323 ( 
.A(n_314),
.B(n_297),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_323),
.B(n_297),
.C(n_315),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_SL g328 ( 
.A(n_326),
.B(n_327),
.Y(n_328)
);

MAJx2_ASAP7_75t_L g327 ( 
.A(n_321),
.B(n_309),
.C(n_316),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_SL g329 ( 
.A(n_324),
.B(n_316),
.Y(n_329)
);

AOI21xp5_ASAP7_75t_L g330 ( 
.A1(n_329),
.A2(n_294),
.B(n_325),
.Y(n_330)
);

OA21x2_ASAP7_75t_L g331 ( 
.A1(n_330),
.A2(n_328),
.B(n_321),
.Y(n_331)
);

HAxp5_ASAP7_75t_SL g332 ( 
.A(n_331),
.B(n_318),
.CON(n_332),
.SN(n_332)
);

XNOR2xp5_ASAP7_75t_L g333 ( 
.A(n_332),
.B(n_5),
.Y(n_333)
);


endmodule