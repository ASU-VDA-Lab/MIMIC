module fake_jpeg_30012_n_325 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_325);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_325;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx13_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_16),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_5),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_11),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_6),
.Y(n_22)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_10),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_7),
.Y(n_26)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_11),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

BUFx2_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

INVx2_ASAP7_75t_SL g35 ( 
.A(n_15),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_1),
.Y(n_36)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_12),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_0),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_1),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_15),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_13),
.Y(n_41)
);

CKINVDCx16_ASAP7_75t_R g42 ( 
.A(n_24),
.Y(n_42)
);

INVx4_ASAP7_75t_SL g101 ( 
.A(n_42),
.Y(n_101)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_28),
.Y(n_43)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_43),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_28),
.B(n_0),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_44),
.B(n_49),
.Y(n_89)
);

INVx1_ASAP7_75t_SL g45 ( 
.A(n_24),
.Y(n_45)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_45),
.B(n_46),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_19),
.B(n_8),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_30),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_47),
.Y(n_83)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_17),
.Y(n_48)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_48),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_28),
.B(n_0),
.Y(n_49)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_30),
.Y(n_50)
);

INVx5_ASAP7_75t_L g86 ( 
.A(n_50),
.Y(n_86)
);

INVx2_ASAP7_75t_SL g51 ( 
.A(n_36),
.Y(n_51)
);

INVx2_ASAP7_75t_SL g97 ( 
.A(n_51),
.Y(n_97)
);

INVx11_ASAP7_75t_L g52 ( 
.A(n_30),
.Y(n_52)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_52),
.Y(n_80)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_30),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_53),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_19),
.B(n_8),
.Y(n_54)
);

OR2x2_ASAP7_75t_L g82 ( 
.A(n_54),
.B(n_57),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_17),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_55),
.Y(n_96)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_18),
.Y(n_56)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_56),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_20),
.B(n_8),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_17),
.Y(n_58)
);

BUFx2_ASAP7_75t_L g98 ( 
.A(n_58),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_29),
.Y(n_59)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_59),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_33),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_60),
.B(n_61),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_20),
.B(n_9),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_29),
.Y(n_62)
);

BUFx12f_ASAP7_75t_L g70 ( 
.A(n_62),
.Y(n_70)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_29),
.Y(n_63)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_63),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_29),
.Y(n_64)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_64),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_46),
.A2(n_41),
.B1(n_25),
.B2(n_26),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_67),
.A2(n_75),
.B1(n_93),
.B2(n_103),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_L g68 ( 
.A1(n_63),
.A2(n_33),
.B1(n_32),
.B2(n_27),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_68),
.A2(n_71),
.B1(n_105),
.B2(n_77),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_L g71 ( 
.A1(n_63),
.A2(n_33),
.B1(n_32),
.B2(n_27),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_54),
.B(n_41),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_74),
.B(n_76),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_50),
.A2(n_35),
.B1(n_33),
.B2(n_23),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_57),
.B(n_22),
.Y(n_76)
);

NAND2x2_ASAP7_75t_L g77 ( 
.A(n_60),
.B(n_35),
.Y(n_77)
);

OA22x2_ASAP7_75t_L g124 ( 
.A1(n_77),
.A2(n_53),
.B1(n_51),
.B2(n_47),
.Y(n_124)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_43),
.Y(n_79)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_79),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_42),
.B(n_22),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_81),
.B(n_84),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_56),
.B(n_31),
.Y(n_84)
);

A2O1A1Ixp33_ASAP7_75t_L g85 ( 
.A1(n_44),
.A2(n_49),
.B(n_21),
.C(n_18),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_SL g117 ( 
.A1(n_85),
.A2(n_35),
.B(n_51),
.Y(n_117)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_45),
.Y(n_87)
);

CKINVDCx16_ASAP7_75t_R g122 ( 
.A(n_87),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_59),
.B(n_31),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_90),
.B(n_91),
.Y(n_133)
);

AOI21xp33_ASAP7_75t_L g91 ( 
.A1(n_48),
.A2(n_21),
.B(n_26),
.Y(n_91)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_55),
.Y(n_92)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_92),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_59),
.A2(n_32),
.B1(n_27),
.B2(n_37),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_62),
.B(n_25),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_94),
.B(n_100),
.Y(n_142)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_55),
.Y(n_95)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_95),
.Y(n_129)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_58),
.Y(n_99)
);

INVx1_ASAP7_75t_SL g121 ( 
.A(n_99),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_48),
.B(n_39),
.Y(n_100)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_58),
.Y(n_102)
);

CKINVDCx16_ASAP7_75t_R g145 ( 
.A(n_102),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_50),
.A2(n_35),
.B1(n_23),
.B2(n_37),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_L g105 ( 
.A1(n_62),
.A2(n_32),
.B1(n_37),
.B2(n_23),
.Y(n_105)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_64),
.Y(n_106)
);

INVx1_ASAP7_75t_SL g123 ( 
.A(n_106),
.Y(n_123)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_52),
.Y(n_108)
);

INVx1_ASAP7_75t_SL g138 ( 
.A(n_108),
.Y(n_138)
);

BUFx10_ASAP7_75t_L g109 ( 
.A(n_48),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_109),
.Y(n_135)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_78),
.Y(n_110)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_110),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_109),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_111),
.B(n_117),
.Y(n_147)
);

BUFx3_ASAP7_75t_L g112 ( 
.A(n_66),
.Y(n_112)
);

INVx4_ASAP7_75t_L g163 ( 
.A(n_112),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_89),
.B(n_107),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_114),
.B(n_115),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_107),
.B(n_39),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_65),
.Y(n_116)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_116),
.Y(n_156)
);

OAI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_77),
.A2(n_64),
.B1(n_47),
.B2(n_53),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_119),
.A2(n_80),
.B1(n_88),
.B2(n_86),
.Y(n_179)
);

AND2x2_ASAP7_75t_L g169 ( 
.A(n_120),
.B(n_124),
.Y(n_169)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_96),
.Y(n_125)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_125),
.Y(n_152)
);

INVx8_ASAP7_75t_L g127 ( 
.A(n_88),
.Y(n_127)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_127),
.Y(n_161)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_96),
.Y(n_130)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_130),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_109),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_131),
.B(n_139),
.Y(n_154)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_73),
.Y(n_132)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_132),
.Y(n_165)
);

BUFx2_ASAP7_75t_L g134 ( 
.A(n_73),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_134),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_83),
.Y(n_136)
);

HB1xp67_ASAP7_75t_L g177 ( 
.A(n_136),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_83),
.Y(n_137)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_137),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_98),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_98),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_140),
.B(n_97),
.Y(n_158)
);

AOI21xp5_ASAP7_75t_L g141 ( 
.A1(n_77),
.A2(n_36),
.B(n_40),
.Y(n_141)
);

AOI21xp5_ASAP7_75t_SL g178 ( 
.A1(n_141),
.A2(n_86),
.B(n_70),
.Y(n_178)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_72),
.Y(n_144)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_144),
.Y(n_172)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_70),
.Y(n_146)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_146),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_143),
.B(n_69),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g186 ( 
.A(n_148),
.B(n_153),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_113),
.B(n_82),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_133),
.B(n_85),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_155),
.B(n_170),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_126),
.A2(n_105),
.B1(n_71),
.B2(n_68),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_157),
.A2(n_159),
.B1(n_124),
.B2(n_138),
.Y(n_198)
);

INVxp67_ASAP7_75t_L g197 ( 
.A(n_158),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_141),
.A2(n_103),
.B1(n_75),
.B2(n_82),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_L g160 ( 
.A1(n_120),
.A2(n_101),
.B1(n_80),
.B2(n_104),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_160),
.A2(n_121),
.B1(n_132),
.B2(n_134),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_142),
.B(n_101),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_162),
.B(n_164),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_122),
.B(n_34),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g166 ( 
.A(n_114),
.B(n_97),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_166),
.B(n_118),
.C(n_144),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_112),
.Y(n_167)
);

OR2x2_ASAP7_75t_L g189 ( 
.A(n_167),
.B(n_176),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_110),
.B(n_104),
.Y(n_170)
);

AND2x2_ASAP7_75t_L g171 ( 
.A(n_124),
.B(n_115),
.Y(n_171)
);

AND2x2_ASAP7_75t_L g183 ( 
.A(n_171),
.B(n_178),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_117),
.B(n_38),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_174),
.B(n_180),
.Y(n_191)
);

OR2x2_ASAP7_75t_L g176 ( 
.A(n_135),
.B(n_38),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_179),
.A2(n_140),
.B1(n_139),
.B2(n_123),
.Y(n_207)
);

OAI32xp33_ASAP7_75t_L g180 ( 
.A1(n_124),
.A2(n_34),
.A3(n_70),
.B1(n_40),
.B2(n_36),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_116),
.Y(n_181)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_181),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_138),
.B(n_34),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_182),
.B(n_135),
.Y(n_192)
);

INVx1_ASAP7_75t_SL g184 ( 
.A(n_163),
.Y(n_184)
);

INVxp67_ASAP7_75t_SL g233 ( 
.A(n_184),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_154),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_185),
.B(n_194),
.Y(n_226)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_149),
.Y(n_188)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_188),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_192),
.B(n_201),
.Y(n_223)
);

INVx4_ASAP7_75t_L g193 ( 
.A(n_163),
.Y(n_193)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_193),
.Y(n_217)
);

NOR2x1_ASAP7_75t_L g194 ( 
.A(n_171),
.B(n_155),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_176),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_195),
.B(n_204),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_159),
.A2(n_171),
.B1(n_169),
.B2(n_157),
.Y(n_196)
);

INVxp67_ASAP7_75t_L g224 ( 
.A(n_196),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_198),
.A2(n_215),
.B1(n_1),
.B2(n_2),
.Y(n_240)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_152),
.Y(n_199)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_199),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_200),
.B(n_203),
.Y(n_229)
);

AO22x1_ASAP7_75t_L g201 ( 
.A1(n_169),
.A2(n_147),
.B1(n_180),
.B2(n_178),
.Y(n_201)
);

INVx3_ASAP7_75t_L g202 ( 
.A(n_167),
.Y(n_202)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_202),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_166),
.B(n_151),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_151),
.B(n_145),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_170),
.B(n_118),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_205),
.B(n_208),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_207),
.A2(n_209),
.B1(n_212),
.B2(n_150),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_149),
.B(n_123),
.Y(n_208)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_152),
.Y(n_210)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_210),
.Y(n_228)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_156),
.Y(n_211)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_211),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_169),
.A2(n_121),
.B1(n_137),
.B2(n_136),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_182),
.B(n_129),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_213),
.B(n_214),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_175),
.B(n_34),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_179),
.A2(n_127),
.B1(n_129),
.B2(n_128),
.Y(n_215)
);

AOI21xp5_ASAP7_75t_L g216 ( 
.A1(n_183),
.A2(n_175),
.B(n_150),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_216),
.B(n_240),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_203),
.B(n_181),
.C(n_156),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_222),
.B(n_200),
.C(n_197),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_189),
.B(n_165),
.Y(n_227)
);

CKINVDCx14_ASAP7_75t_R g253 ( 
.A(n_227),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_198),
.A2(n_172),
.B1(n_177),
.B2(n_165),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_L g244 ( 
.A1(n_230),
.A2(n_231),
.B1(n_239),
.B2(n_215),
.Y(n_244)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_211),
.Y(n_232)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_232),
.Y(n_250)
);

AOI322xp5_ASAP7_75t_L g235 ( 
.A1(n_191),
.A2(n_34),
.A3(n_172),
.B1(n_161),
.B2(n_173),
.C1(n_125),
.C2(n_130),
.Y(n_235)
);

OAI321xp33_ASAP7_75t_L g245 ( 
.A1(n_235),
.A2(n_192),
.A3(n_190),
.B1(n_212),
.B2(n_213),
.C(n_208),
.Y(n_245)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_187),
.Y(n_237)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_237),
.Y(n_252)
);

OAI32xp33_ASAP7_75t_L g238 ( 
.A1(n_190),
.A2(n_161),
.A3(n_173),
.B1(n_168),
.B2(n_128),
.Y(n_238)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_238),
.Y(n_256)
);

AOI22x1_ASAP7_75t_SL g239 ( 
.A1(n_201),
.A2(n_168),
.B1(n_146),
.B2(n_40),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_SL g241 ( 
.A(n_201),
.B(n_9),
.C(n_14),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_241),
.B(n_189),
.Y(n_243)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_217),
.Y(n_242)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_242),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_243),
.B(n_249),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_244),
.A2(n_245),
.B1(n_239),
.B2(n_240),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_247),
.B(n_248),
.C(n_251),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_229),
.B(n_196),
.C(n_183),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_234),
.B(n_186),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_229),
.B(n_183),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_222),
.B(n_194),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_254),
.B(n_262),
.C(n_224),
.Y(n_268)
);

A2O1A1O1Ixp25_ASAP7_75t_L g255 ( 
.A1(n_223),
.A2(n_206),
.B(n_205),
.C(n_197),
.D(n_209),
.Y(n_255)
);

OAI21xp5_ASAP7_75t_L g275 ( 
.A1(n_255),
.A2(n_228),
.B(n_220),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_226),
.B(n_193),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_257),
.Y(n_274)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_219),
.Y(n_258)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_258),
.Y(n_263)
);

CKINVDCx16_ASAP7_75t_R g259 ( 
.A(n_221),
.Y(n_259)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_259),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_223),
.B(n_202),
.Y(n_260)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_260),
.Y(n_265)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_218),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_261),
.B(n_225),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_224),
.B(n_184),
.C(n_210),
.Y(n_262)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_267),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_268),
.B(n_5),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_246),
.B(n_225),
.Y(n_269)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_269),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_271),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_256),
.A2(n_231),
.B1(n_241),
.B2(n_236),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_272),
.A2(n_273),
.B1(n_277),
.B2(n_255),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_256),
.A2(n_216),
.B1(n_238),
.B2(n_221),
.Y(n_273)
);

AOI21x1_ASAP7_75t_L g282 ( 
.A1(n_275),
.A2(n_262),
.B(n_251),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_246),
.A2(n_217),
.B1(n_228),
.B2(n_220),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_248),
.B(n_199),
.C(n_233),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_278),
.B(n_250),
.C(n_9),
.Y(n_285)
);

AOI22xp33_ASAP7_75t_L g280 ( 
.A1(n_275),
.A2(n_253),
.B1(n_261),
.B2(n_252),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_280),
.B(n_281),
.Y(n_292)
);

OAI21xp5_ASAP7_75t_L g296 ( 
.A1(n_282),
.A2(n_268),
.B(n_278),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_266),
.B(n_254),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_283),
.B(n_289),
.Y(n_300)
);

AOI321xp33_ASAP7_75t_L g284 ( 
.A1(n_276),
.A2(n_247),
.A3(n_250),
.B1(n_258),
.B2(n_252),
.C(n_242),
.Y(n_284)
);

OAI211xp5_ASAP7_75t_L g297 ( 
.A1(n_284),
.A2(n_288),
.B(n_267),
.C(n_263),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_285),
.B(n_286),
.C(n_274),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_266),
.B(n_6),
.C(n_14),
.Y(n_286)
);

INVxp67_ASAP7_75t_L g287 ( 
.A(n_277),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_287),
.B(n_270),
.Y(n_302)
);

AOI21xp5_ASAP7_75t_L g288 ( 
.A1(n_274),
.A2(n_11),
.B(n_14),
.Y(n_288)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_293),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_291),
.A2(n_272),
.B1(n_265),
.B2(n_263),
.Y(n_294)
);

INVxp67_ASAP7_75t_L g307 ( 
.A(n_294),
.Y(n_307)
);

OAI21xp33_ASAP7_75t_L g295 ( 
.A1(n_290),
.A2(n_269),
.B(n_265),
.Y(n_295)
);

AOI21xp5_ASAP7_75t_L g310 ( 
.A1(n_295),
.A2(n_296),
.B(n_302),
.Y(n_310)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_297),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_287),
.A2(n_264),
.B1(n_271),
.B2(n_273),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_298),
.A2(n_5),
.B1(n_13),
.B2(n_3),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_281),
.B(n_264),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_SL g309 ( 
.A(n_299),
.B(n_3),
.Y(n_309)
);

O2A1O1Ixp33_ASAP7_75t_L g301 ( 
.A1(n_279),
.A2(n_270),
.B(n_285),
.C(n_283),
.Y(n_301)
);

OAI21xp5_ASAP7_75t_L g305 ( 
.A1(n_301),
.A2(n_286),
.B(n_289),
.Y(n_305)
);

XOR2xp5_ASAP7_75t_L g314 ( 
.A(n_305),
.B(n_300),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_296),
.B(n_300),
.C(n_292),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_SL g315 ( 
.A(n_306),
.B(n_308),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_309),
.B(n_13),
.Y(n_312)
);

NOR2xp67_ASAP7_75t_SL g311 ( 
.A(n_306),
.B(n_301),
.Y(n_311)
);

AOI21xp5_ASAP7_75t_L g318 ( 
.A1(n_311),
.A2(n_313),
.B(n_307),
.Y(n_318)
);

OR2x2_ASAP7_75t_L g320 ( 
.A(n_312),
.B(n_316),
.Y(n_320)
);

OAI21xp5_ASAP7_75t_SL g313 ( 
.A1(n_304),
.A2(n_293),
.B(n_295),
.Y(n_313)
);

XOR2xp5_ASAP7_75t_L g319 ( 
.A(n_314),
.B(n_12),
.Y(n_319)
);

OAI321xp33_ASAP7_75t_L g316 ( 
.A1(n_310),
.A2(n_3),
.A3(n_4),
.B1(n_12),
.B2(n_16),
.C(n_1),
.Y(n_316)
);

OAI21xp5_ASAP7_75t_SL g317 ( 
.A1(n_315),
.A2(n_303),
.B(n_307),
.Y(n_317)
);

INVxp67_ASAP7_75t_L g322 ( 
.A(n_317),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_318),
.B(n_319),
.Y(n_321)
);

XOR2xp5_ASAP7_75t_L g323 ( 
.A(n_321),
.B(n_320),
.Y(n_323)
);

OAI21x1_ASAP7_75t_L g324 ( 
.A1(n_323),
.A2(n_322),
.B(n_320),
.Y(n_324)
);

AOI21xp5_ASAP7_75t_L g325 ( 
.A1(n_324),
.A2(n_4),
.B(n_2),
.Y(n_325)
);


endmodule