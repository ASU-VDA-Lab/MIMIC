module fake_jpeg_13030_n_137 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_137);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_137;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_11),
.B(n_3),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_16),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_1),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_24),
.Y(n_44)
);

INVx11_ASAP7_75t_L g45 ( 
.A(n_19),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_29),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_7),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_31),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_13),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_40),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_35),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_14),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_1),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_3),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_8),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_10),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_2),
.Y(n_57)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_45),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_58),
.B(n_59),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_45),
.Y(n_59)
);

BUFx4f_ASAP7_75t_SL g60 ( 
.A(n_42),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_60),
.B(n_64),
.Y(n_77)
);

BUFx4f_ASAP7_75t_L g61 ( 
.A(n_47),
.Y(n_61)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_61),
.Y(n_81)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_43),
.Y(n_62)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_62),
.Y(n_73)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_47),
.Y(n_63)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_63),
.Y(n_76)
);

OR2x4_ASAP7_75t_L g64 ( 
.A(n_41),
.B(n_0),
.Y(n_64)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_44),
.Y(n_65)
);

NAND2xp33_ASAP7_75t_SL g78 ( 
.A(n_65),
.B(n_66),
.Y(n_78)
);

INVx8_ASAP7_75t_L g66 ( 
.A(n_44),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_55),
.B(n_57),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_67),
.B(n_68),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_46),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_68),
.A2(n_46),
.B1(n_48),
.B2(n_54),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_70),
.B(n_79),
.Y(n_89)
);

OA22x2_ASAP7_75t_L g71 ( 
.A1(n_66),
.A2(n_48),
.B1(n_51),
.B2(n_50),
.Y(n_71)
);

OA22x2_ASAP7_75t_SL g94 ( 
.A1(n_71),
.A2(n_75),
.B1(n_5),
.B2(n_6),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_67),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_74),
.B(n_5),
.Y(n_91)
);

OAI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_61),
.A2(n_57),
.B1(n_56),
.B2(n_54),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_58),
.B(n_52),
.Y(n_79)
);

OAI32xp33_ASAP7_75t_L g80 ( 
.A1(n_58),
.A2(n_53),
.A3(n_49),
.B1(n_43),
.B2(n_56),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_80),
.B(n_60),
.Y(n_86)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_81),
.Y(n_82)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_82),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_77),
.B(n_49),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_83),
.B(n_85),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_78),
.A2(n_53),
.B1(n_2),
.B2(n_4),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_84),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_72),
.B(n_0),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_86),
.A2(n_94),
.B1(n_96),
.B2(n_71),
.Y(n_97)
);

INVx1_ASAP7_75t_SL g87 ( 
.A(n_76),
.Y(n_87)
);

CKINVDCx5p33_ASAP7_75t_R g99 ( 
.A(n_87),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_69),
.Y(n_88)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_88),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_73),
.B(n_4),
.Y(n_90)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_90),
.Y(n_106)
);

OR2x2_ASAP7_75t_L g103 ( 
.A(n_91),
.B(n_92),
.Y(n_103)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_79),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_81),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_93),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_72),
.B(n_71),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_95),
.B(n_9),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_L g96 ( 
.A1(n_71),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_97),
.A2(n_107),
.B1(n_109),
.B2(n_20),
.Y(n_122)
);

HAxp5_ASAP7_75t_SL g101 ( 
.A(n_94),
.B(n_80),
.CON(n_101),
.SN(n_101)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_101),
.B(n_111),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_SL g104 ( 
.A1(n_88),
.A2(n_78),
.B(n_10),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_104),
.B(n_110),
.C(n_12),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_89),
.A2(n_9),
.B1(n_11),
.B2(n_12),
.Y(n_107)
);

OAI32xp33_ASAP7_75t_L g109 ( 
.A1(n_89),
.A2(n_26),
.A3(n_38),
.B1(n_37),
.B2(n_15),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_87),
.B(n_25),
.C(n_36),
.Y(n_110)
);

AOI21xp5_ASAP7_75t_SL g124 ( 
.A1(n_112),
.A2(n_114),
.B(n_115),
.Y(n_124)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_98),
.Y(n_113)
);

HB1xp67_ASAP7_75t_L g127 ( 
.A(n_113),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_108),
.B(n_102),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_100),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_111),
.B(n_82),
.C(n_94),
.Y(n_116)
);

A2O1A1O1Ixp25_ASAP7_75t_L g126 ( 
.A1(n_116),
.A2(n_117),
.B(n_119),
.C(n_120),
.D(n_121),
.Y(n_126)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_99),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_101),
.A2(n_13),
.B1(n_17),
.B2(n_18),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_118),
.A2(n_122),
.B1(n_103),
.B2(n_106),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_104),
.B(n_105),
.C(n_103),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_99),
.Y(n_120)
);

NAND3xp33_ASAP7_75t_L g130 ( 
.A(n_123),
.B(n_39),
.C(n_23),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_116),
.A2(n_105),
.B1(n_109),
.B2(n_110),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_L g128 ( 
.A1(n_125),
.A2(n_126),
.B(n_119),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_128),
.B(n_129),
.C(n_127),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_124),
.B(n_112),
.C(n_22),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_130),
.B(n_21),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_131),
.B(n_132),
.C(n_27),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_133),
.B(n_28),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_L g135 ( 
.A1(n_134),
.A2(n_30),
.B(n_32),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_135),
.B(n_33),
.C(n_34),
.Y(n_136)
);

XOR2xp5_ASAP7_75t_L g137 ( 
.A(n_136),
.B(n_127),
.Y(n_137)
);


endmodule