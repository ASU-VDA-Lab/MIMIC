module fake_jpeg_15021_n_239 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_239);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_239;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_182;
wire n_19;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_122;
wire n_75;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx3_ASAP7_75t_L g16 ( 
.A(n_14),
.Y(n_16)
);

INVx8_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

INVx8_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

CKINVDCx16_ASAP7_75t_R g19 ( 
.A(n_6),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

INVx5_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_2),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

INVx8_ASAP7_75t_SL g33 ( 
.A(n_1),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_30),
.B(n_9),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_34),
.B(n_35),
.Y(n_43)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_20),
.Y(n_35)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_20),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_36),
.Y(n_56)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_33),
.Y(n_37)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_20),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_38),
.B(n_31),
.Y(n_52)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_20),
.Y(n_39)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_39),
.Y(n_44)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_22),
.Y(n_40)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_40),
.Y(n_45)
);

INVx4_ASAP7_75t_SL g41 ( 
.A(n_33),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_41),
.B(n_16),
.Y(n_46)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_22),
.Y(n_42)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_42),
.Y(n_51)
);

INVxp67_ASAP7_75t_L g73 ( 
.A(n_46),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g47 ( 
.A1(n_40),
.A2(n_24),
.B1(n_18),
.B2(n_17),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_47),
.A2(n_49),
.B1(n_53),
.B2(n_58),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_39),
.B(n_26),
.Y(n_48)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_48),
.B(n_0),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_L g49 ( 
.A1(n_40),
.A2(n_24),
.B1(n_18),
.B2(n_17),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_34),
.B(n_27),
.Y(n_50)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_50),
.Y(n_66)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_52),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_41),
.A2(n_24),
.B1(n_18),
.B2(n_17),
.Y(n_53)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

INVx5_ASAP7_75t_L g81 ( 
.A(n_55),
.Y(n_81)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_37),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_57),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g58 ( 
.A1(n_42),
.A2(n_25),
.B1(n_26),
.B2(n_27),
.Y(n_58)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_36),
.Y(n_59)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_59),
.Y(n_62)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_36),
.Y(n_60)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_60),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_54),
.A2(n_41),
.B1(n_19),
.B2(n_35),
.Y(n_63)
);

AOI21xp5_ASAP7_75t_L g103 ( 
.A1(n_63),
.A2(n_83),
.B(n_4),
.Y(n_103)
);

A2O1A1Ixp33_ASAP7_75t_L g64 ( 
.A1(n_43),
.A2(n_30),
.B(n_21),
.C(n_25),
.Y(n_64)
);

AO21x1_ASAP7_75t_L g104 ( 
.A1(n_64),
.A2(n_85),
.B(n_91),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_48),
.A2(n_42),
.B1(n_35),
.B2(n_37),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_67),
.A2(n_76),
.B1(n_95),
.B2(n_3),
.Y(n_99)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_51),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_68),
.B(n_71),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_43),
.B(n_50),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_69),
.B(n_70),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_58),
.B(n_29),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_46),
.B(n_29),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_44),
.B(n_21),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_72),
.B(n_93),
.Y(n_120)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_74),
.B(n_0),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_45),
.A2(n_37),
.B1(n_38),
.B2(n_19),
.Y(n_76)
);

OAI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_59),
.A2(n_28),
.B1(n_32),
.B2(n_22),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_L g97 ( 
.A1(n_77),
.A2(n_86),
.B1(n_23),
.B2(n_16),
.Y(n_97)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_44),
.Y(n_78)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_78),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_54),
.B(n_31),
.Y(n_80)
);

CKINVDCx16_ASAP7_75t_R g105 ( 
.A(n_80),
.Y(n_105)
);

INVx2_ASAP7_75t_SL g82 ( 
.A(n_57),
.Y(n_82)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_82),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_59),
.A2(n_41),
.B1(n_32),
.B2(n_28),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_47),
.B(n_0),
.Y(n_84)
);

XOR2xp5_ASAP7_75t_L g100 ( 
.A(n_84),
.B(n_90),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_56),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_45),
.A2(n_32),
.B1(n_28),
.B2(n_23),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_60),
.B(n_16),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_87),
.Y(n_106)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_56),
.Y(n_88)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_88),
.Y(n_116)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_57),
.Y(n_89)
);

BUFx5_ASAP7_75t_L g108 ( 
.A(n_89),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_57),
.B(n_38),
.C(n_31),
.Y(n_90)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_51),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_56),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_92),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_55),
.B(n_0),
.Y(n_93)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_60),
.Y(n_94)
);

HB1xp67_ASAP7_75t_L g121 ( 
.A(n_94),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_55),
.A2(n_23),
.B1(n_1),
.B2(n_3),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_L g127 ( 
.A1(n_96),
.A2(n_102),
.B(n_110),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_L g139 ( 
.A1(n_97),
.A2(n_99),
.B1(n_103),
.B2(n_81),
.Y(n_139)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_82),
.Y(n_101)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_101),
.Y(n_123)
);

AND2x2_ASAP7_75t_L g102 ( 
.A(n_93),
.B(n_3),
.Y(n_102)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_88),
.Y(n_107)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_107),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_65),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_109),
.A2(n_112),
.B1(n_118),
.B2(n_119),
.Y(n_131)
);

AOI21xp5_ASAP7_75t_L g110 ( 
.A1(n_84),
.A2(n_6),
.B(n_8),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_70),
.A2(n_67),
.B1(n_73),
.B2(n_69),
.Y(n_112)
);

AOI32xp33_ASAP7_75t_L g115 ( 
.A1(n_73),
.A2(n_8),
.A3(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_115),
.B(n_13),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_95),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_84),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_119)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_82),
.Y(n_122)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_122),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_117),
.B(n_66),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_124),
.B(n_128),
.Y(n_159)
);

A2O1A1Ixp33_ASAP7_75t_SL g126 ( 
.A1(n_103),
.A2(n_76),
.B(n_72),
.C(n_91),
.Y(n_126)
);

AOI21xp5_ASAP7_75t_SL g157 ( 
.A1(n_126),
.A2(n_116),
.B(n_114),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_117),
.B(n_74),
.Y(n_128)
);

AOI21xp5_ASAP7_75t_L g129 ( 
.A1(n_100),
.A2(n_94),
.B(n_81),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_SL g161 ( 
.A1(n_129),
.A2(n_130),
.B(n_138),
.Y(n_161)
);

AO21x1_ASAP7_75t_L g130 ( 
.A1(n_104),
.A2(n_61),
.B(n_78),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g150 ( 
.A(n_132),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_113),
.B(n_61),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_133),
.B(n_134),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_112),
.B(n_74),
.Y(n_134)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_98),
.Y(n_136)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_136),
.Y(n_148)
);

AND2x6_ASAP7_75t_L g137 ( 
.A(n_104),
.B(n_64),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_137),
.B(n_147),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_120),
.A2(n_100),
.B1(n_99),
.B2(n_109),
.Y(n_138)
);

INVxp67_ASAP7_75t_L g160 ( 
.A(n_139),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_98),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_140),
.B(n_143),
.Y(n_165)
);

O2A1O1Ixp33_ASAP7_75t_L g141 ( 
.A1(n_113),
.A2(n_89),
.B(n_90),
.C(n_62),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_L g167 ( 
.A1(n_141),
.A2(n_145),
.B(n_105),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_120),
.A2(n_62),
.B1(n_75),
.B2(n_79),
.Y(n_142)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_142),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_111),
.B(n_75),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_SL g144 ( 
.A(n_110),
.B(n_14),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_144),
.B(n_118),
.Y(n_155)
);

AOI21xp5_ASAP7_75t_L g145 ( 
.A1(n_106),
.A2(n_79),
.B(n_14),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_107),
.Y(n_146)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_146),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_102),
.B(n_106),
.Y(n_147)
);

CKINVDCx16_ASAP7_75t_R g151 ( 
.A(n_123),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_151),
.B(n_135),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_125),
.B(n_121),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_153),
.B(n_164),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g154 ( 
.A(n_129),
.B(n_119),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_154),
.B(n_131),
.C(n_144),
.Y(n_178)
);

AOI21xp33_ASAP7_75t_L g179 ( 
.A1(n_155),
.A2(n_126),
.B(n_146),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_138),
.B(n_102),
.Y(n_156)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_156),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_SL g170 ( 
.A1(n_157),
.A2(n_169),
.B(n_145),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_130),
.B(n_96),
.Y(n_162)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_162),
.Y(n_185)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_136),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_130),
.B(n_96),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_166),
.B(n_127),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_L g180 ( 
.A1(n_167),
.A2(n_126),
.B1(n_125),
.B2(n_122),
.Y(n_180)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_123),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_168),
.B(n_108),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_L g169 ( 
.A1(n_127),
.A2(n_114),
.B(n_116),
.Y(n_169)
);

AOI21xp5_ASAP7_75t_L g198 ( 
.A1(n_170),
.A2(n_171),
.B(n_182),
.Y(n_198)
);

AOI21xp5_ASAP7_75t_L g171 ( 
.A1(n_161),
.A2(n_126),
.B(n_140),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_163),
.B(n_142),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_SL g197 ( 
.A(n_174),
.B(n_175),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_152),
.A2(n_126),
.B1(n_137),
.B2(n_141),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_176),
.A2(n_157),
.B1(n_166),
.B2(n_155),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_154),
.B(n_131),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_177),
.B(n_178),
.C(n_183),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_179),
.A2(n_180),
.B1(n_165),
.B2(n_148),
.Y(n_192)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_181),
.Y(n_190)
);

AOI21xp5_ASAP7_75t_L g182 ( 
.A1(n_161),
.A2(n_135),
.B(n_108),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g183 ( 
.A(n_156),
.B(n_101),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_184),
.B(n_158),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_160),
.A2(n_152),
.B1(n_157),
.B2(n_149),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_186),
.A2(n_167),
.B1(n_169),
.B2(n_162),
.Y(n_188)
);

CKINVDCx14_ASAP7_75t_R g211 ( 
.A(n_188),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_183),
.B(n_163),
.C(n_159),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_189),
.B(n_173),
.C(n_185),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_SL g207 ( 
.A1(n_191),
.A2(n_195),
.B(n_199),
.Y(n_207)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_192),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_172),
.B(n_165),
.Y(n_193)
);

CKINVDCx16_ASAP7_75t_R g209 ( 
.A(n_193),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_172),
.B(n_158),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_194),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_184),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_196),
.B(n_200),
.Y(n_203)
);

AOI21x1_ASAP7_75t_SL g199 ( 
.A1(n_171),
.A2(n_148),
.B(n_164),
.Y(n_199)
);

CKINVDCx16_ASAP7_75t_R g200 ( 
.A(n_182),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_187),
.B(n_177),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_201),
.B(n_202),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_187),
.B(n_178),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_188),
.B(n_189),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_205),
.B(n_210),
.C(n_212),
.Y(n_218)
);

NAND3xp33_ASAP7_75t_L g208 ( 
.A(n_199),
.B(n_175),
.C(n_150),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_208),
.B(n_176),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_191),
.B(n_186),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_211),
.A2(n_198),
.B1(n_173),
.B2(n_185),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_213),
.A2(n_214),
.B1(n_220),
.B2(n_210),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_SL g215 ( 
.A1(n_207),
.A2(n_198),
.B(n_170),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_215),
.B(n_207),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_206),
.B(n_195),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_216),
.B(n_217),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_209),
.B(n_197),
.Y(n_217)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_203),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_L g225 ( 
.A1(n_219),
.A2(n_190),
.B(n_197),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_204),
.A2(n_174),
.B1(n_196),
.B2(n_190),
.Y(n_220)
);

AOI21xp5_ASAP7_75t_L g229 ( 
.A1(n_222),
.A2(n_223),
.B(n_225),
.Y(n_229)
);

AOI21x1_ASAP7_75t_L g223 ( 
.A1(n_215),
.A2(n_203),
.B(n_212),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_226),
.B(n_227),
.Y(n_231)
);

NAND4xp25_ASAP7_75t_SL g227 ( 
.A(n_220),
.B(n_151),
.C(n_168),
.D(n_15),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_SL g228 ( 
.A1(n_224),
.A2(n_218),
.B(n_205),
.Y(n_228)
);

AO21x1_ASAP7_75t_L g234 ( 
.A1(n_228),
.A2(n_221),
.B(n_201),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_222),
.B(n_218),
.C(n_221),
.Y(n_230)
);

INVxp67_ASAP7_75t_SL g233 ( 
.A(n_230),
.Y(n_233)
);

OAI21x1_ASAP7_75t_L g232 ( 
.A1(n_229),
.A2(n_227),
.B(n_213),
.Y(n_232)
);

AOI21xp5_ASAP7_75t_L g235 ( 
.A1(n_232),
.A2(n_234),
.B(n_231),
.Y(n_235)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_235),
.Y(n_237)
);

A2O1A1Ixp33_ASAP7_75t_SL g236 ( 
.A1(n_233),
.A2(n_159),
.B(n_202),
.C(n_15),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_237),
.B(n_236),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_238),
.B(n_15),
.Y(n_239)
);


endmodule