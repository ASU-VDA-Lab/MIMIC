module fake_netlist_5_2539_n_109 (n_16, n_0, n_12, n_9, n_18, n_1, n_8, n_10, n_4, n_11, n_17, n_19, n_7, n_15, n_5, n_14, n_2, n_13, n_3, n_6, n_109);

input n_16;
input n_0;
input n_12;
input n_9;
input n_18;
input n_1;
input n_8;
input n_10;
input n_4;
input n_11;
input n_17;
input n_19;
input n_7;
input n_15;
input n_5;
input n_14;
input n_2;
input n_13;
input n_3;
input n_6;

output n_109;

wire n_91;
wire n_82;
wire n_24;
wire n_86;
wire n_83;
wire n_61;
wire n_90;
wire n_75;
wire n_101;
wire n_65;
wire n_78;
wire n_74;
wire n_57;
wire n_96;
wire n_37;
wire n_108;
wire n_31;
wire n_66;
wire n_98;
wire n_60;
wire n_43;
wire n_107;
wire n_58;
wire n_69;
wire n_42;
wire n_22;
wire n_45;
wire n_46;
wire n_21;
wire n_94;
wire n_38;
wire n_105;
wire n_80;
wire n_35;
wire n_73;
wire n_92;
wire n_30;
wire n_33;
wire n_84;
wire n_23;
wire n_29;
wire n_79;
wire n_47;
wire n_25;
wire n_53;
wire n_44;
wire n_40;
wire n_34;
wire n_100;
wire n_62;
wire n_71;
wire n_85;
wire n_95;
wire n_59;
wire n_26;
wire n_55;
wire n_99;
wire n_49;
wire n_20;
wire n_39;
wire n_54;
wire n_67;
wire n_36;
wire n_76;
wire n_87;
wire n_27;
wire n_77;
wire n_64;
wire n_102;
wire n_106;
wire n_81;
wire n_28;
wire n_89;
wire n_70;
wire n_68;
wire n_93;
wire n_72;
wire n_32;
wire n_41;
wire n_104;
wire n_103;
wire n_56;
wire n_51;
wire n_63;
wire n_97;
wire n_48;
wire n_50;
wire n_52;
wire n_88;

INVx1_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

INVx1_ASAP7_75t_SL g21 ( 
.A(n_12),
.Y(n_21)
);

INVx1_ASAP7_75t_SL g22 ( 
.A(n_0),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_1),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_3),
.Y(n_24)
);

INVxp67_ASAP7_75t_L g25 ( 
.A(n_18),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_17),
.Y(n_30)
);

HB1xp67_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

INVxp67_ASAP7_75t_SL g32 ( 
.A(n_2),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_11),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_3),
.Y(n_35)
);

BUFx2_ASAP7_75t_L g36 ( 
.A(n_23),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

CKINVDCx8_ASAP7_75t_R g38 ( 
.A(n_23),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_28),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_29),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_20),
.Y(n_43)
);

NAND2xp33_ASAP7_75t_SL g44 ( 
.A(n_24),
.B(n_1),
.Y(n_44)
);

CKINVDCx5p33_ASAP7_75t_R g45 ( 
.A(n_31),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_26),
.Y(n_46)
);

AND2x4_ASAP7_75t_L g47 ( 
.A(n_30),
.B(n_2),
.Y(n_47)
);

NAND2xp33_ASAP7_75t_SL g48 ( 
.A(n_24),
.B(n_4),
.Y(n_48)
);

AND2x2_ASAP7_75t_L g49 ( 
.A(n_45),
.B(n_21),
.Y(n_49)
);

INVxp33_ASAP7_75t_SL g50 ( 
.A(n_36),
.Y(n_50)
);

AO22x2_ASAP7_75t_L g51 ( 
.A1(n_47),
.A2(n_35),
.B1(n_32),
.B2(n_22),
.Y(n_51)
);

AO22x2_ASAP7_75t_L g52 ( 
.A1(n_47),
.A2(n_34),
.B1(n_33),
.B2(n_27),
.Y(n_52)
);

AO22x2_ASAP7_75t_L g53 ( 
.A1(n_37),
.A2(n_25),
.B1(n_5),
.B2(n_6),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

INVx1_ASAP7_75t_SL g58 ( 
.A(n_49),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g59 ( 
.A(n_51),
.B(n_39),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_54),
.B(n_41),
.Y(n_60)
);

BUFx4f_ASAP7_75t_L g61 ( 
.A(n_56),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_55),
.Y(n_62)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_57),
.Y(n_63)
);

A2O1A1Ixp33_ASAP7_75t_L g64 ( 
.A1(n_59),
.A2(n_44),
.B(n_48),
.C(n_42),
.Y(n_64)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_58),
.B(n_51),
.Y(n_65)
);

INVxp67_ASAP7_75t_L g66 ( 
.A(n_59),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_60),
.A2(n_51),
.B1(n_53),
.B2(n_52),
.Y(n_67)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_63),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_62),
.B(n_38),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_68),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_66),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_69),
.Y(n_72)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_65),
.B(n_52),
.Y(n_73)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_67),
.Y(n_74)
);

OA21x2_ASAP7_75t_L g75 ( 
.A1(n_74),
.A2(n_62),
.B(n_63),
.Y(n_75)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_70),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_71),
.Y(n_77)
);

BUFx2_ASAP7_75t_L g78 ( 
.A(n_72),
.Y(n_78)
);

INVx5_ASAP7_75t_SL g79 ( 
.A(n_76),
.Y(n_79)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_76),
.Y(n_80)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_77),
.Y(n_81)
);

AOI21xp5_ASAP7_75t_L g82 ( 
.A1(n_75),
.A2(n_61),
.B(n_74),
.Y(n_82)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_80),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_81),
.B(n_78),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_79),
.B(n_73),
.Y(n_85)
);

NOR2x1_ASAP7_75t_L g86 ( 
.A(n_82),
.B(n_78),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_79),
.B(n_64),
.Y(n_87)
);

BUFx2_ASAP7_75t_L g88 ( 
.A(n_81),
.Y(n_88)
);

HB1xp67_ASAP7_75t_L g89 ( 
.A(n_88),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_85),
.B(n_50),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_84),
.B(n_73),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_83),
.B(n_53),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_89),
.B(n_90),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_91),
.B(n_86),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_92),
.A2(n_87),
.B1(n_48),
.B2(n_44),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_89),
.B(n_87),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_89),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_94),
.B(n_39),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_93),
.B(n_50),
.Y(n_99)
);

NOR3xp33_ASAP7_75t_SL g100 ( 
.A(n_94),
.B(n_67),
.C(n_46),
.Y(n_100)
);

NOR3xp33_ASAP7_75t_L g101 ( 
.A(n_95),
.B(n_43),
.C(n_53),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_98),
.B(n_97),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_99),
.B(n_96),
.Y(n_103)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_100),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_104),
.A2(n_101),
.B1(n_52),
.B2(n_75),
.Y(n_105)
);

NAND4xp25_ASAP7_75t_L g106 ( 
.A(n_105),
.B(n_103),
.C(n_102),
.D(n_4),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_106),
.B(n_6),
.Y(n_107)
);

HB1xp67_ASAP7_75t_L g108 ( 
.A(n_107),
.Y(n_108)
);

AOI221xp5_ASAP7_75t_L g109 ( 
.A1(n_108),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.C(n_19),
.Y(n_109)
);


endmodule