module fake_jpeg_24193_n_331 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_331);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_331;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx3_ASAP7_75t_L g16 ( 
.A(n_14),
.Y(n_16)
);

HB1xp67_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_9),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_15),
.Y(n_20)
);

INVx6_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

INVx6_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

BUFx16f_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

INVxp67_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_0),
.Y(n_30)
);

INVx8_ASAP7_75t_SL g31 ( 
.A(n_2),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_12),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

INVx6_ASAP7_75t_SL g35 ( 
.A(n_4),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_31),
.Y(n_36)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_30),
.Y(n_37)
);

AND2x2_ASAP7_75t_L g50 ( 
.A(n_37),
.B(n_43),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_22),
.Y(n_38)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_27),
.B(n_15),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_39),
.A2(n_28),
.B1(n_19),
.B2(n_33),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_22),
.Y(n_40)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_22),
.Y(n_41)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_41),
.Y(n_62)
);

BUFx12_ASAP7_75t_L g42 ( 
.A(n_27),
.Y(n_42)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_42),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_18),
.B(n_0),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_22),
.Y(n_44)
);

BUFx2_ASAP7_75t_L g70 ( 
.A(n_44),
.Y(n_70)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_16),
.Y(n_45)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_45),
.Y(n_59)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_16),
.Y(n_46)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_46),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_18),
.B(n_0),
.Y(n_47)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_47),
.B(n_0),
.Y(n_61)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_44),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_48),
.B(n_49),
.Y(n_85)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_42),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_46),
.A2(n_21),
.B1(n_23),
.B2(n_20),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_52),
.A2(n_56),
.B1(n_55),
.B2(n_62),
.Y(n_97)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_54),
.B(n_57),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_46),
.A2(n_21),
.B1(n_23),
.B2(n_20),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_42),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_44),
.Y(n_60)
);

INVx5_ASAP7_75t_L g94 ( 
.A(n_60),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_61),
.B(n_9),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_43),
.A2(n_17),
.B1(n_29),
.B2(n_33),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_63),
.A2(n_71),
.B1(n_73),
.B2(n_35),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_44),
.Y(n_64)
);

INVx8_ASAP7_75t_L g92 ( 
.A(n_64),
.Y(n_92)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_42),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_65),
.B(n_68),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_44),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_67),
.Y(n_80)
);

INVx4_ASAP7_75t_SL g68 ( 
.A(n_36),
.Y(n_68)
);

OR2x2_ASAP7_75t_SL g109 ( 
.A(n_69),
.B(n_24),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_47),
.A2(n_30),
.B1(n_29),
.B2(n_19),
.Y(n_71)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_44),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_72),
.B(n_36),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_43),
.A2(n_28),
.B1(n_32),
.B2(n_24),
.Y(n_73)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_60),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_74),
.B(n_75),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_69),
.A2(n_47),
.B1(n_45),
.B2(n_37),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_50),
.B(n_37),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_76),
.B(n_79),
.Y(n_117)
);

AND2x2_ASAP7_75t_L g122 ( 
.A(n_77),
.B(n_12),
.Y(n_122)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_70),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_78),
.B(n_81),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_50),
.B(n_39),
.Y(n_79)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_53),
.Y(n_81)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_53),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_82),
.B(n_88),
.Y(n_118)
);

FAx1_ASAP7_75t_SL g133 ( 
.A(n_83),
.B(n_11),
.CI(n_10),
.CON(n_133),
.SN(n_133)
);

AOI21xp5_ASAP7_75t_L g84 ( 
.A1(n_50),
.A2(n_45),
.B(n_32),
.Y(n_84)
);

AOI21xp5_ASAP7_75t_L g119 ( 
.A1(n_84),
.A2(n_91),
.B(n_10),
.Y(n_119)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_68),
.Y(n_86)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_86),
.Y(n_115)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_59),
.Y(n_88)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_70),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_89),
.B(n_96),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_55),
.A2(n_15),
.B1(n_9),
.B2(n_11),
.Y(n_91)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_93),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_71),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_95),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_64),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_97),
.A2(n_103),
.B1(n_109),
.B2(n_34),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_58),
.Y(n_98)
);

INVx8_ASAP7_75t_L g123 ( 
.A(n_98),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_58),
.Y(n_99)
);

CKINVDCx16_ASAP7_75t_R g139 ( 
.A(n_99),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_61),
.B(n_36),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_100),
.B(n_101),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_61),
.B(n_27),
.Y(n_101)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_62),
.Y(n_102)
);

BUFx2_ASAP7_75t_L g137 ( 
.A(n_102),
.Y(n_137)
);

AO22x2_ASAP7_75t_SL g103 ( 
.A1(n_66),
.A2(n_41),
.B1(n_38),
.B2(n_40),
.Y(n_103)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_67),
.Y(n_104)
);

CKINVDCx14_ASAP7_75t_R g124 ( 
.A(n_104),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_48),
.B(n_25),
.Y(n_105)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_105),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_72),
.B(n_25),
.Y(n_106)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_106),
.Y(n_134)
);

BUFx3_ASAP7_75t_L g107 ( 
.A(n_49),
.Y(n_107)
);

INVx4_ASAP7_75t_L g116 ( 
.A(n_107),
.Y(n_116)
);

NAND2x1p5_ASAP7_75t_L g108 ( 
.A(n_54),
.B(n_35),
.Y(n_108)
);

AOI21xp5_ASAP7_75t_SL g114 ( 
.A1(n_108),
.A2(n_41),
.B(n_40),
.Y(n_114)
);

CKINVDCx16_ASAP7_75t_R g110 ( 
.A(n_57),
.Y(n_110)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_110),
.Y(n_136)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_51),
.Y(n_111)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_111),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_51),
.Y(n_112)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_112),
.Y(n_140)
);

AO21x1_ASAP7_75t_L g159 ( 
.A1(n_114),
.A2(n_42),
.B(n_98),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_L g167 ( 
.A1(n_119),
.A2(n_92),
.B1(n_94),
.B2(n_4),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_120),
.A2(n_133),
.B1(n_74),
.B2(n_3),
.Y(n_168)
);

MAJx2_ASAP7_75t_L g121 ( 
.A(n_84),
.B(n_41),
.C(n_40),
.Y(n_121)
);

MAJx2_ASAP7_75t_L g151 ( 
.A(n_121),
.B(n_103),
.C(n_107),
.Y(n_151)
);

OAI21xp33_ASAP7_75t_SL g163 ( 
.A1(n_122),
.A2(n_1),
.B(n_2),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_75),
.B(n_38),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_125),
.B(n_131),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_109),
.A2(n_34),
.B1(n_26),
.B2(n_38),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g165 ( 
.A(n_130),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_77),
.B(n_26),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_87),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_141),
.Y(n_164)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_90),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_142),
.B(n_115),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_143),
.B(n_145),
.Y(n_180)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_118),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_129),
.B(n_77),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_146),
.B(n_147),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_129),
.B(n_83),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_125),
.B(n_108),
.Y(n_148)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_148),
.Y(n_179)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_118),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_149),
.B(n_152),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_120),
.A2(n_103),
.B1(n_108),
.B2(n_102),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_150),
.A2(n_153),
.B1(n_168),
.B2(n_138),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_SL g182 ( 
.A1(n_151),
.A2(n_159),
.B(n_162),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_128),
.B(n_85),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_135),
.A2(n_81),
.B1(n_88),
.B2(n_104),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_115),
.B(n_86),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_154),
.B(n_157),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_128),
.A2(n_92),
.B1(n_96),
.B2(n_94),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_155),
.A2(n_167),
.B1(n_172),
.B2(n_173),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_132),
.B(n_112),
.Y(n_156)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_156),
.Y(n_190)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_123),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_132),
.B(n_99),
.Y(n_158)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_158),
.Y(n_205)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_113),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_160),
.B(n_166),
.Y(n_189)
);

FAx1_ASAP7_75t_SL g161 ( 
.A(n_121),
.B(n_111),
.CI(n_2),
.CON(n_161),
.SN(n_161)
);

XNOR2x1_ASAP7_75t_SL g208 ( 
.A(n_161),
.B(n_5),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_134),
.B(n_1),
.Y(n_162)
);

OAI21xp33_ASAP7_75t_L g196 ( 
.A1(n_163),
.A2(n_1),
.B(n_3),
.Y(n_196)
);

BUFx2_ASAP7_75t_L g166 ( 
.A(n_126),
.Y(n_166)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_113),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_169),
.B(n_170),
.Y(n_197)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_137),
.Y(n_170)
);

INVx1_ASAP7_75t_SL g171 ( 
.A(n_119),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_171),
.B(n_174),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_121),
.A2(n_80),
.B1(n_3),
.B2(n_4),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_L g173 ( 
.A1(n_133),
.A2(n_80),
.B1(n_3),
.B2(n_4),
.Y(n_173)
);

INVx4_ASAP7_75t_L g174 ( 
.A(n_141),
.Y(n_174)
);

AND2x2_ASAP7_75t_L g175 ( 
.A(n_131),
.B(n_1),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_SL g184 ( 
.A1(n_175),
.A2(n_114),
.B(n_117),
.Y(n_184)
);

BUFx24_ASAP7_75t_SL g176 ( 
.A(n_117),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_176),
.B(n_126),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_171),
.A2(n_147),
.B1(n_172),
.B2(n_165),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_177),
.A2(n_181),
.B1(n_195),
.B2(n_198),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_165),
.A2(n_130),
.B1(n_114),
.B2(n_133),
.Y(n_181)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_155),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_183),
.B(n_191),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_SL g214 ( 
.A(n_184),
.B(n_186),
.C(n_196),
.Y(n_214)
);

OA21x2_ASAP7_75t_L g186 ( 
.A1(n_159),
.A2(n_137),
.B(n_127),
.Y(n_186)
);

INVxp67_ASAP7_75t_L g191 ( 
.A(n_156),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_L g192 ( 
.A1(n_148),
.A2(n_138),
.B(n_134),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_L g212 ( 
.A1(n_192),
.A2(n_199),
.B(n_175),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_L g223 ( 
.A1(n_193),
.A2(n_170),
.B1(n_166),
.B2(n_8),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_144),
.B(n_142),
.C(n_136),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_194),
.B(n_207),
.C(n_209),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_144),
.A2(n_123),
.B1(n_139),
.B2(n_127),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_151),
.A2(n_123),
.B1(n_139),
.B2(n_136),
.Y(n_198)
);

AND2x2_ASAP7_75t_L g199 ( 
.A(n_150),
.B(n_124),
.Y(n_199)
);

A2O1A1Ixp33_ASAP7_75t_SL g200 ( 
.A1(n_161),
.A2(n_137),
.B(n_6),
.C(n_7),
.Y(n_200)
);

OAI22x1_ASAP7_75t_L g216 ( 
.A1(n_200),
.A2(n_208),
.B1(n_186),
.B2(n_184),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_202),
.B(n_209),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_174),
.B(n_116),
.Y(n_203)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_203),
.Y(n_219)
);

BUFx6f_ASAP7_75t_L g204 ( 
.A(n_157),
.Y(n_204)
);

BUFx6f_ASAP7_75t_L g229 ( 
.A(n_204),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_161),
.A2(n_140),
.B1(n_116),
.B2(n_122),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_206),
.A2(n_6),
.B1(n_8),
.B2(n_181),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_146),
.B(n_140),
.C(n_122),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_SL g217 ( 
.A(n_208),
.B(n_175),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_162),
.B(n_5),
.Y(n_209)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_204),
.Y(n_210)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_210),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_182),
.A2(n_158),
.B1(n_164),
.B2(n_169),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_211),
.A2(n_223),
.B1(n_225),
.B2(n_185),
.Y(n_251)
);

MAJx2_ASAP7_75t_L g259 ( 
.A(n_212),
.B(n_192),
.C(n_199),
.Y(n_259)
);

INVx13_ASAP7_75t_L g213 ( 
.A(n_204),
.Y(n_213)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_213),
.Y(n_239)
);

BUFx5_ASAP7_75t_L g215 ( 
.A(n_186),
.Y(n_215)
);

CKINVDCx16_ASAP7_75t_R g253 ( 
.A(n_215),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_L g243 ( 
.A1(n_216),
.A2(n_200),
.B1(n_193),
.B2(n_199),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_SL g249 ( 
.A(n_217),
.B(n_227),
.Y(n_249)
);

OAI21xp5_ASAP7_75t_L g220 ( 
.A1(n_201),
.A2(n_160),
.B(n_153),
.Y(n_220)
);

AOI21xp5_ASAP7_75t_L g246 ( 
.A1(n_220),
.A2(n_231),
.B(n_235),
.Y(n_246)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_189),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_221),
.B(n_222),
.Y(n_237)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_197),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_191),
.B(n_5),
.Y(n_224)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_224),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_183),
.A2(n_5),
.B1(n_6),
.B2(n_8),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_188),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_226),
.B(n_228),
.Y(n_250)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_180),
.Y(n_228)
);

NOR2xp67_ASAP7_75t_SL g230 ( 
.A(n_200),
.B(n_8),
.Y(n_230)
);

AOI21xp33_ASAP7_75t_L g256 ( 
.A1(n_230),
.A2(n_214),
.B(n_217),
.Y(n_256)
);

AOI21xp5_ASAP7_75t_SL g231 ( 
.A1(n_182),
.A2(n_179),
.B(n_178),
.Y(n_231)
);

INVxp67_ASAP7_75t_L g233 ( 
.A(n_177),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_233),
.B(n_236),
.Y(n_257)
);

OAI21xp5_ASAP7_75t_L g235 ( 
.A1(n_179),
.A2(n_178),
.B(n_200),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_234),
.B(n_207),
.C(n_194),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_240),
.B(n_241),
.C(n_248),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_234),
.B(n_212),
.C(n_218),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_243),
.A2(n_254),
.B1(n_229),
.B2(n_253),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_211),
.B(n_206),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_244),
.B(n_249),
.Y(n_275)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_232),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_245),
.B(n_255),
.Y(n_276)
);

NAND3xp33_ASAP7_75t_L g247 ( 
.A(n_216),
.B(n_190),
.C(n_205),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_247),
.B(n_251),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_218),
.B(n_190),
.C(n_205),
.Y(n_248)
);

NAND3xp33_ASAP7_75t_L g252 ( 
.A(n_214),
.B(n_200),
.C(n_187),
.Y(n_252)
);

OAI21xp5_ASAP7_75t_SL g264 ( 
.A1(n_252),
.A2(n_256),
.B(n_258),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_233),
.A2(n_215),
.B1(n_227),
.B2(n_231),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_224),
.Y(n_255)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_220),
.Y(n_258)
);

MAJx2_ASAP7_75t_L g274 ( 
.A(n_259),
.B(n_249),
.C(n_246),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_241),
.B(n_235),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_260),
.B(n_274),
.Y(n_279)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_237),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_261),
.B(n_263),
.Y(n_287)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_237),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_240),
.B(n_219),
.C(n_195),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_265),
.B(n_266),
.C(n_267),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_248),
.B(n_222),
.C(n_210),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_258),
.B(n_229),
.C(n_213),
.Y(n_267)
);

HB1xp67_ASAP7_75t_L g268 ( 
.A(n_239),
.Y(n_268)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_268),
.Y(n_282)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_250),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_269),
.B(n_270),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_SL g271 ( 
.A(n_250),
.B(n_257),
.Y(n_271)
);

CKINVDCx14_ASAP7_75t_R g289 ( 
.A(n_271),
.Y(n_289)
);

INVxp67_ASAP7_75t_L g273 ( 
.A(n_257),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_273),
.B(n_278),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_275),
.B(n_277),
.Y(n_291)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_244),
.B(n_246),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_254),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_276),
.B(n_242),
.Y(n_284)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_284),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_273),
.B(n_242),
.Y(n_285)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_285),
.Y(n_302)
);

BUFx12_ASAP7_75t_L g286 ( 
.A(n_274),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_286),
.B(n_288),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_267),
.Y(n_288)
);

OAI22x1_ASAP7_75t_L g290 ( 
.A1(n_277),
.A2(n_264),
.B1(n_259),
.B2(n_251),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_290),
.A2(n_281),
.B1(n_284),
.B2(n_287),
.Y(n_303)
);

INVx5_ASAP7_75t_L g292 ( 
.A(n_266),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_292),
.B(n_293),
.Y(n_305)
);

BUFx2_ASAP7_75t_L g293 ( 
.A(n_272),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_279),
.B(n_262),
.Y(n_295)
);

XOR2xp5_ASAP7_75t_L g314 ( 
.A(n_295),
.B(n_303),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_L g297 ( 
.A1(n_290),
.A2(n_245),
.B1(n_265),
.B2(n_255),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_297),
.B(n_300),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_280),
.B(n_262),
.C(n_275),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_298),
.B(n_299),
.C(n_304),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_280),
.B(n_260),
.C(n_238),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_SL g300 ( 
.A(n_289),
.B(n_283),
.Y(n_300)
);

OR2x2_ASAP7_75t_L g301 ( 
.A(n_281),
.B(n_285),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_301),
.B(n_306),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_279),
.B(n_292),
.C(n_282),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g306 ( 
.A(n_291),
.B(n_286),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_294),
.A2(n_286),
.B1(n_291),
.B2(n_293),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_L g321 ( 
.A1(n_307),
.A2(n_312),
.B1(n_311),
.B2(n_309),
.Y(n_321)
);

INVx11_ASAP7_75t_L g311 ( 
.A(n_301),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_311),
.A2(n_309),
.B1(n_315),
.B2(n_313),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_SL g312 ( 
.A1(n_296),
.A2(n_302),
.B1(n_304),
.B2(n_305),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_299),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_313),
.B(n_315),
.C(n_295),
.Y(n_319)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_306),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_SL g316 ( 
.A(n_314),
.B(n_307),
.Y(n_316)
);

AOI21xp5_ASAP7_75t_L g322 ( 
.A1(n_316),
.A2(n_319),
.B(n_320),
.Y(n_322)
);

INVxp67_ASAP7_75t_L g324 ( 
.A(n_317),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_L g318 ( 
.A(n_314),
.B(n_298),
.Y(n_318)
);

CKINVDCx16_ASAP7_75t_R g323 ( 
.A(n_318),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_310),
.B(n_308),
.Y(n_320)
);

INVxp33_ASAP7_75t_L g325 ( 
.A(n_322),
.Y(n_325)
);

AO221x1_ASAP7_75t_L g327 ( 
.A1(n_325),
.A2(n_326),
.B1(n_310),
.B2(n_319),
.C(n_324),
.Y(n_327)
);

HB1xp67_ASAP7_75t_L g326 ( 
.A(n_323),
.Y(n_326)
);

INVxp67_ASAP7_75t_L g328 ( 
.A(n_327),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_328),
.Y(n_329)
);

OAI21xp5_ASAP7_75t_L g330 ( 
.A1(n_329),
.A2(n_317),
.B(n_321),
.Y(n_330)
);

XOR2xp5_ASAP7_75t_L g331 ( 
.A(n_330),
.B(n_312),
.Y(n_331)
);


endmodule