module fake_jpeg_28101_n_133 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_133);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_133;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_131;
wire n_56;
wire n_79;
wire n_12;
wire n_132;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

INVx8_ASAP7_75t_L g11 ( 
.A(n_4),
.Y(n_11)
);

BUFx3_ASAP7_75t_L g12 ( 
.A(n_3),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_3),
.Y(n_13)
);

INVx6_ASAP7_75t_L g14 ( 
.A(n_10),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_7),
.Y(n_15)
);

INVx4_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

BUFx3_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

BUFx10_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

BUFx8_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_2),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_10),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_8),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_L g24 ( 
.A1(n_14),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_24)
);

OAI22xp33_ASAP7_75t_SL g40 ( 
.A1(n_24),
.A2(n_14),
.B1(n_21),
.B2(n_23),
.Y(n_40)
);

INVx5_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_25),
.Y(n_35)
);

AOI22xp5_ASAP7_75t_SL g26 ( 
.A1(n_14),
.A2(n_16),
.B1(n_13),
.B2(n_19),
.Y(n_26)
);

AOI21xp5_ASAP7_75t_SL g33 ( 
.A1(n_26),
.A2(n_31),
.B(n_13),
.Y(n_33)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_16),
.Y(n_27)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_16),
.Y(n_28)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_SL g37 ( 
.A(n_29),
.B(n_13),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g30 ( 
.A(n_15),
.B(n_0),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_30),
.B(n_15),
.Y(n_34)
);

AOI21xp33_ASAP7_75t_L g31 ( 
.A1(n_15),
.A2(n_0),
.B(n_1),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_30),
.B(n_23),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_32),
.B(n_33),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_34),
.B(n_37),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_27),
.B(n_23),
.Y(n_39)
);

CKINVDCx14_ASAP7_75t_R g48 ( 
.A(n_39),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_40),
.A2(n_22),
.B1(n_21),
.B2(n_19),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_26),
.B(n_18),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_41),
.B(n_24),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_26),
.B(n_22),
.Y(n_42)
);

BUFx24_ASAP7_75t_SL g44 ( 
.A(n_42),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g43 ( 
.A1(n_41),
.A2(n_14),
.B1(n_28),
.B2(n_27),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_43),
.A2(n_29),
.B1(n_25),
.B2(n_11),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_35),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g59 ( 
.A(n_45),
.B(n_54),
.Y(n_59)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_46),
.Y(n_63)
);

INVx13_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_50),
.B(n_56),
.Y(n_61)
);

BUFx10_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_51),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_52),
.B(n_38),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_33),
.B(n_28),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_53),
.B(n_55),
.Y(n_58)
);

NAND3xp33_ASAP7_75t_L g54 ( 
.A(n_34),
.B(n_31),
.C(n_4),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_36),
.B(n_18),
.Y(n_55)
);

CKINVDCx16_ASAP7_75t_R g56 ( 
.A(n_36),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_57),
.A2(n_21),
.B1(n_22),
.B2(n_19),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_60),
.B(n_64),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_62),
.B(n_68),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_53),
.B(n_38),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_65),
.A2(n_73),
.B1(n_50),
.B2(n_46),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_48),
.B(n_17),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_66),
.B(n_69),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_49),
.B(n_17),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_49),
.B(n_17),
.Y(n_69)
);

O2A1O1Ixp33_ASAP7_75t_L g70 ( 
.A1(n_52),
.A2(n_25),
.B(n_11),
.C(n_20),
.Y(n_70)
);

OAI21xp5_ASAP7_75t_SL g87 ( 
.A1(n_70),
.A2(n_73),
.B(n_60),
.Y(n_87)
);

XOR2xp5_ASAP7_75t_L g71 ( 
.A(n_47),
.B(n_17),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_71),
.B(n_20),
.C(n_51),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_47),
.B(n_12),
.Y(n_72)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_72),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_57),
.A2(n_18),
.B1(n_20),
.B2(n_12),
.Y(n_73)
);

AO22x1_ASAP7_75t_L g74 ( 
.A1(n_70),
.A2(n_43),
.B1(n_55),
.B2(n_44),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_74),
.B(n_78),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_75),
.A2(n_82),
.B1(n_51),
.B2(n_20),
.Y(n_95)
);

CKINVDCx16_ASAP7_75t_R g76 ( 
.A(n_61),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_76),
.B(n_83),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_58),
.B(n_56),
.Y(n_78)
);

AOI21xp5_ASAP7_75t_L g80 ( 
.A1(n_58),
.A2(n_45),
.B(n_50),
.Y(n_80)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_80),
.Y(n_99)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_63),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_81),
.B(n_63),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_64),
.A2(n_46),
.B1(n_18),
.B2(n_20),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_65),
.Y(n_83)
);

XNOR2xp5_ASAP7_75t_L g93 ( 
.A(n_86),
.B(n_67),
.Y(n_93)
);

OAI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_87),
.A2(n_59),
.B1(n_18),
.B2(n_20),
.Y(n_96)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_88),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_L g89 ( 
.A1(n_83),
.A2(n_62),
.B1(n_71),
.B2(n_68),
.Y(n_89)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_89),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_85),
.B(n_76),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_91),
.B(n_94),
.Y(n_102)
);

XNOR2xp5_ASAP7_75t_L g106 ( 
.A(n_93),
.B(n_98),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_85),
.B(n_67),
.Y(n_94)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_95),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_L g105 ( 
.A1(n_96),
.A2(n_80),
.B(n_86),
.Y(n_105)
);

AOI322xp5_ASAP7_75t_SL g97 ( 
.A1(n_79),
.A2(n_59),
.A3(n_5),
.B1(n_6),
.B2(n_7),
.C1(n_8),
.C2(n_9),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_97),
.Y(n_100)
);

A2O1A1O1Ixp25_ASAP7_75t_L g98 ( 
.A1(n_87),
.A2(n_18),
.B(n_12),
.C(n_51),
.D(n_7),
.Y(n_98)
);

HB1xp67_ASAP7_75t_L g101 ( 
.A(n_92),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_L g115 ( 
.A(n_101),
.B(n_82),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_105),
.A2(n_108),
.B1(n_99),
.B2(n_95),
.Y(n_109)
);

AOI21xp5_ASAP7_75t_L g108 ( 
.A1(n_99),
.A2(n_78),
.B(n_75),
.Y(n_108)
);

XOR2xp5_ASAP7_75t_L g117 ( 
.A(n_109),
.B(n_114),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_104),
.A2(n_90),
.B1(n_84),
.B2(n_91),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_110),
.B(n_111),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_106),
.B(n_93),
.C(n_105),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_106),
.B(n_92),
.C(n_77),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_112),
.B(n_113),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_103),
.B(n_84),
.C(n_77),
.Y(n_113)
);

XOR2xp5_ASAP7_75t_L g114 ( 
.A(n_108),
.B(n_90),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_L g120 ( 
.A1(n_115),
.A2(n_107),
.B(n_81),
.Y(n_120)
);

OAI21x1_ASAP7_75t_L g119 ( 
.A1(n_114),
.A2(n_102),
.B(n_98),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_L g122 ( 
.A(n_119),
.B(n_120),
.Y(n_122)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_117),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_121),
.B(n_123),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_SL g123 ( 
.A1(n_116),
.A2(n_100),
.B(n_111),
.Y(n_123)
);

MAJx2_ASAP7_75t_L g124 ( 
.A(n_117),
.B(n_112),
.C(n_74),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_124),
.B(n_51),
.C(n_9),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_118),
.A2(n_74),
.B1(n_5),
.B2(n_6),
.Y(n_125)
);

AOI322xp5_ASAP7_75t_L g126 ( 
.A1(n_125),
.A2(n_74),
.A3(n_5),
.B1(n_8),
.B2(n_9),
.C1(n_10),
.C2(n_18),
.Y(n_126)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_126),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_127),
.B(n_129),
.C(n_124),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_122),
.B(n_0),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_131),
.B(n_128),
.C(n_130),
.Y(n_132)
);

FAx1_ASAP7_75t_SL g133 ( 
.A(n_132),
.B(n_128),
.CI(n_131),
.CON(n_133),
.SN(n_133)
);


endmodule