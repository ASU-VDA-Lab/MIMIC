module fake_ariane_1842_n_187 (n_8, n_24, n_7, n_22, n_1, n_6, n_13, n_20, n_17, n_4, n_2, n_18, n_9, n_11, n_3, n_14, n_0, n_19, n_16, n_5, n_12, n_15, n_21, n_23, n_10, n_25, n_187);

input n_8;
input n_24;
input n_7;
input n_22;
input n_1;
input n_6;
input n_13;
input n_20;
input n_17;
input n_4;
input n_2;
input n_18;
input n_9;
input n_11;
input n_3;
input n_14;
input n_0;
input n_19;
input n_16;
input n_5;
input n_12;
input n_15;
input n_21;
input n_23;
input n_10;
input n_25;

output n_187;

wire n_83;
wire n_56;
wire n_60;
wire n_170;
wire n_160;
wire n_64;
wire n_180;
wire n_179;
wire n_119;
wire n_124;
wire n_167;
wire n_90;
wire n_38;
wire n_47;
wire n_110;
wire n_153;
wire n_86;
wire n_75;
wire n_89;
wire n_67;
wire n_176;
wire n_149;
wire n_34;
wire n_158;
wire n_172;
wire n_69;
wire n_95;
wire n_175;
wire n_92;
wire n_143;
wire n_183;
wire n_150;
wire n_98;
wire n_74;
wire n_113;
wire n_114;
wire n_33;
wire n_40;
wire n_181;
wire n_152;
wire n_120;
wire n_169;
wire n_106;
wire n_53;
wire n_173;
wire n_111;
wire n_115;
wire n_133;
wire n_66;
wire n_71;
wire n_109;
wire n_96;
wire n_156;
wire n_49;
wire n_174;
wire n_100;
wire n_50;
wire n_132;
wire n_62;
wire n_147;
wire n_51;
wire n_166;
wire n_76;
wire n_103;
wire n_79;
wire n_26;
wire n_46;
wire n_84;
wire n_36;
wire n_91;
wire n_159;
wire n_107;
wire n_72;
wire n_105;
wire n_128;
wire n_44;
wire n_30;
wire n_82;
wire n_178;
wire n_31;
wire n_42;
wire n_57;
wire n_131;
wire n_70;
wire n_117;
wire n_139;
wire n_165;
wire n_85;
wire n_130;
wire n_144;
wire n_48;
wire n_94;
wire n_101;
wire n_134;
wire n_185;
wire n_32;
wire n_37;
wire n_58;
wire n_65;
wire n_123;
wire n_138;
wire n_112;
wire n_45;
wire n_162;
wire n_129;
wire n_126;
wire n_137;
wire n_122;
wire n_148;
wire n_164;
wire n_52;
wire n_157;
wire n_184;
wire n_177;
wire n_135;
wire n_73;
wire n_77;
wire n_171;
wire n_118;
wire n_93;
wire n_121;
wire n_61;
wire n_108;
wire n_102;
wire n_182;
wire n_125;
wire n_168;
wire n_43;
wire n_81;
wire n_87;
wire n_27;
wire n_29;
wire n_41;
wire n_140;
wire n_55;
wire n_151;
wire n_136;
wire n_28;
wire n_80;
wire n_146;
wire n_97;
wire n_154;
wire n_142;
wire n_161;
wire n_163;
wire n_88;
wire n_186;
wire n_141;
wire n_68;
wire n_116;
wire n_104;
wire n_145;
wire n_78;
wire n_39;
wire n_59;
wire n_63;
wire n_99;
wire n_155;
wire n_127;
wire n_35;
wire n_54;

INVx1_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_16),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_21),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_22),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_19),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_18),
.Y(n_32)
);

INVxp67_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

BUFx2_ASAP7_75t_L g35 ( 
.A(n_6),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_3),
.Y(n_36)
);

CKINVDCx16_ASAP7_75t_R g37 ( 
.A(n_7),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_15),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_13),
.Y(n_39)
);

NOR2xp67_ASAP7_75t_L g40 ( 
.A(n_10),
.B(n_9),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_23),
.Y(n_41)
);

HB1xp67_ASAP7_75t_L g42 ( 
.A(n_24),
.Y(n_42)
);

INVx1_ASAP7_75t_SL g43 ( 
.A(n_13),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_25),
.Y(n_44)
);

CKINVDCx5p33_ASAP7_75t_R g45 ( 
.A(n_17),
.Y(n_45)
);

BUFx2_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

INVxp67_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_27),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_27),
.Y(n_49)
);

AND2x4_ASAP7_75t_L g50 ( 
.A(n_31),
.B(n_0),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_37),
.B(n_0),
.Y(n_51)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_28),
.Y(n_52)
);

OR2x2_ASAP7_75t_SL g53 ( 
.A(n_42),
.B(n_1),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_28),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_30),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_30),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_32),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_32),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_44),
.B(n_1),
.Y(n_59)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_44),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_31),
.Y(n_61)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_34),
.B(n_2),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_38),
.B(n_2),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_34),
.Y(n_64)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_41),
.Y(n_65)
);

AND2x4_ASAP7_75t_L g66 ( 
.A(n_36),
.B(n_3),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_57),
.Y(n_67)
);

AO22x2_ASAP7_75t_L g68 ( 
.A1(n_53),
.A2(n_36),
.B1(n_26),
.B2(n_39),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_57),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_57),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_48),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_47),
.B(n_45),
.Y(n_72)
);

INVxp67_ASAP7_75t_L g73 ( 
.A(n_46),
.Y(n_73)
);

INVx2_ASAP7_75t_SL g74 ( 
.A(n_46),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_48),
.Y(n_75)
);

NAND2x1p5_ASAP7_75t_L g76 ( 
.A(n_62),
.B(n_43),
.Y(n_76)
);

NAND3xp33_ASAP7_75t_SL g77 ( 
.A(n_51),
.B(n_33),
.C(n_29),
.Y(n_77)
);

BUFx8_ASAP7_75t_L g78 ( 
.A(n_62),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_49),
.Y(n_79)
);

AO22x2_ASAP7_75t_L g80 ( 
.A1(n_53),
.A2(n_40),
.B1(n_6),
.B2(n_7),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_49),
.Y(n_81)
);

AO22x2_ASAP7_75t_L g82 ( 
.A1(n_53),
.A2(n_5),
.B1(n_8),
.B2(n_9),
.Y(n_82)
);

A2O1A1Ixp33_ASAP7_75t_L g83 ( 
.A1(n_50),
.A2(n_45),
.B(n_8),
.C(n_11),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_71),
.B(n_62),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_75),
.B(n_56),
.Y(n_85)
);

NAND2x1p5_ASAP7_75t_L g86 ( 
.A(n_67),
.B(n_60),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_69),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_79),
.B(n_64),
.Y(n_88)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_70),
.Y(n_89)
);

INVxp33_ASAP7_75t_SL g90 ( 
.A(n_68),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_81),
.B(n_56),
.Y(n_91)
);

BUFx8_ASAP7_75t_L g92 ( 
.A(n_74),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_83),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_72),
.B(n_55),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_76),
.A2(n_47),
.B1(n_59),
.B2(n_63),
.Y(n_95)
);

HB1xp67_ASAP7_75t_L g96 ( 
.A(n_93),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_93),
.B(n_68),
.Y(n_97)
);

OR2x2_ASAP7_75t_L g98 ( 
.A(n_95),
.B(n_73),
.Y(n_98)
);

CKINVDCx6p67_ASAP7_75t_R g99 ( 
.A(n_94),
.Y(n_99)
);

OAI21x1_ASAP7_75t_SL g100 ( 
.A1(n_85),
.A2(n_59),
.B(n_63),
.Y(n_100)
);

BUFx12f_ASAP7_75t_L g101 ( 
.A(n_92),
.Y(n_101)
);

AND2x4_ASAP7_75t_L g102 ( 
.A(n_84),
.B(n_50),
.Y(n_102)
);

CKINVDCx5p33_ASAP7_75t_R g103 ( 
.A(n_92),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_96),
.B(n_84),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_98),
.A2(n_95),
.B1(n_90),
.B2(n_68),
.Y(n_105)
);

AND2x4_ASAP7_75t_L g106 ( 
.A(n_102),
.B(n_88),
.Y(n_106)
);

OR2x2_ASAP7_75t_L g107 ( 
.A(n_98),
.B(n_76),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_L g108 ( 
.A1(n_97),
.A2(n_77),
.B1(n_80),
.B2(n_82),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_96),
.B(n_88),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_L g110 ( 
.A1(n_102),
.A2(n_86),
.B(n_87),
.Y(n_110)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_104),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_104),
.Y(n_112)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_109),
.Y(n_113)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_106),
.Y(n_114)
);

OR2x2_ASAP7_75t_L g115 ( 
.A(n_107),
.B(n_98),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_115),
.B(n_105),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_111),
.Y(n_117)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_112),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_113),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_115),
.B(n_107),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_114),
.Y(n_121)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_114),
.Y(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_114),
.Y(n_123)
);

AND4x1_ASAP7_75t_L g124 ( 
.A(n_111),
.B(n_108),
.C(n_82),
.D(n_80),
.Y(n_124)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_111),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_113),
.B(n_106),
.Y(n_126)
);

INVx1_ASAP7_75t_SL g127 ( 
.A(n_120),
.Y(n_127)
);

AND2x2_ASAP7_75t_L g128 ( 
.A(n_118),
.B(n_82),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_117),
.Y(n_129)
);

INVx1_ASAP7_75t_SL g130 ( 
.A(n_126),
.Y(n_130)
);

OR2x2_ASAP7_75t_L g131 ( 
.A(n_116),
.B(n_97),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_116),
.B(n_80),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_119),
.B(n_106),
.Y(n_133)
);

AND2x2_ASAP7_75t_L g134 ( 
.A(n_118),
.B(n_110),
.Y(n_134)
);

BUFx2_ASAP7_75t_L g135 ( 
.A(n_129),
.Y(n_135)
);

OR2x2_ASAP7_75t_L g136 ( 
.A(n_127),
.B(n_119),
.Y(n_136)
);

NOR2x1p5_ASAP7_75t_SL g137 ( 
.A(n_129),
.B(n_122),
.Y(n_137)
);

NAND2x1_ASAP7_75t_L g138 ( 
.A(n_134),
.B(n_121),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_127),
.B(n_122),
.Y(n_139)
);

INVx1_ASAP7_75t_SL g140 ( 
.A(n_130),
.Y(n_140)
);

OR2x2_ASAP7_75t_L g141 ( 
.A(n_131),
.B(n_117),
.Y(n_141)
);

AND2x2_ASAP7_75t_L g142 ( 
.A(n_134),
.B(n_125),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_128),
.B(n_124),
.Y(n_143)
);

AOI21xp5_ASAP7_75t_L g144 ( 
.A1(n_133),
.A2(n_121),
.B(n_100),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_132),
.B(n_123),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_142),
.B(n_128),
.Y(n_146)
);

AND2x4_ASAP7_75t_SL g147 ( 
.A(n_145),
.B(n_99),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_135),
.B(n_55),
.Y(n_148)
);

AOI21xp5_ASAP7_75t_L g149 ( 
.A1(n_138),
.A2(n_100),
.B(n_77),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_145),
.B(n_58),
.Y(n_150)
);

AND2x2_ASAP7_75t_L g151 ( 
.A(n_141),
.B(n_131),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_136),
.B(n_58),
.Y(n_152)
);

OR2x2_ASAP7_75t_L g153 ( 
.A(n_140),
.B(n_65),
.Y(n_153)
);

INVx1_ASAP7_75t_SL g154 ( 
.A(n_139),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_137),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_151),
.B(n_144),
.Y(n_156)
);

NAND4xp25_ASAP7_75t_L g157 ( 
.A(n_148),
.B(n_144),
.C(n_66),
.D(n_50),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_155),
.Y(n_158)
);

NAND3xp33_ASAP7_75t_L g159 ( 
.A(n_150),
.B(n_58),
.C(n_54),
.Y(n_159)
);

AND2x2_ASAP7_75t_L g160 ( 
.A(n_146),
.B(n_143),
.Y(n_160)
);

INVx1_ASAP7_75t_SL g161 ( 
.A(n_153),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_154),
.Y(n_162)
);

AND2x2_ASAP7_75t_L g163 ( 
.A(n_150),
.B(n_64),
.Y(n_163)
);

HB1xp67_ASAP7_75t_L g164 ( 
.A(n_152),
.Y(n_164)
);

NAND3xp33_ASAP7_75t_L g165 ( 
.A(n_158),
.B(n_152),
.C(n_149),
.Y(n_165)
);

NOR2x1p5_ASAP7_75t_L g166 ( 
.A(n_156),
.B(n_101),
.Y(n_166)
);

AOI221xp5_ASAP7_75t_L g167 ( 
.A1(n_158),
.A2(n_50),
.B1(n_66),
.B2(n_54),
.C(n_58),
.Y(n_167)
);

OR2x2_ASAP7_75t_L g168 ( 
.A(n_164),
.B(n_147),
.Y(n_168)
);

OAI22xp33_ASAP7_75t_SL g169 ( 
.A1(n_161),
.A2(n_103),
.B1(n_61),
.B2(n_65),
.Y(n_169)
);

OAI321xp33_ASAP7_75t_L g170 ( 
.A1(n_157),
.A2(n_61),
.A3(n_58),
.B1(n_65),
.B2(n_91),
.C(n_78),
.Y(n_170)
);

NAND3xp33_ASAP7_75t_L g171 ( 
.A(n_162),
.B(n_58),
.C(n_52),
.Y(n_171)
);

OAI22x1_ASAP7_75t_L g172 ( 
.A1(n_160),
.A2(n_66),
.B1(n_50),
.B2(n_52),
.Y(n_172)
);

OAI211xp5_ASAP7_75t_SL g173 ( 
.A1(n_165),
.A2(n_168),
.B(n_167),
.C(n_171),
.Y(n_173)
);

NOR2x1_ASAP7_75t_L g174 ( 
.A(n_166),
.B(n_163),
.Y(n_174)
);

NAND4xp75_ASAP7_75t_L g175 ( 
.A(n_169),
.B(n_163),
.C(n_160),
.D(n_101),
.Y(n_175)
);

AOI221xp5_ASAP7_75t_L g176 ( 
.A1(n_170),
.A2(n_66),
.B1(n_58),
.B2(n_60),
.C(n_52),
.Y(n_176)
);

OAI211xp5_ASAP7_75t_L g177 ( 
.A1(n_172),
.A2(n_159),
.B(n_60),
.C(n_52),
.Y(n_177)
);

OAI22x1_ASAP7_75t_SL g178 ( 
.A1(n_169),
.A2(n_92),
.B1(n_60),
.B2(n_101),
.Y(n_178)
);

OR2x2_ASAP7_75t_L g179 ( 
.A(n_168),
.B(n_5),
.Y(n_179)
);

AOI211xp5_ASAP7_75t_L g180 ( 
.A1(n_165),
.A2(n_66),
.B(n_12),
.C(n_14),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_180),
.A2(n_102),
.B1(n_14),
.B2(n_11),
.Y(n_181)
);

AND4x1_ASAP7_75t_L g182 ( 
.A(n_174),
.B(n_89),
.C(n_87),
.D(n_100),
.Y(n_182)
);

AOI221xp5_ASAP7_75t_L g183 ( 
.A1(n_173),
.A2(n_89),
.B1(n_102),
.B2(n_86),
.C(n_99),
.Y(n_183)
);

AOI221xp5_ASAP7_75t_L g184 ( 
.A1(n_176),
.A2(n_102),
.B1(n_86),
.B2(n_99),
.C(n_20),
.Y(n_184)
);

AOI21xp5_ASAP7_75t_L g185 ( 
.A1(n_181),
.A2(n_177),
.B(n_178),
.Y(n_185)
);

AOI21xp33_ASAP7_75t_L g186 ( 
.A1(n_185),
.A2(n_183),
.B(n_179),
.Y(n_186)
);

AOI221xp5_ASAP7_75t_L g187 ( 
.A1(n_186),
.A2(n_184),
.B1(n_182),
.B2(n_175),
.C(n_102),
.Y(n_187)
);


endmodule