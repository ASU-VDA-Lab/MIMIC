module fake_jpeg_28923_n_210 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_210);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_210;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_13),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_14),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_0),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

BUFx16f_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_2),
.Y(n_25)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_0),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_6),
.B(n_3),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_3),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_7),
.Y(n_32)
);

BUFx24_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_8),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_2),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_12),
.Y(n_37)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_31),
.Y(n_38)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_38),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_23),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_39),
.B(n_51),
.Y(n_71)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_33),
.Y(n_40)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_40),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_31),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_41),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_28),
.B(n_15),
.Y(n_42)
);

AND2x2_ASAP7_75t_L g60 ( 
.A(n_42),
.B(n_20),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_31),
.Y(n_43)
);

BUFx2_ASAP7_75t_L g70 ( 
.A(n_43),
.Y(n_70)
);

INVx4_ASAP7_75t_SL g44 ( 
.A(n_33),
.Y(n_44)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_44),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_26),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_45),
.Y(n_65)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_46),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_37),
.Y(n_47)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_47),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_48),
.Y(n_79)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_17),
.Y(n_49)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_49),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_26),
.Y(n_50)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_50),
.Y(n_81)
);

BUFx12_ASAP7_75t_L g51 ( 
.A(n_23),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_23),
.Y(n_52)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_52),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_19),
.B(n_25),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_53),
.B(n_35),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_34),
.Y(n_54)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_54),
.Y(n_83)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_33),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_55),
.B(n_57),
.Y(n_80)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_18),
.Y(n_56)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_56),
.Y(n_58)
);

OR2x2_ASAP7_75t_L g57 ( 
.A(n_19),
.B(n_0),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_44),
.A2(n_40),
.B1(n_55),
.B2(n_54),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_59),
.A2(n_67),
.B1(n_72),
.B2(n_74),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_60),
.B(n_62),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_L g61 ( 
.A1(n_47),
.A2(n_36),
.B1(n_29),
.B2(n_18),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_61),
.A2(n_75),
.B1(n_87),
.B2(n_1),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_57),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_40),
.A2(n_34),
.B1(n_36),
.B2(n_33),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_68),
.B(n_84),
.Y(n_90)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_46),
.Y(n_69)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_69),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_55),
.A2(n_36),
.B1(n_35),
.B2(n_32),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_48),
.B(n_32),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_73),
.B(n_30),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_L g75 ( 
.A1(n_41),
.A2(n_29),
.B1(n_22),
.B2(n_27),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_50),
.B(n_16),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_76),
.B(n_13),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_51),
.B(n_16),
.Y(n_84)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_43),
.Y(n_86)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_86),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_38),
.A2(n_30),
.B1(n_27),
.B2(n_25),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_52),
.B(n_22),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_88),
.B(n_24),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_89),
.B(n_95),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_85),
.B(n_21),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_91),
.B(n_96),
.Y(n_117)
);

AND2x4_ASAP7_75t_L g92 ( 
.A(n_67),
.B(n_51),
.Y(n_92)
);

AOI21xp5_ASAP7_75t_L g119 ( 
.A1(n_92),
.A2(n_110),
.B(n_59),
.Y(n_119)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_77),
.Y(n_93)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_93),
.Y(n_136)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_64),
.Y(n_94)
);

BUFx3_ASAP7_75t_L g121 ( 
.A(n_94),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_58),
.B(n_24),
.Y(n_96)
);

CKINVDCx16_ASAP7_75t_R g122 ( 
.A(n_97),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_80),
.B(n_21),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_98),
.B(n_100),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_88),
.B(n_20),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_71),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_103),
.B(n_107),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_60),
.B(n_17),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_104),
.B(n_108),
.Y(n_120)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_75),
.Y(n_105)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_105),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_72),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_106),
.B(n_115),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_66),
.B(n_70),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_70),
.Y(n_109)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_109),
.Y(n_129)
);

NAND2xp33_ASAP7_75t_SL g110 ( 
.A(n_65),
.B(n_45),
.Y(n_110)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_61),
.Y(n_111)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_111),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_112),
.A2(n_79),
.B1(n_78),
.B2(n_83),
.Y(n_133)
);

INVx11_ASAP7_75t_L g113 ( 
.A(n_64),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_113),
.B(n_65),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_82),
.B(n_10),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g134 ( 
.A(n_114),
.B(n_1),
.Y(n_134)
);

BUFx3_ASAP7_75t_L g115 ( 
.A(n_63),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_SL g141 ( 
.A1(n_119),
.A2(n_92),
.B(n_110),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_126),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_90),
.B(n_99),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_127),
.B(n_128),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_99),
.B(n_82),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_96),
.B(n_81),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_131),
.B(n_89),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_105),
.A2(n_81),
.B1(n_79),
.B2(n_78),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_132),
.A2(n_135),
.B1(n_109),
.B2(n_116),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_133),
.A2(n_101),
.B1(n_94),
.B2(n_113),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_SL g145 ( 
.A(n_134),
.B(n_137),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_111),
.A2(n_66),
.B1(n_83),
.B2(n_4),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_98),
.B(n_1),
.Y(n_137)
);

INVxp67_ASAP7_75t_L g164 ( 
.A(n_139),
.Y(n_164)
);

AND2x2_ASAP7_75t_L g165 ( 
.A(n_140),
.B(n_141),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_L g142 ( 
.A1(n_116),
.A2(n_112),
.B1(n_92),
.B2(n_93),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_142),
.A2(n_146),
.B1(n_155),
.B2(n_126),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g143 ( 
.A(n_117),
.B(n_100),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_143),
.B(n_144),
.C(n_120),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_SL g144 ( 
.A1(n_119),
.A2(n_92),
.B(n_91),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_122),
.A2(n_92),
.B1(n_102),
.B2(n_103),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_129),
.Y(n_147)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_147),
.Y(n_158)
);

OR2x4_ASAP7_75t_L g148 ( 
.A(n_130),
.B(n_102),
.Y(n_148)
);

HAxp5_ASAP7_75t_SL g169 ( 
.A(n_148),
.B(n_149),
.CON(n_169),
.SN(n_169)
);

AND2x4_ASAP7_75t_L g149 ( 
.A(n_117),
.B(n_108),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_150),
.A2(n_151),
.B1(n_153),
.B2(n_156),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_122),
.A2(n_104),
.B1(n_114),
.B2(n_107),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_SL g152 ( 
.A(n_125),
.B(n_101),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_152),
.B(n_154),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_133),
.A2(n_115),
.B1(n_4),
.B2(n_5),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_127),
.B(n_9),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_131),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_159),
.B(n_144),
.Y(n_174)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_148),
.Y(n_160)
);

CKINVDCx14_ASAP7_75t_R g173 ( 
.A(n_160),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_L g161 ( 
.A1(n_146),
.A2(n_123),
.B(n_128),
.Y(n_161)
);

AND2x2_ASAP7_75t_L g183 ( 
.A(n_161),
.B(n_162),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_L g162 ( 
.A1(n_141),
.A2(n_130),
.B(n_120),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_163),
.B(n_167),
.Y(n_175)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_140),
.Y(n_166)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_166),
.Y(n_172)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_156),
.Y(n_167)
);

AOI322xp5_ASAP7_75t_SL g168 ( 
.A1(n_145),
.A2(n_134),
.A3(n_125),
.B1(n_124),
.B2(n_118),
.C1(n_135),
.C2(n_132),
.Y(n_168)
);

NOR3xp33_ASAP7_75t_L g177 ( 
.A(n_168),
.B(n_118),
.C(n_124),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_170),
.B(n_171),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_138),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_174),
.B(n_179),
.C(n_180),
.Y(n_186)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_158),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_176),
.B(n_182),
.Y(n_185)
);

OAI322xp33_ASAP7_75t_L g190 ( 
.A1(n_177),
.A2(n_169),
.A3(n_164),
.B1(n_149),
.B2(n_160),
.C1(n_161),
.C2(n_170),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_SL g178 ( 
.A1(n_165),
.A2(n_149),
.B(n_136),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_178),
.B(n_173),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_159),
.B(n_143),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_165),
.B(n_149),
.C(n_129),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_157),
.B(n_155),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_172),
.A2(n_166),
.B1(n_163),
.B2(n_165),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_184),
.A2(n_167),
.B1(n_180),
.B2(n_183),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_178),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_187),
.B(n_189),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_SL g188 ( 
.A(n_174),
.B(n_162),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_188),
.B(n_179),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_181),
.B(n_164),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_190),
.B(n_183),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_191),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_SL g192 ( 
.A1(n_185),
.A2(n_175),
.B(n_183),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_192),
.B(n_194),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_196),
.A2(n_121),
.B1(n_136),
.B2(n_8),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_197),
.B(n_188),
.C(n_186),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_198),
.B(n_199),
.C(n_202),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_194),
.B(n_186),
.C(n_184),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_195),
.B(n_158),
.Y(n_201)
);

AOI21xp5_ASAP7_75t_L g205 ( 
.A1(n_201),
.A2(n_192),
.B(n_196),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_SL g203 ( 
.A(n_201),
.B(n_193),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_203),
.B(n_205),
.Y(n_207)
);

AO21x1_ASAP7_75t_L g206 ( 
.A1(n_204),
.A2(n_200),
.B(n_121),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_L g208 ( 
.A1(n_206),
.A2(n_6),
.B(n_7),
.Y(n_208)
);

AOI21xp5_ASAP7_75t_L g209 ( 
.A1(n_208),
.A2(n_207),
.B(n_8),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_209),
.B(n_9),
.Y(n_210)
);


endmodule