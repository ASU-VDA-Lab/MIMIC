module fake_jpeg_30654_n_108 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_108);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_108;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_106;
wire n_44;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_100;
wire n_82;
wire n_96;

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_31),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_20),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_34),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_19),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_32),
.Y(n_40)
);

BUFx10_ASAP7_75t_L g41 ( 
.A(n_12),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_26),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_21),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_2),
.Y(n_44)
);

INVxp67_ASAP7_75t_L g45 ( 
.A(n_22),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_9),
.Y(n_46)
);

A2O1A1Ixp33_ASAP7_75t_L g47 ( 
.A1(n_45),
.A2(n_14),
.B(n_30),
.C(n_29),
.Y(n_47)
);

NOR2x1_ASAP7_75t_L g55 ( 
.A(n_47),
.B(n_41),
.Y(n_55)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_48),
.B(n_51),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_L g49 ( 
.A1(n_35),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_49),
.B(n_50),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_45),
.B(n_46),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_44),
.B(n_0),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_37),
.B(n_1),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_52),
.B(n_3),
.Y(n_62)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_53),
.Y(n_65)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_43),
.Y(n_54)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_54),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_55),
.B(n_59),
.Y(n_74)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_54),
.Y(n_58)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_58),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_51),
.B(n_41),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_48),
.B(n_41),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_60),
.B(n_63),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_62),
.B(n_66),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_53),
.B(n_44),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_47),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_64),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_51),
.B(n_44),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_56),
.A2(n_35),
.B1(n_40),
.B2(n_39),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_69),
.A2(n_70),
.B1(n_73),
.B2(n_10),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_64),
.A2(n_42),
.B1(n_15),
.B2(n_17),
.Y(n_70)
);

INVx2_ASAP7_75t_R g71 ( 
.A(n_55),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_71),
.B(n_72),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_57),
.B(n_3),
.Y(n_72)
);

OAI21xp33_ASAP7_75t_SL g73 ( 
.A1(n_59),
.A2(n_13),
.B(n_28),
.Y(n_73)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_65),
.Y(n_75)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_75),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_65),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_76),
.A2(n_77),
.B1(n_79),
.B2(n_71),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_61),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_77)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_77),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_61),
.B(n_23),
.C(n_27),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_80),
.B(n_25),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_68),
.B(n_58),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_81),
.B(n_82),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_67),
.B(n_7),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_74),
.B(n_7),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_84),
.B(n_87),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_88),
.Y(n_96)
);

XNOR2xp5_ASAP7_75t_L g95 ( 
.A(n_89),
.B(n_90),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_78),
.B(n_8),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_73),
.A2(n_80),
.B1(n_8),
.B2(n_18),
.Y(n_91)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_91),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_79),
.B(n_11),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_93),
.B(n_85),
.Y(n_98)
);

XOR2xp5_ASAP7_75t_L g101 ( 
.A(n_98),
.B(n_99),
.Y(n_101)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_94),
.B(n_92),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_95),
.B(n_83),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_101),
.B(n_100),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_102),
.B(n_95),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_103),
.A2(n_96),
.B1(n_97),
.B2(n_86),
.Y(n_104)
);

XNOR2xp5_ASAP7_75t_L g105 ( 
.A(n_104),
.B(n_86),
.Y(n_105)
);

HB1xp67_ASAP7_75t_L g106 ( 
.A(n_105),
.Y(n_106)
);

XOR2xp5_ASAP7_75t_L g107 ( 
.A(n_106),
.B(n_24),
.Y(n_107)
);

XOR2xp5_ASAP7_75t_L g108 ( 
.A(n_107),
.B(n_33),
.Y(n_108)
);


endmodule