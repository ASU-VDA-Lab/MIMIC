module real_jpeg_10320_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_247;
wire n_146;
wire n_78;
wire n_83;
wire n_249;
wire n_166;
wire n_176;
wire n_215;
wire n_221;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_271;
wire n_163;
wire n_276;
wire n_22;
wire n_237;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_173;
wire n_105;
wire n_255;
wire n_243;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_275;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_172;
wire n_160;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_148;
wire n_19;
wire n_262;
wire n_222;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_205;
wire n_195;
wire n_258;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_228;
wire n_150;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_278;
wire n_130;
wire n_241;
wire n_103;
wire n_225;
wire n_259;
wire n_232;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_277;
wire n_226;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_216;
wire n_128;
wire n_213;
wire n_167;
wire n_179;
wire n_202;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_274;
wire n_256;
wire n_182;
wire n_253;
wire n_96;
wire n_269;
wire n_273;
wire n_89;

BUFx24_ASAP7_75t_L g58 ( 
.A(n_0),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_1),
.A2(n_52),
.B1(n_60),
.B2(n_61),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_1),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_1),
.A2(n_57),
.B1(n_58),
.B2(n_61),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_1),
.A2(n_26),
.B1(n_29),
.B2(n_61),
.Y(n_208)
);

AOI22xp33_ASAP7_75t_SL g245 ( 
.A1(n_1),
.A2(n_37),
.B1(n_38),
.B2(n_61),
.Y(n_245)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_2),
.A2(n_52),
.B1(n_60),
.B2(n_100),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_2),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g169 ( 
.A1(n_2),
.A2(n_57),
.B1(n_58),
.B2(n_100),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_SL g206 ( 
.A1(n_2),
.A2(n_26),
.B1(n_29),
.B2(n_100),
.Y(n_206)
);

AOI22xp33_ASAP7_75t_SL g237 ( 
.A1(n_2),
.A2(n_37),
.B1(n_38),
.B2(n_100),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g36 ( 
.A1(n_3),
.A2(n_37),
.B1(n_38),
.B2(n_40),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_3),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_3),
.A2(n_40),
.B1(n_57),
.B2(n_58),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_3),
.A2(n_26),
.B1(n_29),
.B2(n_40),
.Y(n_151)
);

BUFx12_ASAP7_75t_L g54 ( 
.A(n_4),
.Y(n_54)
);

BUFx10_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

BUFx10_ASAP7_75t_L g42 ( 
.A(n_7),
.Y(n_42)
);

BUFx6f_ASAP7_75t_SL g69 ( 
.A(n_8),
.Y(n_69)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_9),
.Y(n_39)
);

OAI22xp33_ASAP7_75t_SL g25 ( 
.A1(n_10),
.A2(n_26),
.B1(n_28),
.B2(n_29),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_10),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_10),
.A2(n_28),
.B1(n_57),
.B2(n_58),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_L g86 ( 
.A1(n_10),
.A2(n_28),
.B1(n_37),
.B2(n_38),
.Y(n_86)
);

OAI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_10),
.A2(n_28),
.B1(n_52),
.B2(n_60),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_L g143 ( 
.A1(n_11),
.A2(n_52),
.B1(n_60),
.B2(n_144),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_11),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_11),
.A2(n_57),
.B1(n_58),
.B2(n_144),
.Y(n_192)
);

AOI22xp33_ASAP7_75t_SL g214 ( 
.A1(n_11),
.A2(n_37),
.B1(n_38),
.B2(n_144),
.Y(n_214)
);

AOI22xp33_ASAP7_75t_SL g224 ( 
.A1(n_11),
.A2(n_26),
.B1(n_29),
.B2(n_144),
.Y(n_224)
);

BUFx10_ASAP7_75t_L g52 ( 
.A(n_12),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_13),
.A2(n_37),
.B1(n_38),
.B2(n_47),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_13),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_13),
.A2(n_26),
.B1(n_29),
.B2(n_47),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_13),
.A2(n_47),
.B1(n_57),
.B2(n_58),
.Y(n_118)
);

OAI22xp33_ASAP7_75t_SL g33 ( 
.A1(n_14),
.A2(n_26),
.B1(n_29),
.B2(n_34),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_14),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_14),
.A2(n_34),
.B1(n_52),
.B2(n_60),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_14),
.A2(n_34),
.B1(n_57),
.B2(n_58),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_14),
.A2(n_34),
.B1(n_37),
.B2(n_38),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_15),
.Y(n_148)
);

AOI21xp33_ASAP7_75t_L g149 ( 
.A1(n_15),
.A2(n_54),
.B(n_58),
.Y(n_149)
);

OAI22xp33_ASAP7_75t_SL g172 ( 
.A1(n_15),
.A2(n_52),
.B1(n_60),
.B2(n_148),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_15),
.B(n_64),
.Y(n_193)
);

AOI21xp5_ASAP7_75t_L g212 ( 
.A1(n_15),
.A2(n_37),
.B(n_213),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_15),
.B(n_37),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_15),
.A2(n_80),
.B1(n_81),
.B2(n_224),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_127),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_SL g17 ( 
.A(n_18),
.B(n_125),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_104),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_19),
.B(n_104),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_77),
.C(n_88),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_20),
.A2(n_21),
.B1(n_77),
.B2(n_154),
.Y(n_153)
);

CKINVDCx16_ASAP7_75t_R g20 ( 
.A(n_21),
.Y(n_20)
);

XOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_48),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_22),
.B(n_49),
.C(n_76),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_35),
.Y(n_22)
);

XNOR2xp5_ASAP7_75t_L g133 ( 
.A(n_23),
.B(n_35),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_32),
.Y(n_23)
);

OAI21xp5_ASAP7_75t_L g195 ( 
.A1(n_24),
.A2(n_81),
.B(n_151),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g24 ( 
.A(n_25),
.B(n_30),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_25),
.B(n_31),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_26),
.Y(n_29)
);

AOI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_26),
.A2(n_29),
.B1(n_42),
.B2(n_45),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_26),
.A2(n_216),
.B1(n_217),
.B2(n_218),
.Y(n_215)
);

BUFx24_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_SL g30 ( 
.A(n_29),
.B(n_31),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_SL g216 ( 
.A(n_29),
.B(n_45),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_SL g227 ( 
.A(n_29),
.B(n_228),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_30),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_30),
.A2(n_31),
.B1(n_205),
.B2(n_207),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_31),
.B(n_33),
.Y(n_32)
);

CKINVDCx16_ASAP7_75t_R g81 ( 
.A(n_31),
.Y(n_81)
);

OAI21xp5_ASAP7_75t_SL g238 ( 
.A1(n_32),
.A2(n_80),
.B(n_208),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_33),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g35 ( 
.A1(n_36),
.A2(n_41),
.B1(n_44),
.B2(n_46),
.Y(n_35)
);

OAI21xp5_ASAP7_75t_L g93 ( 
.A1(n_36),
.A2(n_44),
.B(n_94),
.Y(n_93)
);

A2O1A1Ixp33_ASAP7_75t_SL g41 ( 
.A1(n_37),
.A2(n_42),
.B(n_43),
.C(n_44),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_37),
.B(n_42),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_37),
.A2(n_38),
.B1(n_68),
.B2(n_69),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g252 ( 
.A(n_37),
.B(n_68),
.Y(n_252)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_L g251 ( 
.A1(n_38),
.A2(n_73),
.B1(n_247),
.B2(n_252),
.Y(n_251)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

OAI21xp5_ASAP7_75t_SL g83 ( 
.A1(n_41),
.A2(n_46),
.B(n_84),
.Y(n_83)
);

CKINVDCx16_ASAP7_75t_R g96 ( 
.A(n_41),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_41),
.A2(n_44),
.B1(n_212),
.B2(n_214),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_41),
.A2(n_44),
.B1(n_214),
.B2(n_237),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g244 ( 
.A1(n_41),
.A2(n_44),
.B1(n_237),
.B2(n_245),
.Y(n_244)
);

OAI21xp5_ASAP7_75t_SL g267 ( 
.A1(n_41),
.A2(n_120),
.B(n_245),
.Y(n_267)
);

CKINVDCx16_ASAP7_75t_R g45 ( 
.A(n_42),
.Y(n_45)
);

INVxp67_ASAP7_75t_L g218 ( 
.A(n_43),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_44),
.B(n_86),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_44),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g222 ( 
.A(n_44),
.B(n_148),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_49),
.A2(n_50),
.B1(n_65),
.B2(n_76),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_50),
.Y(n_49)
);

OAI21xp5_ASAP7_75t_SL g50 ( 
.A1(n_51),
.A2(n_59),
.B(n_62),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_51),
.A2(n_56),
.B1(n_59),
.B2(n_99),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_SL g109 ( 
.A1(n_51),
.A2(n_110),
.B(n_111),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_51),
.A2(n_56),
.B1(n_99),
.B2(n_143),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_51),
.Y(n_171)
);

A2O1A1Ixp33_ASAP7_75t_L g51 ( 
.A1(n_52),
.A2(n_53),
.B(n_55),
.C(n_56),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_52),
.B(n_53),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_52),
.Y(n_60)
);

A2O1A1Ixp33_ASAP7_75t_L g147 ( 
.A1(n_52),
.A2(n_53),
.B(n_148),
.C(n_149),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g56 ( 
.A1(n_53),
.A2(n_54),
.B1(n_57),
.B2(n_58),
.Y(n_56)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_56),
.Y(n_64)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

O2A1O1Ixp33_ASAP7_75t_L g72 ( 
.A1(n_58),
.A2(n_67),
.B(n_68),
.C(n_73),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_58),
.B(n_68),
.Y(n_73)
);

HAxp5_ASAP7_75t_SL g247 ( 
.A(n_58),
.B(n_148),
.CON(n_247),
.SN(n_247)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_63),
.B(n_64),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_63),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_64),
.B(n_112),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_64),
.A2(n_171),
.B1(n_172),
.B2(n_173),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_65),
.Y(n_76)
);

OAI21xp5_ASAP7_75t_L g65 ( 
.A1(n_66),
.A2(n_70),
.B(n_71),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_66),
.B(n_75),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_66),
.A2(n_138),
.B1(n_139),
.B2(n_169),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_66),
.A2(n_138),
.B1(n_169),
.B2(n_191),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_66),
.B(n_148),
.Y(n_235)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_67),
.A2(n_72),
.B1(n_117),
.B2(n_118),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_67),
.B(n_102),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_67),
.A2(n_72),
.B1(n_192),
.B2(n_247),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_69),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_70),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_72),
.B(n_74),
.Y(n_71)
);

AOI21xp5_ASAP7_75t_L g101 ( 
.A1(n_72),
.A2(n_102),
.B(n_103),
.Y(n_101)
);

CKINVDCx16_ASAP7_75t_R g138 ( 
.A(n_72),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_75),
.Y(n_74)
);

CKINVDCx14_ASAP7_75t_R g154 ( 
.A(n_77),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_78),
.A2(n_79),
.B1(n_83),
.B2(n_87),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_78),
.A2(n_79),
.B1(n_108),
.B2(n_109),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_79),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_79),
.B(n_83),
.Y(n_113)
);

AOI21xp5_ASAP7_75t_L g79 ( 
.A1(n_80),
.A2(n_81),
.B(n_82),
.Y(n_79)
);

OAI21xp5_ASAP7_75t_SL g90 ( 
.A1(n_80),
.A2(n_91),
.B(n_92),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_80),
.A2(n_81),
.B1(n_91),
.B2(n_151),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_80),
.A2(n_81),
.B1(n_206),
.B2(n_224),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_SL g253 ( 
.A1(n_80),
.A2(n_82),
.B(n_92),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_81),
.B(n_148),
.Y(n_228)
);

CKINVDCx14_ASAP7_75t_R g87 ( 
.A(n_83),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_85),
.Y(n_84)
);

AOI21xp5_ASAP7_75t_L g174 ( 
.A1(n_85),
.A2(n_96),
.B(n_122),
.Y(n_174)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_86),
.Y(n_95)
);

XOR2xp5_ASAP7_75t_L g152 ( 
.A(n_88),
.B(n_153),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_97),
.C(n_101),
.Y(n_88)
);

XOR2xp5_ASAP7_75t_L g130 ( 
.A(n_89),
.B(n_131),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_93),
.Y(n_89)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_90),
.B(n_93),
.Y(n_164)
);

AND2x2_ASAP7_75t_L g119 ( 
.A(n_94),
.B(n_120),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_96),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_97),
.A2(n_98),
.B1(n_101),
.B2(n_132),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_98),
.Y(n_97)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_101),
.Y(n_132)
);

BUFx24_ASAP7_75t_SL g279 ( 
.A(n_104),
.Y(n_279)
);

FAx1_ASAP7_75t_SL g104 ( 
.A(n_105),
.B(n_115),
.CI(n_124),
.CON(n_104),
.SN(n_104)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_106),
.A2(n_107),
.B1(n_113),
.B2(n_114),
.Y(n_105)
);

CKINVDCx16_ASAP7_75t_R g106 ( 
.A(n_107),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_109),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_113),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_L g115 ( 
.A1(n_116),
.A2(n_119),
.B(n_123),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_116),
.B(n_119),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_122),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_L g127 ( 
.A1(n_128),
.A2(n_155),
.B(n_278),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_152),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_129),
.B(n_152),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_133),
.C(n_134),
.Y(n_129)
);

XOR2xp5_ASAP7_75t_L g176 ( 
.A(n_130),
.B(n_133),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_134),
.A2(n_135),
.B1(n_176),
.B2(n_177),
.Y(n_175)
);

CKINVDCx14_ASAP7_75t_R g134 ( 
.A(n_135),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_141),
.C(n_145),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_136),
.A2(n_137),
.B1(n_141),
.B2(n_142),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_137),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_SL g137 ( 
.A1(n_138),
.A2(n_139),
.B(n_140),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_142),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_143),
.Y(n_173)
);

XOR2xp5_ASAP7_75t_L g161 ( 
.A(n_145),
.B(n_162),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_150),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_146),
.A2(n_147),
.B1(n_150),
.B2(n_186),
.Y(n_185)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_150),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_197),
.Y(n_155)
);

INVxp33_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

AOI21xp5_ASAP7_75t_L g157 ( 
.A1(n_158),
.A2(n_178),
.B(n_196),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

NOR3xp33_ASAP7_75t_L g197 ( 
.A(n_159),
.B(n_198),
.C(n_277),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_175),
.Y(n_159)
);

AND2x2_ASAP7_75t_L g196 ( 
.A(n_160),
.B(n_175),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_163),
.C(n_165),
.Y(n_160)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_161),
.B(n_180),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_163),
.A2(n_164),
.B1(n_165),
.B2(n_166),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_164),
.Y(n_163)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_170),
.C(n_174),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_167),
.A2(n_168),
.B1(n_174),
.B2(n_184),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_168),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_170),
.B(n_183),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_174),
.Y(n_184)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_176),
.Y(n_177)
);

AND2x2_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_181),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_179),
.B(n_181),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_185),
.C(n_187),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_182),
.B(n_274),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_L g274 ( 
.A1(n_185),
.A2(n_187),
.B1(n_188),
.B2(n_275),
.Y(n_274)
);

CKINVDCx16_ASAP7_75t_R g275 ( 
.A(n_185),
.Y(n_275)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_193),
.C(n_194),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_189),
.A2(n_190),
.B1(n_261),
.B2(n_262),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_190),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_192),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_193),
.A2(n_194),
.B1(n_195),
.B2(n_263),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_193),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_195),
.Y(n_194)
);

AOI21xp5_ASAP7_75t_L g198 ( 
.A1(n_199),
.A2(n_271),
.B(n_276),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_SL g199 ( 
.A1(n_200),
.A2(n_256),
.B(n_270),
.Y(n_199)
);

AOI21xp5_ASAP7_75t_L g200 ( 
.A1(n_201),
.A2(n_240),
.B(n_255),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_SL g201 ( 
.A1(n_202),
.A2(n_231),
.B(n_239),
.Y(n_201)
);

AOI21xp5_ASAP7_75t_L g202 ( 
.A1(n_203),
.A2(n_220),
.B(n_230),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_209),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_SL g230 ( 
.A(n_204),
.B(n_209),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_206),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_208),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_210),
.A2(n_211),
.B1(n_215),
.B2(n_219),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_SL g232 ( 
.A(n_210),
.B(n_219),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_211),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_213),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_215),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_SL g220 ( 
.A1(n_221),
.A2(n_225),
.B(n_229),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_223),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_222),
.B(n_223),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_226),
.B(n_227),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_233),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_232),
.B(n_233),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_234),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_234),
.B(n_241),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_SL g255 ( 
.A(n_234),
.B(n_241),
.Y(n_255)
);

FAx1_ASAP7_75t_SL g234 ( 
.A(n_235),
.B(n_236),
.CI(n_238),
.CON(n_234),
.SN(n_234)
);

AOI22xp33_ASAP7_75t_SL g241 ( 
.A1(n_242),
.A2(n_243),
.B1(n_250),
.B2(n_254),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_L g243 ( 
.A1(n_244),
.A2(n_246),
.B1(n_248),
.B2(n_249),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_244),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_246),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_246),
.B(n_249),
.C(n_254),
.Y(n_257)
);

CKINVDCx14_ASAP7_75t_R g254 ( 
.A(n_250),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_253),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_251),
.B(n_253),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_257),
.B(n_258),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_257),
.B(n_258),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_259),
.A2(n_260),
.B1(n_264),
.B2(n_265),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_259),
.B(n_267),
.C(n_268),
.Y(n_272)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_266),
.A2(n_267),
.B1(n_268),
.B2(n_269),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_266),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_267),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_273),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_SL g276 ( 
.A(n_272),
.B(n_273),
.Y(n_276)
);


endmodule