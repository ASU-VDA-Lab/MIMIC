module fake_netlist_5_584_n_1511 (n_91, n_82, n_122, n_10, n_24, n_124, n_86, n_83, n_61, n_90, n_127, n_75, n_101, n_65, n_78, n_74, n_114, n_57, n_96, n_37, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_60, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_105, n_80, n_4, n_125, n_35, n_128, n_73, n_17, n_92, n_19, n_120, n_30, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_29, n_79, n_47, n_25, n_53, n_8, n_44, n_40, n_34, n_100, n_62, n_71, n_109, n_112, n_85, n_95, n_119, n_59, n_26, n_55, n_99, n_2, n_3, n_49, n_20, n_6, n_39, n_54, n_12, n_67, n_121, n_36, n_76, n_87, n_27, n_64, n_77, n_102, n_106, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_32, n_41, n_104, n_103, n_56, n_51, n_63, n_97, n_11, n_7, n_15, n_48, n_50, n_52, n_88, n_110, n_1511);

input n_91;
input n_82;
input n_122;
input n_10;
input n_24;
input n_124;
input n_86;
input n_83;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_65;
input n_78;
input n_74;
input n_114;
input n_57;
input n_96;
input n_37;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_60;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_105;
input n_80;
input n_4;
input n_125;
input n_35;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_120;
input n_30;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_29;
input n_79;
input n_47;
input n_25;
input n_53;
input n_8;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_71;
input n_109;
input n_112;
input n_85;
input n_95;
input n_119;
input n_59;
input n_26;
input n_55;
input n_99;
input n_2;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_27;
input n_64;
input n_77;
input n_102;
input n_106;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_32;
input n_41;
input n_104;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_11;
input n_7;
input n_15;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_1511;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1166;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1150;
wire n_226;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_155;
wire n_552;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1021;
wire n_551;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1353;
wire n_800;
wire n_1347;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_864;
wire n_173;
wire n_859;
wire n_951;
wire n_1264;
wire n_447;
wire n_247;
wire n_1494;
wire n_292;
wire n_625;
wire n_854;
wire n_1462;
wire n_674;
wire n_417;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_606;
wire n_275;
wire n_877;
wire n_755;
wire n_1118;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1359;
wire n_530;
wire n_150;
wire n_1107;
wire n_556;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_929;
wire n_1124;
wire n_902;
wire n_191;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1257;
wire n_171;
wire n_1182;
wire n_579;
wire n_1261;
wire n_938;
wire n_1098;
wire n_320;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_406;
wire n_519;
wire n_1016;
wire n_1243;
wire n_546;
wire n_1280;
wire n_281;
wire n_240;
wire n_291;
wire n_231;
wire n_257;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_709;
wire n_1490;
wire n_317;
wire n_1236;
wire n_569;
wire n_227;
wire n_920;
wire n_1289;
wire n_335;
wire n_370;
wire n_976;
wire n_343;
wire n_1449;
wire n_308;
wire n_297;
wire n_156;
wire n_1078;
wire n_775;
wire n_219;
wire n_157;
wire n_600;
wire n_1484;
wire n_1374;
wire n_1328;
wire n_223;
wire n_264;
wire n_955;
wire n_163;
wire n_339;
wire n_1146;
wire n_882;
wire n_183;
wire n_243;
wire n_1036;
wire n_1097;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_215;
wire n_350;
wire n_196;
wire n_798;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_290;
wire n_580;
wire n_1040;
wire n_578;
wire n_926;
wire n_344;
wire n_1218;
wire n_422;
wire n_475;
wire n_777;
wire n_1070;
wire n_1030;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_496;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_521;
wire n_663;
wire n_845;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_680;
wire n_1473;
wire n_395;
wire n_164;
wire n_553;
wire n_901;
wire n_813;
wire n_1284;
wire n_214;
wire n_675;
wire n_888;
wire n_1167;
wire n_637;
wire n_1384;
wire n_184;
wire n_446;
wire n_1064;
wire n_144;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_468;
wire n_213;
wire n_342;
wire n_464;
wire n_363;
wire n_197;
wire n_1069;
wire n_1075;
wire n_1450;
wire n_1322;
wire n_1471;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_477;
wire n_571;
wire n_461;
wire n_1211;
wire n_1197;
wire n_907;
wire n_1447;
wire n_1377;
wire n_190;
wire n_989;
wire n_1039;
wire n_228;
wire n_283;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_1463;
wire n_310;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1248;
wire n_230;
wire n_1331;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_476;
wire n_534;
wire n_884;
wire n_345;
wire n_944;
wire n_182;
wire n_143;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_857;
wire n_832;
wire n_207;
wire n_561;
wire n_1319;
wire n_1387;
wire n_1027;
wire n_971;
wire n_1156;
wire n_326;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1199;
wire n_352;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_887;
wire n_154;
wire n_300;
wire n_809;
wire n_870;
wire n_931;
wire n_599;
wire n_1481;
wire n_434;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1293;
wire n_965;
wire n_935;
wire n_1175;
wire n_817;
wire n_360;
wire n_1479;
wire n_759;
wire n_806;
wire n_1477;
wire n_324;
wire n_187;
wire n_1189;
wire n_1259;
wire n_706;
wire n_746;
wire n_747;
wire n_784;
wire n_1244;
wire n_431;
wire n_1194;
wire n_615;
wire n_851;
wire n_843;
wire n_523;
wire n_913;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_776;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_284;
wire n_1128;
wire n_139;
wire n_744;
wire n_590;
wire n_629;
wire n_1308;
wire n_254;
wire n_1233;
wire n_526;
wire n_293;
wire n_372;
wire n_677;
wire n_244;
wire n_1333;
wire n_1121;
wire n_314;
wire n_368;
wire n_433;
wire n_604;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1001;
wire n_1503;
wire n_498;
wire n_1468;
wire n_689;
wire n_738;
wire n_640;
wire n_1510;
wire n_252;
wire n_624;
wire n_1380;
wire n_295;
wire n_133;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_610;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_259;
wire n_448;
wire n_758;
wire n_999;
wire n_1158;
wire n_1509;
wire n_563;
wire n_1145;
wire n_878;
wire n_524;
wire n_204;
wire n_394;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1306;
wire n_1068;
wire n_331;
wire n_906;
wire n_1163;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_658;
wire n_1362;
wire n_456;
wire n_959;
wire n_535;
wire n_152;
wire n_940;
wire n_1445;
wire n_1492;
wire n_592;
wire n_1169;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1269;
wire n_1095;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_1431;
wire n_484;
wire n_1033;
wire n_442;
wire n_131;
wire n_636;
wire n_660;
wire n_1009;
wire n_1148;
wire n_750;
wire n_742;
wire n_995;
wire n_454;
wire n_374;
wire n_185;
wire n_396;
wire n_1383;
wire n_1073;
wire n_255;
wire n_662;
wire n_459;
wire n_218;
wire n_962;
wire n_1215;
wire n_1171;
wire n_723;
wire n_1065;
wire n_1336;
wire n_473;
wire n_1309;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_168;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_208;
wire n_142;
wire n_743;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_1240;
wire n_829;
wire n_1416;
wire n_361;
wire n_1237;
wire n_700;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1006;
wire n_329;
wire n_274;
wire n_1270;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_309;
wire n_512;
wire n_322;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1349;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_224;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_239;
wire n_630;
wire n_504;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_1304;
wire n_1324;
wire n_987;
wire n_261;
wire n_174;
wire n_1455;
wire n_767;
wire n_993;
wire n_1407;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_729;
wire n_1131;
wire n_1084;
wire n_970;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_340;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_233;
wire n_572;
wire n_366;
wire n_815;
wire n_327;
wire n_135;
wire n_1381;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_426;
wire n_1438;
wire n_1082;
wire n_589;
wire n_716;
wire n_562;
wire n_1436;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_531;
wire n_890;
wire n_764;
wire n_1056;
wire n_1424;
wire n_162;
wire n_960;
wire n_222;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_634;
wire n_199;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_256;
wire n_950;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1060;
wire n_1141;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_136;
wire n_146;
wire n_912;
wire n_315;
wire n_968;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_683;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_983;
wire n_280;
wire n_1305;
wire n_873;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_690;
wire n_583;
wire n_302;
wire n_1343;
wire n_1203;
wire n_821;
wire n_321;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1288;
wire n_385;
wire n_212;
wire n_507;
wire n_330;
wire n_1228;
wire n_972;
wire n_692;
wire n_820;
wire n_1200;
wire n_1301;
wire n_1363;
wire n_1185;
wire n_991;
wire n_828;
wire n_779;
wire n_576;
wire n_1143;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_945;
wire n_492;
wire n_153;
wire n_1504;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_286;
wire n_883;
wire n_470;
wire n_325;
wire n_449;
wire n_132;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_856;
wire n_918;
wire n_942;
wire n_189;
wire n_1147;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_195;
wire n_356;
wire n_894;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1470;
wire n_1096;
wire n_234;
wire n_833;
wire n_225;
wire n_1307;
wire n_988;
wire n_814;
wire n_192;
wire n_1201;
wire n_1114;
wire n_655;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_387;
wire n_1149;
wire n_398;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_211;
wire n_1219;
wire n_1204;
wire n_178;
wire n_1035;
wire n_287;
wire n_555;
wire n_783;
wire n_1188;
wire n_661;
wire n_849;
wire n_336;
wire n_584;
wire n_681;
wire n_430;
wire n_510;
wire n_216;
wire n_311;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_445;
wire n_749;
wire n_1134;
wire n_1358;
wire n_717;
wire n_165;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_249;
wire n_304;
wire n_1338;
wire n_577;
wire n_1419;
wire n_338;
wire n_149;
wire n_693;
wire n_1506;
wire n_836;
wire n_990;
wire n_1389;
wire n_975;
wire n_1256;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_151;
wire n_306;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1164;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_876;
wire n_1190;
wire n_601;
wire n_917;
wire n_966;
wire n_253;
wire n_1116;
wire n_1212;
wire n_172;
wire n_206;
wire n_217;
wire n_726;
wire n_982;
wire n_1453;
wire n_818;
wire n_861;
wire n_1183;
wire n_899;
wire n_1253;
wire n_210;
wire n_774;
wire n_1335;
wire n_1059;
wire n_1345;
wire n_176;
wire n_1133;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_1168;
wire n_707;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_665;
wire n_1440;
wire n_177;
wire n_421;
wire n_1356;
wire n_910;
wire n_768;
wire n_1475;
wire n_1302;
wire n_205;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_179;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_735;
wire n_232;
wire n_1109;
wire n_895;
wire n_1310;
wire n_202;
wire n_427;
wire n_1399;
wire n_791;
wire n_732;
wire n_193;
wire n_808;
wire n_797;
wire n_1025;
wire n_500;
wire n_1067;
wire n_148;
wire n_435;
wire n_159;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_594;
wire n_200;
wire n_1291;
wire n_1297;
wire n_1155;
wire n_1418;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_985;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1352;
wire n_626;
wire n_1144;
wire n_1137;
wire n_1170;
wire n_305;
wire n_137;
wire n_676;
wire n_294;
wire n_318;
wire n_653;
wire n_642;
wire n_194;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_268;
wire n_664;
wire n_503;
wire n_235;
wire n_1372;
wire n_605;
wire n_1273;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_840;
wire n_1334;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_581;
wire n_382;
wire n_554;
wire n_898;
wire n_1013;
wire n_1452;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_198;
wire n_714;
wire n_909;
wire n_1497;
wire n_997;
wire n_932;
wire n_612;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_508;
wire n_506;
wire n_1320;
wire n_737;
wire n_986;
wire n_509;
wire n_1317;
wire n_147;
wire n_1281;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_209;
wire n_733;
wire n_1489;
wire n_1376;
wire n_941;
wire n_981;
wire n_867;
wire n_186;
wire n_134;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_518;
wire n_505;
wire n_282;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_381;
wire n_220;
wire n_390;
wire n_1330;
wire n_481;
wire n_769;
wire n_1046;
wire n_271;
wire n_934;
wire n_826;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_167;
wire n_379;
wire n_428;
wire n_1341;
wire n_570;
wire n_1361;
wire n_853;
wire n_377;
wire n_751;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_158;
wire n_704;
wire n_787;
wire n_138;
wire n_961;
wire n_771;
wire n_276;
wire n_1225;
wire n_169;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_181;
wire n_1411;
wire n_221;
wire n_622;
wire n_1087;
wire n_386;
wire n_994;
wire n_848;
wire n_1498;
wire n_1223;
wire n_1272;
wire n_682;
wire n_141;
wire n_1247;
wire n_922;
wire n_816;
wire n_591;
wire n_145;
wire n_1344;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_432;
wire n_839;
wire n_1210;
wire n_1364;
wire n_328;
wire n_140;
wire n_1250;
wire n_369;
wire n_871;
wire n_598;
wire n_685;
wire n_928;
wire n_608;
wire n_1367;
wire n_1460;
wire n_772;
wire n_499;
wire n_517;
wire n_402;
wire n_413;
wire n_1086;
wire n_796;
wire n_236;
wire n_1502;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_903;
wire n_740;
wire n_203;
wire n_384;
wire n_1404;
wire n_1315;
wire n_277;
wire n_1061;
wire n_333;
wire n_1298;
wire n_462;
wire n_1193;
wire n_1255;
wire n_258;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_188;
wire n_844;
wire n_201;
wire n_471;
wire n_852;
wire n_1487;
wire n_1028;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1245;
wire n_846;
wire n_465;
wire n_362;
wire n_1321;
wire n_170;
wire n_161;
wire n_273;
wire n_585;
wire n_270;
wire n_616;
wire n_745;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_641;
wire n_730;
wire n_1325;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_180;
wire n_656;
wire n_1220;
wire n_229;
wire n_437;
wire n_453;
wire n_403;
wire n_1130;
wire n_720;
wire n_863;
wire n_805;
wire n_1275;
wire n_712;
wire n_246;
wire n_1042;
wire n_1402;
wire n_269;
wire n_285;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_251;
wire n_160;
wire n_566;
wire n_565;
wire n_1448;
wire n_1507;
wire n_1398;
wire n_597;
wire n_1181;
wire n_1505;
wire n_1196;
wire n_651;
wire n_1340;
wire n_334;
wire n_811;
wire n_807;
wire n_835;
wire n_175;
wire n_666;
wire n_262;
wire n_1433;
wire n_1254;
wire n_1026;
wire n_1234;
wire n_319;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_242;
wire n_1018;
wire n_438;
wire n_713;
wire n_904;
wire n_166;
wire n_1180;
wire n_1271;
wire n_533;
wire n_1251;
wire n_278;

CKINVDCx5p33_ASAP7_75t_R g131 ( 
.A(n_72),
.Y(n_131)
);

CKINVDCx5p33_ASAP7_75t_R g132 ( 
.A(n_75),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_85),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_0),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_107),
.Y(n_135)
);

CKINVDCx5p33_ASAP7_75t_R g136 ( 
.A(n_65),
.Y(n_136)
);

BUFx3_ASAP7_75t_L g137 ( 
.A(n_68),
.Y(n_137)
);

CKINVDCx5p33_ASAP7_75t_R g138 ( 
.A(n_76),
.Y(n_138)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_82),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_69),
.Y(n_140)
);

CKINVDCx5p33_ASAP7_75t_R g141 ( 
.A(n_84),
.Y(n_141)
);

CKINVDCx5p33_ASAP7_75t_R g142 ( 
.A(n_126),
.Y(n_142)
);

CKINVDCx5p33_ASAP7_75t_R g143 ( 
.A(n_61),
.Y(n_143)
);

INVx2_ASAP7_75t_SL g144 ( 
.A(n_20),
.Y(n_144)
);

CKINVDCx5p33_ASAP7_75t_R g145 ( 
.A(n_11),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_122),
.Y(n_146)
);

CKINVDCx5p33_ASAP7_75t_R g147 ( 
.A(n_8),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_36),
.Y(n_148)
);

CKINVDCx5p33_ASAP7_75t_R g149 ( 
.A(n_23),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_15),
.Y(n_150)
);

CKINVDCx16_ASAP7_75t_R g151 ( 
.A(n_26),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_129),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_124),
.Y(n_153)
);

CKINVDCx5p33_ASAP7_75t_R g154 ( 
.A(n_97),
.Y(n_154)
);

CKINVDCx5p33_ASAP7_75t_R g155 ( 
.A(n_7),
.Y(n_155)
);

CKINVDCx5p33_ASAP7_75t_R g156 ( 
.A(n_77),
.Y(n_156)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_112),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_94),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_40),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_55),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_44),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_115),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_21),
.Y(n_163)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_67),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_51),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_52),
.Y(n_166)
);

INVx2_ASAP7_75t_SL g167 ( 
.A(n_70),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_102),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_39),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_95),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_29),
.Y(n_171)
);

BUFx10_ASAP7_75t_L g172 ( 
.A(n_12),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_125),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_100),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_89),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_103),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_92),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_113),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_62),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_111),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_40),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_130),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_41),
.Y(n_183)
);

BUFx5_ASAP7_75t_L g184 ( 
.A(n_10),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_13),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_33),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_91),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_53),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_60),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_5),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_63),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_5),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_81),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_119),
.Y(n_194)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_64),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_90),
.Y(n_196)
);

BUFx5_ASAP7_75t_L g197 ( 
.A(n_47),
.Y(n_197)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_19),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_66),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_57),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_118),
.Y(n_201)
);

HB1xp67_ASAP7_75t_L g202 ( 
.A(n_48),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_58),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_49),
.Y(n_204)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_43),
.Y(n_205)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_117),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_39),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_7),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_12),
.Y(n_209)
);

BUFx6f_ASAP7_75t_L g210 ( 
.A(n_27),
.Y(n_210)
);

INVx1_ASAP7_75t_SL g211 ( 
.A(n_99),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_8),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_87),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_98),
.Y(n_214)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_35),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_106),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_43),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_1),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_59),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_86),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_11),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_108),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_120),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_109),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_83),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_32),
.Y(n_226)
);

CKINVDCx14_ASAP7_75t_R g227 ( 
.A(n_20),
.Y(n_227)
);

CKINVDCx16_ASAP7_75t_R g228 ( 
.A(n_46),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_14),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_105),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_23),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_18),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_4),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_14),
.Y(n_234)
);

INVxp67_ASAP7_75t_L g235 ( 
.A(n_88),
.Y(n_235)
);

INVx1_ASAP7_75t_SL g236 ( 
.A(n_127),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_22),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_56),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_93),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_54),
.Y(n_240)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_79),
.Y(n_241)
);

BUFx6f_ASAP7_75t_L g242 ( 
.A(n_50),
.Y(n_242)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_2),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_96),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_38),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_46),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_4),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_153),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_156),
.Y(n_249)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_184),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_184),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_227),
.B(n_167),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_167),
.B(n_0),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_184),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_184),
.Y(n_255)
);

BUFx2_ASAP7_75t_L g256 ( 
.A(n_145),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_184),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_184),
.Y(n_258)
);

INVxp67_ASAP7_75t_SL g259 ( 
.A(n_137),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_184),
.Y(n_260)
);

HB1xp67_ASAP7_75t_L g261 ( 
.A(n_151),
.Y(n_261)
);

CKINVDCx16_ASAP7_75t_R g262 ( 
.A(n_228),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_184),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_165),
.Y(n_264)
);

INVxp67_ASAP7_75t_L g265 ( 
.A(n_202),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_197),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_162),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_170),
.Y(n_268)
);

INVxp33_ASAP7_75t_SL g269 ( 
.A(n_145),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_173),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_188),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_235),
.B(n_2),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_174),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_197),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_197),
.Y(n_275)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_197),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_197),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_197),
.Y(n_278)
);

HB1xp67_ASAP7_75t_L g279 ( 
.A(n_147),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_197),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_197),
.Y(n_281)
);

INVxp67_ASAP7_75t_SL g282 ( 
.A(n_137),
.Y(n_282)
);

INVxp33_ASAP7_75t_SL g283 ( 
.A(n_147),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_175),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_176),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_179),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_210),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_182),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_187),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_210),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_189),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_210),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_210),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_210),
.Y(n_294)
);

CKINVDCx14_ASAP7_75t_R g295 ( 
.A(n_172),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_191),
.Y(n_296)
);

HB1xp67_ASAP7_75t_L g297 ( 
.A(n_149),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_198),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_198),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_193),
.Y(n_300)
);

NOR2xp67_ASAP7_75t_L g301 ( 
.A(n_144),
.B(n_3),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_194),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_196),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_205),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_205),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_199),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_215),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_139),
.B(n_6),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_215),
.Y(n_309)
);

INVx2_ASAP7_75t_L g310 ( 
.A(n_243),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_139),
.B(n_9),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_200),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_201),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_203),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_204),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_243),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_287),
.Y(n_317)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_250),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_R g319 ( 
.A(n_295),
.B(n_131),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_287),
.Y(n_320)
);

NOR2xp67_ASAP7_75t_L g321 ( 
.A(n_251),
.B(n_135),
.Y(n_321)
);

INVx3_ASAP7_75t_L g322 ( 
.A(n_250),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_R g323 ( 
.A(n_273),
.B(n_291),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_249),
.Y(n_324)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_276),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_259),
.B(n_131),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_290),
.Y(n_327)
);

INVx3_ASAP7_75t_L g328 ( 
.A(n_276),
.Y(n_328)
);

AND2x4_ASAP7_75t_L g329 ( 
.A(n_292),
.B(n_157),
.Y(n_329)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_251),
.Y(n_330)
);

AND2x4_ASAP7_75t_L g331 ( 
.A(n_292),
.B(n_157),
.Y(n_331)
);

BUFx6f_ASAP7_75t_L g332 ( 
.A(n_254),
.Y(n_332)
);

INVx2_ASAP7_75t_L g333 ( 
.A(n_254),
.Y(n_333)
);

INVx2_ASAP7_75t_L g334 ( 
.A(n_255),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_293),
.Y(n_335)
);

INVx2_ASAP7_75t_L g336 ( 
.A(n_255),
.Y(n_336)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_257),
.Y(n_337)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_257),
.Y(n_338)
);

BUFx8_ASAP7_75t_L g339 ( 
.A(n_256),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_282),
.B(n_132),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_293),
.Y(n_341)
);

INVx2_ASAP7_75t_L g342 ( 
.A(n_258),
.Y(n_342)
);

BUFx3_ASAP7_75t_L g343 ( 
.A(n_294),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_253),
.B(n_132),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g345 ( 
.A(n_248),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_294),
.Y(n_346)
);

BUFx2_ASAP7_75t_L g347 ( 
.A(n_261),
.Y(n_347)
);

INVx2_ASAP7_75t_L g348 ( 
.A(n_258),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_260),
.B(n_136),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_310),
.Y(n_350)
);

AND2x2_ASAP7_75t_L g351 ( 
.A(n_310),
.B(n_164),
.Y(n_351)
);

BUFx2_ASAP7_75t_L g352 ( 
.A(n_256),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_260),
.B(n_136),
.Y(n_353)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_263),
.Y(n_354)
);

INVx2_ASAP7_75t_L g355 ( 
.A(n_263),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_264),
.Y(n_356)
);

BUFx3_ASAP7_75t_L g357 ( 
.A(n_266),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_268),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_270),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_284),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_285),
.Y(n_361)
);

AND2x2_ASAP7_75t_L g362 ( 
.A(n_266),
.B(n_164),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_274),
.Y(n_363)
);

CKINVDCx6p67_ASAP7_75t_R g364 ( 
.A(n_262),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_274),
.Y(n_365)
);

INVxp67_ASAP7_75t_L g366 ( 
.A(n_279),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_275),
.Y(n_367)
);

BUFx6f_ASAP7_75t_L g368 ( 
.A(n_275),
.Y(n_368)
);

HB1xp67_ASAP7_75t_L g369 ( 
.A(n_297),
.Y(n_369)
);

BUFx6f_ASAP7_75t_L g370 ( 
.A(n_277),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_277),
.Y(n_371)
);

CKINVDCx20_ASAP7_75t_R g372 ( 
.A(n_267),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_278),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_278),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_280),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_R g376 ( 
.A(n_296),
.B(n_138),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_R g377 ( 
.A(n_303),
.B(n_138),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_286),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_280),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_R g380 ( 
.A(n_288),
.B(n_141),
.Y(n_380)
);

OA21x2_ASAP7_75t_L g381 ( 
.A1(n_281),
.A2(n_299),
.B(n_298),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_289),
.Y(n_382)
);

INVx2_ASAP7_75t_L g383 ( 
.A(n_318),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_L g384 ( 
.A(n_344),
.B(n_300),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_SL g385 ( 
.A(n_349),
.B(n_195),
.Y(n_385)
);

INVx2_ASAP7_75t_SL g386 ( 
.A(n_326),
.Y(n_386)
);

AOI22xp33_ASAP7_75t_L g387 ( 
.A1(n_344),
.A2(n_252),
.B1(n_311),
.B2(n_308),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_357),
.Y(n_388)
);

INVx2_ASAP7_75t_SL g389 ( 
.A(n_326),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_363),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_L g391 ( 
.A(n_340),
.B(n_302),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_353),
.B(n_312),
.Y(n_392)
);

INVx3_ASAP7_75t_L g393 ( 
.A(n_322),
.Y(n_393)
);

AOI22xp5_ASAP7_75t_L g394 ( 
.A1(n_366),
.A2(n_306),
.B1(n_315),
.B2(n_314),
.Y(n_394)
);

INVx4_ASAP7_75t_L g395 ( 
.A(n_332),
.Y(n_395)
);

BUFx10_ASAP7_75t_L g396 ( 
.A(n_324),
.Y(n_396)
);

BUFx2_ASAP7_75t_L g397 ( 
.A(n_376),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_363),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_365),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_365),
.Y(n_400)
);

AND2x2_ASAP7_75t_L g401 ( 
.A(n_351),
.B(n_316),
.Y(n_401)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_318),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_367),
.Y(n_403)
);

AND2x4_ASAP7_75t_L g404 ( 
.A(n_351),
.B(n_298),
.Y(n_404)
);

INVx2_ASAP7_75t_L g405 ( 
.A(n_318),
.Y(n_405)
);

AOI22xp33_ASAP7_75t_L g406 ( 
.A1(n_362),
.A2(n_301),
.B1(n_272),
.B2(n_265),
.Y(n_406)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_325),
.Y(n_407)
);

NOR2xp33_ASAP7_75t_L g408 ( 
.A(n_340),
.B(n_313),
.Y(n_408)
);

BUFx6f_ASAP7_75t_L g409 ( 
.A(n_343),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_SL g410 ( 
.A(n_362),
.B(n_206),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_367),
.Y(n_411)
);

AOI22xp33_ASAP7_75t_L g412 ( 
.A1(n_371),
.A2(n_301),
.B1(n_269),
.B2(n_283),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_SL g413 ( 
.A(n_380),
.B(n_241),
.Y(n_413)
);

INVx6_ASAP7_75t_L g414 ( 
.A(n_332),
.Y(n_414)
);

INVx2_ASAP7_75t_L g415 ( 
.A(n_325),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_SL g416 ( 
.A(n_380),
.B(n_133),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_SL g417 ( 
.A(n_377),
.B(n_133),
.Y(n_417)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_325),
.Y(n_418)
);

AND2x2_ASAP7_75t_SL g419 ( 
.A(n_381),
.B(n_133),
.Y(n_419)
);

INVx3_ASAP7_75t_L g420 ( 
.A(n_322),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_373),
.Y(n_421)
);

AND2x4_ASAP7_75t_L g422 ( 
.A(n_351),
.B(n_299),
.Y(n_422)
);

OR2x2_ASAP7_75t_L g423 ( 
.A(n_352),
.B(n_316),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_SL g424 ( 
.A(n_356),
.B(n_133),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_374),
.Y(n_425)
);

AND2x6_ASAP7_75t_L g426 ( 
.A(n_375),
.B(n_133),
.Y(n_426)
);

NOR2xp33_ASAP7_75t_L g427 ( 
.A(n_358),
.B(n_359),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_375),
.B(n_211),
.Y(n_428)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_322),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_379),
.Y(n_430)
);

BUFx3_ASAP7_75t_L g431 ( 
.A(n_381),
.Y(n_431)
);

INVx3_ASAP7_75t_L g432 ( 
.A(n_328),
.Y(n_432)
);

BUFx3_ASAP7_75t_L g433 ( 
.A(n_381),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_343),
.Y(n_434)
);

INVx5_ASAP7_75t_L g435 ( 
.A(n_332),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_343),
.Y(n_436)
);

XNOR2xp5_ASAP7_75t_SL g437 ( 
.A(n_352),
.B(n_9),
.Y(n_437)
);

AND2x2_ASAP7_75t_SL g438 ( 
.A(n_381),
.B(n_242),
.Y(n_438)
);

BUFx3_ASAP7_75t_L g439 ( 
.A(n_381),
.Y(n_439)
);

BUFx10_ASAP7_75t_L g440 ( 
.A(n_360),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_L g441 ( 
.A(n_361),
.B(n_271),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_330),
.B(n_236),
.Y(n_442)
);

OR2x2_ASAP7_75t_L g443 ( 
.A(n_369),
.B(n_309),
.Y(n_443)
);

AND2x2_ASAP7_75t_L g444 ( 
.A(n_350),
.B(n_309),
.Y(n_444)
);

NOR2xp33_ASAP7_75t_L g445 ( 
.A(n_378),
.B(n_141),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_SL g446 ( 
.A(n_382),
.B(n_242),
.Y(n_446)
);

AND2x6_ASAP7_75t_L g447 ( 
.A(n_330),
.B(n_242),
.Y(n_447)
);

AND2x4_ASAP7_75t_L g448 ( 
.A(n_329),
.B(n_331),
.Y(n_448)
);

INVx2_ASAP7_75t_L g449 ( 
.A(n_328),
.Y(n_449)
);

INVx3_ASAP7_75t_L g450 ( 
.A(n_328),
.Y(n_450)
);

INVx2_ASAP7_75t_L g451 ( 
.A(n_328),
.Y(n_451)
);

NAND2x1p5_ASAP7_75t_L g452 ( 
.A(n_329),
.B(n_140),
.Y(n_452)
);

BUFx3_ASAP7_75t_L g453 ( 
.A(n_329),
.Y(n_453)
);

INVx2_ASAP7_75t_SL g454 ( 
.A(n_369),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_323),
.Y(n_455)
);

BUFx4f_ASAP7_75t_L g456 ( 
.A(n_332),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_333),
.Y(n_457)
);

INVx5_ASAP7_75t_L g458 ( 
.A(n_332),
.Y(n_458)
);

AND2x4_ASAP7_75t_L g459 ( 
.A(n_329),
.B(n_331),
.Y(n_459)
);

AOI22xp33_ASAP7_75t_L g460 ( 
.A1(n_331),
.A2(n_181),
.B1(n_134),
.B2(n_183),
.Y(n_460)
);

INVx3_ASAP7_75t_L g461 ( 
.A(n_368),
.Y(n_461)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_334),
.Y(n_462)
);

BUFx6f_ASAP7_75t_L g463 ( 
.A(n_368),
.Y(n_463)
);

INVx3_ASAP7_75t_L g464 ( 
.A(n_368),
.Y(n_464)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_334),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_334),
.Y(n_466)
);

NOR2xp33_ASAP7_75t_L g467 ( 
.A(n_347),
.B(n_142),
.Y(n_467)
);

INVx6_ASAP7_75t_L g468 ( 
.A(n_368),
.Y(n_468)
);

INVx2_ASAP7_75t_L g469 ( 
.A(n_336),
.Y(n_469)
);

NOR2xp33_ASAP7_75t_L g470 ( 
.A(n_347),
.B(n_317),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_336),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_337),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_337),
.Y(n_473)
);

OAI221xp5_ASAP7_75t_L g474 ( 
.A1(n_321),
.A2(n_186),
.B1(n_148),
.B2(n_150),
.C(n_245),
.Y(n_474)
);

AND2x4_ASAP7_75t_L g475 ( 
.A(n_331),
.B(n_304),
.Y(n_475)
);

INVx2_ASAP7_75t_SL g476 ( 
.A(n_319),
.Y(n_476)
);

BUFx6f_ASAP7_75t_L g477 ( 
.A(n_368),
.Y(n_477)
);

AOI22xp33_ASAP7_75t_L g478 ( 
.A1(n_338),
.A2(n_342),
.B1(n_348),
.B2(n_354),
.Y(n_478)
);

INVx3_ASAP7_75t_L g479 ( 
.A(n_368),
.Y(n_479)
);

AND2x2_ASAP7_75t_L g480 ( 
.A(n_350),
.B(n_307),
.Y(n_480)
);

OR2x6_ASAP7_75t_L g481 ( 
.A(n_364),
.B(n_159),
.Y(n_481)
);

INVxp67_ASAP7_75t_L g482 ( 
.A(n_339),
.Y(n_482)
);

OAI22xp33_ASAP7_75t_L g483 ( 
.A1(n_364),
.A2(n_171),
.B1(n_192),
.B2(n_185),
.Y(n_483)
);

AOI22xp33_ASAP7_75t_L g484 ( 
.A1(n_338),
.A2(n_190),
.B1(n_163),
.B2(n_207),
.Y(n_484)
);

BUFx3_ASAP7_75t_L g485 ( 
.A(n_370),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g486 ( 
.A(n_338),
.B(n_146),
.Y(n_486)
);

INVx6_ASAP7_75t_L g487 ( 
.A(n_370),
.Y(n_487)
);

AOI22xp5_ASAP7_75t_L g488 ( 
.A1(n_364),
.A2(n_142),
.B1(n_143),
.B2(n_213),
.Y(n_488)
);

INVx2_ASAP7_75t_L g489 ( 
.A(n_342),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_348),
.Y(n_490)
);

BUFx3_ASAP7_75t_L g491 ( 
.A(n_370),
.Y(n_491)
);

AND2x2_ASAP7_75t_L g492 ( 
.A(n_317),
.B(n_307),
.Y(n_492)
);

BUFx3_ASAP7_75t_L g493 ( 
.A(n_370),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_354),
.Y(n_494)
);

BUFx2_ASAP7_75t_L g495 ( 
.A(n_339),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_SL g496 ( 
.A(n_370),
.B(n_242),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_355),
.Y(n_497)
);

INVx1_ASAP7_75t_SL g498 ( 
.A(n_345),
.Y(n_498)
);

INVx1_ASAP7_75t_SL g499 ( 
.A(n_372),
.Y(n_499)
);

AND2x4_ASAP7_75t_L g500 ( 
.A(n_320),
.B(n_304),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_386),
.B(n_370),
.Y(n_501)
);

AOI22xp33_ASAP7_75t_L g502 ( 
.A1(n_431),
.A2(n_355),
.B1(n_177),
.B2(n_178),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_386),
.B(n_355),
.Y(n_503)
);

INVx2_ASAP7_75t_L g504 ( 
.A(n_431),
.Y(n_504)
);

NOR2xp33_ASAP7_75t_L g505 ( 
.A(n_389),
.B(n_154),
.Y(n_505)
);

INVx2_ASAP7_75t_L g506 ( 
.A(n_433),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_453),
.Y(n_507)
);

OAI22xp5_ASAP7_75t_L g508 ( 
.A1(n_389),
.A2(n_219),
.B1(n_158),
.B2(n_160),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_384),
.B(n_391),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_408),
.B(n_392),
.Y(n_510)
);

INVxp67_ASAP7_75t_SL g511 ( 
.A(n_439),
.Y(n_511)
);

BUFx3_ASAP7_75t_L g512 ( 
.A(n_453),
.Y(n_512)
);

A2O1A1Ixp33_ASAP7_75t_L g513 ( 
.A1(n_387),
.A2(n_223),
.B(n_166),
.C(n_168),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_388),
.B(n_320),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_401),
.Y(n_515)
);

NOR2xp33_ASAP7_75t_SL g516 ( 
.A(n_455),
.B(n_339),
.Y(n_516)
);

NOR2xp33_ASAP7_75t_L g517 ( 
.A(n_423),
.B(n_154),
.Y(n_517)
);

BUFx2_ASAP7_75t_L g518 ( 
.A(n_454),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_390),
.B(n_327),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_398),
.B(n_327),
.Y(n_520)
);

INVxp67_ASAP7_75t_L g521 ( 
.A(n_467),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_399),
.B(n_335),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_L g523 ( 
.A(n_400),
.B(n_335),
.Y(n_523)
);

INVx3_ASAP7_75t_L g524 ( 
.A(n_404),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_403),
.B(n_411),
.Y(n_525)
);

BUFx3_ASAP7_75t_L g526 ( 
.A(n_448),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_404),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_SL g528 ( 
.A(n_419),
.B(n_339),
.Y(n_528)
);

INVx2_ASAP7_75t_L g529 ( 
.A(n_383),
.Y(n_529)
);

AND2x2_ASAP7_75t_L g530 ( 
.A(n_454),
.B(n_172),
.Y(n_530)
);

NOR2xp33_ASAP7_75t_L g531 ( 
.A(n_423),
.B(n_213),
.Y(n_531)
);

INVx2_ASAP7_75t_L g532 ( 
.A(n_383),
.Y(n_532)
);

INVx2_ASAP7_75t_L g533 ( 
.A(n_402),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_SL g534 ( 
.A(n_419),
.B(n_152),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_421),
.B(n_341),
.Y(n_535)
);

NOR2xp33_ASAP7_75t_L g536 ( 
.A(n_470),
.B(n_214),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_425),
.B(n_341),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_SL g538 ( 
.A(n_438),
.B(n_180),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_430),
.B(n_346),
.Y(n_539)
);

NOR2xp67_ASAP7_75t_L g540 ( 
.A(n_476),
.B(n_346),
.Y(n_540)
);

OR2x6_ASAP7_75t_L g541 ( 
.A(n_495),
.B(n_481),
.Y(n_541)
);

NOR2xp33_ASAP7_75t_L g542 ( 
.A(n_445),
.B(n_222),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_SL g543 ( 
.A(n_412),
.B(n_238),
.Y(n_543)
);

INVx4_ASAP7_75t_L g544 ( 
.A(n_409),
.Y(n_544)
);

BUFx6f_ASAP7_75t_L g545 ( 
.A(n_409),
.Y(n_545)
);

NOR2xp33_ASAP7_75t_SL g546 ( 
.A(n_455),
.B(n_218),
.Y(n_546)
);

INVx2_ASAP7_75t_L g547 ( 
.A(n_405),
.Y(n_547)
);

NAND3xp33_ASAP7_75t_L g548 ( 
.A(n_406),
.B(n_155),
.C(n_161),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_422),
.Y(n_549)
);

BUFx6f_ASAP7_75t_L g550 ( 
.A(n_409),
.Y(n_550)
);

AOI22xp33_ASAP7_75t_L g551 ( 
.A1(n_385),
.A2(n_220),
.B1(n_216),
.B2(n_224),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_SL g552 ( 
.A(n_428),
.B(n_238),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_SL g553 ( 
.A(n_438),
.B(n_225),
.Y(n_553)
);

BUFx3_ASAP7_75t_L g554 ( 
.A(n_448),
.Y(n_554)
);

INVx2_ASAP7_75t_L g555 ( 
.A(n_407),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_L g556 ( 
.A(n_434),
.B(n_436),
.Y(n_556)
);

AND2x2_ASAP7_75t_L g557 ( 
.A(n_397),
.B(n_305),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_L g558 ( 
.A(n_459),
.B(n_230),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_L g559 ( 
.A(n_459),
.B(n_239),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_L g560 ( 
.A(n_459),
.B(n_244),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_475),
.Y(n_561)
);

NOR2xp33_ASAP7_75t_L g562 ( 
.A(n_443),
.B(n_240),
.Y(n_562)
);

OR2x6_ASAP7_75t_L g563 ( 
.A(n_481),
.B(n_231),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_SL g564 ( 
.A(n_393),
.B(n_240),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_475),
.Y(n_565)
);

BUFx2_ASAP7_75t_L g566 ( 
.A(n_481),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_407),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_475),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_L g569 ( 
.A(n_442),
.B(n_169),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_500),
.Y(n_570)
);

NOR2xp33_ASAP7_75t_L g571 ( 
.A(n_424),
.B(n_208),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_SL g572 ( 
.A(n_424),
.B(n_247),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_500),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_415),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_SL g575 ( 
.A(n_446),
.B(n_247),
.Y(n_575)
);

AOI22xp33_ASAP7_75t_L g576 ( 
.A1(n_410),
.A2(n_246),
.B1(n_237),
.B2(n_234),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_L g577 ( 
.A(n_420),
.B(n_246),
.Y(n_577)
);

OR2x6_ASAP7_75t_L g578 ( 
.A(n_481),
.B(n_13),
.Y(n_578)
);

NOR2xp33_ASAP7_75t_L g579 ( 
.A(n_446),
.B(n_234),
.Y(n_579)
);

INVx2_ASAP7_75t_L g580 ( 
.A(n_415),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_SL g581 ( 
.A(n_432),
.B(n_233),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_L g582 ( 
.A(n_432),
.B(n_232),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_500),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_SL g584 ( 
.A(n_450),
.B(n_229),
.Y(n_584)
);

NOR3xp33_ASAP7_75t_L g585 ( 
.A(n_483),
.B(n_217),
.C(n_221),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_L g586 ( 
.A(n_450),
.B(n_226),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_SL g587 ( 
.A(n_394),
.B(n_226),
.Y(n_587)
);

NOR2xp33_ASAP7_75t_L g588 ( 
.A(n_413),
.B(n_212),
.Y(n_588)
);

INVx2_ASAP7_75t_SL g589 ( 
.A(n_417),
.Y(n_589)
);

INVx2_ASAP7_75t_SL g590 ( 
.A(n_417),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_492),
.Y(n_591)
);

INVx2_ASAP7_75t_L g592 ( 
.A(n_418),
.Y(n_592)
);

INVx2_ASAP7_75t_SL g593 ( 
.A(n_416),
.Y(n_593)
);

INVx2_ASAP7_75t_L g594 ( 
.A(n_418),
.Y(n_594)
);

BUFx6f_ASAP7_75t_L g595 ( 
.A(n_485),
.Y(n_595)
);

NOR3x1_ASAP7_75t_L g596 ( 
.A(n_474),
.B(n_209),
.C(n_17),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_L g597 ( 
.A(n_461),
.B(n_128),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_492),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_SL g599 ( 
.A(n_462),
.B(n_123),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_SL g600 ( 
.A(n_462),
.B(n_121),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_L g601 ( 
.A(n_464),
.B(n_116),
.Y(n_601)
);

BUFx3_ASAP7_75t_L g602 ( 
.A(n_396),
.Y(n_602)
);

BUFx3_ASAP7_75t_L g603 ( 
.A(n_396),
.Y(n_603)
);

INVx2_ASAP7_75t_L g604 ( 
.A(n_465),
.Y(n_604)
);

INVx2_ASAP7_75t_L g605 ( 
.A(n_465),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g606 ( 
.A(n_464),
.B(n_114),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_444),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_480),
.Y(n_608)
);

AOI22xp5_ASAP7_75t_L g609 ( 
.A1(n_416),
.A2(n_110),
.B1(n_104),
.B2(n_101),
.Y(n_609)
);

OAI22xp5_ASAP7_75t_L g610 ( 
.A1(n_488),
.A2(n_80),
.B1(n_78),
.B2(n_74),
.Y(n_610)
);

AND2x4_ASAP7_75t_L g611 ( 
.A(n_480),
.B(n_73),
.Y(n_611)
);

NOR2xp33_ASAP7_75t_L g612 ( 
.A(n_427),
.B(n_16),
.Y(n_612)
);

NOR2x1p5_ASAP7_75t_L g613 ( 
.A(n_437),
.B(n_16),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_SL g614 ( 
.A(n_469),
.B(n_489),
.Y(n_614)
);

INVx2_ASAP7_75t_SL g615 ( 
.A(n_396),
.Y(n_615)
);

AND2x2_ASAP7_75t_L g616 ( 
.A(n_440),
.B(n_17),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_429),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_SL g618 ( 
.A(n_469),
.B(n_71),
.Y(n_618)
);

INVx2_ASAP7_75t_L g619 ( 
.A(n_489),
.Y(n_619)
);

NOR2xp67_ASAP7_75t_L g620 ( 
.A(n_482),
.B(n_18),
.Y(n_620)
);

OAI22xp5_ASAP7_75t_L g621 ( 
.A1(n_452),
.A2(n_22),
.B1(n_24),
.B2(n_25),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_429),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_SL g623 ( 
.A(n_479),
.B(n_27),
.Y(n_623)
);

NOR2xp33_ASAP7_75t_L g624 ( 
.A(n_457),
.B(n_28),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_509),
.B(n_466),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_L g626 ( 
.A(n_510),
.B(n_503),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_527),
.Y(n_627)
);

BUFx2_ASAP7_75t_L g628 ( 
.A(n_518),
.Y(n_628)
);

OAI21xp5_ASAP7_75t_L g629 ( 
.A1(n_504),
.A2(n_478),
.B(n_497),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_L g630 ( 
.A(n_511),
.B(n_473),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_L g631 ( 
.A(n_504),
.B(n_472),
.Y(n_631)
);

AOI21xp5_ASAP7_75t_L g632 ( 
.A1(n_544),
.A2(n_395),
.B(n_491),
.Y(n_632)
);

AOI21x1_ASAP7_75t_L g633 ( 
.A1(n_614),
.A2(n_471),
.B(n_494),
.Y(n_633)
);

AOI21xp5_ASAP7_75t_L g634 ( 
.A1(n_534),
.A2(n_493),
.B(n_491),
.Y(n_634)
);

AOI21xp5_ASAP7_75t_L g635 ( 
.A1(n_538),
.A2(n_493),
.B(n_477),
.Y(n_635)
);

AOI21xp5_ASAP7_75t_L g636 ( 
.A1(n_538),
.A2(n_477),
.B(n_463),
.Y(n_636)
);

AND2x4_ASAP7_75t_L g637 ( 
.A(n_526),
.B(n_499),
.Y(n_637)
);

AOI21xp5_ASAP7_75t_L g638 ( 
.A1(n_553),
.A2(n_463),
.B(n_477),
.Y(n_638)
);

OAI22xp5_ASAP7_75t_L g639 ( 
.A1(n_506),
.A2(n_460),
.B1(n_484),
.B2(n_441),
.Y(n_639)
);

OAI21xp5_ASAP7_75t_L g640 ( 
.A1(n_506),
.A2(n_490),
.B(n_486),
.Y(n_640)
);

INVx2_ASAP7_75t_L g641 ( 
.A(n_529),
.Y(n_641)
);

NOR3xp33_ASAP7_75t_L g642 ( 
.A(n_521),
.B(n_498),
.C(n_496),
.Y(n_642)
);

AOI21xp5_ASAP7_75t_L g643 ( 
.A1(n_553),
.A2(n_477),
.B(n_463),
.Y(n_643)
);

O2A1O1Ixp33_ASAP7_75t_L g644 ( 
.A1(n_513),
.A2(n_623),
.B(n_612),
.C(n_584),
.Y(n_644)
);

AOI21xp5_ASAP7_75t_L g645 ( 
.A1(n_556),
.A2(n_463),
.B(n_435),
.Y(n_645)
);

A2O1A1Ixp33_ASAP7_75t_L g646 ( 
.A1(n_579),
.A2(n_479),
.B(n_449),
.C(n_451),
.Y(n_646)
);

AOI21xp5_ASAP7_75t_L g647 ( 
.A1(n_558),
.A2(n_435),
.B(n_458),
.Y(n_647)
);

NOR2xp33_ASAP7_75t_L g648 ( 
.A(n_542),
.B(n_440),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_542),
.B(n_451),
.Y(n_649)
);

OAI21xp5_ASAP7_75t_L g650 ( 
.A1(n_502),
.A2(n_426),
.B(n_447),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_L g651 ( 
.A(n_505),
.B(n_524),
.Y(n_651)
);

INVx3_ASAP7_75t_SL g652 ( 
.A(n_615),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_L g653 ( 
.A(n_505),
.B(n_487),
.Y(n_653)
);

AOI21xp5_ASAP7_75t_L g654 ( 
.A1(n_559),
.A2(n_435),
.B(n_458),
.Y(n_654)
);

OAI21xp5_ASAP7_75t_L g655 ( 
.A1(n_614),
.A2(n_426),
.B(n_447),
.Y(n_655)
);

INVxp67_ASAP7_75t_L g656 ( 
.A(n_557),
.Y(n_656)
);

INVx1_ASAP7_75t_SL g657 ( 
.A(n_530),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_549),
.Y(n_658)
);

AOI21xp5_ASAP7_75t_L g659 ( 
.A1(n_560),
.A2(n_435),
.B(n_458),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_593),
.B(n_487),
.Y(n_660)
);

NAND3xp33_ASAP7_75t_SL g661 ( 
.A(n_612),
.B(n_437),
.C(n_440),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_L g662 ( 
.A(n_589),
.B(n_468),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_L g663 ( 
.A(n_590),
.B(n_468),
.Y(n_663)
);

BUFx4f_ASAP7_75t_L g664 ( 
.A(n_541),
.Y(n_664)
);

AOI22xp33_ASAP7_75t_L g665 ( 
.A1(n_611),
.A2(n_468),
.B1(n_414),
.B2(n_426),
.Y(n_665)
);

A2O1A1Ixp33_ASAP7_75t_L g666 ( 
.A1(n_588),
.A2(n_458),
.B(n_435),
.C(n_468),
.Y(n_666)
);

NOR3xp33_ASAP7_75t_L g667 ( 
.A(n_587),
.B(n_28),
.C(n_29),
.Y(n_667)
);

AOI21xp5_ASAP7_75t_L g668 ( 
.A1(n_525),
.A2(n_458),
.B(n_414),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_591),
.B(n_414),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_L g670 ( 
.A(n_598),
.B(n_426),
.Y(n_670)
);

AND2x4_ASAP7_75t_L g671 ( 
.A(n_526),
.B(n_30),
.Y(n_671)
);

AOI21xp5_ASAP7_75t_L g672 ( 
.A1(n_545),
.A2(n_447),
.B(n_426),
.Y(n_672)
);

OAI21xp5_ASAP7_75t_L g673 ( 
.A1(n_515),
.A2(n_447),
.B(n_31),
.Y(n_673)
);

AOI21xp5_ASAP7_75t_L g674 ( 
.A1(n_545),
.A2(n_447),
.B(n_31),
.Y(n_674)
);

NOR2xp67_ASAP7_75t_L g675 ( 
.A(n_602),
.B(n_30),
.Y(n_675)
);

AOI21xp5_ASAP7_75t_L g676 ( 
.A1(n_545),
.A2(n_32),
.B(n_33),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_607),
.B(n_34),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_L g678 ( 
.A(n_608),
.B(n_34),
.Y(n_678)
);

AOI21xp5_ASAP7_75t_L g679 ( 
.A1(n_550),
.A2(n_35),
.B(n_36),
.Y(n_679)
);

A2O1A1Ixp33_ASAP7_75t_L g680 ( 
.A1(n_588),
.A2(n_48),
.B(n_41),
.C(n_42),
.Y(n_680)
);

O2A1O1Ixp33_ASAP7_75t_L g681 ( 
.A1(n_623),
.A2(n_37),
.B(n_42),
.C(n_45),
.Y(n_681)
);

AOI21xp5_ASAP7_75t_L g682 ( 
.A1(n_550),
.A2(n_37),
.B(n_45),
.Y(n_682)
);

NOR2xp33_ASAP7_75t_L g683 ( 
.A(n_546),
.B(n_517),
.Y(n_683)
);

INVx4_ASAP7_75t_L g684 ( 
.A(n_554),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_570),
.Y(n_685)
);

OR2x2_ASAP7_75t_L g686 ( 
.A(n_517),
.B(n_531),
.Y(n_686)
);

AOI21xp5_ASAP7_75t_L g687 ( 
.A1(n_514),
.A2(n_611),
.B(n_561),
.Y(n_687)
);

AOI21xp5_ASAP7_75t_L g688 ( 
.A1(n_565),
.A2(n_568),
.B(n_573),
.Y(n_688)
);

OAI22xp5_ASAP7_75t_L g689 ( 
.A1(n_571),
.A2(n_551),
.B1(n_528),
.B2(n_583),
.Y(n_689)
);

OAI21xp5_ASAP7_75t_L g690 ( 
.A1(n_604),
.A2(n_619),
.B(n_605),
.Y(n_690)
);

BUFx3_ASAP7_75t_L g691 ( 
.A(n_602),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_L g692 ( 
.A(n_562),
.B(n_569),
.Y(n_692)
);

NOR3xp33_ASAP7_75t_L g693 ( 
.A(n_543),
.B(n_531),
.C(n_548),
.Y(n_693)
);

OAI21xp5_ASAP7_75t_L g694 ( 
.A1(n_604),
.A2(n_605),
.B(n_619),
.Y(n_694)
);

O2A1O1Ixp33_ASAP7_75t_L g695 ( 
.A1(n_581),
.A2(n_584),
.B(n_508),
.C(n_564),
.Y(n_695)
);

INVxp67_ASAP7_75t_L g696 ( 
.A(n_562),
.Y(n_696)
);

BUFx4f_ASAP7_75t_L g697 ( 
.A(n_541),
.Y(n_697)
);

AOI21x1_ASAP7_75t_L g698 ( 
.A1(n_519),
.A2(n_537),
.B(n_539),
.Y(n_698)
);

AND2x4_ASAP7_75t_L g699 ( 
.A(n_554),
.B(n_512),
.Y(n_699)
);

BUFx6f_ASAP7_75t_L g700 ( 
.A(n_512),
.Y(n_700)
);

INVx3_ASAP7_75t_L g701 ( 
.A(n_595),
.Y(n_701)
);

CKINVDCx8_ASAP7_75t_R g702 ( 
.A(n_566),
.Y(n_702)
);

INVx1_ASAP7_75t_SL g703 ( 
.A(n_603),
.Y(n_703)
);

AOI21xp5_ASAP7_75t_L g704 ( 
.A1(n_520),
.A2(n_522),
.B(n_523),
.Y(n_704)
);

OAI21xp5_ASAP7_75t_L g705 ( 
.A1(n_532),
.A2(n_580),
.B(n_574),
.Y(n_705)
);

AOI21xp5_ASAP7_75t_L g706 ( 
.A1(n_535),
.A2(n_606),
.B(n_601),
.Y(n_706)
);

AND2x4_ASAP7_75t_L g707 ( 
.A(n_507),
.B(n_603),
.Y(n_707)
);

INVx3_ASAP7_75t_L g708 ( 
.A(n_595),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_571),
.B(n_540),
.Y(n_709)
);

NOR2xp33_ASAP7_75t_L g710 ( 
.A(n_552),
.B(n_575),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_L g711 ( 
.A(n_577),
.B(n_582),
.Y(n_711)
);

NAND2x1p5_ASAP7_75t_L g712 ( 
.A(n_595),
.B(n_528),
.Y(n_712)
);

BUFx6f_ASAP7_75t_L g713 ( 
.A(n_595),
.Y(n_713)
);

NOR2xp33_ASAP7_75t_L g714 ( 
.A(n_572),
.B(n_581),
.Y(n_714)
);

AOI21xp5_ASAP7_75t_L g715 ( 
.A1(n_597),
.A2(n_617),
.B(n_622),
.Y(n_715)
);

AOI21xp5_ASAP7_75t_L g716 ( 
.A1(n_586),
.A2(n_580),
.B(n_532),
.Y(n_716)
);

BUFx2_ASAP7_75t_L g717 ( 
.A(n_578),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_L g718 ( 
.A(n_533),
.B(n_574),
.Y(n_718)
);

INVx5_ASAP7_75t_L g719 ( 
.A(n_533),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_547),
.B(n_592),
.Y(n_720)
);

INVx1_ASAP7_75t_SL g721 ( 
.A(n_616),
.Y(n_721)
);

AO21x1_ASAP7_75t_L g722 ( 
.A1(n_621),
.A2(n_618),
.B(n_600),
.Y(n_722)
);

HB1xp67_ASAP7_75t_L g723 ( 
.A(n_596),
.Y(n_723)
);

NOR2xp33_ASAP7_75t_L g724 ( 
.A(n_563),
.B(n_541),
.Y(n_724)
);

INVx2_ASAP7_75t_SL g725 ( 
.A(n_613),
.Y(n_725)
);

AOI21xp5_ASAP7_75t_L g726 ( 
.A1(n_555),
.A2(n_594),
.B(n_567),
.Y(n_726)
);

BUFx10_ASAP7_75t_L g727 ( 
.A(n_624),
.Y(n_727)
);

NOR2xp33_ASAP7_75t_L g728 ( 
.A(n_563),
.B(n_585),
.Y(n_728)
);

HB1xp67_ASAP7_75t_L g729 ( 
.A(n_620),
.Y(n_729)
);

INVx2_ASAP7_75t_L g730 ( 
.A(n_599),
.Y(n_730)
);

INVx2_ASAP7_75t_L g731 ( 
.A(n_600),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_610),
.Y(n_732)
);

A2O1A1Ixp33_ASAP7_75t_L g733 ( 
.A1(n_609),
.A2(n_509),
.B(n_510),
.C(n_579),
.Y(n_733)
);

HB1xp67_ASAP7_75t_L g734 ( 
.A(n_578),
.Y(n_734)
);

BUFx6f_ASAP7_75t_L g735 ( 
.A(n_578),
.Y(n_735)
);

AOI21xp5_ASAP7_75t_L g736 ( 
.A1(n_576),
.A2(n_456),
.B(n_501),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_SL g737 ( 
.A(n_509),
.B(n_510),
.Y(n_737)
);

BUFx6f_ASAP7_75t_L g738 ( 
.A(n_526),
.Y(n_738)
);

NOR2xp33_ASAP7_75t_L g739 ( 
.A(n_509),
.B(n_510),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_L g740 ( 
.A(n_509),
.B(n_510),
.Y(n_740)
);

CKINVDCx6p67_ASAP7_75t_R g741 ( 
.A(n_602),
.Y(n_741)
);

AOI21xp5_ASAP7_75t_L g742 ( 
.A1(n_501),
.A2(n_456),
.B(n_433),
.Y(n_742)
);

INVx2_ASAP7_75t_L g743 ( 
.A(n_529),
.Y(n_743)
);

AOI21xp5_ASAP7_75t_L g744 ( 
.A1(n_501),
.A2(n_456),
.B(n_433),
.Y(n_744)
);

BUFx6f_ASAP7_75t_L g745 ( 
.A(n_526),
.Y(n_745)
);

BUFx12f_ASAP7_75t_L g746 ( 
.A(n_615),
.Y(n_746)
);

A2O1A1Ixp33_ASAP7_75t_L g747 ( 
.A1(n_509),
.A2(n_510),
.B(n_579),
.C(n_588),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_SL g748 ( 
.A(n_509),
.B(n_510),
.Y(n_748)
);

AOI21xp5_ASAP7_75t_L g749 ( 
.A1(n_501),
.A2(n_456),
.B(n_433),
.Y(n_749)
);

AOI21xp5_ASAP7_75t_L g750 ( 
.A1(n_501),
.A2(n_456),
.B(n_433),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_L g751 ( 
.A(n_509),
.B(n_510),
.Y(n_751)
);

BUFx2_ASAP7_75t_L g752 ( 
.A(n_518),
.Y(n_752)
);

AOI21xp5_ASAP7_75t_L g753 ( 
.A1(n_501),
.A2(n_456),
.B(n_433),
.Y(n_753)
);

AOI21xp5_ASAP7_75t_L g754 ( 
.A1(n_501),
.A2(n_456),
.B(n_433),
.Y(n_754)
);

NAND3xp33_ASAP7_75t_L g755 ( 
.A(n_509),
.B(n_536),
.C(n_542),
.Y(n_755)
);

AND2x2_ASAP7_75t_L g756 ( 
.A(n_518),
.B(n_557),
.Y(n_756)
);

CKINVDCx5p33_ASAP7_75t_R g757 ( 
.A(n_602),
.Y(n_757)
);

NOR2xp33_ASAP7_75t_L g758 ( 
.A(n_509),
.B(n_510),
.Y(n_758)
);

O2A1O1Ixp33_ASAP7_75t_L g759 ( 
.A1(n_509),
.A2(n_538),
.B(n_553),
.C(n_534),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_509),
.B(n_510),
.Y(n_760)
);

OAI321xp33_ASAP7_75t_L g761 ( 
.A1(n_509),
.A2(n_612),
.A3(n_536),
.B1(n_621),
.B2(n_513),
.C(n_588),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_SL g762 ( 
.A(n_509),
.B(n_510),
.Y(n_762)
);

NOR2xp33_ASAP7_75t_SL g763 ( 
.A(n_516),
.B(n_455),
.Y(n_763)
);

NOR2xp33_ASAP7_75t_L g764 ( 
.A(n_509),
.B(n_510),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_L g765 ( 
.A(n_739),
.B(n_758),
.Y(n_765)
);

AOI22xp5_ASAP7_75t_L g766 ( 
.A1(n_764),
.A2(n_751),
.B1(n_740),
.B2(n_760),
.Y(n_766)
);

OAI21x1_ASAP7_75t_L g767 ( 
.A1(n_633),
.A2(n_716),
.B(n_715),
.Y(n_767)
);

BUFx2_ASAP7_75t_L g768 ( 
.A(n_628),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_627),
.Y(n_769)
);

OAI21xp33_ASAP7_75t_L g770 ( 
.A1(n_686),
.A2(n_683),
.B(n_755),
.Y(n_770)
);

BUFx6f_ASAP7_75t_L g771 ( 
.A(n_713),
.Y(n_771)
);

OR2x2_ASAP7_75t_L g772 ( 
.A(n_656),
.B(n_756),
.Y(n_772)
);

OAI21x1_ASAP7_75t_L g773 ( 
.A1(n_690),
.A2(n_705),
.B(n_694),
.Y(n_773)
);

INVx5_ASAP7_75t_L g774 ( 
.A(n_713),
.Y(n_774)
);

OAI21xp33_ASAP7_75t_L g775 ( 
.A1(n_747),
.A2(n_648),
.B(n_696),
.Y(n_775)
);

AOI21xp5_ASAP7_75t_L g776 ( 
.A1(n_706),
.A2(n_687),
.B(n_704),
.Y(n_776)
);

INVx3_ASAP7_75t_L g777 ( 
.A(n_713),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_L g778 ( 
.A(n_626),
.B(n_737),
.Y(n_778)
);

AO21x1_ASAP7_75t_L g779 ( 
.A1(n_644),
.A2(n_689),
.B(n_759),
.Y(n_779)
);

OR2x6_ASAP7_75t_L g780 ( 
.A(n_752),
.B(n_735),
.Y(n_780)
);

NOR2x1_ASAP7_75t_L g781 ( 
.A(n_691),
.B(n_684),
.Y(n_781)
);

AOI21xp5_ASAP7_75t_L g782 ( 
.A1(n_748),
.A2(n_762),
.B(n_709),
.Y(n_782)
);

AO31x2_ASAP7_75t_L g783 ( 
.A1(n_666),
.A2(n_646),
.A3(n_689),
.B(n_733),
.Y(n_783)
);

A2O1A1Ixp33_ASAP7_75t_L g784 ( 
.A1(n_695),
.A2(n_692),
.B(n_714),
.C(n_761),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_625),
.B(n_711),
.Y(n_785)
);

INVx1_ASAP7_75t_SL g786 ( 
.A(n_657),
.Y(n_786)
);

OAI21x1_ASAP7_75t_L g787 ( 
.A1(n_726),
.A2(n_750),
.B(n_744),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_658),
.Y(n_788)
);

AO21x1_ASAP7_75t_L g789 ( 
.A1(n_732),
.A2(n_693),
.B(n_736),
.Y(n_789)
);

INVx5_ASAP7_75t_L g790 ( 
.A(n_746),
.Y(n_790)
);

OAI21x1_ASAP7_75t_L g791 ( 
.A1(n_742),
.A2(n_754),
.B(n_753),
.Y(n_791)
);

AND2x4_ASAP7_75t_L g792 ( 
.A(n_699),
.B(n_707),
.Y(n_792)
);

BUFx4f_ASAP7_75t_L g793 ( 
.A(n_741),
.Y(n_793)
);

OAI21x1_ASAP7_75t_L g794 ( 
.A1(n_749),
.A2(n_638),
.B(n_636),
.Y(n_794)
);

OAI21x1_ASAP7_75t_L g795 ( 
.A1(n_643),
.A2(n_635),
.B(n_632),
.Y(n_795)
);

BUFx3_ASAP7_75t_L g796 ( 
.A(n_652),
.Y(n_796)
);

AOI21xp33_ASAP7_75t_L g797 ( 
.A1(n_710),
.A2(n_681),
.B(n_651),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_685),
.Y(n_798)
);

AO31x2_ASAP7_75t_L g799 ( 
.A1(n_649),
.A2(n_680),
.A3(n_731),
.B(n_730),
.Y(n_799)
);

AOI21xp5_ASAP7_75t_L g800 ( 
.A1(n_625),
.A2(n_630),
.B(n_653),
.Y(n_800)
);

AOI221xp5_ASAP7_75t_L g801 ( 
.A1(n_667),
.A2(n_661),
.B1(n_728),
.B2(n_639),
.C(n_723),
.Y(n_801)
);

OAI21x1_ASAP7_75t_L g802 ( 
.A1(n_634),
.A2(n_640),
.B(n_631),
.Y(n_802)
);

INVx2_ASAP7_75t_SL g803 ( 
.A(n_725),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_L g804 ( 
.A(n_631),
.B(n_641),
.Y(n_804)
);

OAI22xp5_ASAP7_75t_L g805 ( 
.A1(n_639),
.A2(n_678),
.B1(n_677),
.B2(n_665),
.Y(n_805)
);

AND2x4_ASAP7_75t_L g806 ( 
.A(n_699),
.B(n_707),
.Y(n_806)
);

OAI21x1_ASAP7_75t_SL g807 ( 
.A1(n_688),
.A2(n_673),
.B(n_682),
.Y(n_807)
);

OAI21x1_ASAP7_75t_L g808 ( 
.A1(n_640),
.A2(n_659),
.B(n_654),
.Y(n_808)
);

INVx4_ASAP7_75t_L g809 ( 
.A(n_700),
.Y(n_809)
);

OAI21x1_ASAP7_75t_L g810 ( 
.A1(n_647),
.A2(n_720),
.B(n_718),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_L g811 ( 
.A(n_743),
.B(n_698),
.Y(n_811)
);

OAI21x1_ASAP7_75t_L g812 ( 
.A1(n_629),
.A2(n_645),
.B(n_668),
.Y(n_812)
);

OAI21x1_ASAP7_75t_L g813 ( 
.A1(n_669),
.A2(n_662),
.B(n_663),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_L g814 ( 
.A(n_721),
.B(n_708),
.Y(n_814)
);

INVx3_ASAP7_75t_L g815 ( 
.A(n_701),
.Y(n_815)
);

INVx4_ASAP7_75t_L g816 ( 
.A(n_700),
.Y(n_816)
);

OAI21x1_ASAP7_75t_L g817 ( 
.A1(n_660),
.A2(n_701),
.B(n_708),
.Y(n_817)
);

OAI21x1_ASAP7_75t_L g818 ( 
.A1(n_712),
.A2(n_670),
.B(n_672),
.Y(n_818)
);

OR2x2_ASAP7_75t_L g819 ( 
.A(n_637),
.B(n_703),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_L g820 ( 
.A(n_738),
.B(n_745),
.Y(n_820)
);

OAI21x1_ASAP7_75t_L g821 ( 
.A1(n_712),
.A2(n_655),
.B(n_650),
.Y(n_821)
);

OAI21x1_ASAP7_75t_L g822 ( 
.A1(n_655),
.A2(n_674),
.B(n_679),
.Y(n_822)
);

AOI21xp5_ASAP7_75t_L g823 ( 
.A1(n_719),
.A2(n_684),
.B(n_738),
.Y(n_823)
);

OAI21x1_ASAP7_75t_L g824 ( 
.A1(n_676),
.A2(n_675),
.B(n_729),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_L g825 ( 
.A(n_738),
.B(n_745),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_671),
.Y(n_826)
);

AOI21xp5_ASAP7_75t_L g827 ( 
.A1(n_745),
.A2(n_700),
.B(n_637),
.Y(n_827)
);

NOR2xp33_ASAP7_75t_L g828 ( 
.A(n_727),
.B(n_763),
.Y(n_828)
);

AO31x2_ASAP7_75t_L g829 ( 
.A1(n_724),
.A2(n_717),
.A3(n_727),
.B(n_671),
.Y(n_829)
);

AND2x2_ASAP7_75t_L g830 ( 
.A(n_642),
.B(n_757),
.Y(n_830)
);

OAI21x1_ASAP7_75t_L g831 ( 
.A1(n_734),
.A2(n_664),
.B(n_697),
.Y(n_831)
);

AND2x2_ASAP7_75t_L g832 ( 
.A(n_735),
.B(n_702),
.Y(n_832)
);

INVxp67_ASAP7_75t_L g833 ( 
.A(n_735),
.Y(n_833)
);

INVx6_ASAP7_75t_L g834 ( 
.A(n_697),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_627),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_L g836 ( 
.A(n_739),
.B(n_758),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_SL g837 ( 
.A(n_686),
.B(n_509),
.Y(n_837)
);

AND2x2_ASAP7_75t_L g838 ( 
.A(n_756),
.B(n_656),
.Y(n_838)
);

AND2x2_ASAP7_75t_L g839 ( 
.A(n_756),
.B(n_656),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_L g840 ( 
.A(n_739),
.B(n_758),
.Y(n_840)
);

BUFx3_ASAP7_75t_L g841 ( 
.A(n_628),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_739),
.B(n_758),
.Y(n_842)
);

INVxp67_ASAP7_75t_L g843 ( 
.A(n_628),
.Y(n_843)
);

AOI22xp5_ASAP7_75t_L g844 ( 
.A1(n_739),
.A2(n_758),
.B1(n_764),
.B2(n_509),
.Y(n_844)
);

AO21x1_ASAP7_75t_L g845 ( 
.A1(n_644),
.A2(n_509),
.B(n_689),
.Y(n_845)
);

NAND2x1p5_ASAP7_75t_L g846 ( 
.A(n_713),
.B(n_684),
.Y(n_846)
);

NOR2xp67_ASAP7_75t_SL g847 ( 
.A(n_755),
.B(n_602),
.Y(n_847)
);

AOI21x1_ASAP7_75t_SL g848 ( 
.A1(n_692),
.A2(n_509),
.B(n_709),
.Y(n_848)
);

BUFx3_ASAP7_75t_L g849 ( 
.A(n_628),
.Y(n_849)
);

AOI22xp5_ASAP7_75t_L g850 ( 
.A1(n_739),
.A2(n_758),
.B1(n_764),
.B2(n_509),
.Y(n_850)
);

A2O1A1Ixp33_ASAP7_75t_L g851 ( 
.A1(n_739),
.A2(n_764),
.B(n_758),
.C(n_509),
.Y(n_851)
);

OAI21xp5_ASAP7_75t_L g852 ( 
.A1(n_747),
.A2(n_733),
.B(n_739),
.Y(n_852)
);

A2O1A1Ixp33_ASAP7_75t_L g853 ( 
.A1(n_739),
.A2(n_764),
.B(n_758),
.C(n_509),
.Y(n_853)
);

INVx4_ASAP7_75t_L g854 ( 
.A(n_713),
.Y(n_854)
);

OAI22x1_ASAP7_75t_L g855 ( 
.A1(n_683),
.A2(n_755),
.B1(n_648),
.B2(n_509),
.Y(n_855)
);

OAI22xp5_ASAP7_75t_L g856 ( 
.A1(n_739),
.A2(n_764),
.B1(n_758),
.B2(n_509),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_739),
.B(n_758),
.Y(n_857)
);

OR2x2_ASAP7_75t_L g858 ( 
.A(n_740),
.B(n_751),
.Y(n_858)
);

OAI21x1_ASAP7_75t_L g859 ( 
.A1(n_633),
.A2(n_716),
.B(n_715),
.Y(n_859)
);

OAI21x1_ASAP7_75t_L g860 ( 
.A1(n_633),
.A2(n_716),
.B(n_715),
.Y(n_860)
);

BUFx2_ASAP7_75t_L g861 ( 
.A(n_628),
.Y(n_861)
);

INVx3_ASAP7_75t_L g862 ( 
.A(n_713),
.Y(n_862)
);

OAI22xp5_ASAP7_75t_L g863 ( 
.A1(n_739),
.A2(n_764),
.B1(n_758),
.B2(n_509),
.Y(n_863)
);

INVx5_ASAP7_75t_L g864 ( 
.A(n_713),
.Y(n_864)
);

NAND2x1p5_ASAP7_75t_L g865 ( 
.A(n_713),
.B(n_684),
.Y(n_865)
);

INVx5_ASAP7_75t_L g866 ( 
.A(n_713),
.Y(n_866)
);

AO31x2_ASAP7_75t_L g867 ( 
.A1(n_722),
.A2(n_666),
.A3(n_646),
.B(n_689),
.Y(n_867)
);

AND2x4_ASAP7_75t_L g868 ( 
.A(n_699),
.B(n_707),
.Y(n_868)
);

AO31x2_ASAP7_75t_L g869 ( 
.A1(n_722),
.A2(n_666),
.A3(n_646),
.B(n_689),
.Y(n_869)
);

OAI21xp5_ASAP7_75t_L g870 ( 
.A1(n_747),
.A2(n_733),
.B(n_739),
.Y(n_870)
);

AOI21xp33_ASAP7_75t_L g871 ( 
.A1(n_686),
.A2(n_509),
.B(n_755),
.Y(n_871)
);

INVx3_ASAP7_75t_L g872 ( 
.A(n_713),
.Y(n_872)
);

INVx3_ASAP7_75t_SL g873 ( 
.A(n_757),
.Y(n_873)
);

AOI21xp5_ASAP7_75t_L g874 ( 
.A1(n_759),
.A2(n_751),
.B(n_740),
.Y(n_874)
);

OAI21x1_ASAP7_75t_L g875 ( 
.A1(n_633),
.A2(n_716),
.B(n_715),
.Y(n_875)
);

INVx4_ASAP7_75t_L g876 ( 
.A(n_713),
.Y(n_876)
);

INVx3_ASAP7_75t_L g877 ( 
.A(n_713),
.Y(n_877)
);

AO21x1_ASAP7_75t_L g878 ( 
.A1(n_644),
.A2(n_509),
.B(n_689),
.Y(n_878)
);

OR2x6_ASAP7_75t_L g879 ( 
.A(n_628),
.B(n_752),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_L g880 ( 
.A(n_739),
.B(n_758),
.Y(n_880)
);

INVx1_ASAP7_75t_SL g881 ( 
.A(n_756),
.Y(n_881)
);

INVx1_ASAP7_75t_SL g882 ( 
.A(n_756),
.Y(n_882)
);

NOR2xp67_ASAP7_75t_L g883 ( 
.A(n_729),
.B(n_615),
.Y(n_883)
);

O2A1O1Ixp33_ASAP7_75t_L g884 ( 
.A1(n_851),
.A2(n_853),
.B(n_856),
.C(n_863),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_L g885 ( 
.A(n_765),
.B(n_836),
.Y(n_885)
);

NAND2x1p5_ASAP7_75t_L g886 ( 
.A(n_774),
.B(n_864),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_L g887 ( 
.A(n_765),
.B(n_840),
.Y(n_887)
);

AOI21xp5_ASAP7_75t_L g888 ( 
.A1(n_776),
.A2(n_870),
.B(n_852),
.Y(n_888)
);

BUFx3_ASAP7_75t_L g889 ( 
.A(n_796),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_L g890 ( 
.A(n_840),
.B(n_842),
.Y(n_890)
);

OR2x6_ASAP7_75t_L g891 ( 
.A(n_834),
.B(n_879),
.Y(n_891)
);

OR2x2_ASAP7_75t_L g892 ( 
.A(n_858),
.B(n_881),
.Y(n_892)
);

NAND2x1p5_ASAP7_75t_L g893 ( 
.A(n_774),
.B(n_864),
.Y(n_893)
);

BUFx3_ASAP7_75t_L g894 ( 
.A(n_841),
.Y(n_894)
);

AOI21xp5_ASAP7_75t_L g895 ( 
.A1(n_852),
.A2(n_870),
.B(n_874),
.Y(n_895)
);

NOR2xp33_ASAP7_75t_L g896 ( 
.A(n_842),
.B(n_857),
.Y(n_896)
);

BUFx3_ASAP7_75t_L g897 ( 
.A(n_849),
.Y(n_897)
);

NOR2xp33_ASAP7_75t_R g898 ( 
.A(n_873),
.B(n_793),
.Y(n_898)
);

CKINVDCx11_ASAP7_75t_R g899 ( 
.A(n_879),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_L g900 ( 
.A(n_857),
.B(n_880),
.Y(n_900)
);

OAI21xp33_ASAP7_75t_L g901 ( 
.A1(n_844),
.A2(n_850),
.B(n_880),
.Y(n_901)
);

BUFx3_ASAP7_75t_L g902 ( 
.A(n_768),
.Y(n_902)
);

AND2x4_ASAP7_75t_L g903 ( 
.A(n_792),
.B(n_806),
.Y(n_903)
);

BUFx2_ASAP7_75t_SL g904 ( 
.A(n_790),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_L g905 ( 
.A(n_766),
.B(n_785),
.Y(n_905)
);

INVx3_ASAP7_75t_L g906 ( 
.A(n_815),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_L g907 ( 
.A(n_766),
.B(n_785),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_788),
.Y(n_908)
);

INVx4_ASAP7_75t_L g909 ( 
.A(n_774),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_798),
.Y(n_910)
);

AND2x4_ASAP7_75t_L g911 ( 
.A(n_792),
.B(n_806),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_835),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_L g913 ( 
.A(n_837),
.B(n_778),
.Y(n_913)
);

NOR2xp67_ASAP7_75t_L g914 ( 
.A(n_843),
.B(n_803),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_L g915 ( 
.A(n_778),
.B(n_770),
.Y(n_915)
);

AND2x4_ASAP7_75t_L g916 ( 
.A(n_868),
.B(n_826),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_SL g917 ( 
.A(n_775),
.B(n_770),
.Y(n_917)
);

INVx1_ASAP7_75t_SL g918 ( 
.A(n_861),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_L g919 ( 
.A(n_871),
.B(n_855),
.Y(n_919)
);

BUFx2_ASAP7_75t_L g920 ( 
.A(n_879),
.Y(n_920)
);

OAI21xp33_ASAP7_75t_L g921 ( 
.A1(n_881),
.A2(n_882),
.B(n_801),
.Y(n_921)
);

NAND2x1_ASAP7_75t_L g922 ( 
.A(n_854),
.B(n_876),
.Y(n_922)
);

NOR2xp33_ASAP7_75t_L g923 ( 
.A(n_871),
.B(n_775),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_L g924 ( 
.A(n_882),
.B(n_838),
.Y(n_924)
);

AOI22xp33_ASAP7_75t_L g925 ( 
.A1(n_845),
.A2(n_878),
.B1(n_779),
.B2(n_801),
.Y(n_925)
);

AND2x4_ASAP7_75t_L g926 ( 
.A(n_868),
.B(n_831),
.Y(n_926)
);

CKINVDCx12_ASAP7_75t_R g927 ( 
.A(n_780),
.Y(n_927)
);

AND2x2_ASAP7_75t_L g928 ( 
.A(n_839),
.B(n_772),
.Y(n_928)
);

INVxp67_ASAP7_75t_L g929 ( 
.A(n_819),
.Y(n_929)
);

AND2x2_ASAP7_75t_L g930 ( 
.A(n_830),
.B(n_786),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_L g931 ( 
.A(n_784),
.B(n_800),
.Y(n_931)
);

BUFx2_ASAP7_75t_L g932 ( 
.A(n_780),
.Y(n_932)
);

BUFx3_ASAP7_75t_L g933 ( 
.A(n_793),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_L g934 ( 
.A(n_804),
.B(n_814),
.Y(n_934)
);

NAND2xp33_ASAP7_75t_L g935 ( 
.A(n_781),
.B(n_820),
.Y(n_935)
);

BUFx6f_ASAP7_75t_L g936 ( 
.A(n_864),
.Y(n_936)
);

AOI22xp33_ASAP7_75t_L g937 ( 
.A1(n_797),
.A2(n_805),
.B1(n_789),
.B2(n_847),
.Y(n_937)
);

INVx2_ASAP7_75t_SL g938 ( 
.A(n_832),
.Y(n_938)
);

NOR2xp67_ASAP7_75t_L g939 ( 
.A(n_809),
.B(n_816),
.Y(n_939)
);

AOI22xp33_ASAP7_75t_L g940 ( 
.A1(n_805),
.A2(n_807),
.B1(n_804),
.B2(n_782),
.Y(n_940)
);

AND2x4_ASAP7_75t_L g941 ( 
.A(n_809),
.B(n_816),
.Y(n_941)
);

OR2x2_ASAP7_75t_L g942 ( 
.A(n_829),
.B(n_820),
.Y(n_942)
);

AND2x2_ASAP7_75t_L g943 ( 
.A(n_829),
.B(n_828),
.Y(n_943)
);

INVx3_ASAP7_75t_SL g944 ( 
.A(n_790),
.Y(n_944)
);

INVx1_ASAP7_75t_L g945 ( 
.A(n_811),
.Y(n_945)
);

NOR2xp33_ASAP7_75t_SL g946 ( 
.A(n_790),
.B(n_834),
.Y(n_946)
);

BUFx3_ASAP7_75t_L g947 ( 
.A(n_780),
.Y(n_947)
);

NOR2xp33_ASAP7_75t_L g948 ( 
.A(n_825),
.B(n_827),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_L g949 ( 
.A(n_825),
.B(n_829),
.Y(n_949)
);

AND2x2_ASAP7_75t_L g950 ( 
.A(n_833),
.B(n_883),
.Y(n_950)
);

AND2x4_ASAP7_75t_L g951 ( 
.A(n_866),
.B(n_876),
.Y(n_951)
);

BUFx6f_ASAP7_75t_L g952 ( 
.A(n_866),
.Y(n_952)
);

BUFx6f_ASAP7_75t_L g953 ( 
.A(n_866),
.Y(n_953)
);

INVx2_ASAP7_75t_SL g954 ( 
.A(n_771),
.Y(n_954)
);

INVx2_ASAP7_75t_SL g955 ( 
.A(n_771),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_SL g956 ( 
.A(n_824),
.B(n_823),
.Y(n_956)
);

OR2x6_ASAP7_75t_SL g957 ( 
.A(n_848),
.B(n_865),
.Y(n_957)
);

AOI22xp33_ASAP7_75t_L g958 ( 
.A1(n_822),
.A2(n_773),
.B1(n_802),
.B2(n_821),
.Y(n_958)
);

AND2x2_ASAP7_75t_L g959 ( 
.A(n_777),
.B(n_877),
.Y(n_959)
);

AND2x2_ASAP7_75t_L g960 ( 
.A(n_777),
.B(n_877),
.Y(n_960)
);

INVx2_ASAP7_75t_L g961 ( 
.A(n_799),
.Y(n_961)
);

INVx3_ASAP7_75t_L g962 ( 
.A(n_854),
.Y(n_962)
);

CKINVDCx6p67_ASAP7_75t_R g963 ( 
.A(n_771),
.Y(n_963)
);

AND2x4_ASAP7_75t_L g964 ( 
.A(n_862),
.B(n_872),
.Y(n_964)
);

HB1xp67_ASAP7_75t_L g965 ( 
.A(n_846),
.Y(n_965)
);

CKINVDCx5p33_ASAP7_75t_R g966 ( 
.A(n_846),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_865),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_817),
.Y(n_968)
);

OR2x6_ASAP7_75t_L g969 ( 
.A(n_818),
.B(n_812),
.Y(n_969)
);

BUFx3_ASAP7_75t_L g970 ( 
.A(n_783),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_L g971 ( 
.A(n_783),
.B(n_869),
.Y(n_971)
);

A2O1A1Ixp33_ASAP7_75t_L g972 ( 
.A1(n_810),
.A2(n_813),
.B(n_859),
.C(n_860),
.Y(n_972)
);

BUFx4f_ASAP7_75t_L g973 ( 
.A(n_867),
.Y(n_973)
);

BUFx2_ASAP7_75t_L g974 ( 
.A(n_869),
.Y(n_974)
);

A2O1A1Ixp33_ASAP7_75t_SL g975 ( 
.A1(n_808),
.A2(n_794),
.B(n_795),
.C(n_767),
.Y(n_975)
);

AND2x2_ASAP7_75t_L g976 ( 
.A(n_875),
.B(n_756),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_769),
.Y(n_977)
);

OAI21x1_ASAP7_75t_L g978 ( 
.A1(n_818),
.A2(n_791),
.B(n_813),
.Y(n_978)
);

INVx2_ASAP7_75t_SL g979 ( 
.A(n_841),
.Y(n_979)
);

AND2x2_ASAP7_75t_L g980 ( 
.A(n_881),
.B(n_756),
.Y(n_980)
);

INVx1_ASAP7_75t_L g981 ( 
.A(n_769),
.Y(n_981)
);

NAND3xp33_ASAP7_75t_L g982 ( 
.A(n_844),
.B(n_509),
.C(n_755),
.Y(n_982)
);

AND2x2_ASAP7_75t_L g983 ( 
.A(n_881),
.B(n_756),
.Y(n_983)
);

INVx1_ASAP7_75t_L g984 ( 
.A(n_769),
.Y(n_984)
);

OAI22xp5_ASAP7_75t_SL g985 ( 
.A1(n_844),
.A2(n_509),
.B1(n_648),
.B2(n_372),
.Y(n_985)
);

AND2x2_ASAP7_75t_L g986 ( 
.A(n_881),
.B(n_756),
.Y(n_986)
);

BUFx2_ASAP7_75t_L g987 ( 
.A(n_879),
.Y(n_987)
);

AOI21xp5_ASAP7_75t_L g988 ( 
.A1(n_776),
.A2(n_509),
.B(n_852),
.Y(n_988)
);

NAND2x1p5_ASAP7_75t_L g989 ( 
.A(n_774),
.B(n_864),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_SL g990 ( 
.A(n_844),
.B(n_850),
.Y(n_990)
);

AOI21xp5_ASAP7_75t_L g991 ( 
.A1(n_776),
.A2(n_509),
.B(n_852),
.Y(n_991)
);

INVx4_ASAP7_75t_L g992 ( 
.A(n_774),
.Y(n_992)
);

AND2x2_ASAP7_75t_L g993 ( 
.A(n_881),
.B(n_756),
.Y(n_993)
);

OAI22xp5_ASAP7_75t_L g994 ( 
.A1(n_844),
.A2(n_850),
.B1(n_509),
.B2(n_836),
.Y(n_994)
);

BUFx6f_ASAP7_75t_L g995 ( 
.A(n_774),
.Y(n_995)
);

OR2x6_ASAP7_75t_L g996 ( 
.A(n_834),
.B(n_879),
.Y(n_996)
);

CKINVDCx5p33_ASAP7_75t_R g997 ( 
.A(n_873),
.Y(n_997)
);

A2O1A1Ixp33_ASAP7_75t_SL g998 ( 
.A1(n_852),
.A2(n_509),
.B(n_612),
.C(n_870),
.Y(n_998)
);

AND2x4_ASAP7_75t_L g999 ( 
.A(n_792),
.B(n_806),
.Y(n_999)
);

INVx1_ASAP7_75t_SL g1000 ( 
.A(n_768),
.Y(n_1000)
);

NAND2x1p5_ASAP7_75t_L g1001 ( 
.A(n_774),
.B(n_864),
.Y(n_1001)
);

NOR2xp33_ASAP7_75t_L g1002 ( 
.A(n_765),
.B(n_509),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_L g1003 ( 
.A(n_765),
.B(n_739),
.Y(n_1003)
);

BUFx10_ASAP7_75t_L g1004 ( 
.A(n_828),
.Y(n_1004)
);

INVxp33_ASAP7_75t_L g1005 ( 
.A(n_768),
.Y(n_1005)
);

NOR2xp33_ASAP7_75t_L g1006 ( 
.A(n_765),
.B(n_509),
.Y(n_1006)
);

AND2x2_ASAP7_75t_L g1007 ( 
.A(n_881),
.B(n_756),
.Y(n_1007)
);

AND2x4_ASAP7_75t_L g1008 ( 
.A(n_792),
.B(n_806),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_769),
.Y(n_1009)
);

HB1xp67_ASAP7_75t_L g1010 ( 
.A(n_881),
.Y(n_1010)
);

AND2x2_ASAP7_75t_L g1011 ( 
.A(n_928),
.B(n_980),
.Y(n_1011)
);

CKINVDCx20_ASAP7_75t_R g1012 ( 
.A(n_899),
.Y(n_1012)
);

BUFx5_ASAP7_75t_L g1013 ( 
.A(n_968),
.Y(n_1013)
);

INVx1_ASAP7_75t_L g1014 ( 
.A(n_908),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_910),
.Y(n_1015)
);

INVx1_ASAP7_75t_L g1016 ( 
.A(n_912),
.Y(n_1016)
);

INVx2_ASAP7_75t_SL g1017 ( 
.A(n_889),
.Y(n_1017)
);

INVx1_ASAP7_75t_L g1018 ( 
.A(n_977),
.Y(n_1018)
);

AOI21x1_ASAP7_75t_L g1019 ( 
.A1(n_956),
.A2(n_917),
.B(n_931),
.Y(n_1019)
);

OAI22xp33_ASAP7_75t_L g1020 ( 
.A1(n_1003),
.A2(n_900),
.B1(n_890),
.B2(n_885),
.Y(n_1020)
);

NAND2x1p5_ASAP7_75t_L g1021 ( 
.A(n_909),
.B(n_992),
.Y(n_1021)
);

BUFx3_ASAP7_75t_L g1022 ( 
.A(n_894),
.Y(n_1022)
);

INVxp67_ASAP7_75t_L g1023 ( 
.A(n_930),
.Y(n_1023)
);

AOI22xp33_ASAP7_75t_L g1024 ( 
.A1(n_990),
.A2(n_901),
.B1(n_985),
.B2(n_994),
.Y(n_1024)
);

CKINVDCx20_ASAP7_75t_R g1025 ( 
.A(n_899),
.Y(n_1025)
);

INVx1_ASAP7_75t_L g1026 ( 
.A(n_981),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_984),
.Y(n_1027)
);

OAI22xp5_ASAP7_75t_L g1028 ( 
.A1(n_1002),
.A2(n_1006),
.B1(n_896),
.B2(n_887),
.Y(n_1028)
);

CKINVDCx11_ASAP7_75t_R g1029 ( 
.A(n_944),
.Y(n_1029)
);

INVx2_ASAP7_75t_L g1030 ( 
.A(n_1009),
.Y(n_1030)
);

INVx2_ASAP7_75t_SL g1031 ( 
.A(n_889),
.Y(n_1031)
);

INVx3_ASAP7_75t_L g1032 ( 
.A(n_906),
.Y(n_1032)
);

INVxp33_ASAP7_75t_L g1033 ( 
.A(n_983),
.Y(n_1033)
);

INVx2_ASAP7_75t_L g1034 ( 
.A(n_945),
.Y(n_1034)
);

OAI21xp5_ASAP7_75t_L g1035 ( 
.A1(n_982),
.A2(n_1006),
.B(n_1002),
.Y(n_1035)
);

AND2x2_ASAP7_75t_L g1036 ( 
.A(n_986),
.B(n_993),
.Y(n_1036)
);

AND2x2_ASAP7_75t_L g1037 ( 
.A(n_1007),
.B(n_892),
.Y(n_1037)
);

BUFx3_ASAP7_75t_L g1038 ( 
.A(n_897),
.Y(n_1038)
);

AOI22xp33_ASAP7_75t_L g1039 ( 
.A1(n_923),
.A2(n_925),
.B1(n_921),
.B2(n_895),
.Y(n_1039)
);

AOI22xp5_ASAP7_75t_L g1040 ( 
.A1(n_926),
.A2(n_938),
.B1(n_943),
.B2(n_916),
.Y(n_1040)
);

BUFx6f_ASAP7_75t_L g1041 ( 
.A(n_936),
.Y(n_1041)
);

INVx3_ASAP7_75t_L g1042 ( 
.A(n_906),
.Y(n_1042)
);

NAND2xp5_ASAP7_75t_L g1043 ( 
.A(n_913),
.B(n_924),
.Y(n_1043)
);

AOI22xp33_ASAP7_75t_L g1044 ( 
.A1(n_925),
.A2(n_895),
.B1(n_937),
.B2(n_919),
.Y(n_1044)
);

INVx11_ASAP7_75t_L g1045 ( 
.A(n_963),
.Y(n_1045)
);

AOI22xp33_ASAP7_75t_L g1046 ( 
.A1(n_937),
.A2(n_888),
.B1(n_915),
.B2(n_991),
.Y(n_1046)
);

NOR2xp33_ASAP7_75t_L g1047 ( 
.A(n_929),
.B(n_1005),
.Y(n_1047)
);

INVx2_ASAP7_75t_SL g1048 ( 
.A(n_902),
.Y(n_1048)
);

AOI22xp33_ASAP7_75t_L g1049 ( 
.A1(n_888),
.A2(n_991),
.B1(n_988),
.B2(n_1010),
.Y(n_1049)
);

INVx1_ASAP7_75t_SL g1050 ( 
.A(n_918),
.Y(n_1050)
);

NAND2x1p5_ASAP7_75t_L g1051 ( 
.A(n_909),
.B(n_992),
.Y(n_1051)
);

AND2x2_ASAP7_75t_L g1052 ( 
.A(n_903),
.B(n_911),
.Y(n_1052)
);

AOI22xp5_ASAP7_75t_L g1053 ( 
.A1(n_926),
.A2(n_916),
.B1(n_946),
.B2(n_920),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_1010),
.Y(n_1054)
);

AND2x2_ASAP7_75t_L g1055 ( 
.A(n_903),
.B(n_911),
.Y(n_1055)
);

INVx4_ASAP7_75t_L g1056 ( 
.A(n_936),
.Y(n_1056)
);

CKINVDCx11_ASAP7_75t_R g1057 ( 
.A(n_944),
.Y(n_1057)
);

AOI22xp33_ASAP7_75t_L g1058 ( 
.A1(n_929),
.A2(n_940),
.B1(n_976),
.B2(n_934),
.Y(n_1058)
);

INVxp33_ASAP7_75t_L g1059 ( 
.A(n_1005),
.Y(n_1059)
);

OR2x6_ASAP7_75t_L g1060 ( 
.A(n_891),
.B(n_996),
.Y(n_1060)
);

OAI21xp33_ASAP7_75t_L g1061 ( 
.A1(n_884),
.A2(n_940),
.B(n_948),
.Y(n_1061)
);

OAI22xp5_ASAP7_75t_L g1062 ( 
.A1(n_1000),
.A2(n_891),
.B1(n_996),
.B2(n_966),
.Y(n_1062)
);

BUFx3_ASAP7_75t_L g1063 ( 
.A(n_902),
.Y(n_1063)
);

AOI22xp33_ASAP7_75t_L g1064 ( 
.A1(n_948),
.A2(n_973),
.B1(n_970),
.B2(n_1004),
.Y(n_1064)
);

CKINVDCx6p67_ASAP7_75t_R g1065 ( 
.A(n_933),
.Y(n_1065)
);

INVx1_ASAP7_75t_L g1066 ( 
.A(n_949),
.Y(n_1066)
);

BUFx6f_ASAP7_75t_L g1067 ( 
.A(n_952),
.Y(n_1067)
);

AOI21x1_ASAP7_75t_L g1068 ( 
.A1(n_969),
.A2(n_961),
.B(n_971),
.Y(n_1068)
);

AND2x2_ASAP7_75t_L g1069 ( 
.A(n_999),
.B(n_1008),
.Y(n_1069)
);

INVx1_ASAP7_75t_L g1070 ( 
.A(n_942),
.Y(n_1070)
);

INVx2_ASAP7_75t_L g1071 ( 
.A(n_970),
.Y(n_1071)
);

OA21x2_ASAP7_75t_L g1072 ( 
.A1(n_972),
.A2(n_958),
.B(n_974),
.Y(n_1072)
);

INVx1_ASAP7_75t_L g1073 ( 
.A(n_959),
.Y(n_1073)
);

AOI22xp33_ASAP7_75t_L g1074 ( 
.A1(n_973),
.A2(n_1004),
.B1(n_987),
.B2(n_932),
.Y(n_1074)
);

AOI22xp33_ASAP7_75t_L g1075 ( 
.A1(n_891),
.A2(n_996),
.B1(n_947),
.B2(n_998),
.Y(n_1075)
);

OAI21x1_ASAP7_75t_L g1076 ( 
.A1(n_975),
.A2(n_967),
.B(n_893),
.Y(n_1076)
);

INVx1_ASAP7_75t_L g1077 ( 
.A(n_960),
.Y(n_1077)
);

AOI22xp33_ASAP7_75t_L g1078 ( 
.A1(n_999),
.A2(n_1008),
.B1(n_935),
.B2(n_904),
.Y(n_1078)
);

INVx1_ASAP7_75t_L g1079 ( 
.A(n_965),
.Y(n_1079)
);

OAI22xp33_ASAP7_75t_SL g1080 ( 
.A1(n_957),
.A2(n_979),
.B1(n_969),
.B2(n_1001),
.Y(n_1080)
);

INVx2_ASAP7_75t_L g1081 ( 
.A(n_969),
.Y(n_1081)
);

CKINVDCx16_ASAP7_75t_R g1082 ( 
.A(n_898),
.Y(n_1082)
);

AOI22xp33_ASAP7_75t_L g1083 ( 
.A1(n_950),
.A2(n_898),
.B1(n_964),
.B2(n_997),
.Y(n_1083)
);

OAI221xp5_ASAP7_75t_L g1084 ( 
.A1(n_914),
.A2(n_939),
.B1(n_922),
.B2(n_893),
.C(n_886),
.Y(n_1084)
);

AND2x4_ASAP7_75t_L g1085 ( 
.A(n_964),
.B(n_941),
.Y(n_1085)
);

INVx1_ASAP7_75t_L g1086 ( 
.A(n_954),
.Y(n_1086)
);

INVx6_ASAP7_75t_L g1087 ( 
.A(n_952),
.Y(n_1087)
);

AOI22xp33_ASAP7_75t_L g1088 ( 
.A1(n_941),
.A2(n_962),
.B1(n_995),
.B2(n_952),
.Y(n_1088)
);

AND2x2_ASAP7_75t_L g1089 ( 
.A(n_955),
.B(n_951),
.Y(n_1089)
);

AOI22xp33_ASAP7_75t_L g1090 ( 
.A1(n_962),
.A2(n_953),
.B1(n_995),
.B2(n_951),
.Y(n_1090)
);

AOI21xp33_ASAP7_75t_L g1091 ( 
.A1(n_953),
.A2(n_995),
.B(n_989),
.Y(n_1091)
);

BUFx2_ASAP7_75t_L g1092 ( 
.A(n_953),
.Y(n_1092)
);

CKINVDCx11_ASAP7_75t_R g1093 ( 
.A(n_953),
.Y(n_1093)
);

BUFx8_ASAP7_75t_L g1094 ( 
.A(n_927),
.Y(n_1094)
);

BUFx2_ASAP7_75t_SL g1095 ( 
.A(n_1001),
.Y(n_1095)
);

INVx3_ASAP7_75t_L g1096 ( 
.A(n_886),
.Y(n_1096)
);

INVx2_ASAP7_75t_SL g1097 ( 
.A(n_889),
.Y(n_1097)
);

NAND2x1p5_ASAP7_75t_L g1098 ( 
.A(n_909),
.B(n_992),
.Y(n_1098)
);

HB1xp67_ASAP7_75t_L g1099 ( 
.A(n_1010),
.Y(n_1099)
);

BUFx4f_ASAP7_75t_SL g1100 ( 
.A(n_889),
.Y(n_1100)
);

CKINVDCx11_ASAP7_75t_R g1101 ( 
.A(n_944),
.Y(n_1101)
);

OAI21x1_ASAP7_75t_L g1102 ( 
.A1(n_978),
.A2(n_791),
.B(n_787),
.Y(n_1102)
);

INVx6_ASAP7_75t_L g1103 ( 
.A(n_936),
.Y(n_1103)
);

BUFx6f_ASAP7_75t_L g1104 ( 
.A(n_936),
.Y(n_1104)
);

AND2x2_ASAP7_75t_L g1105 ( 
.A(n_928),
.B(n_980),
.Y(n_1105)
);

AND2x2_ASAP7_75t_L g1106 ( 
.A(n_928),
.B(n_980),
.Y(n_1106)
);

INVxp33_ASAP7_75t_L g1107 ( 
.A(n_980),
.Y(n_1107)
);

NAND2xp5_ASAP7_75t_L g1108 ( 
.A(n_1002),
.B(n_739),
.Y(n_1108)
);

CKINVDCx12_ASAP7_75t_R g1109 ( 
.A(n_891),
.Y(n_1109)
);

OAI21x1_ASAP7_75t_SL g1110 ( 
.A1(n_905),
.A2(n_907),
.B(n_789),
.Y(n_1110)
);

HB1xp67_ASAP7_75t_L g1111 ( 
.A(n_1010),
.Y(n_1111)
);

AOI22xp33_ASAP7_75t_SL g1112 ( 
.A1(n_985),
.A2(n_509),
.B1(n_683),
.B2(n_648),
.Y(n_1112)
);

OAI22xp5_ASAP7_75t_L g1113 ( 
.A1(n_1003),
.A2(n_844),
.B1(n_850),
.B2(n_509),
.Y(n_1113)
);

INVx2_ASAP7_75t_SL g1114 ( 
.A(n_889),
.Y(n_1114)
);

HB1xp67_ASAP7_75t_L g1115 ( 
.A(n_1010),
.Y(n_1115)
);

INVxp33_ASAP7_75t_L g1116 ( 
.A(n_1011),
.Y(n_1116)
);

OR2x2_ASAP7_75t_L g1117 ( 
.A(n_1070),
.B(n_1066),
.Y(n_1117)
);

INVx2_ASAP7_75t_L g1118 ( 
.A(n_1013),
.Y(n_1118)
);

HB1xp67_ASAP7_75t_L g1119 ( 
.A(n_1099),
.Y(n_1119)
);

INVx3_ASAP7_75t_L g1120 ( 
.A(n_1081),
.Y(n_1120)
);

INVx2_ASAP7_75t_L g1121 ( 
.A(n_1013),
.Y(n_1121)
);

AOI21x1_ASAP7_75t_L g1122 ( 
.A1(n_1019),
.A2(n_1068),
.B(n_1102),
.Y(n_1122)
);

BUFx3_ASAP7_75t_L g1123 ( 
.A(n_1060),
.Y(n_1123)
);

INVx3_ASAP7_75t_L g1124 ( 
.A(n_1081),
.Y(n_1124)
);

OAI21x1_ASAP7_75t_SL g1125 ( 
.A1(n_1110),
.A2(n_1024),
.B(n_1035),
.Y(n_1125)
);

INVx2_ASAP7_75t_L g1126 ( 
.A(n_1013),
.Y(n_1126)
);

NOR2xp33_ASAP7_75t_SL g1127 ( 
.A(n_1082),
.B(n_1061),
.Y(n_1127)
);

HB1xp67_ASAP7_75t_L g1128 ( 
.A(n_1111),
.Y(n_1128)
);

HB1xp67_ASAP7_75t_L g1129 ( 
.A(n_1115),
.Y(n_1129)
);

AO21x2_ASAP7_75t_L g1130 ( 
.A1(n_1076),
.A2(n_1071),
.B(n_1113),
.Y(n_1130)
);

BUFx4f_ASAP7_75t_L g1131 ( 
.A(n_1060),
.Y(n_1131)
);

AND2x2_ASAP7_75t_L g1132 ( 
.A(n_1044),
.B(n_1049),
.Y(n_1132)
);

HB1xp67_ASAP7_75t_L g1133 ( 
.A(n_1054),
.Y(n_1133)
);

OR2x2_ASAP7_75t_L g1134 ( 
.A(n_1049),
.B(n_1044),
.Y(n_1134)
);

AND2x4_ASAP7_75t_L g1135 ( 
.A(n_1060),
.B(n_1034),
.Y(n_1135)
);

OA21x2_ASAP7_75t_L g1136 ( 
.A1(n_1046),
.A2(n_1039),
.B(n_1076),
.Y(n_1136)
);

NAND2xp5_ASAP7_75t_L g1137 ( 
.A(n_1028),
.B(n_1020),
.Y(n_1137)
);

INVx2_ASAP7_75t_L g1138 ( 
.A(n_1072),
.Y(n_1138)
);

AO21x1_ASAP7_75t_SL g1139 ( 
.A1(n_1024),
.A2(n_1046),
.B(n_1039),
.Y(n_1139)
);

INVx2_ASAP7_75t_L g1140 ( 
.A(n_1072),
.Y(n_1140)
);

OAI21x1_ASAP7_75t_L g1141 ( 
.A1(n_1072),
.A2(n_1075),
.B(n_1030),
.Y(n_1141)
);

BUFx3_ASAP7_75t_L g1142 ( 
.A(n_1094),
.Y(n_1142)
);

OAI21x1_ASAP7_75t_L g1143 ( 
.A1(n_1075),
.A2(n_1064),
.B(n_1042),
.Y(n_1143)
);

AND2x4_ASAP7_75t_L g1144 ( 
.A(n_1032),
.B(n_1042),
.Y(n_1144)
);

AO21x2_ASAP7_75t_L g1145 ( 
.A1(n_1014),
.A2(n_1018),
.B(n_1026),
.Y(n_1145)
);

INVx1_ASAP7_75t_L g1146 ( 
.A(n_1015),
.Y(n_1146)
);

INVx2_ASAP7_75t_L g1147 ( 
.A(n_1016),
.Y(n_1147)
);

HB1xp67_ASAP7_75t_L g1148 ( 
.A(n_1079),
.Y(n_1148)
);

INVx1_ASAP7_75t_L g1149 ( 
.A(n_1027),
.Y(n_1149)
);

AND2x2_ASAP7_75t_L g1150 ( 
.A(n_1037),
.B(n_1033),
.Y(n_1150)
);

INVxp67_ASAP7_75t_L g1151 ( 
.A(n_1047),
.Y(n_1151)
);

INVxp67_ASAP7_75t_L g1152 ( 
.A(n_1047),
.Y(n_1152)
);

AND2x2_ASAP7_75t_L g1153 ( 
.A(n_1033),
.B(n_1107),
.Y(n_1153)
);

OR2x2_ASAP7_75t_L g1154 ( 
.A(n_1058),
.B(n_1023),
.Y(n_1154)
);

HB1xp67_ASAP7_75t_L g1155 ( 
.A(n_1073),
.Y(n_1155)
);

NAND2xp5_ASAP7_75t_L g1156 ( 
.A(n_1108),
.B(n_1043),
.Y(n_1156)
);

BUFx2_ASAP7_75t_L g1157 ( 
.A(n_1040),
.Y(n_1157)
);

BUFx2_ASAP7_75t_L g1158 ( 
.A(n_1053),
.Y(n_1158)
);

AOI22xp33_ASAP7_75t_SL g1159 ( 
.A1(n_1112),
.A2(n_1094),
.B1(n_1062),
.B2(n_1012),
.Y(n_1159)
);

AND2x2_ASAP7_75t_L g1160 ( 
.A(n_1107),
.B(n_1058),
.Y(n_1160)
);

AOI22xp33_ASAP7_75t_L g1161 ( 
.A1(n_1059),
.A2(n_1074),
.B1(n_1083),
.B2(n_1106),
.Y(n_1161)
);

HB1xp67_ASAP7_75t_L g1162 ( 
.A(n_1077),
.Y(n_1162)
);

HB1xp67_ASAP7_75t_L g1163 ( 
.A(n_1109),
.Y(n_1163)
);

AND2x2_ASAP7_75t_L g1164 ( 
.A(n_1105),
.B(n_1036),
.Y(n_1164)
);

NOR2xp33_ASAP7_75t_L g1165 ( 
.A(n_1059),
.B(n_1050),
.Y(n_1165)
);

OAI21xp5_ASAP7_75t_L g1166 ( 
.A1(n_1078),
.A2(n_1088),
.B(n_1090),
.Y(n_1166)
);

INVxp33_ASAP7_75t_L g1167 ( 
.A(n_1052),
.Y(n_1167)
);

OA21x2_ASAP7_75t_L g1168 ( 
.A1(n_1090),
.A2(n_1083),
.B(n_1086),
.Y(n_1168)
);

INVxp67_ASAP7_75t_L g1169 ( 
.A(n_1063),
.Y(n_1169)
);

INVxp33_ASAP7_75t_L g1170 ( 
.A(n_1055),
.Y(n_1170)
);

OA21x2_ASAP7_75t_L g1171 ( 
.A1(n_1091),
.A2(n_1080),
.B(n_1092),
.Y(n_1171)
);

AND2x2_ASAP7_75t_L g1172 ( 
.A(n_1085),
.B(n_1069),
.Y(n_1172)
);

NAND2xp5_ASAP7_75t_L g1173 ( 
.A(n_1048),
.B(n_1063),
.Y(n_1173)
);

OR2x2_ASAP7_75t_L g1174 ( 
.A(n_1096),
.B(n_1085),
.Y(n_1174)
);

OR2x2_ASAP7_75t_L g1175 ( 
.A(n_1085),
.B(n_1114),
.Y(n_1175)
);

AND2x2_ASAP7_75t_L g1176 ( 
.A(n_1089),
.B(n_1041),
.Y(n_1176)
);

OR2x2_ASAP7_75t_L g1177 ( 
.A(n_1017),
.B(n_1097),
.Y(n_1177)
);

OR2x2_ASAP7_75t_L g1178 ( 
.A(n_1031),
.B(n_1056),
.Y(n_1178)
);

AND2x2_ASAP7_75t_L g1179 ( 
.A(n_1138),
.B(n_1067),
.Y(n_1179)
);

BUFx3_ASAP7_75t_L g1180 ( 
.A(n_1171),
.Y(n_1180)
);

INVxp67_ASAP7_75t_L g1181 ( 
.A(n_1145),
.Y(n_1181)
);

NAND2xp5_ASAP7_75t_L g1182 ( 
.A(n_1137),
.B(n_1041),
.Y(n_1182)
);

BUFx3_ASAP7_75t_L g1183 ( 
.A(n_1171),
.Y(n_1183)
);

NAND2xp5_ASAP7_75t_L g1184 ( 
.A(n_1137),
.B(n_1041),
.Y(n_1184)
);

AND2x2_ASAP7_75t_L g1185 ( 
.A(n_1136),
.B(n_1041),
.Y(n_1185)
);

AND2x2_ASAP7_75t_L g1186 ( 
.A(n_1136),
.B(n_1104),
.Y(n_1186)
);

AND2x2_ASAP7_75t_L g1187 ( 
.A(n_1136),
.B(n_1104),
.Y(n_1187)
);

AND2x2_ASAP7_75t_L g1188 ( 
.A(n_1140),
.B(n_1104),
.Y(n_1188)
);

INVx4_ASAP7_75t_L g1189 ( 
.A(n_1131),
.Y(n_1189)
);

INVx5_ASAP7_75t_L g1190 ( 
.A(n_1118),
.Y(n_1190)
);

BUFx2_ASAP7_75t_L g1191 ( 
.A(n_1141),
.Y(n_1191)
);

BUFx3_ASAP7_75t_L g1192 ( 
.A(n_1171),
.Y(n_1192)
);

HB1xp67_ASAP7_75t_L g1193 ( 
.A(n_1148),
.Y(n_1193)
);

HB1xp67_ASAP7_75t_L g1194 ( 
.A(n_1145),
.Y(n_1194)
);

INVx4_ASAP7_75t_L g1195 ( 
.A(n_1131),
.Y(n_1195)
);

HB1xp67_ASAP7_75t_L g1196 ( 
.A(n_1145),
.Y(n_1196)
);

INVxp67_ASAP7_75t_SL g1197 ( 
.A(n_1133),
.Y(n_1197)
);

BUFx2_ASAP7_75t_L g1198 ( 
.A(n_1141),
.Y(n_1198)
);

NAND2xp5_ASAP7_75t_L g1199 ( 
.A(n_1117),
.B(n_1094),
.Y(n_1199)
);

OR2x2_ASAP7_75t_SL g1200 ( 
.A(n_1134),
.B(n_1087),
.Y(n_1200)
);

INVx2_ASAP7_75t_L g1201 ( 
.A(n_1147),
.Y(n_1201)
);

AND2x2_ASAP7_75t_L g1202 ( 
.A(n_1121),
.B(n_1103),
.Y(n_1202)
);

AND2x4_ASAP7_75t_L g1203 ( 
.A(n_1126),
.B(n_1022),
.Y(n_1203)
);

AND2x2_ASAP7_75t_L g1204 ( 
.A(n_1132),
.B(n_1087),
.Y(n_1204)
);

OAI21x1_ASAP7_75t_SL g1205 ( 
.A1(n_1125),
.A2(n_1095),
.B(n_1084),
.Y(n_1205)
);

AND2x2_ASAP7_75t_L g1206 ( 
.A(n_1132),
.B(n_1087),
.Y(n_1206)
);

NAND3xp33_ASAP7_75t_L g1207 ( 
.A(n_1182),
.B(n_1127),
.C(n_1161),
.Y(n_1207)
);

OAI221xp5_ASAP7_75t_L g1208 ( 
.A1(n_1199),
.A2(n_1159),
.B1(n_1127),
.B2(n_1163),
.C(n_1156),
.Y(n_1208)
);

NAND2xp5_ASAP7_75t_L g1209 ( 
.A(n_1193),
.B(n_1153),
.Y(n_1209)
);

AND2x2_ASAP7_75t_L g1210 ( 
.A(n_1179),
.B(n_1153),
.Y(n_1210)
);

AND2x2_ASAP7_75t_L g1211 ( 
.A(n_1179),
.B(n_1130),
.Y(n_1211)
);

NAND2xp5_ASAP7_75t_L g1212 ( 
.A(n_1193),
.B(n_1119),
.Y(n_1212)
);

AOI221xp5_ASAP7_75t_L g1213 ( 
.A1(n_1182),
.A2(n_1125),
.B1(n_1151),
.B2(n_1152),
.C(n_1116),
.Y(n_1213)
);

NAND2xp5_ASAP7_75t_L g1214 ( 
.A(n_1197),
.B(n_1128),
.Y(n_1214)
);

INVx1_ASAP7_75t_L g1215 ( 
.A(n_1201),
.Y(n_1215)
);

NAND2xp5_ASAP7_75t_L g1216 ( 
.A(n_1197),
.B(n_1129),
.Y(n_1216)
);

OAI21xp33_ASAP7_75t_L g1217 ( 
.A1(n_1180),
.A2(n_1160),
.B(n_1154),
.Y(n_1217)
);

NAND3xp33_ASAP7_75t_L g1218 ( 
.A(n_1184),
.B(n_1154),
.C(n_1166),
.Y(n_1218)
);

OA21x2_ASAP7_75t_L g1219 ( 
.A1(n_1181),
.A2(n_1122),
.B(n_1143),
.Y(n_1219)
);

AOI22xp33_ASAP7_75t_SL g1220 ( 
.A1(n_1189),
.A2(n_1158),
.B1(n_1131),
.B2(n_1157),
.Y(n_1220)
);

NOR3xp33_ASAP7_75t_L g1221 ( 
.A(n_1199),
.B(n_1166),
.C(n_1158),
.Y(n_1221)
);

OAI21xp5_ASAP7_75t_SL g1222 ( 
.A1(n_1184),
.A2(n_1134),
.B(n_1157),
.Y(n_1222)
);

NAND4xp25_ASAP7_75t_L g1223 ( 
.A(n_1204),
.B(n_1165),
.C(n_1150),
.D(n_1164),
.Y(n_1223)
);

AOI22xp33_ASAP7_75t_L g1224 ( 
.A1(n_1189),
.A2(n_1139),
.B1(n_1131),
.B2(n_1123),
.Y(n_1224)
);

AND2x2_ASAP7_75t_L g1225 ( 
.A(n_1179),
.B(n_1130),
.Y(n_1225)
);

AOI221xp5_ASAP7_75t_L g1226 ( 
.A1(n_1180),
.A2(n_1150),
.B1(n_1192),
.B2(n_1183),
.C(n_1155),
.Y(n_1226)
);

OAI221xp5_ASAP7_75t_SL g1227 ( 
.A1(n_1180),
.A2(n_1160),
.B1(n_1142),
.B2(n_1123),
.C(n_1169),
.Y(n_1227)
);

OAI22xp5_ASAP7_75t_L g1228 ( 
.A1(n_1200),
.A2(n_1123),
.B1(n_1012),
.B2(n_1025),
.Y(n_1228)
);

AND2x2_ASAP7_75t_L g1229 ( 
.A(n_1179),
.B(n_1130),
.Y(n_1229)
);

NAND2xp5_ASAP7_75t_L g1230 ( 
.A(n_1203),
.B(n_1135),
.Y(n_1230)
);

OAI21xp5_ASAP7_75t_SL g1231 ( 
.A1(n_1206),
.A2(n_1170),
.B(n_1167),
.Y(n_1231)
);

NAND2xp5_ASAP7_75t_L g1232 ( 
.A(n_1203),
.B(n_1135),
.Y(n_1232)
);

NAND2xp5_ASAP7_75t_L g1233 ( 
.A(n_1203),
.B(n_1135),
.Y(n_1233)
);

NAND2xp5_ASAP7_75t_SL g1234 ( 
.A(n_1205),
.B(n_1135),
.Y(n_1234)
);

OAI21xp5_ASAP7_75t_SL g1235 ( 
.A1(n_1206),
.A2(n_1204),
.B(n_1172),
.Y(n_1235)
);

NAND2xp5_ASAP7_75t_L g1236 ( 
.A(n_1203),
.B(n_1146),
.Y(n_1236)
);

NAND2xp5_ASAP7_75t_L g1237 ( 
.A(n_1203),
.B(n_1146),
.Y(n_1237)
);

NAND3xp33_ASAP7_75t_L g1238 ( 
.A(n_1180),
.B(n_1168),
.C(n_1171),
.Y(n_1238)
);

NAND2xp5_ASAP7_75t_L g1239 ( 
.A(n_1203),
.B(n_1206),
.Y(n_1239)
);

NAND2xp5_ASAP7_75t_SL g1240 ( 
.A(n_1205),
.B(n_1144),
.Y(n_1240)
);

AOI22xp33_ASAP7_75t_SL g1241 ( 
.A1(n_1189),
.A2(n_1168),
.B1(n_1142),
.B2(n_1143),
.Y(n_1241)
);

NAND2xp5_ASAP7_75t_L g1242 ( 
.A(n_1206),
.B(n_1149),
.Y(n_1242)
);

OAI22xp5_ASAP7_75t_L g1243 ( 
.A1(n_1200),
.A2(n_1025),
.B1(n_1142),
.B2(n_1175),
.Y(n_1243)
);

OAI21xp5_ASAP7_75t_SL g1244 ( 
.A1(n_1204),
.A2(n_1172),
.B(n_1191),
.Y(n_1244)
);

OAI22xp5_ASAP7_75t_L g1245 ( 
.A1(n_1200),
.A2(n_1175),
.B1(n_1174),
.B2(n_1177),
.Y(n_1245)
);

NOR3xp33_ASAP7_75t_L g1246 ( 
.A(n_1189),
.B(n_1173),
.C(n_1101),
.Y(n_1246)
);

AND2x2_ASAP7_75t_L g1247 ( 
.A(n_1188),
.B(n_1120),
.Y(n_1247)
);

NAND3xp33_ASAP7_75t_L g1248 ( 
.A(n_1183),
.B(n_1168),
.C(n_1162),
.Y(n_1248)
);

OAI22xp5_ASAP7_75t_L g1249 ( 
.A1(n_1189),
.A2(n_1174),
.B1(n_1177),
.B2(n_1168),
.Y(n_1249)
);

AND2x2_ASAP7_75t_L g1250 ( 
.A(n_1185),
.B(n_1120),
.Y(n_1250)
);

NOR2xp33_ASAP7_75t_L g1251 ( 
.A(n_1189),
.B(n_1164),
.Y(n_1251)
);

OAI21xp5_ASAP7_75t_SL g1252 ( 
.A1(n_1191),
.A2(n_1139),
.B(n_1176),
.Y(n_1252)
);

NOR2xp33_ASAP7_75t_R g1253 ( 
.A(n_1195),
.B(n_1093),
.Y(n_1253)
);

AND2x2_ASAP7_75t_L g1254 ( 
.A(n_1185),
.B(n_1124),
.Y(n_1254)
);

NAND2xp5_ASAP7_75t_L g1255 ( 
.A(n_1202),
.B(n_1149),
.Y(n_1255)
);

NAND2xp5_ASAP7_75t_SL g1256 ( 
.A(n_1205),
.B(n_1144),
.Y(n_1256)
);

AND2x4_ASAP7_75t_SL g1257 ( 
.A(n_1246),
.B(n_1195),
.Y(n_1257)
);

INVx1_ASAP7_75t_L g1258 ( 
.A(n_1215),
.Y(n_1258)
);

AND2x2_ASAP7_75t_L g1259 ( 
.A(n_1210),
.B(n_1250),
.Y(n_1259)
);

AND2x2_ASAP7_75t_L g1260 ( 
.A(n_1210),
.B(n_1185),
.Y(n_1260)
);

OR2x2_ASAP7_75t_L g1261 ( 
.A(n_1209),
.B(n_1183),
.Y(n_1261)
);

OR2x2_ASAP7_75t_L g1262 ( 
.A(n_1236),
.B(n_1183),
.Y(n_1262)
);

INVx1_ASAP7_75t_L g1263 ( 
.A(n_1215),
.Y(n_1263)
);

INVx1_ASAP7_75t_L g1264 ( 
.A(n_1255),
.Y(n_1264)
);

INVx1_ASAP7_75t_L g1265 ( 
.A(n_1237),
.Y(n_1265)
);

INVxp67_ASAP7_75t_L g1266 ( 
.A(n_1214),
.Y(n_1266)
);

INVx4_ASAP7_75t_L g1267 ( 
.A(n_1219),
.Y(n_1267)
);

INVx1_ASAP7_75t_L g1268 ( 
.A(n_1216),
.Y(n_1268)
);

NAND2xp5_ASAP7_75t_L g1269 ( 
.A(n_1242),
.B(n_1194),
.Y(n_1269)
);

HB1xp67_ASAP7_75t_L g1270 ( 
.A(n_1212),
.Y(n_1270)
);

AND2x4_ASAP7_75t_L g1271 ( 
.A(n_1240),
.B(n_1192),
.Y(n_1271)
);

OR2x2_ASAP7_75t_L g1272 ( 
.A(n_1239),
.B(n_1192),
.Y(n_1272)
);

INVx1_ASAP7_75t_L g1273 ( 
.A(n_1254),
.Y(n_1273)
);

OR2x2_ASAP7_75t_L g1274 ( 
.A(n_1211),
.B(n_1192),
.Y(n_1274)
);

NOR2xp33_ASAP7_75t_L g1275 ( 
.A(n_1223),
.B(n_1029),
.Y(n_1275)
);

AND2x4_ASAP7_75t_L g1276 ( 
.A(n_1240),
.B(n_1190),
.Y(n_1276)
);

AND2x4_ASAP7_75t_L g1277 ( 
.A(n_1256),
.B(n_1190),
.Y(n_1277)
);

INVx3_ASAP7_75t_L g1278 ( 
.A(n_1211),
.Y(n_1278)
);

INVx1_ASAP7_75t_L g1279 ( 
.A(n_1247),
.Y(n_1279)
);

INVx1_ASAP7_75t_L g1280 ( 
.A(n_1225),
.Y(n_1280)
);

AND2x2_ASAP7_75t_L g1281 ( 
.A(n_1225),
.B(n_1186),
.Y(n_1281)
);

INVx2_ASAP7_75t_L g1282 ( 
.A(n_1229),
.Y(n_1282)
);

NOR2xp33_ASAP7_75t_L g1283 ( 
.A(n_1208),
.B(n_1029),
.Y(n_1283)
);

AND2x2_ASAP7_75t_L g1284 ( 
.A(n_1229),
.B(n_1186),
.Y(n_1284)
);

NOR2xp67_ASAP7_75t_L g1285 ( 
.A(n_1248),
.B(n_1181),
.Y(n_1285)
);

NAND2xp5_ASAP7_75t_L g1286 ( 
.A(n_1226),
.B(n_1217),
.Y(n_1286)
);

INVx2_ASAP7_75t_L g1287 ( 
.A(n_1219),
.Y(n_1287)
);

AND2x2_ASAP7_75t_L g1288 ( 
.A(n_1244),
.B(n_1186),
.Y(n_1288)
);

AND2x2_ASAP7_75t_L g1289 ( 
.A(n_1230),
.B(n_1187),
.Y(n_1289)
);

BUFx6f_ASAP7_75t_L g1290 ( 
.A(n_1219),
.Y(n_1290)
);

INVxp67_ASAP7_75t_L g1291 ( 
.A(n_1251),
.Y(n_1291)
);

INVx1_ASAP7_75t_L g1292 ( 
.A(n_1232),
.Y(n_1292)
);

AND2x2_ASAP7_75t_L g1293 ( 
.A(n_1233),
.B(n_1187),
.Y(n_1293)
);

NAND2xp5_ASAP7_75t_L g1294 ( 
.A(n_1218),
.B(n_1194),
.Y(n_1294)
);

INVx1_ASAP7_75t_L g1295 ( 
.A(n_1258),
.Y(n_1295)
);

OR2x2_ASAP7_75t_L g1296 ( 
.A(n_1294),
.B(n_1238),
.Y(n_1296)
);

NAND2xp5_ASAP7_75t_L g1297 ( 
.A(n_1266),
.B(n_1221),
.Y(n_1297)
);

INVx1_ASAP7_75t_L g1298 ( 
.A(n_1258),
.Y(n_1298)
);

AND2x2_ASAP7_75t_L g1299 ( 
.A(n_1288),
.B(n_1241),
.Y(n_1299)
);

AND2x2_ASAP7_75t_L g1300 ( 
.A(n_1288),
.B(n_1187),
.Y(n_1300)
);

INVx2_ASAP7_75t_L g1301 ( 
.A(n_1287),
.Y(n_1301)
);

INVx2_ASAP7_75t_L g1302 ( 
.A(n_1287),
.Y(n_1302)
);

AOI22xp5_ASAP7_75t_L g1303 ( 
.A1(n_1283),
.A2(n_1207),
.B1(n_1222),
.B2(n_1228),
.Y(n_1303)
);

NAND2xp5_ASAP7_75t_L g1304 ( 
.A(n_1266),
.B(n_1235),
.Y(n_1304)
);

NAND2xp5_ASAP7_75t_L g1305 ( 
.A(n_1268),
.B(n_1213),
.Y(n_1305)
);

OR2x2_ASAP7_75t_L g1306 ( 
.A(n_1294),
.B(n_1249),
.Y(n_1306)
);

NOR2x1p5_ASAP7_75t_SL g1307 ( 
.A(n_1287),
.B(n_1274),
.Y(n_1307)
);

AND2x2_ASAP7_75t_L g1308 ( 
.A(n_1281),
.B(n_1191),
.Y(n_1308)
);

INVx3_ASAP7_75t_L g1309 ( 
.A(n_1276),
.Y(n_1309)
);

INVx1_ASAP7_75t_L g1310 ( 
.A(n_1263),
.Y(n_1310)
);

NAND2xp5_ASAP7_75t_L g1311 ( 
.A(n_1268),
.B(n_1252),
.Y(n_1311)
);

INVxp67_ASAP7_75t_L g1312 ( 
.A(n_1270),
.Y(n_1312)
);

INVx3_ASAP7_75t_R g1313 ( 
.A(n_1271),
.Y(n_1313)
);

INVx1_ASAP7_75t_L g1314 ( 
.A(n_1263),
.Y(n_1314)
);

AND2x4_ASAP7_75t_L g1315 ( 
.A(n_1276),
.B(n_1234),
.Y(n_1315)
);

NAND2xp5_ASAP7_75t_L g1316 ( 
.A(n_1265),
.B(n_1231),
.Y(n_1316)
);

INVx1_ASAP7_75t_L g1317 ( 
.A(n_1265),
.Y(n_1317)
);

INVx2_ASAP7_75t_L g1318 ( 
.A(n_1290),
.Y(n_1318)
);

AND2x2_ASAP7_75t_L g1319 ( 
.A(n_1281),
.B(n_1198),
.Y(n_1319)
);

INVx1_ASAP7_75t_L g1320 ( 
.A(n_1273),
.Y(n_1320)
);

INVx1_ASAP7_75t_SL g1321 ( 
.A(n_1261),
.Y(n_1321)
);

AND2x2_ASAP7_75t_L g1322 ( 
.A(n_1284),
.B(n_1198),
.Y(n_1322)
);

AND2x2_ASAP7_75t_L g1323 ( 
.A(n_1284),
.B(n_1198),
.Y(n_1323)
);

AND2x4_ASAP7_75t_L g1324 ( 
.A(n_1276),
.B(n_1234),
.Y(n_1324)
);

AND2x2_ASAP7_75t_L g1325 ( 
.A(n_1260),
.B(n_1202),
.Y(n_1325)
);

NAND2xp5_ASAP7_75t_L g1326 ( 
.A(n_1292),
.B(n_1202),
.Y(n_1326)
);

INVxp67_ASAP7_75t_L g1327 ( 
.A(n_1275),
.Y(n_1327)
);

INVx1_ASAP7_75t_L g1328 ( 
.A(n_1273),
.Y(n_1328)
);

NAND2xp5_ASAP7_75t_SL g1329 ( 
.A(n_1286),
.B(n_1253),
.Y(n_1329)
);

AND2x2_ASAP7_75t_L g1330 ( 
.A(n_1260),
.B(n_1278),
.Y(n_1330)
);

OR2x2_ASAP7_75t_L g1331 ( 
.A(n_1269),
.B(n_1196),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_1279),
.Y(n_1332)
);

INVx1_ASAP7_75t_L g1333 ( 
.A(n_1295),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_1295),
.Y(n_1334)
);

INVx1_ASAP7_75t_L g1335 ( 
.A(n_1298),
.Y(n_1335)
);

OR2x2_ASAP7_75t_L g1336 ( 
.A(n_1296),
.B(n_1269),
.Y(n_1336)
);

INVx1_ASAP7_75t_L g1337 ( 
.A(n_1298),
.Y(n_1337)
);

AOI21xp33_ASAP7_75t_L g1338 ( 
.A1(n_1296),
.A2(n_1286),
.B(n_1285),
.Y(n_1338)
);

OAI21xp5_ASAP7_75t_L g1339 ( 
.A1(n_1303),
.A2(n_1285),
.B(n_1271),
.Y(n_1339)
);

NAND2xp5_ASAP7_75t_L g1340 ( 
.A(n_1305),
.B(n_1291),
.Y(n_1340)
);

INVx1_ASAP7_75t_L g1341 ( 
.A(n_1310),
.Y(n_1341)
);

OR2x2_ASAP7_75t_L g1342 ( 
.A(n_1306),
.B(n_1282),
.Y(n_1342)
);

INVx1_ASAP7_75t_L g1343 ( 
.A(n_1310),
.Y(n_1343)
);

INVx1_ASAP7_75t_L g1344 ( 
.A(n_1314),
.Y(n_1344)
);

INVx1_ASAP7_75t_L g1345 ( 
.A(n_1314),
.Y(n_1345)
);

INVx1_ASAP7_75t_L g1346 ( 
.A(n_1317),
.Y(n_1346)
);

INVx1_ASAP7_75t_L g1347 ( 
.A(n_1317),
.Y(n_1347)
);

INVx1_ASAP7_75t_L g1348 ( 
.A(n_1320),
.Y(n_1348)
);

AOI221xp5_ASAP7_75t_L g1349 ( 
.A1(n_1297),
.A2(n_1271),
.B1(n_1292),
.B2(n_1264),
.C(n_1267),
.Y(n_1349)
);

OR2x2_ASAP7_75t_L g1350 ( 
.A(n_1306),
.B(n_1282),
.Y(n_1350)
);

NAND2xp5_ASAP7_75t_L g1351 ( 
.A(n_1312),
.B(n_1316),
.Y(n_1351)
);

NAND2x1p5_ASAP7_75t_L g1352 ( 
.A(n_1315),
.B(n_1276),
.Y(n_1352)
);

INVx2_ASAP7_75t_L g1353 ( 
.A(n_1301),
.Y(n_1353)
);

OR2x2_ASAP7_75t_L g1354 ( 
.A(n_1321),
.B(n_1282),
.Y(n_1354)
);

NOR5xp2_ASAP7_75t_L g1355 ( 
.A(n_1327),
.B(n_1227),
.C(n_1313),
.D(n_1307),
.E(n_1332),
.Y(n_1355)
);

NAND2xp5_ASAP7_75t_L g1356 ( 
.A(n_1304),
.B(n_1311),
.Y(n_1356)
);

NAND2xp5_ASAP7_75t_L g1357 ( 
.A(n_1303),
.B(n_1264),
.Y(n_1357)
);

NAND2xp5_ASAP7_75t_L g1358 ( 
.A(n_1325),
.B(n_1289),
.Y(n_1358)
);

INVx1_ASAP7_75t_L g1359 ( 
.A(n_1320),
.Y(n_1359)
);

INVx1_ASAP7_75t_L g1360 ( 
.A(n_1328),
.Y(n_1360)
);

NOR2xp67_ASAP7_75t_L g1361 ( 
.A(n_1309),
.B(n_1315),
.Y(n_1361)
);

INVx1_ASAP7_75t_L g1362 ( 
.A(n_1328),
.Y(n_1362)
);

AND2x2_ASAP7_75t_L g1363 ( 
.A(n_1315),
.B(n_1271),
.Y(n_1363)
);

INVx1_ASAP7_75t_L g1364 ( 
.A(n_1332),
.Y(n_1364)
);

NAND2xp5_ASAP7_75t_L g1365 ( 
.A(n_1325),
.B(n_1289),
.Y(n_1365)
);

INVx1_ASAP7_75t_SL g1366 ( 
.A(n_1329),
.Y(n_1366)
);

INVx2_ASAP7_75t_L g1367 ( 
.A(n_1301),
.Y(n_1367)
);

NAND2xp5_ASAP7_75t_L g1368 ( 
.A(n_1326),
.B(n_1293),
.Y(n_1368)
);

INVx1_ASAP7_75t_L g1369 ( 
.A(n_1301),
.Y(n_1369)
);

INVx1_ASAP7_75t_L g1370 ( 
.A(n_1302),
.Y(n_1370)
);

NOR2xp33_ASAP7_75t_L g1371 ( 
.A(n_1299),
.B(n_1261),
.Y(n_1371)
);

NAND2xp5_ASAP7_75t_L g1372 ( 
.A(n_1299),
.B(n_1293),
.Y(n_1372)
);

NAND2xp5_ASAP7_75t_L g1373 ( 
.A(n_1300),
.B(n_1259),
.Y(n_1373)
);

AND2x2_ASAP7_75t_L g1374 ( 
.A(n_1315),
.B(n_1324),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_1302),
.Y(n_1375)
);

INVx1_ASAP7_75t_L g1376 ( 
.A(n_1333),
.Y(n_1376)
);

OR2x2_ASAP7_75t_L g1377 ( 
.A(n_1336),
.B(n_1331),
.Y(n_1377)
);

AND2x2_ASAP7_75t_L g1378 ( 
.A(n_1374),
.B(n_1324),
.Y(n_1378)
);

NAND2xp5_ASAP7_75t_L g1379 ( 
.A(n_1356),
.B(n_1300),
.Y(n_1379)
);

BUFx2_ASAP7_75t_L g1380 ( 
.A(n_1374),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_1334),
.Y(n_1381)
);

AND2x2_ASAP7_75t_L g1382 ( 
.A(n_1361),
.B(n_1324),
.Y(n_1382)
);

INVx2_ASAP7_75t_L g1383 ( 
.A(n_1353),
.Y(n_1383)
);

NAND2xp5_ASAP7_75t_L g1384 ( 
.A(n_1366),
.B(n_1340),
.Y(n_1384)
);

NAND2x1p5_ASAP7_75t_L g1385 ( 
.A(n_1363),
.B(n_1324),
.Y(n_1385)
);

INVx1_ASAP7_75t_SL g1386 ( 
.A(n_1351),
.Y(n_1386)
);

BUFx3_ASAP7_75t_L g1387 ( 
.A(n_1352),
.Y(n_1387)
);

NOR2xp67_ASAP7_75t_L g1388 ( 
.A(n_1339),
.B(n_1309),
.Y(n_1388)
);

OR2x2_ASAP7_75t_L g1389 ( 
.A(n_1336),
.B(n_1331),
.Y(n_1389)
);

INVx1_ASAP7_75t_L g1390 ( 
.A(n_1335),
.Y(n_1390)
);

INVx1_ASAP7_75t_L g1391 ( 
.A(n_1337),
.Y(n_1391)
);

AND2x2_ASAP7_75t_L g1392 ( 
.A(n_1363),
.B(n_1309),
.Y(n_1392)
);

AND2x4_ASAP7_75t_L g1393 ( 
.A(n_1346),
.B(n_1307),
.Y(n_1393)
);

INVx1_ASAP7_75t_L g1394 ( 
.A(n_1341),
.Y(n_1394)
);

INVx1_ASAP7_75t_L g1395 ( 
.A(n_1343),
.Y(n_1395)
);

INVx1_ASAP7_75t_L g1396 ( 
.A(n_1344),
.Y(n_1396)
);

NAND2xp5_ASAP7_75t_L g1397 ( 
.A(n_1357),
.B(n_1330),
.Y(n_1397)
);

CKINVDCx5p33_ASAP7_75t_R g1398 ( 
.A(n_1371),
.Y(n_1398)
);

INVx1_ASAP7_75t_L g1399 ( 
.A(n_1345),
.Y(n_1399)
);

INVx2_ASAP7_75t_L g1400 ( 
.A(n_1353),
.Y(n_1400)
);

AND2x2_ASAP7_75t_L g1401 ( 
.A(n_1352),
.B(n_1309),
.Y(n_1401)
);

OR2x2_ASAP7_75t_L g1402 ( 
.A(n_1372),
.B(n_1318),
.Y(n_1402)
);

INVx1_ASAP7_75t_L g1403 ( 
.A(n_1348),
.Y(n_1403)
);

OR2x2_ASAP7_75t_L g1404 ( 
.A(n_1342),
.B(n_1318),
.Y(n_1404)
);

INVx4_ASAP7_75t_L g1405 ( 
.A(n_1367),
.Y(n_1405)
);

INVx1_ASAP7_75t_SL g1406 ( 
.A(n_1342),
.Y(n_1406)
);

NAND2xp5_ASAP7_75t_L g1407 ( 
.A(n_1371),
.B(n_1330),
.Y(n_1407)
);

INVx1_ASAP7_75t_L g1408 ( 
.A(n_1347),
.Y(n_1408)
);

AOI22xp33_ASAP7_75t_L g1409 ( 
.A1(n_1338),
.A2(n_1257),
.B1(n_1243),
.B2(n_1220),
.Y(n_1409)
);

NAND2xp5_ASAP7_75t_L g1410 ( 
.A(n_1349),
.B(n_1280),
.Y(n_1410)
);

INVx2_ASAP7_75t_L g1411 ( 
.A(n_1367),
.Y(n_1411)
);

AND2x2_ASAP7_75t_L g1412 ( 
.A(n_1378),
.B(n_1350),
.Y(n_1412)
);

INVx1_ASAP7_75t_L g1413 ( 
.A(n_1376),
.Y(n_1413)
);

INVx1_ASAP7_75t_L g1414 ( 
.A(n_1376),
.Y(n_1414)
);

AOI21xp33_ASAP7_75t_SL g1415 ( 
.A1(n_1398),
.A2(n_1355),
.B(n_1354),
.Y(n_1415)
);

INVx1_ASAP7_75t_L g1416 ( 
.A(n_1381),
.Y(n_1416)
);

OAI32xp33_ASAP7_75t_L g1417 ( 
.A1(n_1398),
.A2(n_1350),
.A3(n_1267),
.B1(n_1318),
.B2(n_1354),
.Y(n_1417)
);

INVx1_ASAP7_75t_L g1418 ( 
.A(n_1381),
.Y(n_1418)
);

OAI32xp33_ASAP7_75t_L g1419 ( 
.A1(n_1386),
.A2(n_1267),
.A3(n_1274),
.B1(n_1359),
.B2(n_1360),
.Y(n_1419)
);

AOI22xp33_ASAP7_75t_L g1420 ( 
.A1(n_1388),
.A2(n_1257),
.B1(n_1224),
.B2(n_1277),
.Y(n_1420)
);

OAI221xp5_ASAP7_75t_L g1421 ( 
.A1(n_1409),
.A2(n_1362),
.B1(n_1364),
.B2(n_1373),
.C(n_1368),
.Y(n_1421)
);

INVx1_ASAP7_75t_SL g1422 ( 
.A(n_1380),
.Y(n_1422)
);

NAND2xp5_ASAP7_75t_L g1423 ( 
.A(n_1384),
.B(n_1358),
.Y(n_1423)
);

HB1xp67_ASAP7_75t_L g1424 ( 
.A(n_1380),
.Y(n_1424)
);

AND2x2_ASAP7_75t_L g1425 ( 
.A(n_1378),
.B(n_1365),
.Y(n_1425)
);

AND2x2_ASAP7_75t_L g1426 ( 
.A(n_1392),
.B(n_1308),
.Y(n_1426)
);

AOI21xp33_ASAP7_75t_L g1427 ( 
.A1(n_1406),
.A2(n_1370),
.B(n_1369),
.Y(n_1427)
);

OAI21xp5_ASAP7_75t_L g1428 ( 
.A1(n_1410),
.A2(n_1375),
.B(n_1256),
.Y(n_1428)
);

NAND2xp5_ASAP7_75t_L g1429 ( 
.A(n_1397),
.B(n_1308),
.Y(n_1429)
);

AOI21xp5_ASAP7_75t_L g1430 ( 
.A1(n_1407),
.A2(n_1257),
.B(n_1277),
.Y(n_1430)
);

AOI22xp33_ASAP7_75t_L g1431 ( 
.A1(n_1387),
.A2(n_1277),
.B1(n_1195),
.B2(n_1245),
.Y(n_1431)
);

OAI322xp33_ASAP7_75t_L g1432 ( 
.A1(n_1402),
.A2(n_1267),
.A3(n_1290),
.B1(n_1302),
.B2(n_1262),
.C1(n_1280),
.C2(n_1272),
.Y(n_1432)
);

NAND2xp5_ASAP7_75t_L g1433 ( 
.A(n_1379),
.B(n_1319),
.Y(n_1433)
);

AND2x2_ASAP7_75t_L g1434 ( 
.A(n_1392),
.B(n_1319),
.Y(n_1434)
);

INVx1_ASAP7_75t_L g1435 ( 
.A(n_1390),
.Y(n_1435)
);

INVx1_ASAP7_75t_L g1436 ( 
.A(n_1390),
.Y(n_1436)
);

INVxp67_ASAP7_75t_SL g1437 ( 
.A(n_1385),
.Y(n_1437)
);

NOR2xp33_ASAP7_75t_L g1438 ( 
.A(n_1423),
.B(n_1387),
.Y(n_1438)
);

INVx1_ASAP7_75t_L g1439 ( 
.A(n_1424),
.Y(n_1439)
);

NAND2xp5_ASAP7_75t_L g1440 ( 
.A(n_1422),
.B(n_1395),
.Y(n_1440)
);

NAND2xp5_ASAP7_75t_L g1441 ( 
.A(n_1415),
.B(n_1396),
.Y(n_1441)
);

NAND2xp5_ASAP7_75t_L g1442 ( 
.A(n_1425),
.B(n_1408),
.Y(n_1442)
);

NAND2xp5_ASAP7_75t_L g1443 ( 
.A(n_1413),
.B(n_1391),
.Y(n_1443)
);

AND2x4_ASAP7_75t_L g1444 ( 
.A(n_1437),
.B(n_1401),
.Y(n_1444)
);

NAND2xp5_ASAP7_75t_L g1445 ( 
.A(n_1425),
.B(n_1412),
.Y(n_1445)
);

NAND2xp5_ASAP7_75t_L g1446 ( 
.A(n_1413),
.B(n_1391),
.Y(n_1446)
);

INVx1_ASAP7_75t_L g1447 ( 
.A(n_1414),
.Y(n_1447)
);

OR2x2_ASAP7_75t_L g1448 ( 
.A(n_1429),
.B(n_1402),
.Y(n_1448)
);

INVx1_ASAP7_75t_L g1449 ( 
.A(n_1414),
.Y(n_1449)
);

NAND2x1_ASAP7_75t_L g1450 ( 
.A(n_1412),
.B(n_1393),
.Y(n_1450)
);

NAND2xp5_ASAP7_75t_L g1451 ( 
.A(n_1416),
.B(n_1394),
.Y(n_1451)
);

HB1xp67_ASAP7_75t_L g1452 ( 
.A(n_1416),
.Y(n_1452)
);

INVx1_ASAP7_75t_L g1453 ( 
.A(n_1418),
.Y(n_1453)
);

AND2x2_ASAP7_75t_L g1454 ( 
.A(n_1426),
.B(n_1385),
.Y(n_1454)
);

INVx1_ASAP7_75t_L g1455 ( 
.A(n_1418),
.Y(n_1455)
);

INVx1_ASAP7_75t_L g1456 ( 
.A(n_1435),
.Y(n_1456)
);

AND2x2_ASAP7_75t_L g1457 ( 
.A(n_1426),
.B(n_1385),
.Y(n_1457)
);

NOR3x1_ASAP7_75t_L g1458 ( 
.A(n_1441),
.B(n_1421),
.C(n_1428),
.Y(n_1458)
);

INVx1_ASAP7_75t_L g1459 ( 
.A(n_1452),
.Y(n_1459)
);

AOI21xp33_ASAP7_75t_SL g1460 ( 
.A1(n_1438),
.A2(n_1427),
.B(n_1417),
.Y(n_1460)
);

NAND2xp5_ASAP7_75t_SL g1461 ( 
.A(n_1444),
.B(n_1420),
.Y(n_1461)
);

AOI221xp5_ASAP7_75t_L g1462 ( 
.A1(n_1439),
.A2(n_1419),
.B1(n_1417),
.B2(n_1432),
.C(n_1435),
.Y(n_1462)
);

OAI222xp33_ASAP7_75t_L g1463 ( 
.A1(n_1450),
.A2(n_1430),
.B1(n_1401),
.B2(n_1382),
.C1(n_1431),
.C2(n_1377),
.Y(n_1463)
);

AOI221xp5_ASAP7_75t_L g1464 ( 
.A1(n_1440),
.A2(n_1419),
.B1(n_1436),
.B2(n_1393),
.C(n_1394),
.Y(n_1464)
);

NOR2x1_ASAP7_75t_L g1465 ( 
.A(n_1447),
.B(n_1436),
.Y(n_1465)
);

O2A1O1Ixp33_ASAP7_75t_L g1466 ( 
.A1(n_1440),
.A2(n_1399),
.B(n_1403),
.C(n_1393),
.Y(n_1466)
);

OAI21xp5_ASAP7_75t_SL g1467 ( 
.A1(n_1445),
.A2(n_1382),
.B(n_1434),
.Y(n_1467)
);

NAND2xp5_ASAP7_75t_L g1468 ( 
.A(n_1444),
.B(n_1434),
.Y(n_1468)
);

OAI22xp5_ASAP7_75t_L g1469 ( 
.A1(n_1468),
.A2(n_1448),
.B1(n_1457),
.B2(n_1454),
.Y(n_1469)
);

INVx1_ASAP7_75t_L g1470 ( 
.A(n_1465),
.Y(n_1470)
);

NOR3xp33_ASAP7_75t_L g1471 ( 
.A(n_1461),
.B(n_1460),
.C(n_1466),
.Y(n_1471)
);

NAND2xp5_ASAP7_75t_L g1472 ( 
.A(n_1467),
.B(n_1442),
.Y(n_1472)
);

AOI21xp5_ASAP7_75t_L g1473 ( 
.A1(n_1464),
.A2(n_1451),
.B(n_1446),
.Y(n_1473)
);

OA22x2_ASAP7_75t_L g1474 ( 
.A1(n_1459),
.A2(n_1456),
.B1(n_1455),
.B2(n_1453),
.Y(n_1474)
);

NAND3xp33_ASAP7_75t_L g1475 ( 
.A(n_1462),
.B(n_1449),
.C(n_1446),
.Y(n_1475)
);

NOR2xp33_ASAP7_75t_L g1476 ( 
.A(n_1463),
.B(n_1443),
.Y(n_1476)
);

NAND4xp25_ASAP7_75t_L g1477 ( 
.A(n_1458),
.B(n_1443),
.C(n_1405),
.D(n_1433),
.Y(n_1477)
);

NAND3xp33_ASAP7_75t_L g1478 ( 
.A(n_1464),
.B(n_1405),
.C(n_1403),
.Y(n_1478)
);

NOR3xp33_ASAP7_75t_L g1479 ( 
.A(n_1471),
.B(n_1101),
.C(n_1057),
.Y(n_1479)
);

A2O1A1Ixp33_ASAP7_75t_L g1480 ( 
.A1(n_1473),
.A2(n_1399),
.B(n_1404),
.C(n_1389),
.Y(n_1480)
);

NAND3xp33_ASAP7_75t_L g1481 ( 
.A(n_1475),
.B(n_1476),
.C(n_1470),
.Y(n_1481)
);

OAI221xp5_ASAP7_75t_SL g1482 ( 
.A1(n_1478),
.A2(n_1377),
.B1(n_1389),
.B2(n_1404),
.C(n_1411),
.Y(n_1482)
);

OAI211xp5_ASAP7_75t_L g1483 ( 
.A1(n_1477),
.A2(n_1057),
.B(n_1405),
.C(n_1093),
.Y(n_1483)
);

NOR2x1_ASAP7_75t_L g1484 ( 
.A(n_1472),
.B(n_1022),
.Y(n_1484)
);

INVx1_ASAP7_75t_L g1485 ( 
.A(n_1480),
.Y(n_1485)
);

AOI22xp5_ASAP7_75t_L g1486 ( 
.A1(n_1481),
.A2(n_1469),
.B1(n_1474),
.B2(n_1400),
.Y(n_1486)
);

AOI22xp5_ASAP7_75t_L g1487 ( 
.A1(n_1479),
.A2(n_1483),
.B1(n_1484),
.B2(n_1383),
.Y(n_1487)
);

AND2x2_ASAP7_75t_L g1488 ( 
.A(n_1482),
.B(n_1411),
.Y(n_1488)
);

INVx1_ASAP7_75t_SL g1489 ( 
.A(n_1484),
.Y(n_1489)
);

CKINVDCx20_ASAP7_75t_R g1490 ( 
.A(n_1481),
.Y(n_1490)
);

NOR2x1_ASAP7_75t_L g1491 ( 
.A(n_1481),
.B(n_1038),
.Y(n_1491)
);

AND2x2_ASAP7_75t_L g1492 ( 
.A(n_1488),
.B(n_1383),
.Y(n_1492)
);

OAI22xp5_ASAP7_75t_L g1493 ( 
.A1(n_1490),
.A2(n_1486),
.B1(n_1487),
.B2(n_1485),
.Y(n_1493)
);

INVx1_ASAP7_75t_L g1494 ( 
.A(n_1491),
.Y(n_1494)
);

AOI22xp5_ASAP7_75t_L g1495 ( 
.A1(n_1489),
.A2(n_1400),
.B1(n_1100),
.B2(n_1065),
.Y(n_1495)
);

NOR2x1_ASAP7_75t_L g1496 ( 
.A(n_1490),
.B(n_1038),
.Y(n_1496)
);

NOR2xp33_ASAP7_75t_SL g1497 ( 
.A(n_1496),
.B(n_1100),
.Y(n_1497)
);

NAND2xp5_ASAP7_75t_L g1498 ( 
.A(n_1492),
.B(n_1290),
.Y(n_1498)
);

INVx3_ASAP7_75t_L g1499 ( 
.A(n_1494),
.Y(n_1499)
);

INVx1_ASAP7_75t_L g1500 ( 
.A(n_1499),
.Y(n_1500)
);

NOR2x2_ASAP7_75t_L g1501 ( 
.A(n_1500),
.B(n_1497),
.Y(n_1501)
);

NOR2xp33_ASAP7_75t_L g1502 ( 
.A(n_1501),
.B(n_1493),
.Y(n_1502)
);

INVx1_ASAP7_75t_L g1503 ( 
.A(n_1501),
.Y(n_1503)
);

INVx1_ASAP7_75t_L g1504 ( 
.A(n_1503),
.Y(n_1504)
);

OAI21xp33_ASAP7_75t_SL g1505 ( 
.A1(n_1502),
.A2(n_1495),
.B(n_1498),
.Y(n_1505)
);

AOI21xp5_ASAP7_75t_L g1506 ( 
.A1(n_1504),
.A2(n_1065),
.B(n_1045),
.Y(n_1506)
);

INVx2_ASAP7_75t_L g1507 ( 
.A(n_1505),
.Y(n_1507)
);

AOI22xp33_ASAP7_75t_L g1508 ( 
.A1(n_1507),
.A2(n_1290),
.B1(n_1277),
.B2(n_1278),
.Y(n_1508)
);

AOI322xp5_ASAP7_75t_L g1509 ( 
.A1(n_1508),
.A2(n_1506),
.A3(n_1290),
.B1(n_1313),
.B2(n_1323),
.C1(n_1322),
.C2(n_1278),
.Y(n_1509)
);

OAI221xp5_ASAP7_75t_R g1510 ( 
.A1(n_1509),
.A2(n_1290),
.B1(n_1051),
.B2(n_1098),
.C(n_1021),
.Y(n_1510)
);

AOI211xp5_ASAP7_75t_L g1511 ( 
.A1(n_1510),
.A2(n_1178),
.B(n_1262),
.C(n_1272),
.Y(n_1511)
);


endmodule