module fake_netlist_1_2729_n_40 (n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_40);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_40;
wire n_20;
wire n_38;
wire n_36;
wire n_37;
wire n_34;
wire n_28;
wire n_23;
wire n_31;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_30;
wire n_33;
wire n_18;
wire n_32;
wire n_35;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_27;
wire n_21;
wire n_29;
wire n_39;
CKINVDCx5p33_ASAP7_75t_R g11 ( .A(n_5), .Y(n_11) );
NAND2xp5_ASAP7_75t_SL g12 ( .A(n_9), .B(n_4), .Y(n_12) );
CKINVDCx20_ASAP7_75t_R g13 ( .A(n_4), .Y(n_13) );
CKINVDCx5p33_ASAP7_75t_R g14 ( .A(n_3), .Y(n_14) );
BUFx6f_ASAP7_75t_L g15 ( .A(n_7), .Y(n_15) );
AND2x4_ASAP7_75t_L g16 ( .A(n_2), .B(n_1), .Y(n_16) );
BUFx6f_ASAP7_75t_L g17 ( .A(n_10), .Y(n_17) );
BUFx2_ASAP7_75t_L g18 ( .A(n_11), .Y(n_18) );
NOR3xp33_ASAP7_75t_SL g19 ( .A(n_14), .B(n_0), .C(n_1), .Y(n_19) );
BUFx4f_ASAP7_75t_L g20 ( .A(n_16), .Y(n_20) );
INVx2_ASAP7_75t_L g21 ( .A(n_17), .Y(n_21) );
NOR3xp33_ASAP7_75t_SL g22 ( .A(n_12), .B(n_0), .C(n_2), .Y(n_22) );
AO31x2_ASAP7_75t_L g23 ( .A1(n_21), .A2(n_16), .A3(n_12), .B(n_3), .Y(n_23) );
INVx1_ASAP7_75t_L g24 ( .A(n_20), .Y(n_24) );
AND2x2_ASAP7_75t_L g25 ( .A(n_18), .B(n_13), .Y(n_25) );
INVx2_ASAP7_75t_L g26 ( .A(n_20), .Y(n_26) );
AOI22xp33_ASAP7_75t_L g27 ( .A1(n_26), .A2(n_15), .B1(n_17), .B2(n_19), .Y(n_27) );
AOI22xp5_ASAP7_75t_L g28 ( .A1(n_24), .A2(n_19), .B1(n_22), .B2(n_15), .Y(n_28) );
AND2x2_ASAP7_75t_L g29 ( .A(n_25), .B(n_5), .Y(n_29) );
INVx1_ASAP7_75t_L g30 ( .A(n_29), .Y(n_30) );
OR2x2_ASAP7_75t_L g31 ( .A(n_28), .B(n_23), .Y(n_31) );
CKINVDCx5p33_ASAP7_75t_R g32 ( .A(n_30), .Y(n_32) );
O2A1O1Ixp33_ASAP7_75t_SL g33 ( .A1(n_31), .A2(n_26), .B(n_23), .C(n_27), .Y(n_33) );
OAI21x1_ASAP7_75t_SL g34 ( .A1(n_33), .A2(n_23), .B(n_8), .Y(n_34) );
AOI22xp5_ASAP7_75t_L g35 ( .A1(n_32), .A2(n_15), .B1(n_17), .B2(n_23), .Y(n_35) );
OA21x2_ASAP7_75t_L g36 ( .A1(n_33), .A2(n_15), .B(n_17), .Y(n_36) );
CKINVDCx5p33_ASAP7_75t_R g37 ( .A(n_35), .Y(n_37) );
NAND2xp5_ASAP7_75t_L g38 ( .A(n_34), .B(n_6), .Y(n_38) );
INVx2_ASAP7_75t_SL g39 ( .A(n_37), .Y(n_39) );
AOI22xp33_ASAP7_75t_L g40 ( .A1(n_39), .A2(n_36), .B1(n_38), .B2(n_37), .Y(n_40) );
endmodule