module fake_jpeg_3681_n_208 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_208);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_208;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_207;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_202;
wire n_75;
wire n_122;
wire n_102;
wire n_121;
wire n_130;
wire n_99;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g51 ( 
.A(n_50),
.Y(n_51)
);

BUFx5_ASAP7_75t_L g52 ( 
.A(n_33),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_46),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_16),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_45),
.Y(n_55)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_2),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_26),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_29),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_35),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_3),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_1),
.Y(n_61)
);

BUFx16f_ASAP7_75t_L g62 ( 
.A(n_28),
.Y(n_62)
);

BUFx5_ASAP7_75t_L g63 ( 
.A(n_10),
.Y(n_63)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_18),
.Y(n_64)
);

BUFx12f_ASAP7_75t_L g65 ( 
.A(n_49),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_27),
.Y(n_66)
);

INVx11_ASAP7_75t_SL g67 ( 
.A(n_22),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_15),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_36),
.Y(n_69)
);

BUFx4f_ASAP7_75t_SL g70 ( 
.A(n_30),
.Y(n_70)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_19),
.Y(n_71)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_20),
.Y(n_72)
);

BUFx8_ASAP7_75t_L g73 ( 
.A(n_4),
.Y(n_73)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_12),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_59),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_75),
.Y(n_86)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_74),
.Y(n_76)
);

INVx2_ASAP7_75t_SL g82 ( 
.A(n_76),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_54),
.B(n_0),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_77),
.B(n_70),
.Y(n_85)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_51),
.Y(n_78)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_78),
.Y(n_87)
);

BUFx12_ASAP7_75t_L g79 ( 
.A(n_62),
.Y(n_79)
);

BUFx3_ASAP7_75t_L g84 ( 
.A(n_79),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_67),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_80),
.B(n_73),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_59),
.Y(n_81)
);

INVx5_ASAP7_75t_L g93 ( 
.A(n_81),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_76),
.B(n_53),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_83),
.B(n_88),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_85),
.B(n_89),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_75),
.A2(n_69),
.B1(n_56),
.B2(n_71),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_80),
.A2(n_73),
.B1(n_61),
.B2(n_60),
.Y(n_90)
);

INVx1_ASAP7_75t_SL g97 ( 
.A(n_90),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_78),
.B(n_58),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_91),
.B(n_79),
.C(n_65),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_81),
.B(n_66),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_92),
.B(n_94),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_79),
.B(n_55),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_L g95 ( 
.A1(n_82),
.A2(n_70),
.B1(n_67),
.B2(n_69),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_95),
.A2(n_102),
.B1(n_63),
.B2(n_2),
.Y(n_124)
);

INVx13_ASAP7_75t_L g96 ( 
.A(n_84),
.Y(n_96)
);

INVx13_ASAP7_75t_L g114 ( 
.A(n_96),
.Y(n_114)
);

BUFx12f_ASAP7_75t_L g98 ( 
.A(n_87),
.Y(n_98)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_98),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_83),
.B(n_60),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_SL g128 ( 
.A1(n_100),
.A2(n_107),
.B(n_108),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_L g102 ( 
.A1(n_82),
.A2(n_68),
.B1(n_57),
.B2(n_62),
.Y(n_102)
);

INVx8_ASAP7_75t_L g103 ( 
.A(n_86),
.Y(n_103)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_103),
.Y(n_113)
);

INVx5_ASAP7_75t_L g105 ( 
.A(n_84),
.Y(n_105)
);

HB1xp67_ASAP7_75t_L g119 ( 
.A(n_105),
.Y(n_119)
);

OR2x2_ASAP7_75t_L g106 ( 
.A(n_87),
.B(n_79),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_106),
.B(n_65),
.Y(n_118)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_91),
.B(n_60),
.Y(n_107)
);

NOR4xp25_ASAP7_75t_SL g108 ( 
.A(n_88),
.B(n_25),
.C(n_48),
.D(n_47),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_93),
.B(n_72),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_109),
.B(n_111),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_110),
.B(n_64),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_93),
.B(n_65),
.Y(n_111)
);

INVx13_ASAP7_75t_L g112 ( 
.A(n_86),
.Y(n_112)
);

INVx13_ASAP7_75t_L g126 ( 
.A(n_112),
.Y(n_126)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_98),
.Y(n_115)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_115),
.Y(n_135)
);

INVx6_ASAP7_75t_SL g117 ( 
.A(n_96),
.Y(n_117)
);

CKINVDCx14_ASAP7_75t_R g149 ( 
.A(n_117),
.Y(n_149)
);

OR2x2_ASAP7_75t_L g145 ( 
.A(n_118),
.B(n_6),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_100),
.B(n_52),
.C(n_64),
.Y(n_120)
);

XOR2xp5_ASAP7_75t_L g143 ( 
.A(n_120),
.B(n_130),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_121),
.B(n_97),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_99),
.B(n_0),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_123),
.B(n_124),
.Y(n_134)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_102),
.Y(n_125)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_125),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_101),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_127),
.A2(n_130),
.B1(n_7),
.B2(n_8),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_104),
.B(n_5),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_129),
.B(n_131),
.Y(n_142)
);

AO21x2_ASAP7_75t_L g130 ( 
.A1(n_95),
.A2(n_23),
.B(n_43),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_107),
.B(n_5),
.Y(n_131)
);

INVx13_ASAP7_75t_L g132 ( 
.A(n_106),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_132),
.Y(n_154)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_103),
.Y(n_133)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_133),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g162 ( 
.A(n_137),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_128),
.B(n_98),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_138),
.B(n_139),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_116),
.B(n_31),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_132),
.A2(n_97),
.B1(n_112),
.B2(n_24),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_141),
.A2(n_151),
.B1(n_155),
.B2(n_11),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_143),
.B(n_32),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_119),
.B(n_6),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_144),
.B(n_146),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_SL g156 ( 
.A1(n_145),
.A2(n_147),
.B(n_114),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_113),
.B(n_44),
.Y(n_146)
);

OR2x2_ASAP7_75t_L g147 ( 
.A(n_120),
.B(n_7),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_119),
.Y(n_148)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_148),
.Y(n_160)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_122),
.Y(n_150)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_150),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_122),
.Y(n_152)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_152),
.Y(n_165)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_130),
.Y(n_153)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_153),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_130),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_156),
.B(n_166),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_L g157 ( 
.A1(n_154),
.A2(n_114),
.B(n_126),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_157),
.A2(n_163),
.B1(n_145),
.B2(n_134),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_138),
.B(n_143),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_158),
.B(n_159),
.C(n_168),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_140),
.B(n_126),
.Y(n_159)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_161),
.B(n_146),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_136),
.A2(n_9),
.B1(n_11),
.B2(n_12),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_149),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_147),
.B(n_37),
.C(n_41),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_170),
.B(n_171),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_139),
.B(n_13),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_135),
.Y(n_172)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_172),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_174),
.B(n_162),
.C(n_169),
.Y(n_187)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_164),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_177),
.B(n_178),
.Y(n_185)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_160),
.Y(n_178)
);

CKINVDCx16_ASAP7_75t_R g180 ( 
.A(n_173),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_180),
.B(n_181),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_158),
.A2(n_141),
.B1(n_152),
.B2(n_142),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_182),
.B(n_184),
.Y(n_189)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_165),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_175),
.B(n_162),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_L g197 ( 
.A1(n_186),
.A2(n_191),
.B(n_185),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_187),
.B(n_190),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_183),
.B(n_168),
.C(n_159),
.Y(n_190)
);

AOI21xp5_ASAP7_75t_L g191 ( 
.A1(n_176),
.A2(n_167),
.B(n_14),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_179),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_192),
.B(n_13),
.Y(n_196)
);

AOI22xp33_ASAP7_75t_SL g193 ( 
.A1(n_186),
.A2(n_182),
.B1(n_183),
.B2(n_174),
.Y(n_193)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_193),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_188),
.B(n_38),
.Y(n_195)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_195),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_196),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_L g201 ( 
.A1(n_198),
.A2(n_193),
.B(n_194),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_SL g202 ( 
.A(n_201),
.B(n_189),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_202),
.A2(n_197),
.B1(n_199),
.B2(n_200),
.Y(n_203)
);

OAI22xp33_ASAP7_75t_SL g204 ( 
.A1(n_203),
.A2(n_17),
.B1(n_21),
.B2(n_34),
.Y(n_204)
);

INVxp67_ASAP7_75t_L g205 ( 
.A(n_204),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_205),
.B(n_39),
.C(n_40),
.Y(n_206)
);

BUFx24_ASAP7_75t_SL g207 ( 
.A(n_206),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_207),
.B(n_42),
.Y(n_208)
);


endmodule