module fake_jpeg_3436_n_171 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_171);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_171;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g42 ( 
.A(n_1),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_37),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_39),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_22),
.Y(n_45)
);

INVx11_ASAP7_75t_L g46 ( 
.A(n_30),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_9),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_11),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_31),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_12),
.Y(n_50)
);

BUFx5_ASAP7_75t_L g51 ( 
.A(n_18),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_19),
.Y(n_52)
);

INVx11_ASAP7_75t_SL g53 ( 
.A(n_20),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_26),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_8),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_33),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_3),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_4),
.Y(n_58)
);

INVx11_ASAP7_75t_L g59 ( 
.A(n_53),
.Y(n_59)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_59),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_47),
.B(n_0),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_60),
.B(n_49),
.Y(n_77)
);

AOI21xp33_ASAP7_75t_L g61 ( 
.A1(n_43),
.A2(n_16),
.B(n_40),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_61),
.B(n_45),
.Y(n_69)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_44),
.Y(n_62)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_62),
.Y(n_67)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_53),
.Y(n_63)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_63),
.Y(n_70)
);

BUFx6f_ASAP7_75t_SL g64 ( 
.A(n_43),
.Y(n_64)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_64),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_56),
.Y(n_65)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_65),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_69),
.B(n_45),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_61),
.B(n_52),
.Y(n_72)
);

XOR2xp5_ASAP7_75t_SL g82 ( 
.A(n_72),
.B(n_57),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_60),
.B(n_58),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_73),
.B(n_74),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_62),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_63),
.B(n_55),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_75),
.B(n_77),
.Y(n_89)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_59),
.Y(n_76)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_76),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_79),
.B(n_82),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_74),
.B(n_42),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_80),
.B(n_83),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_72),
.B(n_67),
.Y(n_83)
);

OA22x2_ASAP7_75t_L g84 ( 
.A1(n_69),
.A2(n_65),
.B1(n_57),
.B2(n_50),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_84),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_67),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_85),
.B(n_1),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_70),
.B(n_54),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_86),
.B(n_0),
.Y(n_103)
);

BUFx12f_ASAP7_75t_L g87 ( 
.A(n_70),
.Y(n_87)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_87),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_71),
.A2(n_65),
.B1(n_50),
.B2(n_56),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_88),
.A2(n_46),
.B1(n_51),
.B2(n_21),
.Y(n_108)
);

HB1xp67_ASAP7_75t_L g90 ( 
.A(n_66),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_90),
.Y(n_104)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_71),
.Y(n_91)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_91),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_SL g92 ( 
.A1(n_68),
.A2(n_48),
.B(n_64),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_SL g111 ( 
.A1(n_92),
.A2(n_2),
.B(n_5),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_68),
.B(n_65),
.C(n_64),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_93),
.B(n_17),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_84),
.A2(n_48),
.B1(n_66),
.B2(n_76),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_95),
.A2(n_98),
.B1(n_108),
.B2(n_110),
.Y(n_115)
);

OAI21xp33_ASAP7_75t_L g96 ( 
.A1(n_82),
.A2(n_84),
.B(n_81),
.Y(n_96)
);

CKINVDCx14_ASAP7_75t_R g128 ( 
.A(n_96),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_L g97 ( 
.A1(n_78),
.A2(n_63),
.B(n_59),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g112 ( 
.A(n_97),
.B(n_109),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_88),
.A2(n_63),
.B1(n_46),
.B2(n_51),
.Y(n_98)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_78),
.Y(n_102)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_102),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_103),
.B(n_32),
.Y(n_130)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_93),
.Y(n_106)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_106),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_107),
.B(n_5),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_89),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_111),
.Y(n_121)
);

OAI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_94),
.A2(n_96),
.B1(n_99),
.B2(n_95),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_116),
.A2(n_127),
.B1(n_13),
.B2(n_14),
.Y(n_144)
);

AO22x1_ASAP7_75t_SL g117 ( 
.A1(n_94),
.A2(n_87),
.B1(n_24),
.B2(n_25),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_117),
.B(n_120),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_100),
.B(n_87),
.C(n_23),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_118),
.B(n_119),
.C(n_29),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_101),
.B(n_15),
.C(n_38),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_104),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_122),
.B(n_125),
.Y(n_135)
);

INVx2_ASAP7_75t_SL g123 ( 
.A(n_105),
.Y(n_123)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_123),
.Y(n_133)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_104),
.Y(n_124)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_124),
.Y(n_140)
);

CKINVDCx16_ASAP7_75t_R g125 ( 
.A(n_97),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_98),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_126),
.A2(n_129),
.B1(n_13),
.B2(n_14),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_94),
.A2(n_6),
.B1(n_7),
.B2(n_9),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_94),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_130),
.B(n_131),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_100),
.B(n_10),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_SL g132 ( 
.A1(n_121),
.A2(n_34),
.B(n_36),
.Y(n_132)
);

AOI21xp5_ASAP7_75t_L g153 ( 
.A1(n_132),
.A2(n_121),
.B(n_41),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_113),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_134),
.Y(n_154)
);

INVxp67_ASAP7_75t_L g136 ( 
.A(n_112),
.Y(n_136)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_136),
.Y(n_148)
);

INVx1_ASAP7_75t_SL g151 ( 
.A(n_137),
.Y(n_151)
);

XNOR2x1_ASAP7_75t_L g138 ( 
.A(n_114),
.B(n_27),
.Y(n_138)
);

XOR2xp5_ASAP7_75t_L g155 ( 
.A(n_138),
.B(n_139),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_128),
.B(n_28),
.C(n_35),
.Y(n_139)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_141),
.Y(n_149)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_112),
.Y(n_143)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_143),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_L g152 ( 
.A1(n_144),
.A2(n_145),
.B(n_146),
.Y(n_152)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_123),
.Y(n_145)
);

CKINVDCx16_ASAP7_75t_R g146 ( 
.A(n_118),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_L g159 ( 
.A1(n_153),
.A2(n_137),
.B(n_139),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_148),
.A2(n_142),
.B1(n_150),
.B2(n_116),
.Y(n_156)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_156),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_149),
.A2(n_135),
.B1(n_115),
.B2(n_143),
.Y(n_157)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_157),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_154),
.B(n_147),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_158),
.B(n_159),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_151),
.B(n_136),
.C(n_140),
.Y(n_160)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_161),
.B(n_160),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_SL g166 ( 
.A1(n_164),
.A2(n_165),
.B(n_163),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_162),
.B(n_151),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_166),
.B(n_160),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_167),
.A2(n_152),
.B1(n_133),
.B2(n_155),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g169 ( 
.A(n_168),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_169),
.B(n_138),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_170),
.B(n_155),
.Y(n_171)
);


endmodule