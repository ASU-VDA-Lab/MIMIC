module fake_jpeg_16167_n_64 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_64);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_64;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_23;
wire n_10;
wire n_27;
wire n_55;
wire n_22;
wire n_51;
wire n_47;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_59;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_62;
wire n_17;
wire n_31;
wire n_25;
wire n_56;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;

NAND2xp5_ASAP7_75t_L g8 ( 
.A(n_4),
.B(n_6),
.Y(n_8)
);

BUFx6f_ASAP7_75t_L g9 ( 
.A(n_1),
.Y(n_9)
);

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_1),
.Y(n_10)
);

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_1),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_4),
.Y(n_12)
);

NOR2xp33_ASAP7_75t_L g13 ( 
.A(n_6),
.B(n_4),
.Y(n_13)
);

BUFx4f_ASAP7_75t_L g14 ( 
.A(n_0),
.Y(n_14)
);

INVx4_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_2),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_18),
.B(n_20),
.Y(n_27)
);

AOI22xp33_ASAP7_75t_SL g19 ( 
.A1(n_15),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_19)
);

OR2x2_ASAP7_75t_L g25 ( 
.A(n_19),
.B(n_23),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

AOI21xp5_ASAP7_75t_L g21 ( 
.A1(n_14),
.A2(n_2),
.B(n_3),
.Y(n_21)
);

OAI21xp5_ASAP7_75t_SL g28 ( 
.A1(n_21),
.A2(n_22),
.B(n_14),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_14),
.A2(n_3),
.B1(n_5),
.B2(n_7),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_21),
.B(n_8),
.Y(n_24)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_24),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_22),
.B(n_8),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_26),
.B(n_12),
.Y(n_34)
);

AOI22xp5_ASAP7_75t_L g40 ( 
.A1(n_28),
.A2(n_10),
.B1(n_11),
.B2(n_16),
.Y(n_40)
);

INVx5_ASAP7_75t_L g29 ( 
.A(n_20),
.Y(n_29)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_29),
.Y(n_33)
);

INVx5_ASAP7_75t_L g30 ( 
.A(n_18),
.Y(n_30)
);

INVxp67_ASAP7_75t_L g36 ( 
.A(n_30),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_SL g31 ( 
.A1(n_26),
.A2(n_15),
.B1(n_17),
.B2(n_11),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_31),
.B(n_38),
.Y(n_45)
);

AND2x2_ASAP7_75t_L g46 ( 
.A(n_34),
.B(n_35),
.Y(n_46)
);

MAJIxp5_ASAP7_75t_L g35 ( 
.A(n_28),
.B(n_17),
.C(n_12),
.Y(n_35)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_27),
.Y(n_37)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_37),
.Y(n_47)
);

BUFx12_ASAP7_75t_L g38 ( 
.A(n_30),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_SL g39 ( 
.A(n_25),
.B(n_13),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_SL g43 ( 
.A(n_39),
.B(n_10),
.Y(n_43)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_40),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_33),
.Y(n_42)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_42),
.Y(n_48)
);

OAI21xp5_ASAP7_75t_SL g49 ( 
.A1(n_43),
.A2(n_44),
.B(n_34),
.Y(n_49)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

XOR2xp5_ASAP7_75t_L g53 ( 
.A(n_49),
.B(n_51),
.Y(n_53)
);

XNOR2xp5_ASAP7_75t_SL g50 ( 
.A(n_46),
.B(n_35),
.Y(n_50)
);

XNOR2xp5_ASAP7_75t_SL g54 ( 
.A(n_50),
.B(n_52),
.Y(n_54)
);

XOR2xp5_ASAP7_75t_L g51 ( 
.A(n_46),
.B(n_45),
.Y(n_51)
);

OAI21xp5_ASAP7_75t_SL g52 ( 
.A1(n_46),
.A2(n_32),
.B(n_40),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g55 ( 
.A1(n_48),
.A2(n_41),
.B1(n_47),
.B2(n_25),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_55),
.A2(n_41),
.B1(n_31),
.B2(n_25),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g56 ( 
.A(n_54),
.B(n_53),
.C(n_50),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_56),
.B(n_57),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_56),
.A2(n_44),
.B1(n_29),
.B2(n_16),
.Y(n_58)
);

OAI21xp5_ASAP7_75t_SL g60 ( 
.A1(n_58),
.A2(n_36),
.B(n_27),
.Y(n_60)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_60),
.B(n_61),
.C(n_54),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_59),
.B(n_38),
.Y(n_61)
);

MAJx2_ASAP7_75t_L g63 ( 
.A(n_62),
.B(n_7),
.C(n_36),
.Y(n_63)
);

XNOR2xp5_ASAP7_75t_L g64 ( 
.A(n_63),
.B(n_38),
.Y(n_64)
);


endmodule