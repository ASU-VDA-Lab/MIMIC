module fake_jpeg_14119_n_343 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_343);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_343;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

BUFx16f_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

INVx1_ASAP7_75t_SL g19 ( 
.A(n_10),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_6),
.Y(n_20)
);

BUFx4f_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_5),
.Y(n_22)
);

INVx11_ASAP7_75t_SL g23 ( 
.A(n_15),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_5),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_1),
.Y(n_26)
);

BUFx12_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

BUFx12_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

INVx1_ASAP7_75t_SL g29 ( 
.A(n_7),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_15),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_11),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_5),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_9),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g36 ( 
.A(n_19),
.B(n_0),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_36),
.B(n_39),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_35),
.Y(n_37)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_21),
.Y(n_38)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g39 ( 
.A(n_19),
.B(n_0),
.Y(n_39)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_17),
.Y(n_40)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_40),
.Y(n_66)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_16),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_41),
.Y(n_73)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_21),
.Y(n_42)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_42),
.Y(n_55)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_30),
.Y(n_43)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_43),
.Y(n_63)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_17),
.Y(n_44)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_44),
.Y(n_72)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_18),
.Y(n_45)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_45),
.Y(n_52)
);

INVx2_ASAP7_75t_SL g46 ( 
.A(n_30),
.Y(n_46)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_46),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_16),
.Y(n_47)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_47),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_16),
.Y(n_48)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_48),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_36),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_51),
.B(n_67),
.Y(n_98)
);

OAI22xp33_ASAP7_75t_L g54 ( 
.A1(n_45),
.A2(n_26),
.B1(n_25),
.B2(n_22),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_54),
.A2(n_59),
.B1(n_61),
.B2(n_23),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_39),
.B(n_46),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_58),
.B(n_70),
.Y(n_76)
);

OAI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_47),
.A2(n_24),
.B1(n_19),
.B2(n_29),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_46),
.A2(n_29),
.B1(n_18),
.B2(n_33),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_60),
.A2(n_25),
.B1(n_26),
.B2(n_30),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_47),
.A2(n_24),
.B1(n_16),
.B2(n_29),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_37),
.B(n_20),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_SL g82 ( 
.A(n_62),
.B(n_65),
.Y(n_82)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_40),
.Y(n_64)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_64),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_37),
.B(n_20),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_37),
.B(n_20),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_L g68 ( 
.A1(n_47),
.A2(n_24),
.B1(n_22),
.B2(n_26),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_68),
.A2(n_46),
.B1(n_22),
.B2(n_25),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_37),
.B(n_32),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_40),
.Y(n_71)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_71),
.Y(n_93)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_53),
.Y(n_74)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_74),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_75),
.A2(n_57),
.B1(n_69),
.B2(n_48),
.Y(n_108)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_66),
.Y(n_77)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_77),
.Y(n_110)
);

INVx5_ASAP7_75t_L g78 ( 
.A(n_50),
.Y(n_78)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_78),
.Y(n_114)
);

AO22x2_ASAP7_75t_L g79 ( 
.A1(n_56),
.A2(n_43),
.B1(n_44),
.B2(n_48),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g123 ( 
.A(n_79),
.B(n_97),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_51),
.B(n_58),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_80),
.B(n_94),
.Y(n_119)
);

AOI21xp5_ASAP7_75t_L g118 ( 
.A1(n_81),
.A2(n_85),
.B(n_92),
.Y(n_118)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_53),
.Y(n_83)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_83),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_L g85 ( 
.A1(n_49),
.A2(n_33),
.B(n_18),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_56),
.B(n_44),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_86),
.B(n_38),
.C(n_73),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_70),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_87),
.B(n_96),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_73),
.Y(n_88)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_88),
.Y(n_133)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_55),
.Y(n_89)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_89),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_61),
.A2(n_33),
.B1(n_30),
.B2(n_41),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_90),
.A2(n_97),
.B1(n_102),
.B2(n_92),
.Y(n_131)
);

A2O1A1Ixp33_ASAP7_75t_L g91 ( 
.A1(n_49),
.A2(n_31),
.B(n_32),
.C(n_17),
.Y(n_91)
);

O2A1O1Ixp33_ASAP7_75t_L g109 ( 
.A1(n_91),
.A2(n_34),
.B(n_17),
.C(n_21),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_52),
.A2(n_23),
.B1(n_31),
.B2(n_43),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_52),
.B(n_42),
.Y(n_94)
);

BUFx3_ASAP7_75t_L g95 ( 
.A(n_66),
.Y(n_95)
);

BUFx24_ASAP7_75t_L g117 ( 
.A(n_95),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_62),
.Y(n_96)
);

AOI32xp33_ASAP7_75t_L g99 ( 
.A1(n_65),
.A2(n_30),
.A3(n_34),
.B1(n_21),
.B2(n_17),
.Y(n_99)
);

XOR2xp5_ASAP7_75t_L g122 ( 
.A(n_99),
.B(n_35),
.Y(n_122)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_72),
.Y(n_100)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_100),
.Y(n_124)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_64),
.Y(n_101)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_101),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_57),
.A2(n_48),
.B1(n_41),
.B2(n_42),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_102),
.A2(n_69),
.B1(n_30),
.B2(n_21),
.Y(n_130)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_55),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_103),
.B(n_105),
.Y(n_120)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_72),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_104),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_67),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_82),
.A2(n_50),
.B1(n_71),
.B2(n_63),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_SL g154 ( 
.A1(n_107),
.A2(n_89),
.B(n_83),
.Y(n_154)
);

OA22x2_ASAP7_75t_L g156 ( 
.A1(n_108),
.A2(n_88),
.B1(n_78),
.B2(n_28),
.Y(n_156)
);

AND2x2_ASAP7_75t_L g149 ( 
.A(n_109),
.B(n_113),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_86),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_116),
.B(n_127),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_98),
.B(n_63),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_121),
.B(n_129),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_122),
.A2(n_131),
.B1(n_132),
.B2(n_79),
.Y(n_141)
);

O2A1O1Ixp33_ASAP7_75t_L g125 ( 
.A1(n_91),
.A2(n_63),
.B(n_73),
.C(n_69),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_L g152 ( 
.A1(n_125),
.A2(n_104),
.B(n_100),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_80),
.B(n_38),
.C(n_24),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_126),
.B(n_93),
.C(n_84),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_86),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_76),
.B(n_10),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_L g161 ( 
.A1(n_130),
.A2(n_28),
.B1(n_27),
.B2(n_2),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_76),
.A2(n_35),
.B1(n_27),
.B2(n_28),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_L g136 ( 
.A(n_119),
.B(n_85),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_136),
.B(n_145),
.C(n_114),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_119),
.A2(n_94),
.B1(n_75),
.B2(n_79),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_137),
.A2(n_160),
.B1(n_110),
.B2(n_114),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_SL g139 ( 
.A(n_106),
.B(n_84),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g188 ( 
.A(n_139),
.B(n_150),
.Y(n_188)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_140),
.B(n_28),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_SL g169 ( 
.A1(n_141),
.A2(n_158),
.B(n_117),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_120),
.B(n_93),
.Y(n_142)
);

CKINVDCx14_ASAP7_75t_R g183 ( 
.A(n_142),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_126),
.B(n_116),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_143),
.B(n_146),
.Y(n_173)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_128),
.Y(n_144)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_144),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_122),
.B(n_74),
.C(n_103),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_127),
.B(n_79),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_128),
.Y(n_147)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_147),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_123),
.A2(n_125),
.B1(n_109),
.B2(n_132),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_148),
.A2(n_157),
.B1(n_161),
.B2(n_2),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_124),
.B(n_95),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_113),
.B(n_107),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_151),
.B(n_156),
.Y(n_174)
);

CKINVDCx16_ASAP7_75t_R g176 ( 
.A(n_152),
.Y(n_176)
);

CKINVDCx16_ASAP7_75t_R g153 ( 
.A(n_118),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_153),
.B(n_155),
.Y(n_175)
);

INVxp67_ASAP7_75t_L g185 ( 
.A(n_154),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_118),
.B(n_77),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_123),
.A2(n_27),
.B1(n_28),
.B2(n_8),
.Y(n_157)
);

OAI21xp33_ASAP7_75t_SL g158 ( 
.A1(n_123),
.A2(n_27),
.B(n_7),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_117),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_159),
.B(n_110),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_108),
.A2(n_130),
.B1(n_111),
.B2(n_133),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_111),
.B(n_0),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_162),
.B(n_165),
.Y(n_177)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_112),
.Y(n_163)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_163),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_124),
.B(n_9),
.Y(n_164)
);

INVxp67_ASAP7_75t_L g193 ( 
.A(n_164),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_112),
.B(n_134),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_115),
.Y(n_166)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_166),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_141),
.A2(n_133),
.B1(n_134),
.B2(n_115),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_167),
.B(n_179),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_SL g207 ( 
.A(n_168),
.B(n_196),
.Y(n_207)
);

INVxp67_ASAP7_75t_L g212 ( 
.A(n_169),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_171),
.A2(n_148),
.B1(n_195),
.B2(n_180),
.Y(n_211)
);

CKINVDCx14_ASAP7_75t_R g202 ( 
.A(n_172),
.Y(n_202)
);

AOI22xp33_ASAP7_75t_L g178 ( 
.A1(n_137),
.A2(n_117),
.B1(n_27),
.B2(n_9),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_178),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_136),
.B(n_117),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_139),
.B(n_7),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_SL g206 ( 
.A(n_181),
.B(n_192),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_140),
.B(n_1),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_182),
.B(n_186),
.Y(n_222)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_163),
.Y(n_184)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_184),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_138),
.B(n_6),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_143),
.B(n_6),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_187),
.B(n_190),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_162),
.B(n_1),
.Y(n_189)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_189),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_146),
.B(n_12),
.Y(n_190)
);

AOI22xp33_ASAP7_75t_SL g191 ( 
.A1(n_155),
.A2(n_12),
.B1(n_14),
.B2(n_13),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_L g213 ( 
.A1(n_191),
.A2(n_154),
.B(n_135),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_135),
.B(n_12),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_194),
.B(n_201),
.C(n_151),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_149),
.B(n_13),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_149),
.B(n_13),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_SL g230 ( 
.A(n_198),
.B(n_14),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_149),
.B(n_1),
.Y(n_199)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_199),
.Y(n_225)
);

AND2x2_ASAP7_75t_L g204 ( 
.A(n_200),
.B(n_156),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_145),
.B(n_14),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_203),
.B(n_230),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_204),
.B(n_171),
.Y(n_237)
);

HAxp5_ASAP7_75t_SL g205 ( 
.A(n_176),
.B(n_153),
.CON(n_205),
.SN(n_205)
);

AOI21xp5_ASAP7_75t_L g231 ( 
.A1(n_205),
.A2(n_215),
.B(n_220),
.Y(n_231)
);

HB1xp67_ASAP7_75t_L g208 ( 
.A(n_173),
.Y(n_208)
);

HB1xp67_ASAP7_75t_L g235 ( 
.A(n_208),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_173),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_210),
.B(n_214),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_211),
.A2(n_167),
.B1(n_176),
.B2(n_174),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_L g245 ( 
.A1(n_213),
.A2(n_227),
.B(n_198),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_177),
.Y(n_214)
);

AOI21xp5_ASAP7_75t_L g215 ( 
.A1(n_175),
.A2(n_152),
.B(n_159),
.Y(n_215)
);

NAND3xp33_ASAP7_75t_L g217 ( 
.A(n_183),
.B(n_147),
.C(n_144),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_217),
.B(n_219),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_177),
.Y(n_219)
);

AOI21xp5_ASAP7_75t_L g220 ( 
.A1(n_175),
.A2(n_160),
.B(n_157),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_168),
.B(n_165),
.C(n_166),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_223),
.B(n_226),
.C(n_201),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_186),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_224),
.B(n_188),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_194),
.B(n_156),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_L g227 ( 
.A1(n_185),
.A2(n_156),
.B(n_3),
.Y(n_227)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_180),
.Y(n_229)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_229),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_207),
.B(n_179),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_232),
.B(n_207),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_233),
.B(n_234),
.C(n_255),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_223),
.B(n_182),
.C(n_174),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g266 ( 
.A1(n_236),
.A2(n_245),
.B1(n_220),
.B2(n_213),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_237),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_221),
.B(n_190),
.Y(n_238)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_238),
.Y(n_264)
);

OA21x2_ASAP7_75t_L g239 ( 
.A1(n_212),
.A2(n_199),
.B(n_169),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_SL g262 ( 
.A1(n_239),
.A2(n_254),
.B(n_215),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_221),
.B(n_187),
.Y(n_240)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_240),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_202),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_241),
.B(n_246),
.Y(n_257)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_243),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_211),
.B(n_195),
.Y(n_244)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_244),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_229),
.B(n_216),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_216),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_248),
.B(n_238),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_206),
.B(n_188),
.Y(n_250)
);

NAND3xp33_ASAP7_75t_L g271 ( 
.A(n_250),
.B(n_256),
.C(n_209),
.Y(n_271)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_228),
.Y(n_251)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_251),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_228),
.B(n_189),
.Y(n_253)
);

CKINVDCx16_ASAP7_75t_R g270 ( 
.A(n_253),
.Y(n_270)
);

OAI21xp5_ASAP7_75t_L g254 ( 
.A1(n_212),
.A2(n_196),
.B(n_197),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_203),
.B(n_197),
.C(n_184),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_224),
.B(n_193),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_SL g289 ( 
.A(n_258),
.B(n_260),
.Y(n_289)
);

XNOR2x1_ASAP7_75t_L g260 ( 
.A(n_239),
.B(n_226),
.Y(n_260)
);

INVxp67_ASAP7_75t_SL g261 ( 
.A(n_243),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_261),
.B(n_271),
.Y(n_294)
);

NAND3xp33_ASAP7_75t_SL g286 ( 
.A(n_262),
.B(n_268),
.C(n_246),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_244),
.A2(n_204),
.B1(n_227),
.B2(n_200),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_265),
.A2(n_236),
.B1(n_237),
.B2(n_231),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_266),
.A2(n_239),
.B1(n_245),
.B2(n_248),
.Y(n_283)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_233),
.B(n_232),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_269),
.B(n_252),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_255),
.B(n_225),
.C(n_222),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_272),
.B(n_235),
.C(n_231),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_241),
.B(n_222),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_SL g291 ( 
.A(n_275),
.B(n_242),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_234),
.B(n_225),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_277),
.B(n_252),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_272),
.B(n_249),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_278),
.B(n_284),
.Y(n_298)
);

XNOR2x1_ASAP7_75t_L g297 ( 
.A(n_279),
.B(n_260),
.Y(n_297)
);

XOR2xp5_ASAP7_75t_L g303 ( 
.A(n_280),
.B(n_292),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_281),
.B(n_263),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_274),
.Y(n_282)
);

AOI21xp5_ASAP7_75t_L g306 ( 
.A1(n_282),
.A2(n_253),
.B(n_242),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_283),
.A2(n_293),
.B1(n_265),
.B2(n_290),
.Y(n_295)
);

CKINVDCx16_ASAP7_75t_R g284 ( 
.A(n_257),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_285),
.B(n_287),
.Y(n_309)
);

OAI21xp5_ASAP7_75t_SL g304 ( 
.A1(n_286),
.A2(n_293),
.B(n_267),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_264),
.A2(n_247),
.B1(n_218),
.B2(n_240),
.Y(n_287)
);

BUFx24_ASAP7_75t_SL g288 ( 
.A(n_277),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_288),
.B(n_263),
.Y(n_296)
);

INVx11_ASAP7_75t_L g290 ( 
.A(n_257),
.Y(n_290)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_290),
.Y(n_301)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_291),
.Y(n_308)
);

XOR2xp5_ASAP7_75t_L g292 ( 
.A(n_269),
.B(n_239),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_276),
.A2(n_204),
.B1(n_254),
.B2(n_218),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_295),
.B(n_302),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_SL g318 ( 
.A(n_296),
.B(n_230),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_L g310 ( 
.A(n_297),
.B(n_300),
.Y(n_310)
);

OAI31xp67_ASAP7_75t_L g299 ( 
.A1(n_282),
.A2(n_262),
.A3(n_270),
.B(n_273),
.Y(n_299)
);

NAND3xp33_ASAP7_75t_L g320 ( 
.A(n_299),
.B(n_304),
.C(n_205),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_294),
.B(n_285),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_292),
.B(n_258),
.C(n_267),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_305),
.B(n_307),
.Y(n_316)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_306),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_281),
.B(n_280),
.C(n_289),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_298),
.B(n_251),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_311),
.B(n_312),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_300),
.B(n_289),
.C(n_259),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_309),
.B(n_308),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_314),
.B(n_317),
.Y(n_329)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_306),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_318),
.B(n_303),
.C(n_170),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_304),
.B(n_259),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_319),
.B(n_295),
.Y(n_322)
);

NAND2x1p5_ASAP7_75t_L g323 ( 
.A(n_320),
.B(n_297),
.Y(n_323)
);

OAI21xp5_ASAP7_75t_L g321 ( 
.A1(n_305),
.A2(n_307),
.B(n_301),
.Y(n_321)
);

XOR2xp5_ASAP7_75t_L g330 ( 
.A(n_321),
.B(n_2),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_322),
.B(n_324),
.Y(n_335)
);

OAI21xp5_ASAP7_75t_L g336 ( 
.A1(n_323),
.A2(n_310),
.B(n_3),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_315),
.B(n_303),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_325),
.B(n_326),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_L g326 ( 
.A1(n_313),
.A2(n_170),
.B1(n_3),
.B2(n_4),
.Y(n_326)
);

INVxp67_ASAP7_75t_L g328 ( 
.A(n_312),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_328),
.B(n_330),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_327),
.B(n_316),
.Y(n_333)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_333),
.Y(n_339)
);

AOI31xp67_ASAP7_75t_L g334 ( 
.A1(n_329),
.A2(n_320),
.A3(n_310),
.B(n_4),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_334),
.B(n_323),
.C(n_4),
.Y(n_337)
);

OAI21xp5_ASAP7_75t_L g338 ( 
.A1(n_336),
.A2(n_328),
.B(n_3),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_337),
.B(n_338),
.Y(n_340)
);

OAI21xp5_ASAP7_75t_SL g341 ( 
.A1(n_340),
.A2(n_339),
.B(n_332),
.Y(n_341)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_341),
.B(n_335),
.C(n_331),
.Y(n_342)
);

XOR2xp5_ASAP7_75t_L g343 ( 
.A(n_342),
.B(n_4),
.Y(n_343)
);


endmodule