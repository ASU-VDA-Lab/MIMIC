module fake_jpeg_1817_n_158 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_158);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_158;

wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_24),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_23),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_5),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

BUFx5_ASAP7_75t_L g45 ( 
.A(n_3),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_12),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_25),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_34),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_8),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_2),
.Y(n_50)
);

BUFx5_ASAP7_75t_L g51 ( 
.A(n_1),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_32),
.Y(n_52)
);

BUFx5_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

INVx13_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

BUFx12_ASAP7_75t_L g55 ( 
.A(n_0),
.Y(n_55)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_52),
.Y(n_56)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_56),
.Y(n_67)
);

OR2x2_ASAP7_75t_L g57 ( 
.A(n_50),
.B(n_0),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_57),
.B(n_49),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_43),
.B(n_1),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_58),
.B(n_62),
.Y(n_63)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_52),
.Y(n_59)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_59),
.Y(n_73)
);

INVx11_ASAP7_75t_L g60 ( 
.A(n_52),
.Y(n_60)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_60),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_54),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_61),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_52),
.B(n_40),
.Y(n_62)
);

OAI22xp33_ASAP7_75t_L g64 ( 
.A1(n_59),
.A2(n_49),
.B1(n_46),
.B2(n_48),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_64),
.A2(n_65),
.B1(n_57),
.B2(n_50),
.Y(n_78)
);

OA22x2_ASAP7_75t_L g65 ( 
.A1(n_61),
.A2(n_54),
.B1(n_47),
.B2(n_44),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_61),
.Y(n_66)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_66),
.Y(n_83)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_58),
.Y(n_68)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_68),
.Y(n_86)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_56),
.Y(n_71)
);

BUFx2_ASAP7_75t_L g80 ( 
.A(n_71),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_72),
.B(n_47),
.Y(n_81)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_56),
.Y(n_74)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_74),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_63),
.B(n_57),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_76),
.B(n_78),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_65),
.B(n_48),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_77),
.B(n_85),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_64),
.B(n_57),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_79),
.B(n_82),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_81),
.B(n_88),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_65),
.B(n_62),
.Y(n_82)
);

INVx5_ASAP7_75t_L g84 ( 
.A(n_70),
.Y(n_84)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_84),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_73),
.B(n_42),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_70),
.B(n_41),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_87),
.B(n_4),
.Y(n_105)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_67),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_69),
.B(n_42),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_89),
.B(n_19),
.Y(n_97)
);

A2O1A1Ixp33_ASAP7_75t_L g91 ( 
.A1(n_79),
.A2(n_44),
.B(n_60),
.C(n_53),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_91),
.B(n_9),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_78),
.A2(n_67),
.B1(n_60),
.B2(n_51),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_92),
.A2(n_98),
.B1(n_100),
.B2(n_101),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_86),
.B(n_2),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_94),
.B(n_103),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_97),
.B(n_104),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_89),
.A2(n_51),
.B1(n_45),
.B2(n_53),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_83),
.B(n_55),
.C(n_18),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_99),
.B(n_11),
.C(n_13),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_75),
.A2(n_45),
.B1(n_55),
.B2(n_5),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_75),
.A2(n_55),
.B1(n_4),
.B2(n_6),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_80),
.B(n_3),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_80),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_105),
.B(n_39),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_SL g106 ( 
.A1(n_88),
.A2(n_6),
.B(n_7),
.Y(n_106)
);

XNOR2xp5_ASAP7_75t_L g118 ( 
.A(n_106),
.B(n_101),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_93),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_107),
.B(n_115),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_95),
.A2(n_84),
.B1(n_8),
.B2(n_9),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_108),
.A2(n_119),
.B1(n_121),
.B2(n_114),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_SL g110 ( 
.A(n_96),
.B(n_21),
.Y(n_110)
);

XNOR2xp5_ASAP7_75t_SL g132 ( 
.A(n_110),
.B(n_118),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_111),
.B(n_117),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_97),
.B(n_7),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_112),
.B(n_121),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_SL g125 ( 
.A1(n_113),
.A2(n_122),
.B(n_123),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_90),
.B(n_10),
.Y(n_115)
);

CKINVDCx10_ASAP7_75t_R g116 ( 
.A(n_102),
.Y(n_116)
);

BUFx5_ASAP7_75t_L g126 ( 
.A(n_116),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_91),
.B(n_10),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_92),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_119)
);

CKINVDCx16_ASAP7_75t_R g120 ( 
.A(n_98),
.Y(n_120)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_120),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_106),
.B(n_14),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_99),
.B(n_14),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_124),
.A2(n_100),
.B1(n_16),
.B2(n_17),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_127),
.A2(n_131),
.B1(n_27),
.B2(n_28),
.Y(n_140)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_116),
.Y(n_129)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_129),
.Y(n_142)
);

AOI21xp5_ASAP7_75t_L g130 ( 
.A1(n_118),
.A2(n_37),
.B(n_20),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_SL g144 ( 
.A1(n_130),
.A2(n_30),
.B(n_31),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_124),
.A2(n_15),
.B1(n_22),
.B2(n_26),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_109),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_134),
.B(n_135),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_128),
.B(n_110),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_138),
.B(n_140),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_L g139 ( 
.A(n_132),
.B(n_133),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_139),
.B(n_130),
.C(n_125),
.Y(n_148)
);

NOR2xp67_ASAP7_75t_L g141 ( 
.A(n_132),
.B(n_29),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_141),
.B(n_144),
.Y(n_147)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_142),
.Y(n_146)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_146),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_148),
.B(n_143),
.Y(n_149)
);

NAND2xp33_ASAP7_75t_SL g152 ( 
.A(n_149),
.B(n_151),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_147),
.B(n_137),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_SL g153 ( 
.A1(n_152),
.A2(n_145),
.B(n_140),
.Y(n_153)
);

AND3x1_ASAP7_75t_L g154 ( 
.A(n_153),
.B(n_131),
.C(n_127),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_154),
.B(n_136),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_155),
.B(n_139),
.C(n_150),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_L g157 ( 
.A1(n_156),
.A2(n_126),
.B(n_33),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_157),
.B(n_126),
.Y(n_158)
);


endmodule