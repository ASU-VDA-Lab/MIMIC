module fake_netlist_1_941_n_147 (n_20, n_2, n_5, n_8, n_11, n_16, n_13, n_3, n_18, n_0, n_1, n_12, n_9, n_17, n_14, n_10, n_15, n_19, n_21, n_6, n_4, n_7, n_147);
input n_20;
input n_2;
input n_5;
input n_8;
input n_11;
input n_16;
input n_13;
input n_3;
input n_18;
input n_0;
input n_1;
input n_12;
input n_9;
input n_17;
input n_14;
input n_10;
input n_15;
input n_19;
input n_21;
input n_6;
input n_4;
input n_7;
output n_147;
wire n_117;
wire n_44;
wire n_133;
wire n_81;
wire n_69;
wire n_22;
wire n_57;
wire n_88;
wire n_52;
wire n_26;
wire n_50;
wire n_33;
wire n_102;
wire n_73;
wire n_49;
wire n_119;
wire n_141;
wire n_115;
wire n_97;
wire n_80;
wire n_107;
wire n_60;
wire n_114;
wire n_121;
wire n_41;
wire n_35;
wire n_94;
wire n_65;
wire n_125;
wire n_130;
wire n_103;
wire n_87;
wire n_137;
wire n_104;
wire n_98;
wire n_74;
wire n_29;
wire n_146;
wire n_45;
wire n_85;
wire n_101;
wire n_62;
wire n_36;
wire n_47;
wire n_37;
wire n_34;
wire n_23;
wire n_91;
wire n_108;
wire n_116;
wire n_139;
wire n_113;
wire n_95;
wire n_124;
wire n_128;
wire n_120;
wire n_129;
wire n_70;
wire n_63;
wire n_71;
wire n_90;
wire n_56;
wire n_135;
wire n_42;
wire n_24;
wire n_78;
wire n_127;
wire n_40;
wire n_111;
wire n_79;
wire n_38;
wire n_64;
wire n_142;
wire n_46;
wire n_31;
wire n_58;
wire n_122;
wire n_138;
wire n_126;
wire n_118;
wire n_32;
wire n_84;
wire n_131;
wire n_112;
wire n_55;
wire n_86;
wire n_143;
wire n_75;
wire n_105;
wire n_72;
wire n_136;
wire n_76;
wire n_43;
wire n_89;
wire n_68;
wire n_144;
wire n_27;
wire n_53;
wire n_67;
wire n_77;
wire n_54;
wire n_123;
wire n_83;
wire n_28;
wire n_48;
wire n_100;
wire n_92;
wire n_25;
wire n_30;
wire n_59;
wire n_110;
wire n_66;
wire n_134;
wire n_82;
wire n_106;
wire n_145;
wire n_61;
wire n_99;
wire n_109;
wire n_93;
wire n_132;
wire n_51;
wire n_140;
wire n_96;
wire n_39;
INVxp67_ASAP7_75t_SL g22 ( .A(n_13), .Y(n_22) );
INVx2_ASAP7_75t_L g23 ( .A(n_14), .Y(n_23) );
INVx2_ASAP7_75t_L g24 ( .A(n_10), .Y(n_24) );
INVxp33_ASAP7_75t_L g25 ( .A(n_6), .Y(n_25) );
BUFx6f_ASAP7_75t_L g26 ( .A(n_11), .Y(n_26) );
INVx1_ASAP7_75t_L g27 ( .A(n_20), .Y(n_27) );
INVx1_ASAP7_75t_L g28 ( .A(n_2), .Y(n_28) );
INVx2_ASAP7_75t_L g29 ( .A(n_16), .Y(n_29) );
BUFx3_ASAP7_75t_L g30 ( .A(n_4), .Y(n_30) );
INVx3_ASAP7_75t_L g31 ( .A(n_17), .Y(n_31) );
INVxp33_ASAP7_75t_SL g32 ( .A(n_19), .Y(n_32) );
INVxp67_ASAP7_75t_SL g33 ( .A(n_18), .Y(n_33) );
BUFx3_ASAP7_75t_L g34 ( .A(n_12), .Y(n_34) );
NAND2xp5_ASAP7_75t_SL g35 ( .A(n_25), .B(n_0), .Y(n_35) );
BUFx6f_ASAP7_75t_L g36 ( .A(n_26), .Y(n_36) );
INVx1_ASAP7_75t_L g37 ( .A(n_27), .Y(n_37) );
INVx3_ASAP7_75t_L g38 ( .A(n_31), .Y(n_38) );
BUFx6f_ASAP7_75t_L g39 ( .A(n_26), .Y(n_39) );
INVx3_ASAP7_75t_L g40 ( .A(n_31), .Y(n_40) );
OAI21x1_ASAP7_75t_L g41 ( .A1(n_31), .A2(n_7), .B(n_5), .Y(n_41) );
OAI21x1_ASAP7_75t_L g42 ( .A1(n_23), .A2(n_9), .B(n_8), .Y(n_42) );
BUFx6f_ASAP7_75t_L g43 ( .A(n_26), .Y(n_43) );
BUFx2_ASAP7_75t_L g44 ( .A(n_30), .Y(n_44) );
INVx1_ASAP7_75t_L g45 ( .A(n_38), .Y(n_45) );
INVx2_ASAP7_75t_L g46 ( .A(n_36), .Y(n_46) );
INVx4_ASAP7_75t_L g47 ( .A(n_38), .Y(n_47) );
BUFx3_ASAP7_75t_L g48 ( .A(n_38), .Y(n_48) );
AND2x6_ASAP7_75t_L g49 ( .A(n_38), .B(n_34), .Y(n_49) );
BUFx3_ASAP7_75t_L g50 ( .A(n_40), .Y(n_50) );
BUFx6f_ASAP7_75t_L g51 ( .A(n_36), .Y(n_51) );
INVx2_ASAP7_75t_L g52 ( .A(n_36), .Y(n_52) );
AND2x4_ASAP7_75t_L g53 ( .A(n_44), .B(n_28), .Y(n_53) );
BUFx4f_ASAP7_75t_L g54 ( .A(n_37), .Y(n_54) );
INVx2_ASAP7_75t_L g55 ( .A(n_36), .Y(n_55) );
BUFx6f_ASAP7_75t_L g56 ( .A(n_36), .Y(n_56) );
INVx2_ASAP7_75t_L g57 ( .A(n_36), .Y(n_57) );
AOI21xp5_ASAP7_75t_L g58 ( .A1(n_54), .A2(n_42), .B(n_41), .Y(n_58) );
INVx2_ASAP7_75t_L g59 ( .A(n_47), .Y(n_59) );
INVx3_ASAP7_75t_L g60 ( .A(n_48), .Y(n_60) );
AND2x4_ASAP7_75t_L g61 ( .A(n_53), .B(n_35), .Y(n_61) );
INVx3_ASAP7_75t_L g62 ( .A(n_50), .Y(n_62) );
OAI21xp5_ASAP7_75t_L g63 ( .A1(n_45), .A2(n_42), .B(n_41), .Y(n_63) );
BUFx6f_ASAP7_75t_L g64 ( .A(n_49), .Y(n_64) );
BUFx2_ASAP7_75t_L g65 ( .A(n_49), .Y(n_65) );
INVx3_ASAP7_75t_L g66 ( .A(n_49), .Y(n_66) );
BUFx2_ASAP7_75t_L g67 ( .A(n_49), .Y(n_67) );
BUFx6f_ASAP7_75t_L g68 ( .A(n_54), .Y(n_68) );
BUFx6f_ASAP7_75t_L g69 ( .A(n_51), .Y(n_69) );
BUFx6f_ASAP7_75t_L g70 ( .A(n_51), .Y(n_70) );
INVx2_ASAP7_75t_L g71 ( .A(n_46), .Y(n_71) );
INVx5_ASAP7_75t_L g72 ( .A(n_51), .Y(n_72) );
INVx2_ASAP7_75t_L g73 ( .A(n_46), .Y(n_73) );
INVx3_ASAP7_75t_L g74 ( .A(n_60), .Y(n_74) );
INVx3_ASAP7_75t_L g75 ( .A(n_60), .Y(n_75) );
BUFx6f_ASAP7_75t_L g76 ( .A(n_64), .Y(n_76) );
NAND2xp5_ASAP7_75t_L g77 ( .A(n_61), .B(n_32), .Y(n_77) );
BUFx6f_ASAP7_75t_L g78 ( .A(n_64), .Y(n_78) );
INVx3_ASAP7_75t_L g79 ( .A(n_62), .Y(n_79) );
AOI21xp5_ASAP7_75t_L g80 ( .A1(n_58), .A2(n_33), .B(n_22), .Y(n_80) );
INVx3_ASAP7_75t_L g81 ( .A(n_62), .Y(n_81) );
HB1xp67_ASAP7_75t_L g82 ( .A(n_65), .Y(n_82) );
INVx1_ASAP7_75t_SL g83 ( .A(n_67), .Y(n_83) );
INVxp67_ASAP7_75t_L g84 ( .A(n_59), .Y(n_84) );
O2A1O1Ixp5_ASAP7_75t_L g85 ( .A1(n_63), .A2(n_24), .B(n_29), .C(n_23), .Y(n_85) );
INVx8_ASAP7_75t_L g86 ( .A(n_68), .Y(n_86) );
BUFx2_ASAP7_75t_L g87 ( .A(n_68), .Y(n_87) );
INVxp67_ASAP7_75t_SL g88 ( .A(n_66), .Y(n_88) );
AOI21xp5_ASAP7_75t_L g89 ( .A1(n_80), .A2(n_73), .B(n_71), .Y(n_89) );
OR2x2_ASAP7_75t_L g90 ( .A(n_77), .B(n_1), .Y(n_90) );
AOI21xp5_ASAP7_75t_L g91 ( .A1(n_80), .A2(n_70), .B(n_69), .Y(n_91) );
OAI21x1_ASAP7_75t_L g92 ( .A1(n_85), .A2(n_52), .B(n_46), .Y(n_92) );
AND2x4_ASAP7_75t_L g93 ( .A(n_82), .B(n_72), .Y(n_93) );
BUFx6f_ASAP7_75t_L g94 ( .A(n_76), .Y(n_94) );
CKINVDCx11_ASAP7_75t_R g95 ( .A(n_86), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_84), .Y(n_96) );
AOI21xp5_ASAP7_75t_L g97 ( .A1(n_88), .A2(n_70), .B(n_69), .Y(n_97) );
OAI22xp5_ASAP7_75t_L g98 ( .A1(n_83), .A2(n_39), .B1(n_43), .B2(n_36), .Y(n_98) );
AOI21xp33_ASAP7_75t_L g99 ( .A1(n_87), .A2(n_39), .B(n_36), .Y(n_99) );
OAI21x1_ASAP7_75t_L g100 ( .A1(n_91), .A2(n_75), .B(n_74), .Y(n_100) );
OAI21x1_ASAP7_75t_L g101 ( .A1(n_91), .A2(n_81), .B(n_79), .Y(n_101) );
AOI21x1_ASAP7_75t_L g102 ( .A1(n_98), .A2(n_55), .B(n_52), .Y(n_102) );
AOI21xp5_ASAP7_75t_L g103 ( .A1(n_89), .A2(n_78), .B(n_76), .Y(n_103) );
OAI21x1_ASAP7_75t_L g104 ( .A1(n_92), .A2(n_55), .B(n_52), .Y(n_104) );
OAI21x1_ASAP7_75t_L g105 ( .A1(n_97), .A2(n_57), .B(n_56), .Y(n_105) );
AOI22xp33_ASAP7_75t_L g106 ( .A1(n_90), .A2(n_56), .B1(n_51), .B2(n_3), .Y(n_106) );
BUFx6f_ASAP7_75t_L g107 ( .A(n_95), .Y(n_107) );
INVx3_ASAP7_75t_L g108 ( .A(n_93), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_96), .Y(n_109) );
BUFx6f_ASAP7_75t_L g110 ( .A(n_94), .Y(n_110) );
AO21x2_ASAP7_75t_L g111 ( .A1(n_99), .A2(n_15), .B(n_21), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_109), .Y(n_112) );
INVx2_ASAP7_75t_L g113 ( .A(n_105), .Y(n_113) );
INVx2_ASAP7_75t_L g114 ( .A(n_100), .Y(n_114) );
INVx2_ASAP7_75t_L g115 ( .A(n_101), .Y(n_115) );
INVx2_ASAP7_75t_L g116 ( .A(n_110), .Y(n_116) );
INVx2_ASAP7_75t_L g117 ( .A(n_104), .Y(n_117) );
OR2x2_ASAP7_75t_L g118 ( .A(n_108), .B(n_107), .Y(n_118) );
INVx2_ASAP7_75t_L g119 ( .A(n_102), .Y(n_119) );
AND2x2_ASAP7_75t_L g120 ( .A(n_112), .B(n_106), .Y(n_120) );
INVx2_ASAP7_75t_L g121 ( .A(n_113), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_119), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_119), .Y(n_123) );
INVx2_ASAP7_75t_L g124 ( .A(n_117), .Y(n_124) );
AO21x2_ASAP7_75t_L g125 ( .A1(n_114), .A2(n_103), .B(n_111), .Y(n_125) );
HB1xp67_ASAP7_75t_L g126 ( .A(n_118), .Y(n_126) );
INVx2_ASAP7_75t_L g127 ( .A(n_116), .Y(n_127) );
INVx2_ASAP7_75t_L g128 ( .A(n_115), .Y(n_128) );
INVx2_ASAP7_75t_L g129 ( .A(n_122), .Y(n_129) );
INVx2_ASAP7_75t_L g130 ( .A(n_123), .Y(n_130) );
NAND2xp5_ASAP7_75t_L g131 ( .A(n_120), .B(n_126), .Y(n_131) );
INVx2_ASAP7_75t_L g132 ( .A(n_121), .Y(n_132) );
INVx2_ASAP7_75t_L g133 ( .A(n_121), .Y(n_133) );
OR2x2_ASAP7_75t_L g134 ( .A(n_131), .B(n_127), .Y(n_134) );
INVx2_ASAP7_75t_L g135 ( .A(n_129), .Y(n_135) );
INVx2_ASAP7_75t_L g136 ( .A(n_129), .Y(n_136) );
INVx1_ASAP7_75t_L g137 ( .A(n_134), .Y(n_137) );
INVx1_ASAP7_75t_L g138 ( .A(n_134), .Y(n_138) );
NAND2xp5_ASAP7_75t_L g139 ( .A(n_138), .B(n_137), .Y(n_139) );
INVx1_ASAP7_75t_L g140 ( .A(n_139), .Y(n_140) );
INVx1_ASAP7_75t_L g141 ( .A(n_140), .Y(n_141) );
HB1xp67_ASAP7_75t_L g142 ( .A(n_141), .Y(n_142) );
INVx1_ASAP7_75t_L g143 ( .A(n_142), .Y(n_143) );
OAI22x1_ASAP7_75t_SL g144 ( .A1(n_143), .A2(n_135), .B1(n_136), .B2(n_130), .Y(n_144) );
XNOR2xp5_ASAP7_75t_L g145 ( .A(n_144), .B(n_125), .Y(n_145) );
OAI22xp5_ASAP7_75t_L g146 ( .A1(n_145), .A2(n_132), .B1(n_133), .B2(n_128), .Y(n_146) );
AOI21xp5_ASAP7_75t_L g147 ( .A1(n_146), .A2(n_133), .B(n_124), .Y(n_147) );
endmodule