module fake_jpeg_21274_n_129 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_129);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_129;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_9),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_11),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_2),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

INVx4_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_0),
.Y(n_20)
);

INVx3_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_9),
.Y(n_22)
);

BUFx10_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_0),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_12),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_26),
.Y(n_27)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_27),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_14),
.B(n_1),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_SL g50 ( 
.A(n_28),
.B(n_29),
.Y(n_50)
);

NOR2xp67_ASAP7_75t_L g29 ( 
.A(n_14),
.B(n_2),
.Y(n_29)
);

CKINVDCx9p33_ASAP7_75t_R g30 ( 
.A(n_23),
.Y(n_30)
);

INVx1_ASAP7_75t_SL g56 ( 
.A(n_30),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_26),
.Y(n_31)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_15),
.B(n_3),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_32),
.B(n_38),
.Y(n_48)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_26),
.Y(n_33)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_33),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_SL g34 ( 
.A(n_15),
.B(n_3),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_34),
.Y(n_49)
);

BUFx4f_ASAP7_75t_SL g35 ( 
.A(n_23),
.Y(n_35)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_35),
.Y(n_57)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

INVx13_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

BUFx4f_ASAP7_75t_SL g37 ( 
.A(n_23),
.Y(n_37)
);

OR2x2_ASAP7_75t_SL g53 ( 
.A(n_37),
.B(n_41),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_16),
.B(n_4),
.Y(n_38)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_39),
.A2(n_40),
.B1(n_18),
.B2(n_21),
.Y(n_45)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_21),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_18),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_31),
.B(n_23),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_44),
.B(n_46),
.Y(n_76)
);

CKINVDCx16_ASAP7_75t_R g64 ( 
.A(n_45),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_33),
.B(n_23),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_L g47 ( 
.A1(n_27),
.A2(n_21),
.B1(n_25),
.B2(n_24),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_47),
.A2(n_54),
.B1(n_37),
.B2(n_5),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_39),
.A2(n_30),
.B1(n_40),
.B2(n_25),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_L g73 ( 
.A1(n_51),
.A2(n_58),
.B1(n_4),
.B2(n_6),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_36),
.A2(n_22),
.B1(n_20),
.B2(n_16),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_35),
.A2(n_24),
.B1(n_22),
.B2(n_20),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_50),
.B(n_19),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_59),
.B(n_60),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_50),
.B(n_19),
.Y(n_60)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_53),
.Y(n_61)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_61),
.Y(n_87)
);

NAND3xp33_ASAP7_75t_L g62 ( 
.A(n_53),
.B(n_17),
.C(n_5),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_62),
.B(n_66),
.Y(n_77)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_54),
.Y(n_63)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_63),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_46),
.B(n_36),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_65),
.B(n_43),
.C(n_52),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_49),
.B(n_17),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_55),
.B(n_41),
.Y(n_67)
);

OAI21xp5_ASAP7_75t_SL g86 ( 
.A1(n_67),
.A2(n_69),
.B(n_71),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_48),
.B(n_41),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_68),
.B(n_75),
.Y(n_85)
);

OAI21xp33_ASAP7_75t_L g69 ( 
.A1(n_44),
.A2(n_37),
.B(n_35),
.Y(n_69)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_55),
.Y(n_70)
);

CKINVDCx16_ASAP7_75t_R g88 ( 
.A(n_70),
.Y(n_88)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_57),
.Y(n_71)
);

FAx1_ASAP7_75t_SL g80 ( 
.A(n_72),
.B(n_48),
.CI(n_56),
.CON(n_80),
.SN(n_80)
);

NAND2x1_ASAP7_75t_SL g89 ( 
.A(n_73),
.B(n_74),
.Y(n_89)
);

INVx2_ASAP7_75t_SL g74 ( 
.A(n_43),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_49),
.B(n_8),
.Y(n_75)
);

XNOR2xp5_ASAP7_75t_L g79 ( 
.A(n_76),
.B(n_61),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_79),
.B(n_81),
.C(n_83),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_80),
.A2(n_72),
.B1(n_64),
.B2(n_56),
.Y(n_92)
);

XNOR2xp5_ASAP7_75t_L g81 ( 
.A(n_65),
.B(n_57),
.Y(n_81)
);

XNOR2x1_ASAP7_75t_L g83 ( 
.A(n_69),
.B(n_42),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_84),
.B(n_67),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_88),
.Y(n_90)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_90),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_92),
.B(n_98),
.Y(n_100)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_82),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_93),
.B(n_94),
.Y(n_103)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_80),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_79),
.B(n_67),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_95),
.B(n_97),
.Y(n_102)
);

XNOR2xp5_ASAP7_75t_L g101 ( 
.A(n_96),
.B(n_84),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_81),
.B(n_42),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_80),
.B(n_85),
.Y(n_98)
);

BUFx12f_ASAP7_75t_L g99 ( 
.A(n_83),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_99),
.Y(n_107)
);

XOR2xp5_ASAP7_75t_L g112 ( 
.A(n_101),
.B(n_91),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_97),
.B(n_87),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_104),
.B(n_86),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_92),
.A2(n_87),
.B1(n_89),
.B2(n_95),
.Y(n_105)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_105),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_101),
.B(n_99),
.C(n_91),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_108),
.B(n_110),
.Y(n_118)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_106),
.Y(n_111)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_111),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_112),
.B(n_113),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_103),
.B(n_78),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_SL g114 ( 
.A(n_102),
.B(n_99),
.Y(n_114)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_114),
.B(n_100),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_116),
.B(n_112),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_109),
.A2(n_104),
.B1(n_107),
.B2(n_102),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_117),
.A2(n_70),
.B1(n_74),
.B2(n_77),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_120),
.B(n_123),
.C(n_115),
.Y(n_124)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_117),
.Y(n_121)
);

OR2x2_ASAP7_75t_L g125 ( 
.A(n_121),
.B(n_122),
.Y(n_125)
);

OAI21x1_ASAP7_75t_L g122 ( 
.A1(n_116),
.A2(n_114),
.B(n_89),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_124),
.B(n_8),
.C(n_11),
.Y(n_127)
);

AOI322xp5_ASAP7_75t_L g126 ( 
.A1(n_125),
.A2(n_119),
.A3(n_118),
.B1(n_52),
.B2(n_90),
.C1(n_74),
.C2(n_12),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_126),
.B(n_127),
.C(n_13),
.Y(n_128)
);

XOR2xp5_ASAP7_75t_L g129 ( 
.A(n_128),
.B(n_13),
.Y(n_129)
);


endmodule