module fake_jpeg_3192_n_175 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_175);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_175;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_93;
wire n_54;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_12),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_4),
.Y(n_14)
);

INVx5_ASAP7_75t_L g15 ( 
.A(n_10),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_5),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_7),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_9),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_11),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_31),
.Y(n_61)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_29),
.Y(n_32)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_32),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_33),
.Y(n_67)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_20),
.Y(n_34)
);

INVx5_ASAP7_75t_L g78 ( 
.A(n_34),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_29),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_35),
.Y(n_54)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_22),
.Y(n_36)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_36),
.Y(n_56)
);

INVx5_ASAP7_75t_L g37 ( 
.A(n_20),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_37),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_18),
.B(n_1),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_38),
.B(n_39),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_18),
.B(n_1),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

INVx1_ASAP7_75t_SL g41 ( 
.A(n_14),
.Y(n_41)
);

AND2x2_ASAP7_75t_L g60 ( 
.A(n_41),
.B(n_23),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_13),
.B(n_8),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_42),
.B(n_1),
.Y(n_76)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_20),
.Y(n_43)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_43),
.Y(n_74)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_30),
.Y(n_44)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_44),
.Y(n_59)
);

INVx5_ASAP7_75t_L g45 ( 
.A(n_15),
.Y(n_45)
);

BUFx5_ASAP7_75t_L g72 ( 
.A(n_45),
.Y(n_72)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_15),
.Y(n_46)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_46),
.Y(n_69)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_22),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_47),
.B(n_21),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_14),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_48),
.Y(n_66)
);

HB1xp67_ASAP7_75t_L g49 ( 
.A(n_28),
.Y(n_49)
);

INVxp67_ASAP7_75t_L g57 ( 
.A(n_49),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_48),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_52),
.B(n_53),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g53 ( 
.A(n_41),
.B(n_27),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_37),
.A2(n_17),
.B1(n_25),
.B2(n_19),
.Y(n_58)
);

OAI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_58),
.A2(n_32),
.B1(n_5),
.B2(n_6),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_60),
.B(n_7),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_43),
.A2(n_28),
.B1(n_25),
.B2(n_19),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_62),
.A2(n_65),
.B1(n_80),
.B2(n_3),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_63),
.B(n_64),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_35),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_43),
.A2(n_17),
.B1(n_26),
.B2(n_24),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_46),
.Y(n_68)
);

INVx2_ASAP7_75t_R g82 ( 
.A(n_68),
.Y(n_82)
);

BUFx12f_ASAP7_75t_L g70 ( 
.A(n_31),
.Y(n_70)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_70),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_45),
.B(n_26),
.Y(n_71)
);

INVxp67_ASAP7_75t_L g84 ( 
.A(n_71),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_40),
.B(n_8),
.Y(n_73)
);

CKINVDCx16_ASAP7_75t_R g85 ( 
.A(n_73),
.Y(n_85)
);

NOR2xp67_ASAP7_75t_SL g83 ( 
.A(n_76),
.B(n_3),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_34),
.B(n_2),
.Y(n_77)
);

CKINVDCx16_ASAP7_75t_R g100 ( 
.A(n_77),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_44),
.B(n_2),
.Y(n_79)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_79),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_33),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_80)
);

INVx13_ASAP7_75t_L g81 ( 
.A(n_74),
.Y(n_81)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_81),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_83),
.B(n_96),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_86),
.B(n_61),
.Y(n_113)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_50),
.Y(n_87)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_87),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_92),
.B(n_93),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_55),
.B(n_6),
.Y(n_93)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_50),
.Y(n_94)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_94),
.Y(n_112)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_66),
.Y(n_95)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_95),
.Y(n_118)
);

BUFx12_ASAP7_75t_L g97 ( 
.A(n_74),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_97),
.B(n_78),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_56),
.B(n_51),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_98),
.B(n_99),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_60),
.B(n_57),
.Y(n_99)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_66),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_101),
.B(n_102),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_57),
.B(n_59),
.Y(n_102)
);

INVx13_ASAP7_75t_L g103 ( 
.A(n_75),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_103),
.B(n_78),
.Y(n_120)
);

AOI21xp5_ASAP7_75t_SL g104 ( 
.A1(n_84),
.A2(n_65),
.B(n_58),
.Y(n_104)
);

AOI21xp5_ASAP7_75t_L g126 ( 
.A1(n_104),
.A2(n_96),
.B(n_82),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_98),
.B(n_69),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_107),
.B(n_108),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_93),
.B(n_54),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_102),
.B(n_54),
.C(n_62),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_L g136 ( 
.A(n_109),
.B(n_117),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_88),
.B(n_84),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_110),
.B(n_114),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_89),
.B(n_75),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_111),
.B(n_90),
.Y(n_123)
);

AND2x2_ASAP7_75t_L g137 ( 
.A(n_113),
.B(n_61),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_100),
.B(n_66),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_85),
.B(n_99),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_119),
.Y(n_130)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_120),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_123),
.B(n_91),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_117),
.B(n_110),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g144 ( 
.A(n_125),
.B(n_128),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_L g140 ( 
.A1(n_126),
.A2(n_127),
.B(n_106),
.Y(n_140)
);

AOI21xp5_ASAP7_75t_L g127 ( 
.A1(n_109),
.A2(n_82),
.B(n_101),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_114),
.B(n_96),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_104),
.A2(n_95),
.B1(n_87),
.B2(n_91),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_129),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_122),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_131),
.B(n_137),
.Y(n_138)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_105),
.Y(n_132)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_132),
.Y(n_145)
);

FAx1_ASAP7_75t_SL g134 ( 
.A(n_116),
.B(n_81),
.CI(n_94),
.CON(n_134),
.SN(n_134)
);

FAx1_ASAP7_75t_SL g148 ( 
.A(n_134),
.B(n_97),
.CI(n_72),
.CON(n_148),
.SN(n_148)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_135),
.A2(n_115),
.B1(n_107),
.B2(n_121),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_139),
.B(n_148),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_SL g154 ( 
.A1(n_140),
.A2(n_141),
.B(n_126),
.Y(n_154)
);

A2O1A1O1Ixp25_ASAP7_75t_L g141 ( 
.A1(n_133),
.A2(n_108),
.B(n_112),
.C(n_118),
.D(n_122),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g142 ( 
.A(n_136),
.B(n_103),
.Y(n_142)
);

XNOR2x1_ASAP7_75t_L g153 ( 
.A(n_142),
.B(n_127),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g149 ( 
.A(n_146),
.B(n_147),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_130),
.B(n_70),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_144),
.B(n_124),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_150),
.B(n_154),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_140),
.B(n_136),
.C(n_130),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_151),
.B(n_155),
.C(n_156),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_SL g161 ( 
.A(n_153),
.B(n_148),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_L g155 ( 
.A(n_142),
.B(n_135),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_139),
.B(n_133),
.C(n_132),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_152),
.A2(n_143),
.B1(n_137),
.B2(n_138),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_158),
.B(n_162),
.Y(n_165)
);

MAJx2_ASAP7_75t_L g159 ( 
.A(n_153),
.B(n_148),
.C(n_143),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_159),
.B(n_161),
.Y(n_164)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_150),
.Y(n_162)
);

AOI21xp5_ASAP7_75t_SL g163 ( 
.A1(n_157),
.A2(n_149),
.B(n_141),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_L g168 ( 
.A1(n_163),
.A2(n_167),
.B(n_129),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_160),
.B(n_145),
.Y(n_166)
);

NAND2xp33_ASAP7_75t_SL g169 ( 
.A(n_166),
.B(n_161),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_159),
.B(n_137),
.Y(n_167)
);

A2O1A1O1Ixp25_ASAP7_75t_SL g171 ( 
.A1(n_168),
.A2(n_169),
.B(n_170),
.C(n_134),
.D(n_164),
.Y(n_171)
);

INVx11_ASAP7_75t_L g170 ( 
.A(n_165),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_171),
.Y(n_173)
);

AOI322xp5_ASAP7_75t_L g172 ( 
.A1(n_170),
.A2(n_67),
.A3(n_70),
.B1(n_72),
.B2(n_97),
.C1(n_134),
.C2(n_165),
.Y(n_172)
);

HB1xp67_ASAP7_75t_L g174 ( 
.A(n_173),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_174),
.B(n_172),
.Y(n_175)
);


endmodule