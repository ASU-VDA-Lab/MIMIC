module real_jpeg_3561_n_13 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_13);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_13;

wire n_108;
wire n_54;
wire n_37;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_83;
wire n_78;
wire n_104;
wire n_64;
wire n_131;
wire n_47;
wire n_22;
wire n_87;
wire n_40;
wire n_105;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_126;
wire n_113;
wire n_120;
wire n_93;
wire n_95;
wire n_65;
wire n_33;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_66;
wire n_136;
wire n_44;
wire n_28;
wire n_62;
wire n_121;
wire n_106;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_69;
wire n_31;
wire n_129;
wire n_135;
wire n_134;
wire n_72;
wire n_100;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_110;
wire n_61;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_30;
wire n_15;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_128;
wire n_133;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_101;
wire n_96;
wire n_89;
wire n_16;

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

O2A1O1Ixp33_ASAP7_75t_L g39 ( 
.A1(n_1),
.A2(n_40),
.B(n_41),
.C(n_44),
.Y(n_39)
);

CKINVDCx16_ASAP7_75t_R g43 ( 
.A(n_1),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_1),
.B(n_71),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_1),
.A2(n_43),
.B1(n_44),
.B2(n_45),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_1),
.B(n_60),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_1),
.B(n_24),
.C(n_27),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_L g112 ( 
.A1(n_1),
.A2(n_21),
.B1(n_22),
.B2(n_43),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_1),
.B(n_50),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_1),
.B(n_35),
.Y(n_127)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_2),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_3),
.Y(n_40)
);

BUFx10_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_5),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_6),
.Y(n_74)
);

OAI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_7),
.A2(n_44),
.B1(n_45),
.B2(n_63),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_7),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_7),
.A2(n_21),
.B1(n_22),
.B2(n_63),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_7),
.A2(n_27),
.B1(n_29),
.B2(n_63),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_SL g31 ( 
.A1(n_8),
.A2(n_21),
.B1(n_22),
.B2(n_32),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_8),
.Y(n_32)
);

AOI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_8),
.A2(n_27),
.B1(n_29),
.B2(n_32),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_9),
.A2(n_27),
.B1(n_29),
.B2(n_52),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_9),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_10),
.A2(n_27),
.B1(n_29),
.B2(n_79),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_10),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g36 ( 
.A1(n_11),
.A2(n_21),
.B1(n_22),
.B2(n_37),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_11),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_L g56 ( 
.A1(n_11),
.A2(n_27),
.B1(n_29),
.B2(n_37),
.Y(n_56)
);

OAI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_11),
.A2(n_37),
.B1(n_44),
.B2(n_45),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

XOR2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_91),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_89),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_SL g15 ( 
.A(n_16),
.B(n_80),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_16),
.B(n_80),
.Y(n_90)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_57),
.Y(n_16)
);

XNOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_38),
.Y(n_17)
);

AOI21xp5_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_30),
.B(n_33),
.Y(n_18)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_19),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_19),
.B(n_36),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_26),
.Y(n_19)
);

OAI22xp33_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_22),
.B1(n_24),
.B2(n_25),
.Y(n_20)
);

OAI21xp33_ASAP7_75t_L g41 ( 
.A1(n_21),
.A2(n_42),
.B(n_43),
.Y(n_41)
);

AO22x2_ASAP7_75t_L g60 ( 
.A1(n_21),
.A2(n_22),
.B1(n_40),
.B2(n_42),
.Y(n_60)
);

INVx5_ASAP7_75t_SL g21 ( 
.A(n_22),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_22),
.B(n_110),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

INVx13_ASAP7_75t_L g25 ( 
.A(n_24),
.Y(n_25)
);

OA22x2_ASAP7_75t_L g26 ( 
.A1(n_24),
.A2(n_25),
.B1(n_27),
.B2(n_29),
.Y(n_26)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_26),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_26),
.A2(n_31),
.B1(n_83),
.B2(n_84),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_L g95 ( 
.A1(n_26),
.A2(n_84),
.B(n_96),
.Y(n_95)
);

INVx5_ASAP7_75t_L g29 ( 
.A(n_27),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_27),
.B(n_49),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_27),
.B(n_121),
.Y(n_120)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVxp67_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVxp67_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

OAI21xp5_ASAP7_75t_SL g111 ( 
.A1(n_34),
.A2(n_83),
.B(n_112),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_35),
.B(n_36),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_39),
.B(n_48),
.Y(n_38)
);

XOR2xp5_ASAP7_75t_L g81 ( 
.A(n_39),
.B(n_48),
.Y(n_81)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_40),
.Y(n_42)
);

O2A1O1Ixp33_ASAP7_75t_L g66 ( 
.A1(n_40),
.A2(n_44),
.B(n_60),
.C(n_67),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_40),
.B(n_44),
.Y(n_67)
);

AOI21xp5_ASAP7_75t_L g122 ( 
.A1(n_43),
.A2(n_102),
.B(n_123),
.Y(n_122)
);

OA22x2_ASAP7_75t_L g72 ( 
.A1(n_44),
.A2(n_45),
.B1(n_73),
.B2(n_75),
.Y(n_72)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

OAI21xp5_ASAP7_75t_L g48 ( 
.A1(n_49),
.A2(n_51),
.B(n_53),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_49),
.A2(n_51),
.B1(n_55),
.B2(n_78),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_49),
.B(n_56),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_49),
.A2(n_55),
.B1(n_100),
.B2(n_131),
.Y(n_130)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

AOI21xp5_ASAP7_75t_L g125 ( 
.A1(n_50),
.A2(n_54),
.B(n_126),
.Y(n_125)
);

INVxp67_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_55),
.B(n_56),
.Y(n_54)
);

OAI21xp5_ASAP7_75t_L g99 ( 
.A1(n_55),
.A2(n_100),
.B(n_101),
.Y(n_99)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_55),
.Y(n_123)
);

XOR2xp5_ASAP7_75t_L g57 ( 
.A(n_58),
.B(n_68),
.Y(n_57)
);

OAI21xp5_ASAP7_75t_SL g58 ( 
.A1(n_59),
.A2(n_61),
.B(n_64),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_60),
.B(n_65),
.Y(n_88)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_65),
.B(n_66),
.Y(n_64)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_66),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_69),
.A2(n_70),
.B1(n_76),
.B2(n_77),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx3_ASAP7_75t_SL g75 ( 
.A(n_73),
.Y(n_75)
);

INVx8_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_82),
.C(n_85),
.Y(n_80)
);

XNOR2xp5_ASAP7_75t_L g103 ( 
.A(n_81),
.B(n_104),
.Y(n_103)
);

XNOR2xp5_ASAP7_75t_L g104 ( 
.A(n_82),
.B(n_85),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_SL g85 ( 
.A1(n_86),
.A2(n_87),
.B(n_88),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_L g91 ( 
.A1(n_92),
.A2(n_105),
.B(n_136),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_103),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_93),
.B(n_103),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_97),
.C(n_98),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_94),
.A2(n_95),
.B1(n_97),
.B2(n_115),
.Y(n_114)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_97),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_98),
.A2(n_99),
.B1(n_114),
.B2(n_116),
.Y(n_113)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

AOI21xp5_ASAP7_75t_L g105 ( 
.A1(n_106),
.A2(n_117),
.B(n_135),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_107),
.B(n_113),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_107),
.B(n_113),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_111),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_108),
.A2(n_109),
.B1(n_111),
.B2(n_133),
.Y(n_132)
);

CKINVDCx16_ASAP7_75t_R g108 ( 
.A(n_109),
.Y(n_108)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_111),
.Y(n_133)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_114),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_L g117 ( 
.A1(n_118),
.A2(n_129),
.B(n_134),
.Y(n_117)
);

AOI21xp5_ASAP7_75t_L g118 ( 
.A1(n_119),
.A2(n_124),
.B(n_128),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_120),
.B(n_122),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_125),
.B(n_127),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_125),
.B(n_127),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_126),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_132),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_130),
.B(n_132),
.Y(n_134)
);


endmodule