module fake_netlist_6_2438_n_1783 (n_52, n_435, n_1, n_91, n_326, n_256, n_209, n_367, n_63, n_223, n_278, n_341, n_362, n_148, n_226, n_161, n_22, n_208, n_68, n_316, n_419, n_28, n_304, n_212, n_50, n_7, n_144, n_365, n_125, n_168, n_384, n_297, n_342, n_77, n_106, n_358, n_160, n_131, n_188, n_310, n_186, n_245, n_0, n_368, n_396, n_350, n_78, n_84, n_392, n_142, n_143, n_382, n_180, n_62, n_349, n_233, n_255, n_284, n_400, n_140, n_337, n_214, n_67, n_15, n_246, n_38, n_289, n_421, n_424, n_59, n_181, n_182, n_238, n_202, n_320, n_108, n_327, n_369, n_280, n_287, n_353, n_389, n_415, n_65, n_230, n_141, n_383, n_200, n_176, n_114, n_86, n_198, n_104, n_222, n_179, n_248, n_300, n_71, n_74, n_229, n_305, n_72, n_173, n_250, n_372, n_111, n_314, n_378, n_413, n_377, n_35, n_183, n_79, n_375, n_338, n_56, n_360, n_119, n_235, n_147, n_191, n_340, n_387, n_39, n_344, n_73, n_428, n_432, n_101, n_167, n_174, n_127, n_153, n_156, n_145, n_42, n_133, n_96, n_8, n_371, n_189, n_405, n_213, n_294, n_302, n_380, n_129, n_197, n_11, n_137, n_17, n_343, n_20, n_397, n_155, n_109, n_425, n_122, n_45, n_34, n_218, n_70, n_234, n_37, n_381, n_82, n_27, n_236, n_112, n_172, n_270, n_239, n_126, n_414, n_97, n_58, n_290, n_220, n_118, n_224, n_48, n_25, n_93, n_80, n_196, n_402, n_352, n_9, n_107, n_6, n_417, n_14, n_89, n_374, n_366, n_407, n_103, n_272, n_185, n_348, n_69, n_376, n_390, n_293, n_31, n_334, n_53, n_370, n_44, n_232, n_16, n_163, n_46, n_330, n_298, n_18, n_281, n_258, n_154, n_98, n_260, n_265, n_313, n_279, n_252, n_228, n_356, n_166, n_184, n_216, n_83, n_363, n_395, n_323, n_393, n_411, n_152, n_92, n_321, n_331, n_105, n_227, n_132, n_406, n_102, n_204, n_261, n_420, n_312, n_394, n_32, n_66, n_130, n_164, n_292, n_100, n_121, n_307, n_433, n_23, n_2, n_291, n_219, n_357, n_150, n_264, n_263, n_325, n_329, n_33, n_408, n_61, n_237, n_244, n_399, n_76, n_243, n_124, n_94, n_282, n_436, n_116, n_211, n_117, n_175, n_322, n_345, n_409, n_231, n_354, n_40, n_240, n_139, n_319, n_41, n_134, n_273, n_95, n_311, n_10, n_403, n_253, n_123, n_136, n_249, n_201, n_386, n_159, n_157, n_162, n_115, n_128, n_241, n_30, n_275, n_43, n_276, n_221, n_423, n_146, n_318, n_303, n_306, n_21, n_193, n_269, n_359, n_346, n_88, n_3, n_416, n_277, n_418, n_113, n_4, n_199, n_138, n_266, n_296, n_268, n_271, n_404, n_158, n_217, n_49, n_210, n_299, n_206, n_5, n_333, n_215, n_178, n_247, n_225, n_308, n_309, n_355, n_426, n_317, n_149, n_431, n_90, n_347, n_24, n_54, n_328, n_429, n_373, n_87, n_195, n_285, n_85, n_99, n_257, n_13, n_203, n_286, n_254, n_207, n_242, n_19, n_47, n_29, n_75, n_401, n_324, n_335, n_430, n_205, n_120, n_251, n_301, n_274, n_110, n_151, n_412, n_81, n_36, n_26, n_55, n_267, n_339, n_315, n_434, n_64, n_288, n_427, n_422, n_135, n_165, n_351, n_437, n_259, n_177, n_391, n_364, n_295, n_385, n_388, n_190, n_262, n_187, n_60, n_361, n_379, n_170, n_332, n_336, n_12, n_398, n_410, n_194, n_171, n_192, n_57, n_169, n_51, n_283, n_1783);

input n_52;
input n_435;
input n_1;
input n_91;
input n_326;
input n_256;
input n_209;
input n_367;
input n_63;
input n_223;
input n_278;
input n_341;
input n_362;
input n_148;
input n_226;
input n_161;
input n_22;
input n_208;
input n_68;
input n_316;
input n_419;
input n_28;
input n_304;
input n_212;
input n_50;
input n_7;
input n_144;
input n_365;
input n_125;
input n_168;
input n_384;
input n_297;
input n_342;
input n_77;
input n_106;
input n_358;
input n_160;
input n_131;
input n_188;
input n_310;
input n_186;
input n_245;
input n_0;
input n_368;
input n_396;
input n_350;
input n_78;
input n_84;
input n_392;
input n_142;
input n_143;
input n_382;
input n_180;
input n_62;
input n_349;
input n_233;
input n_255;
input n_284;
input n_400;
input n_140;
input n_337;
input n_214;
input n_67;
input n_15;
input n_246;
input n_38;
input n_289;
input n_421;
input n_424;
input n_59;
input n_181;
input n_182;
input n_238;
input n_202;
input n_320;
input n_108;
input n_327;
input n_369;
input n_280;
input n_287;
input n_353;
input n_389;
input n_415;
input n_65;
input n_230;
input n_141;
input n_383;
input n_200;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_179;
input n_248;
input n_300;
input n_71;
input n_74;
input n_229;
input n_305;
input n_72;
input n_173;
input n_250;
input n_372;
input n_111;
input n_314;
input n_378;
input n_413;
input n_377;
input n_35;
input n_183;
input n_79;
input n_375;
input n_338;
input n_56;
input n_360;
input n_119;
input n_235;
input n_147;
input n_191;
input n_340;
input n_387;
input n_39;
input n_344;
input n_73;
input n_428;
input n_432;
input n_101;
input n_167;
input n_174;
input n_127;
input n_153;
input n_156;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_371;
input n_189;
input n_405;
input n_213;
input n_294;
input n_302;
input n_380;
input n_129;
input n_197;
input n_11;
input n_137;
input n_17;
input n_343;
input n_20;
input n_397;
input n_155;
input n_109;
input n_425;
input n_122;
input n_45;
input n_34;
input n_218;
input n_70;
input n_234;
input n_37;
input n_381;
input n_82;
input n_27;
input n_236;
input n_112;
input n_172;
input n_270;
input n_239;
input n_126;
input n_414;
input n_97;
input n_58;
input n_290;
input n_220;
input n_118;
input n_224;
input n_48;
input n_25;
input n_93;
input n_80;
input n_196;
input n_402;
input n_352;
input n_9;
input n_107;
input n_6;
input n_417;
input n_14;
input n_89;
input n_374;
input n_366;
input n_407;
input n_103;
input n_272;
input n_185;
input n_348;
input n_69;
input n_376;
input n_390;
input n_293;
input n_31;
input n_334;
input n_53;
input n_370;
input n_44;
input n_232;
input n_16;
input n_163;
input n_46;
input n_330;
input n_298;
input n_18;
input n_281;
input n_258;
input n_154;
input n_98;
input n_260;
input n_265;
input n_313;
input n_279;
input n_252;
input n_228;
input n_356;
input n_166;
input n_184;
input n_216;
input n_83;
input n_363;
input n_395;
input n_323;
input n_393;
input n_411;
input n_152;
input n_92;
input n_321;
input n_331;
input n_105;
input n_227;
input n_132;
input n_406;
input n_102;
input n_204;
input n_261;
input n_420;
input n_312;
input n_394;
input n_32;
input n_66;
input n_130;
input n_164;
input n_292;
input n_100;
input n_121;
input n_307;
input n_433;
input n_23;
input n_2;
input n_291;
input n_219;
input n_357;
input n_150;
input n_264;
input n_263;
input n_325;
input n_329;
input n_33;
input n_408;
input n_61;
input n_237;
input n_244;
input n_399;
input n_76;
input n_243;
input n_124;
input n_94;
input n_282;
input n_436;
input n_116;
input n_211;
input n_117;
input n_175;
input n_322;
input n_345;
input n_409;
input n_231;
input n_354;
input n_40;
input n_240;
input n_139;
input n_319;
input n_41;
input n_134;
input n_273;
input n_95;
input n_311;
input n_10;
input n_403;
input n_253;
input n_123;
input n_136;
input n_249;
input n_201;
input n_386;
input n_159;
input n_157;
input n_162;
input n_115;
input n_128;
input n_241;
input n_30;
input n_275;
input n_43;
input n_276;
input n_221;
input n_423;
input n_146;
input n_318;
input n_303;
input n_306;
input n_21;
input n_193;
input n_269;
input n_359;
input n_346;
input n_88;
input n_3;
input n_416;
input n_277;
input n_418;
input n_113;
input n_4;
input n_199;
input n_138;
input n_266;
input n_296;
input n_268;
input n_271;
input n_404;
input n_158;
input n_217;
input n_49;
input n_210;
input n_299;
input n_206;
input n_5;
input n_333;
input n_215;
input n_178;
input n_247;
input n_225;
input n_308;
input n_309;
input n_355;
input n_426;
input n_317;
input n_149;
input n_431;
input n_90;
input n_347;
input n_24;
input n_54;
input n_328;
input n_429;
input n_373;
input n_87;
input n_195;
input n_285;
input n_85;
input n_99;
input n_257;
input n_13;
input n_203;
input n_286;
input n_254;
input n_207;
input n_242;
input n_19;
input n_47;
input n_29;
input n_75;
input n_401;
input n_324;
input n_335;
input n_430;
input n_205;
input n_120;
input n_251;
input n_301;
input n_274;
input n_110;
input n_151;
input n_412;
input n_81;
input n_36;
input n_26;
input n_55;
input n_267;
input n_339;
input n_315;
input n_434;
input n_64;
input n_288;
input n_427;
input n_422;
input n_135;
input n_165;
input n_351;
input n_437;
input n_259;
input n_177;
input n_391;
input n_364;
input n_295;
input n_385;
input n_388;
input n_190;
input n_262;
input n_187;
input n_60;
input n_361;
input n_379;
input n_170;
input n_332;
input n_336;
input n_12;
input n_398;
input n_410;
input n_194;
input n_171;
input n_192;
input n_57;
input n_169;
input n_51;
input n_283;

output n_1783;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_1212;
wire n_726;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_1738;
wire n_798;
wire n_1575;
wire n_509;
wire n_1342;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_1739;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1688;
wire n_1691;
wire n_1009;
wire n_1743;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_830;
wire n_461;
wire n_873;
wire n_1285;
wire n_1371;
wire n_447;
wire n_1172;
wire n_852;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1704;
wire n_1078;
wire n_544;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_616;
wire n_658;
wire n_1119;
wire n_1433;
wire n_1620;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_953;
wire n_1094;
wire n_1345;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1644;
wire n_1558;
wire n_1732;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_813;
wire n_1481;
wire n_606;
wire n_1441;
wire n_818;
wire n_1309;
wire n_1123;
wire n_513;
wire n_645;
wire n_1381;
wire n_1699;
wire n_916;
wire n_483;
wire n_608;
wire n_630;
wire n_541;
wire n_512;
wire n_792;
wire n_476;
wire n_1328;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_982;
wire n_549;
wire n_1762;
wire n_1075;
wire n_932;
wire n_1697;
wire n_979;
wire n_905;
wire n_1680;
wire n_993;
wire n_689;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1233;
wire n_1289;
wire n_487;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_1701;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_530;
wire n_1563;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_1335;
wire n_1760;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_1165;
wire n_702;
wire n_1175;
wire n_1386;
wire n_1747;
wire n_1012;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1504;
wire n_1655;
wire n_835;
wire n_928;
wire n_1214;
wire n_850;
wire n_690;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_701;
wire n_950;
wire n_484;
wire n_1709;
wire n_1757;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_595;
wire n_627;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_963;
wire n_639;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_1765;
wire n_605;
wire n_1514;
wire n_826;
wire n_1646;
wire n_1139;
wire n_872;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_996;
wire n_532;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_622;
wire n_1469;
wire n_1766;
wire n_1776;
wire n_581;
wire n_765;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_899;
wire n_738;
wire n_1304;
wire n_1035;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1577;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_1717;
wire n_926;
wire n_927;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_552;
wire n_1358;
wire n_1388;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_931;
wire n_1021;
wire n_527;
wire n_474;
wire n_683;
wire n_811;
wire n_1207;
wire n_1368;
wire n_1418;
wire n_958;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_1483;
wire n_1372;
wire n_1457;
wire n_505;
wire n_1719;
wire n_1339;
wire n_537;
wire n_1427;
wire n_1466;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_1769;
wire n_1220;
wire n_556;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_1159;
wire n_1092;
wire n_441;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1223;
wire n_511;
wire n_1286;
wire n_1775;
wire n_1773;
wire n_1053;
wire n_1681;
wire n_520;
wire n_1093;
wire n_1533;
wire n_1597;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_1745;
wire n_914;
wire n_759;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_1617;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1267;
wire n_1281;
wire n_983;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_1731;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_778;
wire n_1668;
wire n_1134;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_793;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_1744;
wire n_828;
wire n_607;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_1254;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_1468;
wire n_1095;
wire n_1595;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_597;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1024;
wire n_1768;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_750;
wire n_1115;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_1126;
wire n_710;
wire n_1108;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_1694;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_1262;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_782;
wire n_1539;
wire n_490;
wire n_809;
wire n_1043;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1361;
wire n_1491;
wire n_662;
wire n_1152;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_1695;
wire n_650;
wire n_1046;
wire n_1145;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_1406;
wire n_456;
wire n_1332;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_1222;
wire n_599;
wire n_776;
wire n_1720;
wire n_934;
wire n_482;
wire n_1637;
wire n_1407;
wire n_1341;
wire n_1456;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_1640;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_1676;
wire n_833;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_799;
wire n_1548;
wire n_1155;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1282;
wire n_550;
wire n_652;
wire n_560;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_1758;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_1373;
wire n_1292;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_1248;
wire n_1556;
wire n_902;
wire n_1047;
wire n_1385;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1236;
wire n_1559;
wire n_1725;
wire n_834;
wire n_743;
wire n_766;
wire n_1741;
wire n_1325;
wire n_1002;
wire n_1746;
wire n_545;
wire n_489;
wire n_1727;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_1098;
wire n_1329;
wire n_817;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1118;
wire n_1076;
wire n_1007;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1631;
wire n_591;
wire n_1377;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_1074;
wire n_698;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_955;
wire n_1379;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_573;
wire n_769;
wire n_676;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_814;
wire n_1643;
wire n_1729;
wire n_669;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_1408;
wire n_1196;
wire n_1598;
wire n_863;
wire n_601;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1147;
wire n_763;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1464;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_1028;
wire n_576;
wire n_472;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_712;
wire n_1276;
wire n_1148;
wire n_1161;
wire n_1085;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_1582;
wire n_492;
wire n_1149;
wire n_1184;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_1090;
wire n_592;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_984;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_735;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_1144;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1574;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_1552;
wire n_583;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_973;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_1260;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_1632;
wire n_1557;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_784;
wire n_1059;
wire n_1197;
wire n_722;
wire n_862;
wire n_540;
wire n_1423;
wire n_457;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_827;
wire n_531;
wire n_1025;
wire n_1013;
wire n_1259;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx20_ASAP7_75t_R g438 ( 
.A(n_212),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_332),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_355),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_188),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_221),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_345),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_429),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_85),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_132),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_135),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_382),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_172),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_195),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_223),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_32),
.Y(n_452)
);

BUFx2_ASAP7_75t_L g453 ( 
.A(n_51),
.Y(n_453)
);

BUFx3_ASAP7_75t_L g454 ( 
.A(n_433),
.Y(n_454)
);

CKINVDCx20_ASAP7_75t_R g455 ( 
.A(n_138),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_74),
.Y(n_456)
);

BUFx6f_ASAP7_75t_L g457 ( 
.A(n_57),
.Y(n_457)
);

CKINVDCx5p33_ASAP7_75t_R g458 ( 
.A(n_283),
.Y(n_458)
);

INVx2_ASAP7_75t_L g459 ( 
.A(n_417),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_309),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_47),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_374),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_153),
.Y(n_463)
);

BUFx2_ASAP7_75t_L g464 ( 
.A(n_237),
.Y(n_464)
);

CKINVDCx5p33_ASAP7_75t_R g465 ( 
.A(n_239),
.Y(n_465)
);

BUFx3_ASAP7_75t_L g466 ( 
.A(n_375),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_411),
.Y(n_467)
);

CKINVDCx5p33_ASAP7_75t_R g468 ( 
.A(n_21),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_70),
.Y(n_469)
);

CKINVDCx5p33_ASAP7_75t_R g470 ( 
.A(n_140),
.Y(n_470)
);

INVx2_ASAP7_75t_L g471 ( 
.A(n_182),
.Y(n_471)
);

CKINVDCx5p33_ASAP7_75t_R g472 ( 
.A(n_159),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_31),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_118),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_409),
.Y(n_475)
);

CKINVDCx5p33_ASAP7_75t_R g476 ( 
.A(n_302),
.Y(n_476)
);

CKINVDCx5p33_ASAP7_75t_R g477 ( 
.A(n_336),
.Y(n_477)
);

INVx2_ASAP7_75t_L g478 ( 
.A(n_16),
.Y(n_478)
);

INVx2_ASAP7_75t_SL g479 ( 
.A(n_431),
.Y(n_479)
);

HB1xp67_ASAP7_75t_L g480 ( 
.A(n_410),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_241),
.Y(n_481)
);

CKINVDCx5p33_ASAP7_75t_R g482 ( 
.A(n_193),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_42),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_362),
.Y(n_484)
);

INVx2_ASAP7_75t_L g485 ( 
.A(n_66),
.Y(n_485)
);

CKINVDCx5p33_ASAP7_75t_R g486 ( 
.A(n_197),
.Y(n_486)
);

CKINVDCx5p33_ASAP7_75t_R g487 ( 
.A(n_170),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_295),
.Y(n_488)
);

BUFx2_ASAP7_75t_L g489 ( 
.A(n_247),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_395),
.Y(n_490)
);

INVx2_ASAP7_75t_L g491 ( 
.A(n_192),
.Y(n_491)
);

CKINVDCx5p33_ASAP7_75t_R g492 ( 
.A(n_257),
.Y(n_492)
);

CKINVDCx5p33_ASAP7_75t_R g493 ( 
.A(n_338),
.Y(n_493)
);

CKINVDCx5p33_ASAP7_75t_R g494 ( 
.A(n_67),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_422),
.Y(n_495)
);

BUFx2_ASAP7_75t_L g496 ( 
.A(n_83),
.Y(n_496)
);

CKINVDCx5p33_ASAP7_75t_R g497 ( 
.A(n_404),
.Y(n_497)
);

CKINVDCx20_ASAP7_75t_R g498 ( 
.A(n_113),
.Y(n_498)
);

CKINVDCx5p33_ASAP7_75t_R g499 ( 
.A(n_351),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_432),
.Y(n_500)
);

CKINVDCx5p33_ASAP7_75t_R g501 ( 
.A(n_155),
.Y(n_501)
);

CKINVDCx20_ASAP7_75t_R g502 ( 
.A(n_392),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_326),
.Y(n_503)
);

CKINVDCx20_ASAP7_75t_R g504 ( 
.A(n_33),
.Y(n_504)
);

CKINVDCx5p33_ASAP7_75t_R g505 ( 
.A(n_201),
.Y(n_505)
);

CKINVDCx5p33_ASAP7_75t_R g506 ( 
.A(n_73),
.Y(n_506)
);

CKINVDCx5p33_ASAP7_75t_R g507 ( 
.A(n_152),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_68),
.Y(n_508)
);

CKINVDCx5p33_ASAP7_75t_R g509 ( 
.A(n_370),
.Y(n_509)
);

CKINVDCx5p33_ASAP7_75t_R g510 ( 
.A(n_279),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_314),
.Y(n_511)
);

CKINVDCx5p33_ASAP7_75t_R g512 ( 
.A(n_368),
.Y(n_512)
);

CKINVDCx5p33_ASAP7_75t_R g513 ( 
.A(n_333),
.Y(n_513)
);

CKINVDCx5p33_ASAP7_75t_R g514 ( 
.A(n_154),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_144),
.Y(n_515)
);

CKINVDCx5p33_ASAP7_75t_R g516 ( 
.A(n_251),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_208),
.Y(n_517)
);

CKINVDCx5p33_ASAP7_75t_R g518 ( 
.A(n_214),
.Y(n_518)
);

CKINVDCx5p33_ASAP7_75t_R g519 ( 
.A(n_115),
.Y(n_519)
);

CKINVDCx5p33_ASAP7_75t_R g520 ( 
.A(n_181),
.Y(n_520)
);

CKINVDCx5p33_ASAP7_75t_R g521 ( 
.A(n_50),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_396),
.Y(n_522)
);

CKINVDCx5p33_ASAP7_75t_R g523 ( 
.A(n_426),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_323),
.Y(n_524)
);

CKINVDCx5p33_ASAP7_75t_R g525 ( 
.A(n_235),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_380),
.Y(n_526)
);

BUFx6f_ASAP7_75t_L g527 ( 
.A(n_32),
.Y(n_527)
);

CKINVDCx5p33_ASAP7_75t_R g528 ( 
.A(n_298),
.Y(n_528)
);

CKINVDCx5p33_ASAP7_75t_R g529 ( 
.A(n_142),
.Y(n_529)
);

CKINVDCx5p33_ASAP7_75t_R g530 ( 
.A(n_271),
.Y(n_530)
);

CKINVDCx5p33_ASAP7_75t_R g531 ( 
.A(n_296),
.Y(n_531)
);

CKINVDCx5p33_ASAP7_75t_R g532 ( 
.A(n_365),
.Y(n_532)
);

CKINVDCx20_ASAP7_75t_R g533 ( 
.A(n_76),
.Y(n_533)
);

CKINVDCx5p33_ASAP7_75t_R g534 ( 
.A(n_413),
.Y(n_534)
);

BUFx10_ASAP7_75t_L g535 ( 
.A(n_420),
.Y(n_535)
);

CKINVDCx5p33_ASAP7_75t_R g536 ( 
.A(n_176),
.Y(n_536)
);

CKINVDCx16_ASAP7_75t_R g537 ( 
.A(n_307),
.Y(n_537)
);

CKINVDCx5p33_ASAP7_75t_R g538 ( 
.A(n_238),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_416),
.Y(n_539)
);

INVx2_ASAP7_75t_SL g540 ( 
.A(n_305),
.Y(n_540)
);

CKINVDCx5p33_ASAP7_75t_R g541 ( 
.A(n_169),
.Y(n_541)
);

CKINVDCx20_ASAP7_75t_R g542 ( 
.A(n_51),
.Y(n_542)
);

CKINVDCx5p33_ASAP7_75t_R g543 ( 
.A(n_408),
.Y(n_543)
);

CKINVDCx5p33_ASAP7_75t_R g544 ( 
.A(n_348),
.Y(n_544)
);

CKINVDCx5p33_ASAP7_75t_R g545 ( 
.A(n_11),
.Y(n_545)
);

CKINVDCx14_ASAP7_75t_R g546 ( 
.A(n_175),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_82),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_291),
.Y(n_548)
);

INVx2_ASAP7_75t_L g549 ( 
.A(n_297),
.Y(n_549)
);

INVx2_ASAP7_75t_SL g550 ( 
.A(n_62),
.Y(n_550)
);

BUFx6f_ASAP7_75t_L g551 ( 
.A(n_149),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_340),
.Y(n_552)
);

CKINVDCx5p33_ASAP7_75t_R g553 ( 
.A(n_322),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_277),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_150),
.Y(n_555)
);

CKINVDCx20_ASAP7_75t_R g556 ( 
.A(n_312),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_275),
.Y(n_557)
);

CKINVDCx5p33_ASAP7_75t_R g558 ( 
.A(n_196),
.Y(n_558)
);

BUFx6f_ASAP7_75t_L g559 ( 
.A(n_421),
.Y(n_559)
);

CKINVDCx20_ASAP7_75t_R g560 ( 
.A(n_94),
.Y(n_560)
);

INVx2_ASAP7_75t_L g561 ( 
.A(n_106),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_253),
.Y(n_562)
);

INVxp67_ASAP7_75t_L g563 ( 
.A(n_299),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_425),
.Y(n_564)
);

CKINVDCx5p33_ASAP7_75t_R g565 ( 
.A(n_346),
.Y(n_565)
);

CKINVDCx14_ASAP7_75t_R g566 ( 
.A(n_423),
.Y(n_566)
);

CKINVDCx5p33_ASAP7_75t_R g567 ( 
.A(n_407),
.Y(n_567)
);

INVx1_ASAP7_75t_SL g568 ( 
.A(n_80),
.Y(n_568)
);

CKINVDCx5p33_ASAP7_75t_R g569 ( 
.A(n_183),
.Y(n_569)
);

BUFx5_ASAP7_75t_L g570 ( 
.A(n_414),
.Y(n_570)
);

CKINVDCx5p33_ASAP7_75t_R g571 ( 
.A(n_415),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_139),
.Y(n_572)
);

CKINVDCx5p33_ASAP7_75t_R g573 ( 
.A(n_116),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_282),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_211),
.Y(n_575)
);

CKINVDCx5p33_ASAP7_75t_R g576 ( 
.A(n_405),
.Y(n_576)
);

CKINVDCx5p33_ASAP7_75t_R g577 ( 
.A(n_393),
.Y(n_577)
);

CKINVDCx5p33_ASAP7_75t_R g578 ( 
.A(n_4),
.Y(n_578)
);

INVx2_ASAP7_75t_L g579 ( 
.A(n_12),
.Y(n_579)
);

CKINVDCx5p33_ASAP7_75t_R g580 ( 
.A(n_315),
.Y(n_580)
);

CKINVDCx5p33_ASAP7_75t_R g581 ( 
.A(n_218),
.Y(n_581)
);

CKINVDCx5p33_ASAP7_75t_R g582 ( 
.A(n_134),
.Y(n_582)
);

CKINVDCx5p33_ASAP7_75t_R g583 ( 
.A(n_66),
.Y(n_583)
);

CKINVDCx5p33_ASAP7_75t_R g584 ( 
.A(n_427),
.Y(n_584)
);

CKINVDCx5p33_ASAP7_75t_R g585 ( 
.A(n_337),
.Y(n_585)
);

BUFx10_ASAP7_75t_L g586 ( 
.A(n_424),
.Y(n_586)
);

INVxp67_ASAP7_75t_L g587 ( 
.A(n_41),
.Y(n_587)
);

CKINVDCx5p33_ASAP7_75t_R g588 ( 
.A(n_161),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_264),
.Y(n_589)
);

CKINVDCx5p33_ASAP7_75t_R g590 ( 
.A(n_133),
.Y(n_590)
);

CKINVDCx5p33_ASAP7_75t_R g591 ( 
.A(n_2),
.Y(n_591)
);

CKINVDCx5p33_ASAP7_75t_R g592 ( 
.A(n_419),
.Y(n_592)
);

BUFx4f_ASAP7_75t_SL g593 ( 
.A(n_12),
.Y(n_593)
);

INVx1_ASAP7_75t_SL g594 ( 
.A(n_156),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_96),
.Y(n_595)
);

CKINVDCx5p33_ASAP7_75t_R g596 ( 
.A(n_352),
.Y(n_596)
);

BUFx2_ASAP7_75t_L g597 ( 
.A(n_366),
.Y(n_597)
);

CKINVDCx5p33_ASAP7_75t_R g598 ( 
.A(n_311),
.Y(n_598)
);

CKINVDCx16_ASAP7_75t_R g599 ( 
.A(n_329),
.Y(n_599)
);

CKINVDCx5p33_ASAP7_75t_R g600 ( 
.A(n_189),
.Y(n_600)
);

BUFx3_ASAP7_75t_L g601 ( 
.A(n_255),
.Y(n_601)
);

CKINVDCx16_ASAP7_75t_R g602 ( 
.A(n_244),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_104),
.Y(n_603)
);

HB1xp67_ASAP7_75t_L g604 ( 
.A(n_418),
.Y(n_604)
);

CKINVDCx5p33_ASAP7_75t_R g605 ( 
.A(n_435),
.Y(n_605)
);

INVx1_ASAP7_75t_SL g606 ( 
.A(n_210),
.Y(n_606)
);

INVxp33_ASAP7_75t_R g607 ( 
.A(n_400),
.Y(n_607)
);

CKINVDCx5p33_ASAP7_75t_R g608 ( 
.A(n_399),
.Y(n_608)
);

CKINVDCx20_ASAP7_75t_R g609 ( 
.A(n_328),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_412),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_316),
.Y(n_611)
);

CKINVDCx20_ASAP7_75t_R g612 ( 
.A(n_33),
.Y(n_612)
);

CKINVDCx5p33_ASAP7_75t_R g613 ( 
.A(n_360),
.Y(n_613)
);

CKINVDCx20_ASAP7_75t_R g614 ( 
.A(n_438),
.Y(n_614)
);

INVxp67_ASAP7_75t_L g615 ( 
.A(n_453),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_457),
.Y(n_616)
);

BUFx3_ASAP7_75t_L g617 ( 
.A(n_535),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_457),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_457),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_457),
.Y(n_620)
);

CKINVDCx5p33_ASAP7_75t_R g621 ( 
.A(n_439),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_527),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_527),
.Y(n_623)
);

CKINVDCx20_ASAP7_75t_R g624 ( 
.A(n_455),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_527),
.Y(n_625)
);

BUFx2_ASAP7_75t_L g626 ( 
.A(n_452),
.Y(n_626)
);

INVx2_ASAP7_75t_L g627 ( 
.A(n_527),
.Y(n_627)
);

BUFx2_ASAP7_75t_SL g628 ( 
.A(n_498),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_469),
.Y(n_629)
);

HB1xp67_ASAP7_75t_L g630 ( 
.A(n_461),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_473),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_483),
.Y(n_632)
);

CKINVDCx16_ASAP7_75t_R g633 ( 
.A(n_537),
.Y(n_633)
);

INVxp67_ASAP7_75t_SL g634 ( 
.A(n_587),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_440),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_443),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_447),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_456),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_462),
.Y(n_639)
);

INVx3_ASAP7_75t_L g640 ( 
.A(n_478),
.Y(n_640)
);

CKINVDCx20_ASAP7_75t_R g641 ( 
.A(n_502),
.Y(n_641)
);

CKINVDCx5p33_ASAP7_75t_R g642 ( 
.A(n_441),
.Y(n_642)
);

INVxp67_ASAP7_75t_SL g643 ( 
.A(n_587),
.Y(n_643)
);

BUFx3_ASAP7_75t_L g644 ( 
.A(n_535),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_467),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_474),
.Y(n_646)
);

BUFx3_ASAP7_75t_L g647 ( 
.A(n_586),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_475),
.Y(n_648)
);

BUFx2_ASAP7_75t_L g649 ( 
.A(n_468),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_481),
.Y(n_650)
);

BUFx6f_ASAP7_75t_L g651 ( 
.A(n_551),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_484),
.Y(n_652)
);

CKINVDCx20_ASAP7_75t_R g653 ( 
.A(n_533),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_488),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_490),
.Y(n_655)
);

HB1xp67_ASAP7_75t_L g656 ( 
.A(n_485),
.Y(n_656)
);

INVxp67_ASAP7_75t_SL g657 ( 
.A(n_508),
.Y(n_657)
);

HB1xp67_ASAP7_75t_L g658 ( 
.A(n_579),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_495),
.Y(n_659)
);

NOR2xp67_ASAP7_75t_L g660 ( 
.A(n_480),
.B(n_0),
.Y(n_660)
);

BUFx3_ASAP7_75t_L g661 ( 
.A(n_586),
.Y(n_661)
);

CKINVDCx20_ASAP7_75t_R g662 ( 
.A(n_556),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_500),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_503),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_511),
.Y(n_665)
);

INVxp33_ASAP7_75t_SL g666 ( 
.A(n_480),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_515),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_517),
.Y(n_668)
);

INVxp67_ASAP7_75t_SL g669 ( 
.A(n_550),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_522),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_524),
.Y(n_671)
);

CKINVDCx20_ASAP7_75t_R g672 ( 
.A(n_560),
.Y(n_672)
);

CKINVDCx5p33_ASAP7_75t_R g673 ( 
.A(n_442),
.Y(n_673)
);

INVxp67_ASAP7_75t_L g674 ( 
.A(n_494),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_526),
.Y(n_675)
);

INVxp67_ASAP7_75t_SL g676 ( 
.A(n_563),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_539),
.Y(n_677)
);

CKINVDCx5p33_ASAP7_75t_R g678 ( 
.A(n_444),
.Y(n_678)
);

CKINVDCx5p33_ASAP7_75t_R g679 ( 
.A(n_445),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_547),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_548),
.Y(n_681)
);

INVxp67_ASAP7_75t_SL g682 ( 
.A(n_563),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_552),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_554),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_555),
.Y(n_685)
);

INVx2_ASAP7_75t_L g686 ( 
.A(n_570),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_557),
.Y(n_687)
);

INVxp67_ASAP7_75t_L g688 ( 
.A(n_521),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_562),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_564),
.Y(n_690)
);

CKINVDCx20_ASAP7_75t_R g691 ( 
.A(n_609),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_572),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_574),
.Y(n_693)
);

CKINVDCx5p33_ASAP7_75t_R g694 ( 
.A(n_446),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_575),
.Y(n_695)
);

CKINVDCx5p33_ASAP7_75t_R g696 ( 
.A(n_448),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_589),
.Y(n_697)
);

INVxp67_ASAP7_75t_SL g698 ( 
.A(n_604),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_595),
.Y(n_699)
);

BUFx3_ASAP7_75t_L g700 ( 
.A(n_454),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_603),
.Y(n_701)
);

CKINVDCx5p33_ASAP7_75t_R g702 ( 
.A(n_449),
.Y(n_702)
);

INVxp67_ASAP7_75t_SL g703 ( 
.A(n_551),
.Y(n_703)
);

HB1xp67_ASAP7_75t_L g704 ( 
.A(n_545),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_610),
.Y(n_705)
);

INVxp33_ASAP7_75t_SL g706 ( 
.A(n_578),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_611),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_466),
.Y(n_708)
);

CKINVDCx5p33_ASAP7_75t_R g709 ( 
.A(n_450),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_601),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_459),
.Y(n_711)
);

CKINVDCx5p33_ASAP7_75t_R g712 ( 
.A(n_451),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_471),
.Y(n_713)
);

INVxp67_ASAP7_75t_SL g714 ( 
.A(n_551),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_491),
.Y(n_715)
);

AND2x4_ASAP7_75t_L g716 ( 
.A(n_700),
.B(n_464),
.Y(n_716)
);

BUFx6f_ASAP7_75t_L g717 ( 
.A(n_651),
.Y(n_717)
);

BUFx6f_ASAP7_75t_L g718 ( 
.A(n_651),
.Y(n_718)
);

AND2x4_ASAP7_75t_L g719 ( 
.A(n_669),
.B(n_489),
.Y(n_719)
);

HB1xp67_ASAP7_75t_L g720 ( 
.A(n_704),
.Y(n_720)
);

BUFx2_ASAP7_75t_L g721 ( 
.A(n_617),
.Y(n_721)
);

OAI21x1_ASAP7_75t_L g722 ( 
.A1(n_686),
.A2(n_561),
.B(n_549),
.Y(n_722)
);

BUFx2_ASAP7_75t_L g723 ( 
.A(n_644),
.Y(n_723)
);

BUFx6f_ASAP7_75t_L g724 ( 
.A(n_651),
.Y(n_724)
);

BUFx6f_ASAP7_75t_L g725 ( 
.A(n_651),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_627),
.Y(n_726)
);

INVx6_ASAP7_75t_L g727 ( 
.A(n_647),
.Y(n_727)
);

BUFx6f_ASAP7_75t_L g728 ( 
.A(n_616),
.Y(n_728)
);

BUFx6f_ASAP7_75t_L g729 ( 
.A(n_618),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_619),
.Y(n_730)
);

BUFx12f_ASAP7_75t_L g731 ( 
.A(n_621),
.Y(n_731)
);

CKINVDCx8_ASAP7_75t_R g732 ( 
.A(n_628),
.Y(n_732)
);

AND2x4_ASAP7_75t_L g733 ( 
.A(n_669),
.B(n_496),
.Y(n_733)
);

BUFx6f_ASAP7_75t_L g734 ( 
.A(n_620),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_L g735 ( 
.A(n_642),
.B(n_546),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_622),
.Y(n_736)
);

CKINVDCx5p33_ASAP7_75t_R g737 ( 
.A(n_673),
.Y(n_737)
);

AOI22xp5_ASAP7_75t_L g738 ( 
.A1(n_666),
.A2(n_566),
.B1(n_602),
.B2(n_599),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_678),
.B(n_479),
.Y(n_739)
);

OAI22xp5_ASAP7_75t_L g740 ( 
.A1(n_615),
.A2(n_591),
.B1(n_583),
.B2(n_597),
.Y(n_740)
);

INVx5_ASAP7_75t_L g741 ( 
.A(n_640),
.Y(n_741)
);

INVx5_ASAP7_75t_L g742 ( 
.A(n_640),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_623),
.Y(n_743)
);

HB1xp67_ASAP7_75t_L g744 ( 
.A(n_704),
.Y(n_744)
);

INVx2_ASAP7_75t_L g745 ( 
.A(n_625),
.Y(n_745)
);

OAI21x1_ASAP7_75t_L g746 ( 
.A1(n_703),
.A2(n_570),
.B(n_540),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_679),
.B(n_458),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_703),
.Y(n_748)
);

XNOR2xp5_ASAP7_75t_L g749 ( 
.A(n_614),
.B(n_504),
.Y(n_749)
);

CKINVDCx5p33_ASAP7_75t_R g750 ( 
.A(n_694),
.Y(n_750)
);

INVx2_ASAP7_75t_L g751 ( 
.A(n_629),
.Y(n_751)
);

BUFx6f_ASAP7_75t_L g752 ( 
.A(n_631),
.Y(n_752)
);

INVx3_ASAP7_75t_L g753 ( 
.A(n_632),
.Y(n_753)
);

BUFx6f_ASAP7_75t_L g754 ( 
.A(n_711),
.Y(n_754)
);

CKINVDCx5p33_ASAP7_75t_R g755 ( 
.A(n_696),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_L g756 ( 
.A(n_702),
.B(n_709),
.Y(n_756)
);

BUFx6f_ASAP7_75t_L g757 ( 
.A(n_713),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_714),
.Y(n_758)
);

OAI21x1_ASAP7_75t_L g759 ( 
.A1(n_714),
.A2(n_636),
.B(n_635),
.Y(n_759)
);

INVx2_ASAP7_75t_L g760 ( 
.A(n_715),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_712),
.B(n_460),
.Y(n_761)
);

AND2x4_ASAP7_75t_L g762 ( 
.A(n_661),
.B(n_568),
.Y(n_762)
);

BUFx6f_ASAP7_75t_L g763 ( 
.A(n_637),
.Y(n_763)
);

OAI21x1_ASAP7_75t_L g764 ( 
.A1(n_638),
.A2(n_570),
.B(n_465),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_639),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_645),
.Y(n_766)
);

AND2x2_ASAP7_75t_L g767 ( 
.A(n_674),
.B(n_594),
.Y(n_767)
);

AND2x4_ASAP7_75t_L g768 ( 
.A(n_674),
.B(n_688),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_L g769 ( 
.A(n_676),
.B(n_463),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_646),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_648),
.Y(n_771)
);

BUFx3_ASAP7_75t_L g772 ( 
.A(n_708),
.Y(n_772)
);

AND2x2_ASAP7_75t_L g773 ( 
.A(n_688),
.B(n_606),
.Y(n_773)
);

AOI22xp5_ASAP7_75t_L g774 ( 
.A1(n_633),
.A2(n_612),
.B1(n_542),
.B2(n_593),
.Y(n_774)
);

INVx2_ASAP7_75t_L g775 ( 
.A(n_650),
.Y(n_775)
);

BUFx2_ASAP7_75t_L g776 ( 
.A(n_626),
.Y(n_776)
);

INVx3_ASAP7_75t_L g777 ( 
.A(n_652),
.Y(n_777)
);

INVx2_ASAP7_75t_L g778 ( 
.A(n_654),
.Y(n_778)
);

AND2x4_ASAP7_75t_L g779 ( 
.A(n_698),
.B(n_551),
.Y(n_779)
);

INVx2_ASAP7_75t_L g780 ( 
.A(n_655),
.Y(n_780)
);

BUFx8_ASAP7_75t_L g781 ( 
.A(n_649),
.Y(n_781)
);

HB1xp67_ASAP7_75t_L g782 ( 
.A(n_630),
.Y(n_782)
);

INVx2_ASAP7_75t_L g783 ( 
.A(n_659),
.Y(n_783)
);

INVx3_ASAP7_75t_L g784 ( 
.A(n_663),
.Y(n_784)
);

AND2x2_ASAP7_75t_L g785 ( 
.A(n_698),
.B(n_470),
.Y(n_785)
);

CKINVDCx5p33_ASAP7_75t_R g786 ( 
.A(n_624),
.Y(n_786)
);

INVx2_ASAP7_75t_L g787 ( 
.A(n_664),
.Y(n_787)
);

INVx2_ASAP7_75t_L g788 ( 
.A(n_665),
.Y(n_788)
);

NOR2xp33_ASAP7_75t_L g789 ( 
.A(n_706),
.B(n_472),
.Y(n_789)
);

INVx2_ASAP7_75t_L g790 ( 
.A(n_667),
.Y(n_790)
);

INVx2_ASAP7_75t_L g791 ( 
.A(n_668),
.Y(n_791)
);

HB1xp67_ASAP7_75t_L g792 ( 
.A(n_615),
.Y(n_792)
);

INVx5_ASAP7_75t_L g793 ( 
.A(n_676),
.Y(n_793)
);

AOI22xp5_ASAP7_75t_L g794 ( 
.A1(n_660),
.A2(n_682),
.B1(n_643),
.B2(n_634),
.Y(n_794)
);

BUFx6f_ASAP7_75t_L g795 ( 
.A(n_670),
.Y(n_795)
);

INVx2_ASAP7_75t_L g796 ( 
.A(n_671),
.Y(n_796)
);

AND2x4_ASAP7_75t_L g797 ( 
.A(n_710),
.B(n_559),
.Y(n_797)
);

INVx2_ASAP7_75t_L g798 ( 
.A(n_707),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_L g799 ( 
.A(n_682),
.B(n_675),
.Y(n_799)
);

OAI22x1_ASAP7_75t_SL g800 ( 
.A1(n_641),
.A2(n_607),
.B1(n_477),
.B2(n_482),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_L g801 ( 
.A(n_677),
.B(n_613),
.Y(n_801)
);

INVx2_ASAP7_75t_L g802 ( 
.A(n_728),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_770),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_765),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_765),
.Y(n_805)
);

NAND2xp33_ASAP7_75t_L g806 ( 
.A(n_793),
.B(n_570),
.Y(n_806)
);

CKINVDCx5p33_ASAP7_75t_R g807 ( 
.A(n_786),
.Y(n_807)
);

INVx2_ASAP7_75t_L g808 ( 
.A(n_728),
.Y(n_808)
);

NAND2xp33_ASAP7_75t_SL g809 ( 
.A(n_767),
.B(n_559),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_766),
.Y(n_810)
);

BUFx3_ASAP7_75t_L g811 ( 
.A(n_748),
.Y(n_811)
);

HB1xp67_ASAP7_75t_L g812 ( 
.A(n_793),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_766),
.Y(n_813)
);

BUFx6f_ASAP7_75t_L g814 ( 
.A(n_717),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_771),
.Y(n_815)
);

INVx2_ASAP7_75t_L g816 ( 
.A(n_745),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_771),
.Y(n_817)
);

INVx3_ASAP7_75t_L g818 ( 
.A(n_717),
.Y(n_818)
);

AND2x2_ASAP7_75t_L g819 ( 
.A(n_793),
.B(n_634),
.Y(n_819)
);

BUFx6f_ASAP7_75t_L g820 ( 
.A(n_717),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_763),
.Y(n_821)
);

BUFx6f_ASAP7_75t_L g822 ( 
.A(n_718),
.Y(n_822)
);

INVx2_ASAP7_75t_L g823 ( 
.A(n_730),
.Y(n_823)
);

BUFx2_ASAP7_75t_L g824 ( 
.A(n_776),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_763),
.Y(n_825)
);

INVx2_ASAP7_75t_L g826 ( 
.A(n_730),
.Y(n_826)
);

BUFx6f_ASAP7_75t_L g827 ( 
.A(n_718),
.Y(n_827)
);

BUFx6f_ASAP7_75t_L g828 ( 
.A(n_718),
.Y(n_828)
);

INVx3_ASAP7_75t_L g829 ( 
.A(n_724),
.Y(n_829)
);

AND2x2_ASAP7_75t_L g830 ( 
.A(n_773),
.B(n_643),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_763),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_795),
.Y(n_832)
);

AND2x4_ASAP7_75t_L g833 ( 
.A(n_779),
.B(n_657),
.Y(n_833)
);

BUFx6f_ASAP7_75t_L g834 ( 
.A(n_724),
.Y(n_834)
);

BUFx6f_ASAP7_75t_L g835 ( 
.A(n_724),
.Y(n_835)
);

INVx2_ASAP7_75t_L g836 ( 
.A(n_726),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_795),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_758),
.B(n_680),
.Y(n_838)
);

AND3x2_ASAP7_75t_L g839 ( 
.A(n_720),
.B(n_658),
.C(n_656),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_795),
.Y(n_840)
);

INVx2_ASAP7_75t_L g841 ( 
.A(n_728),
.Y(n_841)
);

INVx3_ASAP7_75t_L g842 ( 
.A(n_725),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_775),
.Y(n_843)
);

OAI21x1_ASAP7_75t_L g844 ( 
.A1(n_759),
.A2(n_683),
.B(n_681),
.Y(n_844)
);

INVx2_ASAP7_75t_L g845 ( 
.A(n_729),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_778),
.Y(n_846)
);

BUFx3_ASAP7_75t_L g847 ( 
.A(n_727),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_780),
.Y(n_848)
);

AND2x4_ASAP7_75t_L g849 ( 
.A(n_779),
.B(n_657),
.Y(n_849)
);

INVxp67_ASAP7_75t_L g850 ( 
.A(n_792),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_783),
.Y(n_851)
);

AND2x2_ASAP7_75t_L g852 ( 
.A(n_785),
.B(n_656),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_L g853 ( 
.A(n_797),
.B(n_799),
.Y(n_853)
);

INVx2_ASAP7_75t_L g854 ( 
.A(n_729),
.Y(n_854)
);

INVx2_ASAP7_75t_L g855 ( 
.A(n_729),
.Y(n_855)
);

INVx2_ASAP7_75t_L g856 ( 
.A(n_734),
.Y(n_856)
);

INVx2_ASAP7_75t_L g857 ( 
.A(n_736),
.Y(n_857)
);

INVx2_ASAP7_75t_L g858 ( 
.A(n_743),
.Y(n_858)
);

INVx2_ASAP7_75t_L g859 ( 
.A(n_734),
.Y(n_859)
);

AND2x4_ASAP7_75t_L g860 ( 
.A(n_772),
.B(n_658),
.Y(n_860)
);

INVx2_ASAP7_75t_L g861 ( 
.A(n_734),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_787),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_788),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_797),
.B(n_684),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_790),
.Y(n_865)
);

INVx6_ASAP7_75t_L g866 ( 
.A(n_727),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_791),
.Y(n_867)
);

INVxp67_ASAP7_75t_L g868 ( 
.A(n_744),
.Y(n_868)
);

INVx2_ASAP7_75t_L g869 ( 
.A(n_725),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_796),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_798),
.Y(n_871)
);

BUFx6f_ASAP7_75t_L g872 ( 
.A(n_725),
.Y(n_872)
);

AND2x2_ASAP7_75t_L g873 ( 
.A(n_768),
.B(n_685),
.Y(n_873)
);

INVx3_ASAP7_75t_L g874 ( 
.A(n_754),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_752),
.Y(n_875)
);

INVx3_ASAP7_75t_L g876 ( 
.A(n_754),
.Y(n_876)
);

INVx2_ASAP7_75t_L g877 ( 
.A(n_760),
.Y(n_877)
);

AND2x2_ASAP7_75t_L g878 ( 
.A(n_768),
.B(n_687),
.Y(n_878)
);

INVx2_ASAP7_75t_L g879 ( 
.A(n_722),
.Y(n_879)
);

INVx2_ASAP7_75t_L g880 ( 
.A(n_751),
.Y(n_880)
);

BUFx6f_ASAP7_75t_L g881 ( 
.A(n_754),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_752),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_752),
.Y(n_883)
);

BUFx6f_ASAP7_75t_L g884 ( 
.A(n_757),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_777),
.Y(n_885)
);

INVx3_ASAP7_75t_L g886 ( 
.A(n_757),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_777),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_784),
.Y(n_888)
);

INVx2_ASAP7_75t_L g889 ( 
.A(n_757),
.Y(n_889)
);

INVx2_ASAP7_75t_L g890 ( 
.A(n_784),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_753),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_753),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_801),
.Y(n_893)
);

AND2x6_ASAP7_75t_L g894 ( 
.A(n_738),
.B(n_559),
.Y(n_894)
);

INVx3_ASAP7_75t_L g895 ( 
.A(n_746),
.Y(n_895)
);

NOR2xp33_ASAP7_75t_L g896 ( 
.A(n_893),
.B(n_756),
.Y(n_896)
);

AOI22xp33_ASAP7_75t_L g897 ( 
.A1(n_894),
.A2(n_719),
.B1(n_733),
.B2(n_769),
.Y(n_897)
);

NOR2xp33_ASAP7_75t_L g898 ( 
.A(n_850),
.B(n_737),
.Y(n_898)
);

INVx1_ASAP7_75t_SL g899 ( 
.A(n_824),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_SL g900 ( 
.A(n_833),
.B(n_732),
.Y(n_900)
);

INVx2_ASAP7_75t_L g901 ( 
.A(n_880),
.Y(n_901)
);

AOI22xp5_ASAP7_75t_L g902 ( 
.A1(n_830),
.A2(n_739),
.B1(n_733),
.B2(n_719),
.Y(n_902)
);

AOI22xp33_ASAP7_75t_L g903 ( 
.A1(n_894),
.A2(n_794),
.B1(n_740),
.B2(n_716),
.Y(n_903)
);

INVxp67_ASAP7_75t_SL g904 ( 
.A(n_814),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_804),
.Y(n_905)
);

AND2x6_ASAP7_75t_L g906 ( 
.A(n_895),
.B(n_762),
.Y(n_906)
);

INVx2_ASAP7_75t_L g907 ( 
.A(n_880),
.Y(n_907)
);

INVx2_ASAP7_75t_L g908 ( 
.A(n_823),
.Y(n_908)
);

INVx2_ASAP7_75t_L g909 ( 
.A(n_823),
.Y(n_909)
);

BUFx3_ASAP7_75t_L g910 ( 
.A(n_847),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_805),
.Y(n_911)
);

CKINVDCx5p33_ASAP7_75t_R g912 ( 
.A(n_807),
.Y(n_912)
);

INVx3_ASAP7_75t_L g913 ( 
.A(n_890),
.Y(n_913)
);

CKINVDCx20_ASAP7_75t_R g914 ( 
.A(n_807),
.Y(n_914)
);

INVx4_ASAP7_75t_L g915 ( 
.A(n_881),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_810),
.Y(n_916)
);

CKINVDCx6p67_ASAP7_75t_R g917 ( 
.A(n_847),
.Y(n_917)
);

INVx2_ASAP7_75t_L g918 ( 
.A(n_826),
.Y(n_918)
);

BUFx6f_ASAP7_75t_L g919 ( 
.A(n_814),
.Y(n_919)
);

BUFx8_ASAP7_75t_SL g920 ( 
.A(n_860),
.Y(n_920)
);

INVx2_ASAP7_75t_L g921 ( 
.A(n_826),
.Y(n_921)
);

AND3x1_ASAP7_75t_L g922 ( 
.A(n_852),
.B(n_774),
.C(n_782),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_L g923 ( 
.A(n_833),
.B(n_735),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_813),
.Y(n_924)
);

INVx2_ASAP7_75t_L g925 ( 
.A(n_877),
.Y(n_925)
);

INVx2_ASAP7_75t_L g926 ( 
.A(n_877),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_815),
.Y(n_927)
);

BUFx4f_ASAP7_75t_L g928 ( 
.A(n_894),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_SL g929 ( 
.A(n_849),
.B(n_762),
.Y(n_929)
);

AND2x2_ASAP7_75t_L g930 ( 
.A(n_819),
.B(n_716),
.Y(n_930)
);

INVx6_ASAP7_75t_L g931 ( 
.A(n_866),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_L g932 ( 
.A(n_849),
.B(n_789),
.Y(n_932)
);

OR2x2_ASAP7_75t_L g933 ( 
.A(n_850),
.B(n_749),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_L g934 ( 
.A(n_853),
.B(n_747),
.Y(n_934)
);

INVx3_ASAP7_75t_L g935 ( 
.A(n_836),
.Y(n_935)
);

AND2x6_ASAP7_75t_L g936 ( 
.A(n_895),
.B(n_559),
.Y(n_936)
);

AND2x2_ASAP7_75t_L g937 ( 
.A(n_860),
.B(n_812),
.Y(n_937)
);

AND2x6_ASAP7_75t_L g938 ( 
.A(n_879),
.B(n_761),
.Y(n_938)
);

INVxp67_ASAP7_75t_L g939 ( 
.A(n_873),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_817),
.Y(n_940)
);

BUFx3_ASAP7_75t_L g941 ( 
.A(n_866),
.Y(n_941)
);

XOR2xp5_ASAP7_75t_L g942 ( 
.A(n_812),
.B(n_653),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_803),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_SL g944 ( 
.A(n_878),
.B(n_750),
.Y(n_944)
);

OR2x6_ASAP7_75t_L g945 ( 
.A(n_866),
.B(n_731),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_836),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_885),
.Y(n_947)
);

BUFx3_ASAP7_75t_L g948 ( 
.A(n_811),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_887),
.Y(n_949)
);

INVx2_ASAP7_75t_L g950 ( 
.A(n_816),
.Y(n_950)
);

BUFx2_ASAP7_75t_L g951 ( 
.A(n_868),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_888),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_SL g953 ( 
.A(n_853),
.B(n_755),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_L g954 ( 
.A(n_811),
.B(n_689),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_SL g955 ( 
.A(n_809),
.B(n_721),
.Y(n_955)
);

INVx2_ASAP7_75t_L g956 ( 
.A(n_816),
.Y(n_956)
);

BUFx6f_ASAP7_75t_L g957 ( 
.A(n_814),
.Y(n_957)
);

INVx3_ASAP7_75t_R g958 ( 
.A(n_857),
.Y(n_958)
);

INVx2_ASAP7_75t_L g959 ( 
.A(n_857),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_L g960 ( 
.A(n_891),
.B(n_690),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_L g961 ( 
.A(n_892),
.B(n_692),
.Y(n_961)
);

AOI22xp33_ASAP7_75t_L g962 ( 
.A1(n_894),
.A2(n_570),
.B1(n_764),
.B2(n_695),
.Y(n_962)
);

INVx4_ASAP7_75t_SL g963 ( 
.A(n_894),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_L g964 ( 
.A(n_838),
.B(n_693),
.Y(n_964)
);

INVx1_ASAP7_75t_L g965 ( 
.A(n_858),
.Y(n_965)
);

INVx2_ASAP7_75t_L g966 ( 
.A(n_858),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_L g967 ( 
.A(n_838),
.B(n_697),
.Y(n_967)
);

NAND2xp33_ASAP7_75t_SL g968 ( 
.A(n_864),
.B(n_662),
.Y(n_968)
);

INVx3_ASAP7_75t_L g969 ( 
.A(n_859),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_SL g970 ( 
.A(n_809),
.B(n_723),
.Y(n_970)
);

INVx3_ASAP7_75t_L g971 ( 
.A(n_859),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_SL g972 ( 
.A(n_868),
.B(n_781),
.Y(n_972)
);

AND2x2_ASAP7_75t_L g973 ( 
.A(n_864),
.B(n_843),
.Y(n_973)
);

OR2x2_ASAP7_75t_L g974 ( 
.A(n_846),
.B(n_699),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_848),
.Y(n_975)
);

AOI22xp33_ASAP7_75t_L g976 ( 
.A1(n_844),
.A2(n_570),
.B1(n_705),
.B2(n_701),
.Y(n_976)
);

BUFx6f_ASAP7_75t_L g977 ( 
.A(n_814),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_L g978 ( 
.A(n_861),
.B(n_476),
.Y(n_978)
);

BUFx10_ASAP7_75t_L g979 ( 
.A(n_839),
.Y(n_979)
);

AOI22xp33_ASAP7_75t_L g980 ( 
.A1(n_806),
.A2(n_487),
.B1(n_492),
.B2(n_486),
.Y(n_980)
);

INVx2_ASAP7_75t_SL g981 ( 
.A(n_839),
.Y(n_981)
);

AND3x2_ASAP7_75t_L g982 ( 
.A(n_851),
.B(n_800),
.C(n_781),
.Y(n_982)
);

BUFx6f_ASAP7_75t_SL g983 ( 
.A(n_862),
.Y(n_983)
);

BUFx4f_ASAP7_75t_L g984 ( 
.A(n_881),
.Y(n_984)
);

NOR2x1p5_ASAP7_75t_L g985 ( 
.A(n_863),
.B(n_493),
.Y(n_985)
);

INVx4_ASAP7_75t_L g986 ( 
.A(n_881),
.Y(n_986)
);

AND2x2_ASAP7_75t_L g987 ( 
.A(n_865),
.B(n_672),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_SL g988 ( 
.A(n_881),
.B(n_691),
.Y(n_988)
);

INVx4_ASAP7_75t_L g989 ( 
.A(n_884),
.Y(n_989)
);

INVx3_ASAP7_75t_L g990 ( 
.A(n_861),
.Y(n_990)
);

CKINVDCx5p33_ASAP7_75t_R g991 ( 
.A(n_889),
.Y(n_991)
);

AOI22xp33_ASAP7_75t_L g992 ( 
.A1(n_806),
.A2(n_499),
.B1(n_501),
.B2(n_497),
.Y(n_992)
);

OR2x6_ASAP7_75t_L g993 ( 
.A(n_867),
.B(n_870),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_SL g994 ( 
.A(n_884),
.B(n_505),
.Y(n_994)
);

HB1xp67_ASAP7_75t_L g995 ( 
.A(n_899),
.Y(n_995)
);

INVx1_ASAP7_75t_L g996 ( 
.A(n_908),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_909),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_L g998 ( 
.A(n_934),
.B(n_871),
.Y(n_998)
);

INVxp33_ASAP7_75t_L g999 ( 
.A(n_951),
.Y(n_999)
);

NOR2xp33_ASAP7_75t_L g1000 ( 
.A(n_896),
.B(n_932),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_L g1001 ( 
.A(n_923),
.B(n_874),
.Y(n_1001)
);

INVx1_ASAP7_75t_L g1002 ( 
.A(n_918),
.Y(n_1002)
);

AND2x4_ASAP7_75t_L g1003 ( 
.A(n_948),
.B(n_821),
.Y(n_1003)
);

BUFx3_ASAP7_75t_L g1004 ( 
.A(n_910),
.Y(n_1004)
);

INVx1_ASAP7_75t_L g1005 ( 
.A(n_921),
.Y(n_1005)
);

INVx2_ASAP7_75t_L g1006 ( 
.A(n_935),
.Y(n_1006)
);

NOR2xp33_ASAP7_75t_L g1007 ( 
.A(n_898),
.B(n_825),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_L g1008 ( 
.A(n_973),
.B(n_874),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_L g1009 ( 
.A(n_930),
.B(n_876),
.Y(n_1009)
);

INVx2_ASAP7_75t_L g1010 ( 
.A(n_935),
.Y(n_1010)
);

INVx2_ASAP7_75t_L g1011 ( 
.A(n_901),
.Y(n_1011)
);

AND2x2_ASAP7_75t_L g1012 ( 
.A(n_937),
.B(n_831),
.Y(n_1012)
);

AND2x6_ASAP7_75t_L g1013 ( 
.A(n_902),
.B(n_879),
.Y(n_1013)
);

INVx2_ASAP7_75t_L g1014 ( 
.A(n_907),
.Y(n_1014)
);

A2O1A1Ixp33_ASAP7_75t_L g1015 ( 
.A1(n_897),
.A2(n_837),
.B(n_840),
.C(n_832),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_SL g1016 ( 
.A(n_903),
.B(n_875),
.Y(n_1016)
);

AOI22xp5_ASAP7_75t_L g1017 ( 
.A1(n_906),
.A2(n_883),
.B1(n_882),
.B2(n_808),
.Y(n_1017)
);

INVx2_ASAP7_75t_L g1018 ( 
.A(n_925),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_SL g1019 ( 
.A(n_929),
.B(n_884),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_L g1020 ( 
.A(n_964),
.B(n_876),
.Y(n_1020)
);

AOI22xp33_ASAP7_75t_L g1021 ( 
.A1(n_906),
.A2(n_841),
.B1(n_845),
.B2(n_802),
.Y(n_1021)
);

INVx2_ASAP7_75t_L g1022 ( 
.A(n_926),
.Y(n_1022)
);

INVx2_ASAP7_75t_L g1023 ( 
.A(n_950),
.Y(n_1023)
);

OAI22xp5_ASAP7_75t_L g1024 ( 
.A1(n_928),
.A2(n_886),
.B1(n_869),
.B2(n_855),
.Y(n_1024)
);

OAI22xp5_ASAP7_75t_L g1025 ( 
.A1(n_928),
.A2(n_886),
.B1(n_856),
.B2(n_854),
.Y(n_1025)
);

OAI22xp33_ASAP7_75t_L g1026 ( 
.A1(n_939),
.A2(n_884),
.B1(n_507),
.B2(n_509),
.Y(n_1026)
);

INVx2_ASAP7_75t_SL g1027 ( 
.A(n_931),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_SL g1028 ( 
.A(n_953),
.B(n_820),
.Y(n_1028)
);

NAND2xp5_ASAP7_75t_L g1029 ( 
.A(n_967),
.B(n_818),
.Y(n_1029)
);

INVx2_ASAP7_75t_L g1030 ( 
.A(n_956),
.Y(n_1030)
);

INVx2_ASAP7_75t_SL g1031 ( 
.A(n_931),
.Y(n_1031)
);

CKINVDCx5p33_ASAP7_75t_R g1032 ( 
.A(n_912),
.Y(n_1032)
);

NAND2xp5_ASAP7_75t_SL g1033 ( 
.A(n_900),
.B(n_820),
.Y(n_1033)
);

INVx2_ASAP7_75t_SL g1034 ( 
.A(n_987),
.Y(n_1034)
);

NOR2xp67_ASAP7_75t_L g1035 ( 
.A(n_933),
.B(n_913),
.Y(n_1035)
);

AOI22xp33_ASAP7_75t_L g1036 ( 
.A1(n_906),
.A2(n_829),
.B1(n_842),
.B2(n_818),
.Y(n_1036)
);

INVx2_ASAP7_75t_SL g1037 ( 
.A(n_974),
.Y(n_1037)
);

NAND3xp33_ASAP7_75t_L g1038 ( 
.A(n_968),
.B(n_510),
.C(n_506),
.Y(n_1038)
);

NAND2xp5_ASAP7_75t_L g1039 ( 
.A(n_938),
.B(n_829),
.Y(n_1039)
);

NOR2xp67_ASAP7_75t_L g1040 ( 
.A(n_913),
.B(n_842),
.Y(n_1040)
);

INVx2_ASAP7_75t_L g1041 ( 
.A(n_959),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_L g1042 ( 
.A(n_938),
.B(n_820),
.Y(n_1042)
);

NAND2xp5_ASAP7_75t_L g1043 ( 
.A(n_905),
.B(n_820),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_L g1044 ( 
.A(n_911),
.B(n_822),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_L g1045 ( 
.A(n_916),
.B(n_822),
.Y(n_1045)
);

INVx1_ASAP7_75t_L g1046 ( 
.A(n_924),
.Y(n_1046)
);

NAND2xp5_ASAP7_75t_L g1047 ( 
.A(n_927),
.B(n_822),
.Y(n_1047)
);

INVx2_ASAP7_75t_L g1048 ( 
.A(n_966),
.Y(n_1048)
);

NOR2xp33_ASAP7_75t_L g1049 ( 
.A(n_944),
.B(n_822),
.Y(n_1049)
);

NAND2xp5_ASAP7_75t_L g1050 ( 
.A(n_940),
.B(n_827),
.Y(n_1050)
);

INVx1_ASAP7_75t_L g1051 ( 
.A(n_965),
.Y(n_1051)
);

NOR2xp33_ASAP7_75t_L g1052 ( 
.A(n_981),
.B(n_827),
.Y(n_1052)
);

INVx2_ASAP7_75t_L g1053 ( 
.A(n_969),
.Y(n_1053)
);

AND2x2_ASAP7_75t_L g1054 ( 
.A(n_917),
.B(n_741),
.Y(n_1054)
);

NOR2xp33_ASAP7_75t_L g1055 ( 
.A(n_991),
.B(n_827),
.Y(n_1055)
);

INVx1_ASAP7_75t_SL g1056 ( 
.A(n_914),
.Y(n_1056)
);

AND2x2_ASAP7_75t_L g1057 ( 
.A(n_941),
.B(n_741),
.Y(n_1057)
);

INVx2_ASAP7_75t_L g1058 ( 
.A(n_969),
.Y(n_1058)
);

OR2x2_ASAP7_75t_L g1059 ( 
.A(n_988),
.B(n_512),
.Y(n_1059)
);

NAND2xp5_ASAP7_75t_L g1060 ( 
.A(n_938),
.B(n_827),
.Y(n_1060)
);

AND2x4_ASAP7_75t_SL g1061 ( 
.A(n_945),
.B(n_828),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_L g1062 ( 
.A(n_938),
.B(n_828),
.Y(n_1062)
);

NAND2xp5_ASAP7_75t_L g1063 ( 
.A(n_906),
.B(n_828),
.Y(n_1063)
);

INVx1_ASAP7_75t_L g1064 ( 
.A(n_946),
.Y(n_1064)
);

NAND2xp5_ASAP7_75t_L g1065 ( 
.A(n_943),
.B(n_828),
.Y(n_1065)
);

NOR2xp33_ASAP7_75t_L g1066 ( 
.A(n_942),
.B(n_834),
.Y(n_1066)
);

NAND3x1_ASAP7_75t_L g1067 ( 
.A(n_982),
.B(n_0),
.C(n_1),
.Y(n_1067)
);

NAND2xp5_ASAP7_75t_SL g1068 ( 
.A(n_984),
.B(n_834),
.Y(n_1068)
);

INVx2_ASAP7_75t_L g1069 ( 
.A(n_971),
.Y(n_1069)
);

INVx1_ASAP7_75t_L g1070 ( 
.A(n_947),
.Y(n_1070)
);

INVx2_ASAP7_75t_L g1071 ( 
.A(n_971),
.Y(n_1071)
);

NOR3xp33_ASAP7_75t_SL g1072 ( 
.A(n_1066),
.B(n_972),
.C(n_970),
.Y(n_1072)
);

BUFx3_ASAP7_75t_L g1073 ( 
.A(n_1004),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_L g1074 ( 
.A(n_1000),
.B(n_954),
.Y(n_1074)
);

NAND2xp5_ASAP7_75t_L g1075 ( 
.A(n_998),
.B(n_949),
.Y(n_1075)
);

AND2x2_ASAP7_75t_SL g1076 ( 
.A(n_1061),
.B(n_922),
.Y(n_1076)
);

AOI22xp33_ASAP7_75t_L g1077 ( 
.A1(n_1013),
.A2(n_952),
.B1(n_975),
.B2(n_985),
.Y(n_1077)
);

INVx1_ASAP7_75t_L g1078 ( 
.A(n_1046),
.Y(n_1078)
);

INVx1_ASAP7_75t_L g1079 ( 
.A(n_1051),
.Y(n_1079)
);

INVx1_ASAP7_75t_L g1080 ( 
.A(n_1064),
.Y(n_1080)
);

NOR2xp33_ASAP7_75t_L g1081 ( 
.A(n_999),
.B(n_955),
.Y(n_1081)
);

NAND2xp5_ASAP7_75t_L g1082 ( 
.A(n_998),
.B(n_960),
.Y(n_1082)
);

NAND2xp5_ASAP7_75t_L g1083 ( 
.A(n_1007),
.B(n_961),
.Y(n_1083)
);

NAND2xp5_ASAP7_75t_L g1084 ( 
.A(n_1008),
.B(n_990),
.Y(n_1084)
);

INVx2_ASAP7_75t_L g1085 ( 
.A(n_1006),
.Y(n_1085)
);

BUFx3_ASAP7_75t_L g1086 ( 
.A(n_1032),
.Y(n_1086)
);

NAND2xp5_ASAP7_75t_L g1087 ( 
.A(n_1008),
.B(n_990),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_L g1088 ( 
.A(n_1001),
.B(n_963),
.Y(n_1088)
);

NAND2xp5_ASAP7_75t_L g1089 ( 
.A(n_1001),
.B(n_963),
.Y(n_1089)
);

INVx1_ASAP7_75t_L g1090 ( 
.A(n_1070),
.Y(n_1090)
);

OR2x6_ASAP7_75t_L g1091 ( 
.A(n_995),
.B(n_945),
.Y(n_1091)
);

INVx1_ASAP7_75t_L g1092 ( 
.A(n_996),
.Y(n_1092)
);

INVxp67_ASAP7_75t_SL g1093 ( 
.A(n_1055),
.Y(n_1093)
);

NAND2xp5_ASAP7_75t_SL g1094 ( 
.A(n_1035),
.B(n_979),
.Y(n_1094)
);

AOI22xp33_ASAP7_75t_L g1095 ( 
.A1(n_1013),
.A2(n_993),
.B1(n_978),
.B2(n_994),
.Y(n_1095)
);

INVx2_ASAP7_75t_SL g1096 ( 
.A(n_1034),
.Y(n_1096)
);

BUFx6f_ASAP7_75t_L g1097 ( 
.A(n_1003),
.Y(n_1097)
);

AOI22xp33_ASAP7_75t_L g1098 ( 
.A1(n_1013),
.A2(n_993),
.B1(n_983),
.B2(n_992),
.Y(n_1098)
);

INVx1_ASAP7_75t_L g1099 ( 
.A(n_997),
.Y(n_1099)
);

NAND2xp5_ASAP7_75t_L g1100 ( 
.A(n_1020),
.B(n_915),
.Y(n_1100)
);

AOI22xp5_ASAP7_75t_L g1101 ( 
.A1(n_1016),
.A2(n_983),
.B1(n_976),
.B2(n_936),
.Y(n_1101)
);

INVx1_ASAP7_75t_L g1102 ( 
.A(n_1002),
.Y(n_1102)
);

INVx1_ASAP7_75t_L g1103 ( 
.A(n_1005),
.Y(n_1103)
);

NAND2xp5_ASAP7_75t_SL g1104 ( 
.A(n_1037),
.B(n_979),
.Y(n_1104)
);

NAND2xp5_ASAP7_75t_L g1105 ( 
.A(n_1020),
.B(n_915),
.Y(n_1105)
);

AOI22xp33_ASAP7_75t_L g1106 ( 
.A1(n_1013),
.A2(n_980),
.B1(n_962),
.B2(n_936),
.Y(n_1106)
);

BUFx4f_ASAP7_75t_L g1107 ( 
.A(n_1027),
.Y(n_1107)
);

CKINVDCx5p33_ASAP7_75t_R g1108 ( 
.A(n_1056),
.Y(n_1108)
);

INVx1_ASAP7_75t_L g1109 ( 
.A(n_1011),
.Y(n_1109)
);

NAND2xp5_ASAP7_75t_L g1110 ( 
.A(n_1029),
.B(n_986),
.Y(n_1110)
);

INVx1_ASAP7_75t_L g1111 ( 
.A(n_1014),
.Y(n_1111)
);

AND2x2_ASAP7_75t_L g1112 ( 
.A(n_1012),
.B(n_741),
.Y(n_1112)
);

INVx1_ASAP7_75t_L g1113 ( 
.A(n_1018),
.Y(n_1113)
);

INVx1_ASAP7_75t_L g1114 ( 
.A(n_1022),
.Y(n_1114)
);

NAND2xp5_ASAP7_75t_SL g1115 ( 
.A(n_1009),
.B(n_984),
.Y(n_1115)
);

NAND2xp5_ASAP7_75t_L g1116 ( 
.A(n_1029),
.B(n_1049),
.Y(n_1116)
);

NOR2xp33_ASAP7_75t_R g1117 ( 
.A(n_1056),
.B(n_919),
.Y(n_1117)
);

INVx3_ASAP7_75t_L g1118 ( 
.A(n_1010),
.Y(n_1118)
);

INVx4_ASAP7_75t_L g1119 ( 
.A(n_1003),
.Y(n_1119)
);

AND2x2_ASAP7_75t_SL g1120 ( 
.A(n_1059),
.B(n_986),
.Y(n_1120)
);

INVx2_ASAP7_75t_L g1121 ( 
.A(n_1023),
.Y(n_1121)
);

NOR3xp33_ASAP7_75t_L g1122 ( 
.A(n_1033),
.B(n_1038),
.C(n_1026),
.Y(n_1122)
);

BUFx3_ASAP7_75t_L g1123 ( 
.A(n_1031),
.Y(n_1123)
);

AOI22xp5_ASAP7_75t_L g1124 ( 
.A1(n_1041),
.A2(n_936),
.B1(n_514),
.B2(n_516),
.Y(n_1124)
);

NAND2xp5_ASAP7_75t_L g1125 ( 
.A(n_1052),
.B(n_989),
.Y(n_1125)
);

INVx1_ASAP7_75t_L g1126 ( 
.A(n_1030),
.Y(n_1126)
);

INVx3_ASAP7_75t_L g1127 ( 
.A(n_1053),
.Y(n_1127)
);

AOI22xp33_ASAP7_75t_SL g1128 ( 
.A1(n_1054),
.A2(n_936),
.B1(n_518),
.B2(n_519),
.Y(n_1128)
);

INVx1_ASAP7_75t_L g1129 ( 
.A(n_1048),
.Y(n_1129)
);

INVx2_ASAP7_75t_L g1130 ( 
.A(n_1058),
.Y(n_1130)
);

NAND2xp5_ASAP7_75t_L g1131 ( 
.A(n_1065),
.B(n_904),
.Y(n_1131)
);

NAND2xp5_ASAP7_75t_L g1132 ( 
.A(n_1065),
.B(n_989),
.Y(n_1132)
);

AND2x4_ASAP7_75t_L g1133 ( 
.A(n_1057),
.B(n_919),
.Y(n_1133)
);

INVx2_ASAP7_75t_L g1134 ( 
.A(n_1069),
.Y(n_1134)
);

INVx2_ASAP7_75t_L g1135 ( 
.A(n_1071),
.Y(n_1135)
);

INVx1_ASAP7_75t_L g1136 ( 
.A(n_1043),
.Y(n_1136)
);

AOI22xp33_ASAP7_75t_L g1137 ( 
.A1(n_1019),
.A2(n_957),
.B1(n_977),
.B2(n_919),
.Y(n_1137)
);

NAND2xp5_ASAP7_75t_L g1138 ( 
.A(n_1044),
.B(n_957),
.Y(n_1138)
);

INVx2_ASAP7_75t_L g1139 ( 
.A(n_1045),
.Y(n_1139)
);

INVx5_ASAP7_75t_L g1140 ( 
.A(n_1068),
.Y(n_1140)
);

INVx1_ASAP7_75t_L g1141 ( 
.A(n_1078),
.Y(n_1141)
);

NAND2xp5_ASAP7_75t_L g1142 ( 
.A(n_1082),
.B(n_1047),
.Y(n_1142)
);

NAND2xp5_ASAP7_75t_L g1143 ( 
.A(n_1074),
.B(n_1050),
.Y(n_1143)
);

NAND2xp5_ASAP7_75t_L g1144 ( 
.A(n_1075),
.B(n_1015),
.Y(n_1144)
);

INVx1_ASAP7_75t_L g1145 ( 
.A(n_1090),
.Y(n_1145)
);

INVx2_ASAP7_75t_L g1146 ( 
.A(n_1079),
.Y(n_1146)
);

OAI22xp5_ASAP7_75t_L g1147 ( 
.A1(n_1075),
.A2(n_1083),
.B1(n_1106),
.B2(n_1093),
.Y(n_1147)
);

INVx3_ASAP7_75t_L g1148 ( 
.A(n_1118),
.Y(n_1148)
);

AO22x1_ASAP7_75t_L g1149 ( 
.A1(n_1108),
.A2(n_1067),
.B1(n_920),
.B2(n_1039),
.Y(n_1149)
);

NOR2xp67_ASAP7_75t_L g1150 ( 
.A(n_1096),
.B(n_1028),
.Y(n_1150)
);

INVx2_ASAP7_75t_L g1151 ( 
.A(n_1080),
.Y(n_1151)
);

BUFx2_ASAP7_75t_L g1152 ( 
.A(n_1117),
.Y(n_1152)
);

NAND2xp33_ASAP7_75t_L g1153 ( 
.A(n_1122),
.B(n_1063),
.Y(n_1153)
);

INVx2_ASAP7_75t_L g1154 ( 
.A(n_1092),
.Y(n_1154)
);

CKINVDCx20_ASAP7_75t_R g1155 ( 
.A(n_1086),
.Y(n_1155)
);

NAND2xp5_ASAP7_75t_L g1156 ( 
.A(n_1116),
.B(n_1042),
.Y(n_1156)
);

INVx3_ASAP7_75t_L g1157 ( 
.A(n_1118),
.Y(n_1157)
);

NAND2xp5_ASAP7_75t_SL g1158 ( 
.A(n_1120),
.B(n_1040),
.Y(n_1158)
);

INVx2_ASAP7_75t_L g1159 ( 
.A(n_1099),
.Y(n_1159)
);

NAND2xp5_ASAP7_75t_L g1160 ( 
.A(n_1136),
.B(n_1042),
.Y(n_1160)
);

AND2x2_ASAP7_75t_L g1161 ( 
.A(n_1112),
.B(n_742),
.Y(n_1161)
);

INVx1_ASAP7_75t_L g1162 ( 
.A(n_1102),
.Y(n_1162)
);

BUFx4f_ASAP7_75t_L g1163 ( 
.A(n_1091),
.Y(n_1163)
);

INVx2_ASAP7_75t_L g1164 ( 
.A(n_1103),
.Y(n_1164)
);

NAND2xp5_ASAP7_75t_L g1165 ( 
.A(n_1139),
.B(n_1021),
.Y(n_1165)
);

AND2x4_ASAP7_75t_L g1166 ( 
.A(n_1133),
.B(n_1119),
.Y(n_1166)
);

BUFx2_ASAP7_75t_L g1167 ( 
.A(n_1073),
.Y(n_1167)
);

CKINVDCx5p33_ASAP7_75t_R g1168 ( 
.A(n_1123),
.Y(n_1168)
);

CKINVDCx5p33_ASAP7_75t_R g1169 ( 
.A(n_1091),
.Y(n_1169)
);

BUFx3_ASAP7_75t_L g1170 ( 
.A(n_1107),
.Y(n_1170)
);

INVxp67_ASAP7_75t_L g1171 ( 
.A(n_1081),
.Y(n_1171)
);

HB1xp67_ASAP7_75t_L g1172 ( 
.A(n_1097),
.Y(n_1172)
);

INVx1_ASAP7_75t_L g1173 ( 
.A(n_1109),
.Y(n_1173)
);

INVx3_ASAP7_75t_L g1174 ( 
.A(n_1127),
.Y(n_1174)
);

INVx2_ASAP7_75t_SL g1175 ( 
.A(n_1107),
.Y(n_1175)
);

INVx1_ASAP7_75t_L g1176 ( 
.A(n_1111),
.Y(n_1176)
);

CKINVDCx16_ASAP7_75t_R g1177 ( 
.A(n_1091),
.Y(n_1177)
);

NAND2xp5_ASAP7_75t_L g1178 ( 
.A(n_1131),
.B(n_1060),
.Y(n_1178)
);

INVxp33_ASAP7_75t_L g1179 ( 
.A(n_1097),
.Y(n_1179)
);

BUFx3_ASAP7_75t_L g1180 ( 
.A(n_1097),
.Y(n_1180)
);

INVx1_ASAP7_75t_L g1181 ( 
.A(n_1113),
.Y(n_1181)
);

NAND2xp5_ASAP7_75t_SL g1182 ( 
.A(n_1119),
.B(n_1017),
.Y(n_1182)
);

INVx1_ASAP7_75t_L g1183 ( 
.A(n_1114),
.Y(n_1183)
);

BUFx12f_ASAP7_75t_L g1184 ( 
.A(n_1076),
.Y(n_1184)
);

NAND2xp5_ASAP7_75t_L g1185 ( 
.A(n_1131),
.B(n_1060),
.Y(n_1185)
);

AOI221xp5_ASAP7_75t_L g1186 ( 
.A1(n_1072),
.A2(n_1025),
.B1(n_1024),
.B2(n_1039),
.C(n_523),
.Y(n_1186)
);

NAND2xp5_ASAP7_75t_SL g1187 ( 
.A(n_1098),
.B(n_1063),
.Y(n_1187)
);

AOI221xp5_ASAP7_75t_L g1188 ( 
.A1(n_1104),
.A2(n_1025),
.B1(n_1024),
.B2(n_525),
.C(n_528),
.Y(n_1188)
);

BUFx6f_ASAP7_75t_L g1189 ( 
.A(n_1133),
.Y(n_1189)
);

INVx2_ASAP7_75t_L g1190 ( 
.A(n_1121),
.Y(n_1190)
);

CKINVDCx5p33_ASAP7_75t_R g1191 ( 
.A(n_1094),
.Y(n_1191)
);

INVx2_ASAP7_75t_L g1192 ( 
.A(n_1126),
.Y(n_1192)
);

INVx2_ASAP7_75t_L g1193 ( 
.A(n_1129),
.Y(n_1193)
);

NOR2xp33_ASAP7_75t_R g1194 ( 
.A(n_1127),
.B(n_1062),
.Y(n_1194)
);

INVx1_ASAP7_75t_L g1195 ( 
.A(n_1085),
.Y(n_1195)
);

AND2x2_ASAP7_75t_L g1196 ( 
.A(n_1130),
.B(n_742),
.Y(n_1196)
);

INVx2_ASAP7_75t_L g1197 ( 
.A(n_1134),
.Y(n_1197)
);

NAND2xp5_ASAP7_75t_SL g1198 ( 
.A(n_1077),
.B(n_1062),
.Y(n_1198)
);

INVx1_ASAP7_75t_L g1199 ( 
.A(n_1135),
.Y(n_1199)
);

NAND2xp5_ASAP7_75t_L g1200 ( 
.A(n_1100),
.B(n_1036),
.Y(n_1200)
);

BUFx4f_ASAP7_75t_L g1201 ( 
.A(n_1140),
.Y(n_1201)
);

NOR2xp33_ASAP7_75t_L g1202 ( 
.A(n_1115),
.B(n_958),
.Y(n_1202)
);

INVx1_ASAP7_75t_SL g1203 ( 
.A(n_1138),
.Y(n_1203)
);

BUFx2_ASAP7_75t_L g1204 ( 
.A(n_1140),
.Y(n_1204)
);

BUFx6f_ASAP7_75t_L g1205 ( 
.A(n_1140),
.Y(n_1205)
);

NAND2xp5_ASAP7_75t_L g1206 ( 
.A(n_1105),
.B(n_957),
.Y(n_1206)
);

CKINVDCx20_ASAP7_75t_R g1207 ( 
.A(n_1101),
.Y(n_1207)
);

OAI21x1_ASAP7_75t_L g1208 ( 
.A1(n_1206),
.A2(n_1087),
.B(n_1084),
.Y(n_1208)
);

NAND2xp5_ASAP7_75t_L g1209 ( 
.A(n_1171),
.B(n_1095),
.Y(n_1209)
);

OAI21x1_ASAP7_75t_L g1210 ( 
.A1(n_1206),
.A2(n_1144),
.B(n_1156),
.Y(n_1210)
);

AOI21xp5_ASAP7_75t_L g1211 ( 
.A1(n_1142),
.A2(n_1153),
.B(n_1144),
.Y(n_1211)
);

INVx2_ASAP7_75t_L g1212 ( 
.A(n_1146),
.Y(n_1212)
);

NAND2xp5_ASAP7_75t_L g1213 ( 
.A(n_1143),
.B(n_1110),
.Y(n_1213)
);

AOI21x1_ASAP7_75t_SL g1214 ( 
.A1(n_1156),
.A2(n_1125),
.B(n_1089),
.Y(n_1214)
);

OAI21xp5_ASAP7_75t_L g1215 ( 
.A1(n_1147),
.A2(n_1101),
.B(n_1132),
.Y(n_1215)
);

INVx4_ASAP7_75t_L g1216 ( 
.A(n_1168),
.Y(n_1216)
);

AOI21x1_ASAP7_75t_L g1217 ( 
.A1(n_1187),
.A2(n_1132),
.B(n_1088),
.Y(n_1217)
);

NAND2xp5_ASAP7_75t_L g1218 ( 
.A(n_1143),
.B(n_1128),
.Y(n_1218)
);

AOI21x1_ASAP7_75t_L g1219 ( 
.A1(n_1198),
.A2(n_1147),
.B(n_1158),
.Y(n_1219)
);

NOR2xp67_ASAP7_75t_SL g1220 ( 
.A(n_1170),
.B(n_977),
.Y(n_1220)
);

OAI21x1_ASAP7_75t_L g1221 ( 
.A1(n_1178),
.A2(n_1137),
.B(n_1124),
.Y(n_1221)
);

AOI21xp5_ASAP7_75t_L g1222 ( 
.A1(n_1142),
.A2(n_977),
.B(n_1124),
.Y(n_1222)
);

OAI21xp5_ASAP7_75t_L g1223 ( 
.A1(n_1200),
.A2(n_520),
.B(n_513),
.Y(n_1223)
);

AOI21xp5_ASAP7_75t_L g1224 ( 
.A1(n_1178),
.A2(n_835),
.B(n_834),
.Y(n_1224)
);

OAI21xp5_ASAP7_75t_L g1225 ( 
.A1(n_1200),
.A2(n_530),
.B(n_529),
.Y(n_1225)
);

INVx2_ASAP7_75t_SL g1226 ( 
.A(n_1167),
.Y(n_1226)
);

NOR2xp33_ASAP7_75t_L g1227 ( 
.A(n_1207),
.B(n_531),
.Y(n_1227)
);

OAI21xp5_ASAP7_75t_L g1228 ( 
.A1(n_1186),
.A2(n_534),
.B(n_532),
.Y(n_1228)
);

INVx2_ASAP7_75t_L g1229 ( 
.A(n_1151),
.Y(n_1229)
);

AOI21xp5_ASAP7_75t_L g1230 ( 
.A1(n_1185),
.A2(n_835),
.B(n_834),
.Y(n_1230)
);

INVx2_ASAP7_75t_SL g1231 ( 
.A(n_1152),
.Y(n_1231)
);

NAND2xp5_ASAP7_75t_L g1232 ( 
.A(n_1203),
.B(n_742),
.Y(n_1232)
);

OAI21x1_ASAP7_75t_L g1233 ( 
.A1(n_1185),
.A2(n_835),
.B(n_872),
.Y(n_1233)
);

AND2x2_ASAP7_75t_L g1234 ( 
.A(n_1203),
.B(n_536),
.Y(n_1234)
);

A2O1A1Ixp33_ASAP7_75t_L g1235 ( 
.A1(n_1202),
.A2(n_541),
.B(n_543),
.C(n_538),
.Y(n_1235)
);

OAI22xp5_ASAP7_75t_L g1236 ( 
.A1(n_1201),
.A2(n_553),
.B1(n_558),
.B2(n_544),
.Y(n_1236)
);

INVx2_ASAP7_75t_L g1237 ( 
.A(n_1154),
.Y(n_1237)
);

A2O1A1Ixp33_ASAP7_75t_L g1238 ( 
.A1(n_1150),
.A2(n_567),
.B(n_569),
.C(n_565),
.Y(n_1238)
);

A2O1A1Ixp33_ASAP7_75t_L g1239 ( 
.A1(n_1201),
.A2(n_573),
.B(n_576),
.C(n_571),
.Y(n_1239)
);

OAI21x1_ASAP7_75t_L g1240 ( 
.A1(n_1182),
.A2(n_872),
.B(n_835),
.Y(n_1240)
);

AND2x4_ASAP7_75t_L g1241 ( 
.A(n_1166),
.B(n_872),
.Y(n_1241)
);

NOR2xp33_ASAP7_75t_L g1242 ( 
.A(n_1191),
.B(n_577),
.Y(n_1242)
);

NAND2xp5_ASAP7_75t_L g1243 ( 
.A(n_1160),
.B(n_580),
.Y(n_1243)
);

AOI21xp5_ASAP7_75t_L g1244 ( 
.A1(n_1160),
.A2(n_872),
.B(n_582),
.Y(n_1244)
);

HB1xp67_ASAP7_75t_L g1245 ( 
.A(n_1189),
.Y(n_1245)
);

AOI21xp5_ASAP7_75t_L g1246 ( 
.A1(n_1165),
.A2(n_1188),
.B(n_1163),
.Y(n_1246)
);

INVx3_ASAP7_75t_L g1247 ( 
.A(n_1205),
.Y(n_1247)
);

O2A1O1Ixp5_ASAP7_75t_L g1248 ( 
.A1(n_1163),
.A2(n_584),
.B(n_585),
.C(n_581),
.Y(n_1248)
);

AOI21xp5_ASAP7_75t_L g1249 ( 
.A1(n_1159),
.A2(n_1164),
.B(n_1145),
.Y(n_1249)
);

BUFx6f_ASAP7_75t_L g1250 ( 
.A(n_1189),
.Y(n_1250)
);

OAI21xp5_ASAP7_75t_L g1251 ( 
.A1(n_1161),
.A2(n_590),
.B(n_588),
.Y(n_1251)
);

BUFx2_ASAP7_75t_L g1252 ( 
.A(n_1172),
.Y(n_1252)
);

OAI21x1_ASAP7_75t_SL g1253 ( 
.A1(n_1192),
.A2(n_77),
.B(n_75),
.Y(n_1253)
);

NAND2xp5_ASAP7_75t_L g1254 ( 
.A(n_1166),
.B(n_592),
.Y(n_1254)
);

AOI21x1_ASAP7_75t_L g1255 ( 
.A1(n_1204),
.A2(n_598),
.B(n_596),
.Y(n_1255)
);

OAI21x1_ASAP7_75t_L g1256 ( 
.A1(n_1173),
.A2(n_79),
.B(n_78),
.Y(n_1256)
);

NAND2xp5_ASAP7_75t_L g1257 ( 
.A(n_1193),
.B(n_600),
.Y(n_1257)
);

OAI21x1_ASAP7_75t_L g1258 ( 
.A1(n_1176),
.A2(n_84),
.B(n_81),
.Y(n_1258)
);

NAND2xp5_ASAP7_75t_L g1259 ( 
.A(n_1190),
.B(n_605),
.Y(n_1259)
);

AOI21xp5_ASAP7_75t_L g1260 ( 
.A1(n_1141),
.A2(n_608),
.B(n_87),
.Y(n_1260)
);

OAI21x1_ASAP7_75t_L g1261 ( 
.A1(n_1181),
.A2(n_88),
.B(n_86),
.Y(n_1261)
);

BUFx3_ASAP7_75t_L g1262 ( 
.A(n_1155),
.Y(n_1262)
);

OAI21x1_ASAP7_75t_L g1263 ( 
.A1(n_1183),
.A2(n_90),
.B(n_89),
.Y(n_1263)
);

INVx3_ASAP7_75t_L g1264 ( 
.A(n_1205),
.Y(n_1264)
);

NAND2x1p5_ASAP7_75t_L g1265 ( 
.A(n_1180),
.B(n_91),
.Y(n_1265)
);

OAI22xp5_ASAP7_75t_L g1266 ( 
.A1(n_1169),
.A2(n_3),
.B1(n_1),
.B2(n_2),
.Y(n_1266)
);

INVx2_ASAP7_75t_L g1267 ( 
.A(n_1197),
.Y(n_1267)
);

NOR2xp33_ASAP7_75t_SL g1268 ( 
.A(n_1184),
.B(n_92),
.Y(n_1268)
);

OAI21x1_ASAP7_75t_L g1269 ( 
.A1(n_1162),
.A2(n_95),
.B(n_93),
.Y(n_1269)
);

AND2x2_ASAP7_75t_L g1270 ( 
.A(n_1189),
.B(n_3),
.Y(n_1270)
);

INVx6_ASAP7_75t_SL g1271 ( 
.A(n_1177),
.Y(n_1271)
);

NAND2xp5_ASAP7_75t_L g1272 ( 
.A(n_1195),
.B(n_4),
.Y(n_1272)
);

NAND2x1p5_ASAP7_75t_L g1273 ( 
.A(n_1205),
.B(n_97),
.Y(n_1273)
);

NAND2xp5_ASAP7_75t_L g1274 ( 
.A(n_1199),
.B(n_5),
.Y(n_1274)
);

OAI21x1_ASAP7_75t_L g1275 ( 
.A1(n_1148),
.A2(n_99),
.B(n_98),
.Y(n_1275)
);

HB1xp67_ASAP7_75t_L g1276 ( 
.A(n_1148),
.Y(n_1276)
);

INVx1_ASAP7_75t_L g1277 ( 
.A(n_1157),
.Y(n_1277)
);

AOI21x1_ASAP7_75t_SL g1278 ( 
.A1(n_1196),
.A2(n_5),
.B(n_6),
.Y(n_1278)
);

AO31x2_ASAP7_75t_L g1279 ( 
.A1(n_1194),
.A2(n_1157),
.A3(n_1174),
.B(n_1149),
.Y(n_1279)
);

AND2x2_ASAP7_75t_L g1280 ( 
.A(n_1179),
.B(n_1174),
.Y(n_1280)
);

AOI221xp5_ASAP7_75t_SL g1281 ( 
.A1(n_1175),
.A2(n_8),
.B1(n_6),
.B2(n_7),
.C(n_9),
.Y(n_1281)
);

AO31x2_ASAP7_75t_L g1282 ( 
.A1(n_1147),
.A2(n_9),
.A3(n_7),
.B(n_8),
.Y(n_1282)
);

NAND2xp5_ASAP7_75t_L g1283 ( 
.A(n_1171),
.B(n_10),
.Y(n_1283)
);

BUFx6f_ASAP7_75t_L g1284 ( 
.A(n_1189),
.Y(n_1284)
);

BUFx6f_ASAP7_75t_L g1285 ( 
.A(n_1189),
.Y(n_1285)
);

INVxp67_ASAP7_75t_SL g1286 ( 
.A(n_1276),
.Y(n_1286)
);

AOI21xp5_ASAP7_75t_L g1287 ( 
.A1(n_1211),
.A2(n_101),
.B(n_100),
.Y(n_1287)
);

NAND2xp5_ASAP7_75t_L g1288 ( 
.A(n_1218),
.B(n_10),
.Y(n_1288)
);

INVx1_ASAP7_75t_L g1289 ( 
.A(n_1212),
.Y(n_1289)
);

INVx3_ASAP7_75t_SL g1290 ( 
.A(n_1216),
.Y(n_1290)
);

NAND2xp5_ASAP7_75t_L g1291 ( 
.A(n_1213),
.B(n_11),
.Y(n_1291)
);

INVx2_ASAP7_75t_L g1292 ( 
.A(n_1229),
.Y(n_1292)
);

AOI21xp5_ASAP7_75t_L g1293 ( 
.A1(n_1222),
.A2(n_103),
.B(n_102),
.Y(n_1293)
);

AOI21xp5_ASAP7_75t_L g1294 ( 
.A1(n_1246),
.A2(n_107),
.B(n_105),
.Y(n_1294)
);

CKINVDCx20_ASAP7_75t_R g1295 ( 
.A(n_1262),
.Y(n_1295)
);

AND2x4_ASAP7_75t_L g1296 ( 
.A(n_1280),
.B(n_1252),
.Y(n_1296)
);

AND2x2_ASAP7_75t_L g1297 ( 
.A(n_1209),
.B(n_108),
.Y(n_1297)
);

NAND2xp5_ASAP7_75t_SL g1298 ( 
.A(n_1243),
.B(n_109),
.Y(n_1298)
);

NAND2xp5_ASAP7_75t_L g1299 ( 
.A(n_1237),
.B(n_1267),
.Y(n_1299)
);

AOI21xp33_ASAP7_75t_L g1300 ( 
.A1(n_1215),
.A2(n_13),
.B(n_14),
.Y(n_1300)
);

OAI21x1_ASAP7_75t_L g1301 ( 
.A1(n_1233),
.A2(n_111),
.B(n_110),
.Y(n_1301)
);

NAND2xp5_ASAP7_75t_L g1302 ( 
.A(n_1234),
.B(n_13),
.Y(n_1302)
);

INVx1_ASAP7_75t_L g1303 ( 
.A(n_1282),
.Y(n_1303)
);

INVx2_ASAP7_75t_L g1304 ( 
.A(n_1277),
.Y(n_1304)
);

BUFx4f_ASAP7_75t_SL g1305 ( 
.A(n_1271),
.Y(n_1305)
);

AOI22xp5_ASAP7_75t_L g1306 ( 
.A1(n_1227),
.A2(n_1266),
.B1(n_1268),
.B2(n_1281),
.Y(n_1306)
);

NAND2xp5_ASAP7_75t_L g1307 ( 
.A(n_1249),
.B(n_14),
.Y(n_1307)
);

CKINVDCx8_ASAP7_75t_R g1308 ( 
.A(n_1250),
.Y(n_1308)
);

NOR2xp33_ASAP7_75t_L g1309 ( 
.A(n_1242),
.B(n_112),
.Y(n_1309)
);

HB1xp67_ASAP7_75t_L g1310 ( 
.A(n_1279),
.Y(n_1310)
);

INVx1_ASAP7_75t_L g1311 ( 
.A(n_1282),
.Y(n_1311)
);

INVx3_ASAP7_75t_SL g1312 ( 
.A(n_1231),
.Y(n_1312)
);

CKINVDCx20_ASAP7_75t_R g1313 ( 
.A(n_1245),
.Y(n_1313)
);

HB1xp67_ASAP7_75t_L g1314 ( 
.A(n_1279),
.Y(n_1314)
);

BUFx4_ASAP7_75t_SL g1315 ( 
.A(n_1271),
.Y(n_1315)
);

AOI22xp33_ASAP7_75t_L g1316 ( 
.A1(n_1228),
.A2(n_1225),
.B1(n_1223),
.B2(n_1283),
.Y(n_1316)
);

AOI22xp33_ASAP7_75t_L g1317 ( 
.A1(n_1270),
.A2(n_17),
.B1(n_15),
.B2(n_16),
.Y(n_1317)
);

AOI22xp33_ASAP7_75t_L g1318 ( 
.A1(n_1253),
.A2(n_18),
.B1(n_15),
.B2(n_17),
.Y(n_1318)
);

INVx2_ASAP7_75t_L g1319 ( 
.A(n_1250),
.Y(n_1319)
);

AOI21xp5_ASAP7_75t_L g1320 ( 
.A1(n_1224),
.A2(n_1230),
.B(n_1244),
.Y(n_1320)
);

AOI21x1_ASAP7_75t_L g1321 ( 
.A1(n_1217),
.A2(n_117),
.B(n_114),
.Y(n_1321)
);

AOI21xp5_ASAP7_75t_L g1322 ( 
.A1(n_1260),
.A2(n_120),
.B(n_119),
.Y(n_1322)
);

INVx2_ASAP7_75t_L g1323 ( 
.A(n_1285),
.Y(n_1323)
);

INVx2_ASAP7_75t_L g1324 ( 
.A(n_1285),
.Y(n_1324)
);

INVx1_ASAP7_75t_L g1325 ( 
.A(n_1282),
.Y(n_1325)
);

INVx1_ASAP7_75t_SL g1326 ( 
.A(n_1232),
.Y(n_1326)
);

NAND2xp5_ASAP7_75t_L g1327 ( 
.A(n_1210),
.B(n_18),
.Y(n_1327)
);

OAI22xp5_ASAP7_75t_L g1328 ( 
.A1(n_1272),
.A2(n_21),
.B1(n_19),
.B2(n_20),
.Y(n_1328)
);

INVx1_ASAP7_75t_L g1329 ( 
.A(n_1219),
.Y(n_1329)
);

A2O1A1Ixp33_ASAP7_75t_SL g1330 ( 
.A1(n_1220),
.A2(n_22),
.B(n_19),
.C(n_20),
.Y(n_1330)
);

NAND2xp5_ASAP7_75t_L g1331 ( 
.A(n_1226),
.B(n_22),
.Y(n_1331)
);

AND2x2_ASAP7_75t_L g1332 ( 
.A(n_1274),
.B(n_1279),
.Y(n_1332)
);

BUFx3_ASAP7_75t_L g1333 ( 
.A(n_1247),
.Y(n_1333)
);

INVx2_ASAP7_75t_L g1334 ( 
.A(n_1285),
.Y(n_1334)
);

AOI22xp33_ASAP7_75t_L g1335 ( 
.A1(n_1253),
.A2(n_25),
.B1(n_23),
.B2(n_24),
.Y(n_1335)
);

NAND2xp5_ASAP7_75t_L g1336 ( 
.A(n_1257),
.B(n_23),
.Y(n_1336)
);

AND2x4_ASAP7_75t_L g1337 ( 
.A(n_1250),
.B(n_121),
.Y(n_1337)
);

AND2x2_ASAP7_75t_L g1338 ( 
.A(n_1284),
.B(n_122),
.Y(n_1338)
);

INVx3_ASAP7_75t_L g1339 ( 
.A(n_1284),
.Y(n_1339)
);

HB1xp67_ASAP7_75t_L g1340 ( 
.A(n_1284),
.Y(n_1340)
);

AOI21xp5_ASAP7_75t_L g1341 ( 
.A1(n_1221),
.A2(n_124),
.B(n_123),
.Y(n_1341)
);

AOI22xp33_ASAP7_75t_L g1342 ( 
.A1(n_1251),
.A2(n_26),
.B1(n_24),
.B2(n_25),
.Y(n_1342)
);

AND2x2_ASAP7_75t_L g1343 ( 
.A(n_1264),
.B(n_125),
.Y(n_1343)
);

NAND2xp5_ASAP7_75t_L g1344 ( 
.A(n_1259),
.B(n_26),
.Y(n_1344)
);

NAND2xp5_ASAP7_75t_SL g1345 ( 
.A(n_1248),
.B(n_126),
.Y(n_1345)
);

INVx1_ASAP7_75t_SL g1346 ( 
.A(n_1254),
.Y(n_1346)
);

INVx1_ASAP7_75t_L g1347 ( 
.A(n_1208),
.Y(n_1347)
);

AOI21xp5_ASAP7_75t_L g1348 ( 
.A1(n_1240),
.A2(n_128),
.B(n_127),
.Y(n_1348)
);

AOI21xp5_ASAP7_75t_L g1349 ( 
.A1(n_1269),
.A2(n_130),
.B(n_129),
.Y(n_1349)
);

INVx2_ASAP7_75t_L g1350 ( 
.A(n_1241),
.Y(n_1350)
);

BUFx6f_ASAP7_75t_L g1351 ( 
.A(n_1241),
.Y(n_1351)
);

INVx3_ASAP7_75t_L g1352 ( 
.A(n_1265),
.Y(n_1352)
);

OR2x2_ASAP7_75t_L g1353 ( 
.A(n_1273),
.B(n_27),
.Y(n_1353)
);

BUFx3_ASAP7_75t_L g1354 ( 
.A(n_1275),
.Y(n_1354)
);

INVx1_ASAP7_75t_L g1355 ( 
.A(n_1256),
.Y(n_1355)
);

AND2x2_ASAP7_75t_SL g1356 ( 
.A(n_1278),
.B(n_27),
.Y(n_1356)
);

INVx1_ASAP7_75t_L g1357 ( 
.A(n_1258),
.Y(n_1357)
);

NAND2xp5_ASAP7_75t_L g1358 ( 
.A(n_1235),
.B(n_28),
.Y(n_1358)
);

HB1xp67_ASAP7_75t_L g1359 ( 
.A(n_1261),
.Y(n_1359)
);

AOI21xp5_ASAP7_75t_L g1360 ( 
.A1(n_1263),
.A2(n_136),
.B(n_131),
.Y(n_1360)
);

AND2x2_ASAP7_75t_L g1361 ( 
.A(n_1296),
.B(n_1255),
.Y(n_1361)
);

AND2x4_ASAP7_75t_L g1362 ( 
.A(n_1286),
.B(n_1238),
.Y(n_1362)
);

OR2x2_ASAP7_75t_L g1363 ( 
.A(n_1326),
.B(n_1236),
.Y(n_1363)
);

INVx2_ASAP7_75t_SL g1364 ( 
.A(n_1315),
.Y(n_1364)
);

NOR2xp67_ASAP7_75t_L g1365 ( 
.A(n_1344),
.B(n_28),
.Y(n_1365)
);

OA21x2_ASAP7_75t_L g1366 ( 
.A1(n_1341),
.A2(n_1239),
.B(n_1214),
.Y(n_1366)
);

AND2x2_ASAP7_75t_L g1367 ( 
.A(n_1296),
.B(n_29),
.Y(n_1367)
);

HB1xp67_ASAP7_75t_L g1368 ( 
.A(n_1326),
.Y(n_1368)
);

NAND2xp5_ASAP7_75t_L g1369 ( 
.A(n_1346),
.B(n_29),
.Y(n_1369)
);

A2O1A1Ixp33_ASAP7_75t_L g1370 ( 
.A1(n_1306),
.A2(n_34),
.B(n_30),
.C(n_31),
.Y(n_1370)
);

AND2x2_ASAP7_75t_L g1371 ( 
.A(n_1332),
.B(n_30),
.Y(n_1371)
);

AND2x2_ASAP7_75t_L g1372 ( 
.A(n_1346),
.B(n_34),
.Y(n_1372)
);

A2O1A1Ixp33_ASAP7_75t_L g1373 ( 
.A1(n_1306),
.A2(n_37),
.B(n_35),
.C(n_36),
.Y(n_1373)
);

A2O1A1Ixp33_ASAP7_75t_L g1374 ( 
.A1(n_1316),
.A2(n_37),
.B(n_35),
.C(n_36),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_1303),
.Y(n_1375)
);

OA21x2_ASAP7_75t_L g1376 ( 
.A1(n_1311),
.A2(n_38),
.B(n_39),
.Y(n_1376)
);

NAND2xp5_ASAP7_75t_L g1377 ( 
.A(n_1289),
.B(n_1292),
.Y(n_1377)
);

NAND2x1p5_ASAP7_75t_L g1378 ( 
.A(n_1352),
.B(n_137),
.Y(n_1378)
);

AOI21xp5_ASAP7_75t_SL g1379 ( 
.A1(n_1298),
.A2(n_143),
.B(n_141),
.Y(n_1379)
);

BUFx4_ASAP7_75t_R g1380 ( 
.A(n_1333),
.Y(n_1380)
);

BUFx6f_ASAP7_75t_L g1381 ( 
.A(n_1312),
.Y(n_1381)
);

OA22x2_ASAP7_75t_L g1382 ( 
.A1(n_1328),
.A2(n_40),
.B1(n_38),
.B2(n_39),
.Y(n_1382)
);

AND2x2_ASAP7_75t_L g1383 ( 
.A(n_1340),
.B(n_40),
.Y(n_1383)
);

AOI21xp5_ASAP7_75t_SL g1384 ( 
.A1(n_1294),
.A2(n_146),
.B(n_145),
.Y(n_1384)
);

O2A1O1Ixp33_ASAP7_75t_L g1385 ( 
.A1(n_1300),
.A2(n_43),
.B(n_41),
.C(n_42),
.Y(n_1385)
);

INVx2_ASAP7_75t_L g1386 ( 
.A(n_1304),
.Y(n_1386)
);

AOI21xp5_ASAP7_75t_SL g1387 ( 
.A1(n_1345),
.A2(n_148),
.B(n_147),
.Y(n_1387)
);

OR2x2_ASAP7_75t_L g1388 ( 
.A(n_1325),
.B(n_43),
.Y(n_1388)
);

AOI21xp5_ASAP7_75t_L g1389 ( 
.A1(n_1320),
.A2(n_157),
.B(n_151),
.Y(n_1389)
);

A2O1A1Ixp33_ASAP7_75t_L g1390 ( 
.A1(n_1309),
.A2(n_46),
.B(n_44),
.C(n_45),
.Y(n_1390)
);

OR2x2_ASAP7_75t_L g1391 ( 
.A(n_1310),
.B(n_44),
.Y(n_1391)
);

INVx1_ASAP7_75t_L g1392 ( 
.A(n_1314),
.Y(n_1392)
);

AND2x2_ASAP7_75t_L g1393 ( 
.A(n_1319),
.B(n_45),
.Y(n_1393)
);

INVx3_ASAP7_75t_L g1394 ( 
.A(n_1308),
.Y(n_1394)
);

INVx1_ASAP7_75t_SL g1395 ( 
.A(n_1313),
.Y(n_1395)
);

NOR2xp33_ASAP7_75t_L g1396 ( 
.A(n_1295),
.B(n_46),
.Y(n_1396)
);

AOI21xp5_ASAP7_75t_L g1397 ( 
.A1(n_1287),
.A2(n_160),
.B(n_158),
.Y(n_1397)
);

AOI21xp5_ASAP7_75t_L g1398 ( 
.A1(n_1322),
.A2(n_163),
.B(n_162),
.Y(n_1398)
);

A2O1A1Ixp33_ASAP7_75t_SL g1399 ( 
.A1(n_1300),
.A2(n_49),
.B(n_47),
.C(n_48),
.Y(n_1399)
);

A2O1A1Ixp33_ASAP7_75t_L g1400 ( 
.A1(n_1342),
.A2(n_50),
.B(n_48),
.C(n_49),
.Y(n_1400)
);

AND2x2_ASAP7_75t_L g1401 ( 
.A(n_1323),
.B(n_52),
.Y(n_1401)
);

INVx3_ASAP7_75t_L g1402 ( 
.A(n_1339),
.Y(n_1402)
);

INVx2_ASAP7_75t_SL g1403 ( 
.A(n_1290),
.Y(n_1403)
);

O2A1O1Ixp5_ASAP7_75t_L g1404 ( 
.A1(n_1328),
.A2(n_54),
.B(n_52),
.C(n_53),
.Y(n_1404)
);

AOI21xp5_ASAP7_75t_SL g1405 ( 
.A1(n_1307),
.A2(n_165),
.B(n_164),
.Y(n_1405)
);

INVx2_ASAP7_75t_L g1406 ( 
.A(n_1299),
.Y(n_1406)
);

INVx2_ASAP7_75t_L g1407 ( 
.A(n_1324),
.Y(n_1407)
);

INVxp33_ASAP7_75t_L g1408 ( 
.A(n_1302),
.Y(n_1408)
);

AND2x2_ASAP7_75t_L g1409 ( 
.A(n_1334),
.B(n_53),
.Y(n_1409)
);

NAND2xp5_ASAP7_75t_L g1410 ( 
.A(n_1288),
.B(n_54),
.Y(n_1410)
);

OAI22xp5_ASAP7_75t_L g1411 ( 
.A1(n_1318),
.A2(n_57),
.B1(n_55),
.B2(n_56),
.Y(n_1411)
);

OR2x2_ASAP7_75t_L g1412 ( 
.A(n_1327),
.B(n_55),
.Y(n_1412)
);

A2O1A1Ixp33_ASAP7_75t_SL g1413 ( 
.A1(n_1329),
.A2(n_59),
.B(n_56),
.C(n_58),
.Y(n_1413)
);

AND2x4_ASAP7_75t_L g1414 ( 
.A(n_1339),
.B(n_437),
.Y(n_1414)
);

INVx2_ASAP7_75t_L g1415 ( 
.A(n_1347),
.Y(n_1415)
);

AND2x2_ASAP7_75t_L g1416 ( 
.A(n_1297),
.B(n_58),
.Y(n_1416)
);

NOR2xp33_ASAP7_75t_L g1417 ( 
.A(n_1336),
.B(n_59),
.Y(n_1417)
);

BUFx2_ASAP7_75t_L g1418 ( 
.A(n_1351),
.Y(n_1418)
);

INVx1_ASAP7_75t_L g1419 ( 
.A(n_1359),
.Y(n_1419)
);

BUFx4f_ASAP7_75t_L g1420 ( 
.A(n_1351),
.Y(n_1420)
);

A2O1A1Ixp33_ASAP7_75t_L g1421 ( 
.A1(n_1358),
.A2(n_60),
.B(n_61),
.C(n_62),
.Y(n_1421)
);

NAND2xp5_ASAP7_75t_L g1422 ( 
.A(n_1291),
.B(n_60),
.Y(n_1422)
);

AND2x2_ASAP7_75t_L g1423 ( 
.A(n_1350),
.B(n_61),
.Y(n_1423)
);

AOI21x1_ASAP7_75t_SL g1424 ( 
.A1(n_1358),
.A2(n_63),
.B(n_64),
.Y(n_1424)
);

HB1xp67_ASAP7_75t_L g1425 ( 
.A(n_1355),
.Y(n_1425)
);

A2O1A1Ixp33_ASAP7_75t_SL g1426 ( 
.A1(n_1352),
.A2(n_63),
.B(n_64),
.C(n_65),
.Y(n_1426)
);

HB1xp67_ASAP7_75t_L g1427 ( 
.A(n_1357),
.Y(n_1427)
);

AND2x2_ASAP7_75t_L g1428 ( 
.A(n_1338),
.B(n_65),
.Y(n_1428)
);

AOI21xp5_ASAP7_75t_L g1429 ( 
.A1(n_1293),
.A2(n_167),
.B(n_166),
.Y(n_1429)
);

CKINVDCx16_ASAP7_75t_R g1430 ( 
.A(n_1353),
.Y(n_1430)
);

INVx1_ASAP7_75t_L g1431 ( 
.A(n_1291),
.Y(n_1431)
);

NOR2xp33_ASAP7_75t_R g1432 ( 
.A(n_1305),
.B(n_168),
.Y(n_1432)
);

INVx1_ASAP7_75t_L g1433 ( 
.A(n_1375),
.Y(n_1433)
);

AND2x2_ASAP7_75t_L g1434 ( 
.A(n_1425),
.B(n_1356),
.Y(n_1434)
);

INVx1_ASAP7_75t_L g1435 ( 
.A(n_1368),
.Y(n_1435)
);

INVx3_ASAP7_75t_L g1436 ( 
.A(n_1407),
.Y(n_1436)
);

INVx2_ASAP7_75t_L g1437 ( 
.A(n_1415),
.Y(n_1437)
);

OR2x2_ASAP7_75t_L g1438 ( 
.A(n_1392),
.B(n_1331),
.Y(n_1438)
);

INVx1_ASAP7_75t_L g1439 ( 
.A(n_1375),
.Y(n_1439)
);

AND2x2_ASAP7_75t_L g1440 ( 
.A(n_1427),
.B(n_1354),
.Y(n_1440)
);

OAI21x1_ASAP7_75t_L g1441 ( 
.A1(n_1419),
.A2(n_1321),
.B(n_1301),
.Y(n_1441)
);

OR2x2_ASAP7_75t_L g1442 ( 
.A(n_1431),
.B(n_1330),
.Y(n_1442)
);

BUFx2_ASAP7_75t_L g1443 ( 
.A(n_1361),
.Y(n_1443)
);

INVx2_ASAP7_75t_L g1444 ( 
.A(n_1386),
.Y(n_1444)
);

INVx1_ASAP7_75t_L g1445 ( 
.A(n_1377),
.Y(n_1445)
);

AND2x2_ASAP7_75t_L g1446 ( 
.A(n_1371),
.B(n_1351),
.Y(n_1446)
);

AOI21xp5_ASAP7_75t_L g1447 ( 
.A1(n_1389),
.A2(n_1360),
.B(n_1349),
.Y(n_1447)
);

INVx2_ASAP7_75t_L g1448 ( 
.A(n_1406),
.Y(n_1448)
);

HB1xp67_ASAP7_75t_L g1449 ( 
.A(n_1391),
.Y(n_1449)
);

INVx1_ASAP7_75t_L g1450 ( 
.A(n_1376),
.Y(n_1450)
);

INVx1_ASAP7_75t_L g1451 ( 
.A(n_1376),
.Y(n_1451)
);

AO21x2_ASAP7_75t_L g1452 ( 
.A1(n_1413),
.A2(n_1348),
.B(n_1343),
.Y(n_1452)
);

INVx2_ASAP7_75t_L g1453 ( 
.A(n_1402),
.Y(n_1453)
);

INVx2_ASAP7_75t_L g1454 ( 
.A(n_1402),
.Y(n_1454)
);

BUFx2_ASAP7_75t_L g1455 ( 
.A(n_1418),
.Y(n_1455)
);

INVx1_ASAP7_75t_L g1456 ( 
.A(n_1388),
.Y(n_1456)
);

INVx1_ASAP7_75t_L g1457 ( 
.A(n_1412),
.Y(n_1457)
);

AND2x2_ASAP7_75t_L g1458 ( 
.A(n_1430),
.B(n_1335),
.Y(n_1458)
);

INVx1_ASAP7_75t_L g1459 ( 
.A(n_1369),
.Y(n_1459)
);

INVx2_ASAP7_75t_L g1460 ( 
.A(n_1366),
.Y(n_1460)
);

INVx1_ASAP7_75t_L g1461 ( 
.A(n_1372),
.Y(n_1461)
);

INVx2_ASAP7_75t_L g1462 ( 
.A(n_1366),
.Y(n_1462)
);

INVx2_ASAP7_75t_L g1463 ( 
.A(n_1393),
.Y(n_1463)
);

INVx2_ASAP7_75t_SL g1464 ( 
.A(n_1381),
.Y(n_1464)
);

INVx2_ASAP7_75t_L g1465 ( 
.A(n_1401),
.Y(n_1465)
);

INVx1_ASAP7_75t_L g1466 ( 
.A(n_1363),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_1409),
.Y(n_1467)
);

INVx1_ASAP7_75t_L g1468 ( 
.A(n_1422),
.Y(n_1468)
);

INVx2_ASAP7_75t_L g1469 ( 
.A(n_1423),
.Y(n_1469)
);

INVx3_ASAP7_75t_L g1470 ( 
.A(n_1362),
.Y(n_1470)
);

INVx1_ASAP7_75t_L g1471 ( 
.A(n_1383),
.Y(n_1471)
);

INVx1_ASAP7_75t_L g1472 ( 
.A(n_1367),
.Y(n_1472)
);

INVx3_ASAP7_75t_L g1473 ( 
.A(n_1362),
.Y(n_1473)
);

INVx1_ASAP7_75t_L g1474 ( 
.A(n_1410),
.Y(n_1474)
);

INVx2_ASAP7_75t_L g1475 ( 
.A(n_1414),
.Y(n_1475)
);

BUFx6f_ASAP7_75t_L g1476 ( 
.A(n_1420),
.Y(n_1476)
);

INVx1_ASAP7_75t_L g1477 ( 
.A(n_1404),
.Y(n_1477)
);

OAI21xp5_ASAP7_75t_L g1478 ( 
.A1(n_1374),
.A2(n_1317),
.B(n_1337),
.Y(n_1478)
);

AND2x2_ASAP7_75t_L g1479 ( 
.A(n_1408),
.B(n_1428),
.Y(n_1479)
);

INVx1_ASAP7_75t_L g1480 ( 
.A(n_1385),
.Y(n_1480)
);

AND2x4_ASAP7_75t_L g1481 ( 
.A(n_1403),
.B(n_1394),
.Y(n_1481)
);

INVx3_ASAP7_75t_L g1482 ( 
.A(n_1381),
.Y(n_1482)
);

HB1xp67_ASAP7_75t_L g1483 ( 
.A(n_1380),
.Y(n_1483)
);

INVx2_ASAP7_75t_L g1484 ( 
.A(n_1414),
.Y(n_1484)
);

HB1xp67_ASAP7_75t_L g1485 ( 
.A(n_1433),
.Y(n_1485)
);

INVx1_ASAP7_75t_L g1486 ( 
.A(n_1433),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_1439),
.Y(n_1487)
);

INVx3_ASAP7_75t_L g1488 ( 
.A(n_1436),
.Y(n_1488)
);

OR2x2_ASAP7_75t_L g1489 ( 
.A(n_1443),
.B(n_1395),
.Y(n_1489)
);

AOI22xp33_ASAP7_75t_L g1490 ( 
.A1(n_1480),
.A2(n_1382),
.B1(n_1411),
.B2(n_1417),
.Y(n_1490)
);

AND2x4_ASAP7_75t_L g1491 ( 
.A(n_1470),
.B(n_1381),
.Y(n_1491)
);

OAI22xp5_ASAP7_75t_L g1492 ( 
.A1(n_1480),
.A2(n_1370),
.B1(n_1373),
.B2(n_1390),
.Y(n_1492)
);

INVx1_ASAP7_75t_L g1493 ( 
.A(n_1444),
.Y(n_1493)
);

OAI22xp33_ASAP7_75t_L g1494 ( 
.A1(n_1478),
.A2(n_1365),
.B1(n_1394),
.B2(n_1396),
.Y(n_1494)
);

INVx2_ASAP7_75t_L g1495 ( 
.A(n_1436),
.Y(n_1495)
);

OR2x2_ASAP7_75t_L g1496 ( 
.A(n_1443),
.B(n_1416),
.Y(n_1496)
);

AOI22xp33_ASAP7_75t_SL g1497 ( 
.A1(n_1458),
.A2(n_1432),
.B1(n_1424),
.B2(n_1421),
.Y(n_1497)
);

AOI22xp33_ASAP7_75t_L g1498 ( 
.A1(n_1477),
.A2(n_1397),
.B1(n_1398),
.B2(n_1429),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_1444),
.Y(n_1499)
);

BUFx4f_ASAP7_75t_SL g1500 ( 
.A(n_1481),
.Y(n_1500)
);

HB1xp67_ASAP7_75t_L g1501 ( 
.A(n_1450),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_1437),
.Y(n_1502)
);

OAI21xp33_ASAP7_75t_L g1503 ( 
.A1(n_1442),
.A2(n_1400),
.B(n_1405),
.Y(n_1503)
);

OR2x6_ASAP7_75t_L g1504 ( 
.A(n_1470),
.B(n_1384),
.Y(n_1504)
);

INVx3_ASAP7_75t_L g1505 ( 
.A(n_1436),
.Y(n_1505)
);

AND2x2_ASAP7_75t_L g1506 ( 
.A(n_1466),
.B(n_1364),
.Y(n_1506)
);

NAND2xp5_ASAP7_75t_L g1507 ( 
.A(n_1445),
.B(n_1448),
.Y(n_1507)
);

AND2x2_ASAP7_75t_L g1508 ( 
.A(n_1455),
.B(n_1420),
.Y(n_1508)
);

AND2x2_ASAP7_75t_L g1509 ( 
.A(n_1455),
.B(n_1378),
.Y(n_1509)
);

INVx2_ASAP7_75t_L g1510 ( 
.A(n_1453),
.Y(n_1510)
);

BUFx4f_ASAP7_75t_L g1511 ( 
.A(n_1476),
.Y(n_1511)
);

AND2x2_ASAP7_75t_L g1512 ( 
.A(n_1449),
.B(n_1337),
.Y(n_1512)
);

AND2x2_ASAP7_75t_L g1513 ( 
.A(n_1435),
.B(n_1387),
.Y(n_1513)
);

OR2x2_ASAP7_75t_L g1514 ( 
.A(n_1456),
.B(n_1399),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_1437),
.Y(n_1515)
);

NAND2xp5_ASAP7_75t_L g1516 ( 
.A(n_1448),
.B(n_1426),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_1438),
.Y(n_1517)
);

AND2x4_ASAP7_75t_L g1518 ( 
.A(n_1470),
.B(n_67),
.Y(n_1518)
);

AND2x2_ASAP7_75t_L g1519 ( 
.A(n_1473),
.B(n_1379),
.Y(n_1519)
);

AND2x2_ASAP7_75t_L g1520 ( 
.A(n_1473),
.B(n_68),
.Y(n_1520)
);

AOI22xp33_ASAP7_75t_L g1521 ( 
.A1(n_1473),
.A2(n_69),
.B1(n_70),
.B2(n_71),
.Y(n_1521)
);

INVxp67_ASAP7_75t_SL g1522 ( 
.A(n_1450),
.Y(n_1522)
);

AND2x2_ASAP7_75t_L g1523 ( 
.A(n_1479),
.B(n_69),
.Y(n_1523)
);

INVx1_ASAP7_75t_L g1524 ( 
.A(n_1438),
.Y(n_1524)
);

AND2x2_ASAP7_75t_L g1525 ( 
.A(n_1491),
.B(n_1457),
.Y(n_1525)
);

INVx2_ASAP7_75t_L g1526 ( 
.A(n_1488),
.Y(n_1526)
);

AND2x2_ASAP7_75t_L g1527 ( 
.A(n_1491),
.B(n_1479),
.Y(n_1527)
);

AND2x2_ASAP7_75t_L g1528 ( 
.A(n_1508),
.B(n_1481),
.Y(n_1528)
);

INVx1_ASAP7_75t_L g1529 ( 
.A(n_1485),
.Y(n_1529)
);

INVx2_ASAP7_75t_L g1530 ( 
.A(n_1488),
.Y(n_1530)
);

AOI22xp33_ASAP7_75t_L g1531 ( 
.A1(n_1492),
.A2(n_1458),
.B1(n_1452),
.B2(n_1468),
.Y(n_1531)
);

INVx1_ASAP7_75t_L g1532 ( 
.A(n_1485),
.Y(n_1532)
);

BUFx2_ASAP7_75t_SL g1533 ( 
.A(n_1518),
.Y(n_1533)
);

HB1xp67_ASAP7_75t_L g1534 ( 
.A(n_1501),
.Y(n_1534)
);

AO31x2_ASAP7_75t_L g1535 ( 
.A1(n_1516),
.A2(n_1451),
.A3(n_1462),
.B(n_1460),
.Y(n_1535)
);

AOI22xp5_ASAP7_75t_L g1536 ( 
.A1(n_1492),
.A2(n_1452),
.B1(n_1434),
.B2(n_1483),
.Y(n_1536)
);

AND2x2_ASAP7_75t_L g1537 ( 
.A(n_1496),
.B(n_1481),
.Y(n_1537)
);

AOI22xp5_ASAP7_75t_L g1538 ( 
.A1(n_1503),
.A2(n_1452),
.B1(n_1434),
.B2(n_1474),
.Y(n_1538)
);

AOI21xp5_ASAP7_75t_SL g1539 ( 
.A1(n_1504),
.A2(n_1494),
.B(n_1518),
.Y(n_1539)
);

INVxp67_ASAP7_75t_SL g1540 ( 
.A(n_1501),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_1486),
.Y(n_1541)
);

AND2x4_ASAP7_75t_L g1542 ( 
.A(n_1517),
.B(n_1440),
.Y(n_1542)
);

INVx1_ASAP7_75t_L g1543 ( 
.A(n_1487),
.Y(n_1543)
);

OR2x2_ASAP7_75t_L g1544 ( 
.A(n_1524),
.B(n_1469),
.Y(n_1544)
);

AND2x4_ASAP7_75t_L g1545 ( 
.A(n_1509),
.B(n_1440),
.Y(n_1545)
);

OR2x2_ASAP7_75t_L g1546 ( 
.A(n_1489),
.B(n_1469),
.Y(n_1546)
);

INVx2_ASAP7_75t_L g1547 ( 
.A(n_1505),
.Y(n_1547)
);

OR2x2_ASAP7_75t_L g1548 ( 
.A(n_1507),
.B(n_1463),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_1507),
.Y(n_1549)
);

BUFx2_ASAP7_75t_L g1550 ( 
.A(n_1527),
.Y(n_1550)
);

AND2x2_ASAP7_75t_L g1551 ( 
.A(n_1542),
.B(n_1506),
.Y(n_1551)
);

INVx1_ASAP7_75t_L g1552 ( 
.A(n_1543),
.Y(n_1552)
);

AND2x2_ASAP7_75t_L g1553 ( 
.A(n_1542),
.B(n_1519),
.Y(n_1553)
);

AND2x2_ASAP7_75t_L g1554 ( 
.A(n_1545),
.B(n_1512),
.Y(n_1554)
);

NAND2xp5_ASAP7_75t_L g1555 ( 
.A(n_1549),
.B(n_1514),
.Y(n_1555)
);

OR2x2_ASAP7_75t_L g1556 ( 
.A(n_1546),
.B(n_1516),
.Y(n_1556)
);

AND2x2_ASAP7_75t_L g1557 ( 
.A(n_1545),
.B(n_1482),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_1541),
.Y(n_1558)
);

INVx2_ASAP7_75t_SL g1559 ( 
.A(n_1534),
.Y(n_1559)
);

HB1xp67_ASAP7_75t_L g1560 ( 
.A(n_1534),
.Y(n_1560)
);

AND2x4_ASAP7_75t_L g1561 ( 
.A(n_1529),
.B(n_1522),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1532),
.Y(n_1562)
);

NAND2xp5_ASAP7_75t_L g1563 ( 
.A(n_1540),
.B(n_1522),
.Y(n_1563)
);

BUFx2_ASAP7_75t_L g1564 ( 
.A(n_1537),
.Y(n_1564)
);

OR2x2_ASAP7_75t_L g1565 ( 
.A(n_1548),
.B(n_1463),
.Y(n_1565)
);

AND2x2_ASAP7_75t_L g1566 ( 
.A(n_1525),
.B(n_1482),
.Y(n_1566)
);

INVx1_ASAP7_75t_SL g1567 ( 
.A(n_1533),
.Y(n_1567)
);

NAND2xp5_ASAP7_75t_L g1568 ( 
.A(n_1540),
.B(n_1538),
.Y(n_1568)
);

AND2x2_ASAP7_75t_L g1569 ( 
.A(n_1526),
.B(n_1505),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_1544),
.Y(n_1570)
);

AND2x2_ASAP7_75t_L g1571 ( 
.A(n_1528),
.B(n_1539),
.Y(n_1571)
);

OR2x2_ASAP7_75t_L g1572 ( 
.A(n_1536),
.B(n_1538),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_1535),
.Y(n_1573)
);

NAND3xp33_ASAP7_75t_SL g1574 ( 
.A(n_1572),
.B(n_1536),
.C(n_1531),
.Y(n_1574)
);

INVx5_ASAP7_75t_L g1575 ( 
.A(n_1559),
.Y(n_1575)
);

AO21x2_ASAP7_75t_L g1576 ( 
.A1(n_1568),
.A2(n_1494),
.B(n_1520),
.Y(n_1576)
);

OR2x2_ASAP7_75t_L g1577 ( 
.A(n_1556),
.B(n_1531),
.Y(n_1577)
);

BUFx3_ASAP7_75t_L g1578 ( 
.A(n_1567),
.Y(n_1578)
);

INVx1_ASAP7_75t_L g1579 ( 
.A(n_1560),
.Y(n_1579)
);

AND2x2_ASAP7_75t_L g1580 ( 
.A(n_1571),
.B(n_1482),
.Y(n_1580)
);

OAI22xp5_ASAP7_75t_L g1581 ( 
.A1(n_1568),
.A2(n_1497),
.B1(n_1490),
.B2(n_1498),
.Y(n_1581)
);

OAI321xp33_ASAP7_75t_L g1582 ( 
.A1(n_1555),
.A2(n_1563),
.A3(n_1559),
.B1(n_1562),
.B2(n_1550),
.C(n_1573),
.Y(n_1582)
);

OAI21x1_ASAP7_75t_L g1583 ( 
.A1(n_1563),
.A2(n_1547),
.B(n_1530),
.Y(n_1583)
);

INVx1_ASAP7_75t_L g1584 ( 
.A(n_1560),
.Y(n_1584)
);

INVx1_ASAP7_75t_L g1585 ( 
.A(n_1558),
.Y(n_1585)
);

AND2x2_ASAP7_75t_L g1586 ( 
.A(n_1557),
.B(n_1464),
.Y(n_1586)
);

INVx1_ASAP7_75t_L g1587 ( 
.A(n_1552),
.Y(n_1587)
);

INVx1_ASAP7_75t_L g1588 ( 
.A(n_1565),
.Y(n_1588)
);

INVx1_ASAP7_75t_L g1589 ( 
.A(n_1570),
.Y(n_1589)
);

AND2x2_ASAP7_75t_L g1590 ( 
.A(n_1578),
.B(n_1553),
.Y(n_1590)
);

AND2x2_ASAP7_75t_L g1591 ( 
.A(n_1580),
.B(n_1564),
.Y(n_1591)
);

OR2x2_ASAP7_75t_L g1592 ( 
.A(n_1577),
.B(n_1555),
.Y(n_1592)
);

INVx1_ASAP7_75t_L g1593 ( 
.A(n_1579),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_1584),
.Y(n_1594)
);

OR2x6_ASAP7_75t_SL g1595 ( 
.A(n_1581),
.B(n_1459),
.Y(n_1595)
);

NAND2xp5_ASAP7_75t_L g1596 ( 
.A(n_1589),
.B(n_1561),
.Y(n_1596)
);

HB1xp67_ASAP7_75t_L g1597 ( 
.A(n_1575),
.Y(n_1597)
);

AND2x2_ASAP7_75t_L g1598 ( 
.A(n_1586),
.B(n_1554),
.Y(n_1598)
);

INVx2_ASAP7_75t_L g1599 ( 
.A(n_1575),
.Y(n_1599)
);

INVx1_ASAP7_75t_L g1600 ( 
.A(n_1585),
.Y(n_1600)
);

OR2x2_ASAP7_75t_L g1601 ( 
.A(n_1576),
.B(n_1588),
.Y(n_1601)
);

NAND2x1_ASAP7_75t_L g1602 ( 
.A(n_1599),
.B(n_1582),
.Y(n_1602)
);

AND2x2_ASAP7_75t_L g1603 ( 
.A(n_1590),
.B(n_1551),
.Y(n_1603)
);

INVx1_ASAP7_75t_L g1604 ( 
.A(n_1597),
.Y(n_1604)
);

NAND3xp33_ASAP7_75t_L g1605 ( 
.A(n_1601),
.B(n_1575),
.C(n_1589),
.Y(n_1605)
);

AND2x4_ASAP7_75t_L g1606 ( 
.A(n_1597),
.B(n_1587),
.Y(n_1606)
);

NAND2xp5_ASAP7_75t_L g1607 ( 
.A(n_1593),
.B(n_1588),
.Y(n_1607)
);

OR2x2_ASAP7_75t_L g1608 ( 
.A(n_1592),
.B(n_1574),
.Y(n_1608)
);

AND2x2_ASAP7_75t_L g1609 ( 
.A(n_1591),
.B(n_1566),
.Y(n_1609)
);

INVx1_ASAP7_75t_L g1610 ( 
.A(n_1594),
.Y(n_1610)
);

AND2x2_ASAP7_75t_L g1611 ( 
.A(n_1598),
.B(n_1569),
.Y(n_1611)
);

INVx2_ASAP7_75t_SL g1612 ( 
.A(n_1596),
.Y(n_1612)
);

AND2x2_ASAP7_75t_L g1613 ( 
.A(n_1596),
.B(n_1569),
.Y(n_1613)
);

OR2x2_ASAP7_75t_L g1614 ( 
.A(n_1608),
.B(n_1612),
.Y(n_1614)
);

OAI221xp5_ASAP7_75t_L g1615 ( 
.A1(n_1602),
.A2(n_1600),
.B1(n_1497),
.B2(n_1595),
.C(n_1521),
.Y(n_1615)
);

O2A1O1Ixp33_ASAP7_75t_SL g1616 ( 
.A1(n_1605),
.A2(n_1464),
.B(n_1442),
.C(n_1461),
.Y(n_1616)
);

INVx1_ASAP7_75t_L g1617 ( 
.A(n_1604),
.Y(n_1617)
);

NAND2xp5_ASAP7_75t_L g1618 ( 
.A(n_1603),
.B(n_1561),
.Y(n_1618)
);

AND2x2_ASAP7_75t_L g1619 ( 
.A(n_1609),
.B(n_1583),
.Y(n_1619)
);

OR2x2_ASAP7_75t_L g1620 ( 
.A(n_1607),
.B(n_1561),
.Y(n_1620)
);

AND2x2_ASAP7_75t_L g1621 ( 
.A(n_1613),
.B(n_1611),
.Y(n_1621)
);

INVx1_ASAP7_75t_SL g1622 ( 
.A(n_1606),
.Y(n_1622)
);

INVx1_ASAP7_75t_L g1623 ( 
.A(n_1606),
.Y(n_1623)
);

INVx1_ASAP7_75t_L g1624 ( 
.A(n_1610),
.Y(n_1624)
);

OR2x2_ASAP7_75t_L g1625 ( 
.A(n_1614),
.B(n_1610),
.Y(n_1625)
);

AND2x2_ASAP7_75t_L g1626 ( 
.A(n_1621),
.B(n_1523),
.Y(n_1626)
);

INVxp67_ASAP7_75t_SL g1627 ( 
.A(n_1623),
.Y(n_1627)
);

AND2x2_ASAP7_75t_L g1628 ( 
.A(n_1622),
.B(n_1472),
.Y(n_1628)
);

INVxp33_ASAP7_75t_L g1629 ( 
.A(n_1618),
.Y(n_1629)
);

NAND2xp5_ASAP7_75t_L g1630 ( 
.A(n_1622),
.B(n_1535),
.Y(n_1630)
);

NOR2xp67_ASAP7_75t_L g1631 ( 
.A(n_1620),
.B(n_1617),
.Y(n_1631)
);

NAND2xp5_ASAP7_75t_L g1632 ( 
.A(n_1624),
.B(n_1619),
.Y(n_1632)
);

NOR2xp33_ASAP7_75t_SL g1633 ( 
.A(n_1615),
.B(n_1511),
.Y(n_1633)
);

AND2x2_ASAP7_75t_L g1634 ( 
.A(n_1616),
.B(n_1471),
.Y(n_1634)
);

INVx1_ASAP7_75t_L g1635 ( 
.A(n_1622),
.Y(n_1635)
);

OAI22xp5_ASAP7_75t_L g1636 ( 
.A1(n_1629),
.A2(n_1500),
.B1(n_1511),
.B2(n_1504),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_1627),
.Y(n_1637)
);

INVx1_ASAP7_75t_L g1638 ( 
.A(n_1635),
.Y(n_1638)
);

OAI22xp5_ASAP7_75t_L g1639 ( 
.A1(n_1625),
.A2(n_1504),
.B1(n_1467),
.B2(n_1465),
.Y(n_1639)
);

O2A1O1Ixp33_ASAP7_75t_L g1640 ( 
.A1(n_1632),
.A2(n_1447),
.B(n_1451),
.C(n_1460),
.Y(n_1640)
);

INVx1_ASAP7_75t_L g1641 ( 
.A(n_1628),
.Y(n_1641)
);

NAND2xp5_ASAP7_75t_L g1642 ( 
.A(n_1626),
.B(n_1535),
.Y(n_1642)
);

NAND2x1_ASAP7_75t_L g1643 ( 
.A(n_1631),
.B(n_1513),
.Y(n_1643)
);

AOI22xp5_ASAP7_75t_L g1644 ( 
.A1(n_1633),
.A2(n_1476),
.B1(n_1465),
.B2(n_1462),
.Y(n_1644)
);

OAI221xp5_ASAP7_75t_SL g1645 ( 
.A1(n_1630),
.A2(n_1475),
.B1(n_1484),
.B2(n_1446),
.C(n_1499),
.Y(n_1645)
);

OAI221xp5_ASAP7_75t_L g1646 ( 
.A1(n_1633),
.A2(n_1476),
.B1(n_1475),
.B2(n_1484),
.C(n_1493),
.Y(n_1646)
);

AND2x2_ASAP7_75t_L g1647 ( 
.A(n_1634),
.B(n_1446),
.Y(n_1647)
);

AOI222xp33_ASAP7_75t_L g1648 ( 
.A1(n_1631),
.A2(n_1515),
.B1(n_1502),
.B2(n_1476),
.C1(n_1510),
.C2(n_1495),
.Y(n_1648)
);

NAND2xp5_ASAP7_75t_L g1649 ( 
.A(n_1637),
.B(n_1453),
.Y(n_1649)
);

INVx1_ASAP7_75t_L g1650 ( 
.A(n_1638),
.Y(n_1650)
);

AND2x2_ASAP7_75t_L g1651 ( 
.A(n_1641),
.B(n_1454),
.Y(n_1651)
);

INVx1_ASAP7_75t_L g1652 ( 
.A(n_1647),
.Y(n_1652)
);

INVx1_ASAP7_75t_SL g1653 ( 
.A(n_1643),
.Y(n_1653)
);

INVx1_ASAP7_75t_L g1654 ( 
.A(n_1642),
.Y(n_1654)
);

NOR2xp33_ASAP7_75t_L g1655 ( 
.A(n_1646),
.B(n_71),
.Y(n_1655)
);

INVx1_ASAP7_75t_SL g1656 ( 
.A(n_1644),
.Y(n_1656)
);

NAND2xp5_ASAP7_75t_L g1657 ( 
.A(n_1648),
.B(n_1454),
.Y(n_1657)
);

NAND2xp5_ASAP7_75t_L g1658 ( 
.A(n_1639),
.B(n_72),
.Y(n_1658)
);

INVx3_ASAP7_75t_L g1659 ( 
.A(n_1645),
.Y(n_1659)
);

OAI21xp33_ASAP7_75t_L g1660 ( 
.A1(n_1636),
.A2(n_1476),
.B(n_1441),
.Y(n_1660)
);

AND2x2_ASAP7_75t_L g1661 ( 
.A(n_1640),
.B(n_72),
.Y(n_1661)
);

NOR2xp33_ASAP7_75t_L g1662 ( 
.A(n_1637),
.B(n_171),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_1637),
.Y(n_1663)
);

INVx1_ASAP7_75t_L g1664 ( 
.A(n_1637),
.Y(n_1664)
);

INVx1_ASAP7_75t_L g1665 ( 
.A(n_1637),
.Y(n_1665)
);

AND2x2_ASAP7_75t_L g1666 ( 
.A(n_1652),
.B(n_1441),
.Y(n_1666)
);

NOR2xp33_ASAP7_75t_L g1667 ( 
.A(n_1653),
.B(n_173),
.Y(n_1667)
);

INVxp67_ASAP7_75t_L g1668 ( 
.A(n_1655),
.Y(n_1668)
);

NAND2xp5_ASAP7_75t_L g1669 ( 
.A(n_1663),
.B(n_174),
.Y(n_1669)
);

INVxp67_ASAP7_75t_L g1670 ( 
.A(n_1661),
.Y(n_1670)
);

INVx2_ASAP7_75t_L g1671 ( 
.A(n_1664),
.Y(n_1671)
);

AND2x2_ASAP7_75t_L g1672 ( 
.A(n_1656),
.B(n_177),
.Y(n_1672)
);

INVx1_ASAP7_75t_L g1673 ( 
.A(n_1665),
.Y(n_1673)
);

INVx1_ASAP7_75t_L g1674 ( 
.A(n_1658),
.Y(n_1674)
);

AOI21xp33_ASAP7_75t_SL g1675 ( 
.A1(n_1650),
.A2(n_436),
.B(n_178),
.Y(n_1675)
);

INVx1_ASAP7_75t_L g1676 ( 
.A(n_1649),
.Y(n_1676)
);

OR2x2_ASAP7_75t_L g1677 ( 
.A(n_1659),
.B(n_179),
.Y(n_1677)
);

NAND2xp5_ASAP7_75t_L g1678 ( 
.A(n_1672),
.B(n_1659),
.Y(n_1678)
);

NAND2xp5_ASAP7_75t_L g1679 ( 
.A(n_1670),
.B(n_1662),
.Y(n_1679)
);

INVx2_ASAP7_75t_L g1680 ( 
.A(n_1671),
.Y(n_1680)
);

NOR3xp33_ASAP7_75t_L g1681 ( 
.A(n_1668),
.B(n_1654),
.C(n_1660),
.Y(n_1681)
);

INVx1_ASAP7_75t_L g1682 ( 
.A(n_1677),
.Y(n_1682)
);

NAND2xp5_ASAP7_75t_L g1683 ( 
.A(n_1667),
.B(n_1651),
.Y(n_1683)
);

NOR4xp25_ASAP7_75t_L g1684 ( 
.A(n_1673),
.B(n_1657),
.C(n_184),
.D(n_185),
.Y(n_1684)
);

NOR2xp33_ASAP7_75t_L g1685 ( 
.A(n_1674),
.B(n_180),
.Y(n_1685)
);

NOR2x1_ASAP7_75t_L g1686 ( 
.A(n_1669),
.B(n_186),
.Y(n_1686)
);

OAI211xp5_ASAP7_75t_L g1687 ( 
.A1(n_1676),
.A2(n_187),
.B(n_190),
.C(n_191),
.Y(n_1687)
);

NAND2xp5_ASAP7_75t_SL g1688 ( 
.A(n_1684),
.B(n_1675),
.Y(n_1688)
);

AOI211xp5_ASAP7_75t_L g1689 ( 
.A1(n_1681),
.A2(n_1666),
.B(n_198),
.C(n_199),
.Y(n_1689)
);

O2A1O1Ixp5_ASAP7_75t_SL g1690 ( 
.A1(n_1682),
.A2(n_194),
.B(n_200),
.C(n_202),
.Y(n_1690)
);

INVx1_ASAP7_75t_L g1691 ( 
.A(n_1678),
.Y(n_1691)
);

NAND4xp75_ASAP7_75t_L g1692 ( 
.A(n_1686),
.B(n_203),
.C(n_204),
.D(n_205),
.Y(n_1692)
);

A2O1A1O1Ixp25_ASAP7_75t_L g1693 ( 
.A1(n_1679),
.A2(n_206),
.B(n_207),
.C(n_209),
.D(n_213),
.Y(n_1693)
);

A2O1A1Ixp33_ASAP7_75t_L g1694 ( 
.A1(n_1685),
.A2(n_215),
.B(n_216),
.C(n_217),
.Y(n_1694)
);

NOR3x1_ASAP7_75t_L g1695 ( 
.A(n_1683),
.B(n_219),
.C(n_220),
.Y(n_1695)
);

NAND3x1_ASAP7_75t_L g1696 ( 
.A(n_1680),
.B(n_222),
.C(n_224),
.Y(n_1696)
);

NAND2xp5_ASAP7_75t_L g1697 ( 
.A(n_1687),
.B(n_225),
.Y(n_1697)
);

NAND2xp5_ASAP7_75t_L g1698 ( 
.A(n_1682),
.B(n_226),
.Y(n_1698)
);

OAI21xp33_ASAP7_75t_SL g1699 ( 
.A1(n_1678),
.A2(n_227),
.B(n_228),
.Y(n_1699)
);

O2A1O1Ixp33_ASAP7_75t_L g1700 ( 
.A1(n_1678),
.A2(n_229),
.B(n_230),
.C(n_231),
.Y(n_1700)
);

AOI221xp5_ASAP7_75t_L g1701 ( 
.A1(n_1688),
.A2(n_232),
.B1(n_233),
.B2(n_234),
.C(n_236),
.Y(n_1701)
);

INVx1_ASAP7_75t_L g1702 ( 
.A(n_1698),
.Y(n_1702)
);

NAND4xp75_ASAP7_75t_L g1703 ( 
.A(n_1699),
.B(n_240),
.C(n_242),
.D(n_243),
.Y(n_1703)
);

INVx1_ASAP7_75t_L g1704 ( 
.A(n_1691),
.Y(n_1704)
);

AOI22xp5_ASAP7_75t_L g1705 ( 
.A1(n_1697),
.A2(n_245),
.B1(n_246),
.B2(n_248),
.Y(n_1705)
);

AOI22xp33_ASAP7_75t_L g1706 ( 
.A1(n_1693),
.A2(n_249),
.B1(n_250),
.B2(n_252),
.Y(n_1706)
);

NAND2xp5_ASAP7_75t_SL g1707 ( 
.A(n_1689),
.B(n_254),
.Y(n_1707)
);

INVx1_ASAP7_75t_L g1708 ( 
.A(n_1695),
.Y(n_1708)
);

O2A1O1Ixp33_ASAP7_75t_L g1709 ( 
.A1(n_1700),
.A2(n_256),
.B(n_258),
.C(n_259),
.Y(n_1709)
);

INVx2_ASAP7_75t_L g1710 ( 
.A(n_1692),
.Y(n_1710)
);

NAND3xp33_ASAP7_75t_L g1711 ( 
.A(n_1690),
.B(n_260),
.C(n_261),
.Y(n_1711)
);

INVx1_ASAP7_75t_SL g1712 ( 
.A(n_1696),
.Y(n_1712)
);

INVx1_ASAP7_75t_L g1713 ( 
.A(n_1694),
.Y(n_1713)
);

NAND2xp5_ASAP7_75t_L g1714 ( 
.A(n_1695),
.B(n_262),
.Y(n_1714)
);

AOI211xp5_ASAP7_75t_L g1715 ( 
.A1(n_1699),
.A2(n_434),
.B(n_265),
.C(n_266),
.Y(n_1715)
);

NAND4xp75_ASAP7_75t_L g1716 ( 
.A(n_1704),
.B(n_263),
.C(n_267),
.D(n_268),
.Y(n_1716)
);

OR2x2_ASAP7_75t_L g1717 ( 
.A(n_1712),
.B(n_269),
.Y(n_1717)
);

INVx2_ASAP7_75t_L g1718 ( 
.A(n_1703),
.Y(n_1718)
);

NOR2x1_ASAP7_75t_L g1719 ( 
.A(n_1711),
.B(n_270),
.Y(n_1719)
);

NOR2x1_ASAP7_75t_L g1720 ( 
.A(n_1714),
.B(n_430),
.Y(n_1720)
);

OR2x2_ASAP7_75t_L g1721 ( 
.A(n_1708),
.B(n_272),
.Y(n_1721)
);

AND2x2_ASAP7_75t_L g1722 ( 
.A(n_1710),
.B(n_1713),
.Y(n_1722)
);

NOR2xp33_ASAP7_75t_R g1723 ( 
.A(n_1702),
.B(n_273),
.Y(n_1723)
);

AND3x4_ASAP7_75t_L g1724 ( 
.A(n_1715),
.B(n_1707),
.C(n_1706),
.Y(n_1724)
);

NOR3xp33_ASAP7_75t_L g1725 ( 
.A(n_1701),
.B(n_274),
.C(n_276),
.Y(n_1725)
);

INVx1_ASAP7_75t_L g1726 ( 
.A(n_1705),
.Y(n_1726)
);

INVx1_ASAP7_75t_L g1727 ( 
.A(n_1709),
.Y(n_1727)
);

AND2x2_ASAP7_75t_L g1728 ( 
.A(n_1712),
.B(n_278),
.Y(n_1728)
);

OAI21xp33_ASAP7_75t_SL g1729 ( 
.A1(n_1712),
.A2(n_280),
.B(n_281),
.Y(n_1729)
);

NAND2x1_ASAP7_75t_L g1730 ( 
.A(n_1708),
.B(n_284),
.Y(n_1730)
);

NOR3xp33_ASAP7_75t_L g1731 ( 
.A(n_1704),
.B(n_285),
.C(n_286),
.Y(n_1731)
);

AOI21xp5_ASAP7_75t_L g1732 ( 
.A1(n_1707),
.A2(n_287),
.B(n_288),
.Y(n_1732)
);

NOR2x1_ASAP7_75t_L g1733 ( 
.A(n_1703),
.B(n_289),
.Y(n_1733)
);

NOR2xp67_ASAP7_75t_L g1734 ( 
.A(n_1711),
.B(n_428),
.Y(n_1734)
);

NOR3xp33_ASAP7_75t_L g1735 ( 
.A(n_1704),
.B(n_290),
.C(n_292),
.Y(n_1735)
);

NAND2xp33_ASAP7_75t_SL g1736 ( 
.A(n_1730),
.B(n_293),
.Y(n_1736)
);

AOI22xp5_ASAP7_75t_L g1737 ( 
.A1(n_1724),
.A2(n_294),
.B1(n_300),
.B2(n_301),
.Y(n_1737)
);

NAND4xp75_ASAP7_75t_L g1738 ( 
.A(n_1720),
.B(n_303),
.C(n_304),
.D(n_306),
.Y(n_1738)
);

AND3x4_ASAP7_75t_L g1739 ( 
.A(n_1733),
.B(n_308),
.C(n_310),
.Y(n_1739)
);

NOR3xp33_ASAP7_75t_L g1740 ( 
.A(n_1722),
.B(n_313),
.C(n_317),
.Y(n_1740)
);

NAND3xp33_ASAP7_75t_SL g1741 ( 
.A(n_1717),
.B(n_318),
.C(n_319),
.Y(n_1741)
);

NAND2x1_ASAP7_75t_SL g1742 ( 
.A(n_1719),
.B(n_320),
.Y(n_1742)
);

NOR3xp33_ASAP7_75t_L g1743 ( 
.A(n_1729),
.B(n_1728),
.C(n_1727),
.Y(n_1743)
);

AND2x2_ASAP7_75t_L g1744 ( 
.A(n_1718),
.B(n_1734),
.Y(n_1744)
);

INVx1_ASAP7_75t_L g1745 ( 
.A(n_1721),
.Y(n_1745)
);

AOI221xp5_ASAP7_75t_L g1746 ( 
.A1(n_1725),
.A2(n_321),
.B1(n_324),
.B2(n_325),
.C(n_327),
.Y(n_1746)
);

AOI22xp5_ASAP7_75t_L g1747 ( 
.A1(n_1726),
.A2(n_330),
.B1(n_331),
.B2(n_334),
.Y(n_1747)
);

HB1xp67_ASAP7_75t_L g1748 ( 
.A(n_1738),
.Y(n_1748)
);

HB1xp67_ASAP7_75t_L g1749 ( 
.A(n_1739),
.Y(n_1749)
);

NOR2xp67_ASAP7_75t_L g1750 ( 
.A(n_1741),
.B(n_1732),
.Y(n_1750)
);

INVx2_ASAP7_75t_L g1751 ( 
.A(n_1742),
.Y(n_1751)
);

HB1xp67_ASAP7_75t_L g1752 ( 
.A(n_1745),
.Y(n_1752)
);

AOI22xp5_ASAP7_75t_L g1753 ( 
.A1(n_1743),
.A2(n_1735),
.B1(n_1731),
.B2(n_1716),
.Y(n_1753)
);

AND2x4_ASAP7_75t_L g1754 ( 
.A(n_1744),
.B(n_1723),
.Y(n_1754)
);

HB1xp67_ASAP7_75t_L g1755 ( 
.A(n_1740),
.Y(n_1755)
);

OAI22xp5_ASAP7_75t_L g1756 ( 
.A1(n_1753),
.A2(n_1737),
.B1(n_1746),
.B2(n_1747),
.Y(n_1756)
);

NAND2xp5_ASAP7_75t_L g1757 ( 
.A(n_1752),
.B(n_1736),
.Y(n_1757)
);

INVx5_ASAP7_75t_L g1758 ( 
.A(n_1754),
.Y(n_1758)
);

NAND2xp5_ASAP7_75t_L g1759 ( 
.A(n_1749),
.B(n_335),
.Y(n_1759)
);

NAND4xp75_ASAP7_75t_L g1760 ( 
.A(n_1757),
.B(n_1750),
.C(n_1751),
.D(n_1748),
.Y(n_1760)
);

INVx2_ASAP7_75t_L g1761 ( 
.A(n_1758),
.Y(n_1761)
);

OAI322xp33_ASAP7_75t_L g1762 ( 
.A1(n_1761),
.A2(n_1756),
.A3(n_1759),
.B1(n_1755),
.B2(n_343),
.C1(n_344),
.C2(n_347),
.Y(n_1762)
);

OAI21x1_ASAP7_75t_L g1763 ( 
.A1(n_1760),
.A2(n_339),
.B(n_341),
.Y(n_1763)
);

OAI22xp33_ASAP7_75t_L g1764 ( 
.A1(n_1762),
.A2(n_342),
.B1(n_349),
.B2(n_350),
.Y(n_1764)
);

NAND4xp25_ASAP7_75t_L g1765 ( 
.A(n_1763),
.B(n_353),
.C(n_354),
.D(n_356),
.Y(n_1765)
);

INVx1_ASAP7_75t_L g1766 ( 
.A(n_1765),
.Y(n_1766)
);

INVx4_ASAP7_75t_L g1767 ( 
.A(n_1764),
.Y(n_1767)
);

INVx2_ASAP7_75t_L g1768 ( 
.A(n_1767),
.Y(n_1768)
);

OAI22xp5_ASAP7_75t_SL g1769 ( 
.A1(n_1766),
.A2(n_357),
.B1(n_358),
.B2(n_359),
.Y(n_1769)
);

AOI21xp5_ASAP7_75t_L g1770 ( 
.A1(n_1768),
.A2(n_361),
.B(n_363),
.Y(n_1770)
);

OAI22xp5_ASAP7_75t_L g1771 ( 
.A1(n_1769),
.A2(n_364),
.B1(n_367),
.B2(n_369),
.Y(n_1771)
);

OAI31xp33_ASAP7_75t_SL g1772 ( 
.A1(n_1771),
.A2(n_371),
.A3(n_372),
.B(n_373),
.Y(n_1772)
);

OAI222xp33_ASAP7_75t_L g1773 ( 
.A1(n_1770),
.A2(n_376),
.B1(n_377),
.B2(n_378),
.C1(n_379),
.C2(n_381),
.Y(n_1773)
);

OAI21xp5_ASAP7_75t_L g1774 ( 
.A1(n_1771),
.A2(n_383),
.B(n_384),
.Y(n_1774)
);

OAI22xp5_ASAP7_75t_L g1775 ( 
.A1(n_1771),
.A2(n_385),
.B1(n_386),
.B2(n_387),
.Y(n_1775)
);

HB1xp67_ASAP7_75t_L g1776 ( 
.A(n_1774),
.Y(n_1776)
);

INVx4_ASAP7_75t_L g1777 ( 
.A(n_1772),
.Y(n_1777)
);

HB1xp67_ASAP7_75t_L g1778 ( 
.A(n_1775),
.Y(n_1778)
);

NOR3xp33_ASAP7_75t_L g1779 ( 
.A(n_1777),
.B(n_1773),
.C(n_389),
.Y(n_1779)
);

OR2x6_ASAP7_75t_L g1780 ( 
.A(n_1776),
.B(n_388),
.Y(n_1780)
);

AOI221xp5_ASAP7_75t_L g1781 ( 
.A1(n_1778),
.A2(n_390),
.B1(n_391),
.B2(n_394),
.C(n_397),
.Y(n_1781)
);

AOI221xp5_ASAP7_75t_L g1782 ( 
.A1(n_1779),
.A2(n_398),
.B1(n_401),
.B2(n_402),
.C(n_403),
.Y(n_1782)
);

AOI211xp5_ASAP7_75t_L g1783 ( 
.A1(n_1782),
.A2(n_1781),
.B(n_1780),
.C(n_406),
.Y(n_1783)
);


endmodule