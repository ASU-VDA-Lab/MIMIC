module fake_jpeg_12053_n_38 (n_3, n_2, n_1, n_0, n_4, n_5, n_38);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_38;

wire n_13;
wire n_21;
wire n_33;
wire n_10;
wire n_23;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_19;
wire n_20;
wire n_18;
wire n_35;
wire n_34;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_31;
wire n_25;
wire n_29;
wire n_37;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

INVx8_ASAP7_75t_L g6 ( 
.A(n_5),
.Y(n_6)
);

CKINVDCx20_ASAP7_75t_R g7 ( 
.A(n_1),
.Y(n_7)
);

HB1xp67_ASAP7_75t_L g8 ( 
.A(n_1),
.Y(n_8)
);

BUFx6f_ASAP7_75t_L g9 ( 
.A(n_0),
.Y(n_9)
);

INVx3_ASAP7_75t_L g10 ( 
.A(n_5),
.Y(n_10)
);

INVx2_ASAP7_75t_L g11 ( 
.A(n_0),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_0),
.Y(n_12)
);

BUFx12f_ASAP7_75t_L g13 ( 
.A(n_2),
.Y(n_13)
);

OAI22xp5_ASAP7_75t_L g14 ( 
.A1(n_10),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_14)
);

OAI22xp5_ASAP7_75t_L g24 ( 
.A1(n_14),
.A2(n_15),
.B1(n_16),
.B2(n_17),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g15 ( 
.A1(n_11),
.A2(n_3),
.B1(n_4),
.B2(n_9),
.Y(n_15)
);

AO21x1_ASAP7_75t_L g16 ( 
.A1(n_11),
.A2(n_8),
.B(n_7),
.Y(n_16)
);

OR2x4_ASAP7_75t_L g17 ( 
.A(n_13),
.B(n_12),
.Y(n_17)
);

XNOR2xp5_ASAP7_75t_SL g26 ( 
.A(n_17),
.B(n_20),
.Y(n_26)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_18),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_7),
.B(n_13),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_19),
.B(n_21),
.Y(n_25)
);

AND2x2_ASAP7_75t_L g20 ( 
.A(n_13),
.B(n_6),
.Y(n_20)
);

AND2x2_ASAP7_75t_L g21 ( 
.A(n_6),
.B(n_9),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_22),
.B(n_23),
.Y(n_27)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

NAND2xp33_ASAP7_75t_SL g32 ( 
.A(n_24),
.B(n_28),
.Y(n_32)
);

A2O1A1O1Ixp25_ASAP7_75t_L g28 ( 
.A1(n_16),
.A2(n_21),
.B(n_15),
.C(n_20),
.D(n_22),
.Y(n_28)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_29),
.Y(n_30)
);

AOI22xp33_ASAP7_75t_L g34 ( 
.A1(n_30),
.A2(n_31),
.B1(n_25),
.B2(n_26),
.Y(n_34)
);

BUFx12_ASAP7_75t_L g31 ( 
.A(n_29),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_L g33 ( 
.A1(n_32),
.A2(n_28),
.B1(n_27),
.B2(n_26),
.Y(n_33)
);

AOI21xp5_ASAP7_75t_L g35 ( 
.A1(n_33),
.A2(n_34),
.B(n_31),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_35),
.Y(n_36)
);

INVxp67_ASAP7_75t_L g37 ( 
.A(n_36),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_37),
.B(n_34),
.Y(n_38)
);


endmodule