module real_aes_6318_n_101 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_101);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_101;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_578;
wire n_528;
wire n_202;
wire n_495;
wire n_370;
wire n_744;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_178;
wire n_409;
wire n_748;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_310;
wire n_455;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_363;
wire n_182;
wire n_417;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_527;
wire n_502;
wire n_434;
wire n_505;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_402;
wire n_602;
wire n_552;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_633;
wire n_520;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_420;
wire n_336;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_741;
wire n_314;
wire n_283;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_103;
wire n_541;
wire n_166;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
INVx1_ASAP7_75t_L g110 ( .A(n_0), .Y(n_110) );
INVx1_ASAP7_75t_L g495 ( .A(n_1), .Y(n_495) );
INVx1_ASAP7_75t_L g266 ( .A(n_2), .Y(n_266) );
AOI22xp33_ASAP7_75t_L g522 ( .A1(n_3), .A2(n_36), .B1(n_185), .B2(n_523), .Y(n_522) );
AOI21xp33_ASAP7_75t_L g173 ( .A1(n_4), .A2(n_174), .B(n_175), .Y(n_173) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_5), .B(n_172), .Y(n_472) );
AND2x6_ASAP7_75t_L g147 ( .A(n_6), .B(n_148), .Y(n_147) );
AOI21xp5_ASAP7_75t_L g241 ( .A1(n_7), .A2(n_242), .B(n_243), .Y(n_241) );
INVx1_ASAP7_75t_L g107 ( .A(n_8), .Y(n_107) );
NOR2xp33_ASAP7_75t_L g126 ( .A(n_8), .B(n_37), .Y(n_126) );
INVx1_ASAP7_75t_L g182 ( .A(n_9), .Y(n_182) );
NAND2xp5_ASAP7_75t_L g233 ( .A(n_10), .B(n_234), .Y(n_233) );
INVx1_ASAP7_75t_L g144 ( .A(n_11), .Y(n_144) );
INVx1_ASAP7_75t_L g491 ( .A(n_12), .Y(n_491) );
INVx1_ASAP7_75t_L g248 ( .A(n_13), .Y(n_248) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_14), .B(n_150), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_15), .B(n_140), .Y(n_500) );
AO32x2_ASAP7_75t_L g520 ( .A1(n_16), .A2(n_139), .A3(n_172), .B1(n_483), .B2(n_521), .Y(n_520) );
NAND2xp5_ASAP7_75t_SL g532 ( .A(n_17), .B(n_185), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g220 ( .A(n_18), .B(n_193), .Y(n_220) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_19), .B(n_140), .Y(n_497) );
AOI22xp33_ASAP7_75t_L g524 ( .A1(n_20), .A2(n_48), .B1(n_185), .B2(n_523), .Y(n_524) );
NAND2xp5_ASAP7_75t_SL g202 ( .A(n_21), .B(n_174), .Y(n_202) );
AOI22xp33_ASAP7_75t_SL g543 ( .A1(n_22), .A2(n_74), .B1(n_150), .B2(n_185), .Y(n_543) );
NAND2xp5_ASAP7_75t_SL g515 ( .A(n_23), .B(n_185), .Y(n_515) );
NAND2xp5_ASAP7_75t_L g196 ( .A(n_24), .B(n_170), .Y(n_196) );
A2O1A1Ixp33_ASAP7_75t_L g245 ( .A1(n_25), .A2(n_246), .B(n_247), .C(n_249), .Y(n_245) );
BUFx6f_ASAP7_75t_L g155 ( .A(n_26), .Y(n_155) );
NAND2xp5_ASAP7_75t_L g484 ( .A(n_27), .B(n_187), .Y(n_484) );
NAND2xp5_ASAP7_75t_L g267 ( .A(n_28), .B(n_180), .Y(n_267) );
INVx1_ASAP7_75t_L g158 ( .A(n_29), .Y(n_158) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_30), .B(n_187), .Y(n_517) );
INVx2_ASAP7_75t_L g152 ( .A(n_31), .Y(n_152) );
NAND2xp5_ASAP7_75t_SL g477 ( .A(n_32), .B(n_185), .Y(n_477) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_33), .B(n_187), .Y(n_534) );
AOI22xp5_ASAP7_75t_L g129 ( .A1(n_34), .A2(n_40), .B1(n_130), .B2(n_131), .Y(n_129) );
CKINVDCx20_ASAP7_75t_R g131 ( .A(n_34), .Y(n_131) );
A2O1A1Ixp33_ASAP7_75t_L g203 ( .A1(n_35), .A2(n_147), .B(n_159), .C(n_204), .Y(n_203) );
NAND2xp5_ASAP7_75t_L g106 ( .A(n_37), .B(n_107), .Y(n_106) );
INVx1_ASAP7_75t_L g156 ( .A(n_38), .Y(n_156) );
NAND2xp5_ASAP7_75t_SL g219 ( .A(n_39), .B(n_180), .Y(n_219) );
CKINVDCx20_ASAP7_75t_R g130 ( .A(n_40), .Y(n_130) );
NAND2xp5_ASAP7_75t_SL g465 ( .A(n_41), .B(n_185), .Y(n_465) );
AOI22xp33_ASAP7_75t_L g542 ( .A1(n_42), .A2(n_87), .B1(n_210), .B2(n_523), .Y(n_542) );
NAND2xp5_ASAP7_75t_SL g468 ( .A(n_43), .B(n_185), .Y(n_468) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_44), .B(n_185), .Y(n_492) );
CKINVDCx16_ASAP7_75t_R g162 ( .A(n_45), .Y(n_162) );
NAND2xp5_ASAP7_75t_L g469 ( .A(n_46), .B(n_470), .Y(n_469) );
NAND2xp5_ASAP7_75t_L g236 ( .A(n_47), .B(n_174), .Y(n_236) );
AOI22xp33_ASAP7_75t_SL g504 ( .A1(n_49), .A2(n_59), .B1(n_150), .B2(n_185), .Y(n_504) );
AOI22xp5_ASAP7_75t_L g149 ( .A1(n_50), .A2(n_150), .B1(n_153), .B2(n_159), .Y(n_149) );
CKINVDCx20_ASAP7_75t_R g213 ( .A(n_51), .Y(n_213) );
NAND2xp5_ASAP7_75t_SL g482 ( .A(n_52), .B(n_185), .Y(n_482) );
CKINVDCx16_ASAP7_75t_R g263 ( .A(n_53), .Y(n_263) );
NAND2xp5_ASAP7_75t_SL g528 ( .A(n_54), .B(n_185), .Y(n_528) );
A2O1A1Ixp33_ASAP7_75t_L g178 ( .A1(n_55), .A2(n_179), .B(n_181), .C(n_184), .Y(n_178) );
AOI22xp33_ASAP7_75t_L g101 ( .A1(n_56), .A2(n_102), .B1(n_115), .B2(n_748), .Y(n_101) );
CKINVDCx20_ASAP7_75t_R g223 ( .A(n_57), .Y(n_223) );
INVx1_ASAP7_75t_L g176 ( .A(n_58), .Y(n_176) );
INVx1_ASAP7_75t_L g148 ( .A(n_60), .Y(n_148) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_61), .B(n_185), .Y(n_496) );
INVx1_ASAP7_75t_L g143 ( .A(n_62), .Y(n_143) );
CKINVDCx20_ASAP7_75t_R g120 ( .A(n_63), .Y(n_120) );
AO32x2_ASAP7_75t_L g540 ( .A1(n_64), .A2(n_172), .A3(n_228), .B1(n_483), .B2(n_541), .Y(n_540) );
INVx1_ASAP7_75t_L g480 ( .A(n_65), .Y(n_480) );
INVx1_ASAP7_75t_L g512 ( .A(n_66), .Y(n_512) );
A2O1A1Ixp33_ASAP7_75t_SL g192 ( .A1(n_67), .A2(n_184), .B(n_193), .C(n_194), .Y(n_192) );
INVxp67_ASAP7_75t_L g195 ( .A(n_68), .Y(n_195) );
NAND2xp5_ASAP7_75t_SL g513 ( .A(n_69), .B(n_150), .Y(n_513) );
INVx1_ASAP7_75t_L g114 ( .A(n_70), .Y(n_114) );
CKINVDCx20_ASAP7_75t_R g167 ( .A(n_71), .Y(n_167) );
INVx1_ASAP7_75t_L g216 ( .A(n_72), .Y(n_216) );
OAI22xp5_ASAP7_75t_L g738 ( .A1(n_73), .A2(n_99), .B1(n_739), .B2(n_740), .Y(n_738) );
CKINVDCx20_ASAP7_75t_R g739 ( .A(n_73), .Y(n_739) );
A2O1A1Ixp33_ASAP7_75t_L g217 ( .A1(n_75), .A2(n_147), .B(n_159), .C(n_218), .Y(n_217) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_76), .B(n_523), .Y(n_533) );
NAND2xp5_ASAP7_75t_SL g516 ( .A(n_77), .B(n_150), .Y(n_516) );
NAND2xp5_ASAP7_75t_SL g205 ( .A(n_78), .B(n_206), .Y(n_205) );
INVx2_ASAP7_75t_L g141 ( .A(n_79), .Y(n_141) );
NAND2xp5_ASAP7_75t_L g207 ( .A(n_80), .B(n_193), .Y(n_207) );
AOI222xp33_ASAP7_75t_L g449 ( .A1(n_81), .A2(n_450), .B1(n_738), .B2(n_741), .C1(n_742), .C2(n_744), .Y(n_449) );
NAND2xp5_ASAP7_75t_L g466 ( .A(n_82), .B(n_150), .Y(n_466) );
A2O1A1Ixp33_ASAP7_75t_L g264 ( .A1(n_83), .A2(n_147), .B(n_159), .C(n_265), .Y(n_264) );
INVx2_ASAP7_75t_L g111 ( .A(n_84), .Y(n_111) );
OR2x2_ASAP7_75t_L g123 ( .A(n_84), .B(n_124), .Y(n_123) );
OR2x2_ASAP7_75t_L g453 ( .A(n_84), .B(n_125), .Y(n_453) );
NAND2xp5_ASAP7_75t_L g445 ( .A(n_85), .B(n_446), .Y(n_445) );
AOI22xp33_ASAP7_75t_L g503 ( .A1(n_86), .A2(n_100), .B1(n_150), .B2(n_151), .Y(n_503) );
NAND2xp5_ASAP7_75t_L g186 ( .A(n_88), .B(n_187), .Y(n_186) );
CKINVDCx20_ASAP7_75t_R g270 ( .A(n_89), .Y(n_270) );
A2O1A1Ixp33_ASAP7_75t_L g230 ( .A1(n_90), .A2(n_147), .B(n_159), .C(n_231), .Y(n_230) );
CKINVDCx20_ASAP7_75t_R g238 ( .A(n_91), .Y(n_238) );
INVx1_ASAP7_75t_L g191 ( .A(n_92), .Y(n_191) );
CKINVDCx16_ASAP7_75t_R g244 ( .A(n_93), .Y(n_244) );
NAND2xp5_ASAP7_75t_SL g232 ( .A(n_94), .B(n_206), .Y(n_232) );
NAND2xp5_ASAP7_75t_L g478 ( .A(n_95), .B(n_150), .Y(n_478) );
NAND2xp5_ASAP7_75t_L g250 ( .A(n_96), .B(n_172), .Y(n_250) );
NAND2xp5_ASAP7_75t_L g113 ( .A(n_97), .B(n_114), .Y(n_113) );
AOI21xp5_ASAP7_75t_L g189 ( .A1(n_98), .A2(n_174), .B(n_190), .Y(n_189) );
CKINVDCx16_ASAP7_75t_R g740 ( .A(n_99), .Y(n_740) );
CKINVDCx20_ASAP7_75t_R g102 ( .A(n_103), .Y(n_102) );
CKINVDCx16_ASAP7_75t_R g103 ( .A(n_104), .Y(n_103) );
INVx2_ASAP7_75t_L g750 ( .A(n_104), .Y(n_750) );
AND2x2_ASAP7_75t_L g104 ( .A(n_105), .B(n_108), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
CKINVDCx14_ASAP7_75t_R g108 ( .A(n_109), .Y(n_108) );
NAND3xp33_ASAP7_75t_SL g109 ( .A(n_110), .B(n_111), .C(n_112), .Y(n_109) );
AND2x2_ASAP7_75t_L g125 ( .A(n_110), .B(n_126), .Y(n_125) );
OR2x2_ASAP7_75t_L g737 ( .A(n_111), .B(n_125), .Y(n_737) );
NOR2x2_ASAP7_75t_L g746 ( .A(n_111), .B(n_124), .Y(n_746) );
INVx1_ASAP7_75t_SL g112 ( .A(n_113), .Y(n_112) );
OA21x2_ASAP7_75t_L g115 ( .A1(n_116), .A2(n_121), .B(n_448), .Y(n_115) );
BUFx2_ASAP7_75t_SL g116 ( .A(n_117), .Y(n_116) );
CKINVDCx20_ASAP7_75t_R g117 ( .A(n_118), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
INVx2_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
INVx1_ASAP7_75t_L g747 ( .A(n_120), .Y(n_747) );
OAI21xp5_ASAP7_75t_L g121 ( .A1(n_122), .A2(n_127), .B(n_445), .Y(n_121) );
INVx1_ASAP7_75t_SL g122 ( .A(n_123), .Y(n_122) );
BUFx2_ASAP7_75t_L g447 ( .A(n_123), .Y(n_447) );
INVx2_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
AOI22xp33_ASAP7_75t_L g127 ( .A1(n_128), .A2(n_129), .B1(n_132), .B2(n_444), .Y(n_127) );
CKINVDCx20_ASAP7_75t_R g128 ( .A(n_129), .Y(n_128) );
INVx1_ASAP7_75t_L g444 ( .A(n_132), .Y(n_444) );
OAI22xp5_ASAP7_75t_SL g450 ( .A1(n_132), .A2(n_451), .B1(n_454), .B2(n_735), .Y(n_450) );
AND3x1_ASAP7_75t_L g132 ( .A(n_133), .B(n_369), .C(n_418), .Y(n_132) );
NOR3xp33_ASAP7_75t_SL g133 ( .A(n_134), .B(n_276), .C(n_314), .Y(n_133) );
OAI222xp33_ASAP7_75t_L g134 ( .A1(n_135), .A2(n_197), .B1(n_251), .B2(n_257), .C1(n_271), .C2(n_274), .Y(n_134) );
NAND2xp5_ASAP7_75t_L g135 ( .A(n_136), .B(n_168), .Y(n_135) );
NAND2xp5_ASAP7_75t_L g343 ( .A(n_136), .B(n_344), .Y(n_343) );
NAND2xp5_ASAP7_75t_L g410 ( .A(n_136), .B(n_319), .Y(n_410) );
BUFx2_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
OR2x2_ASAP7_75t_L g287 ( .A(n_137), .B(n_188), .Y(n_287) );
NAND2xp5_ASAP7_75t_L g295 ( .A(n_137), .B(n_169), .Y(n_295) );
AND2x2_ASAP7_75t_L g330 ( .A(n_137), .B(n_307), .Y(n_330) );
OR2x2_ASAP7_75t_L g354 ( .A(n_137), .B(n_169), .Y(n_354) );
OR2x2_ASAP7_75t_L g362 ( .A(n_137), .B(n_261), .Y(n_362) );
AND2x2_ASAP7_75t_L g365 ( .A(n_137), .B(n_188), .Y(n_365) );
INVx3_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
OR2x2_ASAP7_75t_L g259 ( .A(n_138), .B(n_260), .Y(n_259) );
AND2x2_ASAP7_75t_L g273 ( .A(n_138), .B(n_188), .Y(n_273) );
AND2x2_ASAP7_75t_L g323 ( .A(n_138), .B(n_261), .Y(n_323) );
AND2x2_ASAP7_75t_L g336 ( .A(n_138), .B(n_169), .Y(n_336) );
NOR2xp33_ASAP7_75t_L g443 ( .A(n_138), .B(n_422), .Y(n_443) );
AO21x2_ASAP7_75t_L g138 ( .A1(n_139), .A2(n_145), .B(n_166), .Y(n_138) );
NOR2xp33_ASAP7_75t_L g166 ( .A(n_139), .B(n_167), .Y(n_166) );
INVx2_ASAP7_75t_L g211 ( .A(n_139), .Y(n_211) );
AO21x2_ASAP7_75t_L g261 ( .A1(n_139), .A2(n_262), .B(n_269), .Y(n_261) );
INVx1_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
BUFx6f_ASAP7_75t_L g172 ( .A(n_140), .Y(n_172) );
AND2x2_ASAP7_75t_L g140 ( .A(n_141), .B(n_142), .Y(n_140) );
AND2x2_ASAP7_75t_SL g187 ( .A(n_141), .B(n_142), .Y(n_187) );
NAND2xp5_ASAP7_75t_L g142 ( .A(n_143), .B(n_144), .Y(n_142) );
OAI22xp33_ASAP7_75t_L g145 ( .A1(n_146), .A2(n_149), .B1(n_162), .B2(n_163), .Y(n_145) );
O2A1O1Ixp33_ASAP7_75t_L g175 ( .A1(n_146), .A2(n_176), .B(n_177), .C(n_178), .Y(n_175) );
O2A1O1Ixp33_ASAP7_75t_L g190 ( .A1(n_146), .A2(n_177), .B(n_191), .C(n_192), .Y(n_190) );
O2A1O1Ixp33_ASAP7_75t_L g243 ( .A1(n_146), .A2(n_177), .B(n_244), .C(n_245), .Y(n_243) );
INVx4_ASAP7_75t_SL g146 ( .A(n_147), .Y(n_146) );
NAND2x1p5_ASAP7_75t_L g163 ( .A(n_147), .B(n_164), .Y(n_163) );
AND2x4_ASAP7_75t_L g174 ( .A(n_147), .B(n_164), .Y(n_174) );
OAI21xp5_ASAP7_75t_L g463 ( .A1(n_147), .A2(n_464), .B(n_467), .Y(n_463) );
BUFx3_ASAP7_75t_L g483 ( .A(n_147), .Y(n_483) );
OAI21xp5_ASAP7_75t_L g489 ( .A1(n_147), .A2(n_490), .B(n_494), .Y(n_489) );
OAI21xp5_ASAP7_75t_L g510 ( .A1(n_147), .A2(n_511), .B(n_514), .Y(n_510) );
OAI21xp5_ASAP7_75t_L g526 ( .A1(n_147), .A2(n_527), .B(n_531), .Y(n_526) );
INVx2_ASAP7_75t_L g268 ( .A(n_150), .Y(n_268) );
INVx3_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
INVx1_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
INVx2_ASAP7_75t_L g160 ( .A(n_152), .Y(n_160) );
INVx1_ASAP7_75t_L g165 ( .A(n_152), .Y(n_165) );
OAI22xp5_ASAP7_75t_SL g153 ( .A1(n_154), .A2(n_156), .B1(n_157), .B2(n_158), .Y(n_153) );
INVx2_ASAP7_75t_L g157 ( .A(n_154), .Y(n_157) );
INVx4_ASAP7_75t_L g246 ( .A(n_154), .Y(n_246) );
BUFx6f_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
INVx1_ASAP7_75t_L g161 ( .A(n_155), .Y(n_161) );
AND2x2_ASAP7_75t_L g164 ( .A(n_155), .B(n_165), .Y(n_164) );
BUFx6f_ASAP7_75t_L g180 ( .A(n_155), .Y(n_180) );
INVx3_ASAP7_75t_L g183 ( .A(n_155), .Y(n_183) );
INVx1_ASAP7_75t_L g193 ( .A(n_155), .Y(n_193) );
INVx5_ASAP7_75t_L g177 ( .A(n_159), .Y(n_177) );
AND2x6_ASAP7_75t_L g159 ( .A(n_160), .B(n_161), .Y(n_159) );
BUFx6f_ASAP7_75t_L g185 ( .A(n_160), .Y(n_185) );
BUFx3_ASAP7_75t_L g210 ( .A(n_160), .Y(n_210) );
INVx1_ASAP7_75t_L g523 ( .A(n_160), .Y(n_523) );
OAI21xp5_ASAP7_75t_L g215 ( .A1(n_163), .A2(n_216), .B(n_217), .Y(n_215) );
OAI21xp5_ASAP7_75t_L g262 ( .A1(n_163), .A2(n_263), .B(n_264), .Y(n_262) );
INVx1_ASAP7_75t_L g470 ( .A(n_165), .Y(n_470) );
O2A1O1Ixp33_ASAP7_75t_L g361 ( .A1(n_168), .A2(n_362), .B(n_363), .C(n_366), .Y(n_361) );
NAND2xp5_ASAP7_75t_L g390 ( .A(n_168), .B(n_391), .Y(n_390) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_168), .B(n_306), .Y(n_428) );
AND2x2_ASAP7_75t_L g168 ( .A(n_169), .B(n_188), .Y(n_168) );
AND2x2_ASAP7_75t_SL g272 ( .A(n_169), .B(n_273), .Y(n_272) );
INVx2_ASAP7_75t_L g286 ( .A(n_169), .Y(n_286) );
AND2x2_ASAP7_75t_L g313 ( .A(n_169), .B(n_307), .Y(n_313) );
INVx1_ASAP7_75t_SL g321 ( .A(n_169), .Y(n_321) );
AND2x2_ASAP7_75t_L g344 ( .A(n_169), .B(n_345), .Y(n_344) );
BUFx2_ASAP7_75t_L g422 ( .A(n_169), .Y(n_422) );
OA21x2_ASAP7_75t_L g169 ( .A1(n_170), .A2(n_173), .B(n_186), .Y(n_169) );
INVx3_ASAP7_75t_L g170 ( .A(n_171), .Y(n_170) );
NOR2xp33_ASAP7_75t_SL g212 ( .A(n_171), .B(n_213), .Y(n_212) );
NAND3xp33_ASAP7_75t_L g501 ( .A(n_171), .B(n_483), .C(n_502), .Y(n_501) );
AO21x1_ASAP7_75t_L g546 ( .A1(n_171), .A2(n_502), .B(n_547), .Y(n_546) );
INVx4_ASAP7_75t_L g171 ( .A(n_172), .Y(n_171) );
OA21x2_ASAP7_75t_L g188 ( .A1(n_172), .A2(n_189), .B(n_196), .Y(n_188) );
OA21x2_ASAP7_75t_L g462 ( .A1(n_172), .A2(n_463), .B(n_472), .Y(n_462) );
BUFx2_ASAP7_75t_L g242 ( .A(n_174), .Y(n_242) );
O2A1O1Ixp5_ASAP7_75t_L g479 ( .A1(n_179), .A2(n_480), .B(n_481), .C(n_482), .Y(n_479) );
AOI21xp5_ASAP7_75t_L g531 ( .A1(n_179), .A2(n_532), .B(n_533), .Y(n_531) );
INVx2_ASAP7_75t_L g179 ( .A(n_180), .Y(n_179) );
INVx4_ASAP7_75t_L g234 ( .A(n_180), .Y(n_234) );
OAI22xp5_ASAP7_75t_L g502 ( .A1(n_180), .A2(n_471), .B1(n_503), .B2(n_504), .Y(n_502) );
OAI22xp5_ASAP7_75t_L g521 ( .A1(n_180), .A2(n_471), .B1(n_522), .B2(n_524), .Y(n_521) );
OAI22xp5_ASAP7_75t_SL g541 ( .A1(n_180), .A2(n_183), .B1(n_542), .B2(n_543), .Y(n_541) );
NOR2xp33_ASAP7_75t_L g181 ( .A(n_182), .B(n_183), .Y(n_181) );
NOR2xp33_ASAP7_75t_L g194 ( .A(n_183), .B(n_195), .Y(n_194) );
INVx5_ASAP7_75t_L g206 ( .A(n_183), .Y(n_206) );
O2A1O1Ixp5_ASAP7_75t_SL g511 ( .A1(n_184), .A2(n_206), .B(n_512), .C(n_513), .Y(n_511) );
INVx3_ASAP7_75t_L g184 ( .A(n_185), .Y(n_184) );
HB1xp67_ASAP7_75t_L g235 ( .A(n_185), .Y(n_235) );
INVx1_ASAP7_75t_L g224 ( .A(n_187), .Y(n_224) );
INVx2_ASAP7_75t_L g228 ( .A(n_187), .Y(n_228) );
OA21x2_ASAP7_75t_L g240 ( .A1(n_187), .A2(n_241), .B(n_250), .Y(n_240) );
OA21x2_ASAP7_75t_L g509 ( .A1(n_187), .A2(n_510), .B(n_517), .Y(n_509) );
OA21x2_ASAP7_75t_L g525 ( .A1(n_187), .A2(n_526), .B(n_534), .Y(n_525) );
BUFx2_ASAP7_75t_L g258 ( .A(n_188), .Y(n_258) );
INVx1_ASAP7_75t_L g320 ( .A(n_188), .Y(n_320) );
INVx3_ASAP7_75t_L g345 ( .A(n_188), .Y(n_345) );
INVx1_ASAP7_75t_L g530 ( .A(n_193), .Y(n_530) );
NAND2xp5_ASAP7_75t_SL g278 ( .A(n_197), .B(n_279), .Y(n_278) );
OR2x2_ASAP7_75t_L g197 ( .A(n_198), .B(n_225), .Y(n_197) );
INVx1_ASAP7_75t_L g341 ( .A(n_198), .Y(n_341) );
OAI32xp33_ASAP7_75t_L g347 ( .A1(n_198), .A2(n_286), .A3(n_348), .B1(n_349), .B2(n_350), .Y(n_347) );
OAI22xp5_ASAP7_75t_L g351 ( .A1(n_198), .A2(n_352), .B1(n_355), .B2(n_360), .Y(n_351) );
INVx4_ASAP7_75t_L g198 ( .A(n_199), .Y(n_198) );
AND2x2_ASAP7_75t_L g289 ( .A(n_199), .B(n_290), .Y(n_289) );
AND2x2_ASAP7_75t_L g367 ( .A(n_199), .B(n_368), .Y(n_367) );
AND2x2_ASAP7_75t_L g437 ( .A(n_199), .B(n_383), .Y(n_437) );
AND2x2_ASAP7_75t_L g199 ( .A(n_200), .B(n_214), .Y(n_199) );
AND2x2_ASAP7_75t_L g252 ( .A(n_200), .B(n_253), .Y(n_252) );
INVx2_ASAP7_75t_L g282 ( .A(n_200), .Y(n_282) );
INVx1_ASAP7_75t_L g301 ( .A(n_200), .Y(n_301) );
OR2x2_ASAP7_75t_L g309 ( .A(n_200), .B(n_310), .Y(n_309) );
AND2x2_ASAP7_75t_L g316 ( .A(n_200), .B(n_290), .Y(n_316) );
NOR2xp33_ASAP7_75t_L g324 ( .A(n_200), .B(n_325), .Y(n_324) );
AND2x2_ASAP7_75t_L g337 ( .A(n_200), .B(n_255), .Y(n_337) );
INVx3_ASAP7_75t_L g359 ( .A(n_200), .Y(n_359) );
AND2x2_ASAP7_75t_L g384 ( .A(n_200), .B(n_256), .Y(n_384) );
NOR2xp33_ASAP7_75t_L g432 ( .A(n_200), .B(n_349), .Y(n_432) );
OR2x6_ASAP7_75t_L g200 ( .A(n_201), .B(n_212), .Y(n_200) );
AOI21xp5_ASAP7_75t_SL g201 ( .A1(n_202), .A2(n_203), .B(n_211), .Y(n_201) );
AOI21xp5_ASAP7_75t_L g204 ( .A1(n_205), .A2(n_207), .B(n_208), .Y(n_204) );
O2A1O1Ixp33_ASAP7_75t_L g265 ( .A1(n_206), .A2(n_266), .B(n_267), .C(n_268), .Y(n_265) );
AOI21xp5_ASAP7_75t_L g464 ( .A1(n_206), .A2(n_465), .B(n_466), .Y(n_464) );
INVx2_ASAP7_75t_L g471 ( .A(n_206), .Y(n_471) );
AOI21xp5_ASAP7_75t_L g476 ( .A1(n_206), .A2(n_477), .B(n_478), .Y(n_476) );
AOI21xp5_ASAP7_75t_L g218 ( .A1(n_208), .A2(n_219), .B(n_220), .Y(n_218) );
INVx2_ASAP7_75t_L g208 ( .A(n_209), .Y(n_208) );
INVx2_ASAP7_75t_L g209 ( .A(n_210), .Y(n_209) );
INVx1_ASAP7_75t_L g249 ( .A(n_210), .Y(n_249) );
INVx1_ASAP7_75t_L g221 ( .A(n_211), .Y(n_221) );
OA21x2_ASAP7_75t_L g474 ( .A1(n_211), .A2(n_475), .B(n_484), .Y(n_474) );
OA21x2_ASAP7_75t_L g488 ( .A1(n_211), .A2(n_489), .B(n_497), .Y(n_488) );
INVx2_ASAP7_75t_L g256 ( .A(n_214), .Y(n_256) );
AND2x2_ASAP7_75t_L g388 ( .A(n_214), .B(n_226), .Y(n_388) );
AO21x2_ASAP7_75t_L g214 ( .A1(n_215), .A2(n_221), .B(n_222), .Y(n_214) );
NOR2xp33_ASAP7_75t_L g222 ( .A(n_223), .B(n_224), .Y(n_222) );
NOR2xp33_ASAP7_75t_L g237 ( .A(n_224), .B(n_238), .Y(n_237) );
NOR2xp33_ASAP7_75t_L g269 ( .A(n_224), .B(n_270), .Y(n_269) );
INVx2_ASAP7_75t_L g430 ( .A(n_225), .Y(n_430) );
OR2x2_ASAP7_75t_L g225 ( .A(n_226), .B(n_239), .Y(n_225) );
INVx1_ASAP7_75t_L g275 ( .A(n_226), .Y(n_275) );
AND2x2_ASAP7_75t_L g302 ( .A(n_226), .B(n_303), .Y(n_302) );
NAND2xp5_ASAP7_75t_L g310 ( .A(n_226), .B(n_256), .Y(n_310) );
AND2x2_ASAP7_75t_L g368 ( .A(n_226), .B(n_291), .Y(n_368) );
INVx2_ASAP7_75t_L g226 ( .A(n_227), .Y(n_226) );
INVx1_ASAP7_75t_L g254 ( .A(n_227), .Y(n_254) );
AND2x2_ASAP7_75t_L g281 ( .A(n_227), .B(n_282), .Y(n_281) );
AND2x2_ASAP7_75t_L g290 ( .A(n_227), .B(n_291), .Y(n_290) );
NAND2xp5_ASAP7_75t_L g356 ( .A(n_227), .B(n_256), .Y(n_356) );
AO21x2_ASAP7_75t_L g227 ( .A1(n_228), .A2(n_229), .B(n_237), .Y(n_227) );
NAND2xp5_ASAP7_75t_L g229 ( .A(n_230), .B(n_236), .Y(n_229) );
AOI21xp5_ASAP7_75t_L g231 ( .A1(n_232), .A2(n_233), .B(n_235), .Y(n_231) );
NAND2xp5_ASAP7_75t_L g283 ( .A(n_239), .B(n_284), .Y(n_283) );
INVx2_ASAP7_75t_L g303 ( .A(n_239), .Y(n_303) );
NAND2xp5_ASAP7_75t_L g349 ( .A(n_239), .B(n_256), .Y(n_349) );
AND2x2_ASAP7_75t_L g358 ( .A(n_239), .B(n_359), .Y(n_358) );
INVx1_ASAP7_75t_L g383 ( .A(n_239), .Y(n_383) );
INVx2_ASAP7_75t_L g239 ( .A(n_240), .Y(n_239) );
AND2x2_ASAP7_75t_L g255 ( .A(n_240), .B(n_256), .Y(n_255) );
INVx1_ASAP7_75t_L g291 ( .A(n_240), .Y(n_291) );
NOR2xp33_ASAP7_75t_L g247 ( .A(n_246), .B(n_248), .Y(n_247) );
INVx1_ASAP7_75t_L g493 ( .A(n_246), .Y(n_493) );
AOI21xp5_ASAP7_75t_L g514 ( .A1(n_246), .A2(n_515), .B(n_516), .Y(n_514) );
OAI22xp5_ASAP7_75t_L g419 ( .A1(n_251), .A2(n_261), .B1(n_420), .B2(n_423), .Y(n_419) );
INVx1_ASAP7_75t_SL g251 ( .A(n_252), .Y(n_251) );
OAI21xp5_ASAP7_75t_SL g442 ( .A1(n_253), .A2(n_364), .B(n_443), .Y(n_442) );
AND2x2_ASAP7_75t_L g253 ( .A(n_254), .B(n_255), .Y(n_253) );
NOR2xp33_ASAP7_75t_L g376 ( .A(n_254), .B(n_359), .Y(n_376) );
INVx1_ASAP7_75t_L g401 ( .A(n_254), .Y(n_401) );
NAND2xp5_ASAP7_75t_L g274 ( .A(n_255), .B(n_275), .Y(n_274) );
AND2x2_ASAP7_75t_L g328 ( .A(n_255), .B(n_281), .Y(n_328) );
INVx2_ASAP7_75t_L g284 ( .A(n_256), .Y(n_284) );
INVx1_ASAP7_75t_L g334 ( .A(n_256), .Y(n_334) );
OAI221xp5_ASAP7_75t_L g425 ( .A1(n_257), .A2(n_409), .B1(n_426), .B2(n_429), .C(n_431), .Y(n_425) );
OR2x2_ASAP7_75t_L g257 ( .A(n_258), .B(n_259), .Y(n_257) );
INVx1_ASAP7_75t_L g296 ( .A(n_258), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g348 ( .A(n_258), .B(n_307), .Y(n_348) );
NOR2xp33_ASAP7_75t_L g317 ( .A(n_259), .B(n_318), .Y(n_317) );
OR2x2_ASAP7_75t_L g350 ( .A(n_259), .B(n_296), .Y(n_350) );
INVx3_ASAP7_75t_SL g391 ( .A(n_259), .Y(n_391) );
AND2x2_ASAP7_75t_L g335 ( .A(n_260), .B(n_336), .Y(n_335) );
AND2x2_ASAP7_75t_L g364 ( .A(n_260), .B(n_365), .Y(n_364) );
NAND2xp5_ASAP7_75t_L g379 ( .A(n_260), .B(n_273), .Y(n_379) );
NAND2xp5_ASAP7_75t_L g405 ( .A(n_260), .B(n_319), .Y(n_405) );
INVx3_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
INVx3_ASAP7_75t_L g307 ( .A(n_261), .Y(n_307) );
OAI322xp33_ASAP7_75t_L g402 ( .A1(n_261), .A2(n_333), .A3(n_355), .B1(n_403), .B2(n_405), .C1(n_406), .C2(n_407), .Y(n_402) );
O2A1O1Ixp33_ASAP7_75t_L g490 ( .A1(n_268), .A2(n_491), .B(n_492), .C(n_493), .Y(n_490) );
INVx1_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
AOI21xp33_ASAP7_75t_L g426 ( .A1(n_272), .A2(n_275), .B(n_427), .Y(n_426) );
NOR2xp33_ASAP7_75t_SL g352 ( .A(n_273), .B(n_353), .Y(n_352) );
AND2x2_ASAP7_75t_L g374 ( .A(n_273), .B(n_286), .Y(n_374) );
NAND2xp5_ASAP7_75t_L g389 ( .A(n_273), .B(n_313), .Y(n_389) );
INVxp67_ASAP7_75t_L g340 ( .A(n_275), .Y(n_340) );
AOI211xp5_ASAP7_75t_L g346 ( .A1(n_275), .A2(n_347), .B(n_351), .C(n_361), .Y(n_346) );
OAI221xp5_ASAP7_75t_SL g276 ( .A1(n_277), .A2(n_285), .B1(n_288), .B2(n_292), .C(n_297), .Y(n_276) );
INVxp67_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
OR2x2_ASAP7_75t_L g279 ( .A(n_280), .B(n_283), .Y(n_279) );
INVx1_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
AND2x2_ASAP7_75t_L g300 ( .A(n_284), .B(n_301), .Y(n_300) );
INVx1_ASAP7_75t_L g417 ( .A(n_284), .Y(n_417) );
OAI221xp5_ASAP7_75t_L g433 ( .A1(n_285), .A2(n_434), .B1(n_439), .B2(n_440), .C(n_442), .Y(n_433) );
OR2x2_ASAP7_75t_L g285 ( .A(n_286), .B(n_287), .Y(n_285) );
NAND2xp5_ASAP7_75t_L g329 ( .A(n_286), .B(n_330), .Y(n_329) );
INVx1_ASAP7_75t_SL g333 ( .A(n_286), .Y(n_333) );
NAND2xp5_ASAP7_75t_L g371 ( .A(n_286), .B(n_364), .Y(n_371) );
AND2x2_ASAP7_75t_L g413 ( .A(n_286), .B(n_391), .Y(n_413) );
NOR2xp33_ASAP7_75t_L g311 ( .A(n_287), .B(n_312), .Y(n_311) );
OAI22xp33_ASAP7_75t_L g408 ( .A1(n_287), .A2(n_299), .B1(n_409), .B2(n_410), .Y(n_408) );
OR2x2_ASAP7_75t_L g439 ( .A(n_287), .B(n_307), .Y(n_439) );
CKINVDCx16_ASAP7_75t_R g288 ( .A(n_289), .Y(n_288) );
INVx1_ASAP7_75t_L g416 ( .A(n_290), .Y(n_416) );
AND2x2_ASAP7_75t_L g441 ( .A(n_290), .B(n_384), .Y(n_441) );
INVxp67_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
NOR2xp33_ASAP7_75t_SL g293 ( .A(n_294), .B(n_296), .Y(n_293) );
INVx1_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
OR2x2_ASAP7_75t_L g305 ( .A(n_295), .B(n_306), .Y(n_305) );
AOI22xp5_ASAP7_75t_L g297 ( .A1(n_298), .A2(n_304), .B1(n_308), .B2(n_311), .Y(n_297) );
INVx1_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
NAND2xp5_ASAP7_75t_L g299 ( .A(n_300), .B(n_302), .Y(n_299) );
INVx1_ASAP7_75t_L g372 ( .A(n_300), .Y(n_372) );
NAND2xp5_ASAP7_75t_L g407 ( .A(n_300), .B(n_340), .Y(n_407) );
AOI322xp5_ASAP7_75t_L g331 ( .A1(n_302), .A2(n_332), .A3(n_334), .B1(n_335), .B2(n_337), .C1(n_338), .C2(n_342), .Y(n_331) );
INVxp67_ASAP7_75t_L g325 ( .A(n_303), .Y(n_325) );
INVx1_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
OAI22xp5_ASAP7_75t_L g326 ( .A1(n_305), .A2(n_310), .B1(n_327), .B2(n_329), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g406 ( .A(n_306), .B(n_319), .Y(n_406) );
INVx1_ASAP7_75t_SL g306 ( .A(n_307), .Y(n_306) );
NOR2xp33_ASAP7_75t_L g415 ( .A(n_307), .B(n_345), .Y(n_415) );
NOR2xp33_ASAP7_75t_L g421 ( .A(n_307), .B(n_422), .Y(n_421) );
INVx1_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
OR2x2_ASAP7_75t_L g403 ( .A(n_309), .B(n_404), .Y(n_403) );
INVx1_ASAP7_75t_SL g312 ( .A(n_313), .Y(n_312) );
NAND3xp33_ASAP7_75t_SL g314 ( .A(n_315), .B(n_331), .C(n_346), .Y(n_314) );
AOI221xp5_ASAP7_75t_L g315 ( .A1(n_316), .A2(n_317), .B1(n_322), .B2(n_324), .C(n_326), .Y(n_315) );
AND2x2_ASAP7_75t_L g322 ( .A(n_318), .B(n_323), .Y(n_322) );
INVx3_ASAP7_75t_SL g318 ( .A(n_319), .Y(n_318) );
AND2x4_ASAP7_75t_L g319 ( .A(n_320), .B(n_321), .Y(n_319) );
AND2x2_ASAP7_75t_L g332 ( .A(n_323), .B(n_333), .Y(n_332) );
HB1xp67_ASAP7_75t_L g404 ( .A(n_325), .Y(n_404) );
INVx1_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g360 ( .A(n_330), .B(n_344), .Y(n_360) );
NAND2xp5_ASAP7_75t_L g397 ( .A(n_333), .B(n_391), .Y(n_397) );
NOR2xp33_ASAP7_75t_L g393 ( .A(n_334), .B(n_394), .Y(n_393) );
INVx1_ASAP7_75t_SL g409 ( .A(n_337), .Y(n_409) );
AND2x2_ASAP7_75t_L g424 ( .A(n_337), .B(n_401), .Y(n_424) );
INVx1_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
NAND2xp5_ASAP7_75t_L g339 ( .A(n_340), .B(n_341), .Y(n_339) );
INVx1_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
AOI211xp5_ASAP7_75t_L g418 ( .A1(n_348), .A2(n_419), .B(n_425), .C(n_433), .Y(n_418) );
INVx1_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
OR2x2_ASAP7_75t_L g355 ( .A(n_356), .B(n_357), .Y(n_355) );
INVx1_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
AND2x2_ASAP7_75t_L g387 ( .A(n_358), .B(n_388), .Y(n_387) );
NAND2x1_ASAP7_75t_SL g429 ( .A(n_359), .B(n_430), .Y(n_429) );
CKINVDCx16_ASAP7_75t_R g399 ( .A(n_362), .Y(n_399) );
INVx1_ASAP7_75t_SL g363 ( .A(n_364), .Y(n_363) );
INVx1_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
INVx1_ASAP7_75t_L g394 ( .A(n_368), .Y(n_394) );
AND2x2_ASAP7_75t_L g398 ( .A(n_368), .B(n_384), .Y(n_398) );
NOR5xp2_ASAP7_75t_L g369 ( .A(n_370), .B(n_385), .C(n_402), .D(n_408), .E(n_411), .Y(n_369) );
OAI221xp5_ASAP7_75t_L g370 ( .A1(n_371), .A2(n_372), .B1(n_373), .B2(n_375), .C(n_377), .Y(n_370) );
INVx2_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_374), .B(n_432), .Y(n_431) );
INVxp67_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
NAND2xp5_ASAP7_75t_L g377 ( .A(n_378), .B(n_380), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
INVx1_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
NAND2xp5_ASAP7_75t_L g381 ( .A(n_382), .B(n_384), .Y(n_381) );
INVx1_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
AND2x2_ASAP7_75t_L g400 ( .A(n_384), .B(n_401), .Y(n_400) );
OAI221xp5_ASAP7_75t_SL g385 ( .A1(n_386), .A2(n_389), .B1(n_390), .B2(n_392), .C(n_395), .Y(n_385) );
INVx1_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
INVx1_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
AOI22xp33_ASAP7_75t_L g395 ( .A1(n_396), .A2(n_398), .B1(n_399), .B2(n_400), .Y(n_395) );
INVx1_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
INVx1_ASAP7_75t_L g438 ( .A(n_398), .Y(n_438) );
AOI211xp5_ASAP7_75t_SL g411 ( .A1(n_412), .A2(n_414), .B(n_416), .C(n_417), .Y(n_411) );
INVx1_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
INVx1_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
INVx1_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
INVx1_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
INVx1_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
INVxp67_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
NAND2xp5_ASAP7_75t_L g435 ( .A(n_436), .B(n_438), .Y(n_435) );
INVx1_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
CKINVDCx14_ASAP7_75t_R g440 ( .A(n_441), .Y(n_440) );
OAI22xp5_ASAP7_75t_SL g742 ( .A1(n_444), .A2(n_451), .B1(n_455), .B2(n_743), .Y(n_742) );
NAND3xp33_ASAP7_75t_L g448 ( .A(n_445), .B(n_449), .C(n_747), .Y(n_448) );
INVx1_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
INVx2_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
INVx1_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
INVx2_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
NAND2x1p5_ASAP7_75t_L g455 ( .A(n_456), .B(n_659), .Y(n_455) );
AND2x2_ASAP7_75t_SL g456 ( .A(n_457), .B(n_617), .Y(n_456) );
NOR4xp25_ASAP7_75t_L g457 ( .A(n_458), .B(n_557), .C(n_593), .D(n_607), .Y(n_457) );
OAI221xp5_ASAP7_75t_SL g458 ( .A1(n_459), .A2(n_505), .B1(n_535), .B2(n_544), .C(n_548), .Y(n_458) );
NAND2xp5_ASAP7_75t_SL g691 ( .A(n_459), .B(n_692), .Y(n_691) );
OR2x2_ASAP7_75t_L g459 ( .A(n_460), .B(n_485), .Y(n_459) );
INVx1_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
AND2x2_ASAP7_75t_L g461 ( .A(n_462), .B(n_473), .Y(n_461) );
AND2x2_ASAP7_75t_L g554 ( .A(n_462), .B(n_474), .Y(n_554) );
INVx3_ASAP7_75t_L g562 ( .A(n_462), .Y(n_562) );
AND2x2_ASAP7_75t_L g616 ( .A(n_462), .B(n_488), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g652 ( .A(n_462), .B(n_487), .Y(n_652) );
AND2x2_ASAP7_75t_L g710 ( .A(n_462), .B(n_572), .Y(n_710) );
AOI21xp5_ASAP7_75t_L g467 ( .A1(n_468), .A2(n_469), .B(n_471), .Y(n_467) );
INVx2_ASAP7_75t_L g481 ( .A(n_470), .Y(n_481) );
O2A1O1Ixp33_ASAP7_75t_L g494 ( .A1(n_471), .A2(n_481), .B(n_495), .C(n_496), .Y(n_494) );
AND2x2_ASAP7_75t_L g545 ( .A(n_473), .B(n_546), .Y(n_545) );
AND2x2_ASAP7_75t_L g559 ( .A(n_473), .B(n_488), .Y(n_559) );
INVx2_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
NAND2xp5_ASAP7_75t_L g574 ( .A(n_474), .B(n_488), .Y(n_574) );
AND2x2_ASAP7_75t_L g586 ( .A(n_474), .B(n_562), .Y(n_586) );
OR2x2_ASAP7_75t_L g588 ( .A(n_474), .B(n_546), .Y(n_588) );
AND2x2_ASAP7_75t_L g623 ( .A(n_474), .B(n_546), .Y(n_623) );
HB1xp67_ASAP7_75t_L g668 ( .A(n_474), .Y(n_668) );
INVx1_ASAP7_75t_L g676 ( .A(n_474), .Y(n_676) );
OAI21xp5_ASAP7_75t_L g475 ( .A1(n_476), .A2(n_479), .B(n_483), .Y(n_475) );
OAI221xp5_ASAP7_75t_L g593 ( .A1(n_485), .A2(n_594), .B1(n_598), .B2(n_602), .C(n_603), .Y(n_593) );
INVx1_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
AND2x2_ASAP7_75t_L g553 ( .A(n_486), .B(n_554), .Y(n_553) );
AND2x2_ASAP7_75t_L g486 ( .A(n_487), .B(n_498), .Y(n_486) );
INVx2_ASAP7_75t_L g552 ( .A(n_487), .Y(n_552) );
AND2x2_ASAP7_75t_L g605 ( .A(n_487), .B(n_606), .Y(n_605) );
AND2x2_ASAP7_75t_L g624 ( .A(n_487), .B(n_562), .Y(n_624) );
INVx2_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
AND2x2_ASAP7_75t_L g687 ( .A(n_488), .B(n_562), .Y(n_687) );
AND2x2_ASAP7_75t_L g609 ( .A(n_498), .B(n_554), .Y(n_609) );
OAI322xp33_ASAP7_75t_L g677 ( .A1(n_498), .A2(n_633), .A3(n_678), .B1(n_680), .B2(n_683), .C1(n_685), .C2(n_689), .Y(n_677) );
INVx3_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
NOR2x1_ASAP7_75t_L g560 ( .A(n_499), .B(n_561), .Y(n_560) );
INVx2_ASAP7_75t_L g573 ( .A(n_499), .Y(n_573) );
AND2x2_ASAP7_75t_L g682 ( .A(n_499), .B(n_562), .Y(n_682) );
AND2x2_ASAP7_75t_L g714 ( .A(n_499), .B(n_586), .Y(n_714) );
OR2x2_ASAP7_75t_L g717 ( .A(n_499), .B(n_718), .Y(n_717) );
AND2x4_ASAP7_75t_L g499 ( .A(n_500), .B(n_501), .Y(n_499) );
INVx1_ASAP7_75t_L g547 ( .A(n_500), .Y(n_547) );
INVx1_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
AND2x2_ASAP7_75t_L g506 ( .A(n_507), .B(n_518), .Y(n_506) );
INVx1_ASAP7_75t_L g730 ( .A(n_507), .Y(n_730) );
INVx1_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
OR2x2_ASAP7_75t_L g537 ( .A(n_508), .B(n_525), .Y(n_537) );
INVx2_ASAP7_75t_L g570 ( .A(n_508), .Y(n_570) );
INVx2_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
INVx2_ASAP7_75t_L g592 ( .A(n_509), .Y(n_592) );
HB1xp67_ASAP7_75t_L g600 ( .A(n_509), .Y(n_600) );
OR2x2_ASAP7_75t_L g724 ( .A(n_509), .B(n_725), .Y(n_724) );
AND2x2_ASAP7_75t_L g549 ( .A(n_518), .B(n_550), .Y(n_549) );
AND2x2_ASAP7_75t_L g589 ( .A(n_518), .B(n_590), .Y(n_589) );
AND2x2_ASAP7_75t_L g641 ( .A(n_518), .B(n_642), .Y(n_641) );
AND2x2_ASAP7_75t_L g518 ( .A(n_519), .B(n_525), .Y(n_518) );
AND2x2_ASAP7_75t_L g538 ( .A(n_519), .B(n_539), .Y(n_538) );
NOR2xp67_ASAP7_75t_L g596 ( .A(n_519), .B(n_597), .Y(n_596) );
AND2x2_ASAP7_75t_L g650 ( .A(n_519), .B(n_540), .Y(n_650) );
OR2x2_ASAP7_75t_L g658 ( .A(n_519), .B(n_592), .Y(n_658) );
INVx2_ASAP7_75t_L g519 ( .A(n_520), .Y(n_519) );
BUFx2_ASAP7_75t_L g567 ( .A(n_520), .Y(n_567) );
AND2x2_ASAP7_75t_L g577 ( .A(n_520), .B(n_578), .Y(n_577) );
AND2x2_ASAP7_75t_L g601 ( .A(n_520), .B(n_525), .Y(n_601) );
AND2x2_ASAP7_75t_L g665 ( .A(n_520), .B(n_540), .Y(n_665) );
NOR2xp33_ASAP7_75t_L g555 ( .A(n_525), .B(n_556), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g569 ( .A(n_525), .B(n_570), .Y(n_569) );
INVx2_ASAP7_75t_L g578 ( .A(n_525), .Y(n_578) );
INVx1_ASAP7_75t_L g583 ( .A(n_525), .Y(n_583) );
AND2x2_ASAP7_75t_L g595 ( .A(n_525), .B(n_596), .Y(n_595) );
HB1xp67_ASAP7_75t_L g673 ( .A(n_525), .Y(n_673) );
INVx1_ASAP7_75t_L g725 ( .A(n_525), .Y(n_725) );
AOI21xp5_ASAP7_75t_L g527 ( .A1(n_528), .A2(n_529), .B(n_530), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g535 ( .A(n_536), .B(n_538), .Y(n_535) );
AND2x2_ASAP7_75t_L g702 ( .A(n_536), .B(n_611), .Y(n_702) );
INVx2_ASAP7_75t_SL g536 ( .A(n_537), .Y(n_536) );
AND2x2_ASAP7_75t_L g629 ( .A(n_538), .B(n_630), .Y(n_629) );
AND2x2_ASAP7_75t_L g728 ( .A(n_538), .B(n_663), .Y(n_728) );
INVx1_ASAP7_75t_L g550 ( .A(n_539), .Y(n_550) );
AND2x2_ASAP7_75t_L g576 ( .A(n_539), .B(n_570), .Y(n_576) );
BUFx2_ASAP7_75t_L g635 ( .A(n_539), .Y(n_635) );
INVx1_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
BUFx6f_ASAP7_75t_L g556 ( .A(n_540), .Y(n_556) );
INVx1_ASAP7_75t_L g566 ( .A(n_540), .Y(n_566) );
NOR2xp67_ASAP7_75t_L g704 ( .A(n_544), .B(n_551), .Y(n_704) );
INVx2_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
AOI32xp33_ASAP7_75t_L g548 ( .A1(n_545), .A2(n_549), .A3(n_551), .B1(n_553), .B2(n_555), .Y(n_548) );
AND2x2_ASAP7_75t_L g688 ( .A(n_545), .B(n_561), .Y(n_688) );
AND2x2_ASAP7_75t_L g726 ( .A(n_545), .B(n_624), .Y(n_726) );
INVx1_ASAP7_75t_L g606 ( .A(n_546), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g720 ( .A(n_550), .B(n_612), .Y(n_720) );
NAND2xp5_ASAP7_75t_L g585 ( .A(n_551), .B(n_586), .Y(n_585) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_551), .B(n_554), .Y(n_602) );
NAND2xp5_ASAP7_75t_SL g705 ( .A(n_551), .B(n_623), .Y(n_705) );
OR2x2_ASAP7_75t_L g719 ( .A(n_551), .B(n_588), .Y(n_719) );
INVx3_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
AND2x2_ASAP7_75t_L g646 ( .A(n_552), .B(n_554), .Y(n_646) );
OR2x2_ASAP7_75t_L g655 ( .A(n_552), .B(n_642), .Y(n_655) );
NAND2xp5_ASAP7_75t_L g627 ( .A(n_554), .B(n_605), .Y(n_627) );
INVx2_ASAP7_75t_L g642 ( .A(n_556), .Y(n_642) );
OR2x2_ASAP7_75t_L g657 ( .A(n_556), .B(n_658), .Y(n_657) );
AND2x2_ASAP7_75t_L g672 ( .A(n_556), .B(n_673), .Y(n_672) );
A2O1A1Ixp33_ASAP7_75t_L g729 ( .A1(n_556), .A2(n_649), .B(n_730), .C(n_731), .Y(n_729) );
OAI321xp33_ASAP7_75t_L g557 ( .A1(n_558), .A2(n_563), .A3(n_568), .B1(n_571), .B2(n_575), .C(n_579), .Y(n_557) );
INVx1_ASAP7_75t_L g670 ( .A(n_558), .Y(n_670) );
NAND2x1p5_ASAP7_75t_L g558 ( .A(n_559), .B(n_560), .Y(n_558) );
AND2x2_ASAP7_75t_L g681 ( .A(n_559), .B(n_682), .Y(n_681) );
INVx1_ASAP7_75t_L g633 ( .A(n_561), .Y(n_633) );
INVx2_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g693 ( .A(n_562), .B(n_676), .Y(n_693) );
OAI221xp5_ASAP7_75t_L g700 ( .A1(n_563), .A2(n_701), .B1(n_703), .B2(n_705), .C(n_706), .Y(n_700) );
INVx1_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
AND2x2_ASAP7_75t_L g564 ( .A(n_565), .B(n_567), .Y(n_564) );
AND2x2_ASAP7_75t_L g638 ( .A(n_565), .B(n_612), .Y(n_638) );
HB1xp67_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g591 ( .A(n_566), .B(n_592), .Y(n_591) );
INVx2_ASAP7_75t_L g611 ( .A(n_567), .Y(n_611) );
A2O1A1Ixp33_ASAP7_75t_L g653 ( .A1(n_568), .A2(n_609), .B(n_654), .C(n_656), .Y(n_653) );
INVx1_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
AND2x2_ASAP7_75t_L g620 ( .A(n_570), .B(n_577), .Y(n_620) );
BUFx2_ASAP7_75t_L g630 ( .A(n_570), .Y(n_630) );
INVx1_ASAP7_75t_L g645 ( .A(n_570), .Y(n_645) );
INVx1_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
NOR2xp33_ASAP7_75t_L g572 ( .A(n_573), .B(n_574), .Y(n_572) );
OR2x2_ASAP7_75t_L g651 ( .A(n_573), .B(n_652), .Y(n_651) );
INVx1_ASAP7_75t_L g734 ( .A(n_573), .Y(n_734) );
INVx1_ASAP7_75t_L g727 ( .A(n_574), .Y(n_727) );
NAND2xp5_ASAP7_75t_L g575 ( .A(n_576), .B(n_577), .Y(n_575) );
AND2x2_ASAP7_75t_L g580 ( .A(n_576), .B(n_581), .Y(n_580) );
AND2x2_ASAP7_75t_L g684 ( .A(n_576), .B(n_601), .Y(n_684) );
INVx1_ASAP7_75t_L g613 ( .A(n_577), .Y(n_613) );
AOI22xp5_ASAP7_75t_L g579 ( .A1(n_580), .A2(n_584), .B1(n_587), .B2(n_589), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g696 ( .A(n_581), .B(n_697), .Y(n_696) );
INVxp67_ASAP7_75t_L g581 ( .A(n_582), .Y(n_581) );
AND2x4_ASAP7_75t_L g649 ( .A(n_582), .B(n_650), .Y(n_649) );
BUFx3_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
AND2x2_ASAP7_75t_SL g612 ( .A(n_583), .B(n_592), .Y(n_612) );
INVx1_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
AND2x2_ASAP7_75t_L g604 ( .A(n_586), .B(n_605), .Y(n_604) );
INVx1_ASAP7_75t_SL g587 ( .A(n_588), .Y(n_587) );
OR2x2_ASAP7_75t_L g614 ( .A(n_588), .B(n_615), .Y(n_614) );
INVx1_ASAP7_75t_SL g590 ( .A(n_591), .Y(n_590) );
OAI221xp5_ASAP7_75t_L g708 ( .A1(n_591), .A2(n_709), .B1(n_711), .B2(n_712), .C(n_713), .Y(n_708) );
INVx1_ASAP7_75t_L g597 ( .A(n_592), .Y(n_597) );
HB1xp67_ASAP7_75t_L g663 ( .A(n_592), .Y(n_663) );
INVx1_ASAP7_75t_SL g594 ( .A(n_595), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g713 ( .A(n_595), .B(n_714), .Y(n_713) );
OAI21xp5_ASAP7_75t_L g603 ( .A1(n_596), .A2(n_601), .B(n_604), .Y(n_603) );
INVx1_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
NAND2xp5_ASAP7_75t_L g706 ( .A(n_599), .B(n_609), .Y(n_706) );
AND2x2_ASAP7_75t_L g599 ( .A(n_600), .B(n_601), .Y(n_599) );
INVx1_ASAP7_75t_L g675 ( .A(n_600), .Y(n_675) );
AND2x2_ASAP7_75t_L g634 ( .A(n_601), .B(n_635), .Y(n_634) );
INVx2_ASAP7_75t_L g723 ( .A(n_601), .Y(n_723) );
INVx1_ASAP7_75t_L g639 ( .A(n_604), .Y(n_639) );
INVx1_ASAP7_75t_L g694 ( .A(n_605), .Y(n_694) );
OAI22xp5_ASAP7_75t_L g607 ( .A1(n_608), .A2(n_610), .B1(n_613), .B2(n_614), .Y(n_607) );
INVx1_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g610 ( .A(n_611), .B(n_612), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g644 ( .A(n_611), .B(n_645), .Y(n_644) );
INVx2_ASAP7_75t_L g679 ( .A(n_612), .Y(n_679) );
NAND2xp5_ASAP7_75t_SL g716 ( .A(n_612), .B(n_650), .Y(n_716) );
OR2x2_ASAP7_75t_L g689 ( .A(n_613), .B(n_642), .Y(n_689) );
INVx1_ASAP7_75t_L g628 ( .A(n_614), .Y(n_628) );
INVx1_ASAP7_75t_SL g615 ( .A(n_616), .Y(n_615) );
NAND2xp5_ASAP7_75t_L g666 ( .A(n_616), .B(n_667), .Y(n_666) );
NOR3xp33_ASAP7_75t_L g617 ( .A(n_618), .B(n_636), .C(n_647), .Y(n_617) );
OAI211xp5_ASAP7_75t_L g618 ( .A1(n_619), .A2(n_621), .B(n_625), .C(n_631), .Y(n_618) );
INVxp67_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
AOI221xp5_ASAP7_75t_L g690 ( .A1(n_620), .A2(n_691), .B1(n_695), .B2(n_698), .C(n_700), .Y(n_690) );
INVx1_ASAP7_75t_SL g621 ( .A(n_622), .Y(n_621) );
AND2x2_ASAP7_75t_L g622 ( .A(n_623), .B(n_624), .Y(n_622) );
AND2x2_ASAP7_75t_L g632 ( .A(n_623), .B(n_633), .Y(n_632) );
AND2x2_ASAP7_75t_L g686 ( .A(n_623), .B(n_687), .Y(n_686) );
OAI211xp5_ASAP7_75t_L g671 ( .A1(n_624), .A2(n_672), .B(n_674), .C(n_676), .Y(n_671) );
INVx2_ASAP7_75t_L g718 ( .A(n_624), .Y(n_718) );
OAI21xp5_ASAP7_75t_SL g625 ( .A1(n_626), .A2(n_628), .B(n_629), .Y(n_625) );
INVx1_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
AND2x2_ASAP7_75t_L g697 ( .A(n_630), .B(n_650), .Y(n_697) );
NAND2xp5_ASAP7_75t_L g631 ( .A(n_632), .B(n_634), .Y(n_631) );
OAI21xp5_ASAP7_75t_SL g636 ( .A1(n_637), .A2(n_639), .B(n_640), .Y(n_636) );
INVxp67_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
OAI21xp5_ASAP7_75t_SL g640 ( .A1(n_641), .A2(n_643), .B(n_646), .Y(n_640) );
NAND2xp5_ASAP7_75t_L g669 ( .A(n_641), .B(n_670), .Y(n_669) );
INVxp67_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g732 ( .A(n_646), .B(n_733), .Y(n_732) );
OAI21xp33_ASAP7_75t_L g647 ( .A1(n_648), .A2(n_651), .B(n_653), .Y(n_647) );
INVx1_ASAP7_75t_SL g648 ( .A(n_649), .Y(n_648) );
AND2x2_ASAP7_75t_L g674 ( .A(n_650), .B(n_675), .Y(n_674) );
INVx1_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
INVx1_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
AND4x1_ASAP7_75t_L g659 ( .A(n_660), .B(n_690), .C(n_707), .D(n_729), .Y(n_659) );
NOR2xp33_ASAP7_75t_L g660 ( .A(n_661), .B(n_677), .Y(n_660) );
OAI211xp5_ASAP7_75t_SL g661 ( .A1(n_662), .A2(n_666), .B(n_669), .C(n_671), .Y(n_661) );
OR2x2_ASAP7_75t_L g662 ( .A(n_663), .B(n_664), .Y(n_662) );
INVx1_ASAP7_75t_SL g664 ( .A(n_665), .Y(n_664) );
NAND2xp5_ASAP7_75t_L g678 ( .A(n_665), .B(n_679), .Y(n_678) );
INVx1_ASAP7_75t_L g667 ( .A(n_668), .Y(n_667) );
NOR2xp33_ASAP7_75t_L g698 ( .A(n_676), .B(n_699), .Y(n_698) );
INVx1_ASAP7_75t_L g680 ( .A(n_681), .Y(n_680) );
INVx1_ASAP7_75t_L g683 ( .A(n_684), .Y(n_683) );
NOR2xp33_ASAP7_75t_L g685 ( .A(n_686), .B(n_688), .Y(n_685) );
INVx1_ASAP7_75t_L g711 ( .A(n_686), .Y(n_711) );
INVx2_ASAP7_75t_SL g699 ( .A(n_687), .Y(n_699) );
OR2x2_ASAP7_75t_L g692 ( .A(n_693), .B(n_694), .Y(n_692) );
INVx1_ASAP7_75t_L g695 ( .A(n_696), .Y(n_695) );
INVx1_ASAP7_75t_L g712 ( .A(n_697), .Y(n_712) );
INVx1_ASAP7_75t_L g701 ( .A(n_702), .Y(n_701) );
INVx1_ASAP7_75t_L g703 ( .A(n_704), .Y(n_703) );
NOR2xp33_ASAP7_75t_SL g707 ( .A(n_708), .B(n_715), .Y(n_707) );
INVx1_ASAP7_75t_SL g709 ( .A(n_710), .Y(n_709) );
OAI221xp5_ASAP7_75t_SL g715 ( .A1(n_716), .A2(n_717), .B1(n_719), .B2(n_720), .C(n_721), .Y(n_715) );
AOI22xp5_ASAP7_75t_L g721 ( .A1(n_722), .A2(n_726), .B1(n_727), .B2(n_728), .Y(n_721) );
NAND2xp5_ASAP7_75t_SL g722 ( .A(n_723), .B(n_724), .Y(n_722) );
INVx1_ASAP7_75t_L g731 ( .A(n_732), .Y(n_731) );
INVx1_ASAP7_75t_L g733 ( .A(n_734), .Y(n_733) );
INVx2_ASAP7_75t_L g735 ( .A(n_736), .Y(n_735) );
INVx2_ASAP7_75t_L g743 ( .A(n_736), .Y(n_743) );
INVx1_ASAP7_75t_L g736 ( .A(n_737), .Y(n_736) );
CKINVDCx14_ASAP7_75t_R g741 ( .A(n_738), .Y(n_741) );
INVx2_ASAP7_75t_L g744 ( .A(n_745), .Y(n_744) );
INVx2_ASAP7_75t_L g745 ( .A(n_746), .Y(n_745) );
INVx1_ASAP7_75t_L g748 ( .A(n_749), .Y(n_748) );
INVx1_ASAP7_75t_L g749 ( .A(n_750), .Y(n_749) );
endmodule