module fake_jpeg_18392_n_131 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_131);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_131;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_57;
wire n_21;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

NOR2xp33_ASAP7_75t_L g13 ( 
.A(n_9),
.B(n_7),
.Y(n_13)
);

INVx2_ASAP7_75t_SL g14 ( 
.A(n_5),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_9),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_12),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_12),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_8),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_4),
.Y(n_27)
);

BUFx16f_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_13),
.B(n_8),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_29),
.B(n_30),
.Y(n_40)
);

INVx6_ASAP7_75t_SL g30 ( 
.A(n_28),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_23),
.Y(n_31)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_31),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_24),
.Y(n_32)
);

INVx1_ASAP7_75t_SL g42 ( 
.A(n_32),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_24),
.Y(n_33)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_33),
.Y(n_41)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_23),
.Y(n_34)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

AND2x2_ASAP7_75t_L g35 ( 
.A(n_28),
.B(n_0),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_35),
.B(n_14),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_24),
.Y(n_36)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_36),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_23),
.Y(n_38)
);

OR2x2_ASAP7_75t_L g39 ( 
.A(n_38),
.B(n_14),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_39),
.B(n_51),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_35),
.B(n_18),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g65 ( 
.A(n_45),
.B(n_46),
.Y(n_65)
);

A2O1A1Ixp33_ASAP7_75t_L g46 ( 
.A1(n_35),
.A2(n_13),
.B(n_20),
.C(n_15),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g47 ( 
.A1(n_38),
.A2(n_14),
.B1(n_27),
.B2(n_17),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_47),
.B(n_33),
.Y(n_54)
);

AOI21xp33_ASAP7_75t_L g63 ( 
.A1(n_48),
.A2(n_52),
.B(n_25),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_37),
.B(n_26),
.Y(n_51)
);

AND2x2_ASAP7_75t_L g52 ( 
.A(n_32),
.B(n_28),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_53),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_54),
.A2(n_41),
.B1(n_22),
.B2(n_17),
.Y(n_79)
);

CKINVDCx16_ASAP7_75t_R g55 ( 
.A(n_39),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_55),
.B(n_58),
.Y(n_72)
);

OA22x2_ASAP7_75t_L g56 ( 
.A1(n_39),
.A2(n_30),
.B1(n_34),
.B2(n_32),
.Y(n_56)
);

OA21x2_ASAP7_75t_L g85 ( 
.A1(n_56),
.A2(n_33),
.B(n_19),
.Y(n_85)
);

OR2x2_ASAP7_75t_L g57 ( 
.A(n_47),
.B(n_27),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_57),
.B(n_61),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_40),
.B(n_26),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_49),
.B(n_18),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_59),
.B(n_60),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_49),
.B(n_15),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_46),
.B(n_25),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_63),
.B(n_66),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_50),
.B(n_21),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_50),
.B(n_20),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_67),
.B(n_22),
.Y(n_81)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_52),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_68),
.B(n_70),
.Y(n_77)
);

BUFx2_ASAP7_75t_L g69 ( 
.A(n_42),
.Y(n_69)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_69),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_44),
.B(n_21),
.Y(n_70)
);

AND2x6_ASAP7_75t_L g73 ( 
.A(n_68),
.B(n_52),
.Y(n_73)
);

XOR2x2_ASAP7_75t_SL g89 ( 
.A(n_73),
.B(n_85),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_54),
.A2(n_53),
.B1(n_43),
.B2(n_44),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_74),
.A2(n_75),
.B1(n_85),
.B2(n_56),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_57),
.A2(n_43),
.B1(n_41),
.B2(n_42),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_79),
.A2(n_57),
.B1(n_61),
.B2(n_67),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_62),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_80),
.B(n_81),
.Y(n_93)
);

BUFx2_ASAP7_75t_L g82 ( 
.A(n_69),
.Y(n_82)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_82),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_62),
.Y(n_83)
);

AOI21xp5_ASAP7_75t_L g94 ( 
.A1(n_83),
.A2(n_56),
.B(n_69),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_73),
.A2(n_55),
.B1(n_85),
.B2(n_64),
.Y(n_86)
);

XNOR2xp5_ASAP7_75t_SL g100 ( 
.A(n_86),
.B(n_89),
.Y(n_100)
);

XOR2xp5_ASAP7_75t_L g87 ( 
.A(n_71),
.B(n_64),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_87),
.B(n_92),
.C(n_95),
.Y(n_103)
);

INVxp33_ASAP7_75t_L g90 ( 
.A(n_82),
.Y(n_90)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_90),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_91),
.A2(n_97),
.B1(n_77),
.B2(n_72),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_76),
.B(n_65),
.C(n_56),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_94),
.B(n_80),
.Y(n_106)
);

XOR2xp5_ASAP7_75t_L g95 ( 
.A(n_71),
.B(n_65),
.Y(n_95)
);

AOI22x1_ASAP7_75t_L g96 ( 
.A1(n_75),
.A2(n_56),
.B1(n_19),
.B2(n_16),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_96),
.A2(n_79),
.B1(n_84),
.B2(n_78),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_93),
.B(n_81),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_98),
.B(n_102),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_101),
.A2(n_106),
.B1(n_107),
.B2(n_0),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_87),
.B(n_95),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_92),
.B(n_74),
.C(n_83),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_104),
.B(n_89),
.C(n_96),
.Y(n_108)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_88),
.Y(n_105)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_105),
.Y(n_109)
);

XOR2xp5_ASAP7_75t_L g119 ( 
.A(n_108),
.B(n_111),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_103),
.B(n_84),
.C(n_16),
.Y(n_111)
);

AOI21xp5_ASAP7_75t_SL g112 ( 
.A1(n_100),
.A2(n_90),
.B(n_16),
.Y(n_112)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_112),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_101),
.B(n_10),
.Y(n_113)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_113),
.B(n_114),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_109),
.A2(n_104),
.B1(n_100),
.B2(n_103),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_116),
.A2(n_7),
.B1(n_5),
.B2(n_6),
.Y(n_124)
);

AOI21xp5_ASAP7_75t_L g118 ( 
.A1(n_110),
.A2(n_102),
.B(n_99),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_SL g122 ( 
.A1(n_118),
.A2(n_120),
.B(n_2),
.Y(n_122)
);

AOI21xp5_ASAP7_75t_L g120 ( 
.A1(n_110),
.A2(n_0),
.B(n_1),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_117),
.B(n_2),
.Y(n_121)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_121),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_122),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_115),
.B(n_2),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_L g127 ( 
.A1(n_123),
.A2(n_124),
.B(n_3),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_127),
.B(n_124),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_128),
.B(n_129),
.C(n_125),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_L g129 ( 
.A1(n_126),
.A2(n_122),
.B(n_116),
.Y(n_129)
);

AOI221xp5_ASAP7_75t_L g131 ( 
.A1(n_130),
.A2(n_3),
.B1(n_6),
.B2(n_119),
.C(n_129),
.Y(n_131)
);


endmodule