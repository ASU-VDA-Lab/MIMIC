module fake_jpeg_13962_n_107 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_8, n_15, n_7, n_107);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_8;
input n_15;
input n_7;

output n_107;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_106;
wire n_44;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_10),
.Y(n_32)
);

OR2x2_ASAP7_75t_SL g33 ( 
.A(n_30),
.B(n_1),
.Y(n_33)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

INVx11_ASAP7_75t_L g35 ( 
.A(n_11),
.Y(n_35)
);

BUFx16f_ASAP7_75t_L g36 ( 
.A(n_8),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_18),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_14),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_23),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_17),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_SL g41 ( 
.A(n_25),
.B(n_19),
.Y(n_41)
);

AND2x2_ASAP7_75t_SL g42 ( 
.A(n_9),
.B(n_31),
.Y(n_42)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_21),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_42),
.B(n_0),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_44),
.B(n_45),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_42),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_43),
.Y(n_46)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_46),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_42),
.B(n_0),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_47),
.B(n_49),
.Y(n_62)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_34),
.Y(n_48)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_48),
.B(n_50),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_36),
.B(n_1),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

OR2x2_ASAP7_75t_L g51 ( 
.A(n_33),
.B(n_2),
.Y(n_51)
);

OR2x2_ASAP7_75t_L g54 ( 
.A(n_51),
.B(n_33),
.Y(n_54)
);

CKINVDCx16_ASAP7_75t_R g53 ( 
.A(n_49),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_53),
.B(n_57),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_54),
.B(n_3),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_44),
.B(n_38),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_55),
.B(n_2),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_46),
.Y(n_56)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_56),
.Y(n_68)
);

OR2x2_ASAP7_75t_L g57 ( 
.A(n_51),
.B(n_41),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_46),
.Y(n_59)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_59),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g60 ( 
.A1(n_45),
.A2(n_35),
.B1(n_40),
.B2(n_39),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_60),
.A2(n_36),
.B1(n_4),
.B2(n_5),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_45),
.A2(n_37),
.B1(n_40),
.B2(n_35),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_61),
.A2(n_37),
.B1(n_36),
.B2(n_43),
.Y(n_65)
);

INVxp33_ASAP7_75t_L g64 ( 
.A(n_63),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_64),
.B(n_72),
.Y(n_78)
);

AOI21xp5_ASAP7_75t_L g86 ( 
.A1(n_65),
.A2(n_66),
.B(n_15),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g66 ( 
.A(n_58),
.B(n_32),
.C(n_37),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_67),
.B(n_62),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_69),
.B(n_70),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_63),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_58),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_71),
.B(n_73),
.Y(n_82)
);

CKINVDCx14_ASAP7_75t_R g72 ( 
.A(n_55),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_62),
.A2(n_52),
.B1(n_6),
.B2(n_7),
.Y(n_73)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_75),
.B(n_12),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_79),
.B(n_80),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_76),
.B(n_6),
.Y(n_80)
);

OAI21xp5_ASAP7_75t_L g81 ( 
.A1(n_64),
.A2(n_7),
.B(n_8),
.Y(n_81)
);

CKINVDCx16_ASAP7_75t_R g91 ( 
.A(n_81),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_SL g96 ( 
.A1(n_83),
.A2(n_84),
.B(n_86),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_66),
.B(n_13),
.Y(n_84)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_68),
.Y(n_85)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_85),
.Y(n_93)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_74),
.Y(n_87)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_87),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_75),
.B(n_20),
.Y(n_88)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_88),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_78),
.B(n_77),
.C(n_65),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_90),
.B(n_29),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_82),
.A2(n_22),
.B1(n_24),
.B2(n_26),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_SL g97 ( 
.A1(n_92),
.A2(n_80),
.B(n_78),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_97),
.B(n_98),
.Y(n_102)
);

CKINVDCx16_ASAP7_75t_R g98 ( 
.A(n_89),
.Y(n_98)
);

AOI21xp5_ASAP7_75t_L g99 ( 
.A1(n_90),
.A2(n_27),
.B(n_28),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_SL g101 ( 
.A(n_99),
.B(n_100),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_102),
.A2(n_91),
.B1(n_94),
.B2(n_92),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_103),
.B(n_96),
.Y(n_104)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_104),
.Y(n_105)
);

MAJx2_ASAP7_75t_L g106 ( 
.A(n_105),
.B(n_101),
.C(n_95),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_106),
.B(n_93),
.Y(n_107)
);


endmodule