module fake_netlist_6_4360_n_199 (n_16, n_1, n_9, n_8, n_18, n_10, n_21, n_24, n_6, n_15, n_27, n_3, n_14, n_0, n_4, n_22, n_26, n_13, n_11, n_28, n_17, n_23, n_12, n_20, n_7, n_30, n_2, n_5, n_19, n_29, n_31, n_25, n_199);

input n_16;
input n_1;
input n_9;
input n_8;
input n_18;
input n_10;
input n_21;
input n_24;
input n_6;
input n_15;
input n_27;
input n_3;
input n_14;
input n_0;
input n_4;
input n_22;
input n_26;
input n_13;
input n_11;
input n_28;
input n_17;
input n_23;
input n_12;
input n_20;
input n_7;
input n_30;
input n_2;
input n_5;
input n_19;
input n_29;
input n_31;
input n_25;

output n_199;

wire n_52;
wire n_91;
wire n_119;
wire n_46;
wire n_146;
wire n_163;
wire n_193;
wire n_147;
wire n_154;
wire n_191;
wire n_88;
wire n_98;
wire n_113;
wire n_63;
wire n_39;
wire n_73;
wire n_148;
wire n_138;
wire n_161;
wire n_68;
wire n_166;
wire n_184;
wire n_50;
wire n_158;
wire n_49;
wire n_83;
wire n_101;
wire n_167;
wire n_144;
wire n_174;
wire n_127;
wire n_125;
wire n_153;
wire n_168;
wire n_178;
wire n_77;
wire n_156;
wire n_149;
wire n_152;
wire n_106;
wire n_92;
wire n_145;
wire n_42;
wire n_133;
wire n_96;
wire n_90;
wire n_160;
wire n_105;
wire n_131;
wire n_54;
wire n_132;
wire n_188;
wire n_102;
wire n_186;
wire n_87;
wire n_195;
wire n_189;
wire n_32;
wire n_66;
wire n_99;
wire n_85;
wire n_78;
wire n_84;
wire n_130;
wire n_164;
wire n_100;
wire n_129;
wire n_121;
wire n_197;
wire n_137;
wire n_142;
wire n_143;
wire n_180;
wire n_47;
wire n_62;
wire n_155;
wire n_75;
wire n_109;
wire n_150;
wire n_122;
wire n_45;
wire n_34;
wire n_140;
wire n_70;
wire n_120;
wire n_37;
wire n_67;
wire n_33;
wire n_82;
wire n_38;
wire n_110;
wire n_151;
wire n_61;
wire n_112;
wire n_172;
wire n_81;
wire n_59;
wire n_181;
wire n_76;
wire n_36;
wire n_182;
wire n_124;
wire n_55;
wire n_126;
wire n_97;
wire n_94;
wire n_108;
wire n_58;
wire n_116;
wire n_64;
wire n_117;
wire n_118;
wire n_175;
wire n_48;
wire n_65;
wire n_40;
wire n_93;
wire n_80;
wire n_141;
wire n_135;
wire n_196;
wire n_165;
wire n_139;
wire n_41;
wire n_134;
wire n_177;
wire n_176;
wire n_114;
wire n_86;
wire n_198;
wire n_104;
wire n_95;
wire n_179;
wire n_107;
wire n_71;
wire n_74;
wire n_190;
wire n_123;
wire n_136;
wire n_72;
wire n_187;
wire n_89;
wire n_173;
wire n_103;
wire n_111;
wire n_60;
wire n_159;
wire n_157;
wire n_162;
wire n_170;
wire n_185;
wire n_35;
wire n_183;
wire n_115;
wire n_69;
wire n_128;
wire n_79;
wire n_43;
wire n_194;
wire n_171;
wire n_192;
wire n_57;
wire n_169;
wire n_53;
wire n_51;
wire n_44;
wire n_56;

CKINVDCx14_ASAP7_75t_R g32 ( 
.A(n_17),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_19),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_28),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_31),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_7),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_5),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_25),
.Y(n_39)
);

INVxp67_ASAP7_75t_SL g40 ( 
.A(n_15),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_27),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_5),
.Y(n_42)
);

CKINVDCx5p33_ASAP7_75t_R g43 ( 
.A(n_30),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_26),
.Y(n_44)
);

CKINVDCx5p33_ASAP7_75t_R g45 ( 
.A(n_22),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_2),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_21),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_16),
.Y(n_48)
);

CKINVDCx5p33_ASAP7_75t_R g49 ( 
.A(n_23),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_29),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_20),
.Y(n_51)
);

INVxp67_ASAP7_75t_SL g52 ( 
.A(n_7),
.Y(n_52)
);

INVxp33_ASAP7_75t_SL g53 ( 
.A(n_1),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_8),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_3),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_33),
.Y(n_56)
);

CKINVDCx5p33_ASAP7_75t_R g57 ( 
.A(n_43),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_33),
.Y(n_58)
);

CKINVDCx5p33_ASAP7_75t_R g59 ( 
.A(n_45),
.Y(n_59)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_46),
.Y(n_60)
);

CKINVDCx5p33_ASAP7_75t_R g61 ( 
.A(n_49),
.Y(n_61)
);

CKINVDCx5p33_ASAP7_75t_R g62 ( 
.A(n_32),
.Y(n_62)
);

AND2x4_ASAP7_75t_L g63 ( 
.A(n_35),
.B(n_24),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_R g64 ( 
.A(n_32),
.B(n_14),
.Y(n_64)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_33),
.Y(n_65)
);

CKINVDCx5p33_ASAP7_75t_R g66 ( 
.A(n_53),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_33),
.B(n_0),
.Y(n_67)
);

INVxp67_ASAP7_75t_L g68 ( 
.A(n_34),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_38),
.Y(n_69)
);

BUFx2_ASAP7_75t_L g70 ( 
.A(n_42),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_46),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_R g72 ( 
.A(n_54),
.B(n_18),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_46),
.Y(n_73)
);

CKINVDCx5p33_ASAP7_75t_R g74 ( 
.A(n_42),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_R g75 ( 
.A(n_36),
.B(n_12),
.Y(n_75)
);

CKINVDCx5p33_ASAP7_75t_R g76 ( 
.A(n_46),
.Y(n_76)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_60),
.Y(n_77)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_76),
.B(n_37),
.Y(n_78)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_60),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_71),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_66),
.A2(n_52),
.B1(n_55),
.B2(n_40),
.Y(n_81)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_71),
.Y(n_82)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_60),
.Y(n_83)
);

AND2x4_ASAP7_75t_L g84 ( 
.A(n_63),
.B(n_51),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_73),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_69),
.Y(n_86)
);

NAND3xp33_ASAP7_75t_SL g87 ( 
.A(n_74),
.B(n_50),
.C(n_48),
.Y(n_87)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_60),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_57),
.B(n_44),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_73),
.Y(n_90)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_67),
.Y(n_91)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_63),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_68),
.B(n_47),
.Y(n_93)
);

AND2x4_ASAP7_75t_L g94 ( 
.A(n_92),
.B(n_63),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_91),
.B(n_89),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_91),
.B(n_61),
.Y(n_96)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_83),
.Y(n_97)
);

BUFx3_ASAP7_75t_L g98 ( 
.A(n_83),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_84),
.B(n_63),
.Y(n_99)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_90),
.Y(n_100)
);

AND2x2_ASAP7_75t_SL g101 ( 
.A(n_84),
.B(n_39),
.Y(n_101)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_83),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_84),
.B(n_65),
.Y(n_103)
);

AO31x2_ASAP7_75t_L g104 ( 
.A1(n_81),
.A2(n_58),
.A3(n_56),
.B(n_65),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_78),
.B(n_59),
.Y(n_105)
);

BUFx2_ASAP7_75t_SL g106 ( 
.A(n_97),
.Y(n_106)
);

O2A1O1Ixp33_ASAP7_75t_L g107 ( 
.A1(n_95),
.A2(n_93),
.B(n_87),
.C(n_78),
.Y(n_107)
);

OAI21x1_ASAP7_75t_L g108 ( 
.A1(n_99),
.A2(n_58),
.B(n_56),
.Y(n_108)
);

AOI222xp33_ASAP7_75t_L g109 ( 
.A1(n_96),
.A2(n_70),
.B1(n_93),
.B2(n_41),
.C1(n_62),
.C2(n_86),
.Y(n_109)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_103),
.Y(n_110)
);

AND2x4_ASAP7_75t_L g111 ( 
.A(n_94),
.B(n_80),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_101),
.A2(n_85),
.B1(n_82),
.B2(n_80),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_L g113 ( 
.A1(n_103),
.A2(n_88),
.B(n_79),
.Y(n_113)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_111),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_111),
.Y(n_115)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_111),
.Y(n_116)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_111),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_110),
.B(n_101),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_110),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_106),
.B(n_101),
.Y(n_120)
);

BUFx2_ASAP7_75t_L g121 ( 
.A(n_114),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_116),
.Y(n_122)
);

INVx2_ASAP7_75t_SL g123 ( 
.A(n_117),
.Y(n_123)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_119),
.Y(n_124)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_115),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_124),
.Y(n_126)
);

NOR2xp67_ASAP7_75t_L g127 ( 
.A(n_123),
.B(n_105),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_L g128 ( 
.A1(n_121),
.A2(n_109),
.B1(n_122),
.B2(n_123),
.Y(n_128)
);

HB1xp67_ASAP7_75t_L g129 ( 
.A(n_121),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_124),
.B(n_118),
.Y(n_130)
);

HB1xp67_ASAP7_75t_L g131 ( 
.A(n_122),
.Y(n_131)
);

AND2x4_ASAP7_75t_SL g132 ( 
.A(n_122),
.B(n_86),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_125),
.B(n_70),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_125),
.Y(n_134)
);

AND2x2_ASAP7_75t_L g135 ( 
.A(n_122),
.B(n_118),
.Y(n_135)
);

AND2x2_ASAP7_75t_L g136 ( 
.A(n_122),
.B(n_104),
.Y(n_136)
);

AND2x2_ASAP7_75t_L g137 ( 
.A(n_135),
.B(n_104),
.Y(n_137)
);

OR2x2_ASAP7_75t_L g138 ( 
.A(n_135),
.B(n_120),
.Y(n_138)
);

HB1xp67_ASAP7_75t_L g139 ( 
.A(n_129),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_133),
.B(n_107),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_SL g141 ( 
.A1(n_132),
.A2(n_120),
.B(n_72),
.Y(n_141)
);

HB1xp67_ASAP7_75t_L g142 ( 
.A(n_131),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_126),
.Y(n_143)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_139),
.Y(n_144)
);

INVx1_ASAP7_75t_SL g145 ( 
.A(n_142),
.Y(n_145)
);

OAI22xp33_ASAP7_75t_L g146 ( 
.A1(n_140),
.A2(n_127),
.B1(n_130),
.B2(n_126),
.Y(n_146)
);

AND2x2_ASAP7_75t_L g147 ( 
.A(n_138),
.B(n_136),
.Y(n_147)
);

AND2x2_ASAP7_75t_L g148 ( 
.A(n_138),
.B(n_136),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_141),
.B(n_132),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_143),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_137),
.B(n_134),
.Y(n_151)
);

NAND3xp33_ASAP7_75t_L g152 ( 
.A(n_137),
.B(n_128),
.C(n_100),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_140),
.B(n_134),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_150),
.Y(n_154)
);

BUFx2_ASAP7_75t_L g155 ( 
.A(n_144),
.Y(n_155)
);

INVx1_ASAP7_75t_SL g156 ( 
.A(n_145),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_153),
.B(n_33),
.Y(n_157)
);

NOR2x1_ASAP7_75t_L g158 ( 
.A(n_146),
.B(n_85),
.Y(n_158)
);

AND2x4_ASAP7_75t_SL g159 ( 
.A(n_147),
.B(n_100),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_152),
.B(n_33),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_150),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_151),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_L g163 ( 
.A1(n_160),
.A2(n_149),
.B(n_56),
.Y(n_163)
);

OAI221xp5_ASAP7_75t_L g164 ( 
.A1(n_160),
.A2(n_82),
.B1(n_58),
.B2(n_112),
.C(n_148),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_162),
.B(n_148),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_156),
.B(n_147),
.Y(n_166)
);

OAI211xp5_ASAP7_75t_L g167 ( 
.A1(n_157),
.A2(n_75),
.B(n_64),
.C(n_3),
.Y(n_167)
);

OAI211xp5_ASAP7_75t_SL g168 ( 
.A1(n_158),
.A2(n_0),
.B(n_2),
.C(n_4),
.Y(n_168)
);

O2A1O1Ixp33_ASAP7_75t_L g169 ( 
.A1(n_155),
.A2(n_4),
.B(n_6),
.C(n_8),
.Y(n_169)
);

AOI221xp5_ASAP7_75t_L g170 ( 
.A1(n_154),
.A2(n_161),
.B1(n_159),
.B2(n_10),
.C(n_9),
.Y(n_170)
);

NAND4xp25_ASAP7_75t_SL g171 ( 
.A(n_159),
.B(n_6),
.C(n_9),
.D(n_10),
.Y(n_171)
);

OAI211xp5_ASAP7_75t_SL g172 ( 
.A1(n_169),
.A2(n_77),
.B(n_79),
.C(n_88),
.Y(n_172)
);

OAI21xp33_ASAP7_75t_L g173 ( 
.A1(n_171),
.A2(n_77),
.B(n_99),
.Y(n_173)
);

O2A1O1Ixp5_ASAP7_75t_L g174 ( 
.A1(n_163),
.A2(n_113),
.B(n_94),
.C(n_13),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_165),
.B(n_11),
.Y(n_175)
);

INVx1_ASAP7_75t_SL g176 ( 
.A(n_166),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_170),
.Y(n_177)
);

OAI221xp5_ASAP7_75t_L g178 ( 
.A1(n_168),
.A2(n_106),
.B1(n_104),
.B2(n_98),
.C(n_102),
.Y(n_178)
);

OAI32xp33_ASAP7_75t_L g179 ( 
.A1(n_164),
.A2(n_104),
.A3(n_97),
.B1(n_102),
.B2(n_98),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_176),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_177),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_175),
.Y(n_182)
);

NOR3xp33_ASAP7_75t_SL g183 ( 
.A(n_178),
.B(n_167),
.C(n_104),
.Y(n_183)
);

BUFx2_ASAP7_75t_SL g184 ( 
.A(n_173),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_172),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_174),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_181),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_186),
.B(n_179),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_186),
.A2(n_179),
.B1(n_94),
.B2(n_108),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_180),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_183),
.A2(n_184),
.B1(n_185),
.B2(n_182),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_187),
.B(n_104),
.Y(n_192)
);

HB1xp67_ASAP7_75t_L g193 ( 
.A(n_188),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_190),
.B(n_108),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_193),
.A2(n_191),
.B1(n_189),
.B2(n_94),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_194),
.B(n_98),
.Y(n_196)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_192),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_195),
.A2(n_97),
.B1(n_102),
.B2(n_197),
.Y(n_198)
);

NOR3xp33_ASAP7_75t_L g199 ( 
.A(n_198),
.B(n_196),
.C(n_97),
.Y(n_199)
);


endmodule