module fake_jpeg_9640_n_341 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_341);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_341;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_13),
.Y(n_16)
);

INVx3_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

BUFx12_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

INVx6_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

INVx11_ASAP7_75t_SL g20 ( 
.A(n_0),
.Y(n_20)
);

INVx6_ASAP7_75t_SL g21 ( 
.A(n_10),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

CKINVDCx16_ASAP7_75t_R g23 ( 
.A(n_14),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_3),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_15),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_9),
.Y(n_35)
);

INVx5_ASAP7_75t_L g36 ( 
.A(n_9),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_16),
.B(n_15),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_SL g49 ( 
.A(n_37),
.B(n_27),
.Y(n_49)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_36),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_38),
.B(n_41),
.Y(n_67)
);

INVx3_ASAP7_75t_SL g39 ( 
.A(n_32),
.Y(n_39)
);

BUFx2_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_34),
.Y(n_40)
);

INVx11_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_36),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_34),
.Y(n_42)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_42),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_35),
.Y(n_43)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_43),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_44),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_45),
.Y(n_53)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

BUFx2_ASAP7_75t_L g63 ( 
.A(n_46),
.Y(n_63)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_47),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_38),
.A2(n_19),
.B1(n_17),
.B2(n_32),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_48),
.A2(n_29),
.B1(n_22),
.B2(n_26),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_49),
.B(n_27),
.Y(n_68)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

INVx11_ASAP7_75t_L g88 ( 
.A(n_55),
.Y(n_88)
);

OR2x2_ASAP7_75t_L g56 ( 
.A(n_37),
.B(n_30),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_56),
.B(n_64),
.Y(n_79)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_58),
.Y(n_70)
);

MAJIxp5_ASAP7_75t_L g60 ( 
.A(n_40),
.B(n_32),
.C(n_35),
.Y(n_60)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_60),
.B(n_61),
.Y(n_74)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_46),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_62),
.B(n_65),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_40),
.B(n_29),
.Y(n_64)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_42),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_42),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_66),
.B(n_34),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_68),
.B(n_69),
.Y(n_106)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_64),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_55),
.A2(n_19),
.B1(n_17),
.B2(n_23),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_71),
.A2(n_76),
.B1(n_87),
.B2(n_93),
.Y(n_118)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_67),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_72),
.B(n_73),
.Y(n_126)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_67),
.Y(n_73)
);

BUFx2_ASAP7_75t_L g75 ( 
.A(n_54),
.Y(n_75)
);

INVx3_ASAP7_75t_SL g122 ( 
.A(n_75),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_60),
.A2(n_19),
.B1(n_17),
.B2(n_30),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_48),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_77),
.B(n_81),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g78 ( 
.A(n_51),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_78),
.Y(n_116)
);

HB1xp67_ASAP7_75t_L g80 ( 
.A(n_63),
.Y(n_80)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_80),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_63),
.Y(n_81)
);

AND2x4_ASAP7_75t_L g82 ( 
.A(n_55),
.B(n_21),
.Y(n_82)
);

OR2x4_ASAP7_75t_L g110 ( 
.A(n_82),
.B(n_85),
.Y(n_110)
);

INVx5_ASAP7_75t_L g83 ( 
.A(n_53),
.Y(n_83)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_83),
.Y(n_114)
);

BUFx12f_ASAP7_75t_L g84 ( 
.A(n_59),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_84),
.B(n_86),
.Y(n_135)
);

NOR2x1_ASAP7_75t_L g85 ( 
.A(n_56),
.B(n_21),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_49),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_58),
.A2(n_23),
.B1(n_47),
.B2(n_16),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_89),
.A2(n_24),
.B1(n_31),
.B2(n_28),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_63),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_90),
.B(n_99),
.Y(n_113)
);

HB1xp67_ASAP7_75t_L g92 ( 
.A(n_50),
.Y(n_92)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_92),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_L g93 ( 
.A1(n_61),
.A2(n_22),
.B1(n_26),
.B2(n_28),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_L g94 ( 
.A1(n_62),
.A2(n_31),
.B1(n_28),
.B2(n_24),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_94),
.A2(n_28),
.B1(n_24),
.B2(n_31),
.Y(n_127)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_52),
.Y(n_95)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_95),
.Y(n_107)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_96),
.Y(n_111)
);

BUFx8_ASAP7_75t_L g97 ( 
.A(n_51),
.Y(n_97)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_97),
.Y(n_134)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_54),
.Y(n_98)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_98),
.Y(n_128)
);

OR2x2_ASAP7_75t_L g99 ( 
.A(n_56),
.B(n_13),
.Y(n_99)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_52),
.Y(n_100)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_100),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_51),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_101),
.B(n_50),
.Y(n_119)
);

BUFx12f_ASAP7_75t_L g102 ( 
.A(n_59),
.Y(n_102)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_102),
.Y(n_129)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_65),
.Y(n_103)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_103),
.Y(n_130)
);

BUFx10_ASAP7_75t_L g104 ( 
.A(n_50),
.Y(n_104)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_104),
.Y(n_133)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_66),
.Y(n_105)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_105),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_77),
.A2(n_53),
.B1(n_57),
.B2(n_15),
.Y(n_109)
);

OAI22xp33_ASAP7_75t_SL g157 ( 
.A1(n_109),
.A2(n_112),
.B1(n_10),
.B2(n_12),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_82),
.A2(n_57),
.B1(n_14),
.B2(n_11),
.Y(n_112)
);

AOI21xp5_ASAP7_75t_L g115 ( 
.A1(n_74),
.A2(n_18),
.B(n_33),
.Y(n_115)
);

A2O1A1Ixp33_ASAP7_75t_L g137 ( 
.A1(n_115),
.A2(n_85),
.B(n_74),
.C(n_78),
.Y(n_137)
);

O2A1O1Ixp33_ASAP7_75t_L g117 ( 
.A1(n_82),
.A2(n_33),
.B(n_25),
.C(n_20),
.Y(n_117)
);

OAI32xp33_ASAP7_75t_L g143 ( 
.A1(n_117),
.A2(n_95),
.A3(n_100),
.B1(n_105),
.B2(n_97),
.Y(n_143)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_119),
.Y(n_138)
);

OAI22xp33_ASAP7_75t_L g123 ( 
.A1(n_74),
.A2(n_83),
.B1(n_82),
.B2(n_73),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_123),
.A2(n_25),
.B1(n_33),
.B2(n_84),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_69),
.B(n_45),
.C(n_44),
.Y(n_124)
);

AND2x2_ASAP7_75t_L g165 ( 
.A(n_124),
.B(n_104),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_125),
.A2(n_70),
.B1(n_88),
.B2(n_103),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_127),
.A2(n_90),
.B1(n_81),
.B2(n_98),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_136),
.A2(n_137),
.B1(n_150),
.B2(n_151),
.Y(n_171)
);

BUFx16f_ASAP7_75t_L g139 ( 
.A(n_122),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_139),
.B(n_149),
.Y(n_189)
);

MAJx2_ASAP7_75t_L g140 ( 
.A(n_110),
.B(n_79),
.C(n_72),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_140),
.B(n_11),
.C(n_8),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_113),
.B(n_86),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_141),
.B(n_156),
.Y(n_170)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_119),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_142),
.B(n_144),
.Y(n_186)
);

OAI22xp33_ASAP7_75t_SL g175 ( 
.A1(n_143),
.A2(n_155),
.B1(n_162),
.B2(n_166),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_134),
.B(n_101),
.Y(n_144)
);

AOI32xp33_ASAP7_75t_L g145 ( 
.A1(n_110),
.A2(n_70),
.A3(n_91),
.B1(n_43),
.B2(n_97),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_SL g190 ( 
.A1(n_145),
.A2(n_152),
.B(n_158),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_146),
.A2(n_160),
.B1(n_116),
.B2(n_120),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_126),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_147),
.B(n_148),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_134),
.B(n_84),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_131),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_123),
.A2(n_89),
.B1(n_88),
.B2(n_44),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_127),
.A2(n_45),
.B1(n_24),
.B2(n_31),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_135),
.Y(n_152)
);

INVxp67_ASAP7_75t_L g167 ( 
.A(n_153),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_108),
.B(n_102),
.Y(n_154)
);

CKINVDCx14_ASAP7_75t_R g178 ( 
.A(n_154),
.Y(n_178)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_122),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_113),
.B(n_99),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_157),
.A2(n_107),
.B1(n_111),
.B2(n_132),
.Y(n_177)
);

O2A1O1Ixp33_ASAP7_75t_L g158 ( 
.A1(n_118),
.A2(n_20),
.B(n_25),
.C(n_84),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_121),
.B(n_102),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_159),
.B(n_165),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_125),
.A2(n_104),
.B1(n_75),
.B2(n_102),
.Y(n_160)
);

NOR3xp33_ASAP7_75t_L g161 ( 
.A(n_115),
.B(n_104),
.C(n_18),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_161),
.Y(n_173)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_122),
.Y(n_162)
);

INVx8_ASAP7_75t_L g163 ( 
.A(n_114),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_SL g174 ( 
.A1(n_163),
.A2(n_128),
.B1(n_108),
.B2(n_120),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_SL g164 ( 
.A1(n_114),
.A2(n_12),
.B1(n_11),
.B2(n_10),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_164),
.A2(n_116),
.B1(n_128),
.B2(n_133),
.Y(n_181)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_124),
.Y(n_166)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_159),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_168),
.B(n_176),
.Y(n_206)
);

FAx1_ASAP7_75t_L g169 ( 
.A(n_150),
.B(n_117),
.CI(n_121),
.CON(n_169),
.SN(n_169)
);

OAI21xp5_ASAP7_75t_SL g219 ( 
.A1(n_169),
.A2(n_182),
.B(n_195),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_174),
.A2(n_177),
.B1(n_180),
.B2(n_7),
.Y(n_215)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_139),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_138),
.B(n_132),
.Y(n_179)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_179),
.Y(n_201)
);

OA22x2_ASAP7_75t_L g221 ( 
.A1(n_181),
.A2(n_191),
.B1(n_197),
.B2(n_3),
.Y(n_221)
);

AOI21xp5_ASAP7_75t_L g182 ( 
.A1(n_137),
.A2(n_129),
.B(n_130),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_139),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_183),
.B(n_184),
.Y(n_208)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_136),
.Y(n_184)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_163),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_185),
.B(n_187),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_141),
.Y(n_187)
);

OA22x2_ASAP7_75t_L g191 ( 
.A1(n_143),
.A2(n_130),
.B1(n_133),
.B2(n_18),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_166),
.A2(n_111),
.B1(n_106),
.B2(n_129),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_192),
.A2(n_199),
.B1(n_156),
.B2(n_151),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_193),
.B(n_140),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_153),
.B(n_18),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_194),
.B(n_152),
.C(n_142),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_SL g195 ( 
.A1(n_138),
.A2(n_18),
.B(n_1),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_149),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_196),
.B(n_200),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_146),
.Y(n_197)
);

NOR2x1_ASAP7_75t_L g198 ( 
.A(n_145),
.B(n_0),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_SL g224 ( 
.A(n_198),
.B(n_4),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_158),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_160),
.Y(n_200)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_179),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_202),
.B(n_209),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_204),
.B(n_212),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_205),
.B(n_207),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_196),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_200),
.A2(n_165),
.B1(n_147),
.B2(n_162),
.Y(n_210)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_210),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_L g211 ( 
.A1(n_182),
.A2(n_165),
.B(n_155),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_SL g248 ( 
.A1(n_211),
.A2(n_220),
.B(n_221),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_172),
.B(n_163),
.C(n_1),
.Y(n_212)
);

INVx1_ASAP7_75t_SL g213 ( 
.A(n_172),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_213),
.B(n_214),
.Y(n_247)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_186),
.Y(n_214)
);

CKINVDCx16_ASAP7_75t_R g251 ( 
.A(n_215),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_168),
.B(n_0),
.C(n_2),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_216),
.B(n_199),
.Y(n_255)
);

CKINVDCx16_ASAP7_75t_R g217 ( 
.A(n_189),
.Y(n_217)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_217),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_167),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_218),
.A2(n_225),
.B1(n_228),
.B2(n_230),
.Y(n_231)
);

HB1xp67_ASAP7_75t_SL g220 ( 
.A(n_198),
.Y(n_220)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_188),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_223),
.B(n_224),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_167),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_184),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_226)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_226),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_197),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_227)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_227),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_173),
.A2(n_175),
.B1(n_169),
.B2(n_171),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_SL g229 ( 
.A(n_187),
.B(n_192),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_229),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_185),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_211),
.B(n_190),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_233),
.B(n_243),
.Y(n_256)
);

AOI21xp5_ASAP7_75t_L g234 ( 
.A1(n_219),
.A2(n_190),
.B(n_195),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_234),
.B(n_210),
.Y(n_257)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_208),
.Y(n_236)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_236),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_222),
.A2(n_180),
.B1(n_177),
.B2(n_173),
.Y(n_237)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_237),
.Y(n_261)
);

OA21x2_ASAP7_75t_SL g241 ( 
.A1(n_213),
.A2(n_170),
.B(n_191),
.Y(n_241)
);

XOR2x2_ASAP7_75t_L g262 ( 
.A(n_241),
.B(n_191),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_219),
.B(n_170),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_L g245 ( 
.A1(n_222),
.A2(n_228),
.B1(n_208),
.B2(n_225),
.Y(n_245)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_245),
.Y(n_264)
);

INVxp67_ASAP7_75t_L g246 ( 
.A(n_203),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_246),
.B(n_178),
.Y(n_275)
);

BUFx3_ASAP7_75t_L g249 ( 
.A(n_223),
.Y(n_249)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_249),
.Y(n_266)
);

AND2x2_ASAP7_75t_L g253 ( 
.A(n_201),
.B(n_194),
.Y(n_253)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_253),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_204),
.B(n_193),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_254),
.B(n_206),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_255),
.B(n_169),
.Y(n_274)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_257),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_233),
.B(n_209),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_258),
.B(n_263),
.C(n_267),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_240),
.B(n_176),
.Y(n_259)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_259),
.Y(n_290)
);

AND3x1_ASAP7_75t_L g282 ( 
.A(n_262),
.B(n_241),
.C(n_248),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_240),
.B(n_183),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_265),
.B(n_270),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_235),
.B(n_232),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_243),
.B(n_206),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_269),
.B(n_271),
.C(n_272),
.Y(n_289)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_247),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_235),
.B(n_212),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_232),
.B(n_205),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_247),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_273),
.B(n_275),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_274),
.B(n_262),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_234),
.B(n_216),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_276),
.B(n_255),
.C(n_248),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_266),
.B(n_226),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_277),
.B(n_283),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_SL g295 ( 
.A(n_278),
.B(n_282),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_264),
.A2(n_251),
.B1(n_239),
.B2(n_238),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_280),
.A2(n_293),
.B1(n_294),
.B2(n_201),
.Y(n_302)
);

HB1xp67_ASAP7_75t_L g283 ( 
.A(n_260),
.Y(n_283)
);

XOR2x2_ASAP7_75t_L g286 ( 
.A(n_268),
.B(n_236),
.Y(n_286)
);

AOI21xp5_ASAP7_75t_L g296 ( 
.A1(n_286),
.A2(n_291),
.B(n_282),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_267),
.B(n_254),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_287),
.B(n_258),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_261),
.A2(n_239),
.B1(n_252),
.B2(n_244),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_288),
.B(n_218),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_272),
.B(n_246),
.Y(n_291)
);

XOR2xp5_ASAP7_75t_L g299 ( 
.A(n_292),
.B(n_256),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_276),
.A2(n_252),
.B1(n_244),
.B2(n_227),
.Y(n_293)
);

INVx3_ASAP7_75t_L g294 ( 
.A(n_269),
.Y(n_294)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_296),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_284),
.B(n_263),
.C(n_271),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_297),
.B(n_301),
.C(n_305),
.Y(n_314)
);

BUFx24_ASAP7_75t_SL g298 ( 
.A(n_290),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_298),
.B(n_307),
.Y(n_315)
);

XOR2xp5_ASAP7_75t_L g311 ( 
.A(n_299),
.B(n_303),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_284),
.B(n_289),
.C(n_292),
.Y(n_301)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_302),
.Y(n_317)
);

FAx1_ASAP7_75t_SL g304 ( 
.A(n_286),
.B(n_250),
.CI(n_253),
.CON(n_304),
.SN(n_304)
);

NAND2xp5_ASAP7_75t_SL g313 ( 
.A(n_304),
.B(n_306),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_289),
.B(n_256),
.C(n_202),
.Y(n_305)
);

OAI21xp5_ASAP7_75t_SL g306 ( 
.A1(n_281),
.A2(n_250),
.B(n_242),
.Y(n_306)
);

FAx1_ASAP7_75t_SL g307 ( 
.A(n_285),
.B(n_253),
.CI(n_249),
.CON(n_307),
.SN(n_307)
);

XNOR2xp5_ASAP7_75t_L g308 ( 
.A(n_279),
.B(n_231),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_308),
.B(n_288),
.C(n_221),
.Y(n_318)
);

XOR2xp5_ASAP7_75t_L g319 ( 
.A(n_309),
.B(n_221),
.Y(n_319)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_295),
.A2(n_294),
.B1(n_214),
.B2(n_242),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_310),
.B(n_312),
.Y(n_321)
);

INVx6_ASAP7_75t_L g312 ( 
.A(n_307),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_318),
.B(n_305),
.Y(n_326)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_319),
.Y(n_324)
);

NOR2xp67_ASAP7_75t_L g320 ( 
.A(n_304),
.B(n_221),
.Y(n_320)
);

XOR2x2_ASAP7_75t_L g325 ( 
.A(n_320),
.B(n_300),
.Y(n_325)
);

A2O1A1Ixp33_ASAP7_75t_SL g322 ( 
.A1(n_313),
.A2(n_309),
.B(n_295),
.C(n_191),
.Y(n_322)
);

OAI21x1_ASAP7_75t_L g332 ( 
.A1(n_322),
.A2(n_319),
.B(n_318),
.Y(n_332)
);

XNOR2xp5_ASAP7_75t_L g323 ( 
.A(n_314),
.B(n_301),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_323),
.B(n_327),
.Y(n_330)
);

OAI21x1_ASAP7_75t_L g333 ( 
.A1(n_325),
.A2(n_317),
.B(n_311),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_326),
.B(n_328),
.C(n_314),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_SL g327 ( 
.A(n_312),
.B(n_297),
.Y(n_327)
);

AOI21xp5_ASAP7_75t_L g328 ( 
.A1(n_316),
.A2(n_299),
.B(n_315),
.Y(n_328)
);

INVx6_ASAP7_75t_L g329 ( 
.A(n_321),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_329),
.B(n_331),
.Y(n_334)
);

OAI21xp5_ASAP7_75t_SL g335 ( 
.A1(n_332),
.A2(n_333),
.B(n_324),
.Y(n_335)
);

BUFx24_ASAP7_75t_SL g336 ( 
.A(n_335),
.Y(n_336)
);

AOI21xp5_ASAP7_75t_L g337 ( 
.A1(n_336),
.A2(n_334),
.B(n_330),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_337),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_SL g339 ( 
.A(n_338),
.B(n_329),
.Y(n_339)
);

AOI21xp5_ASAP7_75t_SL g340 ( 
.A1(n_339),
.A2(n_322),
.B(n_324),
.Y(n_340)
);

XOR2xp5_ASAP7_75t_L g341 ( 
.A(n_340),
.B(n_311),
.Y(n_341)
);


endmodule