module fake_ibex_1517_n_1202 (n_21, n_116, n_179, n_12, n_219, n_50, n_54, n_89, n_120, n_48, n_95, n_200, n_158, n_42, n_167, n_8, n_112, n_40, n_156, n_86, n_109, n_47, n_67, n_79, n_113, n_10, n_59, n_46, n_123, n_11, n_88, n_152, n_160, n_188, n_215, n_201, n_82, n_204, n_221, n_26, n_138, n_87, n_178, n_192, n_55, n_171, n_103, n_96, n_27, n_164, n_117, n_33, n_170, n_34, n_190, n_22, n_198, n_169, n_203, n_25, n_29, n_5, n_122, n_2, n_99, n_124, n_196, n_136, n_72, n_181, n_66, n_28, n_102, n_77, n_176, n_62, n_126, n_74, n_173, n_185, n_161, n_197, n_71, n_104, n_213, n_24, n_172, n_31, n_194, n_76, n_148, n_1, n_153, n_141, n_177, n_118, n_166, n_146, n_191, n_207, n_155, n_100, n_220, n_110, n_151, n_222, n_41, n_0, n_174, n_83, n_125, n_45, n_129, n_36, n_58, n_132, n_90, n_216, n_128, n_154, n_206, n_127, n_52, n_115, n_106, n_214, n_193, n_32, n_150, n_111, n_18, n_64, n_211, n_205, n_131, n_4, n_81, n_114, n_16, n_19, n_44, n_94, n_168, n_6, n_60, n_182, n_147, n_202, n_93, n_121, n_140, n_70, n_78, n_69, n_195, n_97, n_39, n_130, n_98, n_63, n_142, n_189, n_38, n_49, n_159, n_15, n_43, n_14, n_84, n_143, n_13, n_165, n_183, n_20, n_51, n_68, n_9, n_80, n_208, n_217, n_137, n_37, n_75, n_107, n_119, n_7, n_133, n_186, n_91, n_199, n_187, n_135, n_73, n_17, n_210, n_175, n_134, n_92, n_139, n_212, n_3, n_108, n_157, n_180, n_65, n_85, n_145, n_35, n_184, n_57, n_61, n_149, n_105, n_218, n_56, n_144, n_53, n_23, n_163, n_162, n_209, n_30, n_101, n_1202);

input n_21;
input n_116;
input n_179;
input n_12;
input n_219;
input n_50;
input n_54;
input n_89;
input n_120;
input n_48;
input n_95;
input n_200;
input n_158;
input n_42;
input n_167;
input n_8;
input n_112;
input n_40;
input n_156;
input n_86;
input n_109;
input n_47;
input n_67;
input n_79;
input n_113;
input n_10;
input n_59;
input n_46;
input n_123;
input n_11;
input n_88;
input n_152;
input n_160;
input n_188;
input n_215;
input n_201;
input n_82;
input n_204;
input n_221;
input n_26;
input n_138;
input n_87;
input n_178;
input n_192;
input n_55;
input n_171;
input n_103;
input n_96;
input n_27;
input n_164;
input n_117;
input n_33;
input n_170;
input n_34;
input n_190;
input n_22;
input n_198;
input n_169;
input n_203;
input n_25;
input n_29;
input n_5;
input n_122;
input n_2;
input n_99;
input n_124;
input n_196;
input n_136;
input n_72;
input n_181;
input n_66;
input n_28;
input n_102;
input n_77;
input n_176;
input n_62;
input n_126;
input n_74;
input n_173;
input n_185;
input n_161;
input n_197;
input n_71;
input n_104;
input n_213;
input n_24;
input n_172;
input n_31;
input n_194;
input n_76;
input n_148;
input n_1;
input n_153;
input n_141;
input n_177;
input n_118;
input n_166;
input n_146;
input n_191;
input n_207;
input n_155;
input n_100;
input n_220;
input n_110;
input n_151;
input n_222;
input n_41;
input n_0;
input n_174;
input n_83;
input n_125;
input n_45;
input n_129;
input n_36;
input n_58;
input n_132;
input n_90;
input n_216;
input n_128;
input n_154;
input n_206;
input n_127;
input n_52;
input n_115;
input n_106;
input n_214;
input n_193;
input n_32;
input n_150;
input n_111;
input n_18;
input n_64;
input n_211;
input n_205;
input n_131;
input n_4;
input n_81;
input n_114;
input n_16;
input n_19;
input n_44;
input n_94;
input n_168;
input n_6;
input n_60;
input n_182;
input n_147;
input n_202;
input n_93;
input n_121;
input n_140;
input n_70;
input n_78;
input n_69;
input n_195;
input n_97;
input n_39;
input n_130;
input n_98;
input n_63;
input n_142;
input n_189;
input n_38;
input n_49;
input n_159;
input n_15;
input n_43;
input n_14;
input n_84;
input n_143;
input n_13;
input n_165;
input n_183;
input n_20;
input n_51;
input n_68;
input n_9;
input n_80;
input n_208;
input n_217;
input n_137;
input n_37;
input n_75;
input n_107;
input n_119;
input n_7;
input n_133;
input n_186;
input n_91;
input n_199;
input n_187;
input n_135;
input n_73;
input n_17;
input n_210;
input n_175;
input n_134;
input n_92;
input n_139;
input n_212;
input n_3;
input n_108;
input n_157;
input n_180;
input n_65;
input n_85;
input n_145;
input n_35;
input n_184;
input n_57;
input n_61;
input n_149;
input n_105;
input n_218;
input n_56;
input n_144;
input n_53;
input n_23;
input n_163;
input n_162;
input n_209;
input n_30;
input n_101;

output n_1202;



endmodule