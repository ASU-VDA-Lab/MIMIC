module fake_jpeg_125_n_660 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_660);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_660;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_19;
wire n_182;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_657;
wire n_27;
wire n_365;
wire n_179;
wire n_620;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_479;
wire n_415;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_643;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_647;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_641;
wire n_48;
wire n_465;
wire n_638;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_637;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_646;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_658;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_639;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_645;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_92;
wire n_332;
wire n_640;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_653;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_642;
wire n_101;
wire n_226;
wire n_509;
wire n_644;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_656;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_649;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_615;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_648;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_650;
wire n_218;
wire n_63;
wire n_652;
wire n_599;
wire n_239;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_655;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_659;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_654;
wire n_445;
wire n_443;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_651;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_16),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_16),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_8),
.Y(n_22)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_18),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_5),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_18),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_8),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_12),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_3),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_6),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_0),
.Y(n_36)
);

BUFx10_ASAP7_75t_L g37 ( 
.A(n_1),
.Y(n_37)
);

CKINVDCx14_ASAP7_75t_R g38 ( 
.A(n_13),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_2),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_8),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_17),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_13),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_10),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_17),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_3),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_12),
.Y(n_46)
);

BUFx5_ASAP7_75t_L g47 ( 
.A(n_3),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_7),
.Y(n_48)
);

BUFx5_ASAP7_75t_L g49 ( 
.A(n_13),
.Y(n_49)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_15),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_14),
.Y(n_51)
);

BUFx5_ASAP7_75t_L g52 ( 
.A(n_18),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_6),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_15),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_1),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_8),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_16),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_16),
.Y(n_58)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_47),
.Y(n_59)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_59),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_19),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_60),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_19),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g175 ( 
.A(n_61),
.Y(n_175)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_19),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g176 ( 
.A(n_62),
.Y(n_176)
);

INVx11_ASAP7_75t_L g63 ( 
.A(n_56),
.Y(n_63)
);

INVx4_ASAP7_75t_L g136 ( 
.A(n_63),
.Y(n_136)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_32),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g131 ( 
.A(n_64),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_22),
.B(n_18),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_65),
.B(n_69),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_19),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g182 ( 
.A(n_66),
.Y(n_182)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_23),
.Y(n_67)
);

INVx3_ASAP7_75t_L g152 ( 
.A(n_67),
.Y(n_152)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_26),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g198 ( 
.A(n_68),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_22),
.B(n_24),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_26),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g200 ( 
.A(n_70),
.Y(n_200)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_28),
.Y(n_71)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_71),
.Y(n_145)
);

BUFx12_ASAP7_75t_L g72 ( 
.A(n_37),
.Y(n_72)
);

BUFx2_ASAP7_75t_R g188 ( 
.A(n_72),
.Y(n_188)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_28),
.Y(n_73)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_73),
.Y(n_146)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_23),
.Y(n_74)
);

INVx3_ASAP7_75t_L g183 ( 
.A(n_74),
.Y(n_183)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_27),
.Y(n_75)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_75),
.Y(n_142)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_47),
.Y(n_76)
);

INVx3_ASAP7_75t_L g185 ( 
.A(n_76),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_26),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g220 ( 
.A(n_77),
.Y(n_220)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_26),
.Y(n_78)
);

INVx6_ASAP7_75t_L g140 ( 
.A(n_78),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_42),
.Y(n_79)
);

INVx6_ASAP7_75t_L g143 ( 
.A(n_79),
.Y(n_143)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_27),
.Y(n_80)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_80),
.Y(n_156)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_30),
.Y(n_81)
);

BUFx3_ASAP7_75t_L g139 ( 
.A(n_81),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_42),
.Y(n_82)
);

INVx3_ASAP7_75t_SL g205 ( 
.A(n_82),
.Y(n_205)
);

INVx3_ASAP7_75t_SL g83 ( 
.A(n_32),
.Y(n_83)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_83),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_38),
.B(n_9),
.Y(n_84)
);

OR2x2_ASAP7_75t_L g216 ( 
.A(n_84),
.B(n_86),
.Y(n_216)
);

INVx6_ASAP7_75t_L g85 ( 
.A(n_42),
.Y(n_85)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_85),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_38),
.B(n_9),
.Y(n_86)
);

BUFx3_ASAP7_75t_L g87 ( 
.A(n_30),
.Y(n_87)
);

BUFx3_ASAP7_75t_L g147 ( 
.A(n_87),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_42),
.Y(n_88)
);

BUFx3_ASAP7_75t_L g180 ( 
.A(n_88),
.Y(n_180)
);

HB1xp67_ASAP7_75t_L g89 ( 
.A(n_23),
.Y(n_89)
);

CKINVDCx16_ASAP7_75t_R g133 ( 
.A(n_89),
.Y(n_133)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_27),
.Y(n_90)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_90),
.Y(n_169)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_50),
.Y(n_91)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_91),
.Y(n_171)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_47),
.Y(n_92)
);

INVx3_ASAP7_75t_L g191 ( 
.A(n_92),
.Y(n_191)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_48),
.Y(n_93)
);

BUFx3_ASAP7_75t_L g206 ( 
.A(n_93),
.Y(n_206)
);

INVx5_ASAP7_75t_L g94 ( 
.A(n_32),
.Y(n_94)
);

INVx4_ASAP7_75t_L g181 ( 
.A(n_94),
.Y(n_181)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_50),
.Y(n_95)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_95),
.Y(n_174)
);

INVx13_ASAP7_75t_L g96 ( 
.A(n_49),
.Y(n_96)
);

CKINVDCx14_ASAP7_75t_R g137 ( 
.A(n_96),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_50),
.B(n_9),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_97),
.B(n_110),
.Y(n_199)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_44),
.Y(n_98)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_98),
.Y(n_154)
);

BUFx3_ASAP7_75t_L g99 ( 
.A(n_30),
.Y(n_99)
);

INVx5_ASAP7_75t_L g130 ( 
.A(n_99),
.Y(n_130)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_58),
.Y(n_100)
);

INVx3_ASAP7_75t_L g208 ( 
.A(n_100),
.Y(n_208)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_58),
.Y(n_101)
);

INVx3_ASAP7_75t_L g212 ( 
.A(n_101),
.Y(n_212)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_48),
.Y(n_102)
);

INVx5_ASAP7_75t_L g161 ( 
.A(n_102),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_48),
.Y(n_103)
);

INVx5_ASAP7_75t_L g204 ( 
.A(n_103),
.Y(n_204)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_58),
.Y(n_104)
);

INVx3_ASAP7_75t_L g217 ( 
.A(n_104),
.Y(n_217)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_56),
.Y(n_105)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_105),
.Y(n_177)
);

INVx2_ASAP7_75t_SL g106 ( 
.A(n_56),
.Y(n_106)
);

INVx4_ASAP7_75t_L g150 ( 
.A(n_106),
.Y(n_150)
);

INVx2_ASAP7_75t_SL g107 ( 
.A(n_56),
.Y(n_107)
);

INVx4_ASAP7_75t_L g153 ( 
.A(n_107),
.Y(n_153)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_56),
.B(n_44),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_108),
.B(n_127),
.Y(n_149)
);

INVx2_ASAP7_75t_SL g109 ( 
.A(n_56),
.Y(n_109)
);

INVx4_ASAP7_75t_L g155 ( 
.A(n_109),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_51),
.B(n_9),
.Y(n_110)
);

INVx5_ASAP7_75t_L g111 ( 
.A(n_32),
.Y(n_111)
);

INVx4_ASAP7_75t_L g159 ( 
.A(n_111),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_57),
.B(n_17),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_112),
.B(n_17),
.Y(n_141)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_36),
.Y(n_113)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_113),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_48),
.Y(n_114)
);

INVx4_ASAP7_75t_L g172 ( 
.A(n_114),
.Y(n_172)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_36),
.Y(n_115)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_115),
.Y(n_195)
);

INVx4_ASAP7_75t_L g116 ( 
.A(n_49),
.Y(n_116)
);

INVx4_ASAP7_75t_L g173 ( 
.A(n_116),
.Y(n_173)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_36),
.Y(n_117)
);

INVx4_ASAP7_75t_L g178 ( 
.A(n_117),
.Y(n_178)
);

INVx4_ASAP7_75t_L g118 ( 
.A(n_49),
.Y(n_118)
);

INVx4_ASAP7_75t_L g186 ( 
.A(n_118),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_36),
.Y(n_119)
);

INVx4_ASAP7_75t_L g190 ( 
.A(n_119),
.Y(n_190)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_45),
.Y(n_120)
);

INVx4_ASAP7_75t_L g214 ( 
.A(n_120),
.Y(n_214)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_45),
.Y(n_121)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_121),
.Y(n_197)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_45),
.Y(n_122)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_122),
.Y(n_201)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_45),
.Y(n_123)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_123),
.Y(n_207)
);

INVx6_ASAP7_75t_L g124 ( 
.A(n_37),
.Y(n_124)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_124),
.Y(n_210)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_51),
.Y(n_125)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_125),
.Y(n_194)
);

INVx4_ASAP7_75t_L g126 ( 
.A(n_52),
.Y(n_126)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_126),
.Y(n_218)
);

OR2x2_ASAP7_75t_L g127 ( 
.A(n_20),
.B(n_7),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_20),
.Y(n_128)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_128),
.Y(n_222)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_20),
.Y(n_129)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_129),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_97),
.A2(n_25),
.B1(n_43),
.B2(n_41),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g246 ( 
.A1(n_134),
.A2(n_135),
.B1(n_164),
.B2(n_166),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_110),
.A2(n_25),
.B1(n_43),
.B2(n_41),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_141),
.B(n_162),
.Y(n_239)
);

AND2x4_ASAP7_75t_L g144 ( 
.A(n_108),
.B(n_128),
.Y(n_144)
);

INVx1_ASAP7_75t_SL g254 ( 
.A(n_144),
.Y(n_254)
);

NAND2xp33_ASAP7_75t_SL g151 ( 
.A(n_89),
.B(n_39),
.Y(n_151)
);

AND2x2_ASAP7_75t_L g268 ( 
.A(n_151),
.B(n_173),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_84),
.B(n_24),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_SL g227 ( 
.A(n_157),
.B(n_158),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_86),
.B(n_57),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_60),
.A2(n_40),
.B1(n_33),
.B2(n_35),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_160),
.A2(n_184),
.B1(n_187),
.B2(n_209),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_106),
.B(n_40),
.Y(n_162)
);

AOI21xp33_ASAP7_75t_SL g163 ( 
.A1(n_72),
.A2(n_35),
.B(n_33),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_163),
.B(n_37),
.C(n_52),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_61),
.A2(n_29),
.B1(n_54),
.B2(n_53),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_62),
.A2(n_29),
.B1(n_54),
.B2(n_53),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_L g168 ( 
.A1(n_119),
.A2(n_21),
.B1(n_54),
.B2(n_53),
.Y(n_168)
);

OA22x2_ASAP7_75t_L g289 ( 
.A1(n_168),
.A2(n_189),
.B1(n_211),
.B2(n_2),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_107),
.B(n_46),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_170),
.B(n_179),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_109),
.B(n_46),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_66),
.A2(n_102),
.B1(n_78),
.B2(n_79),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_70),
.A2(n_21),
.B1(n_31),
.B2(n_46),
.Y(n_187)
);

AOI22xp33_ASAP7_75t_L g189 ( 
.A1(n_120),
.A2(n_31),
.B1(n_21),
.B2(n_34),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_129),
.B(n_31),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_192),
.B(n_203),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_121),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_202),
.B(n_221),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_83),
.B(n_55),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_77),
.A2(n_55),
.B1(n_39),
.B2(n_34),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_82),
.A2(n_55),
.B1(n_39),
.B2(n_34),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_123),
.B(n_10),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_213),
.B(n_219),
.Y(n_283)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_93),
.Y(n_215)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_215),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_103),
.B(n_10),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_114),
.Y(n_221)
);

INVx5_ASAP7_75t_L g224 ( 
.A(n_139),
.Y(n_224)
);

INVx4_ASAP7_75t_L g336 ( 
.A(n_224),
.Y(n_336)
);

INVxp67_ASAP7_75t_SL g225 ( 
.A(n_137),
.Y(n_225)
);

INVxp67_ASAP7_75t_L g351 ( 
.A(n_225),
.Y(n_351)
);

INVx11_ASAP7_75t_L g228 ( 
.A(n_137),
.Y(n_228)
);

INVx4_ASAP7_75t_L g340 ( 
.A(n_228),
.Y(n_340)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_167),
.Y(n_229)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_229),
.Y(n_309)
);

NAND3xp33_ASAP7_75t_L g310 ( 
.A(n_230),
.B(n_232),
.C(n_271),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_138),
.B(n_7),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_SL g338 ( 
.A(n_231),
.B(n_242),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_161),
.Y(n_232)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_197),
.Y(n_233)
);

INVx2_ASAP7_75t_L g324 ( 
.A(n_233),
.Y(n_324)
);

AOI22xp33_ASAP7_75t_SL g234 ( 
.A1(n_144),
.A2(n_37),
.B1(n_52),
.B2(n_11),
.Y(n_234)
);

INVxp67_ASAP7_75t_L g353 ( 
.A(n_234),
.Y(n_353)
);

INVx2_ASAP7_75t_SL g235 ( 
.A(n_150),
.Y(n_235)
);

INVx2_ASAP7_75t_SL g343 ( 
.A(n_235),
.Y(n_343)
);

INVx11_ASAP7_75t_L g236 ( 
.A(n_188),
.Y(n_236)
);

INVx11_ASAP7_75t_L g323 ( 
.A(n_236),
.Y(n_323)
);

BUFx2_ASAP7_75t_L g237 ( 
.A(n_150),
.Y(n_237)
);

INVx2_ASAP7_75t_L g332 ( 
.A(n_237),
.Y(n_332)
);

INVx3_ASAP7_75t_L g238 ( 
.A(n_153),
.Y(n_238)
);

BUFx4f_ASAP7_75t_SL g308 ( 
.A(n_238),
.Y(n_308)
);

AOI22xp33_ASAP7_75t_L g240 ( 
.A1(n_196),
.A2(n_37),
.B1(n_6),
.B2(n_11),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_L g316 ( 
.A1(n_240),
.A2(n_267),
.B1(n_273),
.B2(n_143),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_145),
.B(n_6),
.Y(n_242)
);

BUFx6f_ASAP7_75t_L g243 ( 
.A(n_148),
.Y(n_243)
);

INVx5_ASAP7_75t_L g314 ( 
.A(n_243),
.Y(n_314)
);

AOI22xp33_ASAP7_75t_SL g245 ( 
.A1(n_144),
.A2(n_37),
.B1(n_11),
.B2(n_12),
.Y(n_245)
);

AOI22xp33_ASAP7_75t_SL g339 ( 
.A1(n_245),
.A2(n_255),
.B1(n_289),
.B2(n_292),
.Y(n_339)
);

BUFx3_ASAP7_75t_L g247 ( 
.A(n_130),
.Y(n_247)
);

INVx3_ASAP7_75t_L g315 ( 
.A(n_247),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_146),
.B(n_4),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_248),
.B(n_259),
.Y(n_302)
);

INVx3_ASAP7_75t_L g249 ( 
.A(n_153),
.Y(n_249)
);

INVx3_ASAP7_75t_L g348 ( 
.A(n_249),
.Y(n_348)
);

INVx3_ASAP7_75t_L g250 ( 
.A(n_155),
.Y(n_250)
);

INVx2_ASAP7_75t_L g335 ( 
.A(n_250),
.Y(n_335)
);

INVx4_ASAP7_75t_L g251 ( 
.A(n_155),
.Y(n_251)
);

INVx2_ASAP7_75t_L g349 ( 
.A(n_251),
.Y(n_349)
);

INVx3_ASAP7_75t_L g252 ( 
.A(n_165),
.Y(n_252)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_252),
.Y(n_305)
);

AND2x2_ASAP7_75t_SL g253 ( 
.A(n_199),
.B(n_0),
.Y(n_253)
);

AND2x2_ASAP7_75t_L g329 ( 
.A(n_253),
.B(n_264),
.Y(n_329)
);

AOI22xp33_ASAP7_75t_SL g255 ( 
.A1(n_149),
.A2(n_4),
.B1(n_14),
.B2(n_13),
.Y(n_255)
);

INVx1_ASAP7_75t_SL g256 ( 
.A(n_173),
.Y(n_256)
);

INVx5_ASAP7_75t_SL g345 ( 
.A(n_256),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_216),
.B(n_0),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_SL g311 ( 
.A(n_257),
.B(n_279),
.Y(n_311)
);

INVx3_ASAP7_75t_L g258 ( 
.A(n_159),
.Y(n_258)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_258),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_154),
.B(n_194),
.Y(n_259)
);

CKINVDCx16_ASAP7_75t_R g260 ( 
.A(n_216),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_260),
.B(n_262),
.Y(n_307)
);

INVx5_ASAP7_75t_L g261 ( 
.A(n_139),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_261),
.Y(n_313)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_222),
.Y(n_262)
);

INVx11_ASAP7_75t_L g263 ( 
.A(n_159),
.Y(n_263)
);

INVx11_ASAP7_75t_L g331 ( 
.A(n_263),
.Y(n_331)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_207),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_171),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_265),
.B(n_269),
.Y(n_318)
);

HB1xp67_ASAP7_75t_L g266 ( 
.A(n_208),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_266),
.Y(n_325)
);

AOI22xp33_ASAP7_75t_L g267 ( 
.A1(n_168),
.A2(n_4),
.B1(n_14),
.B2(n_5),
.Y(n_267)
);

AND2x2_ASAP7_75t_L g356 ( 
.A(n_268),
.B(n_270),
.Y(n_356)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_174),
.Y(n_269)
);

INVx5_ASAP7_75t_L g270 ( 
.A(n_147),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_204),
.Y(n_271)
);

INVxp67_ASAP7_75t_L g272 ( 
.A(n_218),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_272),
.B(n_275),
.Y(n_333)
);

AOI22xp33_ASAP7_75t_L g273 ( 
.A1(n_189),
.A2(n_5),
.B1(n_14),
.B2(n_15),
.Y(n_273)
);

AND2x2_ASAP7_75t_L g274 ( 
.A(n_142),
.B(n_156),
.Y(n_274)
);

AND2x2_ASAP7_75t_L g360 ( 
.A(n_274),
.B(n_276),
.Y(n_360)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_140),
.Y(n_275)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_193),
.Y(n_276)
);

HB1xp67_ASAP7_75t_L g277 ( 
.A(n_212),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g352 ( 
.A(n_277),
.B(n_280),
.Y(n_352)
);

AO22x1_ASAP7_75t_SL g278 ( 
.A1(n_169),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_278),
.B(n_288),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_177),
.B(n_201),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_140),
.Y(n_280)
);

INVx3_ASAP7_75t_L g281 ( 
.A(n_178),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_281),
.B(n_284),
.Y(n_354)
);

O2A1O1Ixp33_ASAP7_75t_L g282 ( 
.A1(n_131),
.A2(n_0),
.B(n_1),
.C(n_2),
.Y(n_282)
);

OAI21xp5_ASAP7_75t_L g322 ( 
.A1(n_282),
.A2(n_286),
.B(n_136),
.Y(n_322)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_195),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_132),
.B(n_15),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g359 ( 
.A(n_285),
.B(n_291),
.Y(n_359)
);

AOI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_147),
.A2(n_2),
.B1(n_3),
.B2(n_217),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_133),
.B(n_183),
.Y(n_288)
);

BUFx6f_ASAP7_75t_L g290 ( 
.A(n_148),
.Y(n_290)
);

INVx8_ASAP7_75t_L g355 ( 
.A(n_290),
.Y(n_355)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_205),
.Y(n_291)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_205),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_185),
.B(n_3),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_SL g330 ( 
.A(n_293),
.B(n_296),
.Y(n_330)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_178),
.Y(n_294)
);

AOI22xp33_ASAP7_75t_SL g358 ( 
.A1(n_294),
.A2(n_299),
.B1(n_300),
.B2(n_301),
.Y(n_358)
);

BUFx2_ASAP7_75t_L g295 ( 
.A(n_131),
.Y(n_295)
);

INVx8_ASAP7_75t_L g357 ( 
.A(n_295),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_152),
.B(n_191),
.Y(n_296)
);

CKINVDCx16_ASAP7_75t_R g297 ( 
.A(n_186),
.Y(n_297)
);

CKINVDCx12_ASAP7_75t_R g347 ( 
.A(n_297),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_186),
.B(n_181),
.C(n_210),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g321 ( 
.A(n_298),
.B(n_200),
.Y(n_321)
);

INVx3_ASAP7_75t_L g299 ( 
.A(n_172),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_172),
.Y(n_300)
);

INVx4_ASAP7_75t_L g301 ( 
.A(n_136),
.Y(n_301)
);

AOI22xp33_ASAP7_75t_L g303 ( 
.A1(n_246),
.A2(n_190),
.B1(n_214),
.B2(n_198),
.Y(n_303)
);

OAI22x1_ASAP7_75t_L g380 ( 
.A1(n_303),
.A2(n_320),
.B1(n_342),
.B2(n_350),
.Y(n_380)
);

OAI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_287),
.A2(n_198),
.B1(n_143),
.B2(n_214),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g393 ( 
.A1(n_304),
.A2(n_334),
.B1(n_337),
.B2(n_346),
.Y(n_393)
);

AND2x2_ASAP7_75t_L g368 ( 
.A(n_316),
.B(n_321),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_244),
.B(n_190),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_SL g366 ( 
.A(n_317),
.B(n_341),
.Y(n_366)
);

AOI22xp5_ASAP7_75t_L g319 ( 
.A1(n_287),
.A2(n_182),
.B1(n_175),
.B2(n_176),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_L g374 ( 
.A1(n_319),
.A2(n_326),
.B1(n_327),
.B2(n_228),
.Y(n_374)
);

AOI22xp33_ASAP7_75t_L g320 ( 
.A1(n_254),
.A2(n_182),
.B1(n_175),
.B2(n_176),
.Y(n_320)
);

CKINVDCx16_ASAP7_75t_R g391 ( 
.A(n_322),
.Y(n_391)
);

AOI22xp5_ASAP7_75t_L g326 ( 
.A1(n_254),
.A2(n_200),
.B1(n_220),
.B2(n_206),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_L g327 ( 
.A1(n_268),
.A2(n_220),
.B1(n_206),
.B2(n_180),
.Y(n_327)
);

OR2x4_ASAP7_75t_L g328 ( 
.A(n_268),
.B(n_180),
.Y(n_328)
);

CKINVDCx14_ASAP7_75t_R g378 ( 
.A(n_328),
.Y(n_378)
);

OAI22xp5_ASAP7_75t_L g334 ( 
.A1(n_230),
.A2(n_283),
.B1(n_289),
.B2(n_257),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_L g337 ( 
.A1(n_289),
.A2(n_241),
.B1(n_286),
.B2(n_288),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_253),
.B(n_279),
.Y(n_341)
);

AOI22xp33_ASAP7_75t_L g342 ( 
.A1(n_289),
.A2(n_223),
.B1(n_226),
.B2(n_299),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_253),
.B(n_278),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_SL g379 ( 
.A(n_344),
.B(n_282),
.Y(n_379)
);

OAI22xp5_ASAP7_75t_L g346 ( 
.A1(n_239),
.A2(n_298),
.B1(n_227),
.B2(n_278),
.Y(n_346)
);

AOI22xp33_ASAP7_75t_L g350 ( 
.A1(n_291),
.A2(n_292),
.B1(n_229),
.B2(n_294),
.Y(n_350)
);

AOI22xp33_ASAP7_75t_SL g361 ( 
.A1(n_236),
.A2(n_258),
.B1(n_247),
.B2(n_281),
.Y(n_361)
);

INVxp67_ASAP7_75t_L g364 ( 
.A(n_361),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g362 ( 
.A(n_307),
.B(n_302),
.Y(n_362)
);

INVxp67_ASAP7_75t_L g416 ( 
.A(n_362),
.Y(n_416)
);

MAJx2_ASAP7_75t_L g363 ( 
.A(n_311),
.B(n_274),
.C(n_284),
.Y(n_363)
);

XOR2xp5_ASAP7_75t_L g420 ( 
.A(n_363),
.B(n_395),
.Y(n_420)
);

INVx2_ASAP7_75t_L g365 ( 
.A(n_343),
.Y(n_365)
);

INVx2_ASAP7_75t_SL g445 ( 
.A(n_365),
.Y(n_445)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_343),
.Y(n_367)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_367),
.Y(n_411)
);

INVx1_ASAP7_75t_SL g369 ( 
.A(n_356),
.Y(n_369)
);

BUFx3_ASAP7_75t_L g429 ( 
.A(n_369),
.Y(n_429)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_343),
.Y(n_370)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_370),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_L g371 ( 
.A(n_346),
.B(n_272),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_SL g447 ( 
.A(n_371),
.B(n_375),
.Y(n_447)
);

INVxp67_ASAP7_75t_L g372 ( 
.A(n_354),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_L g415 ( 
.A(n_372),
.B(n_385),
.Y(n_415)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_360),
.Y(n_373)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_373),
.Y(n_414)
);

AOI22xp33_ASAP7_75t_L g425 ( 
.A1(n_374),
.A2(n_309),
.B1(n_331),
.B2(n_324),
.Y(n_425)
);

NOR2xp33_ASAP7_75t_L g375 ( 
.A(n_338),
.B(n_274),
.Y(n_375)
);

BUFx2_ASAP7_75t_L g376 ( 
.A(n_355),
.Y(n_376)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_376),
.Y(n_418)
);

OAI21xp5_ASAP7_75t_SL g377 ( 
.A1(n_328),
.A2(n_235),
.B(n_238),
.Y(n_377)
);

OAI21xp5_ASAP7_75t_L g413 ( 
.A1(n_377),
.A2(n_378),
.B(n_369),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_SL g440 ( 
.A(n_379),
.B(n_348),
.Y(n_440)
);

INVx4_ASAP7_75t_L g381 ( 
.A(n_357),
.Y(n_381)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_381),
.Y(n_419)
);

AOI22xp5_ASAP7_75t_SL g382 ( 
.A1(n_337),
.A2(n_224),
.B1(n_270),
.B2(n_261),
.Y(n_382)
);

AND2x2_ASAP7_75t_L g433 ( 
.A(n_382),
.B(n_384),
.Y(n_433)
);

OAI22xp5_ASAP7_75t_SL g383 ( 
.A1(n_312),
.A2(n_233),
.B1(n_264),
.B2(n_243),
.Y(n_383)
);

AOI22xp5_ASAP7_75t_L g434 ( 
.A1(n_383),
.A2(n_386),
.B1(n_390),
.B2(n_392),
.Y(n_434)
);

AND2x2_ASAP7_75t_L g384 ( 
.A(n_356),
.B(n_252),
.Y(n_384)
);

INVx2_ASAP7_75t_L g385 ( 
.A(n_308),
.Y(n_385)
);

OAI22xp5_ASAP7_75t_SL g386 ( 
.A1(n_312),
.A2(n_290),
.B1(n_276),
.B2(n_250),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_360),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_L g421 ( 
.A(n_387),
.B(n_388),
.Y(n_421)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_308),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_SL g389 ( 
.A(n_311),
.B(n_249),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_389),
.B(n_398),
.Y(n_409)
);

OAI22xp5_ASAP7_75t_SL g390 ( 
.A1(n_319),
.A2(n_295),
.B1(n_251),
.B2(n_256),
.Y(n_390)
);

OAI22xp5_ASAP7_75t_SL g392 ( 
.A1(n_344),
.A2(n_237),
.B1(n_301),
.B2(n_263),
.Y(n_392)
);

OAI22xp5_ASAP7_75t_SL g394 ( 
.A1(n_339),
.A2(n_317),
.B1(n_334),
.B2(n_330),
.Y(n_394)
);

AOI22xp5_ASAP7_75t_SL g427 ( 
.A1(n_394),
.A2(n_397),
.B1(n_403),
.B2(n_345),
.Y(n_427)
);

MAJx2_ASAP7_75t_L g395 ( 
.A(n_341),
.B(n_330),
.C(n_329),
.Y(n_395)
);

AOI22xp33_ASAP7_75t_SL g396 ( 
.A1(n_353),
.A2(n_356),
.B1(n_304),
.B2(n_323),
.Y(n_396)
);

AOI22xp33_ASAP7_75t_SL g410 ( 
.A1(n_396),
.A2(n_351),
.B1(n_340),
.B2(n_315),
.Y(n_410)
);

OAI22xp5_ASAP7_75t_SL g397 ( 
.A1(n_322),
.A2(n_329),
.B1(n_310),
.B2(n_353),
.Y(n_397)
);

OAI32xp33_ASAP7_75t_L g398 ( 
.A1(n_329),
.A2(n_359),
.A3(n_338),
.B1(n_360),
.B2(n_352),
.Y(n_398)
);

BUFx6f_ASAP7_75t_L g399 ( 
.A(n_314),
.Y(n_399)
);

CKINVDCx20_ASAP7_75t_R g424 ( 
.A(n_399),
.Y(n_424)
);

MAJIxp5_ASAP7_75t_L g400 ( 
.A(n_321),
.B(n_318),
.C(n_333),
.Y(n_400)
);

XNOR2xp5_ASAP7_75t_L g435 ( 
.A(n_400),
.B(n_335),
.Y(n_435)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_324),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_L g426 ( 
.A(n_401),
.B(n_402),
.Y(n_426)
);

INVxp67_ASAP7_75t_L g402 ( 
.A(n_315),
.Y(n_402)
);

OAI22xp5_ASAP7_75t_SL g403 ( 
.A1(n_326),
.A2(n_327),
.B1(n_316),
.B2(n_325),
.Y(n_403)
);

CKINVDCx16_ASAP7_75t_R g404 ( 
.A(n_308),
.Y(n_404)
);

NOR2xp33_ASAP7_75t_L g432 ( 
.A(n_404),
.B(n_406),
.Y(n_432)
);

OAI22xp5_ASAP7_75t_L g405 ( 
.A1(n_325),
.A2(n_313),
.B1(n_323),
.B2(n_314),
.Y(n_405)
);

OAI22xp5_ASAP7_75t_L g430 ( 
.A1(n_405),
.A2(n_408),
.B1(n_331),
.B2(n_348),
.Y(n_430)
);

INVx2_ASAP7_75t_L g406 ( 
.A(n_308),
.Y(n_406)
);

NOR2xp33_ASAP7_75t_L g407 ( 
.A(n_305),
.B(n_306),
.Y(n_407)
);

NOR2xp33_ASAP7_75t_L g438 ( 
.A(n_407),
.B(n_372),
.Y(n_438)
);

AOI22xp5_ASAP7_75t_L g408 ( 
.A1(n_313),
.A2(n_305),
.B1(n_306),
.B2(n_345),
.Y(n_408)
);

OAI21xp5_ASAP7_75t_SL g458 ( 
.A1(n_410),
.A2(n_413),
.B(n_427),
.Y(n_458)
);

CKINVDCx16_ASAP7_75t_R g417 ( 
.A(n_408),
.Y(n_417)
);

NOR2xp33_ASAP7_75t_L g451 ( 
.A(n_417),
.B(n_428),
.Y(n_451)
);

OAI22xp5_ASAP7_75t_SL g422 ( 
.A1(n_393),
.A2(n_358),
.B1(n_355),
.B2(n_309),
.Y(n_422)
);

AOI22xp5_ASAP7_75t_L g469 ( 
.A1(n_422),
.A2(n_439),
.B1(n_403),
.B2(n_374),
.Y(n_469)
);

AOI21xp5_ASAP7_75t_L g423 ( 
.A1(n_377),
.A2(n_351),
.B(n_340),
.Y(n_423)
);

AOI21xp5_ASAP7_75t_L g473 ( 
.A1(n_423),
.A2(n_364),
.B(n_384),
.Y(n_473)
);

OAI22xp5_ASAP7_75t_SL g455 ( 
.A1(n_425),
.A2(n_370),
.B1(n_365),
.B2(n_367),
.Y(n_455)
);

CKINVDCx20_ASAP7_75t_R g428 ( 
.A(n_402),
.Y(n_428)
);

HB1xp67_ASAP7_75t_L g452 ( 
.A(n_430),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_366),
.B(n_336),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_431),
.B(n_441),
.Y(n_459)
);

XOR2xp5_ASAP7_75t_L g450 ( 
.A(n_435),
.B(n_363),
.Y(n_450)
);

AOI22xp5_ASAP7_75t_SL g436 ( 
.A1(n_391),
.A2(n_345),
.B1(n_347),
.B2(n_336),
.Y(n_436)
);

OAI21xp5_ASAP7_75t_SL g471 ( 
.A1(n_436),
.A2(n_364),
.B(n_384),
.Y(n_471)
);

CKINVDCx20_ASAP7_75t_R g437 ( 
.A(n_405),
.Y(n_437)
);

NOR2xp33_ASAP7_75t_L g454 ( 
.A(n_437),
.B(n_446),
.Y(n_454)
);

NOR2xp33_ASAP7_75t_SL g463 ( 
.A(n_438),
.B(n_443),
.Y(n_463)
);

OAI22xp5_ASAP7_75t_L g439 ( 
.A1(n_368),
.A2(n_393),
.B1(n_391),
.B2(n_382),
.Y(n_439)
);

CKINVDCx14_ASAP7_75t_R g466 ( 
.A(n_440),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_366),
.B(n_335),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_368),
.B(n_349),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_442),
.B(n_444),
.Y(n_460)
);

NOR2xp33_ASAP7_75t_L g443 ( 
.A(n_401),
.B(n_349),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_SL g444 ( 
.A(n_400),
.B(n_332),
.Y(n_444)
);

CKINVDCx20_ASAP7_75t_R g446 ( 
.A(n_376),
.Y(n_446)
);

INVxp67_ASAP7_75t_L g448 ( 
.A(n_413),
.Y(n_448)
);

INVx2_ASAP7_75t_L g485 ( 
.A(n_448),
.Y(n_485)
);

OAI21xp5_ASAP7_75t_L g449 ( 
.A1(n_409),
.A2(n_379),
.B(n_397),
.Y(n_449)
);

OAI21xp5_ASAP7_75t_SL g498 ( 
.A1(n_449),
.A2(n_471),
.B(n_472),
.Y(n_498)
);

MAJIxp5_ASAP7_75t_L g513 ( 
.A(n_450),
.B(n_453),
.C(n_457),
.Y(n_513)
);

MAJIxp5_ASAP7_75t_L g453 ( 
.A(n_420),
.B(n_395),
.C(n_389),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_455),
.B(n_464),
.Y(n_506)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_412),
.Y(n_456)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_456),
.Y(n_495)
);

MAJIxp5_ASAP7_75t_L g457 ( 
.A(n_420),
.B(n_368),
.C(n_394),
.Y(n_457)
);

MAJIxp5_ASAP7_75t_L g461 ( 
.A(n_420),
.B(n_387),
.C(n_373),
.Y(n_461)
);

XNOR2xp5_ASAP7_75t_L g487 ( 
.A(n_461),
.B(n_474),
.Y(n_487)
);

CKINVDCx16_ASAP7_75t_R g462 ( 
.A(n_438),
.Y(n_462)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_462),
.Y(n_511)
);

CKINVDCx20_ASAP7_75t_R g464 ( 
.A(n_426),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_412),
.Y(n_465)
);

INVx1_ASAP7_75t_SL g493 ( 
.A(n_465),
.Y(n_493)
);

OAI21xp33_ASAP7_75t_L g467 ( 
.A1(n_409),
.A2(n_423),
.B(n_440),
.Y(n_467)
);

AOI21xp5_ASAP7_75t_L g488 ( 
.A1(n_467),
.A2(n_473),
.B(n_433),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_441),
.B(n_398),
.Y(n_468)
);

CKINVDCx20_ASAP7_75t_R g484 ( 
.A(n_468),
.Y(n_484)
);

OAI22xp5_ASAP7_75t_L g486 ( 
.A1(n_469),
.A2(n_417),
.B1(n_437),
.B2(n_434),
.Y(n_486)
);

NOR2xp33_ASAP7_75t_L g470 ( 
.A(n_416),
.B(n_428),
.Y(n_470)
);

NOR2xp33_ASAP7_75t_SL g499 ( 
.A(n_470),
.B(n_421),
.Y(n_499)
);

OAI21xp5_ASAP7_75t_L g472 ( 
.A1(n_427),
.A2(n_439),
.B(n_433),
.Y(n_472)
);

MAJIxp5_ASAP7_75t_L g474 ( 
.A(n_435),
.B(n_392),
.C(n_386),
.Y(n_474)
);

CKINVDCx20_ASAP7_75t_R g475 ( 
.A(n_426),
.Y(n_475)
);

NOR2xp33_ASAP7_75t_L g514 ( 
.A(n_475),
.B(n_478),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_431),
.B(n_383),
.Y(n_476)
);

CKINVDCx20_ASAP7_75t_R g497 ( 
.A(n_476),
.Y(n_497)
);

OAI21xp5_ASAP7_75t_L g477 ( 
.A1(n_427),
.A2(n_433),
.B(n_436),
.Y(n_477)
);

OAI21xp5_ASAP7_75t_L g503 ( 
.A1(n_477),
.A2(n_479),
.B(n_483),
.Y(n_503)
);

CKINVDCx20_ASAP7_75t_R g478 ( 
.A(n_443),
.Y(n_478)
);

NAND2x1_ASAP7_75t_SL g479 ( 
.A(n_433),
.B(n_442),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_411),
.Y(n_480)
);

INVxp67_ASAP7_75t_L g500 ( 
.A(n_480),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_415),
.B(n_404),
.Y(n_481)
);

CKINVDCx20_ASAP7_75t_R g504 ( 
.A(n_481),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_415),
.B(n_381),
.Y(n_482)
);

CKINVDCx20_ASAP7_75t_R g517 ( 
.A(n_482),
.Y(n_517)
);

OAI21xp5_ASAP7_75t_SL g483 ( 
.A1(n_436),
.A2(n_385),
.B(n_388),
.Y(n_483)
);

AOI22xp5_ASAP7_75t_L g529 ( 
.A1(n_486),
.A2(n_454),
.B1(n_467),
.B2(n_466),
.Y(n_529)
);

CKINVDCx16_ASAP7_75t_R g547 ( 
.A(n_488),
.Y(n_547)
);

NOR2x1p5_ASAP7_75t_SL g489 ( 
.A(n_468),
.B(n_414),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_489),
.B(n_501),
.Y(n_519)
);

XOR2xp5_ASAP7_75t_L g490 ( 
.A(n_457),
.B(n_435),
.Y(n_490)
);

XOR2xp5_ASAP7_75t_L g524 ( 
.A(n_490),
.B(n_492),
.Y(n_524)
);

BUFx3_ASAP7_75t_L g491 ( 
.A(n_470),
.Y(n_491)
);

BUFx2_ASAP7_75t_L g525 ( 
.A(n_491),
.Y(n_525)
);

XOR2xp5_ASAP7_75t_L g492 ( 
.A(n_457),
.B(n_444),
.Y(n_492)
);

XNOR2xp5_ASAP7_75t_SL g494 ( 
.A(n_453),
.B(n_414),
.Y(n_494)
);

XOR2xp5_ASAP7_75t_L g532 ( 
.A(n_494),
.B(n_502),
.Y(n_532)
);

XOR2x2_ASAP7_75t_L g496 ( 
.A(n_453),
.B(n_447),
.Y(n_496)
);

NOR2xp33_ASAP7_75t_L g530 ( 
.A(n_496),
.B(n_463),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_SL g538 ( 
.A(n_499),
.B(n_505),
.Y(n_538)
);

OA21x2_ASAP7_75t_L g501 ( 
.A1(n_472),
.A2(n_477),
.B(n_451),
.Y(n_501)
);

XNOR2xp5_ASAP7_75t_L g502 ( 
.A(n_461),
.B(n_450),
.Y(n_502)
);

CKINVDCx16_ASAP7_75t_R g505 ( 
.A(n_481),
.Y(n_505)
);

AOI22xp5_ASAP7_75t_L g507 ( 
.A1(n_469),
.A2(n_422),
.B1(n_430),
.B2(n_434),
.Y(n_507)
);

OAI22xp5_ASAP7_75t_SL g527 ( 
.A1(n_507),
.A2(n_508),
.B1(n_518),
.B2(n_477),
.Y(n_527)
);

AOI22xp5_ASAP7_75t_L g508 ( 
.A1(n_469),
.A2(n_451),
.B1(n_452),
.B2(n_472),
.Y(n_508)
);

OA22x2_ASAP7_75t_L g509 ( 
.A1(n_452),
.A2(n_425),
.B1(n_410),
.B2(n_429),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_509),
.B(n_483),
.Y(n_521)
);

OAI22xp5_ASAP7_75t_L g510 ( 
.A1(n_462),
.A2(n_447),
.B1(n_466),
.B2(n_463),
.Y(n_510)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_510),
.Y(n_522)
);

XNOR2xp5_ASAP7_75t_L g512 ( 
.A(n_461),
.B(n_421),
.Y(n_512)
);

XOR2xp5_ASAP7_75t_L g534 ( 
.A(n_512),
.B(n_515),
.Y(n_534)
);

XNOR2xp5_ASAP7_75t_L g515 ( 
.A(n_450),
.B(n_449),
.Y(n_515)
);

XOR2xp5_ASAP7_75t_L g516 ( 
.A(n_449),
.B(n_460),
.Y(n_516)
);

XOR2xp5_ASAP7_75t_L g543 ( 
.A(n_516),
.B(n_479),
.Y(n_543)
);

AOI22xp5_ASAP7_75t_SL g518 ( 
.A1(n_464),
.A2(n_429),
.B1(n_380),
.B2(n_432),
.Y(n_518)
);

FAx1_ASAP7_75t_SL g520 ( 
.A(n_484),
.B(n_496),
.CI(n_515),
.CON(n_520),
.SN(n_520)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_520),
.B(n_540),
.Y(n_551)
);

AND2x2_ASAP7_75t_L g550 ( 
.A(n_521),
.B(n_544),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g523 ( 
.A(n_500),
.B(n_475),
.Y(n_523)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_523),
.Y(n_574)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_506),
.Y(n_526)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_526),
.Y(n_553)
);

AOI22xp5_ASAP7_75t_L g568 ( 
.A1(n_527),
.A2(n_498),
.B1(n_458),
.B2(n_479),
.Y(n_568)
);

MAJIxp5_ASAP7_75t_L g528 ( 
.A(n_490),
.B(n_460),
.C(n_474),
.Y(n_528)
);

MAJIxp5_ASAP7_75t_L g554 ( 
.A(n_528),
.B(n_494),
.C(n_512),
.Y(n_554)
);

OAI22xp5_ASAP7_75t_L g557 ( 
.A1(n_529),
.A2(n_544),
.B1(n_508),
.B2(n_521),
.Y(n_557)
);

OAI21xp33_ASAP7_75t_L g555 ( 
.A1(n_530),
.A2(n_513),
.B(n_485),
.Y(n_555)
);

NOR2xp33_ASAP7_75t_L g531 ( 
.A(n_511),
.B(n_478),
.Y(n_531)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_531),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_500),
.B(n_454),
.Y(n_533)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_533),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_506),
.B(n_459),
.Y(n_535)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_535),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_L g536 ( 
.A(n_514),
.B(n_459),
.Y(n_536)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_536),
.Y(n_570)
);

XNOR2xp5_ASAP7_75t_L g537 ( 
.A(n_492),
.B(n_474),
.Y(n_537)
);

XNOR2xp5_ASAP7_75t_L g560 ( 
.A(n_537),
.B(n_543),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_497),
.B(n_482),
.Y(n_539)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_539),
.Y(n_562)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_493),
.Y(n_540)
);

CKINVDCx20_ASAP7_75t_R g541 ( 
.A(n_501),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_L g561 ( 
.A(n_541),
.B(n_542),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_L g542 ( 
.A(n_504),
.B(n_476),
.Y(n_542)
);

AOI22xp5_ASAP7_75t_L g544 ( 
.A1(n_507),
.A2(n_473),
.B1(n_458),
.B2(n_455),
.Y(n_544)
);

CKINVDCx20_ASAP7_75t_R g545 ( 
.A(n_503),
.Y(n_545)
);

NOR2xp33_ASAP7_75t_L g564 ( 
.A(n_545),
.B(n_546),
.Y(n_564)
);

NOR2xp33_ASAP7_75t_L g546 ( 
.A(n_491),
.B(n_419),
.Y(n_546)
);

XNOR2xp5_ASAP7_75t_L g548 ( 
.A(n_487),
.B(n_479),
.Y(n_548)
);

XNOR2xp5_ASAP7_75t_L g569 ( 
.A(n_548),
.B(n_498),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_L g549 ( 
.A(n_517),
.B(n_465),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_L g572 ( 
.A(n_549),
.B(n_456),
.Y(n_572)
);

INVxp33_ASAP7_75t_L g586 ( 
.A(n_550),
.Y(n_586)
);

XOR2xp5_ASAP7_75t_L g552 ( 
.A(n_524),
.B(n_502),
.Y(n_552)
);

XOR2xp5_ASAP7_75t_L g583 ( 
.A(n_552),
.B(n_523),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_SL g589 ( 
.A(n_554),
.B(n_571),
.Y(n_589)
);

OAI22xp5_ASAP7_75t_L g584 ( 
.A1(n_555),
.A2(n_567),
.B1(n_568),
.B2(n_547),
.Y(n_584)
);

XNOR2x1_ASAP7_75t_L g594 ( 
.A(n_557),
.B(n_569),
.Y(n_594)
);

MAJIxp5_ASAP7_75t_L g558 ( 
.A(n_524),
.B(n_487),
.C(n_513),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_L g580 ( 
.A(n_558),
.B(n_559),
.Y(n_580)
);

MAJIxp5_ASAP7_75t_L g559 ( 
.A(n_537),
.B(n_516),
.C(n_501),
.Y(n_559)
);

OAI22xp5_ASAP7_75t_SL g563 ( 
.A1(n_522),
.A2(n_526),
.B1(n_529),
.B2(n_519),
.Y(n_563)
);

HB1xp67_ASAP7_75t_L g575 ( 
.A(n_563),
.Y(n_575)
);

OAI22xp5_ASAP7_75t_SL g566 ( 
.A1(n_522),
.A2(n_518),
.B1(n_488),
.B2(n_503),
.Y(n_566)
);

HB1xp67_ASAP7_75t_L g577 ( 
.A(n_566),
.Y(n_577)
);

OAI22xp5_ASAP7_75t_L g567 ( 
.A1(n_538),
.A2(n_485),
.B1(n_493),
.B2(n_489),
.Y(n_567)
);

MAJIxp5_ASAP7_75t_L g571 ( 
.A(n_528),
.B(n_509),
.C(n_432),
.Y(n_571)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_572),
.Y(n_585)
);

MAJIxp5_ASAP7_75t_L g576 ( 
.A(n_558),
.B(n_534),
.C(n_532),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_SL g601 ( 
.A(n_576),
.B(n_578),
.Y(n_601)
);

MAJIxp5_ASAP7_75t_L g578 ( 
.A(n_554),
.B(n_534),
.C(n_532),
.Y(n_578)
);

XNOR2xp5_ASAP7_75t_L g579 ( 
.A(n_559),
.B(n_571),
.Y(n_579)
);

XNOR2xp5_ASAP7_75t_L g611 ( 
.A(n_579),
.B(n_583),
.Y(n_611)
);

MAJIxp5_ASAP7_75t_L g581 ( 
.A(n_552),
.B(n_560),
.C(n_548),
.Y(n_581)
);

MAJIxp5_ASAP7_75t_L g599 ( 
.A(n_581),
.B(n_587),
.C(n_576),
.Y(n_599)
);

CKINVDCx20_ASAP7_75t_R g582 ( 
.A(n_572),
.Y(n_582)
);

AOI22xp33_ASAP7_75t_SL g609 ( 
.A1(n_582),
.A2(n_584),
.B1(n_520),
.B2(n_495),
.Y(n_609)
);

MAJIxp5_ASAP7_75t_L g587 ( 
.A(n_560),
.B(n_543),
.C(n_541),
.Y(n_587)
);

XNOR2xp5_ASAP7_75t_L g588 ( 
.A(n_564),
.B(n_519),
.Y(n_588)
);

XNOR2xp5_ASAP7_75t_L g612 ( 
.A(n_588),
.B(n_595),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_SL g590 ( 
.A(n_556),
.B(n_570),
.Y(n_590)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_590),
.Y(n_602)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_562),
.Y(n_591)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_591),
.Y(n_608)
);

NOR2xp33_ASAP7_75t_SL g592 ( 
.A(n_551),
.B(n_536),
.Y(n_592)
);

OAI22xp5_ASAP7_75t_L g597 ( 
.A1(n_592),
.A2(n_565),
.B1(n_551),
.B2(n_574),
.Y(n_597)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_562),
.Y(n_593)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_593),
.Y(n_596)
);

XNOR2xp5_ASAP7_75t_L g595 ( 
.A(n_566),
.B(n_527),
.Y(n_595)
);

AOI22xp33_ASAP7_75t_L g622 ( 
.A1(n_597),
.A2(n_613),
.B1(n_578),
.B2(n_429),
.Y(n_622)
);

OAI21xp5_ASAP7_75t_SL g598 ( 
.A1(n_586),
.A2(n_561),
.B(n_568),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_L g616 ( 
.A(n_598),
.B(n_604),
.Y(n_616)
);

XNOR2xp5_ASAP7_75t_L g617 ( 
.A(n_599),
.B(n_581),
.Y(n_617)
);

AOI22xp5_ASAP7_75t_L g600 ( 
.A1(n_575),
.A2(n_563),
.B1(n_553),
.B2(n_573),
.Y(n_600)
);

OAI22xp5_ASAP7_75t_SL g625 ( 
.A1(n_600),
.A2(n_603),
.B1(n_607),
.B2(n_411),
.Y(n_625)
);

AOI22xp5_ASAP7_75t_L g603 ( 
.A1(n_577),
.A2(n_550),
.B1(n_561),
.B2(n_533),
.Y(n_603)
);

OAI21xp5_ASAP7_75t_SL g604 ( 
.A1(n_586),
.A2(n_550),
.B(n_539),
.Y(n_604)
);

MAJIxp5_ASAP7_75t_L g605 ( 
.A(n_583),
.B(n_569),
.C(n_525),
.Y(n_605)
);

MAJIxp5_ASAP7_75t_L g615 ( 
.A(n_605),
.B(n_606),
.C(n_587),
.Y(n_615)
);

MAJIxp5_ASAP7_75t_L g606 ( 
.A(n_579),
.B(n_525),
.C(n_540),
.Y(n_606)
);

AOI22xp5_ASAP7_75t_L g607 ( 
.A1(n_585),
.A2(n_549),
.B1(n_535),
.B2(n_542),
.Y(n_607)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_609),
.Y(n_614)
);

OAI22xp5_ASAP7_75t_SL g610 ( 
.A1(n_595),
.A2(n_520),
.B1(n_509),
.B2(n_480),
.Y(n_610)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_610),
.Y(n_626)
);

INVx1_ASAP7_75t_SL g613 ( 
.A(n_588),
.Y(n_613)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_615),
.Y(n_629)
);

NOR2xp33_ASAP7_75t_SL g638 ( 
.A(n_617),
.B(n_618),
.Y(n_638)
);

NOR2xp33_ASAP7_75t_SL g618 ( 
.A(n_601),
.B(n_589),
.Y(n_618)
);

NOR2xp33_ASAP7_75t_L g619 ( 
.A(n_606),
.B(n_612),
.Y(n_619)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_619),
.Y(n_632)
);

MAJIxp5_ASAP7_75t_L g620 ( 
.A(n_611),
.B(n_580),
.C(n_594),
.Y(n_620)
);

MAJIxp5_ASAP7_75t_L g630 ( 
.A(n_620),
.B(n_599),
.C(n_613),
.Y(n_630)
);

NOR2xp33_ASAP7_75t_L g621 ( 
.A(n_612),
.B(n_594),
.Y(n_621)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_621),
.Y(n_635)
);

NOR2xp33_ASAP7_75t_L g634 ( 
.A(n_622),
.B(n_624),
.Y(n_634)
);

OR2x2_ASAP7_75t_L g623 ( 
.A(n_603),
.B(n_509),
.Y(n_623)
);

AOI21xp5_ASAP7_75t_L g631 ( 
.A1(n_623),
.A2(n_598),
.B(n_604),
.Y(n_631)
);

CKINVDCx20_ASAP7_75t_R g624 ( 
.A(n_607),
.Y(n_624)
);

AOI22xp5_ASAP7_75t_L g628 ( 
.A1(n_625),
.A2(n_610),
.B1(n_596),
.B2(n_600),
.Y(n_628)
);

XOR2xp5_ASAP7_75t_L g627 ( 
.A(n_605),
.B(n_611),
.Y(n_627)
);

NOR2xp33_ASAP7_75t_L g637 ( 
.A(n_627),
.B(n_424),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_L g645 ( 
.A(n_628),
.B(n_630),
.Y(n_645)
);

NOR2xp33_ASAP7_75t_L g642 ( 
.A(n_631),
.B(n_636),
.Y(n_642)
);

AOI21xp5_ASAP7_75t_L g633 ( 
.A1(n_617),
.A2(n_602),
.B(n_596),
.Y(n_633)
);

AOI21xp5_ASAP7_75t_L g641 ( 
.A1(n_633),
.A2(n_620),
.B(n_615),
.Y(n_641)
);

XNOR2xp5_ASAP7_75t_SL g636 ( 
.A(n_616),
.B(n_608),
.Y(n_636)
);

NOR2xp33_ASAP7_75t_L g639 ( 
.A(n_637),
.B(n_635),
.Y(n_639)
);

XNOR2xp5_ASAP7_75t_L g647 ( 
.A(n_639),
.B(n_636),
.Y(n_647)
);

OAI21xp5_ASAP7_75t_SL g640 ( 
.A1(n_629),
.A2(n_616),
.B(n_614),
.Y(n_640)
);

AOI21xp5_ASAP7_75t_L g649 ( 
.A1(n_640),
.A2(n_644),
.B(n_646),
.Y(n_649)
);

OAI321xp33_ASAP7_75t_L g648 ( 
.A1(n_641),
.A2(n_643),
.A3(n_623),
.B1(n_628),
.B2(n_424),
.C(n_419),
.Y(n_648)
);

NOR2xp33_ASAP7_75t_SL g643 ( 
.A(n_632),
.B(n_638),
.Y(n_643)
);

NOR2xp33_ASAP7_75t_L g644 ( 
.A(n_630),
.B(n_627),
.Y(n_644)
);

OAI21xp5_ASAP7_75t_L g646 ( 
.A1(n_634),
.A2(n_626),
.B(n_625),
.Y(n_646)
);

AOI21xp5_ASAP7_75t_L g652 ( 
.A1(n_647),
.A2(n_648),
.B(n_650),
.Y(n_652)
);

AOI21xp5_ASAP7_75t_L g650 ( 
.A1(n_642),
.A2(n_471),
.B(n_446),
.Y(n_650)
);

OAI21xp5_ASAP7_75t_SL g651 ( 
.A1(n_645),
.A2(n_418),
.B(n_445),
.Y(n_651)
);

OAI21xp5_ASAP7_75t_SL g654 ( 
.A1(n_651),
.A2(n_445),
.B(n_406),
.Y(n_654)
);

OAI21xp5_ASAP7_75t_L g653 ( 
.A1(n_649),
.A2(n_639),
.B(n_445),
.Y(n_653)
);

OAI21xp5_ASAP7_75t_SL g655 ( 
.A1(n_653),
.A2(n_654),
.B(n_445),
.Y(n_655)
);

OAI321xp33_ASAP7_75t_L g656 ( 
.A1(n_655),
.A2(n_652),
.A3(n_418),
.B1(n_455),
.B2(n_376),
.C(n_347),
.Y(n_656)
);

AND2x2_ASAP7_75t_L g657 ( 
.A(n_656),
.B(n_399),
.Y(n_657)
);

MAJIxp5_ASAP7_75t_L g658 ( 
.A(n_657),
.B(n_399),
.C(n_390),
.Y(n_658)
);

MAJIxp5_ASAP7_75t_L g659 ( 
.A(n_658),
.B(n_380),
.C(n_332),
.Y(n_659)
);

XNOR2xp5_ASAP7_75t_L g660 ( 
.A(n_659),
.B(n_357),
.Y(n_660)
);


endmodule