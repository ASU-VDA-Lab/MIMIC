module fake_jpeg_22928_n_266 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_266);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_266;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_187;
wire n_21;
wire n_57;
wire n_234;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_33;
wire n_91;
wire n_54;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_258;
wire n_96;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_8),
.Y(n_15)
);

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_8),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_2),
.Y(n_22)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

INVx5_ASAP7_75t_L g32 ( 
.A(n_21),
.Y(n_32)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_32),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_20),
.Y(n_33)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_33),
.Y(n_55)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_34),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_20),
.Y(n_35)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

BUFx2_ASAP7_75t_L g58 ( 
.A(n_36),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_20),
.Y(n_37)
);

INVx11_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_38),
.A2(n_23),
.B1(n_28),
.B2(n_31),
.Y(n_48)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_21),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_39),
.B(n_41),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_20),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_40),
.Y(n_44)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_20),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_23),
.Y(n_42)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_42),
.Y(n_62)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_36),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_43),
.B(n_49),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_41),
.B(n_30),
.Y(n_45)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_45),
.B(n_56),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_36),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_46),
.B(n_52),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_48),
.A2(n_53),
.B1(n_19),
.B2(n_27),
.Y(n_86)
);

CKINVDCx5p33_ASAP7_75t_R g49 ( 
.A(n_34),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_50),
.B(n_59),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_39),
.B(n_19),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_38),
.A2(n_23),
.B1(n_31),
.B2(n_28),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_33),
.B(n_30),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_42),
.B(n_17),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_32),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_60),
.Y(n_77)
);

OAI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_35),
.A2(n_31),
.B1(n_26),
.B2(n_21),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_61),
.A2(n_26),
.B1(n_16),
.B2(n_27),
.Y(n_74)
);

INVx2_ASAP7_75t_SL g64 ( 
.A(n_37),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_64),
.B(n_0),
.Y(n_82)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_59),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_65),
.B(n_68),
.Y(n_93)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_45),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_56),
.Y(n_69)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_69),
.Y(n_88)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_52),
.Y(n_71)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_71),
.Y(n_107)
);

AO22x1_ASAP7_75t_L g72 ( 
.A1(n_63),
.A2(n_16),
.B1(n_26),
.B2(n_28),
.Y(n_72)
);

AO22x2_ASAP7_75t_L g106 ( 
.A1(n_72),
.A2(n_64),
.B1(n_44),
.B2(n_55),
.Y(n_106)
);

AND2x2_ASAP7_75t_SL g73 ( 
.A(n_46),
.B(n_16),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_73),
.B(n_62),
.C(n_63),
.Y(n_87)
);

OAI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_74),
.A2(n_78),
.B1(n_80),
.B2(n_55),
.Y(n_103)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_47),
.Y(n_76)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_76),
.Y(n_109)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_47),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_L g79 ( 
.A1(n_57),
.A2(n_29),
.B1(n_15),
.B2(n_18),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_79),
.A2(n_84),
.B1(n_17),
.B2(n_24),
.Y(n_99)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_58),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_49),
.B(n_29),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_81),
.B(n_60),
.Y(n_89)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_82),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_58),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_83),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_L g84 ( 
.A1(n_57),
.A2(n_29),
.B1(n_15),
.B2(n_18),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_58),
.Y(n_85)
);

NOR3xp33_ASAP7_75t_L g105 ( 
.A(n_85),
.B(n_63),
.C(n_25),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_86),
.A2(n_24),
.B1(n_25),
.B2(n_51),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_87),
.B(n_92),
.C(n_73),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_89),
.B(n_90),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_70),
.B(n_62),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_74),
.A2(n_51),
.B1(n_55),
.B2(n_64),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_91),
.A2(n_84),
.B1(n_79),
.B2(n_85),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_L g92 ( 
.A(n_70),
.B(n_63),
.Y(n_92)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_83),
.Y(n_95)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_95),
.Y(n_124)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_72),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_96),
.B(n_104),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_70),
.B(n_60),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_98),
.B(n_100),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_99),
.A2(n_71),
.B1(n_65),
.B2(n_76),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_70),
.B(n_40),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_69),
.B(n_51),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_101),
.B(n_77),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_102),
.Y(n_128)
);

CKINVDCx16_ASAP7_75t_R g120 ( 
.A(n_103),
.Y(n_120)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_72),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_105),
.B(n_108),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_106),
.A2(n_80),
.B1(n_54),
.B2(n_50),
.Y(n_126)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_75),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_97),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_110),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_89),
.B(n_68),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_111),
.B(n_115),
.Y(n_142)
);

AOI21xp5_ASAP7_75t_L g113 ( 
.A1(n_98),
.A2(n_81),
.B(n_67),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_L g136 ( 
.A1(n_113),
.A2(n_118),
.B(n_129),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_117),
.B(n_88),
.C(n_94),
.Y(n_143)
);

AOI21xp5_ASAP7_75t_L g118 ( 
.A1(n_96),
.A2(n_67),
.B(n_75),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_121),
.A2(n_77),
.B1(n_43),
.B2(n_44),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_90),
.B(n_100),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_122),
.B(n_99),
.Y(n_151)
);

INVx8_ASAP7_75t_L g123 ( 
.A(n_106),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_123),
.B(n_106),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_125),
.A2(n_126),
.B1(n_131),
.B2(n_91),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_109),
.B(n_66),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_127),
.B(n_109),
.Y(n_138)
);

OR2x2_ASAP7_75t_SL g129 ( 
.A(n_106),
.B(n_73),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_101),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_130),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_104),
.A2(n_66),
.B1(n_78),
.B2(n_54),
.Y(n_131)
);

AND2x2_ASAP7_75t_L g132 ( 
.A(n_92),
.B(n_73),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_L g146 ( 
.A1(n_132),
.A2(n_106),
.B(n_107),
.Y(n_146)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_126),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_134),
.B(n_135),
.Y(n_158)
);

CKINVDCx16_ASAP7_75t_R g135 ( 
.A(n_115),
.Y(n_135)
);

INVxp67_ASAP7_75t_L g137 ( 
.A(n_126),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_137),
.B(n_138),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_139),
.A2(n_150),
.B1(n_154),
.B2(n_123),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_117),
.B(n_87),
.C(n_88),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_140),
.B(n_143),
.C(n_145),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_110),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_144),
.B(n_127),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_117),
.B(n_93),
.C(n_107),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_L g164 ( 
.A1(n_146),
.A2(n_152),
.B(n_116),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_124),
.B(n_95),
.Y(n_147)
);

CKINVDCx14_ASAP7_75t_R g175 ( 
.A(n_147),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_124),
.B(n_82),
.Y(n_148)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_148),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_114),
.B(n_122),
.C(n_112),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_149),
.B(n_130),
.C(n_118),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_151),
.B(n_155),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_L g152 ( 
.A1(n_114),
.A2(n_22),
.B(n_1),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_112),
.B(n_77),
.Y(n_153)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_153),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_111),
.B(n_22),
.Y(n_155)
);

A2O1A1O1Ixp25_ASAP7_75t_L g159 ( 
.A1(n_136),
.A2(n_132),
.B(n_129),
.C(n_116),
.D(n_119),
.Y(n_159)
);

MAJx2_ASAP7_75t_L g192 ( 
.A(n_159),
.B(n_132),
.C(n_152),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_139),
.A2(n_128),
.B1(n_120),
.B2(n_123),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_160),
.A2(n_151),
.B1(n_135),
.B2(n_141),
.Y(n_190)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_147),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_161),
.B(n_169),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_140),
.B(n_113),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_162),
.B(n_140),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_163),
.B(n_156),
.C(n_149),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_L g183 ( 
.A1(n_164),
.A2(n_165),
.B(n_146),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_L g165 ( 
.A1(n_136),
.A2(n_129),
.B(n_120),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_166),
.A2(n_177),
.B1(n_150),
.B2(n_131),
.Y(n_179)
);

INVx1_ASAP7_75t_SL g168 ( 
.A(n_138),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_168),
.B(n_176),
.Y(n_182)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_153),
.Y(n_169)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_142),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_171),
.B(n_174),
.Y(n_191)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_172),
.Y(n_187)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_142),
.Y(n_174)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_148),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_154),
.A2(n_125),
.B1(n_119),
.B2(n_121),
.Y(n_177)
);

AND2x2_ASAP7_75t_L g178 ( 
.A(n_175),
.B(n_141),
.Y(n_178)
);

AOI21xp5_ASAP7_75t_L g199 ( 
.A1(n_178),
.A2(n_195),
.B(n_170),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_179),
.A2(n_157),
.B1(n_176),
.B2(n_164),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_158),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_180),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_SL g181 ( 
.A(n_173),
.B(n_133),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_181),
.B(n_194),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_183),
.B(n_186),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_168),
.B(n_144),
.Y(n_184)
);

CKINVDCx14_ASAP7_75t_R g204 ( 
.A(n_184),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_162),
.B(n_143),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_188),
.B(n_189),
.C(n_192),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_156),
.B(n_145),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_190),
.A2(n_197),
.B1(n_161),
.B2(n_7),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_193),
.B(n_163),
.C(n_159),
.Y(n_203)
);

NAND3xp33_ASAP7_75t_L g194 ( 
.A(n_167),
.B(n_132),
.C(n_133),
.Y(n_194)
);

XOR2x2_ASAP7_75t_L g195 ( 
.A(n_165),
.B(n_155),
.Y(n_195)
);

CKINVDCx14_ASAP7_75t_R g196 ( 
.A(n_177),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_196),
.B(n_6),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_160),
.A2(n_44),
.B1(n_1),
.B2(n_2),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_SL g198 ( 
.A(n_182),
.B(n_173),
.Y(n_198)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_198),
.Y(n_215)
);

AOI21xp5_ASAP7_75t_L g218 ( 
.A1(n_199),
.A2(n_202),
.B(n_212),
.Y(n_218)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_185),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_203),
.B(n_200),
.C(n_199),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_178),
.B(n_171),
.Y(n_206)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_206),
.Y(n_225)
);

CKINVDCx14_ASAP7_75t_R g207 ( 
.A(n_191),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_207),
.B(n_209),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_179),
.A2(n_195),
.B1(n_157),
.B2(n_192),
.Y(n_208)
);

CKINVDCx16_ASAP7_75t_R g221 ( 
.A(n_208),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_210),
.B(n_187),
.Y(n_216)
);

CKINVDCx14_ASAP7_75t_R g213 ( 
.A(n_197),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_213),
.B(n_183),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_211),
.B(n_193),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_214),
.B(n_220),
.Y(n_229)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_216),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_219),
.B(n_224),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_200),
.B(n_186),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_222),
.B(n_226),
.Y(n_238)
);

A2O1A1Ixp33_ASAP7_75t_SL g223 ( 
.A1(n_206),
.A2(n_189),
.B(n_188),
.C(n_2),
.Y(n_223)
);

AOI21xp5_ASAP7_75t_L g234 ( 
.A1(n_223),
.A2(n_10),
.B(n_13),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_204),
.B(n_6),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_211),
.B(n_7),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_SL g227 ( 
.A(n_201),
.B(n_5),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_SL g236 ( 
.A(n_227),
.B(n_5),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_225),
.A2(n_208),
.B1(n_202),
.B2(n_205),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_228),
.A2(n_234),
.B1(n_221),
.B2(n_223),
.Y(n_242)
);

AOI322xp5_ASAP7_75t_SL g230 ( 
.A1(n_223),
.A2(n_203),
.A3(n_201),
.B1(n_198),
.B2(n_210),
.C1(n_4),
.C2(n_5),
.Y(n_230)
);

NOR2x1_ASAP7_75t_L g239 ( 
.A(n_230),
.B(n_234),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_SL g231 ( 
.A(n_218),
.B(n_9),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_231),
.Y(n_243)
);

AO221x1_ASAP7_75t_L g232 ( 
.A1(n_223),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.C(n_3),
.Y(n_232)
);

OR2x2_ASAP7_75t_L g246 ( 
.A(n_232),
.B(n_0),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_215),
.B(n_10),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_235),
.B(n_236),
.Y(n_241)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_239),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_237),
.B(n_217),
.Y(n_240)
);

AOI21xp5_ASAP7_75t_L g251 ( 
.A1(n_240),
.A2(n_247),
.B(n_229),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_242),
.B(n_244),
.Y(n_249)
);

AND2x2_ASAP7_75t_L g244 ( 
.A(n_238),
.B(n_222),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_233),
.B(n_226),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_245),
.B(n_246),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_228),
.B(n_214),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_243),
.B(n_238),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_248),
.B(n_253),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_SL g255 ( 
.A(n_251),
.B(n_241),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_240),
.B(n_229),
.Y(n_253)
);

A2O1A1Ixp33_ASAP7_75t_SL g254 ( 
.A1(n_249),
.A2(n_246),
.B(n_244),
.C(n_220),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_L g259 ( 
.A1(n_254),
.A2(n_255),
.B1(n_252),
.B2(n_258),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_248),
.B(n_9),
.C(n_11),
.Y(n_256)
);

OAI21xp5_ASAP7_75t_SL g261 ( 
.A1(n_256),
.A2(n_254),
.B(n_13),
.Y(n_261)
);

OAI21x1_ASAP7_75t_L g257 ( 
.A1(n_250),
.A2(n_9),
.B(n_11),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_257),
.B(n_13),
.Y(n_260)
);

AOI21xp5_ASAP7_75t_L g262 ( 
.A1(n_259),
.A2(n_260),
.B(n_261),
.Y(n_262)
);

AOI21xp5_ASAP7_75t_L g263 ( 
.A1(n_261),
.A2(n_14),
.B(n_0),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_263),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_264),
.B(n_262),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_265),
.B(n_14),
.Y(n_266)
);


endmodule