module fake_jpeg_18339_n_293 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_293);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_293;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_13;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_270;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_265;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

BUFx3_ASAP7_75t_L g13 ( 
.A(n_5),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_11),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_4),
.Y(n_15)
);

INVxp33_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

CKINVDCx16_ASAP7_75t_R g18 ( 
.A(n_4),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_11),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_9),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_1),
.Y(n_24)
);

INVx11_ASAP7_75t_SL g25 ( 
.A(n_12),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

INVx11_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_17),
.Y(n_28)
);

BUFx2_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_22),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_29),
.B(n_30),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_22),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_16),
.B(n_14),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_31),
.B(n_33),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_17),
.Y(n_32)
);

INVx5_ASAP7_75t_L g39 ( 
.A(n_32),
.Y(n_39)
);

INVx5_ASAP7_75t_L g33 ( 
.A(n_17),
.Y(n_33)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_17),
.Y(n_34)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g35 ( 
.A(n_14),
.B(n_12),
.Y(n_35)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_35),
.Y(n_41)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_22),
.Y(n_36)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_17),
.Y(n_37)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g40 ( 
.A1(n_34),
.A2(n_27),
.B1(n_18),
.B2(n_24),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_40),
.A2(n_42),
.B1(n_44),
.B2(n_46),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g42 ( 
.A1(n_34),
.A2(n_27),
.B1(n_15),
.B2(n_24),
.Y(n_42)
);

AOI21xp33_ASAP7_75t_SL g43 ( 
.A1(n_37),
.A2(n_25),
.B(n_16),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g56 ( 
.A(n_43),
.B(n_31),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g44 ( 
.A1(n_34),
.A2(n_27),
.B1(n_18),
.B2(n_24),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_33),
.A2(n_27),
.B1(n_25),
.B2(n_15),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g47 ( 
.A1(n_29),
.A2(n_21),
.B1(n_15),
.B2(n_18),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_47),
.B(n_29),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_49),
.Y(n_52)
);

BUFx2_ASAP7_75t_L g77 ( 
.A(n_52),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_41),
.B(n_35),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_53),
.B(n_54),
.Y(n_76)
);

INVxp33_ASAP7_75t_L g54 ( 
.A(n_46),
.Y(n_54)
);

BUFx2_ASAP7_75t_L g55 ( 
.A(n_49),
.Y(n_55)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_55),
.Y(n_85)
);

AOI21xp5_ASAP7_75t_L g94 ( 
.A1(n_56),
.A2(n_20),
.B(n_12),
.Y(n_94)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_45),
.Y(n_57)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_57),
.Y(n_88)
);

HB1xp67_ASAP7_75t_L g58 ( 
.A(n_45),
.Y(n_58)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_58),
.Y(n_95)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_45),
.Y(n_59)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_59),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_41),
.B(n_35),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_60),
.B(n_65),
.Y(n_78)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_39),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_61),
.A2(n_64),
.B1(n_33),
.B2(n_37),
.Y(n_80)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_38),
.Y(n_62)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_62),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_39),
.Y(n_63)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_63),
.Y(n_96)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_39),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_48),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_48),
.B(n_30),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_66),
.B(n_69),
.Y(n_81)
);

NAND3xp33_ASAP7_75t_SL g86 ( 
.A(n_68),
.B(n_44),
.C(n_36),
.Y(n_86)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_40),
.Y(n_69)
);

BUFx12f_ASAP7_75t_L g70 ( 
.A(n_51),
.Y(n_70)
);

INVx13_ASAP7_75t_L g82 ( 
.A(n_70),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_50),
.B(n_30),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_71),
.B(n_72),
.Y(n_87)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_43),
.Y(n_72)
);

BUFx2_ASAP7_75t_L g73 ( 
.A(n_42),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_73),
.B(n_38),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_67),
.A2(n_51),
.B1(n_50),
.B2(n_47),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_74),
.B(n_79),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_68),
.B(n_51),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_80),
.Y(n_101)
);

AO22x1_ASAP7_75t_SL g83 ( 
.A1(n_69),
.A2(n_73),
.B1(n_72),
.B2(n_56),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_83),
.B(n_84),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_65),
.A2(n_44),
.B1(n_40),
.B2(n_33),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_86),
.B(n_32),
.Y(n_115)
);

OAI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_89),
.A2(n_62),
.B1(n_59),
.B2(n_64),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_54),
.A2(n_36),
.B1(n_21),
.B2(n_14),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_90),
.A2(n_61),
.B1(n_38),
.B2(n_37),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_70),
.B(n_20),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_91),
.B(n_92),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_70),
.B(n_20),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_94),
.B(n_21),
.Y(n_109)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_95),
.Y(n_97)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_97),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_81),
.B(n_70),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_98),
.B(n_110),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_99),
.B(n_117),
.Y(n_120)
);

BUFx3_ASAP7_75t_L g100 ( 
.A(n_88),
.Y(n_100)
);

BUFx2_ASAP7_75t_SL g136 ( 
.A(n_100),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_85),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_102),
.B(n_103),
.Y(n_142)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_88),
.Y(n_103)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_77),
.Y(n_104)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_104),
.Y(n_119)
);

BUFx12f_ASAP7_75t_L g105 ( 
.A(n_88),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_105),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_SL g121 ( 
.A(n_109),
.B(n_90),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_81),
.B(n_55),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_87),
.B(n_57),
.C(n_52),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_111),
.B(n_115),
.Y(n_123)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_95),
.Y(n_112)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_112),
.Y(n_132)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_113),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_93),
.A2(n_63),
.B1(n_57),
.B2(n_23),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_114),
.A2(n_118),
.B1(n_104),
.B2(n_93),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_79),
.B(n_28),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_116),
.B(n_84),
.Y(n_124)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_85),
.Y(n_117)
);

INVx4_ASAP7_75t_SL g118 ( 
.A(n_75),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_SL g164 ( 
.A(n_121),
.B(n_141),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_124),
.B(n_131),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_L g126 ( 
.A1(n_101),
.A2(n_76),
.B(n_83),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_SL g148 ( 
.A1(n_126),
.A2(n_133),
.B(n_74),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_L g128 ( 
.A1(n_113),
.A2(n_89),
.B1(n_86),
.B2(n_76),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_128),
.A2(n_130),
.B1(n_134),
.B2(n_135),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_117),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_129),
.B(n_77),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_108),
.A2(n_74),
.B1(n_115),
.B2(n_107),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_116),
.B(n_78),
.Y(n_131)
);

AOI21xp5_ASAP7_75t_L g133 ( 
.A1(n_108),
.A2(n_83),
.B(n_87),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_103),
.A2(n_96),
.B1(n_80),
.B2(n_75),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_L g137 ( 
.A1(n_107),
.A2(n_90),
.B(n_98),
.Y(n_137)
);

AOI21xp5_ASAP7_75t_L g162 ( 
.A1(n_137),
.A2(n_82),
.B(n_1),
.Y(n_162)
);

INVxp67_ASAP7_75t_L g139 ( 
.A(n_110),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_139),
.B(n_140),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_106),
.B(n_83),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g141 ( 
.A(n_106),
.B(n_78),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_118),
.A2(n_96),
.B1(n_75),
.B2(n_83),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_143),
.A2(n_118),
.B1(n_92),
.B2(n_82),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_142),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_144),
.B(n_152),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_L g145 ( 
.A1(n_126),
.A2(n_94),
.B(n_109),
.Y(n_145)
);

AOI21xp5_ASAP7_75t_L g191 ( 
.A1(n_145),
.A2(n_148),
.B(n_0),
.Y(n_191)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_142),
.Y(n_146)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_146),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_141),
.B(n_100),
.Y(n_147)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_147),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_123),
.B(n_111),
.C(n_112),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_150),
.B(n_154),
.C(n_155),
.Y(n_179)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_125),
.Y(n_151)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_151),
.Y(n_192)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_125),
.Y(n_152)
);

OR2x2_ASAP7_75t_L g153 ( 
.A(n_140),
.B(n_102),
.Y(n_153)
);

INVx1_ASAP7_75t_SL g177 ( 
.A(n_153),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_123),
.B(n_97),
.C(n_105),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_133),
.B(n_105),
.C(n_91),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_156),
.A2(n_159),
.B1(n_28),
.B2(n_19),
.Y(n_190)
);

INVx1_ASAP7_75t_SL g157 ( 
.A(n_132),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_157),
.B(n_165),
.Y(n_188)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_132),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_158),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_143),
.A2(n_77),
.B1(n_82),
.B2(n_38),
.Y(n_159)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_122),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_161),
.Y(n_178)
);

O2A1O1Ixp33_ASAP7_75t_L g189 ( 
.A1(n_162),
.A2(n_169),
.B(n_119),
.C(n_26),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_SL g165 ( 
.A(n_122),
.B(n_131),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_130),
.B(n_137),
.C(n_124),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_166),
.B(n_119),
.C(n_105),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_127),
.B(n_100),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_167),
.B(n_170),
.Y(n_193)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_136),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_168),
.Y(n_185)
);

CKINVDCx16_ASAP7_75t_R g170 ( 
.A(n_120),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_150),
.B(n_137),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g209 ( 
.A(n_171),
.B(n_174),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_166),
.B(n_121),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_155),
.B(n_128),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_175),
.B(n_181),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_170),
.A2(n_120),
.B1(n_138),
.B2(n_135),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_176),
.A2(n_180),
.B1(n_190),
.B2(n_191),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_164),
.A2(n_134),
.B1(n_129),
.B2(n_127),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_154),
.B(n_136),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_182),
.B(n_187),
.C(n_195),
.Y(n_210)
);

FAx1_ASAP7_75t_SL g186 ( 
.A(n_148),
.B(n_26),
.CI(n_13),
.CON(n_186),
.SN(n_186)
);

OR2x2_ASAP7_75t_L g211 ( 
.A(n_186),
.B(n_169),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_163),
.B(n_119),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_189),
.B(n_146),
.Y(n_207)
);

XNOR2x1_ASAP7_75t_L g194 ( 
.A(n_164),
.B(n_26),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_194),
.B(n_162),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_161),
.B(n_32),
.C(n_28),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_177),
.A2(n_160),
.B1(n_156),
.B2(n_159),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_196),
.A2(n_145),
.B1(n_186),
.B2(n_157),
.Y(n_228)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_184),
.Y(n_197)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_197),
.Y(n_225)
);

CKINVDCx16_ASAP7_75t_R g198 ( 
.A(n_188),
.Y(n_198)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_198),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_173),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_199),
.Y(n_232)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_200),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_193),
.Y(n_201)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_201),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_178),
.B(n_165),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g216 ( 
.A1(n_202),
.A2(n_205),
.B1(n_207),
.B2(n_211),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_192),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_SL g230 ( 
.A1(n_204),
.A2(n_206),
.B(n_208),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_183),
.B(n_144),
.Y(n_205)
);

INVxp67_ASAP7_75t_L g206 ( 
.A(n_195),
.Y(n_206)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_187),
.Y(n_208)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_189),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_L g218 ( 
.A1(n_213),
.A2(n_215),
.B1(n_153),
.B2(n_172),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_179),
.B(n_160),
.C(n_163),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_214),
.B(n_182),
.C(n_179),
.Y(n_220)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_177),
.Y(n_215)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_218),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_203),
.A2(n_181),
.B1(n_171),
.B2(n_149),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_219),
.A2(n_224),
.B1(n_229),
.B2(n_211),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_220),
.B(n_222),
.C(n_223),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_214),
.B(n_175),
.C(n_174),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_210),
.B(n_191),
.C(n_185),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_215),
.A2(n_149),
.B1(n_190),
.B2(n_153),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_210),
.B(n_152),
.C(n_151),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_SL g234 ( 
.A(n_227),
.B(n_231),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_228),
.A2(n_207),
.B1(n_197),
.B2(n_208),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_213),
.A2(n_186),
.B1(n_158),
.B2(n_194),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_212),
.B(n_168),
.C(n_32),
.Y(n_231)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_216),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_235),
.B(n_239),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_236),
.A2(n_242),
.B1(n_245),
.B2(n_246),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_238),
.A2(n_23),
.B1(n_13),
.B2(n_19),
.Y(n_257)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_224),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_222),
.B(n_212),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_240),
.B(n_26),
.Y(n_256)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_217),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_241),
.B(n_243),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_L g242 ( 
.A1(n_226),
.A2(n_196),
.B1(n_204),
.B2(n_206),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_225),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_220),
.B(n_209),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_244),
.B(n_240),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_229),
.A2(n_223),
.B1(n_219),
.B2(n_225),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_L g246 ( 
.A1(n_232),
.A2(n_209),
.B1(n_28),
.B2(n_23),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_249),
.B(n_251),
.Y(n_260)
);

AND2x2_ASAP7_75t_L g250 ( 
.A(n_238),
.B(n_221),
.Y(n_250)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_250),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_244),
.B(n_227),
.Y(n_251)
);

AOI21xp5_ASAP7_75t_L g252 ( 
.A1(n_234),
.A2(n_230),
.B(n_228),
.Y(n_252)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_252),
.Y(n_267)
);

OAI21xp5_ASAP7_75t_L g254 ( 
.A1(n_237),
.A2(n_230),
.B(n_231),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_254),
.B(n_256),
.Y(n_259)
);

NAND3xp33_ASAP7_75t_L g255 ( 
.A(n_233),
.B(n_0),
.C(n_1),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_255),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_257),
.B(n_239),
.Y(n_261)
);

MAJx2_ASAP7_75t_L g258 ( 
.A(n_245),
.B(n_13),
.C(n_23),
.Y(n_258)
);

OAI21xp5_ASAP7_75t_L g269 ( 
.A1(n_258),
.A2(n_32),
.B(n_19),
.Y(n_269)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_261),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_250),
.A2(n_236),
.B1(n_237),
.B2(n_3),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_263),
.B(n_2),
.Y(n_273)
);

AOI221xp5_ASAP7_75t_L g264 ( 
.A1(n_248),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.C(n_4),
.Y(n_264)
);

OAI21x1_ASAP7_75t_L g277 ( 
.A1(n_264),
.A2(n_3),
.B(n_6),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_253),
.A2(n_23),
.B1(n_19),
.B2(n_13),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_266),
.A2(n_10),
.B1(n_5),
.B2(n_6),
.Y(n_275)
);

AO221x1_ASAP7_75t_L g268 ( 
.A1(n_255),
.A2(n_19),
.B1(n_32),
.B2(n_5),
.C(n_6),
.Y(n_268)
);

AOI21xp5_ASAP7_75t_L g276 ( 
.A1(n_268),
.A2(n_3),
.B(n_6),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_269),
.B(n_247),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_270),
.B(n_272),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_262),
.B(n_256),
.Y(n_271)
);

AOI21xp5_ASAP7_75t_L g280 ( 
.A1(n_271),
.A2(n_263),
.B(n_259),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_260),
.B(n_258),
.C(n_32),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_273),
.B(n_275),
.Y(n_279)
);

OAI21x1_ASAP7_75t_L g278 ( 
.A1(n_276),
.A2(n_277),
.B(n_264),
.Y(n_278)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_278),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_L g284 ( 
.A1(n_280),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_284)
);

AOI21xp5_ASAP7_75t_L g282 ( 
.A1(n_271),
.A2(n_267),
.B(n_265),
.Y(n_282)
);

OAI21xp5_ASAP7_75t_L g283 ( 
.A1(n_282),
.A2(n_274),
.B(n_269),
.Y(n_283)
);

NOR2x1_ASAP7_75t_L g286 ( 
.A(n_283),
.B(n_284),
.Y(n_286)
);

AOI21xp5_ASAP7_75t_L g287 ( 
.A1(n_286),
.A2(n_285),
.B(n_281),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_287),
.B(n_279),
.C(n_8),
.Y(n_288)
);

OAI21xp5_ASAP7_75t_SL g289 ( 
.A1(n_288),
.A2(n_7),
.B(n_8),
.Y(n_289)
);

A2O1A1O1Ixp25_ASAP7_75t_L g290 ( 
.A1(n_289),
.A2(n_7),
.B(n_8),
.C(n_9),
.D(n_10),
.Y(n_290)
);

AOI21xp5_ASAP7_75t_L g291 ( 
.A1(n_290),
.A2(n_7),
.B(n_9),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_291),
.B(n_10),
.Y(n_292)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_292),
.B(n_10),
.Y(n_293)
);


endmodule