module fake_netlist_6_2939_n_809 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_166, n_28, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_127, n_125, n_153, n_168, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_165, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_159, n_157, n_162, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_809);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_127;
input n_125;
input n_153;
input n_168;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_165;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_809;

wire n_591;
wire n_435;
wire n_793;
wire n_326;
wire n_801;
wire n_256;
wire n_440;
wire n_587;
wire n_695;
wire n_507;
wire n_580;
wire n_762;
wire n_209;
wire n_367;
wire n_465;
wire n_680;
wire n_741;
wire n_760;
wire n_590;
wire n_625;
wire n_661;
wire n_223;
wire n_278;
wire n_362;
wire n_341;
wire n_226;
wire n_208;
wire n_462;
wire n_607;
wire n_671;
wire n_726;
wire n_316;
wire n_419;
wire n_304;
wire n_212;
wire n_700;
wire n_694;
wire n_740;
wire n_578;
wire n_703;
wire n_365;
wire n_384;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_342;
wire n_783;
wire n_725;
wire n_358;
wire n_751;
wire n_449;
wire n_749;
wire n_798;
wire n_188;
wire n_310;
wire n_509;
wire n_186;
wire n_245;
wire n_368;
wire n_575;
wire n_677;
wire n_805;
wire n_396;
wire n_495;
wire n_350;
wire n_585;
wire n_732;
wire n_568;
wire n_392;
wire n_442;
wire n_480;
wire n_724;
wire n_382;
wire n_673;
wire n_180;
wire n_628;
wire n_557;
wire n_349;
wire n_643;
wire n_233;
wire n_617;
wire n_698;
wire n_255;
wire n_807;
wire n_739;
wire n_284;
wire n_400;
wire n_337;
wire n_214;
wire n_485;
wire n_443;
wire n_246;
wire n_768;
wire n_471;
wire n_289;
wire n_421;
wire n_781;
wire n_424;
wire n_789;
wire n_615;
wire n_181;
wire n_182;
wire n_238;
wire n_573;
wire n_769;
wire n_202;
wire n_320;
wire n_639;
wire n_676;
wire n_327;
wire n_794;
wire n_727;
wire n_369;
wire n_597;
wire n_685;
wire n_280;
wire n_287;
wire n_353;
wire n_610;
wire n_555;
wire n_389;
wire n_415;
wire n_230;
wire n_605;
wire n_461;
wire n_383;
wire n_669;
wire n_200;
wire n_447;
wire n_176;
wire n_198;
wire n_300;
wire n_222;
wire n_179;
wire n_248;
wire n_517;
wire n_718;
wire n_747;
wire n_667;
wire n_229;
wire n_542;
wire n_644;
wire n_682;
wire n_621;
wire n_305;
wire n_721;
wire n_750;
wire n_532;
wire n_742;
wire n_173;
wire n_535;
wire n_691;
wire n_250;
wire n_372;
wire n_468;
wire n_544;
wire n_504;
wire n_314;
wire n_378;
wire n_413;
wire n_377;
wire n_791;
wire n_183;
wire n_510;
wire n_375;
wire n_601;
wire n_338;
wire n_522;
wire n_466;
wire n_704;
wire n_748;
wire n_506;
wire n_763;
wire n_360;
wire n_603;
wire n_235;
wire n_536;
wire n_622;
wire n_191;
wire n_340;
wire n_710;
wire n_387;
wire n_452;
wire n_616;
wire n_658;
wire n_744;
wire n_344;
wire n_581;
wire n_428;
wire n_761;
wire n_785;
wire n_746;
wire n_609;
wire n_765;
wire n_432;
wire n_641;
wire n_693;
wire n_631;
wire n_174;
wire n_516;
wire n_758;
wire n_525;
wire n_720;
wire n_611;
wire n_491;
wire n_656;
wire n_772;
wire n_797;
wire n_666;
wire n_371;
wire n_795;
wire n_770;
wire n_567;
wire n_189;
wire n_738;
wire n_405;
wire n_213;
wire n_538;
wire n_294;
wire n_302;
wire n_499;
wire n_380;
wire n_705;
wire n_647;
wire n_197;
wire n_343;
wire n_448;
wire n_494;
wire n_539;
wire n_493;
wire n_397;
wire n_614;
wire n_529;
wire n_445;
wire n_425;
wire n_684;
wire n_454;
wire n_218;
wire n_638;
wire n_234;
wire n_486;
wire n_381;
wire n_236;
wire n_653;
wire n_752;
wire n_172;
wire n_713;
wire n_648;
wire n_657;
wire n_576;
wire n_472;
wire n_270;
wire n_239;
wire n_414;
wire n_563;
wire n_782;
wire n_490;
wire n_803;
wire n_290;
wire n_220;
wire n_224;
wire n_734;
wire n_708;
wire n_196;
wire n_402;
wire n_352;
wire n_668;
wire n_478;
wire n_626;
wire n_574;
wire n_779;
wire n_800;
wire n_460;
wire n_417;
wire n_446;
wire n_498;
wire n_662;
wire n_374;
wire n_659;
wire n_709;
wire n_366;
wire n_777;
wire n_407;
wire n_450;
wire n_808;
wire n_272;
wire n_526;
wire n_185;
wire n_712;
wire n_348;
wire n_711;
wire n_579;
wire n_376;
wire n_390;
wire n_473;
wire n_293;
wire n_334;
wire n_559;
wire n_370;
wire n_458;
wire n_232;
wire n_650;
wire n_717;
wire n_330;
wire n_771;
wire n_470;
wire n_475;
wire n_298;
wire n_492;
wire n_281;
wire n_258;
wire n_551;
wire n_699;
wire n_456;
wire n_564;
wire n_265;
wire n_260;
wire n_313;
wire n_451;
wire n_624;
wire n_279;
wire n_686;
wire n_796;
wire n_252;
wire n_757;
wire n_228;
wire n_565;
wire n_594;
wire n_719;
wire n_356;
wire n_577;
wire n_184;
wire n_552;
wire n_619;
wire n_216;
wire n_455;
wire n_521;
wire n_363;
wire n_572;
wire n_395;
wire n_592;
wire n_745;
wire n_654;
wire n_323;
wire n_606;
wire n_393;
wire n_411;
wire n_503;
wire n_716;
wire n_623;
wire n_599;
wire n_513;
wire n_776;
wire n_321;
wire n_645;
wire n_331;
wire n_227;
wire n_570;
wire n_731;
wire n_406;
wire n_483;
wire n_735;
wire n_204;
wire n_482;
wire n_755;
wire n_474;
wire n_527;
wire n_261;
wire n_683;
wire n_620;
wire n_420;
wire n_608;
wire n_630;
wire n_312;
wire n_394;
wire n_519;
wire n_541;
wire n_512;
wire n_292;
wire n_307;
wire n_469;
wire n_433;
wire n_500;
wire n_792;
wire n_476;
wire n_714;
wire n_291;
wire n_219;
wire n_543;
wire n_357;
wire n_264;
wire n_263;
wire n_589;
wire n_481;
wire n_788;
wire n_325;
wire n_767;
wire n_804;
wire n_329;
wire n_464;
wire n_600;
wire n_802;
wire n_561;
wire n_477;
wire n_549;
wire n_533;
wire n_408;
wire n_806;
wire n_237;
wire n_584;
wire n_244;
wire n_399;
wire n_243;
wire n_548;
wire n_282;
wire n_436;
wire n_211;
wire n_523;
wire n_175;
wire n_322;
wire n_707;
wire n_345;
wire n_409;
wire n_231;
wire n_354;
wire n_689;
wire n_799;
wire n_505;
wire n_240;
wire n_756;
wire n_319;
wire n_547;
wire n_537;
wire n_273;
wire n_558;
wire n_635;
wire n_787;
wire n_311;
wire n_403;
wire n_723;
wire n_253;
wire n_634;
wire n_583;
wire n_596;
wire n_546;
wire n_562;
wire n_249;
wire n_201;
wire n_386;
wire n_764;
wire n_556;
wire n_692;
wire n_733;
wire n_754;
wire n_487;
wire n_550;
wire n_241;
wire n_275;
wire n_553;
wire n_652;
wire n_560;
wire n_753;
wire n_642;
wire n_276;
wire n_569;
wire n_441;
wire n_221;
wire n_444;
wire n_586;
wire n_423;
wire n_737;
wire n_318;
wire n_303;
wire n_511;
wire n_715;
wire n_467;
wire n_306;
wire n_193;
wire n_269;
wire n_359;
wire n_346;
wire n_416;
wire n_530;
wire n_277;
wire n_520;
wire n_418;
wire n_618;
wire n_790;
wire n_582;
wire n_199;
wire n_266;
wire n_296;
wire n_674;
wire n_775;
wire n_571;
wire n_268;
wire n_271;
wire n_404;
wire n_651;
wire n_439;
wire n_217;
wire n_210;
wire n_299;
wire n_518;
wire n_206;
wire n_679;
wire n_453;
wire n_612;
wire n_633;
wire n_665;
wire n_333;
wire n_588;
wire n_215;
wire n_178;
wire n_247;
wire n_225;
wire n_308;
wire n_309;
wire n_759;
wire n_355;
wire n_426;
wire n_317;
wire n_632;
wire n_702;
wire n_431;
wire n_347;
wire n_459;
wire n_502;
wire n_328;
wire n_672;
wire n_534;
wire n_488;
wire n_429;
wire n_373;
wire n_195;
wire n_285;
wire n_497;
wire n_780;
wire n_773;
wire n_675;
wire n_257;
wire n_730;
wire n_655;
wire n_706;
wire n_786;
wire n_670;
wire n_203;
wire n_286;
wire n_254;
wire n_207;
wire n_242;
wire n_690;
wire n_401;
wire n_324;
wire n_743;
wire n_766;
wire n_335;
wire n_430;
wire n_463;
wire n_545;
wire n_489;
wire n_205;
wire n_604;
wire n_251;
wire n_301;
wire n_274;
wire n_636;
wire n_728;
wire n_681;
wire n_729;
wire n_774;
wire n_412;
wire n_640;
wire n_660;
wire n_267;
wire n_438;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_515;
wire n_288;
wire n_427;
wire n_479;
wire n_496;
wire n_598;
wire n_422;
wire n_696;
wire n_688;
wire n_722;
wire n_351;
wire n_437;
wire n_259;
wire n_177;
wire n_540;
wire n_593;
wire n_514;
wire n_646;
wire n_528;
wire n_391;
wire n_457;
wire n_697;
wire n_687;
wire n_364;
wire n_637;
wire n_295;
wire n_385;
wire n_701;
wire n_629;
wire n_388;
wire n_190;
wire n_262;
wire n_484;
wire n_736;
wire n_613;
wire n_187;
wire n_501;
wire n_531;
wire n_361;
wire n_508;
wire n_663;
wire n_379;
wire n_170;
wire n_778;
wire n_332;
wire n_336;
wire n_398;
wire n_410;
wire n_566;
wire n_554;
wire n_602;
wire n_194;
wire n_664;
wire n_171;
wire n_678;
wire n_192;
wire n_169;
wire n_649;
wire n_283;

INVx1_ASAP7_75t_L g169 ( 
.A(n_63),
.Y(n_169)
);

BUFx10_ASAP7_75t_L g170 ( 
.A(n_152),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_88),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_76),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_84),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_5),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_111),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_42),
.Y(n_176)
);

BUFx2_ASAP7_75t_L g177 ( 
.A(n_52),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_97),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_93),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_9),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_12),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_165),
.Y(n_182)
);

INVxp67_ASAP7_75t_SL g183 ( 
.A(n_151),
.Y(n_183)
);

BUFx3_ASAP7_75t_L g184 ( 
.A(n_30),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_119),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_64),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_43),
.Y(n_187)
);

INVx2_ASAP7_75t_SL g188 ( 
.A(n_44),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_37),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_46),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_127),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_102),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_100),
.Y(n_193)
);

INVxp67_ASAP7_75t_SL g194 ( 
.A(n_69),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_135),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_24),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_117),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_55),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_133),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_161),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_159),
.Y(n_201)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_85),
.Y(n_202)
);

INVx1_ASAP7_75t_SL g203 ( 
.A(n_96),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_146),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_81),
.Y(n_205)
);

BUFx6f_ASAP7_75t_L g206 ( 
.A(n_34),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_80),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_137),
.Y(n_208)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_106),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_10),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_0),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_17),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_107),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_125),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_54),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_116),
.Y(n_216)
);

CKINVDCx16_ASAP7_75t_R g217 ( 
.A(n_19),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_101),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_167),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_105),
.Y(n_220)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_50),
.Y(n_221)
);

INVx2_ASAP7_75t_SL g222 ( 
.A(n_75),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_60),
.Y(n_223)
);

HB1xp67_ASAP7_75t_L g224 ( 
.A(n_67),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_14),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_163),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_110),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_72),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_138),
.Y(n_229)
);

HB1xp67_ASAP7_75t_L g230 ( 
.A(n_61),
.Y(n_230)
);

INVx2_ASAP7_75t_SL g231 ( 
.A(n_156),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_166),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_32),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_6),
.Y(n_234)
);

AND2x4_ASAP7_75t_L g235 ( 
.A(n_184),
.B(n_18),
.Y(n_235)
);

AND2x2_ASAP7_75t_L g236 ( 
.A(n_177),
.B(n_0),
.Y(n_236)
);

INVxp67_ASAP7_75t_L g237 ( 
.A(n_174),
.Y(n_237)
);

INVxp67_ASAP7_75t_L g238 ( 
.A(n_180),
.Y(n_238)
);

BUFx6f_ASAP7_75t_L g239 ( 
.A(n_206),
.Y(n_239)
);

BUFx12f_ASAP7_75t_L g240 ( 
.A(n_170),
.Y(n_240)
);

AND2x4_ASAP7_75t_L g241 ( 
.A(n_184),
.B(n_202),
.Y(n_241)
);

HB1xp67_ASAP7_75t_L g242 ( 
.A(n_181),
.Y(n_242)
);

AND2x4_ASAP7_75t_L g243 ( 
.A(n_202),
.B(n_20),
.Y(n_243)
);

AND2x4_ASAP7_75t_L g244 ( 
.A(n_209),
.B(n_21),
.Y(n_244)
);

BUFx6f_ASAP7_75t_L g245 ( 
.A(n_206),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_172),
.Y(n_246)
);

AND2x2_ASAP7_75t_L g247 ( 
.A(n_217),
.B(n_1),
.Y(n_247)
);

AND2x4_ASAP7_75t_L g248 ( 
.A(n_209),
.B(n_22),
.Y(n_248)
);

AND2x2_ASAP7_75t_L g249 ( 
.A(n_224),
.B(n_1),
.Y(n_249)
);

AND2x2_ASAP7_75t_L g250 ( 
.A(n_230),
.B(n_170),
.Y(n_250)
);

INVx3_ASAP7_75t_L g251 ( 
.A(n_170),
.Y(n_251)
);

INVx3_ASAP7_75t_L g252 ( 
.A(n_210),
.Y(n_252)
);

BUFx12f_ASAP7_75t_L g253 ( 
.A(n_178),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_211),
.Y(n_254)
);

BUFx3_ASAP7_75t_L g255 ( 
.A(n_169),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_225),
.Y(n_256)
);

BUFx3_ASAP7_75t_L g257 ( 
.A(n_171),
.Y(n_257)
);

BUFx6f_ASAP7_75t_L g258 ( 
.A(n_206),
.Y(n_258)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_234),
.Y(n_259)
);

AND2x4_ASAP7_75t_L g260 ( 
.A(n_221),
.B(n_23),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_173),
.Y(n_261)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_206),
.Y(n_262)
);

OAI22x1_ASAP7_75t_R g263 ( 
.A1(n_185),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_263)
);

BUFx8_ASAP7_75t_SL g264 ( 
.A(n_185),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_175),
.Y(n_265)
);

AND2x4_ASAP7_75t_L g266 ( 
.A(n_221),
.B(n_25),
.Y(n_266)
);

BUFx6f_ASAP7_75t_L g267 ( 
.A(n_176),
.Y(n_267)
);

BUFx3_ASAP7_75t_L g268 ( 
.A(n_179),
.Y(n_268)
);

HB1xp67_ASAP7_75t_L g269 ( 
.A(n_190),
.Y(n_269)
);

BUFx6f_ASAP7_75t_L g270 ( 
.A(n_193),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_233),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_271)
);

HB1xp67_ASAP7_75t_L g272 ( 
.A(n_199),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_200),
.Y(n_273)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_201),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_213),
.Y(n_275)
);

BUFx6f_ASAP7_75t_L g276 ( 
.A(n_223),
.Y(n_276)
);

INVx4_ASAP7_75t_L g277 ( 
.A(n_178),
.Y(n_277)
);

INVx6_ASAP7_75t_L g278 ( 
.A(n_204),
.Y(n_278)
);

BUFx6f_ASAP7_75t_L g279 ( 
.A(n_229),
.Y(n_279)
);

AND2x6_ASAP7_75t_L g280 ( 
.A(n_232),
.B(n_26),
.Y(n_280)
);

OAI21x1_ASAP7_75t_L g281 ( 
.A1(n_183),
.A2(n_87),
.B(n_164),
.Y(n_281)
);

BUFx8_ASAP7_75t_SL g282 ( 
.A(n_233),
.Y(n_282)
);

INVxp67_ASAP7_75t_L g283 ( 
.A(n_188),
.Y(n_283)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_262),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_274),
.Y(n_285)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_239),
.Y(n_286)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_239),
.Y(n_287)
);

INVx2_ASAP7_75t_L g288 ( 
.A(n_239),
.Y(n_288)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_262),
.Y(n_289)
);

AO21x2_ASAP7_75t_L g290 ( 
.A1(n_243),
.A2(n_194),
.B(n_222),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_SL g291 ( 
.A(n_247),
.B(n_243),
.Y(n_291)
);

AOI21x1_ASAP7_75t_L g292 ( 
.A1(n_243),
.A2(n_231),
.B(n_186),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_274),
.Y(n_293)
);

AND2x2_ASAP7_75t_L g294 ( 
.A(n_250),
.B(n_203),
.Y(n_294)
);

BUFx10_ASAP7_75t_L g295 ( 
.A(n_246),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_261),
.Y(n_296)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_239),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_244),
.B(n_204),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_264),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_277),
.B(n_228),
.Y(n_300)
);

BUFx10_ASAP7_75t_L g301 ( 
.A(n_278),
.Y(n_301)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_245),
.Y(n_302)
);

OR2x6_ASAP7_75t_L g303 ( 
.A(n_240),
.B(n_253),
.Y(n_303)
);

INVx3_ASAP7_75t_L g304 ( 
.A(n_245),
.Y(n_304)
);

INVx2_ASAP7_75t_SL g305 ( 
.A(n_278),
.Y(n_305)
);

INVx2_ASAP7_75t_L g306 ( 
.A(n_258),
.Y(n_306)
);

OAI22xp33_ASAP7_75t_SL g307 ( 
.A1(n_251),
.A2(n_226),
.B1(n_227),
.B2(n_220),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_244),
.B(n_226),
.Y(n_308)
);

AND2x2_ASAP7_75t_L g309 ( 
.A(n_251),
.B(n_182),
.Y(n_309)
);

AND2x6_ASAP7_75t_L g310 ( 
.A(n_244),
.B(n_27),
.Y(n_310)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_258),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_265),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_SL g313 ( 
.A(n_248),
.B(n_187),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_273),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_SL g315 ( 
.A(n_248),
.B(n_189),
.Y(n_315)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_258),
.Y(n_316)
);

NAND2xp33_ASAP7_75t_SL g317 ( 
.A(n_236),
.B(n_191),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_283),
.B(n_249),
.Y(n_318)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_258),
.Y(n_319)
);

OR2x6_ASAP7_75t_L g320 ( 
.A(n_240),
.B(n_5),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_277),
.B(n_248),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_275),
.Y(n_322)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_267),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_SL g324 ( 
.A(n_260),
.B(n_192),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_267),
.Y(n_325)
);

AND2x4_ASAP7_75t_L g326 ( 
.A(n_235),
.B(n_195),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_270),
.Y(n_327)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_270),
.Y(n_328)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_270),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_260),
.B(n_196),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_270),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_291),
.B(n_260),
.Y(n_332)
);

BUFx6f_ASAP7_75t_L g333 ( 
.A(n_304),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_291),
.B(n_266),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_321),
.B(n_266),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_SL g336 ( 
.A(n_294),
.B(n_253),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_321),
.B(n_266),
.Y(n_337)
);

OR2x2_ASAP7_75t_L g338 ( 
.A(n_318),
.B(n_241),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_SL g339 ( 
.A(n_307),
.B(n_235),
.Y(n_339)
);

INVx2_ASAP7_75t_L g340 ( 
.A(n_304),
.Y(n_340)
);

NOR3xp33_ASAP7_75t_L g341 ( 
.A(n_298),
.B(n_271),
.C(n_238),
.Y(n_341)
);

NAND3xp33_ASAP7_75t_L g342 ( 
.A(n_318),
.B(n_272),
.C(n_269),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_309),
.B(n_235),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_296),
.Y(n_344)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_297),
.Y(n_345)
);

INVxp67_ASAP7_75t_L g346 ( 
.A(n_312),
.Y(n_346)
);

NAND3xp33_ASAP7_75t_L g347 ( 
.A(n_298),
.B(n_272),
.C(n_269),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_326),
.B(n_278),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_314),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_326),
.B(n_241),
.Y(n_350)
);

INVx2_ASAP7_75t_SL g351 ( 
.A(n_295),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_330),
.B(n_280),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_300),
.B(n_255),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_322),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_330),
.B(n_313),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_SL g356 ( 
.A(n_295),
.B(n_197),
.Y(n_356)
);

OR2x2_ASAP7_75t_L g357 ( 
.A(n_308),
.B(n_305),
.Y(n_357)
);

NAND2xp33_ASAP7_75t_L g358 ( 
.A(n_310),
.B(n_280),
.Y(n_358)
);

INVxp67_ASAP7_75t_L g359 ( 
.A(n_317),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_313),
.B(n_280),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_315),
.B(n_280),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_315),
.B(n_280),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_324),
.B(n_276),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_L g364 ( 
.A(n_308),
.B(n_255),
.Y(n_364)
);

AOI22xp5_ASAP7_75t_L g365 ( 
.A1(n_317),
.A2(n_198),
.B1(n_205),
.B2(n_207),
.Y(n_365)
);

NAND2xp33_ASAP7_75t_L g366 ( 
.A(n_310),
.B(n_208),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_324),
.B(n_276),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_SL g368 ( 
.A(n_301),
.B(n_212),
.Y(n_368)
);

NOR2xp67_ASAP7_75t_L g369 ( 
.A(n_285),
.B(n_237),
.Y(n_369)
);

INVxp33_ASAP7_75t_L g370 ( 
.A(n_293),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_299),
.Y(n_371)
);

BUFx6f_ASAP7_75t_SL g372 ( 
.A(n_303),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_SL g373 ( 
.A(n_301),
.B(n_214),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_290),
.B(n_276),
.Y(n_374)
);

HB1xp67_ASAP7_75t_L g375 ( 
.A(n_320),
.Y(n_375)
);

NOR3xp33_ASAP7_75t_L g376 ( 
.A(n_292),
.B(n_242),
.C(n_256),
.Y(n_376)
);

BUFx6f_ASAP7_75t_L g377 ( 
.A(n_286),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_290),
.B(n_276),
.Y(n_378)
);

AOI22xp5_ASAP7_75t_L g379 ( 
.A1(n_310),
.A2(n_215),
.B1(n_216),
.B2(n_218),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_L g380 ( 
.A(n_325),
.B(n_257),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_327),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_284),
.B(n_289),
.Y(n_382)
);

AND2x2_ASAP7_75t_L g383 ( 
.A(n_303),
.B(n_257),
.Y(n_383)
);

INVx2_ASAP7_75t_SL g384 ( 
.A(n_320),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_SL g385 ( 
.A(n_323),
.B(n_219),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_SL g386 ( 
.A(n_328),
.B(n_268),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_L g387 ( 
.A(n_331),
.B(n_268),
.Y(n_387)
);

AND2x2_ASAP7_75t_L g388 ( 
.A(n_303),
.B(n_242),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_284),
.B(n_279),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_289),
.B(n_279),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_328),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_332),
.B(n_310),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_344),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_334),
.B(n_310),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_SL g395 ( 
.A(n_355),
.B(n_279),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_334),
.B(n_329),
.Y(n_396)
);

OAI22xp5_ASAP7_75t_L g397 ( 
.A1(n_343),
.A2(n_320),
.B1(n_279),
.B2(n_316),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_335),
.B(n_306),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_349),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_335),
.B(n_337),
.Y(n_400)
);

BUFx6f_ASAP7_75t_L g401 ( 
.A(n_377),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_337),
.B(n_306),
.Y(n_402)
);

A2O1A1Ixp33_ASAP7_75t_L g403 ( 
.A1(n_364),
.A2(n_281),
.B(n_254),
.C(n_252),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_354),
.Y(n_404)
);

AND2x2_ASAP7_75t_L g405 ( 
.A(n_338),
.B(n_252),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_353),
.B(n_316),
.Y(n_406)
);

BUFx6f_ASAP7_75t_L g407 ( 
.A(n_377),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_391),
.Y(n_408)
);

AND2x2_ASAP7_75t_L g409 ( 
.A(n_370),
.B(n_351),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_363),
.B(n_287),
.Y(n_410)
);

AOI21xp5_ASAP7_75t_L g411 ( 
.A1(n_374),
.A2(n_319),
.B(n_311),
.Y(n_411)
);

AOI21xp5_ASAP7_75t_L g412 ( 
.A1(n_360),
.A2(n_302),
.B(n_288),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_R g413 ( 
.A(n_371),
.B(n_28),
.Y(n_413)
);

INVxp33_ASAP7_75t_L g414 ( 
.A(n_388),
.Y(n_414)
);

OAI22xp5_ASAP7_75t_L g415 ( 
.A1(n_359),
.A2(n_259),
.B1(n_263),
.B2(n_264),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_367),
.B(n_259),
.Y(n_416)
);

AOI21xp5_ASAP7_75t_L g417 ( 
.A1(n_361),
.A2(n_90),
.B(n_168),
.Y(n_417)
);

A2O1A1Ixp33_ASAP7_75t_L g418 ( 
.A1(n_362),
.A2(n_6),
.B(n_7),
.C(n_8),
.Y(n_418)
);

NOR2xp33_ASAP7_75t_L g419 ( 
.A(n_357),
.B(n_282),
.Y(n_419)
);

INVx2_ASAP7_75t_L g420 ( 
.A(n_345),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_350),
.Y(n_421)
);

NAND2x1p5_ASAP7_75t_L g422 ( 
.A(n_383),
.B(n_336),
.Y(n_422)
);

AOI21xp5_ASAP7_75t_L g423 ( 
.A1(n_378),
.A2(n_91),
.B(n_162),
.Y(n_423)
);

INVxp67_ASAP7_75t_L g424 ( 
.A(n_342),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_372),
.Y(n_425)
);

AOI21xp5_ASAP7_75t_L g426 ( 
.A1(n_378),
.A2(n_89),
.B(n_160),
.Y(n_426)
);

BUFx6f_ASAP7_75t_L g427 ( 
.A(n_377),
.Y(n_427)
);

OAI21xp5_ASAP7_75t_L g428 ( 
.A1(n_352),
.A2(n_86),
.B(n_158),
.Y(n_428)
);

OAI22xp5_ASAP7_75t_L g429 ( 
.A1(n_379),
.A2(n_282),
.B1(n_83),
.B2(n_92),
.Y(n_429)
);

OAI21xp5_ASAP7_75t_L g430 ( 
.A1(n_358),
.A2(n_79),
.B(n_155),
.Y(n_430)
);

HB1xp67_ASAP7_75t_L g431 ( 
.A(n_348),
.Y(n_431)
);

AOI21xp5_ASAP7_75t_L g432 ( 
.A1(n_366),
.A2(n_78),
.B(n_154),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_382),
.Y(n_433)
);

OAI21xp5_ASAP7_75t_L g434 ( 
.A1(n_339),
.A2(n_77),
.B(n_153),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_376),
.B(n_29),
.Y(n_435)
);

AOI21xp33_ASAP7_75t_L g436 ( 
.A1(n_347),
.A2(n_346),
.B(n_365),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_381),
.B(n_380),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_387),
.B(n_340),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_382),
.Y(n_439)
);

AOI21xp5_ASAP7_75t_L g440 ( 
.A1(n_389),
.A2(n_82),
.B(n_150),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_SL g441 ( 
.A(n_372),
.B(n_7),
.Y(n_441)
);

INVx2_ASAP7_75t_L g442 ( 
.A(n_333),
.Y(n_442)
);

NOR2xp33_ASAP7_75t_L g443 ( 
.A(n_356),
.B(n_8),
.Y(n_443)
);

AOI21xp5_ASAP7_75t_L g444 ( 
.A1(n_389),
.A2(n_94),
.B(n_149),
.Y(n_444)
);

O2A1O1Ixp33_ASAP7_75t_L g445 ( 
.A1(n_386),
.A2(n_9),
.B(n_10),
.C(n_11),
.Y(n_445)
);

BUFx2_ASAP7_75t_SL g446 ( 
.A(n_369),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_390),
.Y(n_447)
);

NOR2xp33_ASAP7_75t_L g448 ( 
.A(n_368),
.B(n_373),
.Y(n_448)
);

NAND2xp33_ASAP7_75t_L g449 ( 
.A(n_341),
.B(n_31),
.Y(n_449)
);

BUFx6f_ASAP7_75t_L g450 ( 
.A(n_333),
.Y(n_450)
);

INVx2_ASAP7_75t_L g451 ( 
.A(n_390),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_385),
.Y(n_452)
);

OR2x6_ASAP7_75t_L g453 ( 
.A(n_384),
.B(n_11),
.Y(n_453)
);

AOI21xp5_ASAP7_75t_L g454 ( 
.A1(n_375),
.A2(n_95),
.B(n_148),
.Y(n_454)
);

O2A1O1Ixp33_ASAP7_75t_L g455 ( 
.A1(n_335),
.A2(n_12),
.B(n_13),
.C(n_14),
.Y(n_455)
);

AO21x2_ASAP7_75t_L g456 ( 
.A1(n_378),
.A2(n_98),
.B(n_147),
.Y(n_456)
);

OAI22x1_ASAP7_75t_L g457 ( 
.A1(n_424),
.A2(n_13),
.B1(n_15),
.B2(n_16),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_393),
.Y(n_458)
);

OAI21x1_ASAP7_75t_L g459 ( 
.A1(n_412),
.A2(n_99),
.B(n_145),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_399),
.Y(n_460)
);

INVx1_ASAP7_75t_SL g461 ( 
.A(n_409),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_404),
.Y(n_462)
);

OAI21xp5_ASAP7_75t_L g463 ( 
.A1(n_400),
.A2(n_74),
.B(n_144),
.Y(n_463)
);

OAI21x1_ASAP7_75t_L g464 ( 
.A1(n_392),
.A2(n_73),
.B(n_143),
.Y(n_464)
);

OAI21x1_ASAP7_75t_L g465 ( 
.A1(n_394),
.A2(n_71),
.B(n_142),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_433),
.B(n_15),
.Y(n_466)
);

INVx2_ASAP7_75t_L g467 ( 
.A(n_420),
.Y(n_467)
);

AOI21xp5_ASAP7_75t_L g468 ( 
.A1(n_396),
.A2(n_70),
.B(n_33),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_439),
.B(n_16),
.Y(n_469)
);

AOI21x1_ASAP7_75t_L g470 ( 
.A1(n_398),
.A2(n_35),
.B(n_36),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_421),
.B(n_38),
.Y(n_471)
);

INVx8_ASAP7_75t_L g472 ( 
.A(n_450),
.Y(n_472)
);

BUFx2_ASAP7_75t_L g473 ( 
.A(n_431),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_447),
.B(n_39),
.Y(n_474)
);

OAI21x1_ASAP7_75t_L g475 ( 
.A1(n_402),
.A2(n_40),
.B(n_41),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_405),
.B(n_45),
.Y(n_476)
);

AOI21xp5_ASAP7_75t_L g477 ( 
.A1(n_410),
.A2(n_47),
.B(n_48),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_451),
.B(n_49),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_437),
.B(n_51),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_416),
.B(n_53),
.Y(n_480)
);

INVx3_ASAP7_75t_L g481 ( 
.A(n_401),
.Y(n_481)
);

AOI21xp5_ASAP7_75t_L g482 ( 
.A1(n_395),
.A2(n_56),
.B(n_57),
.Y(n_482)
);

OAI21xp5_ASAP7_75t_L g483 ( 
.A1(n_403),
.A2(n_58),
.B(n_59),
.Y(n_483)
);

AOI22xp5_ASAP7_75t_L g484 ( 
.A1(n_449),
.A2(n_62),
.B1(n_65),
.B2(n_66),
.Y(n_484)
);

INVx1_ASAP7_75t_SL g485 ( 
.A(n_446),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_408),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_406),
.B(n_68),
.Y(n_487)
);

AOI21xp33_ASAP7_75t_L g488 ( 
.A1(n_443),
.A2(n_103),
.B(n_104),
.Y(n_488)
);

CKINVDCx20_ASAP7_75t_R g489 ( 
.A(n_425),
.Y(n_489)
);

OAI21x1_ASAP7_75t_L g490 ( 
.A1(n_432),
.A2(n_108),
.B(n_109),
.Y(n_490)
);

AND2x2_ASAP7_75t_SL g491 ( 
.A(n_441),
.B(n_112),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_438),
.B(n_113),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_SL g493 ( 
.A(n_436),
.B(n_114),
.Y(n_493)
);

AOI21xp5_ASAP7_75t_L g494 ( 
.A1(n_430),
.A2(n_115),
.B(n_118),
.Y(n_494)
);

AOI21x1_ASAP7_75t_L g495 ( 
.A1(n_435),
.A2(n_120),
.B(n_121),
.Y(n_495)
);

AOI21xp33_ASAP7_75t_L g496 ( 
.A1(n_414),
.A2(n_122),
.B(n_123),
.Y(n_496)
);

AOI21xp5_ASAP7_75t_L g497 ( 
.A1(n_452),
.A2(n_124),
.B(n_126),
.Y(n_497)
);

OAI21x1_ASAP7_75t_SL g498 ( 
.A1(n_434),
.A2(n_428),
.B(n_454),
.Y(n_498)
);

OAI22x1_ASAP7_75t_L g499 ( 
.A1(n_422),
.A2(n_128),
.B1(n_129),
.B2(n_130),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_448),
.B(n_131),
.Y(n_500)
);

AND2x4_ASAP7_75t_L g501 ( 
.A(n_442),
.B(n_132),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_450),
.Y(n_502)
);

NAND2xp33_ASAP7_75t_L g503 ( 
.A(n_450),
.B(n_134),
.Y(n_503)
);

AOI21x1_ASAP7_75t_L g504 ( 
.A1(n_423),
.A2(n_136),
.B(n_139),
.Y(n_504)
);

OAI21x1_ASAP7_75t_L g505 ( 
.A1(n_417),
.A2(n_140),
.B(n_141),
.Y(n_505)
);

OAI21x1_ASAP7_75t_L g506 ( 
.A1(n_426),
.A2(n_157),
.B(n_444),
.Y(n_506)
);

OAI21x1_ASAP7_75t_L g507 ( 
.A1(n_440),
.A2(n_397),
.B(n_429),
.Y(n_507)
);

AOI21xp5_ASAP7_75t_L g508 ( 
.A1(n_401),
.A2(n_407),
.B(n_427),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_401),
.B(n_407),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_466),
.B(n_469),
.Y(n_510)
);

AO21x1_ASAP7_75t_L g511 ( 
.A1(n_483),
.A2(n_494),
.B(n_493),
.Y(n_511)
);

OAI21xp5_ASAP7_75t_L g512 ( 
.A1(n_479),
.A2(n_418),
.B(n_445),
.Y(n_512)
);

INVxp67_ASAP7_75t_L g513 ( 
.A(n_473),
.Y(n_513)
);

CKINVDCx5p33_ASAP7_75t_R g514 ( 
.A(n_489),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_458),
.Y(n_515)
);

INVx2_ASAP7_75t_L g516 ( 
.A(n_467),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_460),
.Y(n_517)
);

NOR2xp33_ASAP7_75t_L g518 ( 
.A(n_461),
.B(n_419),
.Y(n_518)
);

AND2x4_ASAP7_75t_L g519 ( 
.A(n_462),
.B(n_407),
.Y(n_519)
);

HB1xp67_ASAP7_75t_L g520 ( 
.A(n_461),
.Y(n_520)
);

NOR2xp33_ASAP7_75t_L g521 ( 
.A(n_485),
.B(n_415),
.Y(n_521)
);

OAI21x1_ASAP7_75t_L g522 ( 
.A1(n_459),
.A2(n_455),
.B(n_456),
.Y(n_522)
);

NOR2xp33_ASAP7_75t_R g523 ( 
.A(n_485),
.B(n_427),
.Y(n_523)
);

NOR2xp33_ASAP7_75t_L g524 ( 
.A(n_486),
.B(n_453),
.Y(n_524)
);

AO21x2_ASAP7_75t_L g525 ( 
.A1(n_498),
.A2(n_413),
.B(n_453),
.Y(n_525)
);

OAI21x1_ASAP7_75t_L g526 ( 
.A1(n_490),
.A2(n_508),
.B(n_465),
.Y(n_526)
);

NAND2x1p5_ASAP7_75t_L g527 ( 
.A(n_501),
.B(n_481),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_502),
.Y(n_528)
);

OAI21xp5_ASAP7_75t_L g529 ( 
.A1(n_474),
.A2(n_500),
.B(n_471),
.Y(n_529)
);

BUFx2_ASAP7_75t_L g530 ( 
.A(n_472),
.Y(n_530)
);

OAI21x1_ASAP7_75t_L g531 ( 
.A1(n_464),
.A2(n_478),
.B(n_505),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_481),
.B(n_501),
.Y(n_532)
);

OAI21x1_ASAP7_75t_SL g533 ( 
.A1(n_463),
.A2(n_483),
.B(n_476),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_509),
.Y(n_534)
);

OAI21x1_ASAP7_75t_L g535 ( 
.A1(n_504),
.A2(n_475),
.B(n_507),
.Y(n_535)
);

INVx2_ASAP7_75t_L g536 ( 
.A(n_470),
.Y(n_536)
);

OAI21xp5_ASAP7_75t_L g537 ( 
.A1(n_492),
.A2(n_487),
.B(n_480),
.Y(n_537)
);

OAI21x1_ASAP7_75t_L g538 ( 
.A1(n_495),
.A2(n_468),
.B(n_477),
.Y(n_538)
);

OAI21x1_ASAP7_75t_L g539 ( 
.A1(n_497),
.A2(n_482),
.B(n_463),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_491),
.B(n_472),
.Y(n_540)
);

OAI21xp5_ASAP7_75t_L g541 ( 
.A1(n_488),
.A2(n_484),
.B(n_496),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_472),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_499),
.Y(n_543)
);

NOR2xp33_ASAP7_75t_L g544 ( 
.A(n_488),
.B(n_484),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_457),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_503),
.Y(n_546)
);

INVx2_ASAP7_75t_L g547 ( 
.A(n_467),
.Y(n_547)
);

AOI22x1_ASAP7_75t_L g548 ( 
.A1(n_498),
.A2(n_483),
.B1(n_494),
.B2(n_463),
.Y(n_548)
);

INVx1_ASAP7_75t_SL g549 ( 
.A(n_461),
.Y(n_549)
);

INVx2_ASAP7_75t_L g550 ( 
.A(n_467),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_458),
.Y(n_551)
);

AND2x4_ASAP7_75t_L g552 ( 
.A(n_458),
.B(n_460),
.Y(n_552)
);

OAI21x1_ASAP7_75t_L g553 ( 
.A1(n_506),
.A2(n_412),
.B(n_411),
.Y(n_553)
);

AO21x2_ASAP7_75t_L g554 ( 
.A1(n_498),
.A2(n_483),
.B(n_400),
.Y(n_554)
);

AND2x2_ASAP7_75t_L g555 ( 
.A(n_461),
.B(n_294),
.Y(n_555)
);

INVx2_ASAP7_75t_SL g556 ( 
.A(n_461),
.Y(n_556)
);

NAND2x1_ASAP7_75t_L g557 ( 
.A(n_481),
.B(n_401),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_458),
.Y(n_558)
);

OR2x6_ASAP7_75t_L g559 ( 
.A(n_541),
.B(n_544),
.Y(n_559)
);

INVx3_ASAP7_75t_L g560 ( 
.A(n_527),
.Y(n_560)
);

INVx2_ASAP7_75t_L g561 ( 
.A(n_516),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_515),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_547),
.Y(n_563)
);

AO21x1_ASAP7_75t_SL g564 ( 
.A1(n_543),
.A2(n_510),
.B(n_512),
.Y(n_564)
);

CKINVDCx11_ASAP7_75t_R g565 ( 
.A(n_549),
.Y(n_565)
);

INVxp33_ASAP7_75t_L g566 ( 
.A(n_555),
.Y(n_566)
);

HB1xp67_ASAP7_75t_L g567 ( 
.A(n_520),
.Y(n_567)
);

AO21x2_ASAP7_75t_L g568 ( 
.A1(n_533),
.A2(n_544),
.B(n_535),
.Y(n_568)
);

INVxp67_ASAP7_75t_SL g569 ( 
.A(n_520),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_517),
.Y(n_570)
);

INVx2_ASAP7_75t_L g571 ( 
.A(n_547),
.Y(n_571)
);

BUFx2_ASAP7_75t_L g572 ( 
.A(n_513),
.Y(n_572)
);

OAI22xp5_ASAP7_75t_L g573 ( 
.A1(n_548),
.A2(n_527),
.B1(n_532),
.B2(n_540),
.Y(n_573)
);

BUFx2_ASAP7_75t_L g574 ( 
.A(n_513),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_551),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_558),
.Y(n_576)
);

BUFx12f_ASAP7_75t_L g577 ( 
.A(n_514),
.Y(n_577)
);

AOI21x1_ASAP7_75t_L g578 ( 
.A1(n_536),
.A2(n_511),
.B(n_522),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_550),
.Y(n_579)
);

AO21x2_ASAP7_75t_L g580 ( 
.A1(n_537),
.A2(n_529),
.B(n_554),
.Y(n_580)
);

INVx2_ASAP7_75t_L g581 ( 
.A(n_550),
.Y(n_581)
);

AND2x2_ASAP7_75t_L g582 ( 
.A(n_534),
.B(n_552),
.Y(n_582)
);

AND2x2_ASAP7_75t_L g583 ( 
.A(n_552),
.B(n_545),
.Y(n_583)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_552),
.Y(n_584)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_519),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_528),
.Y(n_586)
);

BUFx3_ASAP7_75t_L g587 ( 
.A(n_530),
.Y(n_587)
);

OAI21x1_ASAP7_75t_L g588 ( 
.A1(n_526),
.A2(n_553),
.B(n_531),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_519),
.Y(n_589)
);

BUFx3_ASAP7_75t_L g590 ( 
.A(n_556),
.Y(n_590)
);

INVx2_ASAP7_75t_L g591 ( 
.A(n_554),
.Y(n_591)
);

BUFx6f_ASAP7_75t_L g592 ( 
.A(n_557),
.Y(n_592)
);

INVx2_ASAP7_75t_L g593 ( 
.A(n_538),
.Y(n_593)
);

INVx2_ASAP7_75t_L g594 ( 
.A(n_519),
.Y(n_594)
);

OAI22xp33_ASAP7_75t_L g595 ( 
.A1(n_521),
.A2(n_518),
.B1(n_524),
.B2(n_514),
.Y(n_595)
);

BUFx2_ASAP7_75t_R g596 ( 
.A(n_525),
.Y(n_596)
);

BUFx3_ASAP7_75t_L g597 ( 
.A(n_542),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_L g598 ( 
.A(n_518),
.B(n_521),
.Y(n_598)
);

BUFx3_ASAP7_75t_L g599 ( 
.A(n_525),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_546),
.Y(n_600)
);

BUFx3_ASAP7_75t_L g601 ( 
.A(n_524),
.Y(n_601)
);

BUFx3_ASAP7_75t_L g602 ( 
.A(n_587),
.Y(n_602)
);

AND2x2_ASAP7_75t_L g603 ( 
.A(n_559),
.B(n_539),
.Y(n_603)
);

NOR2xp33_ASAP7_75t_L g604 ( 
.A(n_598),
.B(n_523),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_600),
.Y(n_605)
);

AND2x2_ASAP7_75t_L g606 ( 
.A(n_559),
.B(n_523),
.Y(n_606)
);

AO31x2_ASAP7_75t_L g607 ( 
.A1(n_591),
.A2(n_593),
.A3(n_573),
.B(n_600),
.Y(n_607)
);

INVx2_ASAP7_75t_L g608 ( 
.A(n_561),
.Y(n_608)
);

HB1xp67_ASAP7_75t_L g609 ( 
.A(n_572),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_579),
.Y(n_610)
);

OR2x2_ASAP7_75t_L g611 ( 
.A(n_559),
.B(n_568),
.Y(n_611)
);

BUFx2_ASAP7_75t_L g612 ( 
.A(n_569),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_579),
.Y(n_613)
);

AND2x2_ASAP7_75t_L g614 ( 
.A(n_559),
.B(n_584),
.Y(n_614)
);

INVx2_ASAP7_75t_L g615 ( 
.A(n_561),
.Y(n_615)
);

INVx2_ASAP7_75t_SL g616 ( 
.A(n_590),
.Y(n_616)
);

AND2x2_ASAP7_75t_L g617 ( 
.A(n_559),
.B(n_584),
.Y(n_617)
);

INVx1_ASAP7_75t_SL g618 ( 
.A(n_565),
.Y(n_618)
);

BUFx3_ASAP7_75t_L g619 ( 
.A(n_587),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_562),
.Y(n_620)
);

HB1xp67_ASAP7_75t_L g621 ( 
.A(n_572),
.Y(n_621)
);

INVx2_ASAP7_75t_L g622 ( 
.A(n_563),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_582),
.B(n_566),
.Y(n_623)
);

INVx2_ASAP7_75t_L g624 ( 
.A(n_563),
.Y(n_624)
);

AND2x2_ASAP7_75t_L g625 ( 
.A(n_582),
.B(n_564),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_562),
.Y(n_626)
);

AND2x2_ASAP7_75t_L g627 ( 
.A(n_564),
.B(n_581),
.Y(n_627)
);

AND2x2_ASAP7_75t_L g628 ( 
.A(n_571),
.B(n_581),
.Y(n_628)
);

AND2x2_ASAP7_75t_L g629 ( 
.A(n_571),
.B(n_583),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_570),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_570),
.Y(n_631)
);

NAND3xp33_ASAP7_75t_L g632 ( 
.A(n_595),
.B(n_583),
.C(n_589),
.Y(n_632)
);

INVx2_ASAP7_75t_L g633 ( 
.A(n_575),
.Y(n_633)
);

INVxp67_ASAP7_75t_SL g634 ( 
.A(n_567),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_575),
.Y(n_635)
);

AND2x4_ASAP7_75t_L g636 ( 
.A(n_585),
.B(n_594),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_576),
.Y(n_637)
);

INVx2_ASAP7_75t_L g638 ( 
.A(n_576),
.Y(n_638)
);

HB1xp67_ASAP7_75t_L g639 ( 
.A(n_574),
.Y(n_639)
);

HB1xp67_ASAP7_75t_L g640 ( 
.A(n_574),
.Y(n_640)
);

HB1xp67_ASAP7_75t_L g641 ( 
.A(n_590),
.Y(n_641)
);

INVx2_ASAP7_75t_L g642 ( 
.A(n_586),
.Y(n_642)
);

INVx2_ASAP7_75t_L g643 ( 
.A(n_586),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_589),
.Y(n_644)
);

BUFx2_ASAP7_75t_L g645 ( 
.A(n_590),
.Y(n_645)
);

AND2x2_ASAP7_75t_L g646 ( 
.A(n_585),
.B(n_594),
.Y(n_646)
);

AND2x2_ASAP7_75t_L g647 ( 
.A(n_601),
.B(n_560),
.Y(n_647)
);

AND2x2_ASAP7_75t_L g648 ( 
.A(n_614),
.B(n_568),
.Y(n_648)
);

AND2x2_ASAP7_75t_L g649 ( 
.A(n_614),
.B(n_568),
.Y(n_649)
);

BUFx2_ASAP7_75t_L g650 ( 
.A(n_612),
.Y(n_650)
);

AOI22xp33_ASAP7_75t_L g651 ( 
.A1(n_604),
.A2(n_601),
.B1(n_577),
.B2(n_599),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_626),
.Y(n_652)
);

INVx2_ASAP7_75t_L g653 ( 
.A(n_605),
.Y(n_653)
);

CKINVDCx20_ASAP7_75t_R g654 ( 
.A(n_618),
.Y(n_654)
);

AND2x2_ASAP7_75t_L g655 ( 
.A(n_617),
.B(n_599),
.Y(n_655)
);

AND2x2_ASAP7_75t_L g656 ( 
.A(n_617),
.B(n_599),
.Y(n_656)
);

AND2x2_ASAP7_75t_L g657 ( 
.A(n_629),
.B(n_580),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_605),
.Y(n_658)
);

INVxp67_ASAP7_75t_L g659 ( 
.A(n_609),
.Y(n_659)
);

AND2x2_ASAP7_75t_L g660 ( 
.A(n_629),
.B(n_580),
.Y(n_660)
);

INVx2_ASAP7_75t_SL g661 ( 
.A(n_602),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_L g662 ( 
.A(n_623),
.B(n_601),
.Y(n_662)
);

AND2x2_ASAP7_75t_L g663 ( 
.A(n_625),
.B(n_580),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_621),
.B(n_587),
.Y(n_664)
);

HB1xp67_ASAP7_75t_L g665 ( 
.A(n_612),
.Y(n_665)
);

INVxp67_ASAP7_75t_L g666 ( 
.A(n_639),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_L g667 ( 
.A(n_640),
.B(n_560),
.Y(n_667)
);

INVx2_ASAP7_75t_L g668 ( 
.A(n_633),
.Y(n_668)
);

AND2x2_ASAP7_75t_L g669 ( 
.A(n_625),
.B(n_596),
.Y(n_669)
);

INVx2_ASAP7_75t_SL g670 ( 
.A(n_602),
.Y(n_670)
);

AND2x2_ASAP7_75t_L g671 ( 
.A(n_603),
.B(n_578),
.Y(n_671)
);

INVxp67_ASAP7_75t_L g672 ( 
.A(n_641),
.Y(n_672)
);

AOI22xp33_ASAP7_75t_L g673 ( 
.A1(n_632),
.A2(n_606),
.B1(n_603),
.B2(n_647),
.Y(n_673)
);

INVx2_ASAP7_75t_L g674 ( 
.A(n_633),
.Y(n_674)
);

INVx2_ASAP7_75t_L g675 ( 
.A(n_638),
.Y(n_675)
);

AND2x2_ASAP7_75t_L g676 ( 
.A(n_647),
.B(n_578),
.Y(n_676)
);

OAI22xp5_ASAP7_75t_L g677 ( 
.A1(n_634),
.A2(n_597),
.B1(n_577),
.B2(n_560),
.Y(n_677)
);

BUFx2_ASAP7_75t_L g678 ( 
.A(n_627),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_L g679 ( 
.A(n_646),
.B(n_636),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_626),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_635),
.Y(n_681)
);

AND2x2_ASAP7_75t_L g682 ( 
.A(n_627),
.B(n_593),
.Y(n_682)
);

OR2x2_ASAP7_75t_L g683 ( 
.A(n_611),
.B(n_593),
.Y(n_683)
);

AOI22xp33_ASAP7_75t_L g684 ( 
.A1(n_606),
.A2(n_560),
.B1(n_597),
.B2(n_592),
.Y(n_684)
);

AND2x4_ASAP7_75t_L g685 ( 
.A(n_638),
.B(n_597),
.Y(n_685)
);

NOR2xp67_ASAP7_75t_L g686 ( 
.A(n_616),
.B(n_592),
.Y(n_686)
);

INVx2_ASAP7_75t_L g687 ( 
.A(n_642),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_658),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_658),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_652),
.Y(n_690)
);

OR2x2_ASAP7_75t_L g691 ( 
.A(n_657),
.B(n_611),
.Y(n_691)
);

OR2x2_ASAP7_75t_L g692 ( 
.A(n_657),
.B(n_607),
.Y(n_692)
);

AND2x4_ASAP7_75t_L g693 ( 
.A(n_682),
.B(n_678),
.Y(n_693)
);

HB1xp67_ASAP7_75t_L g694 ( 
.A(n_650),
.Y(n_694)
);

AND2x2_ASAP7_75t_L g695 ( 
.A(n_663),
.B(n_607),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_L g696 ( 
.A(n_662),
.B(n_645),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_659),
.B(n_645),
.Y(n_697)
);

NAND4xp25_ASAP7_75t_L g698 ( 
.A(n_651),
.B(n_631),
.C(n_620),
.D(n_630),
.Y(n_698)
);

AND2x2_ASAP7_75t_L g699 ( 
.A(n_663),
.B(n_607),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_L g700 ( 
.A(n_666),
.B(n_643),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_680),
.Y(n_701)
);

INVx1_ASAP7_75t_SL g702 ( 
.A(n_664),
.Y(n_702)
);

OR2x2_ASAP7_75t_L g703 ( 
.A(n_660),
.B(n_607),
.Y(n_703)
);

AND2x2_ASAP7_75t_L g704 ( 
.A(n_655),
.B(n_616),
.Y(n_704)
);

INVx2_ASAP7_75t_L g705 ( 
.A(n_653),
.Y(n_705)
);

AND2x2_ASAP7_75t_L g706 ( 
.A(n_660),
.B(n_607),
.Y(n_706)
);

AND2x2_ASAP7_75t_L g707 ( 
.A(n_655),
.B(n_656),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_681),
.Y(n_708)
);

NOR2xp33_ASAP7_75t_L g709 ( 
.A(n_677),
.B(n_619),
.Y(n_709)
);

OR2x2_ASAP7_75t_L g710 ( 
.A(n_665),
.B(n_643),
.Y(n_710)
);

AND2x2_ASAP7_75t_L g711 ( 
.A(n_656),
.B(n_619),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_653),
.Y(n_712)
);

HB1xp67_ASAP7_75t_L g713 ( 
.A(n_650),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_668),
.Y(n_714)
);

INVx2_ASAP7_75t_L g715 ( 
.A(n_668),
.Y(n_715)
);

INVx4_ASAP7_75t_L g716 ( 
.A(n_685),
.Y(n_716)
);

INVx2_ASAP7_75t_L g717 ( 
.A(n_674),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_L g718 ( 
.A(n_679),
.B(n_667),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_674),
.Y(n_719)
);

AND2x2_ASAP7_75t_L g720 ( 
.A(n_648),
.B(n_637),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_672),
.B(n_642),
.Y(n_721)
);

INVx1_ASAP7_75t_SL g722 ( 
.A(n_702),
.Y(n_722)
);

INVxp67_ASAP7_75t_L g723 ( 
.A(n_694),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_688),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_L g725 ( 
.A(n_718),
.B(n_673),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_L g726 ( 
.A(n_696),
.B(n_676),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_689),
.Y(n_727)
);

INVx2_ASAP7_75t_L g728 ( 
.A(n_705),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_690),
.Y(n_729)
);

AND2x2_ASAP7_75t_L g730 ( 
.A(n_707),
.B(n_693),
.Y(n_730)
);

AOI33xp33_ASAP7_75t_L g731 ( 
.A1(n_701),
.A2(n_669),
.A3(n_635),
.B1(n_637),
.B2(n_671),
.B3(n_676),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_708),
.Y(n_732)
);

INVx4_ASAP7_75t_L g733 ( 
.A(n_716),
.Y(n_733)
);

INVx2_ASAP7_75t_L g734 ( 
.A(n_705),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_712),
.Y(n_735)
);

AOI21xp33_ASAP7_75t_SL g736 ( 
.A1(n_697),
.A2(n_669),
.B(n_670),
.Y(n_736)
);

AND2x2_ASAP7_75t_L g737 ( 
.A(n_693),
.B(n_678),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_694),
.Y(n_738)
);

INVx2_ASAP7_75t_L g739 ( 
.A(n_715),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_713),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_L g741 ( 
.A(n_700),
.B(n_671),
.Y(n_741)
);

NAND3xp33_ASAP7_75t_L g742 ( 
.A(n_731),
.B(n_698),
.C(n_709),
.Y(n_742)
);

OAI22xp5_ASAP7_75t_L g743 ( 
.A1(n_736),
.A2(n_684),
.B1(n_709),
.B2(n_716),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_724),
.Y(n_744)
);

OAI21xp5_ASAP7_75t_SL g745 ( 
.A1(n_725),
.A2(n_695),
.B(n_699),
.Y(n_745)
);

INVx1_ASAP7_75t_SL g746 ( 
.A(n_722),
.Y(n_746)
);

INVxp67_ASAP7_75t_L g747 ( 
.A(n_738),
.Y(n_747)
);

AND2x2_ASAP7_75t_L g748 ( 
.A(n_730),
.B(n_737),
.Y(n_748)
);

INVx1_ASAP7_75t_SL g749 ( 
.A(n_741),
.Y(n_749)
);

AND2x2_ASAP7_75t_SL g750 ( 
.A(n_731),
.B(n_716),
.Y(n_750)
);

INVx1_ASAP7_75t_SL g751 ( 
.A(n_726),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_L g752 ( 
.A(n_729),
.B(n_732),
.Y(n_752)
);

AND2x2_ASAP7_75t_L g753 ( 
.A(n_740),
.B(n_693),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_727),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_735),
.Y(n_755)
);

AOI22xp5_ASAP7_75t_L g756 ( 
.A1(n_750),
.A2(n_648),
.B1(n_649),
.B2(n_733),
.Y(n_756)
);

OAI221xp5_ASAP7_75t_L g757 ( 
.A1(n_742),
.A2(n_721),
.B1(n_723),
.B2(n_733),
.C(n_691),
.Y(n_757)
);

OAI22xp33_ASAP7_75t_L g758 ( 
.A1(n_745),
.A2(n_692),
.B1(n_703),
.B2(n_723),
.Y(n_758)
);

AOI211xp5_ASAP7_75t_L g759 ( 
.A1(n_743),
.A2(n_713),
.B(n_711),
.C(n_686),
.Y(n_759)
);

XNOR2x1_ASAP7_75t_L g760 ( 
.A(n_746),
.B(n_654),
.Y(n_760)
);

OAI22xp5_ASAP7_75t_L g761 ( 
.A1(n_750),
.A2(n_751),
.B1(n_749),
.B2(n_752),
.Y(n_761)
);

AND2x2_ASAP7_75t_L g762 ( 
.A(n_748),
.B(n_695),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_757),
.B(n_754),
.Y(n_763)
);

NOR2xp33_ASAP7_75t_L g764 ( 
.A(n_760),
.B(n_654),
.Y(n_764)
);

NAND3xp33_ASAP7_75t_SL g765 ( 
.A(n_759),
.B(n_756),
.C(n_761),
.Y(n_765)
);

AOI222xp33_ASAP7_75t_L g766 ( 
.A1(n_758),
.A2(n_747),
.B1(n_744),
.B2(n_755),
.C1(n_699),
.C2(n_706),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_762),
.Y(n_767)
);

NAND4xp25_ASAP7_75t_L g768 ( 
.A(n_759),
.B(n_747),
.C(n_710),
.D(n_704),
.Y(n_768)
);

AOI221xp5_ASAP7_75t_L g769 ( 
.A1(n_765),
.A2(n_753),
.B1(n_728),
.B2(n_734),
.C(n_739),
.Y(n_769)
);

OAI21xp33_ASAP7_75t_L g770 ( 
.A1(n_763),
.A2(n_720),
.B(n_706),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_767),
.Y(n_771)
);

NAND3xp33_ASAP7_75t_L g772 ( 
.A(n_766),
.B(n_670),
.C(n_661),
.Y(n_772)
);

NOR3x1_ASAP7_75t_L g773 ( 
.A(n_768),
.B(n_661),
.C(n_719),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_L g774 ( 
.A(n_771),
.B(n_764),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_769),
.B(n_748),
.Y(n_775)
);

AO22x2_ASAP7_75t_L g776 ( 
.A1(n_772),
.A2(n_734),
.B1(n_728),
.B2(n_739),
.Y(n_776)
);

AOI22x1_ASAP7_75t_L g777 ( 
.A1(n_776),
.A2(n_773),
.B1(n_770),
.B2(n_685),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_774),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_775),
.Y(n_779)
);

CKINVDCx5p33_ASAP7_75t_R g780 ( 
.A(n_778),
.Y(n_780)
);

BUFx3_ASAP7_75t_L g781 ( 
.A(n_779),
.Y(n_781)
);

XOR2xp5_ASAP7_75t_L g782 ( 
.A(n_777),
.B(n_636),
.Y(n_782)
);

HB1xp67_ASAP7_75t_L g783 ( 
.A(n_778),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_778),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_783),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_SL g786 ( 
.A(n_780),
.B(n_685),
.Y(n_786)
);

NOR2xp33_ASAP7_75t_L g787 ( 
.A(n_781),
.B(n_714),
.Y(n_787)
);

AOI22xp5_ASAP7_75t_L g788 ( 
.A1(n_782),
.A2(n_720),
.B1(n_682),
.B2(n_649),
.Y(n_788)
);

AOI22xp5_ASAP7_75t_L g789 ( 
.A1(n_784),
.A2(n_717),
.B1(n_715),
.B2(n_644),
.Y(n_789)
);

XNOR2x1_ASAP7_75t_L g790 ( 
.A(n_783),
.B(n_636),
.Y(n_790)
);

BUFx8_ASAP7_75t_L g791 ( 
.A(n_785),
.Y(n_791)
);

AOI22xp33_ASAP7_75t_L g792 ( 
.A1(n_786),
.A2(n_675),
.B1(n_687),
.B2(n_717),
.Y(n_792)
);

INVx2_ASAP7_75t_L g793 ( 
.A(n_790),
.Y(n_793)
);

AOI22xp5_ASAP7_75t_L g794 ( 
.A1(n_787),
.A2(n_613),
.B1(n_610),
.B2(n_687),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_789),
.Y(n_795)
);

AOI21xp5_ASAP7_75t_L g796 ( 
.A1(n_793),
.A2(n_788),
.B(n_592),
.Y(n_796)
);

OA21x2_ASAP7_75t_L g797 ( 
.A1(n_795),
.A2(n_588),
.B(n_613),
.Y(n_797)
);

AOI21xp5_ASAP7_75t_SL g798 ( 
.A1(n_791),
.A2(n_592),
.B(n_610),
.Y(n_798)
);

AOI21xp33_ASAP7_75t_SL g799 ( 
.A1(n_794),
.A2(n_683),
.B(n_675),
.Y(n_799)
);

INVxp67_ASAP7_75t_SL g800 ( 
.A(n_797),
.Y(n_800)
);

AO22x2_ASAP7_75t_L g801 ( 
.A1(n_796),
.A2(n_792),
.B1(n_615),
.B2(n_622),
.Y(n_801)
);

NOR2x1_ASAP7_75t_L g802 ( 
.A(n_798),
.B(n_592),
.Y(n_802)
);

HB1xp67_ASAP7_75t_L g803 ( 
.A(n_799),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_803),
.Y(n_804)
);

NAND4xp25_ASAP7_75t_L g805 ( 
.A(n_802),
.B(n_646),
.C(n_683),
.D(n_628),
.Y(n_805)
);

NOR2xp67_ASAP7_75t_L g806 ( 
.A(n_804),
.B(n_800),
.Y(n_806)
);

OR2x6_ASAP7_75t_L g807 ( 
.A(n_806),
.B(n_801),
.Y(n_807)
);

OR2x2_ASAP7_75t_L g808 ( 
.A(n_807),
.B(n_805),
.Y(n_808)
);

AOI22xp5_ASAP7_75t_L g809 ( 
.A1(n_808),
.A2(n_628),
.B1(n_608),
.B2(n_624),
.Y(n_809)
);


endmodule