module fake_jpeg_19928_n_78 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_78);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_78;

wire n_10;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_65;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_40;
wire n_71;
wire n_30;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_77;
wire n_61;
wire n_45;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_11;
wire n_56;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_22;
wire n_35;
wire n_48;
wire n_46;
wire n_9;
wire n_36;
wire n_62;
wire n_43;
wire n_32;

INVx1_ASAP7_75t_L g9 ( 
.A(n_0),
.Y(n_9)
);

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_7),
.Y(n_10)
);

INVx8_ASAP7_75t_SL g11 ( 
.A(n_8),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_8),
.Y(n_12)
);

BUFx2_ASAP7_75t_L g13 ( 
.A(n_3),
.Y(n_13)
);

BUFx3_ASAP7_75t_L g14 ( 
.A(n_4),
.Y(n_14)
);

BUFx10_ASAP7_75t_L g15 ( 
.A(n_4),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

INVx3_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_18),
.B(n_19),
.Y(n_28)
);

INVx1_ASAP7_75t_SL g19 ( 
.A(n_9),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

INVx6_ASAP7_75t_L g24 ( 
.A(n_20),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_10),
.B(n_12),
.Y(n_21)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_21),
.Y(n_25)
);

INVxp67_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_22),
.Y(n_29)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_23),
.Y(n_26)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_20),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_27),
.B(n_15),
.Y(n_33)
);

OAI21xp5_ASAP7_75t_L g30 ( 
.A1(n_28),
.A2(n_22),
.B(n_9),
.Y(n_30)
);

XNOR2xp5_ASAP7_75t_L g42 ( 
.A(n_30),
.B(n_38),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_L g31 ( 
.A1(n_24),
.A2(n_23),
.B1(n_18),
.B2(n_19),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_31),
.A2(n_36),
.B1(n_30),
.B2(n_17),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g32 ( 
.A(n_25),
.B(n_12),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_SL g43 ( 
.A(n_32),
.B(n_35),
.Y(n_43)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_33),
.Y(n_45)
);

INVx13_ASAP7_75t_L g34 ( 
.A(n_29),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_34),
.B(n_15),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g35 ( 
.A(n_25),
.B(n_10),
.Y(n_35)
);

AOI22xp5_ASAP7_75t_L g36 ( 
.A1(n_24),
.A2(n_9),
.B1(n_17),
.B2(n_13),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_28),
.B(n_13),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_37),
.B(n_15),
.Y(n_48)
);

AND2x2_ASAP7_75t_L g38 ( 
.A(n_27),
.B(n_15),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_38),
.Y(n_39)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_40),
.B(n_44),
.Y(n_55)
);

OR2x2_ASAP7_75t_L g41 ( 
.A(n_37),
.B(n_29),
.Y(n_41)
);

AOI21xp5_ASAP7_75t_L g51 ( 
.A1(n_41),
.A2(n_47),
.B(n_0),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g56 ( 
.A1(n_46),
.A2(n_48),
.B1(n_1),
.B2(n_2),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_32),
.B(n_15),
.Y(n_47)
);

MAJIxp5_ASAP7_75t_L g49 ( 
.A(n_42),
.B(n_38),
.C(n_31),
.Y(n_49)
);

MAJIxp5_ASAP7_75t_L g57 ( 
.A(n_49),
.B(n_53),
.C(n_56),
.Y(n_57)
);

OAI22xp33_ASAP7_75t_L g50 ( 
.A1(n_45),
.A2(n_36),
.B1(n_26),
.B2(n_16),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_50),
.B(n_51),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_39),
.A2(n_26),
.B1(n_16),
.B2(n_15),
.Y(n_52)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_52),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_48),
.A2(n_16),
.B1(n_14),
.B2(n_3),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_56),
.B(n_43),
.Y(n_58)
);

XNOR2xp5_ASAP7_75t_L g64 ( 
.A(n_58),
.B(n_60),
.Y(n_64)
);

MAJIxp5_ASAP7_75t_L g60 ( 
.A(n_49),
.B(n_42),
.C(n_41),
.Y(n_60)
);

AOI322xp5_ASAP7_75t_SL g62 ( 
.A1(n_52),
.A2(n_46),
.A3(n_7),
.B1(n_6),
.B2(n_5),
.C1(n_4),
.C2(n_2),
.Y(n_62)
);

MAJx2_ASAP7_75t_L g66 ( 
.A(n_62),
.B(n_5),
.C(n_6),
.Y(n_66)
);

BUFx2_ASAP7_75t_L g63 ( 
.A(n_61),
.Y(n_63)
);

A2O1A1Ixp33_ASAP7_75t_SL g68 ( 
.A1(n_63),
.A2(n_65),
.B(n_50),
.C(n_53),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_59),
.Y(n_65)
);

XNOR2xp5_ASAP7_75t_L g69 ( 
.A(n_66),
.B(n_57),
.Y(n_69)
);

AOI21xp5_ASAP7_75t_SL g67 ( 
.A1(n_65),
.A2(n_54),
.B(n_62),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_67),
.B(n_68),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_69),
.B(n_55),
.Y(n_71)
);

XNOR2xp5_ASAP7_75t_SL g70 ( 
.A(n_69),
.B(n_64),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_70),
.B(n_71),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_72),
.B(n_44),
.Y(n_74)
);

BUFx24_ASAP7_75t_SL g75 ( 
.A(n_74),
.Y(n_75)
);

OAI21xp5_ASAP7_75t_SL g76 ( 
.A1(n_75),
.A2(n_73),
.B(n_2),
.Y(n_76)
);

OAI211xp5_ASAP7_75t_L g77 ( 
.A1(n_76),
.A2(n_1),
.B(n_16),
.C(n_14),
.Y(n_77)
);

XNOR2x2_ASAP7_75t_SL g78 ( 
.A(n_77),
.B(n_1),
.Y(n_78)
);


endmodule