module fake_jpeg_27223_n_329 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_329);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_329;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_137;
wire n_74;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx16_ASAP7_75t_R g16 ( 
.A(n_14),
.Y(n_16)
);

BUFx10_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_5),
.Y(n_18)
);

INVx5_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_2),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_11),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_11),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

INVx6_ASAP7_75t_SL g30 ( 
.A(n_7),
.Y(n_30)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_14),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

INVx11_ASAP7_75t_SL g34 ( 
.A(n_6),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_20),
.Y(n_35)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_35),
.Y(n_63)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_34),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_36),
.B(n_38),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_34),
.Y(n_37)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_27),
.Y(n_38)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_20),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_40),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_19),
.Y(n_41)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_30),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_42),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_20),
.B(n_0),
.Y(n_43)
);

AND2x2_ASAP7_75t_L g46 ( 
.A(n_43),
.B(n_33),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_19),
.Y(n_44)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_44),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_19),
.Y(n_45)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_45),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_46),
.B(n_68),
.Y(n_71)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_43),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_50),
.B(n_54),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_35),
.B(n_22),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_51),
.B(n_52),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_40),
.B(n_22),
.Y(n_52)
);

HB1xp67_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_53),
.Y(n_73)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_41),
.B(n_21),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_56),
.B(n_65),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_39),
.A2(n_16),
.B1(n_32),
.B2(n_24),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_58),
.A2(n_70),
.B1(n_16),
.B2(n_25),
.Y(n_75)
);

AND2x2_ASAP7_75t_L g59 ( 
.A(n_41),
.B(n_29),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_59),
.B(n_33),
.Y(n_102)
);

INVx5_ASAP7_75t_L g60 ( 
.A(n_37),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_60),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_36),
.A2(n_31),
.B1(n_30),
.B2(n_28),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_61),
.A2(n_28),
.B1(n_25),
.B2(n_31),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_42),
.B(n_22),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_64),
.B(n_66),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_44),
.B(n_18),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_44),
.B(n_21),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_45),
.B(n_26),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_45),
.A2(n_31),
.B1(n_30),
.B2(n_25),
.Y(n_70)
);

BUFx12f_ASAP7_75t_L g72 ( 
.A(n_60),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_72),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_75),
.A2(n_78),
.B1(n_62),
.B2(n_57),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_76),
.A2(n_98),
.B1(n_70),
.B2(n_57),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_50),
.B(n_26),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_77),
.B(n_80),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_56),
.A2(n_31),
.B1(n_28),
.B2(n_26),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_64),
.B(n_32),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_79),
.B(n_85),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_46),
.B(n_32),
.Y(n_80)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_65),
.Y(n_82)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_82),
.Y(n_110)
);

INVx11_ASAP7_75t_L g83 ( 
.A(n_55),
.Y(n_83)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_83),
.Y(n_134)
);

AOI32xp33_ASAP7_75t_L g84 ( 
.A1(n_51),
.A2(n_24),
.A3(n_23),
.B1(n_27),
.B2(n_33),
.Y(n_84)
);

MAJx2_ASAP7_75t_L g131 ( 
.A(n_84),
.B(n_90),
.C(n_103),
.Y(n_131)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_63),
.Y(n_85)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_63),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_86),
.B(n_91),
.Y(n_126)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_66),
.Y(n_87)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_87),
.Y(n_125)
);

AND2x2_ASAP7_75t_SL g88 ( 
.A(n_46),
.B(n_29),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_88),
.B(n_17),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_48),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_89),
.Y(n_111)
);

OR2x4_ASAP7_75t_L g90 ( 
.A(n_58),
.B(n_17),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_52),
.B(n_24),
.Y(n_91)
);

OR2x2_ASAP7_75t_SL g92 ( 
.A(n_68),
.B(n_21),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_92),
.B(n_93),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_47),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_57),
.A2(n_18),
.B1(n_23),
.B2(n_27),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_94),
.Y(n_109)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_47),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_97),
.B(n_100),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_59),
.A2(n_33),
.B1(n_27),
.B2(n_29),
.Y(n_98)
);

CKINVDCx5p33_ASAP7_75t_R g99 ( 
.A(n_67),
.Y(n_99)
);

AO21x2_ASAP7_75t_L g107 ( 
.A1(n_99),
.A2(n_17),
.B(n_55),
.Y(n_107)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_61),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_102),
.B(n_104),
.Y(n_123)
);

AOI21xp5_ASAP7_75t_L g103 ( 
.A1(n_59),
.A2(n_0),
.B(n_1),
.Y(n_103)
);

AOI21xp5_ASAP7_75t_L g113 ( 
.A1(n_103),
.A2(n_90),
.B(n_75),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_48),
.B(n_18),
.Y(n_104)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_48),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_105),
.Y(n_128)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_55),
.Y(n_106)
);

INVx6_ASAP7_75t_L g115 ( 
.A(n_106),
.Y(n_115)
);

CKINVDCx14_ASAP7_75t_R g160 ( 
.A(n_107),
.Y(n_160)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_81),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_108),
.B(n_132),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_112),
.A2(n_130),
.B1(n_72),
.B2(n_1),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_L g157 ( 
.A1(n_113),
.A2(n_72),
.B(n_15),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_114),
.B(n_78),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_100),
.A2(n_62),
.B1(n_69),
.B2(n_49),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_116),
.A2(n_119),
.B1(n_121),
.B2(n_98),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_88),
.A2(n_69),
.B1(n_49),
.B2(n_54),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_88),
.A2(n_82),
.B1(n_87),
.B2(n_71),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_L g124 ( 
.A1(n_96),
.A2(n_17),
.B1(n_23),
.B2(n_15),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_124),
.A2(n_77),
.B1(n_114),
.B2(n_120),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_96),
.B(n_71),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_127),
.B(n_133),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_88),
.A2(n_17),
.B1(n_67),
.B2(n_2),
.Y(n_130)
);

HAxp5_ASAP7_75t_SL g139 ( 
.A(n_131),
.B(n_113),
.CON(n_139),
.SN(n_139)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_81),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_95),
.B(n_17),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_135),
.B(n_130),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_136),
.A2(n_137),
.B1(n_141),
.B2(n_144),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_111),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_138),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_SL g183 ( 
.A1(n_139),
.A2(n_10),
.B(n_1),
.Y(n_183)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_120),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_140),
.B(n_146),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_109),
.A2(n_76),
.B1(n_102),
.B2(n_80),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g142 ( 
.A(n_121),
.B(n_101),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_142),
.B(n_118),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_109),
.A2(n_97),
.B1(n_101),
.B2(n_84),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_145),
.A2(n_149),
.B1(n_150),
.B2(n_153),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_127),
.B(n_95),
.Y(n_146)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_134),
.Y(n_147)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_147),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_119),
.A2(n_89),
.B1(n_85),
.B2(n_86),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_116),
.A2(n_74),
.B1(n_105),
.B2(n_106),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_151),
.B(n_155),
.Y(n_171)
);

INVxp67_ASAP7_75t_L g152 ( 
.A(n_122),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_152),
.B(n_163),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_131),
.A2(n_74),
.B1(n_73),
.B2(n_83),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_135),
.A2(n_73),
.B1(n_104),
.B2(n_92),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_154),
.A2(n_161),
.B1(n_107),
.B2(n_118),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_133),
.B(n_81),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_126),
.B(n_99),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_156),
.B(n_158),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_L g198 ( 
.A1(n_157),
.A2(n_0),
.B(n_2),
.Y(n_198)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_111),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_110),
.B(n_0),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_159),
.B(n_162),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_110),
.B(n_72),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_128),
.Y(n_163)
);

CKINVDCx16_ASAP7_75t_R g164 ( 
.A(n_107),
.Y(n_164)
);

INVxp67_ASAP7_75t_L g188 ( 
.A(n_164),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_125),
.B(n_123),
.Y(n_165)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_165),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_125),
.B(n_13),
.C(n_12),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_166),
.B(n_167),
.C(n_117),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_123),
.B(n_13),
.C(n_12),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_129),
.B(n_10),
.Y(n_168)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_168),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_169),
.B(n_182),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_176),
.A2(n_137),
.B1(n_141),
.B2(n_168),
.Y(n_211)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_148),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_177),
.B(n_191),
.Y(n_206)
);

AO22x1_ASAP7_75t_SL g178 ( 
.A1(n_164),
.A2(n_107),
.B1(n_112),
.B2(n_115),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_178),
.B(n_200),
.Y(n_205)
);

HB1xp67_ASAP7_75t_L g179 ( 
.A(n_155),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_179),
.Y(n_215)
);

AOI22xp33_ASAP7_75t_L g180 ( 
.A1(n_160),
.A2(n_107),
.B1(n_132),
.B2(n_108),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_180),
.A2(n_201),
.B1(n_144),
.B2(n_165),
.Y(n_203)
);

OAI32xp33_ASAP7_75t_L g181 ( 
.A1(n_151),
.A2(n_115),
.A3(n_134),
.B1(n_128),
.B2(n_10),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_SL g213 ( 
.A1(n_181),
.A2(n_183),
.B(n_186),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_142),
.B(n_117),
.Y(n_182)
);

BUFx2_ASAP7_75t_L g184 ( 
.A(n_148),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_184),
.Y(n_221)
);

AOI21xp5_ASAP7_75t_L g186 ( 
.A1(n_157),
.A2(n_160),
.B(n_138),
.Y(n_186)
);

AOI21xp5_ASAP7_75t_L g189 ( 
.A1(n_158),
.A2(n_153),
.B(n_145),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_L g212 ( 
.A1(n_189),
.A2(n_190),
.B(n_198),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_SL g190 ( 
.A1(n_140),
.A2(n_117),
.B(n_2),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_162),
.Y(n_191)
);

CKINVDCx16_ASAP7_75t_R g194 ( 
.A(n_150),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_194),
.B(n_196),
.Y(n_220)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_147),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_156),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_197),
.B(n_199),
.Y(n_209)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_163),
.Y(n_199)
);

AOI22xp33_ASAP7_75t_L g201 ( 
.A1(n_161),
.A2(n_3),
.B1(n_4),
.B2(n_6),
.Y(n_201)
);

INVxp67_ASAP7_75t_L g202 ( 
.A(n_149),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_202),
.B(n_178),
.Y(n_208)
);

CKINVDCx14_ASAP7_75t_R g236 ( 
.A(n_203),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_187),
.A2(n_136),
.B1(n_143),
.B2(n_146),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_204),
.A2(n_211),
.B1(n_214),
.B2(n_216),
.Y(n_231)
);

INVxp67_ASAP7_75t_L g207 ( 
.A(n_195),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_207),
.B(n_218),
.Y(n_244)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_208),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_182),
.B(n_143),
.C(n_154),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_210),
.B(n_219),
.C(n_205),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_188),
.A2(n_159),
.B1(n_167),
.B2(n_166),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_188),
.A2(n_172),
.B1(n_176),
.B2(n_202),
.Y(n_216)
);

INVx4_ASAP7_75t_L g217 ( 
.A(n_184),
.Y(n_217)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_217),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_170),
.B(n_3),
.Y(n_218)
);

INVx4_ASAP7_75t_L g222 ( 
.A(n_192),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_222),
.B(n_223),
.Y(n_249)
);

INVx1_ASAP7_75t_SL g223 ( 
.A(n_173),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_170),
.B(n_3),
.Y(n_224)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_224),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_172),
.A2(n_3),
.B1(n_4),
.B2(n_6),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_225),
.A2(n_228),
.B1(n_192),
.B2(n_196),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_174),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_226),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_173),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_227),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_187),
.A2(n_4),
.B1(n_7),
.B2(n_8),
.Y(n_228)
);

CKINVDCx14_ASAP7_75t_R g229 ( 
.A(n_175),
.Y(n_229)
);

INVxp67_ASAP7_75t_SL g245 ( 
.A(n_229),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_190),
.Y(n_230)
);

INVxp67_ASAP7_75t_L g248 ( 
.A(n_230),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_232),
.B(n_233),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_219),
.B(n_189),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_210),
.B(n_169),
.C(n_171),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_234),
.B(n_239),
.C(n_251),
.Y(n_255)
);

BUFx2_ASAP7_75t_L g235 ( 
.A(n_222),
.Y(n_235)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_235),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_205),
.B(n_171),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_238),
.B(n_247),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_204),
.B(n_191),
.C(n_200),
.Y(n_239)
);

HB1xp67_ASAP7_75t_L g240 ( 
.A(n_208),
.Y(n_240)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_240),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_SL g242 ( 
.A(n_209),
.B(n_193),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_SL g257 ( 
.A(n_242),
.B(n_209),
.Y(n_257)
);

AOI22x1_ASAP7_75t_L g243 ( 
.A1(n_230),
.A2(n_178),
.B1(n_186),
.B2(n_181),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_243),
.A2(n_203),
.B1(n_223),
.B2(n_228),
.Y(n_259)
);

OA22x2_ASAP7_75t_L g246 ( 
.A1(n_227),
.A2(n_198),
.B1(n_177),
.B2(n_185),
.Y(n_246)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_246),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_211),
.B(n_175),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_216),
.B(n_212),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_253),
.A2(n_217),
.B1(n_221),
.B2(n_215),
.Y(n_260)
);

AOI21xp5_ASAP7_75t_L g256 ( 
.A1(n_248),
.A2(n_243),
.B(n_237),
.Y(n_256)
);

OAI21xp5_ASAP7_75t_L g279 ( 
.A1(n_256),
.A2(n_213),
.B(n_246),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_257),
.B(n_264),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_250),
.B(n_226),
.Y(n_258)
);

INVxp67_ASAP7_75t_L g285 ( 
.A(n_258),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_259),
.A2(n_260),
.B1(n_262),
.B2(n_254),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_236),
.A2(n_220),
.B1(n_221),
.B2(n_215),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_245),
.B(n_220),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_232),
.B(n_206),
.C(n_212),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_267),
.B(n_270),
.C(n_234),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_L g269 ( 
.A1(n_243),
.A2(n_225),
.B1(n_206),
.B2(n_224),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_269),
.A2(n_273),
.B1(n_253),
.B2(n_231),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_239),
.B(n_213),
.C(n_214),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_249),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_271),
.B(n_272),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_252),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_L g273 ( 
.A1(n_248),
.A2(n_244),
.B1(n_241),
.B2(n_218),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g291 ( 
.A(n_274),
.B(n_284),
.Y(n_291)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_275),
.Y(n_290)
);

AND2x2_ASAP7_75t_L g276 ( 
.A(n_260),
.B(n_251),
.Y(n_276)
);

OAI21xp5_ASAP7_75t_L g297 ( 
.A1(n_276),
.A2(n_279),
.B(n_265),
.Y(n_297)
);

BUFx6f_ASAP7_75t_L g277 ( 
.A(n_268),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_277),
.B(n_254),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_255),
.B(n_267),
.C(n_270),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_280),
.B(n_271),
.C(n_265),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_255),
.B(n_233),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_281),
.B(n_286),
.Y(n_298)
);

BUFx2_ASAP7_75t_L g282 ( 
.A(n_256),
.Y(n_282)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_282),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_283),
.B(n_259),
.Y(n_292)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_263),
.B(n_238),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_263),
.B(n_247),
.Y(n_286)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_266),
.B(n_231),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_287),
.B(n_266),
.Y(n_289)
);

XOR2xp5_ASAP7_75t_L g306 ( 
.A(n_289),
.B(n_284),
.Y(n_306)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_292),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_294),
.B(n_295),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_280),
.B(n_261),
.C(n_262),
.Y(n_295)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_296),
.Y(n_311)
);

AOI21xp5_ASAP7_75t_L g305 ( 
.A1(n_297),
.A2(n_276),
.B(n_285),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_282),
.A2(n_261),
.B1(n_246),
.B2(n_235),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_299),
.A2(n_287),
.B1(n_278),
.B2(n_274),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_SL g300 ( 
.A(n_285),
.B(n_246),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_300),
.B(n_301),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_277),
.B(n_183),
.Y(n_301)
);

AND2x2_ASAP7_75t_L g302 ( 
.A(n_295),
.B(n_288),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_302),
.B(n_303),
.Y(n_315)
);

INVxp67_ASAP7_75t_L g303 ( 
.A(n_299),
.Y(n_303)
);

OAI21xp5_ASAP7_75t_SL g314 ( 
.A1(n_305),
.A2(n_293),
.B(n_290),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_306),
.B(n_291),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_307),
.B(n_289),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_294),
.B(n_4),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_309),
.B(n_7),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_312),
.B(n_316),
.Y(n_320)
);

AOI21xp5_ASAP7_75t_L g321 ( 
.A1(n_313),
.A2(n_314),
.B(n_318),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_310),
.B(n_297),
.Y(n_317)
);

CKINVDCx14_ASAP7_75t_R g322 ( 
.A(n_317),
.Y(n_322)
);

OAI21xp5_ASAP7_75t_SL g318 ( 
.A1(n_308),
.A2(n_298),
.B(n_291),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_315),
.B(n_304),
.Y(n_319)
);

OAI211xp5_ASAP7_75t_L g324 ( 
.A1(n_319),
.A2(n_311),
.B(n_303),
.C(n_306),
.Y(n_324)
);

AOI21xp5_ASAP7_75t_SL g323 ( 
.A1(n_321),
.A2(n_312),
.B(n_302),
.Y(n_323)
);

OAI21xp5_ASAP7_75t_SL g325 ( 
.A1(n_323),
.A2(n_324),
.B(n_320),
.Y(n_325)
);

XNOR2xp5_ASAP7_75t_L g326 ( 
.A(n_325),
.B(n_322),
.Y(n_326)
);

OAI21xp5_ASAP7_75t_SL g327 ( 
.A1(n_326),
.A2(n_8),
.B(n_9),
.Y(n_327)
);

MAJx2_ASAP7_75t_L g328 ( 
.A(n_327),
.B(n_8),
.C(n_9),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_L g329 ( 
.A1(n_328),
.A2(n_8),
.B1(n_9),
.B2(n_250),
.Y(n_329)
);


endmodule