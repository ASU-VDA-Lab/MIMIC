module fake_netlist_6_1028_n_876 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_166, n_28, n_184, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_188, n_102, n_186, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_104, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_187, n_89, n_173, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_171, n_31, n_57, n_169, n_53, n_51, n_44, n_56, n_876);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_184;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_188;
input n_102;
input n_186;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_104;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_187;
input n_89;
input n_173;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_171;
input n_31;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_876;

wire n_591;
wire n_435;
wire n_793;
wire n_326;
wire n_801;
wire n_256;
wire n_853;
wire n_440;
wire n_587;
wire n_695;
wire n_507;
wire n_580;
wire n_762;
wire n_875;
wire n_209;
wire n_367;
wire n_465;
wire n_680;
wire n_760;
wire n_741;
wire n_590;
wire n_625;
wire n_661;
wire n_223;
wire n_278;
wire n_341;
wire n_362;
wire n_226;
wire n_828;
wire n_208;
wire n_462;
wire n_607;
wire n_671;
wire n_726;
wire n_316;
wire n_419;
wire n_304;
wire n_212;
wire n_700;
wire n_694;
wire n_740;
wire n_578;
wire n_703;
wire n_365;
wire n_384;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_342;
wire n_820;
wire n_783;
wire n_725;
wire n_358;
wire n_751;
wire n_449;
wire n_749;
wire n_798;
wire n_310;
wire n_509;
wire n_245;
wire n_368;
wire n_575;
wire n_677;
wire n_805;
wire n_396;
wire n_495;
wire n_815;
wire n_350;
wire n_585;
wire n_732;
wire n_568;
wire n_392;
wire n_840;
wire n_442;
wire n_480;
wire n_874;
wire n_724;
wire n_382;
wire n_673;
wire n_628;
wire n_557;
wire n_823;
wire n_349;
wire n_643;
wire n_233;
wire n_617;
wire n_698;
wire n_845;
wire n_255;
wire n_807;
wire n_739;
wire n_284;
wire n_400;
wire n_337;
wire n_865;
wire n_214;
wire n_485;
wire n_443;
wire n_246;
wire n_768;
wire n_471;
wire n_289;
wire n_421;
wire n_781;
wire n_424;
wire n_789;
wire n_615;
wire n_238;
wire n_573;
wire n_769;
wire n_202;
wire n_320;
wire n_639;
wire n_676;
wire n_327;
wire n_794;
wire n_727;
wire n_369;
wire n_597;
wire n_685;
wire n_280;
wire n_287;
wire n_832;
wire n_353;
wire n_610;
wire n_555;
wire n_389;
wire n_814;
wire n_415;
wire n_830;
wire n_230;
wire n_605;
wire n_461;
wire n_873;
wire n_383;
wire n_826;
wire n_669;
wire n_200;
wire n_447;
wire n_872;
wire n_198;
wire n_300;
wire n_222;
wire n_248;
wire n_517;
wire n_718;
wire n_747;
wire n_852;
wire n_667;
wire n_229;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_621;
wire n_305;
wire n_721;
wire n_750;
wire n_532;
wire n_742;
wire n_535;
wire n_691;
wire n_250;
wire n_372;
wire n_468;
wire n_544;
wire n_504;
wire n_314;
wire n_378;
wire n_413;
wire n_377;
wire n_791;
wire n_510;
wire n_837;
wire n_836;
wire n_863;
wire n_375;
wire n_601;
wire n_338;
wire n_522;
wire n_466;
wire n_704;
wire n_748;
wire n_506;
wire n_763;
wire n_360;
wire n_603;
wire n_235;
wire n_536;
wire n_866;
wire n_622;
wire n_191;
wire n_340;
wire n_710;
wire n_387;
wire n_452;
wire n_658;
wire n_616;
wire n_744;
wire n_344;
wire n_581;
wire n_428;
wire n_785;
wire n_761;
wire n_746;
wire n_609;
wire n_765;
wire n_432;
wire n_641;
wire n_822;
wire n_693;
wire n_631;
wire n_516;
wire n_720;
wire n_525;
wire n_758;
wire n_842;
wire n_611;
wire n_491;
wire n_656;
wire n_772;
wire n_843;
wire n_797;
wire n_666;
wire n_371;
wire n_795;
wire n_770;
wire n_567;
wire n_189;
wire n_738;
wire n_405;
wire n_213;
wire n_538;
wire n_294;
wire n_302;
wire n_499;
wire n_380;
wire n_838;
wire n_705;
wire n_647;
wire n_197;
wire n_343;
wire n_844;
wire n_448;
wire n_494;
wire n_539;
wire n_493;
wire n_397;
wire n_614;
wire n_529;
wire n_445;
wire n_425;
wire n_684;
wire n_454;
wire n_218;
wire n_638;
wire n_234;
wire n_486;
wire n_381;
wire n_236;
wire n_653;
wire n_752;
wire n_713;
wire n_648;
wire n_657;
wire n_576;
wire n_472;
wire n_270;
wire n_239;
wire n_414;
wire n_563;
wire n_782;
wire n_490;
wire n_803;
wire n_290;
wire n_220;
wire n_809;
wire n_224;
wire n_839;
wire n_734;
wire n_708;
wire n_196;
wire n_402;
wire n_352;
wire n_668;
wire n_478;
wire n_626;
wire n_574;
wire n_800;
wire n_779;
wire n_460;
wire n_854;
wire n_417;
wire n_446;
wire n_498;
wire n_662;
wire n_374;
wire n_659;
wire n_709;
wire n_870;
wire n_366;
wire n_777;
wire n_407;
wire n_450;
wire n_808;
wire n_867;
wire n_272;
wire n_526;
wire n_712;
wire n_348;
wire n_711;
wire n_579;
wire n_376;
wire n_390;
wire n_473;
wire n_293;
wire n_334;
wire n_559;
wire n_370;
wire n_458;
wire n_232;
wire n_650;
wire n_717;
wire n_330;
wire n_771;
wire n_470;
wire n_475;
wire n_298;
wire n_492;
wire n_281;
wire n_258;
wire n_551;
wire n_699;
wire n_456;
wire n_564;
wire n_265;
wire n_260;
wire n_313;
wire n_451;
wire n_624;
wire n_824;
wire n_279;
wire n_686;
wire n_796;
wire n_252;
wire n_757;
wire n_228;
wire n_565;
wire n_594;
wire n_719;
wire n_356;
wire n_577;
wire n_552;
wire n_619;
wire n_216;
wire n_455;
wire n_521;
wire n_363;
wire n_572;
wire n_395;
wire n_813;
wire n_592;
wire n_745;
wire n_654;
wire n_323;
wire n_829;
wire n_606;
wire n_393;
wire n_818;
wire n_411;
wire n_503;
wire n_716;
wire n_623;
wire n_599;
wire n_513;
wire n_855;
wire n_776;
wire n_321;
wire n_645;
wire n_331;
wire n_227;
wire n_868;
wire n_570;
wire n_731;
wire n_859;
wire n_406;
wire n_483;
wire n_735;
wire n_204;
wire n_482;
wire n_755;
wire n_474;
wire n_527;
wire n_261;
wire n_608;
wire n_620;
wire n_420;
wire n_683;
wire n_630;
wire n_312;
wire n_394;
wire n_519;
wire n_541;
wire n_512;
wire n_292;
wire n_307;
wire n_469;
wire n_433;
wire n_500;
wire n_792;
wire n_476;
wire n_714;
wire n_291;
wire n_219;
wire n_543;
wire n_357;
wire n_264;
wire n_263;
wire n_589;
wire n_860;
wire n_481;
wire n_788;
wire n_819;
wire n_821;
wire n_325;
wire n_767;
wire n_804;
wire n_329;
wire n_464;
wire n_600;
wire n_831;
wire n_802;
wire n_561;
wire n_477;
wire n_549;
wire n_533;
wire n_408;
wire n_806;
wire n_864;
wire n_237;
wire n_584;
wire n_244;
wire n_399;
wire n_243;
wire n_548;
wire n_282;
wire n_436;
wire n_833;
wire n_211;
wire n_523;
wire n_322;
wire n_707;
wire n_345;
wire n_409;
wire n_231;
wire n_354;
wire n_689;
wire n_799;
wire n_505;
wire n_240;
wire n_756;
wire n_319;
wire n_547;
wire n_537;
wire n_273;
wire n_558;
wire n_810;
wire n_635;
wire n_787;
wire n_311;
wire n_403;
wire n_723;
wire n_253;
wire n_634;
wire n_583;
wire n_596;
wire n_546;
wire n_562;
wire n_249;
wire n_201;
wire n_386;
wire n_764;
wire n_556;
wire n_692;
wire n_733;
wire n_754;
wire n_487;
wire n_550;
wire n_241;
wire n_275;
wire n_553;
wire n_652;
wire n_849;
wire n_560;
wire n_753;
wire n_642;
wire n_276;
wire n_569;
wire n_441;
wire n_221;
wire n_811;
wire n_444;
wire n_586;
wire n_423;
wire n_737;
wire n_318;
wire n_303;
wire n_511;
wire n_715;
wire n_467;
wire n_306;
wire n_193;
wire n_269;
wire n_359;
wire n_346;
wire n_416;
wire n_530;
wire n_277;
wire n_520;
wire n_418;
wire n_618;
wire n_790;
wire n_582;
wire n_199;
wire n_266;
wire n_296;
wire n_861;
wire n_674;
wire n_857;
wire n_871;
wire n_775;
wire n_571;
wire n_268;
wire n_271;
wire n_404;
wire n_651;
wire n_439;
wire n_217;
wire n_210;
wire n_299;
wire n_518;
wire n_206;
wire n_679;
wire n_453;
wire n_612;
wire n_633;
wire n_665;
wire n_333;
wire n_588;
wire n_215;
wire n_247;
wire n_225;
wire n_308;
wire n_309;
wire n_759;
wire n_355;
wire n_426;
wire n_317;
wire n_632;
wire n_702;
wire n_431;
wire n_347;
wire n_812;
wire n_459;
wire n_502;
wire n_328;
wire n_672;
wire n_534;
wire n_488;
wire n_429;
wire n_373;
wire n_195;
wire n_285;
wire n_497;
wire n_780;
wire n_773;
wire n_675;
wire n_257;
wire n_730;
wire n_655;
wire n_706;
wire n_786;
wire n_670;
wire n_203;
wire n_286;
wire n_254;
wire n_207;
wire n_834;
wire n_242;
wire n_835;
wire n_690;
wire n_850;
wire n_401;
wire n_324;
wire n_766;
wire n_816;
wire n_743;
wire n_335;
wire n_430;
wire n_463;
wire n_545;
wire n_489;
wire n_205;
wire n_604;
wire n_848;
wire n_251;
wire n_301;
wire n_274;
wire n_636;
wire n_825;
wire n_728;
wire n_681;
wire n_729;
wire n_774;
wire n_412;
wire n_640;
wire n_660;
wire n_267;
wire n_438;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_515;
wire n_288;
wire n_427;
wire n_479;
wire n_496;
wire n_598;
wire n_422;
wire n_696;
wire n_688;
wire n_722;
wire n_862;
wire n_351;
wire n_869;
wire n_437;
wire n_259;
wire n_540;
wire n_593;
wire n_514;
wire n_646;
wire n_528;
wire n_391;
wire n_457;
wire n_697;
wire n_687;
wire n_364;
wire n_637;
wire n_295;
wire n_385;
wire n_701;
wire n_817;
wire n_629;
wire n_388;
wire n_190;
wire n_858;
wire n_262;
wire n_484;
wire n_613;
wire n_736;
wire n_846;
wire n_501;
wire n_841;
wire n_531;
wire n_827;
wire n_361;
wire n_508;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_332;
wire n_336;
wire n_398;
wire n_410;
wire n_566;
wire n_554;
wire n_602;
wire n_194;
wire n_664;
wire n_678;
wire n_192;
wire n_649;
wire n_283;

NOR2xp67_ASAP7_75t_L g189 ( 
.A(n_163),
.B(n_168),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_146),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_110),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_49),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_184),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_17),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g195 ( 
.A(n_123),
.Y(n_195)
);

BUFx6f_ASAP7_75t_L g196 ( 
.A(n_52),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_137),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_67),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_39),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_138),
.Y(n_200)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_160),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_76),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_56),
.Y(n_203)
);

BUFx10_ASAP7_75t_L g204 ( 
.A(n_3),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_154),
.Y(n_205)
);

BUFx3_ASAP7_75t_L g206 ( 
.A(n_18),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_132),
.Y(n_207)
);

INVx2_ASAP7_75t_SL g208 ( 
.A(n_141),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_89),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_134),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_2),
.Y(n_211)
);

BUFx6f_ASAP7_75t_L g212 ( 
.A(n_148),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_158),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_156),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_74),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_14),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_145),
.Y(n_217)
);

CKINVDCx16_ASAP7_75t_R g218 ( 
.A(n_99),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_73),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_159),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_187),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_85),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_61),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_44),
.Y(n_224)
);

BUFx2_ASAP7_75t_L g225 ( 
.A(n_136),
.Y(n_225)
);

CKINVDCx16_ASAP7_75t_R g226 ( 
.A(n_128),
.Y(n_226)
);

CKINVDCx16_ASAP7_75t_R g227 ( 
.A(n_92),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_127),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_63),
.Y(n_229)
);

INVx1_ASAP7_75t_SL g230 ( 
.A(n_139),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_179),
.Y(n_231)
);

BUFx6f_ASAP7_75t_L g232 ( 
.A(n_135),
.Y(n_232)
);

BUFx10_ASAP7_75t_L g233 ( 
.A(n_72),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_150),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_153),
.Y(n_235)
);

BUFx10_ASAP7_75t_L g236 ( 
.A(n_14),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_175),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_54),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_126),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_20),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_174),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_106),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_178),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_96),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_105),
.Y(n_245)
);

INVx2_ASAP7_75t_SL g246 ( 
.A(n_171),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_4),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_25),
.Y(n_248)
);

INVx2_ASAP7_75t_SL g249 ( 
.A(n_119),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_71),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_180),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_97),
.Y(n_252)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_173),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_10),
.Y(n_254)
);

BUFx2_ASAP7_75t_L g255 ( 
.A(n_133),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_176),
.Y(n_256)
);

BUFx3_ASAP7_75t_L g257 ( 
.A(n_182),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_68),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_41),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_131),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_81),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_130),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_177),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_120),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_206),
.Y(n_265)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_216),
.Y(n_266)
);

AND2x2_ASAP7_75t_L g267 ( 
.A(n_225),
.B(n_0),
.Y(n_267)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_240),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_247),
.Y(n_269)
);

BUFx12f_ASAP7_75t_L g270 ( 
.A(n_204),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_194),
.Y(n_271)
);

BUFx2_ASAP7_75t_L g272 ( 
.A(n_211),
.Y(n_272)
);

HB1xp67_ASAP7_75t_L g273 ( 
.A(n_254),
.Y(n_273)
);

AND2x4_ASAP7_75t_L g274 ( 
.A(n_257),
.B(n_21),
.Y(n_274)
);

HB1xp67_ASAP7_75t_L g275 ( 
.A(n_255),
.Y(n_275)
);

INVxp67_ASAP7_75t_L g276 ( 
.A(n_204),
.Y(n_276)
);

BUFx12f_ASAP7_75t_L g277 ( 
.A(n_236),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_191),
.Y(n_278)
);

BUFx6f_ASAP7_75t_L g279 ( 
.A(n_195),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_208),
.B(n_0),
.Y(n_280)
);

AOI22x1_ASAP7_75t_SL g281 ( 
.A1(n_200),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_281)
);

BUFx12f_ASAP7_75t_L g282 ( 
.A(n_236),
.Y(n_282)
);

HB1xp67_ASAP7_75t_L g283 ( 
.A(n_193),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_217),
.Y(n_284)
);

BUFx3_ASAP7_75t_L g285 ( 
.A(n_233),
.Y(n_285)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_195),
.Y(n_286)
);

INVxp33_ASAP7_75t_SL g287 ( 
.A(n_190),
.Y(n_287)
);

INVxp67_ASAP7_75t_L g288 ( 
.A(n_233),
.Y(n_288)
);

OAI21x1_ASAP7_75t_L g289 ( 
.A1(n_201),
.A2(n_1),
.B(n_4),
.Y(n_289)
);

INVx2_ASAP7_75t_SL g290 ( 
.A(n_195),
.Y(n_290)
);

BUFx8_ASAP7_75t_SL g291 ( 
.A(n_252),
.Y(n_291)
);

BUFx6f_ASAP7_75t_L g292 ( 
.A(n_195),
.Y(n_292)
);

AND2x6_ASAP7_75t_L g293 ( 
.A(n_196),
.B(n_22),
.Y(n_293)
);

INVx5_ASAP7_75t_L g294 ( 
.A(n_196),
.Y(n_294)
);

INVx6_ASAP7_75t_L g295 ( 
.A(n_196),
.Y(n_295)
);

AND2x2_ASAP7_75t_L g296 ( 
.A(n_218),
.B(n_5),
.Y(n_296)
);

INVx3_ASAP7_75t_L g297 ( 
.A(n_196),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_226),
.Y(n_298)
);

BUFx12f_ASAP7_75t_L g299 ( 
.A(n_192),
.Y(n_299)
);

BUFx12f_ASAP7_75t_L g300 ( 
.A(n_197),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_246),
.B(n_5),
.Y(n_301)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_212),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_L g303 ( 
.A1(n_227),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_303)
);

BUFx6f_ASAP7_75t_L g304 ( 
.A(n_212),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_SL g305 ( 
.A(n_212),
.B(n_6),
.Y(n_305)
);

INVx2_ASAP7_75t_L g306 ( 
.A(n_212),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_220),
.Y(n_307)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_232),
.Y(n_308)
);

AND2x4_ASAP7_75t_L g309 ( 
.A(n_249),
.B(n_23),
.Y(n_309)
);

OAI21x1_ASAP7_75t_L g310 ( 
.A1(n_253),
.A2(n_7),
.B(n_8),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_222),
.Y(n_311)
);

INVx3_ASAP7_75t_L g312 ( 
.A(n_232),
.Y(n_312)
);

INVx2_ASAP7_75t_SL g313 ( 
.A(n_232),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_223),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_198),
.Y(n_315)
);

BUFx12f_ASAP7_75t_L g316 ( 
.A(n_199),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_295),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_291),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_291),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_315),
.Y(n_320)
);

BUFx2_ASAP7_75t_L g321 ( 
.A(n_271),
.Y(n_321)
);

INVx6_ASAP7_75t_L g322 ( 
.A(n_299),
.Y(n_322)
);

BUFx3_ASAP7_75t_L g323 ( 
.A(n_274),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_315),
.Y(n_324)
);

INVx3_ASAP7_75t_L g325 ( 
.A(n_279),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_295),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_299),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_280),
.B(n_230),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_271),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_300),
.Y(n_330)
);

INVxp67_ASAP7_75t_SL g331 ( 
.A(n_266),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_SL g332 ( 
.A(n_296),
.B(n_232),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_300),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_R g334 ( 
.A(n_298),
.B(n_258),
.Y(n_334)
);

AND2x6_ASAP7_75t_L g335 ( 
.A(n_309),
.B(n_228),
.Y(n_335)
);

INVx3_ASAP7_75t_L g336 ( 
.A(n_279),
.Y(n_336)
);

BUFx2_ASAP7_75t_L g337 ( 
.A(n_298),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_295),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_316),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_316),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_287),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_309),
.B(n_231),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_278),
.Y(n_343)
);

BUFx10_ASAP7_75t_L g344 ( 
.A(n_275),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_284),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_287),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_307),
.Y(n_347)
);

CKINVDCx20_ASAP7_75t_R g348 ( 
.A(n_272),
.Y(n_348)
);

BUFx3_ASAP7_75t_L g349 ( 
.A(n_274),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_R g350 ( 
.A(n_270),
.B(n_262),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_311),
.Y(n_351)
);

CKINVDCx16_ASAP7_75t_R g352 ( 
.A(n_270),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_314),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_277),
.Y(n_354)
);

INVx2_ASAP7_75t_L g355 ( 
.A(n_279),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_277),
.Y(n_356)
);

INVx2_ASAP7_75t_L g357 ( 
.A(n_279),
.Y(n_357)
);

INVx2_ASAP7_75t_L g358 ( 
.A(n_292),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_282),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_282),
.Y(n_360)
);

CKINVDCx20_ASAP7_75t_R g361 ( 
.A(n_273),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_269),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_SL g363 ( 
.A(n_296),
.B(n_189),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_285),
.Y(n_364)
);

INVx2_ASAP7_75t_L g365 ( 
.A(n_292),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_309),
.B(n_244),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_285),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_288),
.Y(n_368)
);

INVx3_ASAP7_75t_L g369 ( 
.A(n_292),
.Y(n_369)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_292),
.Y(n_370)
);

OA21x2_ASAP7_75t_L g371 ( 
.A1(n_289),
.A2(n_251),
.B(n_248),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_283),
.Y(n_372)
);

OR2x6_ASAP7_75t_L g373 ( 
.A(n_322),
.B(n_303),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_331),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_R g375 ( 
.A(n_318),
.B(n_202),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_SL g376 ( 
.A(n_363),
.B(n_267),
.Y(n_376)
);

INVx2_ASAP7_75t_L g377 ( 
.A(n_325),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_L g378 ( 
.A(n_328),
.B(n_267),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_323),
.B(n_274),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_331),
.Y(n_380)
);

BUFx8_ASAP7_75t_L g381 ( 
.A(n_321),
.Y(n_381)
);

NAND2xp33_ASAP7_75t_SL g382 ( 
.A(n_334),
.B(n_305),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_323),
.B(n_290),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_L g384 ( 
.A(n_328),
.B(n_276),
.Y(n_384)
);

INVx2_ASAP7_75t_SL g385 ( 
.A(n_344),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_349),
.B(n_290),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_SL g387 ( 
.A(n_364),
.B(n_301),
.Y(n_387)
);

OAI21xp5_ASAP7_75t_L g388 ( 
.A1(n_342),
.A2(n_310),
.B(n_289),
.Y(n_388)
);

INVx3_ASAP7_75t_L g389 ( 
.A(n_325),
.Y(n_389)
);

OR2x2_ASAP7_75t_L g390 ( 
.A(n_332),
.B(n_265),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_349),
.B(n_313),
.Y(n_391)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_336),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_SL g393 ( 
.A(n_367),
.B(n_203),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_L g394 ( 
.A(n_372),
.B(n_305),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_366),
.B(n_313),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_L g396 ( 
.A(n_368),
.B(n_205),
.Y(n_396)
);

NOR3xp33_ASAP7_75t_L g397 ( 
.A(n_337),
.B(n_260),
.C(n_256),
.Y(n_397)
);

INVxp33_ASAP7_75t_L g398 ( 
.A(n_334),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_SL g399 ( 
.A(n_320),
.B(n_207),
.Y(n_399)
);

NOR3xp33_ASAP7_75t_L g400 ( 
.A(n_332),
.B(n_264),
.C(n_263),
.Y(n_400)
);

INVx2_ASAP7_75t_L g401 ( 
.A(n_336),
.Y(n_401)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_369),
.Y(n_402)
);

INVx2_ASAP7_75t_L g403 ( 
.A(n_369),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_L g404 ( 
.A(n_324),
.B(n_209),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_SL g405 ( 
.A(n_341),
.B(n_210),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_362),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_335),
.B(n_294),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_335),
.B(n_286),
.Y(n_408)
);

INVx2_ASAP7_75t_L g409 ( 
.A(n_355),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_SL g410 ( 
.A(n_346),
.B(n_213),
.Y(n_410)
);

INVxp33_ASAP7_75t_L g411 ( 
.A(n_350),
.Y(n_411)
);

NOR3xp33_ASAP7_75t_L g412 ( 
.A(n_352),
.B(n_268),
.C(n_266),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_335),
.B(n_286),
.Y(n_413)
);

AND2x2_ASAP7_75t_L g414 ( 
.A(n_344),
.B(n_268),
.Y(n_414)
);

BUFx3_ASAP7_75t_L g415 ( 
.A(n_317),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_343),
.Y(n_416)
);

NAND2x1_ASAP7_75t_L g417 ( 
.A(n_335),
.B(n_293),
.Y(n_417)
);

NOR2xp33_ASAP7_75t_L g418 ( 
.A(n_345),
.B(n_214),
.Y(n_418)
);

BUFx6f_ASAP7_75t_SL g419 ( 
.A(n_347),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_SL g420 ( 
.A(n_350),
.B(n_215),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_335),
.B(n_294),
.Y(n_421)
);

BUFx5_ASAP7_75t_L g422 ( 
.A(n_351),
.Y(n_422)
);

AND2x2_ASAP7_75t_L g423 ( 
.A(n_353),
.B(n_302),
.Y(n_423)
);

AOI22xp33_ASAP7_75t_L g424 ( 
.A1(n_371),
.A2(n_310),
.B1(n_293),
.B2(n_297),
.Y(n_424)
);

NOR2xp33_ASAP7_75t_L g425 ( 
.A(n_326),
.B(n_219),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_357),
.B(n_294),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_SL g427 ( 
.A(n_327),
.B(n_221),
.Y(n_427)
);

AOI221xp5_ASAP7_75t_L g428 ( 
.A1(n_361),
.A2(n_245),
.B1(n_229),
.B2(n_234),
.C(n_235),
.Y(n_428)
);

NOR2xp33_ASAP7_75t_L g429 ( 
.A(n_338),
.B(n_224),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_358),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_365),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_370),
.B(n_294),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_SL g433 ( 
.A(n_330),
.B(n_237),
.Y(n_433)
);

A2O1A1Ixp33_ASAP7_75t_L g434 ( 
.A1(n_371),
.A2(n_308),
.B(n_306),
.C(n_302),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_371),
.B(n_306),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_322),
.Y(n_436)
);

AND2x2_ASAP7_75t_L g437 ( 
.A(n_322),
.B(n_308),
.Y(n_437)
);

INVxp67_ASAP7_75t_L g438 ( 
.A(n_354),
.Y(n_438)
);

AOI22xp5_ASAP7_75t_L g439 ( 
.A1(n_348),
.A2(n_259),
.B1(n_239),
.B2(n_241),
.Y(n_439)
);

INVx2_ASAP7_75t_L g440 ( 
.A(n_333),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_339),
.B(n_297),
.Y(n_441)
);

OAI21xp5_ASAP7_75t_L g442 ( 
.A1(n_435),
.A2(n_293),
.B(n_297),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_406),
.Y(n_443)
);

AOI22xp33_ASAP7_75t_L g444 ( 
.A1(n_378),
.A2(n_293),
.B1(n_312),
.B2(n_243),
.Y(n_444)
);

AO22x1_ASAP7_75t_L g445 ( 
.A1(n_394),
.A2(n_293),
.B1(n_340),
.B2(n_238),
.Y(n_445)
);

INVx3_ASAP7_75t_L g446 ( 
.A(n_389),
.Y(n_446)
);

NOR2x2_ASAP7_75t_L g447 ( 
.A(n_373),
.B(n_281),
.Y(n_447)
);

BUFx3_ASAP7_75t_L g448 ( 
.A(n_415),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_416),
.Y(n_449)
);

BUFx3_ASAP7_75t_L g450 ( 
.A(n_381),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_423),
.Y(n_451)
);

INVx2_ASAP7_75t_SL g452 ( 
.A(n_414),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_383),
.Y(n_453)
);

INVx3_ASAP7_75t_L g454 ( 
.A(n_389),
.Y(n_454)
);

NOR2xp33_ASAP7_75t_L g455 ( 
.A(n_384),
.B(n_374),
.Y(n_455)
);

INVx2_ASAP7_75t_SL g456 ( 
.A(n_390),
.Y(n_456)
);

AOI21xp5_ASAP7_75t_L g457 ( 
.A1(n_379),
.A2(n_294),
.B(n_304),
.Y(n_457)
);

INVx2_ASAP7_75t_L g458 ( 
.A(n_409),
.Y(n_458)
);

INVx2_ASAP7_75t_L g459 ( 
.A(n_377),
.Y(n_459)
);

INVx2_ASAP7_75t_SL g460 ( 
.A(n_437),
.Y(n_460)
);

INVx3_ASAP7_75t_L g461 ( 
.A(n_392),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_380),
.B(n_242),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_395),
.B(n_250),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_386),
.Y(n_464)
);

INVx4_ASAP7_75t_L g465 ( 
.A(n_422),
.Y(n_465)
);

OAI22xp5_ASAP7_75t_L g466 ( 
.A1(n_376),
.A2(n_261),
.B1(n_312),
.B2(n_356),
.Y(n_466)
);

HB1xp67_ASAP7_75t_L g467 ( 
.A(n_395),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_422),
.B(n_293),
.Y(n_468)
);

INVx2_ASAP7_75t_SL g469 ( 
.A(n_441),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_391),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_430),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_422),
.B(n_312),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_431),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_422),
.B(n_304),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_401),
.Y(n_475)
);

NOR2xp33_ASAP7_75t_L g476 ( 
.A(n_404),
.B(n_9),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_402),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_422),
.B(n_304),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_403),
.Y(n_479)
);

INVx2_ASAP7_75t_L g480 ( 
.A(n_435),
.Y(n_480)
);

OR2x2_ASAP7_75t_L g481 ( 
.A(n_385),
.B(n_359),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_SL g482 ( 
.A(n_382),
.B(n_360),
.Y(n_482)
);

AOI22xp33_ASAP7_75t_L g483 ( 
.A1(n_388),
.A2(n_304),
.B1(n_329),
.B2(n_319),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_434),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_418),
.B(n_24),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g486 ( 
.A(n_424),
.B(n_26),
.Y(n_486)
);

INVx2_ASAP7_75t_L g487 ( 
.A(n_408),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_SL g488 ( 
.A(n_388),
.B(n_408),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_413),
.Y(n_489)
);

AOI22xp33_ASAP7_75t_L g490 ( 
.A1(n_400),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_490)
);

AOI22xp33_ASAP7_75t_L g491 ( 
.A1(n_413),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_396),
.B(n_27),
.Y(n_492)
);

NAND3xp33_ASAP7_75t_SL g493 ( 
.A(n_428),
.B(n_397),
.C(n_439),
.Y(n_493)
);

CKINVDCx5p33_ASAP7_75t_R g494 ( 
.A(n_375),
.Y(n_494)
);

NOR2xp33_ASAP7_75t_L g495 ( 
.A(n_387),
.B(n_12),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_425),
.B(n_28),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_429),
.B(n_29),
.Y(n_497)
);

HB1xp67_ASAP7_75t_L g498 ( 
.A(n_373),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_441),
.Y(n_499)
);

AOI22xp5_ASAP7_75t_L g500 ( 
.A1(n_399),
.A2(n_101),
.B1(n_186),
.B2(n_185),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_426),
.Y(n_501)
);

INVx2_ASAP7_75t_SL g502 ( 
.A(n_373),
.Y(n_502)
);

INVx2_ASAP7_75t_SL g503 ( 
.A(n_436),
.Y(n_503)
);

CKINVDCx5p33_ASAP7_75t_R g504 ( 
.A(n_381),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_393),
.B(n_30),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_SL g506 ( 
.A(n_398),
.B(n_31),
.Y(n_506)
);

INVx1_ASAP7_75t_SL g507 ( 
.A(n_405),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_432),
.Y(n_508)
);

CKINVDCx5p33_ASAP7_75t_R g509 ( 
.A(n_419),
.Y(n_509)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_417),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_410),
.Y(n_511)
);

NOR2xp33_ASAP7_75t_L g512 ( 
.A(n_455),
.B(n_411),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_L g513 ( 
.A(n_455),
.B(n_420),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_480),
.B(n_412),
.Y(n_514)
);

AOI21xp5_ASAP7_75t_L g515 ( 
.A1(n_465),
.A2(n_421),
.B(n_407),
.Y(n_515)
);

INVx3_ASAP7_75t_L g516 ( 
.A(n_446),
.Y(n_516)
);

O2A1O1Ixp33_ASAP7_75t_L g517 ( 
.A1(n_476),
.A2(n_433),
.B(n_427),
.C(n_440),
.Y(n_517)
);

BUFx6f_ASAP7_75t_L g518 ( 
.A(n_448),
.Y(n_518)
);

BUFx6f_ASAP7_75t_L g519 ( 
.A(n_448),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_443),
.Y(n_520)
);

NOR2xp33_ASAP7_75t_L g521 ( 
.A(n_469),
.B(n_438),
.Y(n_521)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_458),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_L g523 ( 
.A(n_499),
.B(n_13),
.Y(n_523)
);

INVx4_ASAP7_75t_L g524 ( 
.A(n_446),
.Y(n_524)
);

AOI21xp5_ASAP7_75t_L g525 ( 
.A1(n_465),
.A2(n_102),
.B(n_188),
.Y(n_525)
);

A2O1A1Ixp33_ASAP7_75t_L g526 ( 
.A1(n_495),
.A2(n_419),
.B(n_16),
.C(n_17),
.Y(n_526)
);

HB1xp67_ASAP7_75t_L g527 ( 
.A(n_498),
.Y(n_527)
);

INVx1_ASAP7_75t_SL g528 ( 
.A(n_498),
.Y(n_528)
);

AOI21xp5_ASAP7_75t_L g529 ( 
.A1(n_488),
.A2(n_100),
.B(n_181),
.Y(n_529)
);

INVx2_ASAP7_75t_L g530 ( 
.A(n_449),
.Y(n_530)
);

NOR3xp33_ASAP7_75t_L g531 ( 
.A(n_493),
.B(n_15),
.C(n_16),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_489),
.B(n_32),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_SL g533 ( 
.A(n_452),
.B(n_33),
.Y(n_533)
);

A2O1A1Ixp33_ASAP7_75t_L g534 ( 
.A1(n_495),
.A2(n_15),
.B(n_18),
.C(n_19),
.Y(n_534)
);

AND2x2_ASAP7_75t_L g535 ( 
.A(n_456),
.B(n_19),
.Y(n_535)
);

AOI21xp5_ASAP7_75t_L g536 ( 
.A1(n_488),
.A2(n_107),
.B(n_34),
.Y(n_536)
);

O2A1O1Ixp33_ASAP7_75t_L g537 ( 
.A1(n_476),
.A2(n_20),
.B(n_35),
.C(n_36),
.Y(n_537)
);

INVx2_ASAP7_75t_L g538 ( 
.A(n_454),
.Y(n_538)
);

AOI22xp33_ASAP7_75t_L g539 ( 
.A1(n_493),
.A2(n_37),
.B1(n_38),
.B2(n_40),
.Y(n_539)
);

AND2x2_ASAP7_75t_SL g540 ( 
.A(n_491),
.B(n_42),
.Y(n_540)
);

AND2x2_ASAP7_75t_L g541 ( 
.A(n_467),
.B(n_43),
.Y(n_541)
);

NOR2xp33_ASAP7_75t_L g542 ( 
.A(n_467),
.B(n_45),
.Y(n_542)
);

AOI22xp33_ASAP7_75t_L g543 ( 
.A1(n_487),
.A2(n_46),
.B1(n_47),
.B2(n_48),
.Y(n_543)
);

CKINVDCx20_ASAP7_75t_R g544 ( 
.A(n_494),
.Y(n_544)
);

AND2x4_ASAP7_75t_L g545 ( 
.A(n_460),
.B(n_50),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_SL g546 ( 
.A(n_511),
.B(n_51),
.Y(n_546)
);

INVx3_ASAP7_75t_L g547 ( 
.A(n_454),
.Y(n_547)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_459),
.Y(n_548)
);

AOI21xp5_ASAP7_75t_L g549 ( 
.A1(n_486),
.A2(n_53),
.B(n_55),
.Y(n_549)
);

AOI21xp5_ASAP7_75t_L g550 ( 
.A1(n_442),
.A2(n_57),
.B(n_58),
.Y(n_550)
);

AOI21xp5_ASAP7_75t_L g551 ( 
.A1(n_501),
.A2(n_59),
.B(n_60),
.Y(n_551)
);

NOR2xp33_ASAP7_75t_L g552 ( 
.A(n_507),
.B(n_62),
.Y(n_552)
);

OAI21x1_ASAP7_75t_L g553 ( 
.A1(n_468),
.A2(n_64),
.B(n_65),
.Y(n_553)
);

NAND3xp33_ASAP7_75t_SL g554 ( 
.A(n_483),
.B(n_490),
.C(n_491),
.Y(n_554)
);

INVx4_ASAP7_75t_L g555 ( 
.A(n_461),
.Y(n_555)
);

NAND2x1_ASAP7_75t_L g556 ( 
.A(n_510),
.B(n_66),
.Y(n_556)
);

OAI21x1_ASAP7_75t_L g557 ( 
.A1(n_484),
.A2(n_183),
.B(n_70),
.Y(n_557)
);

NOR2xp33_ASAP7_75t_SL g558 ( 
.A(n_502),
.B(n_69),
.Y(n_558)
);

INVx2_ASAP7_75t_SL g559 ( 
.A(n_503),
.Y(n_559)
);

OAI22xp5_ASAP7_75t_L g560 ( 
.A1(n_490),
.A2(n_75),
.B1(n_77),
.B2(n_78),
.Y(n_560)
);

AOI21xp5_ASAP7_75t_L g561 ( 
.A1(n_508),
.A2(n_79),
.B(n_80),
.Y(n_561)
);

AND2x4_ASAP7_75t_L g562 ( 
.A(n_451),
.B(n_82),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_461),
.Y(n_563)
);

AOI21xp5_ASAP7_75t_L g564 ( 
.A1(n_472),
.A2(n_83),
.B(n_84),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_SL g565 ( 
.A(n_483),
.B(n_86),
.Y(n_565)
);

O2A1O1Ixp33_ASAP7_75t_L g566 ( 
.A1(n_506),
.A2(n_462),
.B(n_453),
.C(n_464),
.Y(n_566)
);

NOR2xp33_ASAP7_75t_L g567 ( 
.A(n_470),
.B(n_87),
.Y(n_567)
);

INVx2_ASAP7_75t_L g568 ( 
.A(n_471),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_473),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_L g570 ( 
.A(n_463),
.B(n_88),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_L g571 ( 
.A(n_445),
.B(n_90),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_520),
.Y(n_572)
);

INVx5_ASAP7_75t_L g573 ( 
.A(n_524),
.Y(n_573)
);

BUFx8_ASAP7_75t_L g574 ( 
.A(n_518),
.Y(n_574)
);

INVx1_ASAP7_75t_SL g575 ( 
.A(n_528),
.Y(n_575)
);

OAI21x1_ASAP7_75t_L g576 ( 
.A1(n_557),
.A2(n_478),
.B(n_474),
.Y(n_576)
);

OR2x6_ASAP7_75t_L g577 ( 
.A(n_518),
.B(n_450),
.Y(n_577)
);

OAI21x1_ASAP7_75t_L g578 ( 
.A1(n_553),
.A2(n_485),
.B(n_497),
.Y(n_578)
);

INVx8_ASAP7_75t_L g579 ( 
.A(n_518),
.Y(n_579)
);

NAND2x1p5_ASAP7_75t_L g580 ( 
.A(n_540),
.B(n_506),
.Y(n_580)
);

OAI21x1_ASAP7_75t_L g581 ( 
.A1(n_515),
.A2(n_496),
.B(n_505),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_530),
.Y(n_582)
);

OAI21x1_ASAP7_75t_L g583 ( 
.A1(n_550),
.A2(n_492),
.B(n_457),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_568),
.Y(n_584)
);

AOI22x1_ASAP7_75t_L g585 ( 
.A1(n_549),
.A2(n_538),
.B1(n_516),
.B2(n_547),
.Y(n_585)
);

OAI21x1_ASAP7_75t_L g586 ( 
.A1(n_532),
.A2(n_444),
.B(n_477),
.Y(n_586)
);

INVx3_ASAP7_75t_L g587 ( 
.A(n_524),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_569),
.Y(n_588)
);

INVx2_ASAP7_75t_L g589 ( 
.A(n_516),
.Y(n_589)
);

INVxp67_ASAP7_75t_SL g590 ( 
.A(n_547),
.Y(n_590)
);

OAI21xp5_ASAP7_75t_L g591 ( 
.A1(n_532),
.A2(n_444),
.B(n_475),
.Y(n_591)
);

OAI21x1_ASAP7_75t_L g592 ( 
.A1(n_529),
.A2(n_479),
.B(n_500),
.Y(n_592)
);

AO21x2_ASAP7_75t_L g593 ( 
.A1(n_570),
.A2(n_482),
.B(n_466),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_522),
.Y(n_594)
);

OR2x6_ASAP7_75t_L g595 ( 
.A(n_519),
.B(n_481),
.Y(n_595)
);

OAI21x1_ASAP7_75t_L g596 ( 
.A1(n_536),
.A2(n_482),
.B(n_93),
.Y(n_596)
);

OAI21x1_ASAP7_75t_L g597 ( 
.A1(n_556),
.A2(n_91),
.B(n_94),
.Y(n_597)
);

AO21x2_ASAP7_75t_L g598 ( 
.A1(n_554),
.A2(n_565),
.B(n_513),
.Y(n_598)
);

INVx2_ASAP7_75t_R g599 ( 
.A(n_541),
.Y(n_599)
);

AO21x2_ASAP7_75t_L g600 ( 
.A1(n_566),
.A2(n_95),
.B(n_98),
.Y(n_600)
);

OAI21xp5_ASAP7_75t_L g601 ( 
.A1(n_514),
.A2(n_509),
.B(n_504),
.Y(n_601)
);

OAI21x1_ASAP7_75t_L g602 ( 
.A1(n_525),
.A2(n_103),
.B(n_104),
.Y(n_602)
);

INVx1_ASAP7_75t_SL g603 ( 
.A(n_528),
.Y(n_603)
);

BUFx4f_ASAP7_75t_SL g604 ( 
.A(n_544),
.Y(n_604)
);

CKINVDCx6p67_ASAP7_75t_R g605 ( 
.A(n_519),
.Y(n_605)
);

BUFx3_ASAP7_75t_L g606 ( 
.A(n_519),
.Y(n_606)
);

AO21x2_ASAP7_75t_L g607 ( 
.A1(n_571),
.A2(n_108),
.B(n_109),
.Y(n_607)
);

INVx2_ASAP7_75t_SL g608 ( 
.A(n_527),
.Y(n_608)
);

INVx2_ASAP7_75t_L g609 ( 
.A(n_548),
.Y(n_609)
);

BUFx6f_ASAP7_75t_L g610 ( 
.A(n_562),
.Y(n_610)
);

CKINVDCx5p33_ASAP7_75t_R g611 ( 
.A(n_521),
.Y(n_611)
);

AND2x4_ASAP7_75t_L g612 ( 
.A(n_562),
.B(n_111),
.Y(n_612)
);

BUFx2_ASAP7_75t_L g613 ( 
.A(n_545),
.Y(n_613)
);

INVx3_ASAP7_75t_L g614 ( 
.A(n_555),
.Y(n_614)
);

INVx2_ASAP7_75t_SL g615 ( 
.A(n_559),
.Y(n_615)
);

OAI21x1_ASAP7_75t_L g616 ( 
.A1(n_551),
.A2(n_112),
.B(n_113),
.Y(n_616)
);

AND2x2_ASAP7_75t_L g617 ( 
.A(n_512),
.B(n_447),
.Y(n_617)
);

BUFx3_ASAP7_75t_L g618 ( 
.A(n_545),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_563),
.Y(n_619)
);

AOI21xp5_ASAP7_75t_L g620 ( 
.A1(n_567),
.A2(n_114),
.B(n_115),
.Y(n_620)
);

INVx4_ASAP7_75t_L g621 ( 
.A(n_573),
.Y(n_621)
);

OAI21xp5_ASAP7_75t_L g622 ( 
.A1(n_580),
.A2(n_542),
.B(n_560),
.Y(n_622)
);

AND2x4_ASAP7_75t_L g623 ( 
.A(n_610),
.B(n_555),
.Y(n_623)
);

AND2x2_ASAP7_75t_L g624 ( 
.A(n_580),
.B(n_531),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_572),
.Y(n_625)
);

INVx8_ASAP7_75t_L g626 ( 
.A(n_579),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_609),
.Y(n_627)
);

INVx2_ASAP7_75t_L g628 ( 
.A(n_609),
.Y(n_628)
);

OAI22xp5_ASAP7_75t_L g629 ( 
.A1(n_618),
.A2(n_560),
.B1(n_523),
.B2(n_517),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_590),
.Y(n_630)
);

INVx2_ASAP7_75t_L g631 ( 
.A(n_589),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_590),
.Y(n_632)
);

INVx2_ASAP7_75t_SL g633 ( 
.A(n_579),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_L g634 ( 
.A(n_611),
.B(n_552),
.Y(n_634)
);

AND2x2_ASAP7_75t_L g635 ( 
.A(n_598),
.B(n_535),
.Y(n_635)
);

OAI21x1_ASAP7_75t_L g636 ( 
.A1(n_576),
.A2(n_561),
.B(n_564),
.Y(n_636)
);

INVx2_ASAP7_75t_L g637 ( 
.A(n_589),
.Y(n_637)
);

AOI22xp5_ASAP7_75t_SL g638 ( 
.A1(n_611),
.A2(n_534),
.B1(n_558),
.B2(n_526),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_L g639 ( 
.A(n_612),
.B(n_558),
.Y(n_639)
);

CKINVDCx5p33_ASAP7_75t_R g640 ( 
.A(n_604),
.Y(n_640)
);

INVx2_ASAP7_75t_L g641 ( 
.A(n_582),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_584),
.Y(n_642)
);

HB1xp67_ASAP7_75t_L g643 ( 
.A(n_575),
.Y(n_643)
);

OAI22xp5_ASAP7_75t_L g644 ( 
.A1(n_618),
.A2(n_539),
.B1(n_543),
.B2(n_533),
.Y(n_644)
);

INVx3_ASAP7_75t_L g645 ( 
.A(n_573),
.Y(n_645)
);

INVx4_ASAP7_75t_L g646 ( 
.A(n_573),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_588),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_594),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_612),
.B(n_546),
.Y(n_649)
);

AND2x2_ASAP7_75t_L g650 ( 
.A(n_598),
.B(n_537),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_619),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_587),
.Y(n_652)
);

AOI22xp33_ASAP7_75t_L g653 ( 
.A1(n_617),
.A2(n_116),
.B1(n_117),
.B2(n_118),
.Y(n_653)
);

INVx3_ASAP7_75t_L g654 ( 
.A(n_573),
.Y(n_654)
);

INVx2_ASAP7_75t_L g655 ( 
.A(n_587),
.Y(n_655)
);

INVx2_ASAP7_75t_L g656 ( 
.A(n_614),
.Y(n_656)
);

BUFx8_ASAP7_75t_L g657 ( 
.A(n_613),
.Y(n_657)
);

BUFx3_ASAP7_75t_L g658 ( 
.A(n_574),
.Y(n_658)
);

AND2x2_ASAP7_75t_L g659 ( 
.A(n_612),
.B(n_121),
.Y(n_659)
);

AND2x2_ASAP7_75t_L g660 ( 
.A(n_599),
.B(n_122),
.Y(n_660)
);

AND2x2_ASAP7_75t_L g661 ( 
.A(n_599),
.B(n_610),
.Y(n_661)
);

OAI21xp5_ASAP7_75t_L g662 ( 
.A1(n_591),
.A2(n_124),
.B(n_125),
.Y(n_662)
);

OAI22xp33_ASAP7_75t_L g663 ( 
.A1(n_595),
.A2(n_129),
.B1(n_140),
.B2(n_142),
.Y(n_663)
);

NOR2xp33_ASAP7_75t_R g664 ( 
.A(n_640),
.B(n_604),
.Y(n_664)
);

AND2x2_ASAP7_75t_L g665 ( 
.A(n_624),
.B(n_603),
.Y(n_665)
);

AND2x2_ASAP7_75t_L g666 ( 
.A(n_624),
.B(n_634),
.Y(n_666)
);

OAI22xp5_ASAP7_75t_L g667 ( 
.A1(n_622),
.A2(n_610),
.B1(n_601),
.B2(n_595),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_643),
.B(n_610),
.Y(n_668)
);

AND2x4_ASAP7_75t_L g669 ( 
.A(n_658),
.B(n_606),
.Y(n_669)
);

AND2x4_ASAP7_75t_L g670 ( 
.A(n_658),
.B(n_606),
.Y(n_670)
);

AO31x2_ASAP7_75t_L g671 ( 
.A1(n_629),
.A2(n_644),
.A3(n_630),
.B(n_632),
.Y(n_671)
);

BUFx2_ASAP7_75t_R g672 ( 
.A(n_640),
.Y(n_672)
);

HB1xp67_ASAP7_75t_L g673 ( 
.A(n_625),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_639),
.B(n_608),
.Y(n_674)
);

NOR2x1p5_ASAP7_75t_L g675 ( 
.A(n_649),
.B(n_605),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_625),
.Y(n_676)
);

AND2x2_ASAP7_75t_L g677 ( 
.A(n_659),
.B(n_595),
.Y(n_677)
);

AND2x2_ASAP7_75t_L g678 ( 
.A(n_659),
.B(n_615),
.Y(n_678)
);

OR2x2_ASAP7_75t_L g679 ( 
.A(n_641),
.B(n_605),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_642),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_L g681 ( 
.A(n_638),
.B(n_579),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_642),
.Y(n_682)
);

NAND2xp33_ASAP7_75t_R g683 ( 
.A(n_660),
.B(n_577),
.Y(n_683)
);

AOI21x1_ASAP7_75t_L g684 ( 
.A1(n_650),
.A2(n_586),
.B(n_576),
.Y(n_684)
);

AO31x2_ASAP7_75t_L g685 ( 
.A1(n_630),
.A2(n_620),
.A3(n_600),
.B(n_586),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_L g686 ( 
.A(n_638),
.B(n_574),
.Y(n_686)
);

AOI22xp33_ASAP7_75t_SL g687 ( 
.A1(n_662),
.A2(n_574),
.B1(n_593),
.B2(n_600),
.Y(n_687)
);

INVx2_ASAP7_75t_L g688 ( 
.A(n_641),
.Y(n_688)
);

AND2x2_ASAP7_75t_L g689 ( 
.A(n_647),
.B(n_577),
.Y(n_689)
);

OR2x6_ASAP7_75t_L g690 ( 
.A(n_626),
.B(n_577),
.Y(n_690)
);

AND2x2_ASAP7_75t_L g691 ( 
.A(n_647),
.B(n_593),
.Y(n_691)
);

BUFx6f_ASAP7_75t_L g692 ( 
.A(n_626),
.Y(n_692)
);

NOR2xp33_ASAP7_75t_R g693 ( 
.A(n_626),
.B(n_614),
.Y(n_693)
);

BUFx6f_ASAP7_75t_L g694 ( 
.A(n_626),
.Y(n_694)
);

OR2x6_ASAP7_75t_L g695 ( 
.A(n_633),
.B(n_597),
.Y(n_695)
);

HB1xp67_ASAP7_75t_L g696 ( 
.A(n_657),
.Y(n_696)
);

INVxp67_ASAP7_75t_SL g697 ( 
.A(n_632),
.Y(n_697)
);

BUFx3_ASAP7_75t_L g698 ( 
.A(n_657),
.Y(n_698)
);

HB1xp67_ASAP7_75t_L g699 ( 
.A(n_657),
.Y(n_699)
);

BUFx10_ASAP7_75t_L g700 ( 
.A(n_633),
.Y(n_700)
);

NOR2xp33_ASAP7_75t_R g701 ( 
.A(n_645),
.B(n_143),
.Y(n_701)
);

NOR3xp33_ASAP7_75t_SL g702 ( 
.A(n_663),
.B(n_607),
.C(n_596),
.Y(n_702)
);

AO31x2_ASAP7_75t_L g703 ( 
.A1(n_652),
.A2(n_578),
.A3(n_581),
.B(n_583),
.Y(n_703)
);

AND2x2_ASAP7_75t_L g704 ( 
.A(n_648),
.B(n_607),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_648),
.Y(n_705)
);

BUFx6f_ASAP7_75t_L g706 ( 
.A(n_621),
.Y(n_706)
);

AOI22xp33_ASAP7_75t_SL g707 ( 
.A1(n_660),
.A2(n_616),
.B1(n_596),
.B2(n_602),
.Y(n_707)
);

CKINVDCx5p33_ASAP7_75t_R g708 ( 
.A(n_623),
.Y(n_708)
);

AND2x2_ASAP7_75t_L g709 ( 
.A(n_635),
.B(n_597),
.Y(n_709)
);

A2O1A1Ixp33_ASAP7_75t_L g710 ( 
.A1(n_650),
.A2(n_592),
.B(n_616),
.C(n_602),
.Y(n_710)
);

NOR2x1p5_ASAP7_75t_L g711 ( 
.A(n_651),
.B(n_585),
.Y(n_711)
);

AOI21xp5_ASAP7_75t_L g712 ( 
.A1(n_636),
.A2(n_581),
.B(n_583),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_L g713 ( 
.A(n_635),
.B(n_592),
.Y(n_713)
);

INVx2_ASAP7_75t_L g714 ( 
.A(n_676),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_673),
.Y(n_715)
);

INVx2_ASAP7_75t_L g716 ( 
.A(n_680),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_697),
.Y(n_717)
);

AND2x2_ASAP7_75t_L g718 ( 
.A(n_691),
.B(n_661),
.Y(n_718)
);

NOR2x1_ASAP7_75t_L g719 ( 
.A(n_675),
.B(n_646),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_666),
.B(n_651),
.Y(n_720)
);

HB1xp67_ASAP7_75t_L g721 ( 
.A(n_665),
.Y(n_721)
);

AOI22xp33_ASAP7_75t_L g722 ( 
.A1(n_667),
.A2(n_653),
.B1(n_661),
.B2(n_623),
.Y(n_722)
);

OR2x2_ASAP7_75t_L g723 ( 
.A(n_713),
.B(n_627),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_682),
.Y(n_724)
);

AND2x2_ASAP7_75t_L g725 ( 
.A(n_709),
.B(n_631),
.Y(n_725)
);

AND2x4_ASAP7_75t_L g726 ( 
.A(n_705),
.B(n_627),
.Y(n_726)
);

AND2x2_ASAP7_75t_L g727 ( 
.A(n_704),
.B(n_637),
.Y(n_727)
);

OR2x2_ASAP7_75t_L g728 ( 
.A(n_671),
.B(n_628),
.Y(n_728)
);

OAI22xp5_ASAP7_75t_L g729 ( 
.A1(n_686),
.A2(n_623),
.B1(n_652),
.B2(n_646),
.Y(n_729)
);

INVx2_ASAP7_75t_L g730 ( 
.A(n_688),
.Y(n_730)
);

AND2x2_ASAP7_75t_L g731 ( 
.A(n_671),
.B(n_637),
.Y(n_731)
);

BUFx6f_ASAP7_75t_L g732 ( 
.A(n_692),
.Y(n_732)
);

INVx2_ASAP7_75t_L g733 ( 
.A(n_671),
.Y(n_733)
);

INVx3_ASAP7_75t_L g734 ( 
.A(n_695),
.Y(n_734)
);

OR2x2_ASAP7_75t_L g735 ( 
.A(n_681),
.B(n_628),
.Y(n_735)
);

OR2x2_ASAP7_75t_L g736 ( 
.A(n_703),
.B(n_631),
.Y(n_736)
);

AND2x2_ASAP7_75t_L g737 ( 
.A(n_677),
.B(n_656),
.Y(n_737)
);

HB1xp67_ASAP7_75t_L g738 ( 
.A(n_689),
.Y(n_738)
);

OAI33xp33_ASAP7_75t_L g739 ( 
.A1(n_674),
.A2(n_668),
.A3(n_679),
.B1(n_708),
.B2(n_656),
.B3(n_655),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_711),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_703),
.Y(n_741)
);

OR2x2_ASAP7_75t_L g742 ( 
.A(n_703),
.B(n_685),
.Y(n_742)
);

INVx2_ASAP7_75t_L g743 ( 
.A(n_684),
.Y(n_743)
);

HB1xp67_ASAP7_75t_L g744 ( 
.A(n_683),
.Y(n_744)
);

INVx2_ASAP7_75t_SL g745 ( 
.A(n_700),
.Y(n_745)
);

AND2x2_ASAP7_75t_L g746 ( 
.A(n_678),
.B(n_655),
.Y(n_746)
);

OR2x2_ASAP7_75t_L g747 ( 
.A(n_685),
.B(n_636),
.Y(n_747)
);

AND2x4_ASAP7_75t_L g748 ( 
.A(n_692),
.B(n_654),
.Y(n_748)
);

AND2x2_ASAP7_75t_L g749 ( 
.A(n_685),
.B(n_687),
.Y(n_749)
);

AOI21xp5_ASAP7_75t_L g750 ( 
.A1(n_712),
.A2(n_646),
.B(n_621),
.Y(n_750)
);

INVx2_ASAP7_75t_L g751 ( 
.A(n_695),
.Y(n_751)
);

HB1xp67_ASAP7_75t_L g752 ( 
.A(n_690),
.Y(n_752)
);

INVx2_ASAP7_75t_L g753 ( 
.A(n_706),
.Y(n_753)
);

AND2x2_ASAP7_75t_L g754 ( 
.A(n_710),
.B(n_654),
.Y(n_754)
);

INVx2_ASAP7_75t_L g755 ( 
.A(n_706),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_700),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_720),
.B(n_670),
.Y(n_757)
);

INVx2_ASAP7_75t_L g758 ( 
.A(n_714),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_724),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_715),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_714),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_716),
.Y(n_762)
);

OAI211xp5_ASAP7_75t_L g763 ( 
.A1(n_740),
.A2(n_701),
.B(n_702),
.C(n_707),
.Y(n_763)
);

AND2x2_ASAP7_75t_L g764 ( 
.A(n_718),
.B(n_749),
.Y(n_764)
);

AND2x2_ASAP7_75t_L g765 ( 
.A(n_718),
.B(n_699),
.Y(n_765)
);

AND2x2_ASAP7_75t_L g766 ( 
.A(n_738),
.B(n_669),
.Y(n_766)
);

AND2x4_ASAP7_75t_L g767 ( 
.A(n_751),
.B(n_670),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_716),
.Y(n_768)
);

OAI21xp5_ASAP7_75t_SL g769 ( 
.A1(n_744),
.A2(n_696),
.B(n_669),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_L g770 ( 
.A(n_721),
.B(n_698),
.Y(n_770)
);

INVx2_ASAP7_75t_SL g771 ( 
.A(n_751),
.Y(n_771)
);

OR2x2_ASAP7_75t_L g772 ( 
.A(n_723),
.B(n_690),
.Y(n_772)
);

INVxp67_ASAP7_75t_L g773 ( 
.A(n_746),
.Y(n_773)
);

AOI22xp33_ASAP7_75t_L g774 ( 
.A1(n_739),
.A2(n_664),
.B1(n_694),
.B2(n_692),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_735),
.B(n_706),
.Y(n_775)
);

OAI22xp5_ASAP7_75t_L g776 ( 
.A1(n_722),
.A2(n_672),
.B1(n_694),
.B2(n_621),
.Y(n_776)
);

AND2x2_ASAP7_75t_L g777 ( 
.A(n_749),
.B(n_578),
.Y(n_777)
);

AND2x2_ASAP7_75t_L g778 ( 
.A(n_727),
.B(n_654),
.Y(n_778)
);

AND2x2_ASAP7_75t_L g779 ( 
.A(n_727),
.B(n_645),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_717),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_736),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_L g782 ( 
.A(n_735),
.B(n_694),
.Y(n_782)
);

AND2x2_ASAP7_75t_L g783 ( 
.A(n_764),
.B(n_734),
.Y(n_783)
);

AND2x4_ASAP7_75t_L g784 ( 
.A(n_771),
.B(n_734),
.Y(n_784)
);

INVx2_ASAP7_75t_L g785 ( 
.A(n_758),
.Y(n_785)
);

AND2x2_ASAP7_75t_L g786 ( 
.A(n_764),
.B(n_734),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_759),
.Y(n_787)
);

OR2x2_ASAP7_75t_L g788 ( 
.A(n_781),
.B(n_742),
.Y(n_788)
);

INVx1_ASAP7_75t_SL g789 ( 
.A(n_770),
.Y(n_789)
);

NOR2x1_ASAP7_75t_L g790 ( 
.A(n_769),
.B(n_756),
.Y(n_790)
);

AND2x2_ASAP7_75t_L g791 ( 
.A(n_777),
.B(n_733),
.Y(n_791)
);

AND2x2_ASAP7_75t_L g792 ( 
.A(n_777),
.B(n_733),
.Y(n_792)
);

INVx2_ASAP7_75t_L g793 ( 
.A(n_758),
.Y(n_793)
);

HB1xp67_ASAP7_75t_L g794 ( 
.A(n_771),
.Y(n_794)
);

AND2x2_ASAP7_75t_L g795 ( 
.A(n_765),
.B(n_754),
.Y(n_795)
);

AND2x4_ASAP7_75t_L g796 ( 
.A(n_767),
.B(n_754),
.Y(n_796)
);

AND2x4_ASAP7_75t_L g797 ( 
.A(n_767),
.B(n_731),
.Y(n_797)
);

INVxp67_ASAP7_75t_L g798 ( 
.A(n_765),
.Y(n_798)
);

OR2x2_ASAP7_75t_L g799 ( 
.A(n_798),
.B(n_783),
.Y(n_799)
);

INVx2_ASAP7_75t_L g800 ( 
.A(n_785),
.Y(n_800)
);

OAI22xp33_ASAP7_75t_L g801 ( 
.A1(n_790),
.A2(n_776),
.B1(n_772),
.B2(n_729),
.Y(n_801)
);

OAI22xp5_ASAP7_75t_L g802 ( 
.A1(n_789),
.A2(n_774),
.B1(n_763),
.B2(n_752),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_L g803 ( 
.A(n_795),
.B(n_760),
.Y(n_803)
);

OA222x2_ASAP7_75t_L g804 ( 
.A1(n_788),
.A2(n_728),
.B1(n_742),
.B2(n_780),
.C1(n_762),
.C2(n_768),
.Y(n_804)
);

AOI22xp5_ASAP7_75t_L g805 ( 
.A1(n_796),
.A2(n_774),
.B1(n_767),
.B2(n_773),
.Y(n_805)
);

INVxp67_ASAP7_75t_L g806 ( 
.A(n_794),
.Y(n_806)
);

OAI32xp33_ASAP7_75t_L g807 ( 
.A1(n_788),
.A2(n_757),
.A3(n_782),
.B1(n_775),
.B2(n_761),
.Y(n_807)
);

OAI22xp33_ASAP7_75t_L g808 ( 
.A1(n_787),
.A2(n_723),
.B1(n_753),
.B2(n_755),
.Y(n_808)
);

AOI22xp33_ASAP7_75t_SL g809 ( 
.A1(n_802),
.A2(n_796),
.B1(n_795),
.B2(n_797),
.Y(n_809)
);

AO21x1_ASAP7_75t_L g810 ( 
.A1(n_801),
.A2(n_784),
.B(n_796),
.Y(n_810)
);

CKINVDCx16_ASAP7_75t_R g811 ( 
.A(n_805),
.Y(n_811)
);

BUFx3_ASAP7_75t_L g812 ( 
.A(n_803),
.Y(n_812)
);

OAI221xp5_ASAP7_75t_L g813 ( 
.A1(n_806),
.A2(n_745),
.B1(n_719),
.B2(n_766),
.C(n_785),
.Y(n_813)
);

AOI22xp5_ASAP7_75t_L g814 ( 
.A1(n_810),
.A2(n_808),
.B1(n_797),
.B2(n_783),
.Y(n_814)
);

AOI21xp33_ASAP7_75t_SL g815 ( 
.A1(n_811),
.A2(n_807),
.B(n_745),
.Y(n_815)
);

INVxp33_ASAP7_75t_L g816 ( 
.A(n_809),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_812),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_813),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_L g819 ( 
.A(n_812),
.B(n_786),
.Y(n_819)
);

NOR3x1_ASAP7_75t_L g820 ( 
.A(n_818),
.B(n_804),
.C(n_799),
.Y(n_820)
);

OAI22xp5_ASAP7_75t_L g821 ( 
.A1(n_816),
.A2(n_797),
.B1(n_786),
.B2(n_784),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_L g822 ( 
.A(n_817),
.B(n_800),
.Y(n_822)
);

HB1xp67_ASAP7_75t_L g823 ( 
.A(n_819),
.Y(n_823)
);

AOI22xp5_ASAP7_75t_L g824 ( 
.A1(n_821),
.A2(n_814),
.B1(n_784),
.B2(n_778),
.Y(n_824)
);

NOR2x1_ASAP7_75t_L g825 ( 
.A(n_822),
.B(n_815),
.Y(n_825)
);

NOR2x1_ASAP7_75t_L g826 ( 
.A(n_825),
.B(n_820),
.Y(n_826)
);

AOI21xp33_ASAP7_75t_L g827 ( 
.A1(n_824),
.A2(n_823),
.B(n_753),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_825),
.Y(n_828)
);

INVx2_ASAP7_75t_L g829 ( 
.A(n_828),
.Y(n_829)
);

AOI22xp33_ASAP7_75t_L g830 ( 
.A1(n_826),
.A2(n_779),
.B1(n_778),
.B2(n_748),
.Y(n_830)
);

NOR2xp33_ASAP7_75t_L g831 ( 
.A(n_827),
.B(n_746),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_828),
.Y(n_832)
);

INVxp67_ASAP7_75t_SL g833 ( 
.A(n_828),
.Y(n_833)
);

HB1xp67_ASAP7_75t_L g834 ( 
.A(n_828),
.Y(n_834)
);

OAI22xp5_ASAP7_75t_L g835 ( 
.A1(n_830),
.A2(n_793),
.B1(n_792),
.B2(n_791),
.Y(n_835)
);

NAND4xp25_ASAP7_75t_L g836 ( 
.A(n_832),
.B(n_755),
.C(n_737),
.D(n_748),
.Y(n_836)
);

OR2x2_ASAP7_75t_L g837 ( 
.A(n_829),
.B(n_793),
.Y(n_837)
);

NAND3xp33_ASAP7_75t_L g838 ( 
.A(n_834),
.B(n_732),
.C(n_750),
.Y(n_838)
);

NOR3xp33_ASAP7_75t_L g839 ( 
.A(n_833),
.B(n_737),
.C(n_748),
.Y(n_839)
);

AND4x2_ASAP7_75t_L g840 ( 
.A(n_834),
.B(n_732),
.C(n_693),
.D(n_149),
.Y(n_840)
);

INVx2_ASAP7_75t_L g841 ( 
.A(n_831),
.Y(n_841)
);

OAI22xp5_ASAP7_75t_L g842 ( 
.A1(n_841),
.A2(n_732),
.B1(n_791),
.B2(n_792),
.Y(n_842)
);

AND2x2_ASAP7_75t_L g843 ( 
.A(n_839),
.B(n_779),
.Y(n_843)
);

AOI22xp5_ASAP7_75t_L g844 ( 
.A1(n_836),
.A2(n_732),
.B1(n_726),
.B2(n_731),
.Y(n_844)
);

HB1xp67_ASAP7_75t_L g845 ( 
.A(n_837),
.Y(n_845)
);

NAND4xp75_ASAP7_75t_L g846 ( 
.A(n_840),
.B(n_838),
.C(n_835),
.D(n_741),
.Y(n_846)
);

BUFx2_ASAP7_75t_L g847 ( 
.A(n_841),
.Y(n_847)
);

INVx1_ASAP7_75t_SL g848 ( 
.A(n_837),
.Y(n_848)
);

CKINVDCx20_ASAP7_75t_R g849 ( 
.A(n_847),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_848),
.B(n_845),
.Y(n_850)
);

INVx2_ASAP7_75t_L g851 ( 
.A(n_843),
.Y(n_851)
);

INVx3_ASAP7_75t_L g852 ( 
.A(n_846),
.Y(n_852)
);

NAND2x1_ASAP7_75t_L g853 ( 
.A(n_842),
.B(n_645),
.Y(n_853)
);

OAI22xp5_ASAP7_75t_L g854 ( 
.A1(n_844),
.A2(n_728),
.B1(n_747),
.B2(n_726),
.Y(n_854)
);

CKINVDCx20_ASAP7_75t_R g855 ( 
.A(n_847),
.Y(n_855)
);

OA22x2_ASAP7_75t_L g856 ( 
.A1(n_848),
.A2(n_726),
.B1(n_730),
.B2(n_743),
.Y(n_856)
);

INVx2_ASAP7_75t_L g857 ( 
.A(n_847),
.Y(n_857)
);

OAI31xp33_ASAP7_75t_L g858 ( 
.A1(n_857),
.A2(n_747),
.A3(n_730),
.B(n_743),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_849),
.Y(n_859)
);

OAI31xp33_ASAP7_75t_L g860 ( 
.A1(n_850),
.A2(n_725),
.A3(n_736),
.B(n_151),
.Y(n_860)
);

OAI22xp33_ASAP7_75t_L g861 ( 
.A1(n_855),
.A2(n_725),
.B1(n_147),
.B2(n_152),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_852),
.B(n_144),
.Y(n_862)
);

AOI22xp5_ASAP7_75t_L g863 ( 
.A1(n_851),
.A2(n_155),
.B1(n_157),
.B2(n_161),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_856),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_853),
.B(n_162),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_854),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_859),
.B(n_164),
.Y(n_867)
);

XNOR2x1_ASAP7_75t_L g868 ( 
.A(n_862),
.B(n_165),
.Y(n_868)
);

BUFx2_ASAP7_75t_L g869 ( 
.A(n_865),
.Y(n_869)
);

AND2x2_ASAP7_75t_L g870 ( 
.A(n_866),
.B(n_166),
.Y(n_870)
);

CKINVDCx20_ASAP7_75t_R g871 ( 
.A(n_869),
.Y(n_871)
);

AND2x2_ASAP7_75t_L g872 ( 
.A(n_870),
.B(n_864),
.Y(n_872)
);

OAI21xp5_ASAP7_75t_L g873 ( 
.A1(n_872),
.A2(n_871),
.B(n_867),
.Y(n_873)
);

AOI22xp5_ASAP7_75t_L g874 ( 
.A1(n_873),
.A2(n_868),
.B1(n_861),
.B2(n_863),
.Y(n_874)
);

AOI22xp33_ASAP7_75t_SL g875 ( 
.A1(n_874),
.A2(n_860),
.B1(n_858),
.B2(n_170),
.Y(n_875)
);

AOI22xp33_ASAP7_75t_L g876 ( 
.A1(n_875),
.A2(n_167),
.B1(n_169),
.B2(n_172),
.Y(n_876)
);


endmodule