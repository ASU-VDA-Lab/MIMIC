module fake_netlist_1_7940_n_716 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_716);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_716;
wire n_117;
wire n_663;
wire n_707;
wire n_361;
wire n_513;
wire n_185;
wire n_705;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_701;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_715;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_563;
wire n_540;
wire n_638;
wire n_141;
wire n_119;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_712;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_85;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_711;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_708;
wire n_307;
wire n_191;
wire n_634;
wire n_610;
wire n_696;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_699;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_704;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_706;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_90;
wire n_357;
wire n_653;
wire n_260;
wire n_539;
wire n_201;
wire n_197;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_363;
wire n_409;
wire n_315;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_684;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_714;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_618;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_266;
wire n_84;
wire n_683;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_337;
wire n_159;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_695;
wire n_469;
wire n_585;
wire n_713;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_709;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_109;
wire n_132;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
CKINVDCx16_ASAP7_75t_R g80 ( .A(n_56), .Y(n_80) );
INVx1_ASAP7_75t_L g81 ( .A(n_65), .Y(n_81) );
INVx2_ASAP7_75t_L g82 ( .A(n_54), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_38), .Y(n_83) );
CKINVDCx20_ASAP7_75t_R g84 ( .A(n_15), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_74), .Y(n_85) );
INVxp33_ASAP7_75t_L g86 ( .A(n_15), .Y(n_86) );
INVxp33_ASAP7_75t_SL g87 ( .A(n_51), .Y(n_87) );
INVxp33_ASAP7_75t_SL g88 ( .A(n_57), .Y(n_88) );
INVxp33_ASAP7_75t_SL g89 ( .A(n_14), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_77), .Y(n_90) );
INVxp33_ASAP7_75t_L g91 ( .A(n_22), .Y(n_91) );
INVxp67_ASAP7_75t_SL g92 ( .A(n_41), .Y(n_92) );
INVxp33_ASAP7_75t_SL g93 ( .A(n_21), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_59), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_78), .Y(n_95) );
INVxp67_ASAP7_75t_L g96 ( .A(n_0), .Y(n_96) );
CKINVDCx16_ASAP7_75t_R g97 ( .A(n_39), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_48), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_20), .Y(n_99) );
HB1xp67_ASAP7_75t_L g100 ( .A(n_60), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_12), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_46), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_21), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_34), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_68), .Y(n_105) );
INVxp33_ASAP7_75t_SL g106 ( .A(n_50), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_7), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_70), .Y(n_108) );
NOR2xp67_ASAP7_75t_L g109 ( .A(n_5), .B(n_4), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_73), .Y(n_110) );
INVx2_ASAP7_75t_L g111 ( .A(n_58), .Y(n_111) );
INVxp67_ASAP7_75t_SL g112 ( .A(n_20), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_40), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_72), .Y(n_114) );
INVxp67_ASAP7_75t_SL g115 ( .A(n_11), .Y(n_115) );
BUFx3_ASAP7_75t_L g116 ( .A(n_29), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_79), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_24), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_1), .Y(n_119) );
CKINVDCx5p33_ASAP7_75t_R g120 ( .A(n_6), .Y(n_120) );
CKINVDCx5p33_ASAP7_75t_R g121 ( .A(n_32), .Y(n_121) );
CKINVDCx20_ASAP7_75t_R g122 ( .A(n_18), .Y(n_122) );
BUFx6f_ASAP7_75t_L g123 ( .A(n_11), .Y(n_123) );
BUFx6f_ASAP7_75t_L g124 ( .A(n_18), .Y(n_124) );
INVxp67_ASAP7_75t_SL g125 ( .A(n_0), .Y(n_125) );
BUFx10_ASAP7_75t_L g126 ( .A(n_26), .Y(n_126) );
CKINVDCx16_ASAP7_75t_R g127 ( .A(n_17), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_49), .Y(n_128) );
INVx1_ASAP7_75t_L g129 ( .A(n_81), .Y(n_129) );
BUFx8_ASAP7_75t_L g130 ( .A(n_82), .Y(n_130) );
NAND2xp5_ASAP7_75t_L g131 ( .A(n_100), .B(n_1), .Y(n_131) );
NAND2xp33_ASAP7_75t_SL g132 ( .A(n_86), .B(n_2), .Y(n_132) );
INVx3_ASAP7_75t_L g133 ( .A(n_126), .Y(n_133) );
BUFx2_ASAP7_75t_L g134 ( .A(n_127), .Y(n_134) );
AND2x2_ASAP7_75t_L g135 ( .A(n_91), .B(n_2), .Y(n_135) );
BUFx6f_ASAP7_75t_L g136 ( .A(n_116), .Y(n_136) );
INVx1_ASAP7_75t_L g137 ( .A(n_81), .Y(n_137) );
INVx1_ASAP7_75t_L g138 ( .A(n_83), .Y(n_138) );
INVx3_ASAP7_75t_L g139 ( .A(n_126), .Y(n_139) );
INVx1_ASAP7_75t_L g140 ( .A(n_83), .Y(n_140) );
HB1xp67_ASAP7_75t_L g141 ( .A(n_99), .Y(n_141) );
INVx1_ASAP7_75t_L g142 ( .A(n_85), .Y(n_142) );
INVx2_ASAP7_75t_L g143 ( .A(n_82), .Y(n_143) );
INVx1_ASAP7_75t_L g144 ( .A(n_85), .Y(n_144) );
INVx1_ASAP7_75t_L g145 ( .A(n_90), .Y(n_145) );
NAND2xp5_ASAP7_75t_L g146 ( .A(n_99), .B(n_3), .Y(n_146) );
AND2x4_ASAP7_75t_L g147 ( .A(n_101), .B(n_3), .Y(n_147) );
INVx1_ASAP7_75t_L g148 ( .A(n_90), .Y(n_148) );
INVx2_ASAP7_75t_L g149 ( .A(n_111), .Y(n_149) );
INVx3_ASAP7_75t_L g150 ( .A(n_126), .Y(n_150) );
AND2x2_ASAP7_75t_L g151 ( .A(n_80), .B(n_4), .Y(n_151) );
OA21x2_ASAP7_75t_L g152 ( .A1(n_94), .A2(n_36), .B(n_75), .Y(n_152) );
AND2x2_ASAP7_75t_L g153 ( .A(n_97), .B(n_5), .Y(n_153) );
HB1xp67_ASAP7_75t_L g154 ( .A(n_101), .Y(n_154) );
INVx2_ASAP7_75t_L g155 ( .A(n_111), .Y(n_155) );
AND2x6_ASAP7_75t_L g156 ( .A(n_116), .B(n_35), .Y(n_156) );
INVx2_ASAP7_75t_L g157 ( .A(n_94), .Y(n_157) );
BUFx6f_ASAP7_75t_L g158 ( .A(n_123), .Y(n_158) );
BUFx6f_ASAP7_75t_L g159 ( .A(n_123), .Y(n_159) );
AND2x2_ASAP7_75t_L g160 ( .A(n_103), .B(n_6), .Y(n_160) );
INVx2_ASAP7_75t_L g161 ( .A(n_95), .Y(n_161) );
BUFx6f_ASAP7_75t_L g162 ( .A(n_123), .Y(n_162) );
NAND2xp5_ASAP7_75t_L g163 ( .A(n_103), .B(n_7), .Y(n_163) );
INVx1_ASAP7_75t_L g164 ( .A(n_95), .Y(n_164) );
BUFx2_ASAP7_75t_L g165 ( .A(n_120), .Y(n_165) );
INVx3_ASAP7_75t_L g166 ( .A(n_123), .Y(n_166) );
INVx2_ASAP7_75t_L g167 ( .A(n_98), .Y(n_167) );
INVx1_ASAP7_75t_L g168 ( .A(n_98), .Y(n_168) );
HB1xp67_ASAP7_75t_L g169 ( .A(n_107), .Y(n_169) );
BUFx6f_ASAP7_75t_L g170 ( .A(n_123), .Y(n_170) );
NAND2xp33_ASAP7_75t_L g171 ( .A(n_121), .B(n_42), .Y(n_171) );
INVx1_ASAP7_75t_L g172 ( .A(n_102), .Y(n_172) );
NAND2xp5_ASAP7_75t_L g173 ( .A(n_139), .B(n_96), .Y(n_173) );
BUFx3_ASAP7_75t_L g174 ( .A(n_136), .Y(n_174) );
AND2x4_ASAP7_75t_L g175 ( .A(n_139), .B(n_107), .Y(n_175) );
AND2x2_ASAP7_75t_L g176 ( .A(n_141), .B(n_119), .Y(n_176) );
NAND2xp5_ASAP7_75t_L g177 ( .A(n_139), .B(n_128), .Y(n_177) );
INVx1_ASAP7_75t_L g178 ( .A(n_157), .Y(n_178) );
INVx1_ASAP7_75t_L g179 ( .A(n_157), .Y(n_179) );
INVx1_ASAP7_75t_L g180 ( .A(n_157), .Y(n_180) );
INVx1_ASAP7_75t_L g181 ( .A(n_161), .Y(n_181) );
NOR2xp33_ASAP7_75t_L g182 ( .A(n_133), .B(n_106), .Y(n_182) );
NAND2xp5_ASAP7_75t_L g183 ( .A(n_139), .B(n_128), .Y(n_183) );
BUFx6f_ASAP7_75t_L g184 ( .A(n_158), .Y(n_184) );
NAND2xp5_ASAP7_75t_L g185 ( .A(n_139), .B(n_114), .Y(n_185) );
INVx2_ASAP7_75t_L g186 ( .A(n_136), .Y(n_186) );
INVx1_ASAP7_75t_L g187 ( .A(n_161), .Y(n_187) );
AND2x4_ASAP7_75t_L g188 ( .A(n_150), .B(n_119), .Y(n_188) );
NAND2xp5_ASAP7_75t_L g189 ( .A(n_150), .B(n_113), .Y(n_189) );
NOR2xp33_ASAP7_75t_L g190 ( .A(n_133), .B(n_87), .Y(n_190) );
BUFx6f_ASAP7_75t_L g191 ( .A(n_158), .Y(n_191) );
AND2x2_ASAP7_75t_L g192 ( .A(n_141), .B(n_125), .Y(n_192) );
AND2x6_ASAP7_75t_L g193 ( .A(n_147), .B(n_108), .Y(n_193) );
BUFx6f_ASAP7_75t_L g194 ( .A(n_158), .Y(n_194) );
NAND2xp5_ASAP7_75t_SL g195 ( .A(n_150), .B(n_88), .Y(n_195) );
INVx1_ASAP7_75t_L g196 ( .A(n_161), .Y(n_196) );
BUFx3_ASAP7_75t_L g197 ( .A(n_136), .Y(n_197) );
OR2x2_ASAP7_75t_L g198 ( .A(n_134), .B(n_112), .Y(n_198) );
INVx3_ASAP7_75t_L g199 ( .A(n_147), .Y(n_199) );
INVx2_ASAP7_75t_L g200 ( .A(n_136), .Y(n_200) );
NOR2xp33_ASAP7_75t_L g201 ( .A(n_133), .B(n_93), .Y(n_201) );
AND2x4_ASAP7_75t_L g202 ( .A(n_150), .B(n_109), .Y(n_202) );
INVx2_ASAP7_75t_L g203 ( .A(n_136), .Y(n_203) );
INVx1_ASAP7_75t_L g204 ( .A(n_167), .Y(n_204) );
INVx4_ASAP7_75t_L g205 ( .A(n_156), .Y(n_205) );
AND2x4_ASAP7_75t_L g206 ( .A(n_150), .B(n_110), .Y(n_206) );
NAND2xp5_ASAP7_75t_L g207 ( .A(n_133), .B(n_110), .Y(n_207) );
INVxp67_ASAP7_75t_L g208 ( .A(n_134), .Y(n_208) );
INVx1_ASAP7_75t_L g209 ( .A(n_167), .Y(n_209) );
AND2x2_ASAP7_75t_L g210 ( .A(n_154), .B(n_115), .Y(n_210) );
AND2x6_ASAP7_75t_L g211 ( .A(n_147), .B(n_108), .Y(n_211) );
NOR2xp33_ASAP7_75t_L g212 ( .A(n_165), .B(n_89), .Y(n_212) );
AND2x4_ASAP7_75t_L g213 ( .A(n_154), .B(n_113), .Y(n_213) );
NOR2xp33_ASAP7_75t_L g214 ( .A(n_165), .B(n_105), .Y(n_214) );
BUFx2_ASAP7_75t_L g215 ( .A(n_151), .Y(n_215) );
INVx1_ASAP7_75t_L g216 ( .A(n_167), .Y(n_216) );
AOI22xp33_ASAP7_75t_L g217 ( .A1(n_147), .A2(n_124), .B1(n_105), .B2(n_118), .Y(n_217) );
AND2x6_ASAP7_75t_L g218 ( .A(n_147), .B(n_118), .Y(n_218) );
BUFx3_ASAP7_75t_L g219 ( .A(n_136), .Y(n_219) );
INVx1_ASAP7_75t_L g220 ( .A(n_143), .Y(n_220) );
HB1xp67_ASAP7_75t_L g221 ( .A(n_151), .Y(n_221) );
AND2x4_ASAP7_75t_L g222 ( .A(n_169), .B(n_117), .Y(n_222) );
NAND2xp5_ASAP7_75t_L g223 ( .A(n_135), .B(n_104), .Y(n_223) );
INVx3_ASAP7_75t_L g224 ( .A(n_143), .Y(n_224) );
NAND2x1p5_ASAP7_75t_L g225 ( .A(n_160), .B(n_117), .Y(n_225) );
INVx2_ASAP7_75t_L g226 ( .A(n_136), .Y(n_226) );
INVx2_ASAP7_75t_SL g227 ( .A(n_130), .Y(n_227) );
NAND2xp5_ASAP7_75t_SL g228 ( .A(n_130), .B(n_114), .Y(n_228) );
NAND2xp5_ASAP7_75t_SL g229 ( .A(n_130), .B(n_104), .Y(n_229) );
INVx2_ASAP7_75t_L g230 ( .A(n_158), .Y(n_230) );
INVx4_ASAP7_75t_L g231 ( .A(n_156), .Y(n_231) );
BUFx3_ASAP7_75t_L g232 ( .A(n_130), .Y(n_232) );
INVx1_ASAP7_75t_L g233 ( .A(n_143), .Y(n_233) );
NAND2xp5_ASAP7_75t_SL g234 ( .A(n_130), .B(n_102), .Y(n_234) );
INVx1_ASAP7_75t_L g235 ( .A(n_149), .Y(n_235) );
INVx2_ASAP7_75t_L g236 ( .A(n_158), .Y(n_236) );
INVx1_ASAP7_75t_L g237 ( .A(n_149), .Y(n_237) );
HB1xp67_ASAP7_75t_L g238 ( .A(n_151), .Y(n_238) );
AND2x2_ASAP7_75t_L g239 ( .A(n_169), .B(n_124), .Y(n_239) );
INVxp67_ASAP7_75t_L g240 ( .A(n_221), .Y(n_240) );
AOI22xp33_ASAP7_75t_L g241 ( .A1(n_193), .A2(n_172), .B1(n_148), .B2(n_140), .Y(n_241) );
BUFx6f_ASAP7_75t_L g242 ( .A(n_232), .Y(n_242) );
NAND2xp5_ASAP7_75t_L g243 ( .A(n_213), .B(n_135), .Y(n_243) );
INVx1_ASAP7_75t_L g244 ( .A(n_239), .Y(n_244) );
INVx1_ASAP7_75t_L g245 ( .A(n_239), .Y(n_245) );
INVx2_ASAP7_75t_SL g246 ( .A(n_213), .Y(n_246) );
NAND2xp5_ASAP7_75t_L g247 ( .A(n_213), .B(n_135), .Y(n_247) );
INVx2_ASAP7_75t_L g248 ( .A(n_178), .Y(n_248) );
HB1xp67_ASAP7_75t_L g249 ( .A(n_222), .Y(n_249) );
NOR2x1_ASAP7_75t_L g250 ( .A(n_198), .B(n_131), .Y(n_250) );
AOI22xp33_ASAP7_75t_L g251 ( .A1(n_193), .A2(n_172), .B1(n_129), .B2(n_137), .Y(n_251) );
BUFx6f_ASAP7_75t_L g252 ( .A(n_232), .Y(n_252) );
INVx1_ASAP7_75t_L g253 ( .A(n_175), .Y(n_253) );
NAND2xp5_ASAP7_75t_L g254 ( .A(n_222), .B(n_153), .Y(n_254) );
INVx4_ASAP7_75t_L g255 ( .A(n_193), .Y(n_255) );
INVx1_ASAP7_75t_L g256 ( .A(n_175), .Y(n_256) );
INVx1_ASAP7_75t_L g257 ( .A(n_175), .Y(n_257) );
NAND2xp5_ASAP7_75t_L g258 ( .A(n_222), .B(n_153), .Y(n_258) );
INVx1_ASAP7_75t_L g259 ( .A(n_188), .Y(n_259) );
AND2x2_ASAP7_75t_L g260 ( .A(n_215), .B(n_153), .Y(n_260) );
INVx3_ASAP7_75t_L g261 ( .A(n_188), .Y(n_261) );
INVx1_ASAP7_75t_L g262 ( .A(n_188), .Y(n_262) );
INVxp67_ASAP7_75t_L g263 ( .A(n_238), .Y(n_263) );
BUFx2_ASAP7_75t_L g264 ( .A(n_208), .Y(n_264) );
INVx2_ASAP7_75t_L g265 ( .A(n_178), .Y(n_265) );
INVx4_ASAP7_75t_L g266 ( .A(n_193), .Y(n_266) );
AND2x4_ASAP7_75t_L g267 ( .A(n_176), .B(n_160), .Y(n_267) );
BUFx4f_ASAP7_75t_L g268 ( .A(n_225), .Y(n_268) );
OR2x6_ASAP7_75t_L g269 ( .A(n_215), .B(n_131), .Y(n_269) );
BUFx2_ASAP7_75t_L g270 ( .A(n_198), .Y(n_270) );
OR2x6_ASAP7_75t_L g271 ( .A(n_225), .B(n_160), .Y(n_271) );
AOI21xp5_ASAP7_75t_L g272 ( .A1(n_228), .A2(n_152), .B(n_171), .Y(n_272) );
INVx1_ASAP7_75t_L g273 ( .A(n_225), .Y(n_273) );
HB1xp67_ASAP7_75t_L g274 ( .A(n_176), .Y(n_274) );
INVx1_ASAP7_75t_L g275 ( .A(n_179), .Y(n_275) );
NAND2xp5_ASAP7_75t_L g276 ( .A(n_223), .B(n_137), .Y(n_276) );
INVx1_ASAP7_75t_SL g277 ( .A(n_192), .Y(n_277) );
INVx1_ASAP7_75t_L g278 ( .A(n_179), .Y(n_278) );
INVx1_ASAP7_75t_L g279 ( .A(n_180), .Y(n_279) );
INVx2_ASAP7_75t_L g280 ( .A(n_180), .Y(n_280) );
O2A1O1Ixp33_ASAP7_75t_L g281 ( .A1(n_192), .A2(n_163), .B(n_146), .C(n_148), .Y(n_281) );
NAND2xp5_ASAP7_75t_SL g282 ( .A(n_227), .B(n_205), .Y(n_282) );
NAND2xp5_ASAP7_75t_L g283 ( .A(n_206), .B(n_138), .Y(n_283) );
NOR2x1_ASAP7_75t_L g284 ( .A(n_212), .B(n_146), .Y(n_284) );
AND2x4_ASAP7_75t_L g285 ( .A(n_202), .B(n_163), .Y(n_285) );
BUFx6f_ASAP7_75t_L g286 ( .A(n_227), .Y(n_286) );
AND2x4_ASAP7_75t_L g287 ( .A(n_202), .B(n_142), .Y(n_287) );
INVx1_ASAP7_75t_L g288 ( .A(n_181), .Y(n_288) );
CKINVDCx5p33_ASAP7_75t_R g289 ( .A(n_210), .Y(n_289) );
INVx2_ASAP7_75t_L g290 ( .A(n_181), .Y(n_290) );
NAND2xp5_ASAP7_75t_L g291 ( .A(n_206), .B(n_145), .Y(n_291) );
INVx1_ASAP7_75t_L g292 ( .A(n_187), .Y(n_292) );
INVx2_ASAP7_75t_L g293 ( .A(n_187), .Y(n_293) );
INVx1_ASAP7_75t_SL g294 ( .A(n_210), .Y(n_294) );
BUFx6f_ASAP7_75t_L g295 ( .A(n_205), .Y(n_295) );
AND2x4_ASAP7_75t_L g296 ( .A(n_202), .B(n_142), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g297 ( .A(n_206), .B(n_138), .Y(n_297) );
AND2x2_ASAP7_75t_L g298 ( .A(n_214), .B(n_144), .Y(n_298) );
AND3x1_ASAP7_75t_L g299 ( .A(n_201), .B(n_145), .C(n_168), .Y(n_299) );
OAI22xp5_ASAP7_75t_L g300 ( .A1(n_217), .A2(n_168), .B1(n_164), .B2(n_129), .Y(n_300) );
BUFx4f_ASAP7_75t_L g301 ( .A(n_193), .Y(n_301) );
NAND2x1p5_ASAP7_75t_L g302 ( .A(n_199), .B(n_140), .Y(n_302) );
INVx2_ASAP7_75t_L g303 ( .A(n_196), .Y(n_303) );
NAND3xp33_ASAP7_75t_L g304 ( .A(n_182), .B(n_132), .C(n_144), .Y(n_304) );
INVx4_ASAP7_75t_L g305 ( .A(n_193), .Y(n_305) );
INVx1_ASAP7_75t_L g306 ( .A(n_196), .Y(n_306) );
INVx5_ASAP7_75t_L g307 ( .A(n_193), .Y(n_307) );
NAND2xp5_ASAP7_75t_L g308 ( .A(n_173), .B(n_164), .Y(n_308) );
INVx2_ASAP7_75t_L g309 ( .A(n_204), .Y(n_309) );
CKINVDCx11_ASAP7_75t_R g310 ( .A(n_220), .Y(n_310) );
INVx1_ASAP7_75t_L g311 ( .A(n_248), .Y(n_311) );
BUFx6f_ASAP7_75t_L g312 ( .A(n_242), .Y(n_312) );
INVx2_ASAP7_75t_L g313 ( .A(n_248), .Y(n_313) );
INVx2_ASAP7_75t_L g314 ( .A(n_265), .Y(n_314) );
BUFx3_ASAP7_75t_L g315 ( .A(n_242), .Y(n_315) );
INVx1_ASAP7_75t_SL g316 ( .A(n_310), .Y(n_316) );
INVx3_ASAP7_75t_L g317 ( .A(n_255), .Y(n_317) );
INVx1_ASAP7_75t_SL g318 ( .A(n_310), .Y(n_318) );
INVx3_ASAP7_75t_L g319 ( .A(n_255), .Y(n_319) );
AOI22xp5_ASAP7_75t_L g320 ( .A1(n_271), .A2(n_218), .B1(n_211), .B2(n_190), .Y(n_320) );
INVx2_ASAP7_75t_SL g321 ( .A(n_268), .Y(n_321) );
INVx2_ASAP7_75t_L g322 ( .A(n_265), .Y(n_322) );
BUFx2_ASAP7_75t_L g323 ( .A(n_271), .Y(n_323) );
OAI22xp5_ASAP7_75t_L g324 ( .A1(n_271), .A2(n_199), .B1(n_207), .B2(n_189), .Y(n_324) );
INVx1_ASAP7_75t_L g325 ( .A(n_309), .Y(n_325) );
AND2x4_ASAP7_75t_L g326 ( .A(n_273), .B(n_195), .Y(n_326) );
BUFx3_ASAP7_75t_L g327 ( .A(n_242), .Y(n_327) );
AOI22xp5_ASAP7_75t_L g328 ( .A1(n_246), .A2(n_218), .B1(n_211), .B2(n_234), .Y(n_328) );
OAI22xp5_ASAP7_75t_L g329 ( .A1(n_268), .A2(n_199), .B1(n_185), .B2(n_177), .Y(n_329) );
BUFx12f_ASAP7_75t_L g330 ( .A(n_264), .Y(n_330) );
INVx1_ASAP7_75t_L g331 ( .A(n_309), .Y(n_331) );
INVx2_ASAP7_75t_L g332 ( .A(n_280), .Y(n_332) );
INVx3_ASAP7_75t_L g333 ( .A(n_255), .Y(n_333) );
AND2x4_ASAP7_75t_L g334 ( .A(n_266), .B(n_211), .Y(n_334) );
OAI22xp5_ASAP7_75t_L g335 ( .A1(n_249), .A2(n_183), .B1(n_229), .B2(n_122), .Y(n_335) );
NOR2xp33_ASAP7_75t_R g336 ( .A(n_289), .B(n_84), .Y(n_336) );
INVx1_ASAP7_75t_L g337 ( .A(n_280), .Y(n_337) );
NOR2xp33_ASAP7_75t_L g338 ( .A(n_277), .B(n_211), .Y(n_338) );
BUFx6f_ASAP7_75t_L g339 ( .A(n_242), .Y(n_339) );
INVxp67_ASAP7_75t_L g340 ( .A(n_269), .Y(n_340) );
INVx3_ASAP7_75t_L g341 ( .A(n_266), .Y(n_341) );
CKINVDCx5p33_ASAP7_75t_R g342 ( .A(n_269), .Y(n_342) );
AND2x4_ASAP7_75t_L g343 ( .A(n_266), .B(n_211), .Y(n_343) );
OAI22xp5_ASAP7_75t_L g344 ( .A1(n_249), .A2(n_216), .B1(n_204), .B2(n_209), .Y(n_344) );
CKINVDCx5p33_ASAP7_75t_R g345 ( .A(n_269), .Y(n_345) );
BUFx2_ASAP7_75t_L g346 ( .A(n_305), .Y(n_346) );
BUFx5_ASAP7_75t_L g347 ( .A(n_253), .Y(n_347) );
BUFx2_ASAP7_75t_L g348 ( .A(n_305), .Y(n_348) );
INVx2_ASAP7_75t_L g349 ( .A(n_290), .Y(n_349) );
NOR2xp33_ASAP7_75t_L g350 ( .A(n_294), .B(n_211), .Y(n_350) );
INVx3_ASAP7_75t_L g351 ( .A(n_305), .Y(n_351) );
OAI221xp5_ASAP7_75t_L g352 ( .A1(n_254), .A2(n_209), .B1(n_216), .B2(n_237), .C(n_220), .Y(n_352) );
NAND2xp5_ASAP7_75t_L g353 ( .A(n_267), .B(n_211), .Y(n_353) );
INVx1_ASAP7_75t_L g354 ( .A(n_261), .Y(n_354) );
AND2x2_ASAP7_75t_L g355 ( .A(n_267), .B(n_235), .Y(n_355) );
NAND2xp5_ASAP7_75t_L g356 ( .A(n_267), .B(n_218), .Y(n_356) );
AOI21xp5_ASAP7_75t_L g357 ( .A1(n_272), .A2(n_231), .B(n_205), .Y(n_357) );
OR2x6_ASAP7_75t_L g358 ( .A(n_261), .B(n_231), .Y(n_358) );
BUFx2_ASAP7_75t_L g359 ( .A(n_274), .Y(n_359) );
NAND2xp5_ASAP7_75t_SL g360 ( .A(n_252), .B(n_231), .Y(n_360) );
INVx1_ASAP7_75t_L g361 ( .A(n_290), .Y(n_361) );
NAND2xp5_ASAP7_75t_L g362 ( .A(n_243), .B(n_218), .Y(n_362) );
INVx2_ASAP7_75t_L g363 ( .A(n_293), .Y(n_363) );
INVx2_ASAP7_75t_L g364 ( .A(n_293), .Y(n_364) );
NAND2xp5_ASAP7_75t_L g365 ( .A(n_247), .B(n_218), .Y(n_365) );
AOI22xp33_ASAP7_75t_L g366 ( .A1(n_359), .A2(n_270), .B1(n_289), .B2(n_260), .Y(n_366) );
INVxp67_ASAP7_75t_SL g367 ( .A(n_323), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_311), .Y(n_368) );
AOI211x1_ASAP7_75t_L g369 ( .A1(n_352), .A2(n_304), .B(n_283), .C(n_291), .Y(n_369) );
INVx1_ASAP7_75t_SL g370 ( .A(n_330), .Y(n_370) );
INVx1_ASAP7_75t_SL g371 ( .A(n_330), .Y(n_371) );
AOI22xp33_ASAP7_75t_L g372 ( .A1(n_359), .A2(n_274), .B1(n_250), .B2(n_285), .Y(n_372) );
NOR2xp33_ASAP7_75t_L g373 ( .A(n_342), .B(n_258), .Y(n_373) );
INVx2_ASAP7_75t_L g374 ( .A(n_313), .Y(n_374) );
AOI22xp33_ASAP7_75t_SL g375 ( .A1(n_336), .A2(n_285), .B1(n_298), .B2(n_296), .Y(n_375) );
AOI22xp33_ASAP7_75t_L g376 ( .A1(n_323), .A2(n_285), .B1(n_263), .B2(n_240), .Y(n_376) );
O2A1O1Ixp33_ASAP7_75t_SL g377 ( .A1(n_311), .A2(n_275), .B(n_306), .C(n_278), .Y(n_377) );
INVx2_ASAP7_75t_SL g378 ( .A(n_334), .Y(n_378) );
OAI22xp5_ASAP7_75t_L g379 ( .A1(n_320), .A2(n_241), .B1(n_251), .B2(n_297), .Y(n_379) );
AND2x2_ASAP7_75t_L g380 ( .A(n_355), .B(n_276), .Y(n_380) );
AOI222xp33_ASAP7_75t_L g381 ( .A1(n_316), .A2(n_244), .B1(n_245), .B2(n_284), .C1(n_287), .C2(n_296), .Y(n_381) );
BUFx12f_ASAP7_75t_L g382 ( .A(n_342), .Y(n_382) );
INVx2_ASAP7_75t_SL g383 ( .A(n_334), .Y(n_383) );
NOR2xp33_ASAP7_75t_L g384 ( .A(n_345), .B(n_287), .Y(n_384) );
INVx1_ASAP7_75t_L g385 ( .A(n_325), .Y(n_385) );
AOI22xp33_ASAP7_75t_L g386 ( .A1(n_345), .A2(n_218), .B1(n_296), .B2(n_287), .Y(n_386) );
BUFx6f_ASAP7_75t_L g387 ( .A(n_312), .Y(n_387) );
INVx6_ASAP7_75t_L g388 ( .A(n_347), .Y(n_388) );
NAND2xp5_ASAP7_75t_L g389 ( .A(n_355), .B(n_308), .Y(n_389) );
AOI22xp5_ASAP7_75t_L g390 ( .A1(n_335), .A2(n_299), .B1(n_257), .B2(n_259), .Y(n_390) );
AOI22xp33_ASAP7_75t_L g391 ( .A1(n_340), .A2(n_262), .B1(n_256), .B2(n_241), .Y(n_391) );
OAI22xp33_ASAP7_75t_L g392 ( .A1(n_318), .A2(n_301), .B1(n_302), .B2(n_307), .Y(n_392) );
INVx2_ASAP7_75t_L g393 ( .A(n_313), .Y(n_393) );
A2O1A1Ixp33_ASAP7_75t_L g394 ( .A1(n_362), .A2(n_281), .B(n_251), .C(n_279), .Y(n_394) );
INVx1_ASAP7_75t_SL g395 ( .A(n_347), .Y(n_395) );
INVx1_ASAP7_75t_L g396 ( .A(n_325), .Y(n_396) );
INVx1_ASAP7_75t_L g397 ( .A(n_331), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_331), .Y(n_398) );
AND2x2_ASAP7_75t_L g399 ( .A(n_337), .B(n_303), .Y(n_399) );
AOI22x1_ASAP7_75t_L g400 ( .A1(n_395), .A2(n_337), .B1(n_361), .B2(n_357), .Y(n_400) );
AOI22xp33_ASAP7_75t_L g401 ( .A1(n_375), .A2(n_338), .B1(n_350), .B2(n_326), .Y(n_401) );
OAI22xp33_ASAP7_75t_L g402 ( .A1(n_390), .A2(n_324), .B1(n_321), .B2(n_353), .Y(n_402) );
HB1xp67_ASAP7_75t_L g403 ( .A(n_370), .Y(n_403) );
OAI21xp5_ASAP7_75t_L g404 ( .A1(n_394), .A2(n_365), .B(n_361), .Y(n_404) );
OAI221xp5_ASAP7_75t_L g405 ( .A1(n_366), .A2(n_356), .B1(n_344), .B2(n_329), .C(n_354), .Y(n_405) );
AOI221xp5_ASAP7_75t_L g406 ( .A1(n_373), .A2(n_326), .B1(n_300), .B2(n_321), .C(n_292), .Y(n_406) );
OAI21xp5_ASAP7_75t_L g407 ( .A1(n_379), .A2(n_364), .B(n_363), .Y(n_407) );
OAI221xp5_ASAP7_75t_SL g408 ( .A1(n_376), .A2(n_328), .B1(n_155), .B2(n_149), .C(n_363), .Y(n_408) );
HB1xp67_ASAP7_75t_L g409 ( .A(n_371), .Y(n_409) );
OAI211xp5_ASAP7_75t_SL g410 ( .A1(n_381), .A2(n_155), .B(n_92), .C(n_224), .Y(n_410) );
OAI211xp5_ASAP7_75t_L g411 ( .A1(n_390), .A2(n_155), .B(n_237), .C(n_233), .Y(n_411) );
OAI22xp5_ASAP7_75t_SL g412 ( .A1(n_384), .A2(n_326), .B1(n_314), .B2(n_322), .Y(n_412) );
AOI22xp33_ASAP7_75t_L g413 ( .A1(n_380), .A2(n_347), .B1(n_322), .B2(n_314), .Y(n_413) );
OAI22xp33_ASAP7_75t_L g414 ( .A1(n_389), .A2(n_301), .B1(n_346), .B2(n_348), .Y(n_414) );
AOI22xp33_ASAP7_75t_L g415 ( .A1(n_380), .A2(n_347), .B1(n_349), .B2(n_332), .Y(n_415) );
OAI21x1_ASAP7_75t_L g416 ( .A1(n_374), .A2(n_364), .B(n_332), .Y(n_416) );
OR2x2_ASAP7_75t_L g417 ( .A(n_368), .B(n_385), .Y(n_417) );
NOR2xp33_ASAP7_75t_SL g418 ( .A(n_395), .B(n_334), .Y(n_418) );
AOI22xp33_ASAP7_75t_SL g419 ( .A1(n_367), .A2(n_347), .B1(n_343), .B2(n_346), .Y(n_419) );
AOI22xp33_ASAP7_75t_L g420 ( .A1(n_372), .A2(n_382), .B1(n_398), .B2(n_397), .Y(n_420) );
AOI21x1_ASAP7_75t_L g421 ( .A1(n_368), .A2(n_186), .B(n_200), .Y(n_421) );
OAI22xp5_ASAP7_75t_L g422 ( .A1(n_385), .A2(n_398), .B1(n_397), .B2(n_396), .Y(n_422) );
INVx1_ASAP7_75t_L g423 ( .A(n_396), .Y(n_423) );
AND2x2_ASAP7_75t_L g424 ( .A(n_399), .B(n_349), .Y(n_424) );
AOI221xp5_ASAP7_75t_L g425 ( .A1(n_369), .A2(n_124), .B1(n_288), .B2(n_233), .C(n_235), .Y(n_425) );
OAI211xp5_ASAP7_75t_L g426 ( .A1(n_369), .A2(n_224), .B(n_124), .C(n_152), .Y(n_426) );
AND2x6_ASAP7_75t_SL g427 ( .A(n_382), .B(n_343), .Y(n_427) );
INVx2_ASAP7_75t_L g428 ( .A(n_374), .Y(n_428) );
NAND2xp5_ASAP7_75t_L g429 ( .A(n_423), .B(n_399), .Y(n_429) );
HB1xp67_ASAP7_75t_L g430 ( .A(n_424), .Y(n_430) );
OAI221xp5_ASAP7_75t_SL g431 ( .A1(n_420), .A2(n_386), .B1(n_391), .B2(n_392), .C(n_383), .Y(n_431) );
OAI22xp5_ASAP7_75t_L g432 ( .A1(n_401), .A2(n_388), .B1(n_393), .B2(n_348), .Y(n_432) );
INVx2_ASAP7_75t_L g433 ( .A(n_428), .Y(n_433) );
INVx1_ASAP7_75t_L g434 ( .A(n_423), .Y(n_434) );
AO21x2_ASAP7_75t_L g435 ( .A1(n_426), .A2(n_377), .B(n_393), .Y(n_435) );
AOI22xp33_ASAP7_75t_L g436 ( .A1(n_412), .A2(n_383), .B1(n_378), .B2(n_347), .Y(n_436) );
CKINVDCx20_ASAP7_75t_R g437 ( .A(n_403), .Y(n_437) );
OAI211xp5_ASAP7_75t_SL g438 ( .A1(n_409), .A2(n_224), .B(n_166), .C(n_378), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_422), .Y(n_439) );
NAND2xp5_ASAP7_75t_L g440 ( .A(n_424), .B(n_303), .Y(n_440) );
NOR2xp67_ASAP7_75t_L g441 ( .A(n_422), .B(n_387), .Y(n_441) );
INVx2_ASAP7_75t_L g442 ( .A(n_428), .Y(n_442) );
INVx2_ASAP7_75t_L g443 ( .A(n_428), .Y(n_443) );
AOI221xp5_ASAP7_75t_L g444 ( .A1(n_410), .A2(n_124), .B1(n_166), .B2(n_302), .C(n_158), .Y(n_444) );
AOI221xp5_ASAP7_75t_L g445 ( .A1(n_402), .A2(n_166), .B1(n_158), .B2(n_162), .C(n_170), .Y(n_445) );
OAI211xp5_ASAP7_75t_SL g446 ( .A1(n_406), .A2(n_166), .B(n_186), .C(n_200), .Y(n_446) );
OAI33xp33_ASAP7_75t_L g447 ( .A1(n_412), .A2(n_226), .A3(n_203), .B1(n_230), .B2(n_236), .B3(n_13), .Y(n_447) );
OAI221xp5_ASAP7_75t_SL g448 ( .A1(n_425), .A2(n_358), .B1(n_226), .B2(n_203), .C(n_351), .Y(n_448) );
NAND3xp33_ASAP7_75t_L g449 ( .A(n_425), .B(n_162), .C(n_170), .Y(n_449) );
OAI21xp5_ASAP7_75t_L g450 ( .A1(n_404), .A2(n_360), .B(n_156), .Y(n_450) );
INVx1_ASAP7_75t_L g451 ( .A(n_417), .Y(n_451) );
INVx2_ASAP7_75t_L g452 ( .A(n_416), .Y(n_452) );
NAND2xp5_ASAP7_75t_SL g453 ( .A(n_414), .B(n_387), .Y(n_453) );
NAND3xp33_ASAP7_75t_L g454 ( .A(n_400), .B(n_159), .C(n_162), .Y(n_454) );
NAND2xp5_ASAP7_75t_L g455 ( .A(n_417), .B(n_347), .Y(n_455) );
INVx3_ASAP7_75t_L g456 ( .A(n_416), .Y(n_456) );
OAI22xp33_ASAP7_75t_L g457 ( .A1(n_418), .A2(n_388), .B1(n_317), .B2(n_351), .Y(n_457) );
OA21x2_ASAP7_75t_L g458 ( .A1(n_400), .A2(n_230), .B(n_236), .Y(n_458) );
INVx1_ASAP7_75t_SL g459 ( .A(n_418), .Y(n_459) );
OA21x2_ASAP7_75t_L g460 ( .A1(n_407), .A2(n_282), .B(n_152), .Y(n_460) );
INVx4_ASAP7_75t_L g461 ( .A(n_427), .Y(n_461) );
OAI211xp5_ASAP7_75t_SL g462 ( .A1(n_405), .A2(n_351), .B(n_317), .C(n_319), .Y(n_462) );
OAI21x1_ASAP7_75t_L g463 ( .A1(n_421), .A2(n_152), .B(n_341), .Y(n_463) );
NOR3xp33_ASAP7_75t_L g464 ( .A(n_405), .B(n_333), .C(n_319), .Y(n_464) );
AND2x2_ASAP7_75t_L g465 ( .A(n_407), .B(n_388), .Y(n_465) );
AND2x2_ASAP7_75t_L g466 ( .A(n_434), .B(n_404), .Y(n_466) );
AND2x2_ASAP7_75t_L g467 ( .A(n_434), .B(n_152), .Y(n_467) );
AOI22xp5_ASAP7_75t_L g468 ( .A1(n_461), .A2(n_415), .B1(n_413), .B2(n_419), .Y(n_468) );
AOI22xp33_ASAP7_75t_L g469 ( .A1(n_461), .A2(n_388), .B1(n_347), .B2(n_327), .Y(n_469) );
BUFx2_ASAP7_75t_L g470 ( .A(n_461), .Y(n_470) );
INVx2_ASAP7_75t_L g471 ( .A(n_433), .Y(n_471) );
AOI22xp33_ASAP7_75t_L g472 ( .A1(n_461), .A2(n_315), .B1(n_327), .B2(n_387), .Y(n_472) );
INVx2_ASAP7_75t_L g473 ( .A(n_433), .Y(n_473) );
AOI21xp5_ASAP7_75t_L g474 ( .A1(n_454), .A2(n_387), .B(n_408), .Y(n_474) );
AND2x4_ASAP7_75t_L g475 ( .A(n_441), .B(n_387), .Y(n_475) );
NOR3xp33_ASAP7_75t_L g476 ( .A(n_438), .B(n_411), .C(n_421), .Y(n_476) );
INVx1_ASAP7_75t_L g477 ( .A(n_451), .Y(n_477) );
AND2x4_ASAP7_75t_L g478 ( .A(n_441), .B(n_315), .Y(n_478) );
NAND2xp5_ASAP7_75t_SL g479 ( .A(n_459), .B(n_339), .Y(n_479) );
NAND3xp33_ASAP7_75t_L g480 ( .A(n_444), .B(n_159), .C(n_162), .Y(n_480) );
HB1xp67_ASAP7_75t_L g481 ( .A(n_430), .Y(n_481) );
AND2x2_ASAP7_75t_L g482 ( .A(n_433), .B(n_8), .Y(n_482) );
AND2x2_ASAP7_75t_L g483 ( .A(n_451), .B(n_8), .Y(n_483) );
INVx1_ASAP7_75t_L g484 ( .A(n_429), .Y(n_484) );
AOI22xp33_ASAP7_75t_L g485 ( .A1(n_447), .A2(n_339), .B1(n_312), .B2(n_156), .Y(n_485) );
HB1xp67_ASAP7_75t_L g486 ( .A(n_442), .Y(n_486) );
INVx2_ASAP7_75t_L g487 ( .A(n_442), .Y(n_487) );
INVx1_ASAP7_75t_L g488 ( .A(n_455), .Y(n_488) );
AOI33xp33_ASAP7_75t_L g489 ( .A1(n_439), .A2(n_9), .A3(n_10), .B1(n_12), .B2(n_13), .B3(n_14), .Y(n_489) );
NAND4xp25_ASAP7_75t_L g490 ( .A(n_431), .B(n_436), .C(n_439), .D(n_445), .Y(n_490) );
NAND4xp25_ASAP7_75t_L g491 ( .A(n_464), .B(n_9), .C(n_10), .D(n_16), .Y(n_491) );
AOI22xp5_ASAP7_75t_L g492 ( .A1(n_437), .A2(n_343), .B1(n_156), .B2(n_341), .Y(n_492) );
INVx1_ASAP7_75t_L g493 ( .A(n_440), .Y(n_493) );
INVx1_ASAP7_75t_L g494 ( .A(n_442), .Y(n_494) );
NAND2x1p5_ASAP7_75t_SL g495 ( .A(n_453), .B(n_427), .Y(n_495) );
INVx1_ASAP7_75t_L g496 ( .A(n_443), .Y(n_496) );
INVx1_ASAP7_75t_L g497 ( .A(n_443), .Y(n_497) );
INVx1_ASAP7_75t_L g498 ( .A(n_443), .Y(n_498) );
OAI31xp33_ASAP7_75t_L g499 ( .A1(n_448), .A2(n_317), .A3(n_319), .B(n_333), .Y(n_499) );
AND2x4_ASAP7_75t_L g500 ( .A(n_465), .B(n_67), .Y(n_500) );
INVx2_ASAP7_75t_SL g501 ( .A(n_465), .Y(n_501) );
AND2x2_ASAP7_75t_L g502 ( .A(n_459), .B(n_16), .Y(n_502) );
AOI22xp5_ASAP7_75t_L g503 ( .A1(n_432), .A2(n_156), .B1(n_341), .B2(n_333), .Y(n_503) );
OAI33xp33_ASAP7_75t_L g504 ( .A1(n_446), .A2(n_17), .A3(n_19), .B1(n_170), .B2(n_162), .B3(n_159), .Y(n_504) );
OR2x2_ASAP7_75t_L g505 ( .A(n_452), .B(n_19), .Y(n_505) );
INVx1_ASAP7_75t_L g506 ( .A(n_452), .Y(n_506) );
NAND2xp5_ASAP7_75t_L g507 ( .A(n_449), .B(n_159), .Y(n_507) );
INVx4_ASAP7_75t_L g508 ( .A(n_456), .Y(n_508) );
AND2x2_ASAP7_75t_L g509 ( .A(n_452), .B(n_170), .Y(n_509) );
OR2x2_ASAP7_75t_L g510 ( .A(n_456), .B(n_159), .Y(n_510) );
BUFx2_ASAP7_75t_L g511 ( .A(n_456), .Y(n_511) );
INVx1_ASAP7_75t_L g512 ( .A(n_456), .Y(n_512) );
OAI22xp5_ASAP7_75t_L g513 ( .A1(n_449), .A2(n_339), .B1(n_312), .B2(n_358), .Y(n_513) );
INVx1_ASAP7_75t_L g514 ( .A(n_435), .Y(n_514) );
OAI221xp5_ASAP7_75t_SL g515 ( .A1(n_457), .A2(n_358), .B1(n_219), .B2(n_197), .C(n_174), .Y(n_515) );
INVx1_ASAP7_75t_SL g516 ( .A(n_435), .Y(n_516) );
NAND3xp33_ASAP7_75t_L g517 ( .A(n_454), .B(n_170), .C(n_159), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_435), .B(n_159), .Y(n_518) );
AND2x2_ASAP7_75t_L g519 ( .A(n_501), .B(n_458), .Y(n_519) );
INVxp33_ASAP7_75t_L g520 ( .A(n_481), .Y(n_520) );
NAND3xp33_ASAP7_75t_SL g521 ( .A(n_489), .B(n_450), .C(n_156), .Y(n_521) );
INVx1_ASAP7_75t_L g522 ( .A(n_477), .Y(n_522) );
AND2x2_ASAP7_75t_L g523 ( .A(n_501), .B(n_458), .Y(n_523) );
OAI21xp33_ASAP7_75t_L g524 ( .A1(n_489), .A2(n_162), .B(n_170), .Y(n_524) );
INVx1_ASAP7_75t_L g525 ( .A(n_482), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g526 ( .A(n_484), .B(n_460), .Y(n_526) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_493), .B(n_460), .Y(n_527) );
INVx2_ASAP7_75t_L g528 ( .A(n_471), .Y(n_528) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_488), .B(n_460), .Y(n_529) );
HB1xp67_ASAP7_75t_L g530 ( .A(n_486), .Y(n_530) );
AND2x2_ASAP7_75t_L g531 ( .A(n_466), .B(n_458), .Y(n_531) );
AND2x2_ASAP7_75t_L g532 ( .A(n_466), .B(n_458), .Y(n_532) );
INVx2_ASAP7_75t_SL g533 ( .A(n_470), .Y(n_533) );
OR2x2_ASAP7_75t_L g534 ( .A(n_494), .B(n_170), .Y(n_534) );
OR2x2_ASAP7_75t_L g535 ( .A(n_496), .B(n_162), .Y(n_535) );
NOR3xp33_ASAP7_75t_L g536 ( .A(n_491), .B(n_462), .C(n_450), .Y(n_536) );
OR2x2_ASAP7_75t_L g537 ( .A(n_497), .B(n_460), .Y(n_537) );
NOR2x1_ASAP7_75t_L g538 ( .A(n_505), .B(n_339), .Y(n_538) );
AND2x2_ASAP7_75t_L g539 ( .A(n_471), .B(n_463), .Y(n_539) );
INVx2_ASAP7_75t_L g540 ( .A(n_473), .Y(n_540) );
INVx3_ASAP7_75t_L g541 ( .A(n_508), .Y(n_541) );
INVx1_ASAP7_75t_L g542 ( .A(n_482), .Y(n_542) );
INVx1_ASAP7_75t_L g543 ( .A(n_498), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g544 ( .A(n_483), .B(n_156), .Y(n_544) );
INVx1_ASAP7_75t_L g545 ( .A(n_487), .Y(n_545) );
NOR3xp33_ASAP7_75t_L g546 ( .A(n_504), .B(n_219), .C(n_197), .Y(n_546) );
INVxp67_ASAP7_75t_SL g547 ( .A(n_487), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_502), .B(n_156), .Y(n_548) );
INVx2_ASAP7_75t_L g549 ( .A(n_506), .Y(n_549) );
NOR2x1_ASAP7_75t_L g550 ( .A(n_500), .B(n_508), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g551 ( .A(n_500), .B(n_339), .Y(n_551) );
INVx1_ASAP7_75t_L g552 ( .A(n_509), .Y(n_552) );
AND2x2_ASAP7_75t_L g553 ( .A(n_512), .B(n_23), .Y(n_553) );
INVx1_ASAP7_75t_SL g554 ( .A(n_500), .Y(n_554) );
NAND2xp5_ASAP7_75t_L g555 ( .A(n_490), .B(n_312), .Y(n_555) );
NAND4xp25_ASAP7_75t_L g556 ( .A(n_468), .B(n_174), .C(n_282), .D(n_28), .Y(n_556) );
AND2x2_ASAP7_75t_L g557 ( .A(n_511), .B(n_25), .Y(n_557) );
INVx1_ASAP7_75t_L g558 ( .A(n_495), .Y(n_558) );
INVxp67_ASAP7_75t_SL g559 ( .A(n_510), .Y(n_559) );
INVxp67_ASAP7_75t_SL g560 ( .A(n_479), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_467), .B(n_312), .Y(n_561) );
INVx1_ASAP7_75t_L g562 ( .A(n_495), .Y(n_562) );
INVx1_ASAP7_75t_L g563 ( .A(n_467), .Y(n_563) );
INVx3_ASAP7_75t_L g564 ( .A(n_508), .Y(n_564) );
INVxp67_ASAP7_75t_L g565 ( .A(n_513), .Y(n_565) );
OR2x2_ASAP7_75t_L g566 ( .A(n_479), .B(n_27), .Y(n_566) );
NAND3xp33_ASAP7_75t_L g567 ( .A(n_476), .B(n_184), .C(n_191), .Y(n_567) );
NOR2xp33_ASAP7_75t_L g568 ( .A(n_515), .B(n_30), .Y(n_568) );
NOR2xp33_ASAP7_75t_SL g569 ( .A(n_499), .B(n_307), .Y(n_569) );
INVx1_ASAP7_75t_L g570 ( .A(n_478), .Y(n_570) );
OR2x2_ASAP7_75t_L g571 ( .A(n_478), .B(n_31), .Y(n_571) );
OR2x2_ASAP7_75t_L g572 ( .A(n_478), .B(n_33), .Y(n_572) );
INVx1_ASAP7_75t_L g573 ( .A(n_518), .Y(n_573) );
OR2x2_ASAP7_75t_L g574 ( .A(n_475), .B(n_37), .Y(n_574) );
OAI21xp5_ASAP7_75t_SL g575 ( .A1(n_492), .A2(n_252), .B(n_286), .Y(n_575) );
INVx1_ASAP7_75t_L g576 ( .A(n_514), .Y(n_576) );
INVx2_ASAP7_75t_L g577 ( .A(n_475), .Y(n_577) );
OR2x2_ASAP7_75t_L g578 ( .A(n_530), .B(n_516), .Y(n_578) );
INVx1_ASAP7_75t_L g579 ( .A(n_522), .Y(n_579) );
NAND3xp33_ASAP7_75t_L g580 ( .A(n_558), .B(n_485), .C(n_480), .Y(n_580) );
AND2x2_ASAP7_75t_L g581 ( .A(n_563), .B(n_475), .Y(n_581) );
OAI21xp33_ASAP7_75t_L g582 ( .A1(n_520), .A2(n_485), .B(n_503), .Y(n_582) );
INVx1_ASAP7_75t_L g583 ( .A(n_530), .Y(n_583) );
AND2x2_ASAP7_75t_L g584 ( .A(n_531), .B(n_507), .Y(n_584) );
HB1xp67_ASAP7_75t_L g585 ( .A(n_520), .Y(n_585) );
NAND2xp5_ASAP7_75t_L g586 ( .A(n_525), .B(n_472), .Y(n_586) );
NOR2xp33_ASAP7_75t_SL g587 ( .A(n_550), .B(n_474), .Y(n_587) );
INVx1_ASAP7_75t_L g588 ( .A(n_543), .Y(n_588) );
NAND3xp33_ASAP7_75t_L g589 ( .A(n_562), .B(n_472), .C(n_469), .Y(n_589) );
INVx1_ASAP7_75t_L g590 ( .A(n_549), .Y(n_590) );
AND2x2_ASAP7_75t_L g591 ( .A(n_531), .B(n_469), .Y(n_591) );
INVx1_ASAP7_75t_L g592 ( .A(n_549), .Y(n_592) );
INVx1_ASAP7_75t_L g593 ( .A(n_545), .Y(n_593) );
INVx1_ASAP7_75t_L g594 ( .A(n_547), .Y(n_594) );
NOR2xp33_ASAP7_75t_L g595 ( .A(n_555), .B(n_517), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g596 ( .A(n_542), .B(n_43), .Y(n_596) );
INVxp67_ASAP7_75t_SL g597 ( .A(n_559), .Y(n_597) );
NAND3xp33_ASAP7_75t_L g598 ( .A(n_565), .B(n_194), .C(n_191), .Y(n_598) );
AND2x2_ASAP7_75t_L g599 ( .A(n_532), .B(n_577), .Y(n_599) );
AND2x2_ASAP7_75t_L g600 ( .A(n_532), .B(n_44), .Y(n_600) );
AO221x1_ASAP7_75t_L g601 ( .A1(n_541), .A2(n_252), .B1(n_286), .B2(n_52), .C(n_53), .Y(n_601) );
OR2x2_ASAP7_75t_L g602 ( .A(n_526), .B(n_45), .Y(n_602) );
INVx1_ASAP7_75t_L g603 ( .A(n_533), .Y(n_603) );
NAND2xp5_ASAP7_75t_L g604 ( .A(n_552), .B(n_47), .Y(n_604) );
NOR2xp33_ASAP7_75t_L g605 ( .A(n_556), .B(n_55), .Y(n_605) );
AND2x2_ASAP7_75t_L g606 ( .A(n_577), .B(n_61), .Y(n_606) );
INVx1_ASAP7_75t_L g607 ( .A(n_533), .Y(n_607) );
INVx1_ASAP7_75t_L g608 ( .A(n_576), .Y(n_608) );
AND2x2_ASAP7_75t_L g609 ( .A(n_519), .B(n_62), .Y(n_609) );
AND2x2_ASAP7_75t_L g610 ( .A(n_519), .B(n_63), .Y(n_610) );
AND2x2_ASAP7_75t_L g611 ( .A(n_523), .B(n_64), .Y(n_611) );
INVx1_ASAP7_75t_L g612 ( .A(n_528), .Y(n_612) );
INVx1_ASAP7_75t_SL g613 ( .A(n_554), .Y(n_613) );
INVx1_ASAP7_75t_L g614 ( .A(n_540), .Y(n_614) );
BUFx2_ASAP7_75t_L g615 ( .A(n_541), .Y(n_615) );
OR2x2_ASAP7_75t_L g616 ( .A(n_527), .B(n_66), .Y(n_616) );
AOI221x1_ASAP7_75t_L g617 ( .A1(n_524), .A2(n_194), .B1(n_191), .B2(n_184), .C(n_76), .Y(n_617) );
INVx1_ASAP7_75t_L g618 ( .A(n_534), .Y(n_618) );
NAND3xp33_ASAP7_75t_SL g619 ( .A(n_536), .B(n_69), .C(n_71), .Y(n_619) );
AOI21xp5_ASAP7_75t_L g620 ( .A1(n_575), .A2(n_358), .B(n_307), .Y(n_620) );
INVx1_ASAP7_75t_L g621 ( .A(n_535), .Y(n_621) );
AND2x2_ASAP7_75t_L g622 ( .A(n_523), .B(n_184), .Y(n_622) );
NAND2xp5_ASAP7_75t_L g623 ( .A(n_570), .B(n_184), .Y(n_623) );
NAND4xp75_ASAP7_75t_L g624 ( .A(n_557), .B(n_307), .C(n_252), .D(n_194), .Y(n_624) );
INVxp67_ASAP7_75t_L g625 ( .A(n_557), .Y(n_625) );
NOR3xp33_ASAP7_75t_L g626 ( .A(n_521), .B(n_184), .C(n_191), .Y(n_626) );
AND2x2_ASAP7_75t_L g627 ( .A(n_573), .B(n_191), .Y(n_627) );
XNOR2xp5_ASAP7_75t_L g628 ( .A(n_571), .B(n_286), .Y(n_628) );
INVx1_ASAP7_75t_L g629 ( .A(n_583), .Y(n_629) );
INVx1_ASAP7_75t_SL g630 ( .A(n_613), .Y(n_630) );
NOR2xp33_ASAP7_75t_L g631 ( .A(n_585), .B(n_572), .Y(n_631) );
NAND2xp5_ASAP7_75t_L g632 ( .A(n_597), .B(n_529), .Y(n_632) );
INVx1_ASAP7_75t_L g633 ( .A(n_579), .Y(n_633) );
INVx1_ASAP7_75t_L g634 ( .A(n_588), .Y(n_634) );
NAND2xp5_ASAP7_75t_L g635 ( .A(n_608), .B(n_539), .Y(n_635) );
OAI21xp5_ASAP7_75t_L g636 ( .A1(n_589), .A2(n_605), .B(n_619), .Y(n_636) );
NAND2xp5_ASAP7_75t_SL g637 ( .A(n_587), .B(n_564), .Y(n_637) );
INVx3_ASAP7_75t_L g638 ( .A(n_615), .Y(n_638) );
INVx1_ASAP7_75t_L g639 ( .A(n_593), .Y(n_639) );
OAI22xp5_ASAP7_75t_L g640 ( .A1(n_625), .A2(n_564), .B1(n_541), .B2(n_574), .Y(n_640) );
NAND2xp5_ASAP7_75t_SL g641 ( .A(n_615), .B(n_564), .Y(n_641) );
NAND2xp5_ASAP7_75t_L g642 ( .A(n_591), .B(n_537), .Y(n_642) );
INVx1_ASAP7_75t_SL g643 ( .A(n_603), .Y(n_643) );
OAI22xp33_ASAP7_75t_L g644 ( .A1(n_602), .A2(n_569), .B1(n_566), .B2(n_567), .Y(n_644) );
INVx1_ASAP7_75t_L g645 ( .A(n_590), .Y(n_645) );
INVx1_ASAP7_75t_L g646 ( .A(n_592), .Y(n_646) );
INVx1_ASAP7_75t_SL g647 ( .A(n_607), .Y(n_647) );
AND4x1_ASAP7_75t_L g648 ( .A(n_605), .B(n_568), .C(n_538), .D(n_546), .Y(n_648) );
INVxp67_ASAP7_75t_L g649 ( .A(n_594), .Y(n_649) );
AND2x2_ASAP7_75t_L g650 ( .A(n_591), .B(n_560), .Y(n_650) );
INVx1_ASAP7_75t_L g651 ( .A(n_612), .Y(n_651) );
OR2x2_ASAP7_75t_L g652 ( .A(n_578), .B(n_561), .Y(n_652) );
NAND2xp5_ASAP7_75t_L g653 ( .A(n_618), .B(n_553), .Y(n_653) );
XNOR2xp5_ASAP7_75t_L g654 ( .A(n_628), .B(n_581), .Y(n_654) );
AOI21xp5_ASAP7_75t_L g655 ( .A1(n_601), .A2(n_551), .B(n_566), .Y(n_655) );
INVx1_ASAP7_75t_L g656 ( .A(n_614), .Y(n_656) );
AOI22xp5_ASAP7_75t_L g657 ( .A1(n_582), .A2(n_568), .B1(n_548), .B2(n_544), .Y(n_657) );
NAND3xp33_ASAP7_75t_SL g658 ( .A(n_626), .B(n_286), .C(n_194), .Y(n_658) );
INVx1_ASAP7_75t_L g659 ( .A(n_581), .Y(n_659) );
INVx1_ASAP7_75t_SL g660 ( .A(n_600), .Y(n_660) );
AO22x2_ASAP7_75t_L g661 ( .A1(n_621), .A2(n_194), .B1(n_295), .B2(n_578), .Y(n_661) );
INVx1_ASAP7_75t_L g662 ( .A(n_586), .Y(n_662) );
OAI222xp33_ASAP7_75t_L g663 ( .A1(n_600), .A2(n_295), .B1(n_610), .B2(n_611), .C1(n_609), .C2(n_628), .Y(n_663) );
NAND3xp33_ASAP7_75t_L g664 ( .A(n_595), .B(n_295), .C(n_580), .Y(n_664) );
AOI221xp5_ASAP7_75t_L g665 ( .A1(n_595), .A2(n_295), .B1(n_584), .B2(n_596), .C(n_611), .Y(n_665) );
NOR2xp33_ASAP7_75t_L g666 ( .A(n_604), .B(n_616), .Y(n_666) );
NAND2xp5_ASAP7_75t_L g667 ( .A(n_609), .B(n_610), .Y(n_667) );
OAI211xp5_ASAP7_75t_SL g668 ( .A1(n_602), .A2(n_616), .B(n_623), .C(n_620), .Y(n_668) );
OAI321xp33_ASAP7_75t_L g669 ( .A1(n_598), .A2(n_606), .A3(n_622), .B1(n_627), .B2(n_617), .C(n_624), .Y(n_669) );
NAND2xp5_ASAP7_75t_L g670 ( .A(n_606), .B(n_624), .Y(n_670) );
OAI211xp5_ASAP7_75t_L g671 ( .A1(n_597), .A2(n_562), .B(n_558), .C(n_310), .Y(n_671) );
INVx1_ASAP7_75t_L g672 ( .A(n_579), .Y(n_672) );
NOR2xp33_ASAP7_75t_L g673 ( .A(n_585), .B(n_520), .Y(n_673) );
OAI21xp5_ASAP7_75t_L g674 ( .A1(n_589), .A2(n_524), .B(n_558), .Y(n_674) );
INVxp67_ASAP7_75t_L g675 ( .A(n_585), .Y(n_675) );
AND2x2_ASAP7_75t_L g676 ( .A(n_585), .B(n_599), .Y(n_676) );
INVxp67_ASAP7_75t_L g677 ( .A(n_585), .Y(n_677) );
INVx1_ASAP7_75t_L g678 ( .A(n_579), .Y(n_678) );
NAND2xp5_ASAP7_75t_L g679 ( .A(n_597), .B(n_585), .Y(n_679) );
NAND2xp5_ASAP7_75t_L g680 ( .A(n_597), .B(n_585), .Y(n_680) );
OAI22xp33_ASAP7_75t_L g681 ( .A1(n_638), .A2(n_660), .B1(n_637), .B2(n_641), .Y(n_681) );
INVx2_ASAP7_75t_L g682 ( .A(n_638), .Y(n_682) );
INVx1_ASAP7_75t_L g683 ( .A(n_679), .Y(n_683) );
A2O1A1Ixp33_ASAP7_75t_L g684 ( .A1(n_636), .A2(n_671), .B(n_673), .C(n_637), .Y(n_684) );
INVx1_ASAP7_75t_L g685 ( .A(n_680), .Y(n_685) );
NAND2xp5_ASAP7_75t_L g686 ( .A(n_662), .B(n_677), .Y(n_686) );
OAI22xp5_ASAP7_75t_L g687 ( .A1(n_654), .A2(n_630), .B1(n_638), .B2(n_641), .Y(n_687) );
OAI21xp33_ASAP7_75t_L g688 ( .A1(n_650), .A2(n_675), .B(n_674), .Y(n_688) );
OAI21xp5_ASAP7_75t_L g689 ( .A1(n_664), .A2(n_655), .B(n_663), .Y(n_689) );
HB1xp67_ASAP7_75t_L g690 ( .A(n_649), .Y(n_690) );
XNOR2xp5_ASAP7_75t_L g691 ( .A(n_654), .B(n_657), .Y(n_691) );
AO22x1_ASAP7_75t_SL g692 ( .A1(n_663), .A2(n_678), .B1(n_672), .B2(n_634), .Y(n_692) );
INVxp67_ASAP7_75t_L g693 ( .A(n_661), .Y(n_693) );
AO22x1_ASAP7_75t_L g694 ( .A1(n_643), .A2(n_647), .B1(n_640), .B2(n_670), .Y(n_694) );
NAND2xp5_ASAP7_75t_L g695 ( .A(n_693), .B(n_650), .Y(n_695) );
OAI21xp33_ASAP7_75t_L g696 ( .A1(n_688), .A2(n_632), .B(n_631), .Y(n_696) );
INVx1_ASAP7_75t_L g697 ( .A(n_690), .Y(n_697) );
OAI211xp5_ASAP7_75t_SL g698 ( .A1(n_684), .A2(n_665), .B(n_629), .C(n_633), .Y(n_698) );
AOI21xp5_ASAP7_75t_L g699 ( .A1(n_687), .A2(n_661), .B(n_669), .Y(n_699) );
INVx1_ASAP7_75t_L g700 ( .A(n_690), .Y(n_700) );
OAI21xp5_ASAP7_75t_L g701 ( .A1(n_689), .A2(n_668), .B(n_644), .Y(n_701) );
O2A1O1Ixp33_ASAP7_75t_L g702 ( .A1(n_693), .A2(n_668), .B(n_658), .C(n_629), .Y(n_702) );
NAND4xp25_ASAP7_75t_L g703 ( .A(n_701), .B(n_666), .C(n_686), .D(n_683), .Y(n_703) );
NOR3xp33_ASAP7_75t_L g704 ( .A(n_702), .B(n_694), .C(n_681), .Y(n_704) );
OR3x1_ASAP7_75t_L g705 ( .A(n_698), .B(n_692), .C(n_685), .Y(n_705) );
NAND4xp25_ASAP7_75t_L g706 ( .A(n_699), .B(n_691), .C(n_667), .D(n_682), .Y(n_706) );
INVx1_ASAP7_75t_L g707 ( .A(n_697), .Y(n_707) );
NAND5xp2_ASAP7_75t_L g708 ( .A(n_704), .B(n_700), .C(n_696), .D(n_695), .E(n_648), .Y(n_708) );
XNOR2xp5_ASAP7_75t_L g709 ( .A(n_706), .B(n_661), .Y(n_709) );
AND2x4_ASAP7_75t_L g710 ( .A(n_707), .B(n_676), .Y(n_710) );
OAI22xp5_ASAP7_75t_L g711 ( .A1(n_709), .A2(n_705), .B1(n_703), .B2(n_642), .Y(n_711) );
AOI21xp5_ASAP7_75t_L g712 ( .A1(n_708), .A2(n_639), .B(n_635), .Y(n_712) );
OAI22xp5_ASAP7_75t_SL g713 ( .A1(n_711), .A2(n_710), .B1(n_653), .B2(n_659), .Y(n_713) );
INVx1_ASAP7_75t_L g714 ( .A(n_713), .Y(n_714) );
OAI22xp33_ASAP7_75t_L g715 ( .A1(n_714), .A2(n_712), .B1(n_710), .B2(n_652), .Y(n_715) );
AOI221xp5_ASAP7_75t_L g716 ( .A1(n_715), .A2(n_645), .B1(n_646), .B2(n_656), .C(n_651), .Y(n_716) );
endmodule