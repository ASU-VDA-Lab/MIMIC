module fake_jpeg_6656_n_344 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_344);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_344;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVxp67_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_7),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

BUFx12_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_25),
.Y(n_36)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_36),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_25),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_37),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_38),
.Y(n_62)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_35),
.Y(n_39)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_39),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_40),
.Y(n_71)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_19),
.Y(n_41)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_18),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_42),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_21),
.Y(n_43)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_43),
.Y(n_63)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_19),
.Y(n_44)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_44),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_26),
.B(n_15),
.Y(n_45)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_45),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_30),
.Y(n_46)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_46),
.Y(n_54)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_20),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_47),
.A2(n_27),
.B1(n_31),
.B2(n_33),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_21),
.Y(n_48)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_48),
.Y(n_58)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_46),
.Y(n_49)
);

INVx11_ASAP7_75t_L g77 ( 
.A(n_49),
.Y(n_77)
);

OAI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_41),
.A2(n_33),
.B1(n_27),
.B2(n_31),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_51),
.A2(n_73),
.B1(n_34),
.B2(n_30),
.Y(n_75)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_47),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_52),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g78 ( 
.A(n_53),
.Y(n_78)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_57),
.B(n_61),
.Y(n_76)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_38),
.Y(n_61)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_41),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_64),
.B(n_70),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_39),
.A2(n_29),
.B1(n_26),
.B2(n_32),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_66),
.A2(n_67),
.B1(n_69),
.B2(n_74),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_44),
.A2(n_29),
.B1(n_24),
.B2(n_32),
.Y(n_67)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_40),
.Y(n_68)
);

HB1xp67_ASAP7_75t_L g90 ( 
.A(n_68),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_40),
.A2(n_23),
.B1(n_22),
.B2(n_24),
.Y(n_69)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_42),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_42),
.A2(n_17),
.B1(n_22),
.B2(n_23),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_43),
.A2(n_34),
.B1(n_30),
.B2(n_20),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_L g119 ( 
.A1(n_75),
.A2(n_59),
.B1(n_72),
.B2(n_19),
.Y(n_119)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_73),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_79),
.B(n_80),
.Y(n_109)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_62),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_55),
.B(n_20),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_81),
.B(n_88),
.Y(n_104)
);

BUFx12_ASAP7_75t_L g82 ( 
.A(n_50),
.Y(n_82)
);

CKINVDCx14_ASAP7_75t_R g115 ( 
.A(n_82),
.Y(n_115)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_63),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_83),
.B(n_84),
.Y(n_113)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_62),
.Y(n_84)
);

A2O1A1Ixp33_ASAP7_75t_L g85 ( 
.A1(n_56),
.A2(n_20),
.B(n_37),
.C(n_36),
.Y(n_85)
);

NAND3xp33_ASAP7_75t_L g122 ( 
.A(n_85),
.B(n_35),
.C(n_36),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_55),
.B(n_20),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_68),
.A2(n_48),
.B1(n_43),
.B2(n_21),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_89),
.A2(n_59),
.B1(n_72),
.B2(n_28),
.Y(n_118)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_63),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_91),
.B(n_92),
.Y(n_124)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_71),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_71),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_93),
.B(n_95),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_57),
.A2(n_48),
.B1(n_28),
.B2(n_34),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_94),
.A2(n_79),
.B1(n_75),
.B2(n_85),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_52),
.Y(n_95)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_56),
.Y(n_96)
);

INVx1_ASAP7_75t_SL g116 ( 
.A(n_96),
.Y(n_116)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_50),
.Y(n_97)
);

BUFx2_ASAP7_75t_L g129 ( 
.A(n_97),
.Y(n_129)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_49),
.Y(n_98)
);

INVx4_ASAP7_75t_L g126 ( 
.A(n_98),
.Y(n_126)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_54),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_100),
.A2(n_35),
.B1(n_16),
.B2(n_15),
.Y(n_123)
);

FAx1_ASAP7_75t_SL g101 ( 
.A(n_81),
.B(n_64),
.CI(n_37),
.CON(n_101),
.SN(n_101)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_101),
.B(n_106),
.Y(n_134)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_90),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_102),
.B(n_127),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_103),
.A2(n_111),
.B1(n_89),
.B2(n_91),
.Y(n_131)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_88),
.B(n_99),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_SL g155 ( 
.A1(n_105),
.A2(n_108),
.B(n_114),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_99),
.B(n_65),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_L g107 ( 
.A1(n_78),
.A2(n_60),
.B1(n_70),
.B2(n_61),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_107),
.A2(n_112),
.B1(n_118),
.B2(n_119),
.Y(n_132)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_86),
.B(n_28),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_87),
.Y(n_110)
);

INVxp33_ASAP7_75t_L g150 ( 
.A(n_110),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_78),
.A2(n_60),
.B1(n_65),
.B2(n_58),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_L g112 ( 
.A1(n_96),
.A2(n_58),
.B1(n_54),
.B2(n_59),
.Y(n_112)
);

AND2x2_ASAP7_75t_SL g114 ( 
.A(n_87),
.B(n_52),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_76),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_117),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_86),
.B(n_52),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_120),
.B(n_121),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_76),
.B(n_0),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_L g136 ( 
.A1(n_122),
.A2(n_128),
.B(n_93),
.Y(n_136)
);

CKINVDCx16_ASAP7_75t_R g133 ( 
.A(n_123),
.Y(n_133)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_98),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_95),
.B(n_0),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_L g130 ( 
.A1(n_104),
.A2(n_94),
.B(n_84),
.Y(n_130)
);

MAJx2_ASAP7_75t_L g179 ( 
.A(n_130),
.B(n_116),
.C(n_126),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_131),
.A2(n_142),
.B1(n_147),
.B2(n_149),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_136),
.B(n_137),
.Y(n_173)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_109),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_104),
.B(n_100),
.Y(n_138)
);

CKINVDCx16_ASAP7_75t_R g185 ( 
.A(n_138),
.Y(n_185)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_109),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_139),
.B(n_141),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_114),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_140),
.Y(n_178)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_125),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_103),
.A2(n_83),
.B1(n_77),
.B2(n_97),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_106),
.A2(n_77),
.B1(n_92),
.B2(n_80),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_143),
.A2(n_145),
.B1(n_108),
.B2(n_111),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_105),
.A2(n_82),
.B1(n_35),
.B2(n_2),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_121),
.B(n_82),
.Y(n_146)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_146),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_105),
.A2(n_82),
.B1(n_1),
.B2(n_2),
.Y(n_147)
);

AOI21xp5_ASAP7_75t_L g148 ( 
.A1(n_114),
.A2(n_0),
.B(n_1),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_L g167 ( 
.A1(n_148),
.A2(n_108),
.B(n_113),
.Y(n_167)
);

AO21x2_ASAP7_75t_L g149 ( 
.A1(n_114),
.A2(n_1),
.B(n_2),
.Y(n_149)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_125),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_151),
.B(n_6),
.Y(n_186)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_129),
.Y(n_152)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_152),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_120),
.B(n_1),
.C(n_2),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_153),
.B(n_115),
.C(n_124),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_105),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_154),
.A2(n_107),
.B1(n_118),
.B2(n_112),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_101),
.B(n_4),
.Y(n_157)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_157),
.Y(n_165)
);

NAND2x1_ASAP7_75t_L g159 ( 
.A(n_140),
.B(n_101),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_SL g212 ( 
.A1(n_159),
.A2(n_168),
.B(n_171),
.Y(n_212)
);

BUFx24_ASAP7_75t_SL g161 ( 
.A(n_156),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_161),
.B(n_162),
.Y(n_189)
);

O2A1O1Ixp33_ASAP7_75t_L g163 ( 
.A1(n_149),
.A2(n_101),
.B(n_122),
.C(n_128),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_L g201 ( 
.A1(n_163),
.A2(n_164),
.B(n_167),
.Y(n_201)
);

OR2x2_ASAP7_75t_L g164 ( 
.A(n_149),
.B(n_108),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_166),
.A2(n_177),
.B1(n_181),
.B2(n_184),
.Y(n_196)
);

AND2x2_ASAP7_75t_SL g168 ( 
.A(n_140),
.B(n_126),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_138),
.B(n_113),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_169),
.B(n_170),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_156),
.B(n_127),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_L g171 ( 
.A1(n_134),
.A2(n_124),
.B(n_115),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_135),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_172),
.B(n_174),
.Y(n_209)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_135),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_175),
.B(n_180),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_134),
.A2(n_116),
.B1(n_102),
.B2(n_126),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_SL g195 ( 
.A(n_179),
.B(n_145),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_157),
.B(n_129),
.Y(n_180)
);

OAI22x1_ASAP7_75t_SL g181 ( 
.A1(n_149),
.A2(n_116),
.B1(n_129),
.B2(n_7),
.Y(n_181)
);

OAI32xp33_ASAP7_75t_L g182 ( 
.A1(n_149),
.A2(n_5),
.A3(n_6),
.B1(n_8),
.B2(n_9),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_182),
.B(n_184),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_130),
.A2(n_6),
.B1(n_8),
.B2(n_9),
.Y(n_184)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_186),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_170),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_188),
.B(n_190),
.Y(n_227)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_177),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_SL g192 ( 
.A(n_165),
.B(n_141),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_192),
.B(n_193),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_176),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_194),
.B(n_207),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_195),
.B(n_162),
.Y(n_215)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_168),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_197),
.B(n_198),
.Y(n_235)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_169),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_159),
.B(n_155),
.Y(n_199)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_199),
.B(n_183),
.Y(n_222)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_168),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_200),
.B(n_206),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_159),
.A2(n_149),
.B1(n_133),
.B2(n_155),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_L g216 ( 
.A1(n_202),
.A2(n_163),
.B(n_185),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_L g203 ( 
.A1(n_173),
.A2(n_148),
.B(n_149),
.Y(n_203)
);

AOI21xp5_ASAP7_75t_L g226 ( 
.A1(n_203),
.A2(n_164),
.B(n_158),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_183),
.A2(n_130),
.B1(n_143),
.B2(n_132),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_204),
.A2(n_131),
.B1(n_142),
.B2(n_179),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_160),
.B(n_150),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_205),
.Y(n_232)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_168),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_178),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_171),
.B(n_136),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_210),
.B(n_211),
.C(n_185),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_178),
.B(n_175),
.C(n_167),
.Y(n_211)
);

HB1xp67_ASAP7_75t_L g213 ( 
.A(n_181),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_213),
.B(n_166),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_SL g214 ( 
.A1(n_179),
.A2(n_139),
.B(n_137),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_SL g237 ( 
.A1(n_214),
.A2(n_146),
.B(n_186),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_215),
.B(n_222),
.Y(n_257)
);

AOI21xp5_ASAP7_75t_L g254 ( 
.A1(n_216),
.A2(n_226),
.B(n_237),
.Y(n_254)
);

HB1xp67_ASAP7_75t_L g217 ( 
.A(n_197),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_217),
.B(n_160),
.Y(n_248)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_191),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_218),
.B(n_220),
.Y(n_246)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_191),
.Y(n_220)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_221),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_223),
.B(n_228),
.C(n_231),
.Y(n_265)
);

OAI22xp33_ASAP7_75t_SL g224 ( 
.A1(n_190),
.A2(n_158),
.B1(n_165),
.B2(n_151),
.Y(n_224)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_224),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_SL g225 ( 
.A(n_198),
.B(n_180),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_225),
.B(n_188),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_211),
.B(n_174),
.C(n_172),
.Y(n_228)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_206),
.Y(n_230)
);

INVx11_ASAP7_75t_L g247 ( 
.A(n_230),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_199),
.B(n_147),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_L g233 ( 
.A1(n_200),
.A2(n_164),
.B1(n_133),
.B2(n_154),
.Y(n_233)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_233),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_195),
.B(n_201),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_234),
.B(n_210),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_209),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_236),
.B(n_238),
.Y(n_250)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_196),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_196),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_239),
.B(n_194),
.Y(n_263)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_241),
.Y(n_259)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_242),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_238),
.A2(n_204),
.B1(n_212),
.B2(n_214),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_244),
.A2(n_249),
.B1(n_258),
.B2(n_233),
.Y(n_273)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_248),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_L g249 ( 
.A1(n_239),
.A2(n_230),
.B1(n_229),
.B2(n_240),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_225),
.Y(n_251)
);

AOI21xp5_ASAP7_75t_L g268 ( 
.A1(n_251),
.A2(n_255),
.B(n_260),
.Y(n_268)
);

XNOR2x1_ASAP7_75t_L g252 ( 
.A(n_222),
.B(n_212),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_SL g277 ( 
.A(n_252),
.B(n_203),
.Y(n_277)
);

BUFx2_ASAP7_75t_L g253 ( 
.A(n_232),
.Y(n_253)
);

INVxp67_ASAP7_75t_L g267 ( 
.A(n_253),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_SL g255 ( 
.A(n_236),
.B(n_189),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_221),
.A2(n_202),
.B1(n_201),
.B2(n_208),
.Y(n_258)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_235),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_261),
.B(n_234),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_219),
.Y(n_262)
);

OAI21xp5_ASAP7_75t_SL g283 ( 
.A1(n_262),
.A2(n_263),
.B(n_264),
.Y(n_283)
);

INVxp67_ASAP7_75t_SL g264 ( 
.A(n_232),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_265),
.B(n_228),
.C(n_223),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_266),
.B(n_271),
.C(n_272),
.Y(n_285)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_269),
.B(n_270),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_257),
.B(n_215),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_265),
.B(n_208),
.C(n_231),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_257),
.B(n_218),
.C(n_220),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_273),
.A2(n_250),
.B1(n_245),
.B2(n_259),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_252),
.B(n_227),
.C(n_237),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_274),
.B(n_277),
.C(n_279),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_L g276 ( 
.A1(n_243),
.A2(n_226),
.B1(n_216),
.B2(n_187),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_276),
.A2(n_256),
.B1(n_245),
.B2(n_263),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_243),
.A2(n_187),
.B1(n_182),
.B2(n_132),
.Y(n_278)
);

CKINVDCx16_ASAP7_75t_R g290 ( 
.A(n_278),
.Y(n_290)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_261),
.B(n_153),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_SL g281 ( 
.A(n_262),
.B(n_153),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_SL g299 ( 
.A(n_281),
.B(n_251),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_258),
.B(n_152),
.C(n_144),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_282),
.B(n_284),
.C(n_254),
.Y(n_300)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_244),
.B(n_11),
.Y(n_284)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_268),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_286),
.B(n_288),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_287),
.A2(n_292),
.B1(n_246),
.B2(n_275),
.Y(n_301)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_284),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_267),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_289),
.B(n_291),
.Y(n_308)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_282),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_274),
.A2(n_250),
.B1(n_256),
.B2(n_259),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_267),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_SL g313 ( 
.A(n_293),
.B(n_295),
.Y(n_313)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_294),
.Y(n_305)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_272),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_283),
.A2(n_254),
.B1(n_246),
.B2(n_260),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g314 ( 
.A(n_298),
.B(n_299),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_300),
.B(n_271),
.C(n_266),
.Y(n_303)
);

XOR2xp5_ASAP7_75t_L g317 ( 
.A(n_301),
.B(n_303),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_SL g302 ( 
.A(n_292),
.B(n_280),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_SL g316 ( 
.A(n_302),
.B(n_306),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_SL g306 ( 
.A(n_286),
.B(n_279),
.Y(n_306)
);

AOI22xp33_ASAP7_75t_SL g307 ( 
.A1(n_291),
.A2(n_247),
.B1(n_277),
.B2(n_253),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_SL g323 ( 
.A1(n_307),
.A2(n_294),
.B1(n_10),
.B2(n_9),
.Y(n_323)
);

XOR2xp5_ASAP7_75t_L g309 ( 
.A(n_297),
.B(n_269),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_309),
.B(n_297),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_285),
.B(n_270),
.C(n_247),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_310),
.B(n_296),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_287),
.A2(n_6),
.B1(n_8),
.B2(n_9),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_311),
.B(n_300),
.Y(n_319)
);

NOR2xp67_ASAP7_75t_L g312 ( 
.A(n_298),
.B(n_11),
.Y(n_312)
);

AOI21x1_ASAP7_75t_L g324 ( 
.A1(n_312),
.A2(n_12),
.B(n_13),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_L g331 ( 
.A(n_315),
.B(n_320),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_SL g318 ( 
.A(n_310),
.B(n_290),
.Y(n_318)
);

AOI21xp5_ASAP7_75t_L g326 ( 
.A1(n_318),
.A2(n_321),
.B(n_323),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_SL g329 ( 
.A(n_319),
.B(n_320),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_309),
.B(n_285),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_L g322 ( 
.A(n_303),
.B(n_296),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_SL g328 ( 
.A(n_322),
.B(n_324),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_316),
.B(n_314),
.Y(n_325)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_325),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_317),
.B(n_313),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_327),
.B(n_329),
.Y(n_333)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_317),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_330),
.B(n_332),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_SL g332 ( 
.A(n_315),
.B(n_304),
.Y(n_332)
);

AO21x1_ASAP7_75t_L g334 ( 
.A1(n_329),
.A2(n_305),
.B(n_301),
.Y(n_334)
);

NOR3xp33_ASAP7_75t_L g339 ( 
.A(n_334),
.B(n_335),
.C(n_308),
.Y(n_339)
);

AOI22xp5_ASAP7_75t_L g335 ( 
.A1(n_328),
.A2(n_304),
.B1(n_308),
.B2(n_311),
.Y(n_335)
);

OAI21xp5_ASAP7_75t_SL g338 ( 
.A1(n_336),
.A2(n_326),
.B(n_331),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_SL g340 ( 
.A(n_338),
.B(n_339),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_340),
.B(n_333),
.C(n_337),
.Y(n_341)
);

OAI321xp33_ASAP7_75t_L g342 ( 
.A1(n_341),
.A2(n_336),
.A3(n_13),
.B1(n_14),
.B2(n_16),
.C(n_10),
.Y(n_342)
);

AOI21xp5_ASAP7_75t_SL g343 ( 
.A1(n_342),
.A2(n_14),
.B(n_10),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_343),
.B(n_10),
.Y(n_344)
);


endmodule