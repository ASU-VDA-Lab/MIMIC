module fake_jpeg_21594_n_120 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_120);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_120;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_12),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_33),
.Y(n_40)
);

BUFx12_ASAP7_75t_L g41 ( 
.A(n_4),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_9),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_SL g43 ( 
.A(n_8),
.B(n_37),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_14),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_27),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_5),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_20),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_15),
.Y(n_48)
);

INVx1_ASAP7_75t_SL g49 ( 
.A(n_17),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_26),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_31),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_18),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_34),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_13),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_30),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_55),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_57),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_43),
.B(n_0),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_58),
.B(n_63),
.Y(n_74)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_46),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_59),
.B(n_61),
.Y(n_71)
);

INVx11_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_60),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_52),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_40),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_62),
.B(n_47),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_41),
.B(n_0),
.Y(n_63)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_40),
.Y(n_64)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_64),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_64),
.A2(n_48),
.B1(n_49),
.B2(n_53),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_65),
.A2(n_66),
.B1(n_1),
.B2(n_2),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_L g66 ( 
.A1(n_60),
.A2(n_47),
.B1(n_50),
.B2(n_51),
.Y(n_66)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_57),
.Y(n_67)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_67),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_68),
.B(n_75),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_57),
.B(n_43),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_72),
.B(n_54),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_58),
.B(n_56),
.Y(n_75)
);

INVx13_ASAP7_75t_L g76 ( 
.A(n_70),
.Y(n_76)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_76),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_78),
.B(n_81),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_SL g79 ( 
.A1(n_74),
.A2(n_45),
.B(n_44),
.Y(n_79)
);

XOR2xp5_ASAP7_75t_L g94 ( 
.A(n_79),
.B(n_80),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_71),
.B(n_42),
.C(n_39),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_73),
.A2(n_23),
.B1(n_36),
.B2(n_35),
.Y(n_81)
);

INVx1_ASAP7_75t_SL g83 ( 
.A(n_70),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_83),
.B(n_85),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_84),
.B(n_86),
.Y(n_96)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_66),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_69),
.B(n_1),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_65),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_87),
.B(n_89),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_72),
.B(n_2),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_88),
.B(n_6),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_71),
.Y(n_89)
);

OAI21xp33_ASAP7_75t_L g91 ( 
.A1(n_77),
.A2(n_3),
.B(n_4),
.Y(n_91)
);

AOI21xp5_ASAP7_75t_L g106 ( 
.A1(n_91),
.A2(n_98),
.B(n_99),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_77),
.B(n_3),
.Y(n_92)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_92),
.Y(n_105)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_97),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_86),
.B(n_7),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_82),
.B(n_10),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_76),
.B(n_11),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_100),
.A2(n_101),
.B1(n_24),
.B2(n_25),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_78),
.B(n_16),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_96),
.A2(n_19),
.B1(n_21),
.B2(n_22),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_103),
.B(n_104),
.Y(n_110)
);

HB1xp67_ASAP7_75t_L g104 ( 
.A(n_95),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_107),
.B(n_109),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_102),
.A2(n_93),
.B1(n_90),
.B2(n_94),
.Y(n_109)
);

OA21x2_ASAP7_75t_L g111 ( 
.A1(n_105),
.A2(n_102),
.B(n_29),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_111),
.B(n_28),
.Y(n_113)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_113),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_114),
.B(n_108),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_115),
.B(n_112),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_116),
.B(n_110),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_117),
.B(n_104),
.Y(n_118)
);

XOR2xp5_ASAP7_75t_L g119 ( 
.A(n_118),
.B(n_106),
.Y(n_119)
);

XOR2xp5_ASAP7_75t_L g120 ( 
.A(n_119),
.B(n_32),
.Y(n_120)
);


endmodule