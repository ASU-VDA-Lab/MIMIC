module fake_jpeg_15802_n_294 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_294);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_294;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_252;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_137;
wire n_74;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_187;
wire n_21;
wire n_57;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_91;
wire n_93;
wire n_54;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_270;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_265;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

INVx8_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

BUFx8_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_5),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

BUFx16f_ASAP7_75t_L g25 ( 
.A(n_16),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_11),
.Y(n_26)
);

BUFx10_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

BUFx12_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_SL g33 ( 
.A(n_16),
.B(n_10),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_4),
.Y(n_34)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_12),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_29),
.Y(n_36)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g37 ( 
.A(n_33),
.B(n_8),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_SL g50 ( 
.A(n_37),
.B(n_41),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_21),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_39),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_33),
.B(n_9),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_40),
.B(n_43),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_31),
.B(n_9),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_21),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_42),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_27),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_29),
.Y(n_44)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_44),
.Y(n_57)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_38),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_46),
.B(n_47),
.Y(n_78)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_38),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_39),
.A2(n_31),
.B1(n_35),
.B2(n_23),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_48),
.A2(n_49),
.B1(n_53),
.B2(n_60),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_39),
.A2(n_35),
.B1(n_23),
.B2(n_17),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_39),
.A2(n_35),
.B1(n_23),
.B2(n_17),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_52),
.A2(n_68),
.B1(n_24),
.B2(n_18),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_41),
.A2(n_17),
.B1(n_25),
.B2(n_26),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g55 ( 
.A(n_37),
.B(n_32),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_55),
.B(n_28),
.Y(n_85)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_43),
.Y(n_56)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_56),
.Y(n_81)
);

OR2x2_ASAP7_75t_L g58 ( 
.A(n_43),
.B(n_22),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_58),
.B(n_18),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_36),
.A2(n_25),
.B1(n_20),
.B2(n_26),
.Y(n_60)
);

HB1xp67_ASAP7_75t_L g61 ( 
.A(n_36),
.Y(n_61)
);

BUFx2_ASAP7_75t_L g74 ( 
.A(n_61),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_44),
.A2(n_25),
.B1(n_22),
.B2(n_32),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_62),
.A2(n_64),
.B1(n_18),
.B2(n_28),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_37),
.B(n_22),
.Y(n_63)
);

NAND3xp33_ASAP7_75t_L g79 ( 
.A(n_63),
.B(n_40),
.C(n_29),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_44),
.A2(n_25),
.B1(n_19),
.B2(n_20),
.Y(n_64)
);

AND2x2_ASAP7_75t_SL g65 ( 
.A(n_43),
.B(n_25),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_65),
.B(n_0),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_38),
.Y(n_66)
);

INVx3_ASAP7_75t_SL g72 ( 
.A(n_66),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_42),
.A2(n_19),
.B1(n_30),
.B2(n_34),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_L g70 ( 
.A1(n_48),
.A2(n_42),
.B1(n_21),
.B2(n_34),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_70),
.A2(n_71),
.B1(n_83),
.B2(n_87),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_49),
.A2(n_42),
.B1(n_34),
.B2(n_30),
.Y(n_71)
);

XNOR2xp5_ASAP7_75t_SL g126 ( 
.A(n_73),
.B(n_82),
.Y(n_126)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_67),
.Y(n_75)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_75),
.Y(n_106)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_45),
.Y(n_76)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_76),
.Y(n_112)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_45),
.Y(n_77)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_77),
.Y(n_127)
);

OAI21x1_ASAP7_75t_L g120 ( 
.A1(n_79),
.A2(n_92),
.B(n_95),
.Y(n_120)
);

OA22x2_ASAP7_75t_L g80 ( 
.A1(n_56),
.A2(n_18),
.B1(n_21),
.B2(n_24),
.Y(n_80)
);

OA22x2_ASAP7_75t_L g117 ( 
.A1(n_80),
.A2(n_101),
.B1(n_56),
.B2(n_51),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_SL g82 ( 
.A(n_50),
.B(n_40),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_65),
.A2(n_34),
.B1(n_30),
.B2(n_24),
.Y(n_83)
);

AO22x1_ASAP7_75t_L g84 ( 
.A1(n_46),
.A2(n_18),
.B1(n_24),
.B2(n_30),
.Y(n_84)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_84),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_85),
.B(n_86),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_55),
.B(n_28),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_65),
.A2(n_11),
.B1(n_16),
.B2(n_15),
.Y(n_88)
);

XNOR2xp5_ASAP7_75t_L g102 ( 
.A(n_88),
.B(n_94),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_61),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_89),
.B(n_90),
.Y(n_110)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_51),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_91),
.A2(n_10),
.B1(n_12),
.B2(n_14),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_58),
.B(n_29),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_93),
.B(n_99),
.Y(n_103)
);

XOR2xp5_ASAP7_75t_L g94 ( 
.A(n_54),
.B(n_28),
.Y(n_94)
);

OR2x2_ASAP7_75t_L g95 ( 
.A(n_63),
.B(n_28),
.Y(n_95)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_67),
.Y(n_96)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_96),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_54),
.B(n_27),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_97),
.B(n_98),
.Y(n_113)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_57),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_53),
.B(n_0),
.Y(n_99)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_57),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_100),
.B(n_47),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_L g101 ( 
.A1(n_60),
.A2(n_47),
.B1(n_46),
.B2(n_68),
.Y(n_101)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_78),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_104),
.B(n_115),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_81),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_105),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_L g107 ( 
.A(n_94),
.B(n_52),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_107),
.B(n_69),
.C(n_82),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_93),
.B(n_58),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_114),
.B(n_121),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_81),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g134 ( 
.A(n_117),
.B(n_80),
.Y(n_134)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_98),
.Y(n_118)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_118),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_119),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_92),
.B(n_50),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_92),
.B(n_65),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_SL g144 ( 
.A(n_122),
.B(n_124),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_75),
.B(n_27),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_123),
.B(n_27),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_73),
.B(n_66),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_95),
.B(n_66),
.Y(n_125)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_125),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g140 ( 
.A(n_128),
.Y(n_140)
);

INVx2_ASAP7_75t_SL g129 ( 
.A(n_72),
.Y(n_129)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_129),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_SL g190 ( 
.A(n_130),
.B(n_142),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g131 ( 
.A(n_102),
.B(n_69),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_131),
.B(n_135),
.C(n_155),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_134),
.A2(n_146),
.B1(n_148),
.B2(n_154),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g135 ( 
.A(n_102),
.B(n_99),
.Y(n_135)
);

INVxp33_ASAP7_75t_SL g136 ( 
.A(n_105),
.Y(n_136)
);

INVx1_ASAP7_75t_SL g170 ( 
.A(n_136),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_116),
.A2(n_71),
.B1(n_83),
.B2(n_87),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_137),
.A2(n_158),
.B1(n_124),
.B2(n_107),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_SL g139 ( 
.A1(n_125),
.A2(n_99),
.B(n_89),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g180 ( 
.A(n_139),
.Y(n_180)
);

OAI32xp33_ASAP7_75t_L g142 ( 
.A1(n_103),
.A2(n_88),
.A3(n_80),
.B1(n_84),
.B2(n_100),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_SL g143 ( 
.A1(n_122),
.A2(n_80),
.B(n_84),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_143),
.B(n_147),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_109),
.A2(n_96),
.B1(n_77),
.B2(n_76),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_SL g147 ( 
.A1(n_114),
.A2(n_74),
.B(n_29),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_116),
.A2(n_90),
.B1(n_74),
.B2(n_59),
.Y(n_148)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_118),
.Y(n_150)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_150),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_L g152 ( 
.A1(n_120),
.A2(n_74),
.B(n_27),
.Y(n_152)
);

XOR2xp5_ASAP7_75t_L g176 ( 
.A(n_152),
.B(n_156),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_153),
.B(n_159),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_L g154 ( 
.A1(n_117),
.A2(n_72),
.B1(n_59),
.B2(n_51),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_126),
.B(n_72),
.C(n_59),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_126),
.B(n_29),
.C(n_27),
.Y(n_156)
);

OR2x2_ASAP7_75t_L g157 ( 
.A(n_103),
.B(n_0),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_157),
.B(n_106),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_117),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_113),
.B(n_6),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_108),
.Y(n_160)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_160),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_160),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_162),
.B(n_163),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_149),
.B(n_104),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_SL g199 ( 
.A(n_165),
.B(n_169),
.Y(n_199)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_132),
.Y(n_166)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_166),
.Y(n_206)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_132),
.Y(n_167)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_167),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_150),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_168),
.B(n_173),
.Y(n_198)
);

NOR2x1_ASAP7_75t_L g169 ( 
.A(n_139),
.B(n_111),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_171),
.A2(n_134),
.B1(n_131),
.B2(n_155),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_133),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_145),
.Y(n_174)
);

CKINVDCx16_ASAP7_75t_R g193 ( 
.A(n_174),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_133),
.B(n_110),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_175),
.B(n_181),
.Y(n_212)
);

BUFx24_ASAP7_75t_SL g181 ( 
.A(n_151),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_141),
.B(n_106),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_182),
.B(n_183),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_141),
.B(n_121),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_SL g184 ( 
.A(n_157),
.B(n_117),
.Y(n_184)
);

AOI21xp33_ASAP7_75t_L g210 ( 
.A1(n_184),
.A2(n_127),
.B(n_129),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_145),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_SL g203 ( 
.A1(n_185),
.A2(n_188),
.B(n_112),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_138),
.B(n_115),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_186),
.B(n_187),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_138),
.B(n_108),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_148),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_151),
.B(n_144),
.Y(n_189)
);

FAx1_ASAP7_75t_SL g191 ( 
.A(n_189),
.B(n_130),
.CI(n_135),
.CON(n_191),
.SN(n_191)
);

NOR2xp33_ASAP7_75t_SL g217 ( 
.A(n_191),
.B(n_176),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_194),
.A2(n_209),
.B1(n_170),
.B2(n_173),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_178),
.B(n_156),
.C(n_144),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_195),
.B(n_200),
.C(n_201),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_L g197 ( 
.A1(n_180),
.A2(n_169),
.B(n_184),
.Y(n_197)
);

AOI21xp5_ASAP7_75t_L g226 ( 
.A1(n_197),
.A2(n_207),
.B(n_211),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_178),
.B(n_147),
.C(n_152),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_190),
.B(n_172),
.Y(n_201)
);

XNOR2x1_ASAP7_75t_L g202 ( 
.A(n_190),
.B(n_157),
.Y(n_202)
);

AOI321xp33_ASAP7_75t_L g235 ( 
.A1(n_202),
.A2(n_210),
.A3(n_4),
.B1(n_5),
.B2(n_6),
.C(n_7),
.Y(n_235)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_203),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_180),
.A2(n_146),
.B1(n_140),
.B2(n_134),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_204),
.A2(n_161),
.B1(n_164),
.B2(n_129),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_L g207 ( 
.A1(n_172),
.A2(n_140),
.B(n_142),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_171),
.A2(n_137),
.B1(n_158),
.B2(n_143),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_L g211 ( 
.A1(n_165),
.A2(n_183),
.B(n_182),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_L g213 ( 
.A1(n_188),
.A2(n_1),
.B(n_2),
.Y(n_213)
);

AOI21xp5_ASAP7_75t_L g227 ( 
.A1(n_213),
.A2(n_1),
.B(n_2),
.Y(n_227)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_174),
.Y(n_214)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_214),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_209),
.A2(n_177),
.B1(n_170),
.B2(n_185),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_L g246 ( 
.A1(n_215),
.A2(n_229),
.B1(n_213),
.B2(n_193),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_196),
.B(n_168),
.Y(n_216)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_216),
.Y(n_236)
);

AOI321xp33_ASAP7_75t_L g237 ( 
.A1(n_217),
.A2(n_202),
.A3(n_191),
.B1(n_197),
.B2(n_211),
.C(n_199),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_200),
.B(n_176),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_218),
.B(n_222),
.C(n_232),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_220),
.B(n_214),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_196),
.B(n_162),
.Y(n_221)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_221),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_195),
.B(n_167),
.C(n_166),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_SL g238 ( 
.A(n_223),
.B(n_235),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_201),
.B(n_194),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_224),
.B(n_203),
.Y(n_240)
);

INVxp33_ASAP7_75t_L g225 ( 
.A(n_198),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_225),
.B(n_234),
.Y(n_245)
);

OAI21xp5_ASAP7_75t_SL g249 ( 
.A1(n_227),
.A2(n_206),
.B(n_7),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_192),
.B(n_179),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_SL g251 ( 
.A(n_228),
.B(n_233),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_207),
.A2(n_161),
.B1(n_164),
.B2(n_1),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_191),
.B(n_3),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_SL g233 ( 
.A(n_212),
.B(n_3),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_205),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_237),
.B(n_239),
.Y(n_256)
);

OAI322xp33_ASAP7_75t_L g239 ( 
.A1(n_232),
.A2(n_199),
.A3(n_205),
.B1(n_193),
.B2(n_204),
.C1(n_206),
.C2(n_208),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_240),
.B(n_247),
.C(n_250),
.Y(n_260)
);

OAI322xp33_ASAP7_75t_L g242 ( 
.A1(n_235),
.A2(n_226),
.A3(n_230),
.B1(n_216),
.B2(n_221),
.C1(n_224),
.C2(n_218),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_242),
.B(n_229),
.Y(n_253)
);

INVxp67_ASAP7_75t_L g244 ( 
.A(n_223),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_244),
.B(n_222),
.Y(n_257)
);

CKINVDCx14_ASAP7_75t_R g258 ( 
.A(n_246),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_SL g247 ( 
.A(n_226),
.B(n_208),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_248),
.B(n_13),
.Y(n_263)
);

AOI21xp5_ASAP7_75t_L g264 ( 
.A1(n_249),
.A2(n_13),
.B(n_238),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_219),
.B(n_4),
.Y(n_250)
);

OAI21xp5_ASAP7_75t_L g252 ( 
.A1(n_244),
.A2(n_227),
.B(n_215),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_SL g266 ( 
.A(n_252),
.B(n_253),
.Y(n_266)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_245),
.Y(n_254)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_254),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_251),
.B(n_231),
.Y(n_255)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_255),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_SL g268 ( 
.A(n_257),
.B(n_261),
.Y(n_268)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_236),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_259),
.B(n_248),
.Y(n_272)
);

OAI21xp5_ASAP7_75t_L g261 ( 
.A1(n_243),
.A2(n_225),
.B(n_219),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_241),
.B(n_14),
.C(n_10),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_262),
.B(n_264),
.C(n_238),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_263),
.B(n_256),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_264),
.B(n_256),
.Y(n_274)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_267),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_260),
.B(n_240),
.Y(n_269)
);

AND2x2_ASAP7_75t_L g280 ( 
.A(n_269),
.B(n_275),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_270),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_272),
.B(n_274),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_261),
.B(n_258),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_273),
.B(n_262),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_260),
.B(n_257),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_265),
.B(n_252),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_SL g287 ( 
.A(n_277),
.B(n_279),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_271),
.B(n_249),
.Y(n_279)
);

OAI21xp5_ASAP7_75t_L g283 ( 
.A1(n_282),
.A2(n_241),
.B(n_268),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_283),
.B(n_284),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_281),
.B(n_275),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_276),
.B(n_250),
.Y(n_285)
);

NOR4xp25_ASAP7_75t_L g290 ( 
.A(n_285),
.B(n_287),
.C(n_237),
.D(n_269),
.Y(n_290)
);

OAI21xp5_ASAP7_75t_L g286 ( 
.A1(n_280),
.A2(n_266),
.B(n_268),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_L g288 ( 
.A1(n_286),
.A2(n_278),
.B1(n_276),
.B2(n_266),
.Y(n_288)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_288),
.Y(n_292)
);

AOI21xp5_ASAP7_75t_SL g291 ( 
.A1(n_290),
.A2(n_289),
.B(n_247),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_291),
.B(n_13),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_293),
.B(n_292),
.Y(n_294)
);


endmodule