module real_jpeg_18009_n_19 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_19);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_19;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_541;
wire n_441;
wire n_557;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_553;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_366;
wire n_328;
wire n_456;
wire n_556;
wire n_259;
wire n_57;
wire n_507;
wire n_157;
wire n_560;
wire n_84;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_551;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_464;
wire n_423;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_550;
wire n_233;
wire n_73;
wire n_532;
wire n_516;
wire n_348;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_525;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_544;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_561;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_543;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_533;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_559;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_25;
wire n_480;
wire n_542;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_215;
wire n_176;
wire n_166;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_412;
wire n_120;
wire n_155;
wire n_405;
wire n_548;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_546;
wire n_531;
wire n_112;
wire n_554;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_558;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_330;
wire n_298;
wire n_450;
wire n_333;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_537;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_475;
wire n_74;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_534;
wire n_256;
wire n_520;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_545;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_502;
wire n_418;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_555;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_547;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_368;
wire n_100;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_549;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_468;
wire n_133;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_552;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

AOI21xp5_ASAP7_75t_L g19 ( 
.A1(n_0),
.A2(n_20),
.B(n_560),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g560 ( 
.A(n_0),
.B(n_561),
.Y(n_560)
);

AND2x2_ASAP7_75t_L g59 ( 
.A(n_1),
.B(n_60),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_1),
.B(n_78),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_1),
.B(n_91),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g129 ( 
.A(n_1),
.B(n_130),
.Y(n_129)
);

AOI22x1_ASAP7_75t_L g137 ( 
.A1(n_1),
.A2(n_3),
.B1(n_138),
.B2(n_142),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_1),
.B(n_185),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_1),
.B(n_250),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_1),
.B(n_223),
.Y(n_329)
);

CKINVDCx14_ASAP7_75t_R g357 ( 
.A(n_1),
.Y(n_357)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_2),
.Y(n_135)
);

BUFx5_ASAP7_75t_L g141 ( 
.A(n_2),
.Y(n_141)
);

BUFx5_ASAP7_75t_L g415 ( 
.A(n_2),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_3),
.B(n_193),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_3),
.B(n_202),
.Y(n_201)
);

AND2x2_ASAP7_75t_L g280 ( 
.A(n_3),
.B(n_281),
.Y(n_280)
);

AND2x2_ASAP7_75t_L g348 ( 
.A(n_3),
.B(n_349),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_3),
.B(n_384),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_3),
.B(n_436),
.Y(n_435)
);

AND2x2_ASAP7_75t_L g449 ( 
.A(n_3),
.B(n_450),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_3),
.B(n_475),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_4),
.B(n_168),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_4),
.B(n_368),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_SL g387 ( 
.A(n_4),
.B(n_388),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_4),
.B(n_432),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_4),
.B(n_468),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_SL g482 ( 
.A(n_4),
.B(n_483),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_SL g491 ( 
.A(n_4),
.B(n_492),
.Y(n_491)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_5),
.Y(n_39)
);

BUFx5_ASAP7_75t_L g44 ( 
.A(n_5),
.Y(n_44)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_5),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_5),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g221 ( 
.A(n_5),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_6),
.B(n_51),
.Y(n_127)
);

CKINVDCx16_ASAP7_75t_R g149 ( 
.A(n_6),
.Y(n_149)
);

AND2x4_ASAP7_75t_L g163 ( 
.A(n_6),
.B(n_164),
.Y(n_163)
);

AND2x2_ASAP7_75t_SL g182 ( 
.A(n_6),
.B(n_29),
.Y(n_182)
);

AND2x2_ASAP7_75t_L g209 ( 
.A(n_6),
.B(n_210),
.Y(n_209)
);

AND2x2_ASAP7_75t_L g283 ( 
.A(n_6),
.B(n_175),
.Y(n_283)
);

AND2x2_ASAP7_75t_L g364 ( 
.A(n_6),
.B(n_130),
.Y(n_364)
);

AND2x2_ASAP7_75t_L g414 ( 
.A(n_6),
.B(n_415),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_7),
.B(n_35),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_7),
.B(n_49),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_7),
.B(n_82),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_7),
.B(n_96),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g133 ( 
.A(n_7),
.B(n_134),
.Y(n_133)
);

AND2x2_ASAP7_75t_L g196 ( 
.A(n_7),
.B(n_197),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_7),
.B(n_246),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_7),
.B(n_326),
.Y(n_325)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_8),
.Y(n_109)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_8),
.Y(n_172)
);

BUFx5_ASAP7_75t_L g175 ( 
.A(n_8),
.Y(n_175)
);

BUFx6f_ASAP7_75t_L g187 ( 
.A(n_8),
.Y(n_187)
);

BUFx5_ASAP7_75t_L g246 ( 
.A(n_8),
.Y(n_246)
);

BUFx6f_ASAP7_75t_L g487 ( 
.A(n_8),
.Y(n_487)
);

AND2x2_ASAP7_75t_L g152 ( 
.A(n_9),
.B(n_153),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_9),
.B(n_28),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_9),
.B(n_219),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_9),
.B(n_233),
.Y(n_232)
);

AND2x2_ASAP7_75t_L g284 ( 
.A(n_9),
.B(n_285),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g406 ( 
.A(n_9),
.B(n_407),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_9),
.B(n_412),
.Y(n_411)
);

AND2x2_ASAP7_75t_L g451 ( 
.A(n_9),
.B(n_452),
.Y(n_451)
);

BUFx12f_ASAP7_75t_L g132 ( 
.A(n_10),
.Y(n_132)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_10),
.Y(n_159)
);

BUFx4f_ASAP7_75t_L g199 ( 
.A(n_10),
.Y(n_199)
);

BUFx6f_ASAP7_75t_L g241 ( 
.A(n_10),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_11),
.B(n_28),
.Y(n_27)
);

AND2x2_ASAP7_75t_SL g31 ( 
.A(n_11),
.B(n_32),
.Y(n_31)
);

INVx1_ASAP7_75t_SL g45 ( 
.A(n_11),
.Y(n_45)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_11),
.B(n_70),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g195 ( 
.A(n_11),
.B(n_134),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g555 ( 
.A(n_11),
.B(n_556),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_12),
.B(n_65),
.Y(n_64)
);

INVxp33_ASAP7_75t_L g105 ( 
.A(n_12),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g156 ( 
.A(n_12),
.B(n_157),
.Y(n_156)
);

AND2x2_ASAP7_75t_L g174 ( 
.A(n_12),
.B(n_175),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_12),
.B(n_215),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_12),
.B(n_223),
.Y(n_248)
);

AND2x2_ASAP7_75t_SL g277 ( 
.A(n_12),
.B(n_278),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_SL g312 ( 
.A(n_12),
.B(n_313),
.Y(n_312)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_13),
.Y(n_99)
);

BUFx3_ASAP7_75t_L g155 ( 
.A(n_13),
.Y(n_155)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_13),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g561 ( 
.A(n_14),
.Y(n_561)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_15),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g207 ( 
.A(n_15),
.Y(n_207)
);

BUFx3_ASAP7_75t_L g216 ( 
.A(n_15),
.Y(n_216)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_15),
.Y(n_253)
);

BUFx3_ASAP7_75t_L g285 ( 
.A(n_15),
.Y(n_285)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_15),
.Y(n_328)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_16),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_16),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_17),
.B(n_101),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g170 ( 
.A(n_17),
.B(n_171),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_17),
.B(n_205),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_17),
.B(n_223),
.Y(n_222)
);

AND2x2_ASAP7_75t_L g230 ( 
.A(n_17),
.B(n_29),
.Y(n_230)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_17),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_17),
.B(n_322),
.Y(n_321)
);

AND2x2_ASAP7_75t_L g365 ( 
.A(n_17),
.B(n_141),
.Y(n_365)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_18),
.Y(n_53)
);

BUFx5_ASAP7_75t_L g67 ( 
.A(n_18),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g169 ( 
.A(n_18),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_550),
.Y(n_20)
);

OAI21x1_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_116),
.B(n_549),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_23),
.Y(n_22)
);

NAND2x1p5_ASAP7_75t_R g23 ( 
.A(n_24),
.B(n_73),
.Y(n_23)
);

OR2x2_ASAP7_75t_L g549 ( 
.A(n_24),
.B(n_73),
.Y(n_549)
);

XOR2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_54),
.Y(n_24)
);

XNOR2xp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_40),
.Y(n_25)
);

MAJIxp5_ASAP7_75t_L g558 ( 
.A(n_26),
.B(n_40),
.C(n_54),
.Y(n_558)
);

MAJIxp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_31),
.C(n_34),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g41 ( 
.A1(n_27),
.A2(n_42),
.B1(n_46),
.B2(n_47),
.Y(n_41)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_27),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g57 ( 
.A1(n_27),
.A2(n_31),
.B1(n_46),
.B2(n_58),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_SL g553 ( 
.A(n_27),
.B(n_42),
.C(n_48),
.Y(n_553)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx1_ASAP7_75t_SL g58 ( 
.A(n_31),
.Y(n_58)
);

MAJIxp5_ASAP7_75t_L g63 ( 
.A(n_31),
.B(n_64),
.C(n_68),
.Y(n_63)
);

AOI22x1_ASAP7_75t_SL g111 ( 
.A1(n_31),
.A2(n_58),
.B1(n_68),
.B2(n_69),
.Y(n_111)
);

INVx3_ASAP7_75t_L g224 ( 
.A(n_32),
.Y(n_224)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

XOR2xp5_ASAP7_75t_L g56 ( 
.A(n_34),
.B(n_57),
.Y(n_56)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

HB1xp67_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

XNOR2xp5_ASAP7_75t_L g40 ( 
.A(n_41),
.B(n_48),
.Y(n_40)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_42),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g554 ( 
.A1(n_42),
.A2(n_47),
.B1(n_555),
.B2(n_557),
.Y(n_554)
);

NOR2xp33_ASAP7_75t_SL g42 ( 
.A(n_43),
.B(n_45),
.Y(n_42)
);

BUFx2_ASAP7_75t_L g106 ( 
.A(n_43),
.Y(n_106)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

OR2x2_ASAP7_75t_L g107 ( 
.A(n_45),
.B(n_108),
.Y(n_107)
);

OR2x2_ASAP7_75t_L g239 ( 
.A(n_45),
.B(n_240),
.Y(n_239)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g556 ( 
.A(n_51),
.Y(n_556)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_52),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_53),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g54 ( 
.A(n_55),
.B(n_59),
.C(n_63),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_55),
.A2(n_56),
.B1(n_114),
.B2(n_115),
.Y(n_113)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

XNOR2xp5_ASAP7_75t_SL g115 ( 
.A(n_59),
.B(n_63),
.Y(n_115)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

XOR2x1_ASAP7_75t_L g110 ( 
.A(n_64),
.B(n_111),
.Y(n_110)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

BUFx2_ASAP7_75t_L g193 ( 
.A(n_67),
.Y(n_193)
);

AOI22xp33_ASAP7_75t_SL g516 ( 
.A1(n_68),
.A2(n_69),
.B1(n_107),
.B2(n_310),
.Y(n_516)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_SL g103 ( 
.A(n_69),
.B(n_104),
.C(n_107),
.Y(n_103)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_72),
.Y(n_166)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_72),
.Y(n_386)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_74),
.B(n_112),
.C(n_113),
.Y(n_73)
);

XNOR2xp5_ASAP7_75t_L g523 ( 
.A(n_74),
.B(n_524),
.Y(n_523)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_75),
.B(n_103),
.C(n_110),
.Y(n_74)
);

XOR2xp5_ASAP7_75t_L g521 ( 
.A(n_75),
.B(n_522),
.Y(n_521)
);

XNOR2xp5_ASAP7_75t_L g75 ( 
.A(n_76),
.B(n_88),
.Y(n_75)
);

XNOR2xp5_ASAP7_75t_L g76 ( 
.A(n_77),
.B(n_81),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_77),
.B(n_81),
.C(n_88),
.Y(n_112)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx4_ASAP7_75t_L g203 ( 
.A(n_79),
.Y(n_203)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g389 ( 
.A(n_86),
.Y(n_389)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_87),
.Y(n_93)
);

BUFx5_ASAP7_75t_L g145 ( 
.A(n_87),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g317 ( 
.A(n_87),
.Y(n_317)
);

BUFx6f_ASAP7_75t_L g355 ( 
.A(n_87),
.Y(n_355)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_94),
.C(n_100),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g512 ( 
.A1(n_89),
.A2(n_90),
.B1(n_94),
.B2(n_95),
.Y(n_512)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g434 ( 
.A(n_99),
.Y(n_434)
);

XNOR2x1_ASAP7_75t_L g511 ( 
.A(n_100),
.B(n_512),
.Y(n_511)
);

INVx6_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_L g522 ( 
.A(n_103),
.B(n_110),
.Y(n_522)
);

XNOR2xp5_ASAP7_75t_SL g515 ( 
.A(n_104),
.B(n_516),
.Y(n_515)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_106),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_L g309 ( 
.A1(n_107),
.A2(n_239),
.B1(n_310),
.B2(n_311),
.Y(n_309)
);

INVx1_ASAP7_75t_SL g310 ( 
.A(n_107),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g517 ( 
.A(n_107),
.B(n_311),
.C(n_312),
.Y(n_517)
);

BUFx3_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

XNOR2xp5_ASAP7_75t_L g524 ( 
.A(n_112),
.B(n_113),
.Y(n_524)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

AOI21x1_ASAP7_75t_L g116 ( 
.A1(n_117),
.A2(n_505),
.B(n_544),
.Y(n_116)
);

AO21x2_ASAP7_75t_L g117 ( 
.A1(n_118),
.A2(n_333),
.B(n_502),
.Y(n_117)
);

NOR2xp67_ASAP7_75t_SL g118 ( 
.A(n_119),
.B(n_292),
.Y(n_118)
);

AND2x2_ASAP7_75t_L g119 ( 
.A(n_120),
.B(n_256),
.Y(n_119)
);

OR2x2_ASAP7_75t_L g503 ( 
.A(n_120),
.B(n_256),
.Y(n_503)
);

XNOR2xp5_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_188),
.Y(n_120)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_121),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_160),
.C(n_177),
.Y(n_121)
);

INVxp33_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

XNOR2x1_ASAP7_75t_SL g258 ( 
.A(n_123),
.B(n_259),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_136),
.C(n_146),
.Y(n_123)
);

XNOR2xp5_ASAP7_75t_L g369 ( 
.A(n_124),
.B(n_370),
.Y(n_369)
);

XNOR2xp5_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_128),
.Y(n_124)
);

MAJx2_ASAP7_75t_L g513 ( 
.A(n_125),
.B(n_230),
.C(n_304),
.Y(n_513)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_126),
.B(n_230),
.Y(n_301)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_127),
.B(n_129),
.C(n_133),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_133),
.Y(n_128)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g278 ( 
.A(n_134),
.Y(n_278)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx2_ASAP7_75t_L g361 ( 
.A(n_135),
.Y(n_361)
);

AOI22xp5_ASAP7_75t_SL g370 ( 
.A1(n_136),
.A2(n_137),
.B1(n_146),
.B2(n_371),
.Y(n_370)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

AOI21xp5_ASAP7_75t_L g347 ( 
.A1(n_137),
.A2(n_348),
.B(n_356),
.Y(n_347)
);

INVx4_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVx6_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

BUFx12f_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

HB1xp67_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVx2_ASAP7_75t_SL g144 ( 
.A(n_145),
.Y(n_144)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_146),
.Y(n_371)
);

MAJx2_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_152),
.C(n_156),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_147),
.A2(n_148),
.B1(n_237),
.B2(n_238),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_147),
.A2(n_148),
.B1(n_156),
.B2(n_270),
.Y(n_269)
);

INVx1_ASAP7_75t_SL g147 ( 
.A(n_148),
.Y(n_147)
);

MAJx2_ASAP7_75t_L g302 ( 
.A(n_148),
.B(n_195),
.C(n_239),
.Y(n_302)
);

OR2x2_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_150),
.Y(n_148)
);

INVx6_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

INVx3_ASAP7_75t_L g323 ( 
.A(n_151),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_152),
.B(n_269),
.Y(n_268)
);

INVx3_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_155),
.Y(n_282)
);

INVx11_ASAP7_75t_SL g270 ( 
.A(n_156),
.Y(n_270)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

HB1xp67_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_161),
.A2(n_177),
.B1(n_178),
.B2(n_260),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_161),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_173),
.C(n_176),
.Y(n_161)
);

XOR2x2_ASAP7_75t_L g286 ( 
.A(n_162),
.B(n_287),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_167),
.C(n_170),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_SL g344 ( 
.A1(n_163),
.A2(n_170),
.B1(n_345),
.B2(n_346),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_163),
.Y(n_345)
);

XNOR2xp5_ASAP7_75t_L g445 ( 
.A(n_163),
.B(n_446),
.Y(n_445)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g343 ( 
.A(n_167),
.B(n_344),
.Y(n_343)
);

BUFx6f_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g233 ( 
.A(n_169),
.Y(n_233)
);

INVx13_ASAP7_75t_SL g346 ( 
.A(n_170),
.Y(n_346)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g437 ( 
.A(n_172),
.Y(n_437)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_173),
.A2(n_174),
.B1(n_176),
.B2(n_288),
.Y(n_287)
);

CKINVDCx16_ASAP7_75t_R g173 ( 
.A(n_174),
.Y(n_173)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_175),
.Y(n_408)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_176),
.Y(n_288)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

XNOR2x1_ASAP7_75t_SL g178 ( 
.A(n_179),
.B(n_180),
.Y(n_178)
);

MAJx2_ASAP7_75t_L g226 ( 
.A(n_179),
.B(n_181),
.C(n_184),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_181),
.A2(n_182),
.B1(n_183),
.B2(n_184),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g418 ( 
.A1(n_181),
.A2(n_182),
.B1(n_366),
.B2(n_367),
.Y(n_418)
);

INVx2_ASAP7_75t_SL g181 ( 
.A(n_182),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g362 ( 
.A(n_182),
.B(n_363),
.C(n_366),
.Y(n_362)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

INVx3_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

INVx6_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_189),
.A2(n_235),
.B1(n_254),
.B2(n_255),
.Y(n_188)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_189),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_SL g189 ( 
.A(n_190),
.B(n_225),
.Y(n_189)
);

HB1xp67_ASAP7_75t_L g295 ( 
.A(n_190),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_200),
.C(n_213),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_191),
.B(n_200),
.Y(n_262)
);

XNOR2x1_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_194),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_192),
.B(n_195),
.C(n_196),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_SL g194 ( 
.A(n_195),
.B(n_196),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_195),
.B(n_239),
.Y(n_238)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

INVx2_ASAP7_75t_L g450 ( 
.A(n_198),
.Y(n_450)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_199),
.Y(n_413)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_204),
.C(n_208),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_201),
.A2(n_208),
.B1(n_209),
.B2(n_291),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_201),
.Y(n_291)
);

BUFx6f_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_204),
.B(n_290),
.Y(n_289)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

INVx4_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

INVx4_ASAP7_75t_L g469 ( 
.A(n_207),
.Y(n_469)
);

MAJIxp5_ASAP7_75t_L g382 ( 
.A(n_208),
.B(n_383),
.C(n_387),
.Y(n_382)
);

AOI22xp5_ASAP7_75t_L g440 ( 
.A1(n_208),
.A2(n_209),
.B1(n_387),
.B2(n_441),
.Y(n_440)
);

INVx1_ASAP7_75t_SL g208 ( 
.A(n_209),
.Y(n_208)
);

INVx4_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

BUFx3_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_213),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_217),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_214),
.B(n_218),
.C(n_222),
.Y(n_234)
);

BUFx6f_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_222),
.Y(n_217)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

INVx3_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_227),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_226),
.B(n_295),
.C(n_296),
.Y(n_294)
);

HB1xp67_ASAP7_75t_L g296 ( 
.A(n_227),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_234),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_229),
.A2(n_230),
.B1(n_231),
.B2(n_232),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_229),
.B(n_232),
.C(n_234),
.Y(n_305)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_235),
.Y(n_255)
);

HB1xp67_ASAP7_75t_L g332 ( 
.A(n_235),
.Y(n_332)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_242),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_236),
.B(n_243),
.C(n_244),
.Y(n_306)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

INVx1_ASAP7_75t_SL g311 ( 
.A(n_239),
.Y(n_311)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

INVx3_ASAP7_75t_L g276 ( 
.A(n_241),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_243),
.B(n_244),
.Y(n_242)
);

XNOR2x1_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_247),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_245),
.B(n_248),
.C(n_249),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_249),
.Y(n_247)
);

INVx3_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_254),
.B(n_331),
.C(n_332),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_257),
.B(n_261),
.C(n_264),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g337 ( 
.A(n_258),
.B(n_261),
.Y(n_337)
);

XOR2x2_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_263),
.Y(n_261)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g336 ( 
.A(n_265),
.B(n_337),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_266),
.B(n_286),
.C(n_289),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g340 ( 
.A(n_266),
.B(n_341),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_267),
.B(n_271),
.C(n_279),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g392 ( 
.A(n_268),
.B(n_393),
.Y(n_392)
);

XNOR2xp5_ASAP7_75t_L g393 ( 
.A(n_271),
.B(n_279),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_277),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g391 ( 
.A(n_272),
.B(n_277),
.Y(n_391)
);

NOR2x1_ASAP7_75t_R g272 ( 
.A(n_273),
.B(n_274),
.Y(n_272)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

INVx2_ASAP7_75t_L g494 ( 
.A(n_276),
.Y(n_494)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_280),
.B(n_283),
.C(n_284),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_SL g378 ( 
.A1(n_280),
.A2(n_283),
.B1(n_379),
.B2(n_380),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_280),
.Y(n_379)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_283),
.Y(n_380)
);

MAJIxp5_ASAP7_75t_L g463 ( 
.A(n_283),
.B(n_464),
.C(n_466),
.Y(n_463)
);

OAI22xp5_ASAP7_75t_SL g479 ( 
.A1(n_283),
.A2(n_380),
.B1(n_466),
.B2(n_467),
.Y(n_479)
);

XOR2xp5_ASAP7_75t_L g377 ( 
.A(n_284),
.B(n_378),
.Y(n_377)
);

XNOR2xp5_ASAP7_75t_L g341 ( 
.A(n_286),
.B(n_289),
.Y(n_341)
);

OAI21xp5_ASAP7_75t_L g502 ( 
.A1(n_292),
.A2(n_503),
.B(n_504),
.Y(n_502)
);

AND2x2_ASAP7_75t_SL g292 ( 
.A(n_293),
.B(n_330),
.Y(n_292)
);

OR2x2_ASAP7_75t_L g504 ( 
.A(n_293),
.B(n_330),
.Y(n_504)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_294),
.B(n_297),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g540 ( 
.A(n_294),
.B(n_298),
.C(n_307),
.Y(n_540)
);

XNOR2x1_ASAP7_75t_L g297 ( 
.A(n_298),
.B(n_307),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_299),
.B(n_306),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_300),
.B(n_305),
.Y(n_299)
);

HB1xp67_ASAP7_75t_L g538 ( 
.A(n_300),
.Y(n_538)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_301),
.A2(n_302),
.B1(n_303),
.B2(n_304),
.Y(n_300)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_301),
.Y(n_303)
);

INVx1_ASAP7_75t_SL g304 ( 
.A(n_302),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g536 ( 
.A(n_305),
.B(n_537),
.C(n_538),
.Y(n_536)
);

INVxp67_ASAP7_75t_L g537 ( 
.A(n_306),
.Y(n_537)
);

XNOR2xp5_ASAP7_75t_L g307 ( 
.A(n_308),
.B(n_318),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g510 ( 
.A(n_308),
.B(n_319),
.C(n_320),
.Y(n_510)
);

XOR2xp5_ASAP7_75t_L g308 ( 
.A(n_309),
.B(n_312),
.Y(n_308)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

INVx3_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_L g318 ( 
.A(n_319),
.B(n_320),
.Y(n_318)
);

XOR2xp5_ASAP7_75t_L g320 ( 
.A(n_321),
.B(n_324),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g518 ( 
.A(n_321),
.B(n_325),
.C(n_519),
.Y(n_518)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

INVx3_ASAP7_75t_L g368 ( 
.A(n_323),
.Y(n_368)
);

XNOR2xp5_ASAP7_75t_L g324 ( 
.A(n_325),
.B(n_329),
.Y(n_324)
);

BUFx6f_ASAP7_75t_L g326 ( 
.A(n_327),
.Y(n_326)
);

INVx2_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

HB1xp67_ASAP7_75t_L g519 ( 
.A(n_329),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_334),
.B(n_396),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_335),
.B(n_338),
.C(n_372),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_336),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_336),
.B(n_339),
.Y(n_501)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_339),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_340),
.B(n_342),
.C(n_369),
.Y(n_339)
);

XOR2xp5_ASAP7_75t_L g394 ( 
.A(n_340),
.B(n_395),
.Y(n_394)
);

XNOR2xp5_ASAP7_75t_L g395 ( 
.A(n_342),
.B(n_369),
.Y(n_395)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_343),
.B(n_347),
.C(n_362),
.Y(n_342)
);

XNOR2xp5_ASAP7_75t_L g375 ( 
.A(n_343),
.B(n_347),
.Y(n_375)
);

MAJIxp5_ASAP7_75t_L g430 ( 
.A(n_345),
.B(n_431),
.C(n_435),
.Y(n_430)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_350),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_351),
.Y(n_350)
);

INVx2_ASAP7_75t_L g351 ( 
.A(n_352),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_353),
.Y(n_352)
);

INVx2_ASAP7_75t_L g353 ( 
.A(n_354),
.Y(n_353)
);

INVx3_ASAP7_75t_L g354 ( 
.A(n_355),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_L g356 ( 
.A(n_357),
.B(n_358),
.Y(n_356)
);

INVx2_ASAP7_75t_L g358 ( 
.A(n_359),
.Y(n_358)
);

BUFx6f_ASAP7_75t_L g359 ( 
.A(n_360),
.Y(n_359)
);

BUFx6f_ASAP7_75t_L g360 ( 
.A(n_361),
.Y(n_360)
);

XOR2xp5_ASAP7_75t_L g374 ( 
.A(n_362),
.B(n_375),
.Y(n_374)
);

XNOR2xp5_ASAP7_75t_SL g417 ( 
.A(n_363),
.B(n_418),
.Y(n_417)
);

AND2x2_ASAP7_75t_L g363 ( 
.A(n_364),
.B(n_365),
.Y(n_363)
);

XNOR2xp5_ASAP7_75t_L g405 ( 
.A(n_364),
.B(n_365),
.Y(n_405)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_364),
.Y(n_473)
);

AOI22xp5_ASAP7_75t_L g488 ( 
.A1(n_364),
.A2(n_473),
.B1(n_474),
.B2(n_489),
.Y(n_488)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_367),
.Y(n_366)
);

NOR2xp67_ASAP7_75t_L g372 ( 
.A(n_373),
.B(n_394),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_373),
.B(n_394),
.Y(n_397)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_374),
.B(n_376),
.C(n_392),
.Y(n_373)
);

XNOR2xp5_ASAP7_75t_L g419 ( 
.A(n_374),
.B(n_420),
.Y(n_419)
);

XNOR2xp5_ASAP7_75t_L g420 ( 
.A(n_376),
.B(n_392),
.Y(n_420)
);

MAJIxp5_ASAP7_75t_L g376 ( 
.A(n_377),
.B(n_381),
.C(n_390),
.Y(n_376)
);

XOR2xp5_ASAP7_75t_L g402 ( 
.A(n_377),
.B(n_403),
.Y(n_402)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_382),
.Y(n_381)
);

XNOR2xp5_ASAP7_75t_L g403 ( 
.A(n_382),
.B(n_391),
.Y(n_403)
);

XOR2x2_ASAP7_75t_L g439 ( 
.A(n_383),
.B(n_440),
.Y(n_439)
);

INVx2_ASAP7_75t_L g384 ( 
.A(n_385),
.Y(n_384)
);

INVx2_ASAP7_75t_L g385 ( 
.A(n_386),
.Y(n_385)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_387),
.Y(n_441)
);

INVx4_ASAP7_75t_L g388 ( 
.A(n_389),
.Y(n_388)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_391),
.Y(n_390)
);

NAND3xp33_ASAP7_75t_L g396 ( 
.A(n_397),
.B(n_398),
.C(n_501),
.Y(n_396)
);

OAI21xp5_ASAP7_75t_SL g398 ( 
.A1(n_399),
.A2(n_421),
.B(n_500),
.Y(n_398)
);

NOR2xp67_ASAP7_75t_L g399 ( 
.A(n_400),
.B(n_419),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_400),
.B(n_419),
.Y(n_500)
);

MAJIxp5_ASAP7_75t_L g400 ( 
.A(n_401),
.B(n_404),
.C(n_416),
.Y(n_400)
);

AOI22xp5_ASAP7_75t_L g423 ( 
.A1(n_401),
.A2(n_402),
.B1(n_424),
.B2(n_425),
.Y(n_423)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_402),
.Y(n_401)
);

AOI22xp5_ASAP7_75t_L g425 ( 
.A1(n_404),
.A2(n_416),
.B1(n_417),
.B2(n_426),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_404),
.Y(n_426)
);

MAJx2_ASAP7_75t_L g404 ( 
.A(n_405),
.B(n_406),
.C(n_409),
.Y(n_404)
);

XNOR2xp5_ASAP7_75t_L g429 ( 
.A(n_405),
.B(n_406),
.Y(n_429)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_408),
.Y(n_407)
);

XOR2xp5_ASAP7_75t_L g428 ( 
.A(n_409),
.B(n_429),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_410),
.B(n_414),
.Y(n_409)
);

AO22x1_ASAP7_75t_SL g454 ( 
.A1(n_410),
.A2(n_411),
.B1(n_414),
.B2(n_455),
.Y(n_454)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_411),
.Y(n_410)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_413),
.Y(n_412)
);

INVx1_ASAP7_75t_SL g455 ( 
.A(n_414),
.Y(n_455)
);

INVx2_ASAP7_75t_L g453 ( 
.A(n_415),
.Y(n_453)
);

INVx3_ASAP7_75t_L g476 ( 
.A(n_415),
.Y(n_476)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_417),
.Y(n_416)
);

AOI21xp5_ASAP7_75t_L g421 ( 
.A1(n_422),
.A2(n_442),
.B(n_499),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_SL g422 ( 
.A(n_423),
.B(n_427),
.Y(n_422)
);

NOR2xp67_ASAP7_75t_SL g499 ( 
.A(n_423),
.B(n_427),
.Y(n_499)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_425),
.Y(n_424)
);

MAJIxp5_ASAP7_75t_L g427 ( 
.A(n_428),
.B(n_430),
.C(n_438),
.Y(n_427)
);

XOR2xp5_ASAP7_75t_L g456 ( 
.A(n_428),
.B(n_457),
.Y(n_456)
);

XNOR2xp5_ASAP7_75t_L g457 ( 
.A(n_430),
.B(n_439),
.Y(n_457)
);

XNOR2xp5_ASAP7_75t_L g446 ( 
.A(n_431),
.B(n_435),
.Y(n_446)
);

INVx8_ASAP7_75t_L g432 ( 
.A(n_433),
.Y(n_432)
);

INVx6_ASAP7_75t_L g433 ( 
.A(n_434),
.Y(n_433)
);

INVx8_ASAP7_75t_L g436 ( 
.A(n_437),
.Y(n_436)
);

HB1xp67_ASAP7_75t_L g438 ( 
.A(n_439),
.Y(n_438)
);

OAI21x1_ASAP7_75t_SL g442 ( 
.A1(n_443),
.A2(n_458),
.B(n_498),
.Y(n_442)
);

AND2x2_ASAP7_75t_L g443 ( 
.A(n_444),
.B(n_456),
.Y(n_443)
);

OR2x2_ASAP7_75t_L g498 ( 
.A(n_444),
.B(n_456),
.Y(n_498)
);

MAJIxp5_ASAP7_75t_L g444 ( 
.A(n_445),
.B(n_447),
.C(n_454),
.Y(n_444)
);

XOR2xp5_ASAP7_75t_L g460 ( 
.A(n_445),
.B(n_461),
.Y(n_460)
);

AOI22xp5_ASAP7_75t_L g461 ( 
.A1(n_447),
.A2(n_448),
.B1(n_454),
.B2(n_462),
.Y(n_461)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_448),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_449),
.B(n_451),
.Y(n_448)
);

XNOR2xp5_ASAP7_75t_SL g465 ( 
.A(n_449),
.B(n_451),
.Y(n_465)
);

INVx2_ASAP7_75t_L g452 ( 
.A(n_453),
.Y(n_452)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_454),
.Y(n_462)
);

NOR2xp33_ASAP7_75t_L g490 ( 
.A(n_455),
.B(n_491),
.Y(n_490)
);

AOI21x1_ASAP7_75t_SL g458 ( 
.A1(n_459),
.A2(n_470),
.B(n_497),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_SL g459 ( 
.A(n_460),
.B(n_463),
.Y(n_459)
);

NOR2xp33_ASAP7_75t_L g497 ( 
.A(n_460),
.B(n_463),
.Y(n_497)
);

OAI22xp5_ASAP7_75t_SL g477 ( 
.A1(n_464),
.A2(n_465),
.B1(n_478),
.B2(n_479),
.Y(n_477)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_465),
.Y(n_464)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_467),
.Y(n_466)
);

INVx2_ASAP7_75t_L g468 ( 
.A(n_469),
.Y(n_468)
);

OAI21xp5_ASAP7_75t_SL g470 ( 
.A1(n_471),
.A2(n_480),
.B(n_496),
.Y(n_470)
);

NOR2xp33_ASAP7_75t_L g471 ( 
.A(n_472),
.B(n_477),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_472),
.B(n_477),
.Y(n_496)
);

NOR2xp33_ASAP7_75t_SL g472 ( 
.A(n_473),
.B(n_474),
.Y(n_472)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_474),
.Y(n_489)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_476),
.Y(n_475)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_479),
.Y(n_478)
);

AOI21xp5_ASAP7_75t_L g480 ( 
.A1(n_481),
.A2(n_490),
.B(n_495),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_482),
.B(n_488),
.Y(n_481)
);

NOR2xp33_ASAP7_75t_L g495 ( 
.A(n_482),
.B(n_488),
.Y(n_495)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_484),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_485),
.Y(n_484)
);

INVx3_ASAP7_75t_L g485 ( 
.A(n_486),
.Y(n_485)
);

INVx8_ASAP7_75t_L g486 ( 
.A(n_487),
.Y(n_486)
);

BUFx2_ASAP7_75t_L g492 ( 
.A(n_493),
.Y(n_492)
);

BUFx6f_ASAP7_75t_L g493 ( 
.A(n_494),
.Y(n_493)
);

NOR3xp33_ASAP7_75t_SL g505 ( 
.A(n_506),
.B(n_525),
.C(n_539),
.Y(n_505)
);

OAI21xp5_ASAP7_75t_SL g544 ( 
.A1(n_506),
.A2(n_545),
.B(n_548),
.Y(n_544)
);

NOR2xp67_ASAP7_75t_R g506 ( 
.A(n_507),
.B(n_523),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g548 ( 
.A(n_507),
.B(n_523),
.Y(n_548)
);

MAJIxp5_ASAP7_75t_L g507 ( 
.A(n_508),
.B(n_514),
.C(n_520),
.Y(n_507)
);

XNOR2xp5_ASAP7_75t_L g527 ( 
.A(n_508),
.B(n_528),
.Y(n_527)
);

MAJIxp5_ASAP7_75t_L g508 ( 
.A(n_509),
.B(n_511),
.C(n_513),
.Y(n_508)
);

INVxp67_ASAP7_75t_L g509 ( 
.A(n_510),
.Y(n_509)
);

XNOR2xp5_ASAP7_75t_L g532 ( 
.A(n_510),
.B(n_533),
.Y(n_532)
);

XNOR2xp5_ASAP7_75t_L g533 ( 
.A(n_511),
.B(n_513),
.Y(n_533)
);

AOI22xp5_ASAP7_75t_L g528 ( 
.A1(n_514),
.A2(n_520),
.B1(n_521),
.B2(n_529),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_514),
.Y(n_529)
);

MAJIxp5_ASAP7_75t_L g514 ( 
.A(n_515),
.B(n_517),
.C(n_518),
.Y(n_514)
);

XNOR2x1_ASAP7_75t_L g534 ( 
.A(n_515),
.B(n_535),
.Y(n_534)
);

XNOR2xp5_ASAP7_75t_L g535 ( 
.A(n_517),
.B(n_518),
.Y(n_535)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_521),
.Y(n_520)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_526),
.Y(n_525)
);

AOI21xp5_ASAP7_75t_L g545 ( 
.A1(n_526),
.A2(n_546),
.B(n_547),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_527),
.B(n_530),
.Y(n_526)
);

NOR2xp67_ASAP7_75t_SL g547 ( 
.A(n_527),
.B(n_530),
.Y(n_547)
);

MAJIxp5_ASAP7_75t_L g530 ( 
.A(n_531),
.B(n_534),
.C(n_536),
.Y(n_530)
);

AOI22xp5_ASAP7_75t_L g542 ( 
.A1(n_531),
.A2(n_532),
.B1(n_534),
.B2(n_543),
.Y(n_542)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_532),
.Y(n_531)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_534),
.Y(n_543)
);

XOR2xp5_ASAP7_75t_L g541 ( 
.A(n_536),
.B(n_542),
.Y(n_541)
);

AND2x2_ASAP7_75t_L g539 ( 
.A(n_540),
.B(n_541),
.Y(n_539)
);

NOR2xp33_ASAP7_75t_L g546 ( 
.A(n_540),
.B(n_541),
.Y(n_546)
);

NOR2xp33_ASAP7_75t_SL g550 ( 
.A(n_551),
.B(n_559),
.Y(n_550)
);

NOR2xp67_ASAP7_75t_R g551 ( 
.A(n_552),
.B(n_558),
.Y(n_551)
);

AND2x2_ASAP7_75t_L g559 ( 
.A(n_552),
.B(n_558),
.Y(n_559)
);

XNOR2xp5_ASAP7_75t_L g552 ( 
.A(n_553),
.B(n_554),
.Y(n_552)
);

CKINVDCx20_ASAP7_75t_R g557 ( 
.A(n_555),
.Y(n_557)
);


endmodule