module fake_jpeg_4272_n_69 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_69);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_69;

wire n_61;
wire n_45;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_59;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_65;
wire n_34;
wire n_39;
wire n_42;
wire n_49;
wire n_38;
wire n_56;
wire n_50;
wire n_67;
wire n_57;
wire n_53;
wire n_54;
wire n_40;
wire n_48;
wire n_35;
wire n_46;
wire n_44;
wire n_36;
wire n_62;
wire n_37;
wire n_43;
wire n_66;

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_30),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_25),
.Y(n_35)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_19),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

CKINVDCx5p33_ASAP7_75t_R g38 ( 
.A(n_24),
.Y(n_38)
);

BUFx16f_ASAP7_75t_L g39 ( 
.A(n_16),
.Y(n_39)
);

INVx11_ASAP7_75t_SL g40 ( 
.A(n_10),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_17),
.Y(n_41)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_2),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_4),
.B(n_20),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_31),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_21),
.B(n_13),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_40),
.Y(n_46)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_46),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_45),
.B(n_0),
.Y(n_47)
);

AND2x2_ASAP7_75t_L g53 ( 
.A(n_47),
.B(n_48),
.Y(n_53)
);

AND2x4_ASAP7_75t_L g48 ( 
.A(n_39),
.B(n_0),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_39),
.Y(n_49)
);

OAI22x1_ASAP7_75t_L g56 ( 
.A1(n_49),
.A2(n_38),
.B1(n_15),
.B2(n_5),
.Y(n_56)
);

BUFx4f_ASAP7_75t_SL g50 ( 
.A(n_36),
.Y(n_50)
);

AOI21xp5_ASAP7_75t_L g54 ( 
.A1(n_50),
.A2(n_41),
.B(n_35),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g51 ( 
.A1(n_48),
.A2(n_42),
.B1(n_44),
.B2(n_37),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_51),
.A2(n_55),
.B1(n_1),
.B2(n_54),
.Y(n_60)
);

INVxp67_ASAP7_75t_L g59 ( 
.A(n_54),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_L g55 ( 
.A1(n_48),
.A2(n_34),
.B1(n_2),
.B2(n_3),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_56),
.A2(n_43),
.B1(n_3),
.B2(n_1),
.Y(n_57)
);

OAI21xp5_ASAP7_75t_SL g61 ( 
.A1(n_57),
.A2(n_58),
.B(n_6),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_53),
.B(n_43),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_60),
.B(n_7),
.Y(n_62)
);

NAND3xp33_ASAP7_75t_L g63 ( 
.A(n_61),
.B(n_62),
.C(n_8),
.Y(n_63)
);

MAJIxp5_ASAP7_75t_L g64 ( 
.A(n_63),
.B(n_52),
.C(n_11),
.Y(n_64)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_64),
.B(n_9),
.C(n_12),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_65),
.B(n_14),
.Y(n_66)
);

OAI21xp5_ASAP7_75t_L g67 ( 
.A1(n_66),
.A2(n_59),
.B(n_22),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_67),
.B(n_18),
.Y(n_68)
);

AOI322xp5_ASAP7_75t_L g69 ( 
.A1(n_68),
.A2(n_23),
.A3(n_26),
.B1(n_27),
.B2(n_28),
.C1(n_32),
.C2(n_33),
.Y(n_69)
);


endmodule