module real_aes_15475_n_375 (n_76, n_113, n_187, n_90, n_257, n_65, n_74, n_185, n_285, n_30, n_222, n_61, n_20, n_287, n_357, n_64, n_254, n_207, n_10, n_83, n_181, n_362, n_124, n_191, n_209, n_299, n_322, n_328, n_19, n_40, n_318, n_355, n_239, n_100, n_54, n_112, n_319, n_364, n_35, n_42, n_329, n_132, n_131, n_144, n_169, n_242, n_308, n_172, n_341, n_232, n_6, n_69, n_317, n_353, n_321, n_73, n_320, n_77, n_260, n_37, n_97, n_186, n_138, n_374, n_26, n_235, n_245, n_161, n_189, n_271, n_2, n_145, n_227, n_92, n_330, n_332, n_292, n_116, n_94, n_289, n_280, n_333, n_213, n_356, n_184, n_28, n_372, n_202, n_56, n_370, n_34, n_98, n_121, n_352, n_125, n_216, n_82, n_327, n_47, n_106, n_32, n_263, n_230, n_51, n_248, n_301, n_27, n_343, n_369, n_174, n_18, n_104, n_211, n_281, n_173, n_234, n_284, n_153, n_316, n_75, n_178, n_298, n_49, n_43, n_297, n_9, n_119, n_310, n_164, n_231, n_44, n_102, n_122, n_141, n_128, n_111, n_167, n_80, n_179, n_12, n_68, n_129, n_345, n_304, n_311, n_324, n_25, n_278, n_236, n_367, n_267, n_218, n_48, n_204, n_339, n_89, n_277, n_331, n_93, n_182, n_363, n_323, n_199, n_350, n_142, n_223, n_67, n_368, n_250, n_85, n_45, n_5, n_244, n_118, n_139, n_87, n_171, n_78, n_146, n_17, n_226, n_255, n_286, n_120, n_261, n_238, n_360, n_58, n_165, n_361, n_246, n_176, n_163, n_29, n_52, n_251, n_220, n_197, n_296, n_3, n_41, n_256, n_71, n_302, n_351, n_126, n_200, n_115, n_96, n_110, n_150, n_147, n_288, n_23, n_334, n_274, n_160, n_303, n_95, n_188, n_269, n_201, n_306, n_158, n_4, n_366, n_346, n_193, n_293, n_162, n_358, n_275, n_214, n_46, n_109, n_59, n_203, n_81, n_133, n_273, n_114, n_276, n_295, n_265, n_354, n_154, n_127, n_326, n_24, n_217, n_55, n_62, n_291, n_148, n_88, n_159, n_11, n_108, n_373, n_60, n_233, n_290, n_365, n_155, n_243, n_268, n_136, n_157, n_282, n_101, n_309, n_344, n_229, n_107, n_33, n_53, n_36, n_149, n_190, n_262, n_134, n_349, n_336, n_195, n_300, n_252, n_283, n_314, n_249, n_221, n_156, n_359, n_57, n_66, n_21, n_31, n_8, n_312, n_183, n_266, n_205, n_335, n_177, n_313, n_22, n_140, n_219, n_180, n_212, n_210, n_325, n_338, n_371, n_103, n_166, n_224, n_151, n_130, n_253, n_99, n_15, n_72, n_152, n_198, n_7, n_228, n_272, n_196, n_347, n_315, n_123, n_279, n_79, n_270, n_305, n_117, n_208, n_215, n_135, n_70, n_50, n_170, n_86, n_340, n_13, n_168, n_175, n_241, n_105, n_84, n_294, n_258, n_206, n_307, n_342, n_348, n_14, n_194, n_137, n_225, n_16, n_39, n_337, n_247, n_240, n_38, n_259, n_143, n_192, n_0, n_264, n_63, n_1, n_237, n_91, n_375);
input n_76;
input n_113;
input n_187;
input n_90;
input n_257;
input n_65;
input n_74;
input n_185;
input n_285;
input n_30;
input n_222;
input n_61;
input n_20;
input n_287;
input n_357;
input n_64;
input n_254;
input n_207;
input n_10;
input n_83;
input n_181;
input n_362;
input n_124;
input n_191;
input n_209;
input n_299;
input n_322;
input n_328;
input n_19;
input n_40;
input n_318;
input n_355;
input n_239;
input n_100;
input n_54;
input n_112;
input n_319;
input n_364;
input n_35;
input n_42;
input n_329;
input n_132;
input n_131;
input n_144;
input n_169;
input n_242;
input n_308;
input n_172;
input n_341;
input n_232;
input n_6;
input n_69;
input n_317;
input n_353;
input n_321;
input n_73;
input n_320;
input n_77;
input n_260;
input n_37;
input n_97;
input n_186;
input n_138;
input n_374;
input n_26;
input n_235;
input n_245;
input n_161;
input n_189;
input n_271;
input n_2;
input n_145;
input n_227;
input n_92;
input n_330;
input n_332;
input n_292;
input n_116;
input n_94;
input n_289;
input n_280;
input n_333;
input n_213;
input n_356;
input n_184;
input n_28;
input n_372;
input n_202;
input n_56;
input n_370;
input n_34;
input n_98;
input n_121;
input n_352;
input n_125;
input n_216;
input n_82;
input n_327;
input n_47;
input n_106;
input n_32;
input n_263;
input n_230;
input n_51;
input n_248;
input n_301;
input n_27;
input n_343;
input n_369;
input n_174;
input n_18;
input n_104;
input n_211;
input n_281;
input n_173;
input n_234;
input n_284;
input n_153;
input n_316;
input n_75;
input n_178;
input n_298;
input n_49;
input n_43;
input n_297;
input n_9;
input n_119;
input n_310;
input n_164;
input n_231;
input n_44;
input n_102;
input n_122;
input n_141;
input n_128;
input n_111;
input n_167;
input n_80;
input n_179;
input n_12;
input n_68;
input n_129;
input n_345;
input n_304;
input n_311;
input n_324;
input n_25;
input n_278;
input n_236;
input n_367;
input n_267;
input n_218;
input n_48;
input n_204;
input n_339;
input n_89;
input n_277;
input n_331;
input n_93;
input n_182;
input n_363;
input n_323;
input n_199;
input n_350;
input n_142;
input n_223;
input n_67;
input n_368;
input n_250;
input n_85;
input n_45;
input n_5;
input n_244;
input n_118;
input n_139;
input n_87;
input n_171;
input n_78;
input n_146;
input n_17;
input n_226;
input n_255;
input n_286;
input n_120;
input n_261;
input n_238;
input n_360;
input n_58;
input n_165;
input n_361;
input n_246;
input n_176;
input n_163;
input n_29;
input n_52;
input n_251;
input n_220;
input n_197;
input n_296;
input n_3;
input n_41;
input n_256;
input n_71;
input n_302;
input n_351;
input n_126;
input n_200;
input n_115;
input n_96;
input n_110;
input n_150;
input n_147;
input n_288;
input n_23;
input n_334;
input n_274;
input n_160;
input n_303;
input n_95;
input n_188;
input n_269;
input n_201;
input n_306;
input n_158;
input n_4;
input n_366;
input n_346;
input n_193;
input n_293;
input n_162;
input n_358;
input n_275;
input n_214;
input n_46;
input n_109;
input n_59;
input n_203;
input n_81;
input n_133;
input n_273;
input n_114;
input n_276;
input n_295;
input n_265;
input n_354;
input n_154;
input n_127;
input n_326;
input n_24;
input n_217;
input n_55;
input n_62;
input n_291;
input n_148;
input n_88;
input n_159;
input n_11;
input n_108;
input n_373;
input n_60;
input n_233;
input n_290;
input n_365;
input n_155;
input n_243;
input n_268;
input n_136;
input n_157;
input n_282;
input n_101;
input n_309;
input n_344;
input n_229;
input n_107;
input n_33;
input n_53;
input n_36;
input n_149;
input n_190;
input n_262;
input n_134;
input n_349;
input n_336;
input n_195;
input n_300;
input n_252;
input n_283;
input n_314;
input n_249;
input n_221;
input n_156;
input n_359;
input n_57;
input n_66;
input n_21;
input n_31;
input n_8;
input n_312;
input n_183;
input n_266;
input n_205;
input n_335;
input n_177;
input n_313;
input n_22;
input n_140;
input n_219;
input n_180;
input n_212;
input n_210;
input n_325;
input n_338;
input n_371;
input n_103;
input n_166;
input n_224;
input n_151;
input n_130;
input n_253;
input n_99;
input n_15;
input n_72;
input n_152;
input n_198;
input n_7;
input n_228;
input n_272;
input n_196;
input n_347;
input n_315;
input n_123;
input n_279;
input n_79;
input n_270;
input n_305;
input n_117;
input n_208;
input n_215;
input n_135;
input n_70;
input n_50;
input n_170;
input n_86;
input n_340;
input n_13;
input n_168;
input n_175;
input n_241;
input n_105;
input n_84;
input n_294;
input n_258;
input n_206;
input n_307;
input n_342;
input n_348;
input n_14;
input n_194;
input n_137;
input n_225;
input n_16;
input n_39;
input n_337;
input n_247;
input n_240;
input n_38;
input n_259;
input n_143;
input n_192;
input n_0;
input n_264;
input n_63;
input n_1;
input n_237;
input n_91;
output n_375;
wire n_476;
wire n_599;
wire n_887;
wire n_1314;
wire n_1279;
wire n_830;
wire n_1371;
wire n_624;
wire n_618;
wire n_1797;
wire n_933;
wire n_485;
wire n_822;
wire n_750;
wire n_1641;
wire n_503;
wire n_1781;
wire n_1762;
wire n_1591;
wire n_469;
wire n_1310;
wire n_1376;
wire n_592;
wire n_1621;
wire n_1729;
wire n_1737;
wire n_761;
wire n_421;
wire n_919;
wire n_1888;
wire n_1217;
wire n_1423;
wire n_571;
wire n_549;
wire n_1328;
wire n_1034;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_593;
wire n_989;
wire n_431;
wire n_1044;
wire n_1730;
wire n_1744;
wire n_963;
wire n_551;
wire n_884;
wire n_814;
wire n_944;
wire n_1283;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_1873;
wire n_1313;
wire n_1835;
wire n_1871;
wire n_1468;
wire n_1713;
wire n_870;
wire n_1248;
wire n_1602;
wire n_548;
wire n_1859;
wire n_572;
wire n_815;
wire n_1140;
wire n_1453;
wire n_1520;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_1379;
wire n_400;
wire n_1845;
wire n_1597;
wire n_1415;
wire n_1160;
wire n_1849;
wire n_1287;
wire n_883;
wire n_478;
wire n_1575;
wire n_1687;
wire n_553;
wire n_1805;
wire n_744;
wire n_1367;
wire n_1325;
wire n_1225;
wire n_1382;
wire n_875;
wire n_1199;
wire n_951;
wire n_1441;
wire n_1543;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_1833;
wire n_1477;
wire n_595;
wire n_1893;
wire n_1282;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_962;
wire n_1599;
wire n_755;
wire n_409;
wire n_781;
wire n_576;
wire n_1688;
wire n_956;
wire n_1242;
wire n_1537;
wire n_796;
wire n_874;
wire n_1126;
wire n_383;
wire n_1607;
wire n_455;
wire n_1771;
wire n_1809;
wire n_682;
wire n_1745;
wire n_1820;
wire n_812;
wire n_782;
wire n_817;
wire n_1883;
wire n_608;
wire n_760;
wire n_534;
wire n_1454;
wire n_708;
wire n_1020;
wire n_885;
wire n_950;
wire n_381;
wire n_1196;
wire n_1013;
wire n_808;
wire n_1639;
wire n_1224;
wire n_1872;
wire n_1694;
wire n_688;
wire n_1042;
wire n_1588;
wire n_1317;
wire n_417;
wire n_690;
wire n_1419;
wire n_499;
wire n_1142;
wire n_1731;
wire n_1589;
wire n_947;
wire n_970;
wire n_1677;
wire n_1149;
wire n_527;
wire n_1676;
wire n_1342;
wire n_1440;
wire n_1346;
wire n_552;
wire n_1383;
wire n_1890;
wire n_1675;
wire n_590;
wire n_1293;
wire n_1880;
wire n_432;
wire n_1882;
wire n_1131;
wire n_1008;
wire n_1491;
wire n_1865;
wire n_805;
wire n_1600;
wire n_619;
wire n_1250;
wire n_1095;
wire n_1583;
wire n_1284;
wire n_1465;
wire n_859;
wire n_1486;
wire n_1304;
wire n_685;
wire n_1080;
wire n_917;
wire n_1247;
wire n_488;
wire n_501;
wire n_1380;
wire n_1658;
wire n_1866;
wire n_954;
wire n_702;
wire n_1874;
wire n_1007;
wire n_898;
wire n_562;
wire n_1022;
wire n_1502;
wire n_1073;
wire n_404;
wire n_728;
wire n_1301;
wire n_1632;
wire n_1201;
wire n_997;
wire n_1105;
wire n_1768;
wire n_1243;
wire n_1846;
wire n_1003;
wire n_749;
wire n_1870;
wire n_914;
wire n_1837;
wire n_1286;
wire n_494;
wire n_1661;
wire n_927;
wire n_723;
wire n_1351;
wire n_972;
wire n_1813;
wire n_1628;
wire n_1587;
wire n_1821;
wire n_1570;
wire n_1209;
wire n_411;
wire n_498;
wire n_765;
wire n_1397;
wire n_1554;
wire n_648;
wire n_1487;
wire n_939;
wire n_1825;
wire n_1615;
wire n_1763;
wire n_928;
wire n_1384;
wire n_789;
wire n_1515;
wire n_738;
wire n_1387;
wire n_922;
wire n_1048;
wire n_1422;
wire n_787;
wire n_1214;
wire n_806;
wire n_715;
wire n_1714;
wire n_420;
wire n_1666;
wire n_1490;
wire n_1258;
wire n_873;
wire n_438;
wire n_1814;
wire n_446;
wire n_1281;
wire n_1559;
wire n_1495;
wire n_1510;
wire n_1727;
wire n_712;
wire n_422;
wire n_861;
wire n_1574;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_1742;
wire n_724;
wire n_1648;
wire n_440;
wire n_1231;
wire n_1305;
wire n_1161;
wire n_686;
wire n_1299;
wire n_949;
wire n_586;
wire n_1508;
wire n_1421;
wire n_788;
wire n_441;
wire n_1045;
wire n_1339;
wire n_1793;
wire n_837;
wire n_1349;
wire n_1708;
wire n_1445;
wire n_1631;
wire n_829;
wire n_1030;
wire n_1348;
wire n_1391;
wire n_597;
wire n_1036;
wire n_687;
wire n_1751;
wire n_1765;
wire n_1538;
wire n_652;
wire n_500;
wire n_804;
wire n_1173;
wire n_854;
wire n_1787;
wire n_424;
wire n_877;
wire n_802;
wire n_1876;
wire n_1488;
wire n_1572;
wire n_1514;
wire n_480;
wire n_1652;
wire n_684;
wire n_1178;
wire n_1531;
wire n_821;
wire n_1657;
wire n_1616;
wire n_1828;
wire n_1860;
wire n_1563;
wire n_1018;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_1561;
wire n_635;
wire n_792;
wire n_1542;
wire n_1392;
wire n_665;
wire n_991;
wire n_667;
wire n_1712;
wire n_1556;
wire n_580;
wire n_1004;
wire n_1370;
wire n_1417;
wire n_1703;
wire n_1717;
wire n_1723;
wire n_979;
wire n_445;
wire n_596;
wire n_1740;
wire n_1197;
wire n_657;
wire n_1260;
wire n_1606;
wire n_1129;
wire n_1760;
wire n_1285;
wire n_1014;
wire n_742;
wire n_1385;
wire n_1629;
wire n_1618;
wire n_461;
wire n_1770;
wire n_1047;
wire n_1016;
wire n_1545;
wire n_694;
wire n_1350;
wire n_894;
wire n_1750;
wire n_1852;
wire n_545;
wire n_1459;
wire n_1530;
wire n_401;
wire n_538;
wire n_1830;
wire n_1594;
wire n_1864;
wire n_537;
wire n_1767;
wire n_1651;
wire n_560;
wire n_1094;
wire n_1776;
wire n_1719;
wire n_1220;
wire n_696;
wire n_1147;
wire n_1425;
wire n_1613;
wire n_1504;
wire n_704;
wire n_453;
wire n_647;
wire n_399;
wire n_948;
wire n_1499;
wire n_700;
wire n_1269;
wire n_677;
wire n_378;
wire n_591;
wire n_1635;
wire n_1518;
wire n_1702;
wire n_1366;
wire n_678;
wire n_415;
wire n_1400;
wire n_564;
wire n_638;
wire n_1361;
wire n_510;
wire n_1358;
wire n_1577;
wire n_1839;
wire n_1642;
wire n_1406;
wire n_550;
wire n_966;
wire n_1881;
wire n_1568;
wire n_1368;
wire n_994;
wire n_384;
wire n_1479;
wire n_1612;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_1611;
wire n_992;
wire n_813;
wire n_1338;
wire n_981;
wire n_1884;
wire n_1182;
wire n_872;
wire n_1401;
wire n_1086;
wire n_1070;
wire n_1189;
wire n_1665;
wire n_535;
wire n_882;
wire n_1210;
wire n_1741;
wire n_1456;
wire n_1879;
wire n_746;
wire n_656;
wire n_1614;
wire n_1148;
wire n_748;
wire n_860;
wire n_1261;
wire n_1062;
wire n_1439;
wire n_651;
wire n_1585;
wire n_1500;
wire n_801;
wire n_1271;
wire n_1653;
wire n_529;
wire n_504;
wire n_973;
wire n_1853;
wire n_1364;
wire n_659;
wire n_634;
wire n_903;
wire n_1668;
wire n_565;
wire n_925;
wire n_1389;
wire n_1393;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_1362;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_1553;
wire n_754;
wire n_508;
wire n_1141;
wire n_1769;
wire n_1812;
wire n_1112;
wire n_1485;
wire n_1408;
wire n_1680;
wire n_428;
wire n_783;
wire n_1107;
wire n_1564;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1516;
wire n_1386;
wire n_406;
wire n_1493;
wire n_1579;
wire n_1854;
wire n_617;
wire n_602;
wire n_402;
wire n_733;
wire n_1404;
wire n_1856;
wire n_658;
wire n_676;
wire n_531;
wire n_1848;
wire n_1031;
wire n_1394;
wire n_807;
wire n_1011;
wire n_416;
wire n_1567;
wire n_1569;
wire n_895;
wire n_799;
wire n_490;
wire n_391;
wire n_695;
wire n_1181;
wire n_881;
wire n_1626;
wire n_1145;
wire n_645;
wire n_1529;
wire n_557;
wire n_1681;
wire n_1620;
wire n_777;
wire n_985;
wire n_1659;
wire n_910;
wire n_642;
wire n_613;
wire n_1773;
wire n_1125;
wire n_1347;
wire n_1655;
wire n_1766;
wire n_1522;
wire n_1163;
wire n_1278;
wire n_734;
wire n_1623;
wire n_735;
wire n_1179;
wire n_569;
wire n_1171;
wire n_785;
wire n_1203;
wire n_1716;
wire n_1232;
wire n_471;
wire n_1857;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1580;
wire n_1000;
wire n_1187;
wire n_649;
wire n_1234;
wire n_622;
wire n_1634;
wire n_1002;
wire n_1353;
wire n_1165;
wire n_1551;
wire n_1667;
wire n_1058;
wire n_1216;
wire n_662;
wire n_1862;
wire n_850;
wire n_720;
wire n_1026;
wire n_1756;
wire n_1803;
wire n_492;
wire n_407;
wire n_419;
wire n_1023;
wire n_730;
wire n_1699;
wire n_1794;
wire n_1748;
wire n_643;
wire n_1403;
wire n_486;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_526;
wire n_1513;
wire n_1194;
wire n_389;
wire n_1609;
wire n_1462;
wire n_701;
wire n_809;
wire n_1532;
wire n_520;
wire n_679;
wire n_926;
wire n_1643;
wire n_942;
wire n_1374;
wire n_1120;
wire n_1497;
wire n_1548;
wire n_1784;
wire n_1526;
wire n_689;
wire n_1483;
wire n_946;
wire n_753;
wire n_1409;
wire n_1188;
wire n_623;
wire n_1474;
wire n_1032;
wire n_721;
wire n_1431;
wire n_1806;
wire n_1829;
wire n_1133;
wire n_1775;
wire n_1593;
wire n_739;
wire n_1322;
wire n_1525;
wire n_1732;
wire n_1162;
wire n_1463;
wire n_762;
wire n_1524;
wire n_1298;
wire n_442;
wire n_1633;
wire n_740;
wire n_1686;
wire n_1357;
wire n_639;
wire n_1186;
wire n_1365;
wire n_1807;
wire n_459;
wire n_1172;
wire n_998;
wire n_1689;
wire n_1625;
wire n_1395;
wire n_1276;
wire n_836;
wire n_1733;
wire n_1184;
wire n_583;
wire n_414;
wire n_1336;
wire n_776;
wire n_1138;
wire n_890;
wire n_1306;
wire n_1413;
wire n_1783;
wire n_1759;
wire n_1266;
wire n_497;
wire n_911;
wire n_450;
wire n_1578;
wire n_473;
wire n_1779;
wire n_967;
wire n_1709;
wire n_474;
wire n_1159;
wire n_1315;
wire n_1055;
wire n_611;
wire n_380;
wire n_1576;
wire n_844;
wire n_1840;
wire n_968;
wire n_710;
wire n_1040;
wire n_1185;
wire n_1102;
wire n_661;
wire n_447;
wire n_1795;
wire n_403;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1069;
wire n_1451;
wire n_842;
wire n_1788;
wire n_798;
wire n_1700;
wire n_668;
wire n_862;
wire n_869;
wire n_1816;
wire n_1811;
wire n_1066;
wire n_1377;
wire n_800;
wire n_778;
wire n_1170;
wire n_1175;
wire n_522;
wire n_1475;
wire n_943;
wire n_977;
wire n_905;
wire n_386;
wire n_878;
wire n_1734;
wire n_1333;
wire n_577;
wire n_1610;
wire n_759;
wire n_1235;
wire n_900;
wire n_841;
wire n_1724;
wire n_1218;
wire n_736;
wire n_1706;
wire n_766;
wire n_1113;
wire n_852;
wire n_1268;
wire n_1695;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_1302;
wire n_1289;
wire n_937;
wire n_1442;
wire n_773;
wire n_1446;
wire n_1778;
wire n_865;
wire n_1644;
wire n_1736;
wire n_1707;
wire n_594;
wire n_856;
wire n_1146;
wire n_1685;
wire n_1810;
wire n_1435;
wire n_1800;
wire n_932;
wire n_958;
wire n_1755;
wire n_775;
wire n_763;
wire n_1093;
wire n_427;
wire n_1540;
wire n_519;
wire n_1878;
wire n_1116;
wire n_709;
wire n_1834;
wire n_388;
wire n_1470;
wire n_816;
wire n_625;
wire n_953;
wire n_1565;
wire n_1373;
wire n_1558;
wire n_716;
wire n_1683;
wire n_584;
wire n_896;
wire n_1817;
wire n_1722;
wire n_528;
wire n_1078;
wire n_495;
wire n_1072;
wire n_1638;
wire n_1663;
wire n_935;
wire n_1505;
wire n_467;
wire n_1213;
wire n_1053;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_1168;
wire n_1598;
wire n_1309;
wire n_909;
wire n_523;
wire n_996;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1850;
wire n_1332;
wire n_1263;
wire n_1411;
wire n_1115;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_1726;
wire n_1827;
wire n_1656;
wire n_454;
wire n_1303;
wire n_1471;
wire n_443;
wire n_1029;
wire n_1207;
wire n_1555;
wire n_664;
wire n_1017;
wire n_936;
wire n_581;
wire n_1215;
wire n_582;
wire n_641;
wire n_1738;
wire n_940;
wire n_745;
wire n_1608;
wire n_1167;
wire n_1327;
wire n_609;
wire n_1743;
wire n_1752;
wire n_1792;
wire n_1006;
wire n_1869;
wire n_1259;
wire n_561;
wire n_437;
wire n_1560;
wire n_405;
wire n_1223;
wire n_621;
wire n_1012;
wire n_1241;
wire n_1414;
wire n_1671;
wire n_502;
wire n_434;
wire n_769;
wire n_1212;
wire n_1455;
wire n_1054;
wire n_1669;
wire n_1308;
wire n_1050;
wire n_426;
wire n_1550;
wire n_1134;
wire n_1895;
wire n_1670;
wire n_1319;
wire n_1363;
wire n_616;
wire n_880;
wire n_1103;
wire n_1274;
wire n_832;
wire n_1321;
wire n_1429;
wire n_1660;
wire n_1060;
wire n_1154;
wire n_1786;
wire n_632;
wire n_1344;
wire n_1450;
wire n_1603;
wire n_1720;
wire n_1331;
wire n_714;
wire n_1222;
wire n_1041;
wire n_1764;
wire n_1512;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_1335;
wire n_1405;
wire n_912;
wire n_464;
wire n_1227;
wire n_1509;
wire n_945;
wire n_392;
wire n_563;
wire n_891;
wire n_568;
wire n_1586;
wire n_413;
wire n_1157;
wire n_902;
wire n_1749;
wire n_1158;
wire n_1886;
wire n_1079;
wire n_1330;
wire n_1033;
wire n_1464;
wire n_1028;
wire n_1832;
wire n_727;
wire n_1083;
wire n_397;
wire n_1855;
wire n_1056;
wire n_1592;
wire n_1605;
wire n_1802;
wire n_663;
wire n_588;
wire n_1682;
wire n_1698;
wire n_1448;
wire n_707;
wire n_915;
wire n_1785;
wire n_1774;
wire n_1001;
wire n_1418;
wire n_711;
wire n_864;
wire n_1782;
wire n_1169;
wire n_377;
wire n_1139;
wire n_1482;
wire n_1798;
wire n_1038;
wire n_1085;
wire n_1838;
wire n_845;
wire n_1673;
wire n_1619;
wire n_1127;
wire n_1718;
wire n_484;
wire n_893;
wire n_1068;
wire n_747;
wire n_1672;
wire n_1753;
wire n_1244;
wire n_1581;
wire n_1863;
wire n_697;
wire n_978;
wire n_847;
wire n_1452;
wire n_826;
wire n_628;
wire n_487;
wire n_831;
wire n_1772;
wire n_653;
wire n_1725;
wire n_692;
wire n_1433;
wire n_1051;
wire n_1696;
wire n_1355;
wire n_1494;
wire n_1517;
wire n_827;
wire n_472;
wire n_866;
wire n_452;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_1426;
wire n_858;
wire n_764;
wire n_741;
wire n_1090;
wire n_456;
wire n_1469;
wire n_1164;
wire n_433;
wire n_627;
wire n_1693;
wire n_1791;
wire n_418;
wire n_771;
wire n_524;
wire n_1378;
wire n_1496;
wire n_705;
wire n_1191;
wire n_1206;
wire n_1824;
wire n_1270;
wire n_1566;
wire n_1399;
wire n_546;
wire n_1010;
wire n_1375;
wire n_1015;
wire n_1761;
wire n_863;
wire n_525;
wire n_1226;
wire n_1617;
wire n_1790;
wire n_644;
wire n_1150;
wire n_1861;
wire n_1341;
wire n_833;
wire n_1229;
wire n_1690;
wire n_929;
wire n_1143;
wire n_1190;
wire n_1728;
wire n_543;
wire n_1710;
wire n_585;
wire n_465;
wire n_719;
wire n_1343;
wire n_1457;
wire n_1604;
wire n_1156;
wire n_988;
wire n_1757;
wire n_1466;
wire n_921;
wire n_1396;
wire n_1799;
wire n_640;
wire n_1176;
wire n_1691;
wire n_1721;
wire n_1511;
wire n_1151;
wire n_1501;
wire n_1254;
wire n_1458;
wire n_646;
wire n_650;
wire n_1211;
wire n_743;
wire n_823;
wire n_393;
wire n_1804;
wire n_1480;
wire n_1101;
wire n_1076;
wire n_1251;
wire n_1434;
wire n_1461;
wire n_1449;
wire n_1715;
wire n_1407;
wire n_1104;
wire n_1061;
wire n_849;
wire n_554;
wire n_1153;
wire n_1337;
wire n_797;
wire n_1704;
wire n_1844;
wire n_1177;
wire n_758;
wire n_436;
wire n_390;
wire n_1096;
wire n_1316;
wire n_1590;
wire n_1420;
wire n_1552;
wire n_1544;
wire n_1571;
wire n_1092;
wire n_1841;
wire n_846;
wire n_631;
wire n_673;
wire n_1410;
wire n_1067;
wire n_518;
wire n_1192;
wire n_1292;
wire n_1478;
wire n_1507;
wire n_1240;
wire n_1789;
wire n_987;
wire n_1596;
wire n_1065;
wire n_540;
wire n_1064;
wire n_1075;
wire n_1822;
wire n_718;
wire n_669;
wire n_1091;
wire n_423;
wire n_1221;
wire n_458;
wire n_1200;
wire n_444;
wire n_1777;
wire n_555;
wire n_1295;
wire n_974;
wire n_1329;
wire n_857;
wire n_1424;
wire n_1819;
wire n_1887;
wire n_1674;
wire n_376;
wire n_491;
wire n_1294;
wire n_1110;
wire n_1137;
wire n_1533;
wire n_1889;
wire n_460;
wire n_1679;
wire n_1595;
wire n_1735;
wire n_666;
wire n_660;
wire n_1359;
wire n_886;
wire n_1896;
wire n_767;
wire n_889;
wire n_1398;
wire n_379;
wire n_1847;
wire n_1432;
wire n_1021;
wire n_1297;
wire n_1046;
wire n_1109;
wire n_961;
wire n_1447;
wire n_489;
wire n_1622;
wire n_1381;
wire n_1582;
wire n_1747;
wire n_573;
wire n_1099;
wire n_1654;
wire n_626;
wire n_539;
wire n_462;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_1541;
wire n_1272;
wire n_408;
wire n_1754;
wire n_578;
wire n_892;
wire n_938;
wire n_774;
wire n_466;
wire n_1584;
wire n_559;
wire n_1277;
wire n_1049;
wire n_984;
wire n_726;
wire n_517;
wire n_1851;
wire n_780;
wire n_931;
wire n_530;
wire n_834;
wire n_693;
wire n_496;
wire n_1257;
wire n_1360;
wire n_1082;
wire n_468;
wire n_532;
wire n_1025;
wire n_1875;
wire n_1826;
wire n_1836;
wire n_924;
wire n_1264;
wire n_1858;
wire n_1527;
wire n_1245;
wire n_1152;
wire n_1539;
wire n_1081;
wire n_547;
wire n_1324;
wire n_1198;
wire n_1678;
wire n_1307;
wire n_993;
wire n_819;
wire n_737;
wire n_1489;
wire n_1637;
wire n_1318;
wire n_1290;
wire n_1063;
wire n_1135;
wire n_828;
wire n_770;
wire n_867;
wire n_398;
wire n_1100;
wire n_1519;
wire n_425;
wire n_1650;
wire n_879;
wire n_1640;
wire n_449;
wire n_1340;
wire n_1562;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_1443;
wire n_1818;
wire n_655;
wire n_654;
wire n_1521;
wire n_672;
wire n_567;
wire n_916;
wire n_1354;
wire n_1780;
wire n_1547;
wire n_1823;
wire n_1867;
wire n_1334;
wire n_1291;
wire n_1437;
wire n_1473;
wire n_986;
wire n_451;
wire n_1891;
wire n_1037;
wire n_1267;
wire n_790;
wire n_1262;
wire n_1843;
wire n_410;
wire n_1684;
wire n_1444;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_1506;
wire n_1885;
wire n_1356;
wire n_1646;
wire n_768;
wire n_412;
wire n_542;
wire n_1256;
wire n_1427;
wire n_1077;
wire n_1111;
wire n_1503;
wire n_1249;
wire n_1416;
wire n_387;
wire n_1239;
wire n_1796;
wire n_1662;
wire n_969;
wire n_1535;
wire n_1009;
wire n_1202;
wire n_1498;
wire n_1801;
wire n_1549;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_430;
wire n_1252;
wire n_1647;
wire n_1132;
wire n_1649;
wire n_1275;
wire n_843;
wire n_579;
wire n_533;
wire n_1472;
wire n_385;
wire n_536;
wire n_470;
wire n_851;
wire n_1155;
wire n_934;
wire n_1636;
wire n_1027;
wire n_965;
wire n_1894;
wire n_1296;
wire n_382;
wire n_1484;
wire n_1043;
wire n_435;
wire n_511;
wire n_1808;
wire n_1492;
wire n_1467;
wire n_509;
wire n_1204;
wire n_930;
wire n_1265;
wire n_1057;
wire n_907;
wire n_1430;
wire n_1481;
wire n_1758;
wire n_1005;
wire n_1312;
wire n_1697;
wire n_1877;
wire n_899;
wire n_637;
wire n_544;
wire n_1476;
wire n_1087;
wire n_1842;
wire n_1536;
wire n_1746;
wire n_1711;
wire n_482;
wire n_633;
wire n_1892;
wire n_971;
wire n_1052;
wire n_1071;
wire n_1311;
wire n_1601;
wire n_1438;
wire n_1273;
wire n_959;
wire n_1573;
wire n_1130;
wire n_794;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1624;
wire n_1253;
wire n_1183;
wire n_1831;
wire n_516;
wire n_1460;
wire n_521;
wire n_1195;
wire n_1300;
wire n_575;
wire n_1372;
wire n_698;
wire n_1345;
wire n_587;
wire n_1701;
wire n_1664;
wire n_1428;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_1546;
wire n_1436;
wire n_793;
wire n_1390;
wire n_1815;
wire n_1868;
wire n_1412;
wire n_757;
wire n_1534;
wire n_803;
wire n_514;
wire n_507;
wire n_1557;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1739;
wire n_1088;
wire n_1230;
wire n_1326;
wire n_1402;
wire n_1388;
wire n_483;
wire n_1630;
wire n_394;
wire n_729;
wire n_1352;
wire n_1280;
wire n_1323;
wire n_1369;
wire n_703;
wire n_1097;
wire n_601;
wire n_463;
wire n_396;
wire n_1236;
wire n_1523;
wire n_1528;
wire n_603;
wire n_1692;
wire n_1288;
wire n_868;
wire n_1705;
wire n_1024;
wire n_1144;
wire n_1627;
wire n_475;
wire n_897;
wire n_1320;
wire n_855;
wire n_1645;
wire n_429;
AOI22xp33_ASAP7_75t_SL g582 ( .A1(n_0), .A2(n_335), .B1(n_463), .B2(n_583), .Y(n_582) );
INVxp67_ASAP7_75t_SL g633 ( .A(n_0), .Y(n_633) );
INVx1_ASAP7_75t_L g1817 ( .A(n_1), .Y(n_1817) );
INVx1_ASAP7_75t_L g842 ( .A(n_2), .Y(n_842) );
AO22x1_ASAP7_75t_L g881 ( .A1(n_2), .A2(n_247), .B1(n_515), .B2(n_770), .Y(n_881) );
INVx1_ASAP7_75t_L g391 ( .A(n_3), .Y(n_391) );
AND2x2_ASAP7_75t_L g444 ( .A(n_3), .B(n_272), .Y(n_444) );
AND2x2_ASAP7_75t_L g505 ( .A(n_3), .B(n_506), .Y(n_505) );
NOR2xp33_ASAP7_75t_L g879 ( .A(n_3), .B(n_401), .Y(n_879) );
INVx1_ASAP7_75t_L g854 ( .A(n_4), .Y(n_854) );
AOI22xp33_ASAP7_75t_L g880 ( .A1(n_4), .A2(n_147), .B1(n_520), .B2(n_766), .Y(n_880) );
AOI22xp33_ASAP7_75t_SL g1139 ( .A1(n_5), .A2(n_339), .B1(n_569), .B2(n_583), .Y(n_1139) );
AOI221xp5_ASAP7_75t_L g1154 ( .A1(n_5), .A2(n_6), .B1(n_524), .B2(n_542), .C(n_1155), .Y(n_1154) );
AOI22xp33_ASAP7_75t_SL g1146 ( .A1(n_6), .A2(n_9), .B1(n_465), .B2(n_956), .Y(n_1146) );
AOI22xp33_ASAP7_75t_SL g1093 ( .A1(n_7), .A2(n_334), .B1(n_583), .B2(n_986), .Y(n_1093) );
AOI221xp5_ASAP7_75t_L g1110 ( .A1(n_7), .A2(n_281), .B1(n_773), .B2(n_1111), .C(n_1113), .Y(n_1110) );
AOI22xp5_ASAP7_75t_L g1629 ( .A1(n_8), .A2(n_63), .B1(n_1580), .B2(n_1584), .Y(n_1629) );
A2O1A1Ixp33_ASAP7_75t_L g1160 ( .A1(n_9), .A2(n_1026), .B(n_1161), .C(n_1165), .Y(n_1160) );
OAI22xp5_ASAP7_75t_L g1263 ( .A1(n_10), .A2(n_234), .B1(n_412), .B2(n_1214), .Y(n_1263) );
INVx1_ASAP7_75t_L g1077 ( .A(n_11), .Y(n_1077) );
AOI22xp33_ASAP7_75t_SL g993 ( .A1(n_12), .A2(n_239), .B1(n_994), .B2(n_995), .Y(n_993) );
INVxp67_ASAP7_75t_SL g1024 ( .A(n_12), .Y(n_1024) );
AOI22xp33_ASAP7_75t_L g1183 ( .A1(n_13), .A2(n_311), .B1(n_1181), .B2(n_1184), .Y(n_1183) );
AOI221xp5_ASAP7_75t_L g1189 ( .A1(n_13), .A2(n_95), .B1(n_613), .B2(n_766), .C(n_1190), .Y(n_1189) );
AOI22xp33_ASAP7_75t_L g718 ( .A1(n_14), .A2(n_353), .B1(n_527), .B2(n_719), .Y(n_718) );
INVx1_ASAP7_75t_L g739 ( .A(n_14), .Y(n_739) );
INVx2_ASAP7_75t_L g422 ( .A(n_15), .Y(n_422) );
INVx1_ASAP7_75t_L g1816 ( .A(n_16), .Y(n_1816) );
OAI322xp33_ASAP7_75t_L g1818 ( .A1(n_16), .A2(n_599), .A3(n_735), .B1(n_1400), .B2(n_1819), .C1(n_1824), .C2(n_1829), .Y(n_1818) );
OAI22xp5_ASAP7_75t_SL g1287 ( .A1(n_17), .A2(n_303), .B1(n_682), .B2(n_1288), .Y(n_1287) );
OAI221xp5_ASAP7_75t_L g1299 ( .A1(n_17), .A2(n_303), .B1(n_623), .B2(n_1300), .C(n_1301), .Y(n_1299) );
XNOR2x1_ASAP7_75t_L g1266 ( .A(n_18), .B(n_1267), .Y(n_1266) );
INVx1_ASAP7_75t_L g1037 ( .A(n_19), .Y(n_1037) );
OAI222xp33_ASAP7_75t_L g1061 ( .A1(n_19), .A2(n_178), .B1(n_625), .B2(n_724), .C1(n_1062), .C2(n_1067), .Y(n_1061) );
INVx1_ASAP7_75t_L g1245 ( .A(n_20), .Y(n_1245) );
AOI221xp5_ASAP7_75t_L g1810 ( .A1(n_21), .A2(n_259), .B1(n_1190), .B2(n_1255), .C(n_1811), .Y(n_1810) );
INVx1_ASAP7_75t_L g1828 ( .A(n_21), .Y(n_1828) );
AOI22xp33_ASAP7_75t_L g1182 ( .A1(n_22), .A2(n_244), .B1(n_589), .B2(n_1179), .Y(n_1182) );
AOI22xp33_ASAP7_75t_L g1191 ( .A1(n_22), .A2(n_160), .B1(n_1192), .B2(n_1194), .Y(n_1191) );
AOI22xp33_ASAP7_75t_L g1497 ( .A1(n_23), .A2(n_328), .B1(n_527), .B2(n_1115), .Y(n_1497) );
INVx1_ASAP7_75t_L g1517 ( .A(n_23), .Y(n_1517) );
INVx1_ASAP7_75t_L g965 ( .A(n_24), .Y(n_965) );
OAI22xp33_ASAP7_75t_L g592 ( .A1(n_25), .A2(n_280), .B1(n_593), .B2(n_599), .Y(n_592) );
INVx1_ASAP7_75t_L g617 ( .A(n_25), .Y(n_617) );
INVx1_ASAP7_75t_L g1243 ( .A(n_26), .Y(n_1243) );
AOI22xp33_ASAP7_75t_L g1256 ( .A1(n_26), .A2(n_80), .B1(n_1010), .B2(n_1257), .Y(n_1256) );
INVx1_ASAP7_75t_L g1499 ( .A(n_27), .Y(n_1499) );
INVx1_ASAP7_75t_L g429 ( .A(n_28), .Y(n_429) );
AOI22xp5_ASAP7_75t_L g1611 ( .A1(n_29), .A2(n_236), .B1(n_1587), .B2(n_1590), .Y(n_1611) );
CKINVDCx5p33_ASAP7_75t_R g1217 ( .A(n_30), .Y(n_1217) );
HB1xp67_ASAP7_75t_L g386 ( .A(n_31), .Y(n_386) );
AND2x2_ASAP7_75t_L g1581 ( .A(n_31), .B(n_384), .Y(n_1581) );
INVx1_ASAP7_75t_L g1298 ( .A(n_32), .Y(n_1298) );
AOI22xp5_ASAP7_75t_L g1628 ( .A1(n_33), .A2(n_205), .B1(n_1587), .B2(n_1590), .Y(n_1628) );
OAI211xp5_ASAP7_75t_SL g1547 ( .A1(n_34), .A2(n_607), .B(n_1548), .C(n_1552), .Y(n_1547) );
OAI22xp5_ASAP7_75t_L g1557 ( .A1(n_34), .A2(n_293), .B1(n_412), .B2(n_656), .Y(n_1557) );
OAI22xp5_ASAP7_75t_SL g932 ( .A1(n_35), .A2(n_312), .B1(n_933), .B2(n_934), .Y(n_932) );
INVxp67_ASAP7_75t_SL g969 ( .A(n_35), .Y(n_969) );
AOI22xp33_ASAP7_75t_L g1813 ( .A1(n_36), .A2(n_318), .B1(n_1009), .B2(n_1814), .Y(n_1813) );
INVxp67_ASAP7_75t_L g1823 ( .A(n_36), .Y(n_1823) );
CKINVDCx5p33_ASAP7_75t_R g974 ( .A(n_37), .Y(n_974) );
INVx1_ASAP7_75t_L g1855 ( .A(n_38), .Y(n_1855) );
OAI211xp5_ASAP7_75t_L g1863 ( .A1(n_38), .A2(n_1014), .B(n_1060), .C(n_1864), .Y(n_1863) );
INVxp67_ASAP7_75t_L g1085 ( .A(n_39), .Y(n_1085) );
AOI22xp5_ASAP7_75t_L g1603 ( .A1(n_40), .A2(n_296), .B1(n_1587), .B2(n_1590), .Y(n_1603) );
INVx1_ASAP7_75t_L g1797 ( .A(n_40), .Y(n_1797) );
AOI22xp33_ASAP7_75t_L g1845 ( .A1(n_40), .A2(n_1846), .B1(n_1849), .B2(n_1891), .Y(n_1845) );
CKINVDCx5p33_ASAP7_75t_R g1403 ( .A(n_41), .Y(n_1403) );
AOI22xp33_ASAP7_75t_L g1804 ( .A1(n_42), .A2(n_315), .B1(n_1009), .B2(n_1805), .Y(n_1804) );
AOI22xp33_ASAP7_75t_L g1833 ( .A1(n_42), .A2(n_259), .B1(n_463), .B2(n_1834), .Y(n_1833) );
AOI21xp33_ASAP7_75t_L g1353 ( .A1(n_43), .A2(n_643), .B(n_768), .Y(n_1353) );
AOI22xp33_ASAP7_75t_L g1374 ( .A1(n_43), .A2(n_341), .B1(n_589), .B2(n_807), .Y(n_1374) );
AOI221xp5_ASAP7_75t_L g1492 ( .A1(n_44), .A2(n_132), .B1(n_613), .B2(n_1358), .C(n_1493), .Y(n_1492) );
INVx1_ASAP7_75t_L g1518 ( .A(n_44), .Y(n_1518) );
INVx1_ASAP7_75t_L g1058 ( .A(n_45), .Y(n_1058) );
AOI22xp33_ASAP7_75t_L g1140 ( .A1(n_46), .A2(n_112), .B1(n_1091), .B2(n_1141), .Y(n_1140) );
AOI221xp5_ASAP7_75t_L g1162 ( .A1(n_46), .A2(n_209), .B1(n_644), .B2(n_1113), .C(n_1163), .Y(n_1162) );
NOR2xp33_ASAP7_75t_L g1536 ( .A(n_47), .B(n_431), .Y(n_1536) );
INVx1_ASAP7_75t_L g1366 ( .A(n_48), .Y(n_1366) );
AOI221xp5_ASAP7_75t_L g1876 ( .A1(n_49), .A2(n_331), .B1(n_766), .B2(n_768), .C(n_1190), .Y(n_1876) );
INVxp67_ASAP7_75t_SL g1884 ( .A(n_49), .Y(n_1884) );
AOI22xp5_ASAP7_75t_L g1621 ( .A1(n_50), .A2(n_140), .B1(n_1587), .B2(n_1590), .Y(n_1621) );
INVx1_ASAP7_75t_L g1860 ( .A(n_51), .Y(n_1860) );
OAI22xp5_ASAP7_75t_L g1877 ( .A1(n_51), .A2(n_226), .B1(n_607), .B2(n_1878), .Y(n_1877) );
CKINVDCx5p33_ASAP7_75t_R g1393 ( .A(n_52), .Y(n_1393) );
OAI211xp5_ASAP7_75t_SL g1422 ( .A1(n_53), .A2(n_1202), .B(n_1423), .C(n_1426), .Y(n_1422) );
INVx1_ASAP7_75t_L g1472 ( .A(n_53), .Y(n_1472) );
CKINVDCx5p33_ASAP7_75t_R g1399 ( .A(n_54), .Y(n_1399) );
INVx1_ASAP7_75t_L g722 ( .A(n_55), .Y(n_722) );
AOI22xp33_ASAP7_75t_L g990 ( .A1(n_56), .A2(n_302), .B1(n_588), .B2(n_792), .Y(n_990) );
INVx1_ASAP7_75t_L g1017 ( .A(n_56), .Y(n_1017) );
NAND5xp2_ASAP7_75t_L g757 ( .A(n_57), .B(n_758), .C(n_788), .D(n_803), .E(n_813), .Y(n_757) );
INVx1_ASAP7_75t_L g822 ( .A(n_57), .Y(n_822) );
AOI22xp5_ASAP7_75t_L g1619 ( .A1(n_57), .A2(n_181), .B1(n_1580), .B2(n_1620), .Y(n_1619) );
OAI22xp5_ASAP7_75t_L g603 ( .A1(n_58), .A2(n_163), .B1(n_558), .B2(n_604), .Y(n_603) );
OAI211xp5_ASAP7_75t_SL g606 ( .A1(n_58), .A2(n_607), .B(n_608), .C(n_615), .Y(n_606) );
INVx1_ASAP7_75t_L g721 ( .A(n_59), .Y(n_721) );
INVx1_ASAP7_75t_L g1057 ( .A(n_60), .Y(n_1057) );
INVxp67_ASAP7_75t_SL g1875 ( .A(n_61), .Y(n_1875) );
AOI22xp33_ASAP7_75t_L g1890 ( .A1(n_61), .A2(n_158), .B1(n_1181), .B2(n_1286), .Y(n_1890) );
BUFx6f_ASAP7_75t_L g398 ( .A(n_62), .Y(n_398) );
INVx1_ASAP7_75t_L g1363 ( .A(n_64), .Y(n_1363) );
OAI22xp33_ASAP7_75t_L g1378 ( .A1(n_64), .A2(n_330), .B1(n_805), .B2(n_1379), .Y(n_1378) );
XOR2xp5_ASAP7_75t_L g573 ( .A(n_65), .B(n_574), .Y(n_573) );
INVx1_ASAP7_75t_L g982 ( .A(n_66), .Y(n_982) );
INVx1_ASAP7_75t_L g1172 ( .A(n_67), .Y(n_1172) );
OAI222xp33_ASAP7_75t_L g1200 ( .A1(n_67), .A2(n_372), .B1(n_624), .B2(n_724), .C1(n_1201), .C2(n_1205), .Y(n_1200) );
AOI22xp33_ASAP7_75t_SL g584 ( .A1(n_68), .A2(n_308), .B1(n_585), .B2(n_588), .Y(n_584) );
AOI221xp5_ASAP7_75t_L g639 ( .A1(n_68), .A2(n_275), .B1(n_640), .B2(n_642), .C(n_644), .Y(n_639) );
INVx1_ASAP7_75t_L g1297 ( .A(n_69), .Y(n_1297) );
INVx1_ASAP7_75t_L g1431 ( .A(n_70), .Y(n_1431) );
OAI211xp5_ASAP7_75t_L g1459 ( .A1(n_70), .A2(n_1460), .B(n_1462), .C(n_1464), .Y(n_1459) );
XOR2x2_ASAP7_75t_L g1380 ( .A(n_71), .B(n_1381), .Y(n_1380) );
AOI22xp33_ASAP7_75t_L g1579 ( .A1(n_71), .A2(n_262), .B1(n_1580), .B2(n_1584), .Y(n_1579) );
INVx1_ASAP7_75t_L g1504 ( .A(n_72), .Y(n_1504) );
OAI332xp33_ASAP7_75t_SL g1508 ( .A1(n_72), .A2(n_593), .A3(n_735), .B1(n_798), .B2(n_1509), .B3(n_1515), .C1(n_1521), .C2(n_1525), .Y(n_1508) );
CKINVDCx5p33_ASAP7_75t_R g1199 ( .A(n_73), .Y(n_1199) );
AOI221xp5_ASAP7_75t_L g1549 ( .A1(n_74), .A2(n_134), .B1(n_524), .B2(n_612), .C(n_1550), .Y(n_1549) );
AOI22xp33_ASAP7_75t_L g1566 ( .A1(n_74), .A2(n_268), .B1(n_465), .B2(n_1564), .Y(n_1566) );
AOI221xp5_ASAP7_75t_L g765 ( .A1(n_75), .A2(n_179), .B1(n_520), .B2(n_766), .C(n_768), .Y(n_765) );
AOI22xp33_ASAP7_75t_L g793 ( .A1(n_75), .A2(n_255), .B1(n_589), .B2(n_794), .Y(n_793) );
INVx1_ASAP7_75t_L g493 ( .A(n_76), .Y(n_493) );
CKINVDCx5p33_ASAP7_75t_R g1149 ( .A(n_77), .Y(n_1149) );
AOI22xp33_ASAP7_75t_L g769 ( .A1(n_78), .A2(n_255), .B1(n_719), .B2(n_770), .Y(n_769) );
AOI22xp33_ASAP7_75t_L g791 ( .A1(n_78), .A2(n_179), .B1(n_589), .B2(n_792), .Y(n_791) );
AOI22xp33_ASAP7_75t_L g1097 ( .A1(n_79), .A2(n_171), .B1(n_588), .B2(n_1090), .Y(n_1097) );
AOI21xp33_ASAP7_75t_L g1121 ( .A1(n_79), .A2(n_703), .B(n_1122), .Y(n_1121) );
INVx1_ASAP7_75t_L g1233 ( .A(n_80), .Y(n_1233) );
INVx1_ASAP7_75t_L g1136 ( .A(n_81), .Y(n_1136) );
AOI22xp33_ASAP7_75t_L g1494 ( .A1(n_82), .A2(n_274), .B1(n_527), .B2(n_1115), .Y(n_1494) );
INVx1_ASAP7_75t_L g1524 ( .A(n_82), .Y(n_1524) );
AOI22xp33_ASAP7_75t_L g1354 ( .A1(n_83), .A2(n_113), .B1(n_530), .B2(n_1257), .Y(n_1354) );
AOI22xp33_ASAP7_75t_L g1377 ( .A1(n_83), .A2(n_253), .B1(n_465), .B2(n_994), .Y(n_1377) );
AOI22xp33_ASAP7_75t_SL g462 ( .A1(n_84), .A2(n_309), .B1(n_463), .B2(n_465), .Y(n_462) );
AOI22xp33_ASAP7_75t_L g535 ( .A1(n_84), .A2(n_327), .B1(n_529), .B2(n_536), .Y(n_535) );
AOI22xp33_ASAP7_75t_SL g985 ( .A1(n_85), .A2(n_185), .B1(n_744), .B2(n_986), .Y(n_985) );
INVxp67_ASAP7_75t_SL g1023 ( .A(n_85), .Y(n_1023) );
INVx1_ASAP7_75t_L g1501 ( .A(n_86), .Y(n_1501) );
CKINVDCx5p33_ASAP7_75t_R g1836 ( .A(n_87), .Y(n_1836) );
INVx1_ASAP7_75t_L g1807 ( .A(n_88), .Y(n_1807) );
OAI211xp5_ASAP7_75t_L g1837 ( .A1(n_88), .A2(n_450), .B(n_593), .C(n_1838), .Y(n_1837) );
CKINVDCx5p33_ASAP7_75t_R g1100 ( .A(n_89), .Y(n_1100) );
CKINVDCx5p33_ASAP7_75t_R g779 ( .A(n_90), .Y(n_779) );
OAI21xp5_ASAP7_75t_SL g1127 ( .A1(n_91), .A2(n_558), .B(n_1128), .Y(n_1127) );
CKINVDCx5p33_ASAP7_75t_R g1396 ( .A(n_92), .Y(n_1396) );
AOI22xp33_ASAP7_75t_SL g1096 ( .A1(n_93), .A2(n_281), .B1(n_956), .B2(n_995), .Y(n_1096) );
AOI22xp33_ASAP7_75t_L g1120 ( .A1(n_93), .A2(n_334), .B1(n_690), .B2(n_705), .Y(n_1120) );
OR2x2_ASAP7_75t_L g1858 ( .A(n_94), .B(n_431), .Y(n_1858) );
AOI22xp33_ASAP7_75t_L g1178 ( .A1(n_95), .A2(n_152), .B1(n_1179), .B2(n_1181), .Y(n_1178) );
OAI221xp5_ASAP7_75t_L g1870 ( .A1(n_96), .A2(n_224), .B1(n_1300), .B2(n_1871), .C(n_1872), .Y(n_1870) );
OAI322xp33_ASAP7_75t_L g1882 ( .A1(n_96), .A2(n_599), .A3(n_950), .B1(n_1247), .B2(n_1883), .C1(n_1886), .C2(n_1888), .Y(n_1882) );
AOI22xp33_ASAP7_75t_L g1599 ( .A1(n_97), .A2(n_182), .B1(n_1580), .B2(n_1587), .Y(n_1599) );
AOI22xp33_ASAP7_75t_SL g1323 ( .A1(n_98), .A2(n_217), .B1(n_589), .B2(n_792), .Y(n_1323) );
AOI22xp33_ASAP7_75t_L g1334 ( .A1(n_98), .A2(n_109), .B1(n_527), .B2(n_530), .Y(n_1334) );
OAI21xp5_ASAP7_75t_L g557 ( .A1(n_99), .A2(n_558), .B(n_567), .Y(n_557) );
AOI22xp33_ASAP7_75t_SL g937 ( .A1(n_100), .A2(n_172), .B1(n_515), .B2(n_938), .Y(n_937) );
INVxp67_ASAP7_75t_SL g961 ( .A(n_100), .Y(n_961) );
INVx1_ASAP7_75t_L g1270 ( .A(n_101), .Y(n_1270) );
AOI22xp33_ASAP7_75t_SL g1278 ( .A1(n_102), .A2(n_305), .B1(n_671), .B2(n_963), .Y(n_1278) );
AOI221xp5_ASAP7_75t_L g1293 ( .A1(n_102), .A2(n_111), .B1(n_519), .B2(n_643), .C(n_773), .Y(n_1293) );
INVx1_ASAP7_75t_L g1027 ( .A(n_103), .Y(n_1027) );
AOI22xp33_ASAP7_75t_L g1598 ( .A1(n_104), .A2(n_322), .B1(n_1584), .B2(n_1590), .Y(n_1598) );
AOI22xp33_ASAP7_75t_L g680 ( .A1(n_105), .A2(n_292), .B1(n_463), .B2(n_671), .Y(n_680) );
AOI221xp5_ASAP7_75t_L g688 ( .A1(n_105), .A2(n_288), .B1(n_523), .B2(n_524), .C(n_612), .Y(n_688) );
AOI22xp5_ASAP7_75t_L g1605 ( .A1(n_106), .A2(n_168), .B1(n_1580), .B2(n_1606), .Y(n_1605) );
OAI21xp33_ASAP7_75t_L g1213 ( .A1(n_107), .A2(n_1214), .B(n_1215), .Y(n_1213) );
INVx1_ASAP7_75t_L g1272 ( .A(n_108), .Y(n_1272) );
AOI22xp33_ASAP7_75t_SL g1326 ( .A1(n_109), .A2(n_310), .B1(n_589), .B2(n_792), .Y(n_1326) );
INVx1_ASAP7_75t_L g669 ( .A(n_110), .Y(n_669) );
AOI22xp33_ASAP7_75t_L g689 ( .A1(n_110), .A2(n_320), .B1(n_530), .B2(n_690), .Y(n_689) );
AOI22xp33_ASAP7_75t_L g1285 ( .A1(n_111), .A2(n_199), .B1(n_744), .B2(n_1286), .Y(n_1285) );
AOI22xp33_ASAP7_75t_SL g1156 ( .A1(n_112), .A2(n_157), .B1(n_527), .B2(n_529), .Y(n_1156) );
AOI22xp33_ASAP7_75t_L g1373 ( .A1(n_113), .A2(n_279), .B1(n_452), .B2(n_986), .Y(n_1373) );
AOI22xp33_ASAP7_75t_SL g1047 ( .A1(n_114), .A2(n_346), .B1(n_463), .B2(n_671), .Y(n_1047) );
INVxp67_ASAP7_75t_SL g1052 ( .A(n_114), .Y(n_1052) );
INVx1_ASAP7_75t_L g1242 ( .A(n_115), .Y(n_1242) );
AOI221xp5_ASAP7_75t_L g1251 ( .A1(n_115), .A2(n_242), .B1(n_703), .B2(n_1111), .C(n_1190), .Y(n_1251) );
CKINVDCx5p33_ASAP7_75t_R g1108 ( .A(n_116), .Y(n_1108) );
CKINVDCx5p33_ASAP7_75t_R g1319 ( .A(n_117), .Y(n_1319) );
XNOR2xp5_ASAP7_75t_L g709 ( .A(n_118), .B(n_710), .Y(n_709) );
AOI22xp33_ASAP7_75t_L g466 ( .A1(n_119), .A2(n_337), .B1(n_467), .B2(n_472), .Y(n_466) );
AOI221xp5_ASAP7_75t_L g537 ( .A1(n_119), .A2(n_360), .B1(n_538), .B2(n_542), .C(n_546), .Y(n_537) );
OAI211xp5_ASAP7_75t_L g775 ( .A1(n_120), .A2(n_776), .B(n_777), .C(n_778), .Y(n_775) );
INVx1_ASAP7_75t_L g818 ( .A(n_120), .Y(n_818) );
INVx1_ASAP7_75t_L g1873 ( .A(n_121), .Y(n_1873) );
AOI22xp33_ASAP7_75t_L g1586 ( .A1(n_122), .A2(n_352), .B1(n_1587), .B2(n_1590), .Y(n_1586) );
CKINVDCx5p33_ASAP7_75t_R g1103 ( .A(n_123), .Y(n_1103) );
OAI22xp5_ASAP7_75t_L g1124 ( .A1(n_123), .A2(n_144), .B1(n_549), .B2(n_1125), .Y(n_1124) );
AOI22xp33_ASAP7_75t_L g943 ( .A1(n_124), .A2(n_252), .B1(n_515), .B2(n_692), .Y(n_943) );
AOI22xp33_ASAP7_75t_L g955 ( .A1(n_124), .A2(n_277), .B1(n_486), .B2(n_956), .Y(n_955) );
INVx1_ASAP7_75t_L g1542 ( .A(n_125), .Y(n_1542) );
AOI21xp33_ASAP7_75t_L g730 ( .A1(n_126), .A2(n_523), .B(n_546), .Y(n_730) );
INVx1_ASAP7_75t_L g738 ( .A(n_126), .Y(n_738) );
AOI22xp33_ASAP7_75t_L g485 ( .A1(n_127), .A2(n_327), .B1(n_463), .B2(n_486), .Y(n_485) );
AOI221xp5_ASAP7_75t_L g518 ( .A1(n_127), .A2(n_309), .B1(n_519), .B2(n_522), .C(n_524), .Y(n_518) );
INVx1_ASAP7_75t_L g654 ( .A(n_128), .Y(n_654) );
INVx1_ASAP7_75t_L g924 ( .A(n_129), .Y(n_924) );
INVx1_ASAP7_75t_L g384 ( .A(n_130), .Y(n_384) );
AOI221xp5_ASAP7_75t_L g714 ( .A1(n_131), .A2(n_273), .B1(n_524), .B2(n_715), .C(n_716), .Y(n_714) );
AOI22xp33_ASAP7_75t_L g740 ( .A1(n_131), .A2(n_187), .B1(n_452), .B2(n_463), .Y(n_740) );
INVx1_ASAP7_75t_L g1530 ( .A(n_132), .Y(n_1530) );
INVx1_ASAP7_75t_L g1315 ( .A(n_133), .Y(n_1315) );
AOI22xp33_ASAP7_75t_L g1563 ( .A1(n_134), .A2(n_283), .B1(n_452), .B2(n_1564), .Y(n_1563) );
INVx1_ASAP7_75t_L g1314 ( .A(n_135), .Y(n_1314) );
INVx1_ASAP7_75t_L g1553 ( .A(n_136), .Y(n_1553) );
OAI22xp33_ASAP7_75t_L g1568 ( .A1(n_136), .A2(n_192), .B1(n_593), .B2(n_805), .Y(n_1568) );
AOI22xp33_ASAP7_75t_SL g591 ( .A1(n_137), .A2(n_307), .B1(n_463), .B2(n_465), .Y(n_591) );
INVxp67_ASAP7_75t_SL g638 ( .A(n_137), .Y(n_638) );
AOI221xp5_ASAP7_75t_L g1321 ( .A1(n_138), .A2(n_306), .B1(n_465), .B2(n_1286), .C(n_1322), .Y(n_1321) );
AOI221xp5_ASAP7_75t_L g1333 ( .A1(n_138), .A2(n_250), .B1(n_544), .B2(n_612), .C(n_773), .Y(n_1333) );
AOI22xp33_ASAP7_75t_L g988 ( .A1(n_139), .A2(n_193), .B1(n_792), .B2(n_989), .Y(n_988) );
INVx1_ASAP7_75t_L g1021 ( .A(n_139), .Y(n_1021) );
OAI22xp33_ASAP7_75t_L g1229 ( .A1(n_141), .A2(n_324), .B1(n_593), .B2(n_1230), .Y(n_1229) );
INVx1_ASAP7_75t_L g1259 ( .A(n_141), .Y(n_1259) );
OAI222xp33_ASAP7_75t_L g865 ( .A1(n_142), .A2(n_355), .B1(n_866), .B2(n_868), .C1(n_870), .C2(n_872), .Y(n_865) );
INVx1_ASAP7_75t_L g885 ( .A(n_142), .Y(n_885) );
CKINVDCx5p33_ASAP7_75t_R g1391 ( .A(n_143), .Y(n_1391) );
CKINVDCx5p33_ASAP7_75t_R g1102 ( .A(n_144), .Y(n_1102) );
INVx1_ASAP7_75t_L g1350 ( .A(n_145), .Y(n_1350) );
OAI211xp5_ASAP7_75t_L g1355 ( .A1(n_146), .A2(n_686), .B(n_1356), .C(n_1362), .Y(n_1355) );
OAI22xp5_ASAP7_75t_L g1367 ( .A1(n_146), .A2(n_285), .B1(n_412), .B2(n_656), .Y(n_1367) );
INVx1_ASAP7_75t_L g850 ( .A(n_147), .Y(n_850) );
OAI211xp5_ASAP7_75t_L g926 ( .A1(n_148), .A2(n_927), .B(n_928), .C(n_929), .Y(n_926) );
INVxp33_ASAP7_75t_SL g947 ( .A(n_148), .Y(n_947) );
CKINVDCx5p33_ASAP7_75t_R g676 ( .A(n_149), .Y(n_676) );
INVx1_ASAP7_75t_L g1235 ( .A(n_150), .Y(n_1235) );
AOI221xp5_ASAP7_75t_L g1254 ( .A1(n_150), .A2(n_300), .B1(n_1163), .B2(n_1190), .C(n_1255), .Y(n_1254) );
AOI22xp33_ASAP7_75t_SL g1602 ( .A1(n_151), .A2(n_228), .B1(n_1580), .B2(n_1584), .Y(n_1602) );
INVx1_ASAP7_75t_L g1204 ( .A(n_152), .Y(n_1204) );
INVx1_ASAP7_75t_L g664 ( .A(n_153), .Y(n_664) );
AOI21xp33_ASAP7_75t_L g702 ( .A1(n_153), .A2(n_523), .B(n_703), .Y(n_702) );
INVxp67_ASAP7_75t_SL g1352 ( .A(n_154), .Y(n_1352) );
AOI22xp33_ASAP7_75t_SL g1375 ( .A1(n_154), .A2(n_297), .B1(n_469), .B2(n_589), .Y(n_1375) );
OAI22xp5_ASAP7_75t_L g655 ( .A1(n_155), .A2(n_177), .B1(n_604), .B2(n_656), .Y(n_655) );
OAI211xp5_ASAP7_75t_L g685 ( .A1(n_155), .A2(n_686), .B(n_687), .C(n_693), .Y(n_685) );
INVx1_ASAP7_75t_L g978 ( .A(n_156), .Y(n_978) );
OAI222xp33_ASAP7_75t_L g1013 ( .A1(n_156), .A2(n_222), .B1(n_624), .B2(n_1014), .C1(n_1015), .C2(n_1022), .Y(n_1013) );
AOI22xp33_ASAP7_75t_L g1143 ( .A1(n_157), .A2(n_209), .B1(n_1091), .B2(n_1144), .Y(n_1143) );
AOI221xp5_ASAP7_75t_L g1869 ( .A1(n_158), .A2(n_237), .B1(n_519), .B2(n_524), .C(n_766), .Y(n_1869) );
INVx1_ASAP7_75t_L g1806 ( .A(n_159), .Y(n_1806) );
AOI22xp33_ASAP7_75t_SL g1177 ( .A1(n_160), .A2(n_246), .B1(n_589), .B2(n_994), .Y(n_1177) );
OA21x2_ASAP7_75t_L g1268 ( .A1(n_161), .A2(n_431), .B(n_1269), .Y(n_1268) );
CKINVDCx5p33_ASAP7_75t_R g1430 ( .A(n_162), .Y(n_1430) );
OAI22xp33_ASAP7_75t_L g1444 ( .A1(n_164), .A2(n_325), .B1(n_1445), .B2(n_1446), .Y(n_1444) );
OAI22xp33_ASAP7_75t_L g1452 ( .A1(n_164), .A2(n_325), .B1(n_1453), .B2(n_1456), .Y(n_1452) );
INVx1_ASAP7_75t_L g1000 ( .A(n_165), .Y(n_1000) );
AOI221xp5_ASAP7_75t_L g1803 ( .A1(n_166), .A2(n_231), .B1(n_519), .B2(n_703), .C(n_1118), .Y(n_1803) );
INVxp67_ASAP7_75t_L g1820 ( .A(n_166), .Y(n_1820) );
OAI221xp5_ASAP7_75t_L g723 ( .A1(n_167), .A2(n_363), .B1(n_625), .B2(n_724), .C(n_725), .Y(n_723) );
OAI22xp33_ASAP7_75t_L g746 ( .A1(n_167), .A2(n_363), .B1(n_490), .B2(n_682), .Y(n_746) );
INVx1_ASAP7_75t_L g1218 ( .A(n_168), .Y(n_1218) );
AO22x1_ASAP7_75t_L g1089 ( .A1(n_169), .A2(n_208), .B1(n_1090), .B2(n_1091), .Y(n_1089) );
NAND2xp5_ASAP7_75t_L g1117 ( .A(n_169), .B(n_1118), .Y(n_1117) );
INVx1_ASAP7_75t_L g812 ( .A(n_170), .Y(n_812) );
AOI22xp33_ASAP7_75t_SL g1114 ( .A1(n_171), .A2(n_208), .B1(n_536), .B2(n_1115), .Y(n_1114) );
INVx1_ASAP7_75t_L g954 ( .A(n_172), .Y(n_954) );
CKINVDCx5p33_ASAP7_75t_R g602 ( .A(n_173), .Y(n_602) );
OA22x2_ASAP7_75t_L g1537 ( .A1(n_174), .A2(n_1538), .B1(n_1569), .B2(n_1570), .Y(n_1537) );
CKINVDCx16_ASAP7_75t_R g1569 ( .A(n_174), .Y(n_1569) );
CKINVDCx5p33_ASAP7_75t_R g931 ( .A(n_175), .Y(n_931) );
OAI211xp5_ASAP7_75t_L g1348 ( .A1(n_176), .A2(n_621), .B(n_1349), .C(n_1351), .Y(n_1348) );
INVx1_ASAP7_75t_L g1371 ( .A(n_176), .Y(n_1371) );
INVx1_ASAP7_75t_L g1036 ( .A(n_178), .Y(n_1036) );
INVx1_ASAP7_75t_L g844 ( .A(n_180), .Y(n_844) );
AOI22xp33_ASAP7_75t_L g902 ( .A1(n_180), .A2(n_282), .B1(n_719), .B2(n_770), .Y(n_902) );
INVx1_ASAP7_75t_L g572 ( .A(n_182), .Y(n_572) );
INVx1_ASAP7_75t_L g1556 ( .A(n_183), .Y(n_1556) );
OAI22xp5_ASAP7_75t_L g1434 ( .A1(n_184), .A2(n_294), .B1(n_1435), .B2(n_1439), .Y(n_1434) );
OAI22xp33_ASAP7_75t_L g1473 ( .A1(n_184), .A2(n_294), .B1(n_1474), .B2(n_1477), .Y(n_1473) );
AOI221xp5_ASAP7_75t_L g1007 ( .A1(n_185), .A2(n_239), .B1(n_613), .B2(n_640), .C(n_642), .Y(n_1007) );
CKINVDCx5p33_ASAP7_75t_R g930 ( .A(n_186), .Y(n_930) );
AOI22xp33_ASAP7_75t_SL g731 ( .A1(n_187), .A2(n_333), .B1(n_515), .B2(n_536), .Y(n_731) );
OAI211xp5_ASAP7_75t_L g712 ( .A1(n_188), .A2(n_686), .B(n_713), .C(n_720), .Y(n_712) );
OAI22xp5_ASAP7_75t_L g749 ( .A1(n_188), .A2(n_358), .B1(n_604), .B2(n_656), .Y(n_749) );
INVx1_ASAP7_75t_L g941 ( .A(n_189), .Y(n_941) );
INVx1_ASAP7_75t_L g1277 ( .A(n_190), .Y(n_1277) );
AOI221xp5_ASAP7_75t_L g1307 ( .A1(n_190), .A2(n_241), .B1(n_538), .B2(n_544), .C(n_644), .Y(n_1307) );
OAI211xp5_ASAP7_75t_L g759 ( .A1(n_191), .A2(n_760), .B(n_763), .C(n_774), .Y(n_759) );
NOR2xp33_ASAP7_75t_L g787 ( .A(n_191), .B(n_412), .Y(n_787) );
INVx1_ASAP7_75t_L g1554 ( .A(n_192), .Y(n_1554) );
AOI22xp33_ASAP7_75t_L g1008 ( .A1(n_193), .A2(n_302), .B1(n_1009), .B2(n_1010), .Y(n_1008) );
AOI221xp5_ASAP7_75t_L g1324 ( .A1(n_194), .A2(n_250), .B1(n_744), .B2(n_1286), .C(n_1325), .Y(n_1324) );
AOI22xp33_ASAP7_75t_L g1336 ( .A1(n_194), .A2(n_306), .B1(n_530), .B2(n_938), .Y(n_1336) );
INVx2_ASAP7_75t_L g1583 ( .A(n_195), .Y(n_1583) );
AND2x2_ASAP7_75t_L g1585 ( .A(n_195), .B(n_321), .Y(n_1585) );
AND2x2_ASAP7_75t_L g1591 ( .A(n_195), .B(n_1589), .Y(n_1591) );
AOI22xp33_ASAP7_75t_L g1043 ( .A1(n_196), .A2(n_365), .B1(n_1044), .B2(n_1045), .Y(n_1043) );
INVx1_ASAP7_75t_L g1065 ( .A(n_196), .Y(n_1065) );
CKINVDCx5p33_ASAP7_75t_R g1881 ( .A(n_197), .Y(n_1881) );
INVx1_ASAP7_75t_L g695 ( .A(n_198), .Y(n_695) );
INVx1_ASAP7_75t_L g1306 ( .A(n_199), .Y(n_1306) );
XNOR2xp5_ASAP7_75t_L g1345 ( .A(n_200), .B(n_1346), .Y(n_1345) );
INVx1_ASAP7_75t_L g507 ( .A(n_201), .Y(n_507) );
OAI22xp5_ASAP7_75t_L g1150 ( .A1(n_202), .A2(n_304), .B1(n_412), .B2(n_558), .Y(n_1150) );
OAI211xp5_ASAP7_75t_L g1152 ( .A1(n_202), .A2(n_607), .B(n_1153), .C(n_1157), .Y(n_1152) );
AOI22xp5_ASAP7_75t_L g1613 ( .A1(n_203), .A2(n_269), .B1(n_1580), .B2(n_1590), .Y(n_1613) );
XOR2x2_ASAP7_75t_L g1486 ( .A(n_204), .B(n_1487), .Y(n_1486) );
CKINVDCx5p33_ASAP7_75t_R g1107 ( .A(n_206), .Y(n_1107) );
AOI22xp33_ASAP7_75t_L g477 ( .A1(n_207), .A2(n_360), .B1(n_467), .B2(n_478), .Y(n_477) );
AOI22xp33_ASAP7_75t_L g526 ( .A1(n_207), .A2(n_337), .B1(n_527), .B2(n_529), .Y(n_526) );
INVx1_ASAP7_75t_L g913 ( .A(n_210), .Y(n_913) );
AOI22xp33_ASAP7_75t_L g1614 ( .A1(n_211), .A2(n_219), .B1(n_1587), .B2(n_1606), .Y(n_1614) );
INVx1_ASAP7_75t_L g999 ( .A(n_212), .Y(n_999) );
AOI22xp33_ASAP7_75t_L g764 ( .A1(n_213), .A2(n_299), .B1(n_692), .B2(n_719), .Y(n_764) );
AOI22xp33_ASAP7_75t_SL g795 ( .A1(n_213), .A2(n_319), .B1(n_463), .B2(n_796), .Y(n_795) );
AOI22xp33_ASAP7_75t_SL g670 ( .A1(n_214), .A2(n_288), .B1(n_463), .B2(n_671), .Y(n_670) );
AOI22xp33_ASAP7_75t_SL g704 ( .A1(n_214), .A2(n_292), .B1(n_536), .B2(n_705), .Y(n_704) );
INVx1_ASAP7_75t_L g1076 ( .A(n_215), .Y(n_1076) );
AOI21xp33_ASAP7_75t_L g1545 ( .A1(n_216), .A2(n_546), .B(n_716), .Y(n_1545) );
AOI22xp33_ASAP7_75t_L g1565 ( .A1(n_216), .A2(n_342), .B1(n_589), .B2(n_807), .Y(n_1565) );
AOI221xp5_ASAP7_75t_L g1337 ( .A1(n_217), .A2(n_310), .B1(n_544), .B2(n_703), .C(n_715), .Y(n_1337) );
INVx1_ASAP7_75t_L g1239 ( .A(n_218), .Y(n_1239) );
OAI211xp5_ASAP7_75t_L g1540 ( .A1(n_220), .A2(n_621), .B(n_1541), .C(n_1543), .Y(n_1540) );
INVx1_ASAP7_75t_L g1561 ( .A(n_220), .Y(n_1561) );
INVx1_ASAP7_75t_L g1284 ( .A(n_221), .Y(n_1284) );
AOI22xp33_ASAP7_75t_L g1294 ( .A1(n_221), .A2(n_291), .B1(n_719), .B2(n_1295), .Y(n_1294) );
INVx1_ASAP7_75t_L g979 ( .A(n_222), .Y(n_979) );
INVx1_ASAP7_75t_L g1175 ( .A(n_223), .Y(n_1175) );
OAI211xp5_ASAP7_75t_L g1187 ( .A1(n_223), .A2(n_686), .B(n_1188), .C(n_1196), .Y(n_1187) );
INVx1_ASAP7_75t_L g1854 ( .A(n_224), .Y(n_1854) );
CKINVDCx5p33_ASAP7_75t_R g847 ( .A(n_225), .Y(n_847) );
INVx1_ASAP7_75t_L g1857 ( .A(n_226), .Y(n_1857) );
CKINVDCx5p33_ASAP7_75t_R g726 ( .A(n_227), .Y(n_726) );
CKINVDCx5p33_ASAP7_75t_R g782 ( .A(n_229), .Y(n_782) );
INVx2_ASAP7_75t_L g424 ( .A(n_230), .Y(n_424) );
NAND2xp5_ASAP7_75t_L g439 ( .A(n_230), .B(n_422), .Y(n_439) );
INVx1_ASAP7_75t_L g484 ( .A(n_230), .Y(n_484) );
INVxp67_ASAP7_75t_L g1831 ( .A(n_231), .Y(n_1831) );
CKINVDCx5p33_ASAP7_75t_R g1197 ( .A(n_232), .Y(n_1197) );
AOI22xp5_ASAP7_75t_L g1607 ( .A1(n_233), .A2(n_362), .B1(n_1587), .B2(n_1590), .Y(n_1607) );
OAI211xp5_ASAP7_75t_L g1252 ( .A1(n_234), .A2(n_686), .B(n_1253), .C(n_1258), .Y(n_1252) );
INVx1_ASAP7_75t_L g860 ( .A(n_235), .Y(n_860) );
NAND2xp33_ASAP7_75t_SL g903 ( .A(n_235), .B(n_520), .Y(n_903) );
INVx1_ASAP7_75t_L g1887 ( .A(n_237), .Y(n_1887) );
AOI22xp33_ASAP7_75t_L g1046 ( .A1(n_238), .A2(n_338), .B1(n_675), .B2(n_989), .Y(n_1046) );
INVx1_ASAP7_75t_L g1063 ( .A(n_238), .Y(n_1063) );
AOI22xp33_ASAP7_75t_SL g1041 ( .A1(n_240), .A2(n_267), .B1(n_463), .B2(n_1042), .Y(n_1041) );
INVxp67_ASAP7_75t_SL g1068 ( .A(n_240), .Y(n_1068) );
INVx1_ASAP7_75t_L g1282 ( .A(n_241), .Y(n_1282) );
INVx1_ASAP7_75t_L g1240 ( .A(n_242), .Y(n_1240) );
OAI22xp5_ASAP7_75t_L g785 ( .A1(n_243), .A2(n_326), .B1(n_776), .B2(n_786), .Y(n_785) );
INVx1_ASAP7_75t_L g816 ( .A(n_243), .Y(n_816) );
INVx1_ASAP7_75t_L g1203 ( .A(n_244), .Y(n_1203) );
INVx1_ASAP7_75t_L g1868 ( .A(n_245), .Y(n_1868) );
INVx1_ASAP7_75t_L g1206 ( .A(n_246), .Y(n_1206) );
AOI21xp5_ASAP7_75t_L g861 ( .A1(n_247), .A2(n_799), .B(n_862), .Y(n_861) );
INVx1_ASAP7_75t_L g907 ( .A(n_248), .Y(n_907) );
OAI21xp5_ASAP7_75t_L g1073 ( .A1(n_249), .A2(n_656), .B(n_1074), .Y(n_1073) );
BUFx3_ASAP7_75t_L g416 ( .A(n_251), .Y(n_416) );
AOI22xp33_ASAP7_75t_L g962 ( .A1(n_252), .A2(n_295), .B1(n_486), .B2(n_963), .Y(n_962) );
AOI221xp5_ASAP7_75t_L g1357 ( .A1(n_253), .A2(n_279), .B1(n_612), .B2(n_613), .C(n_1358), .Y(n_1357) );
INVx1_ASAP7_75t_L g1507 ( .A(n_254), .Y(n_1507) );
INVx1_ASAP7_75t_L g1331 ( .A(n_256), .Y(n_1331) );
CKINVDCx20_ASAP7_75t_R g488 ( .A(n_257), .Y(n_488) );
OAI22xp5_ASAP7_75t_L g1227 ( .A1(n_258), .A2(n_261), .B1(n_490), .B2(n_1228), .Y(n_1227) );
OAI221xp5_ASAP7_75t_L g1249 ( .A1(n_258), .A2(n_261), .B1(n_621), .B2(n_624), .C(n_1250), .Y(n_1249) );
INVx1_ASAP7_75t_L g833 ( .A(n_260), .Y(n_833) );
NOR2xp33_ASAP7_75t_L g835 ( .A(n_260), .B(n_836), .Y(n_835) );
AOI21xp33_ASAP7_75t_L g942 ( .A1(n_263), .A2(n_523), .B(n_768), .Y(n_942) );
INVx1_ASAP7_75t_L g952 ( .A(n_263), .Y(n_952) );
INVx1_ASAP7_75t_L g501 ( .A(n_264), .Y(n_501) );
INVx1_ASAP7_75t_L g1224 ( .A(n_265), .Y(n_1224) );
XOR2x2_ASAP7_75t_L g919 ( .A(n_266), .B(n_920), .Y(n_919) );
AOI21xp33_ASAP7_75t_L g1054 ( .A1(n_267), .A2(n_643), .B(n_773), .Y(n_1054) );
AOI22xp33_ASAP7_75t_L g1546 ( .A1(n_268), .A2(n_283), .B1(n_530), .B2(n_1257), .Y(n_1546) );
OAI22xp33_ASAP7_75t_L g1147 ( .A1(n_270), .A2(n_287), .B1(n_593), .B2(n_599), .Y(n_1147) );
INVx1_ASAP7_75t_L g1158 ( .A(n_270), .Y(n_1158) );
CKINVDCx5p33_ASAP7_75t_R g1386 ( .A(n_271), .Y(n_1386) );
BUFx3_ASAP7_75t_L g401 ( .A(n_272), .Y(n_401) );
INVx1_ASAP7_75t_L g506 ( .A(n_272), .Y(n_506) );
AOI22xp33_ASAP7_75t_L g743 ( .A1(n_273), .A2(n_333), .B1(n_463), .B2(n_744), .Y(n_743) );
INVx1_ASAP7_75t_L g1512 ( .A(n_274), .Y(n_1512) );
AOI22xp33_ASAP7_75t_SL g590 ( .A1(n_275), .A2(n_329), .B1(n_585), .B2(n_588), .Y(n_590) );
XNOR2x1_ASAP7_75t_L g1311 ( .A(n_276), .B(n_1312), .Y(n_1311) );
NAND2xp5_ASAP7_75t_SL g936 ( .A(n_277), .B(n_523), .Y(n_936) );
AOI22xp33_ASAP7_75t_L g1551 ( .A1(n_278), .A2(n_342), .B1(n_530), .B2(n_1361), .Y(n_1551) );
AOI22xp33_ASAP7_75t_SL g1567 ( .A1(n_278), .A2(n_354), .B1(n_469), .B2(n_1091), .Y(n_1567) );
INVx1_ASAP7_75t_L g616 ( .A(n_280), .Y(n_616) );
INVx1_ASAP7_75t_L g856 ( .A(n_282), .Y(n_856) );
INVx1_ASAP7_75t_L g1330 ( .A(n_284), .Y(n_1330) );
INVx1_ASAP7_75t_L g1137 ( .A(n_286), .Y(n_1137) );
INVx1_ASAP7_75t_L g1159 ( .A(n_287), .Y(n_1159) );
INVx1_ASAP7_75t_L g1865 ( .A(n_289), .Y(n_1865) );
INVx1_ASAP7_75t_L g694 ( .A(n_290), .Y(n_694) );
NAND2xp33_ASAP7_75t_SL g1279 ( .A(n_291), .B(n_989), .Y(n_1279) );
NAND2xp5_ASAP7_75t_SL g939 ( .A(n_295), .B(n_519), .Y(n_939) );
AOI22xp33_ASAP7_75t_L g1360 ( .A1(n_297), .A2(n_341), .B1(n_530), .B2(n_1361), .Y(n_1360) );
XNOR2x2_ASAP7_75t_L g1131 ( .A(n_298), .B(n_1132), .Y(n_1131) );
AOI22xp33_ASAP7_75t_SL g790 ( .A1(n_299), .A2(n_373), .B1(n_463), .B2(n_671), .Y(n_790) );
INVx1_ASAP7_75t_L g1246 ( .A(n_300), .Y(n_1246) );
INVx1_ASAP7_75t_L g419 ( .A(n_301), .Y(n_419) );
INVx1_ASAP7_75t_L g436 ( .A(n_301), .Y(n_436) );
INVx1_ASAP7_75t_L g1303 ( .A(n_305), .Y(n_1303) );
AOI221xp5_ASAP7_75t_L g609 ( .A1(n_307), .A2(n_335), .B1(n_522), .B2(n_610), .C(n_613), .Y(n_609) );
AOI22xp33_ASAP7_75t_L g614 ( .A1(n_308), .A2(n_329), .B1(n_527), .B2(n_529), .Y(n_614) );
INVx1_ASAP7_75t_L g1212 ( .A(n_311), .Y(n_1212) );
OAI21xp33_ASAP7_75t_L g945 ( .A1(n_312), .A2(n_805), .B(n_946), .Y(n_945) );
INVx1_ASAP7_75t_L g1039 ( .A(n_313), .Y(n_1039) );
AOI22xp5_ASAP7_75t_SL g1610 ( .A1(n_314), .A2(n_370), .B1(n_1580), .B2(n_1606), .Y(n_1610) );
INVxp33_ASAP7_75t_L g1825 ( .A(n_315), .Y(n_1825) );
CKINVDCx5p33_ASAP7_75t_R g831 ( .A(n_316), .Y(n_831) );
CKINVDCx5p33_ASAP7_75t_R g1318 ( .A(n_317), .Y(n_1318) );
INVx1_ASAP7_75t_L g1832 ( .A(n_318), .Y(n_1832) );
AOI221xp5_ASAP7_75t_SL g771 ( .A1(n_319), .A2(n_373), .B1(n_520), .B2(n_772), .C(n_773), .Y(n_771) );
INVx1_ASAP7_75t_L g679 ( .A(n_320), .Y(n_679) );
AND2x2_ASAP7_75t_L g1582 ( .A(n_321), .B(n_1583), .Y(n_1582) );
INVx1_ASAP7_75t_L g1589 ( .A(n_321), .Y(n_1589) );
INVx1_ASAP7_75t_L g1502 ( .A(n_323), .Y(n_1502) );
INVx1_ASAP7_75t_L g1260 ( .A(n_324), .Y(n_1260) );
INVx1_ASAP7_75t_L g802 ( .A(n_326), .Y(n_802) );
INVx1_ASAP7_75t_L g1526 ( .A(n_328), .Y(n_1526) );
INVx1_ASAP7_75t_L g1364 ( .A(n_330), .Y(n_1364) );
INVxp67_ASAP7_75t_SL g1889 ( .A(n_331), .Y(n_1889) );
CKINVDCx16_ASAP7_75t_R g867 ( .A(n_332), .Y(n_867) );
CKINVDCx5p33_ASAP7_75t_R g1402 ( .A(n_336), .Y(n_1402) );
AOI22xp5_ASAP7_75t_L g1055 ( .A1(n_338), .A2(n_365), .B1(n_530), .B2(n_938), .Y(n_1055) );
NAND2xp5_ASAP7_75t_L g1164 ( .A(n_339), .B(n_1070), .Y(n_1164) );
OAI21xp33_ASAP7_75t_L g997 ( .A1(n_340), .A2(n_558), .B(n_998), .Y(n_997) );
OAI21xp5_ASAP7_75t_SL g1338 ( .A1(n_343), .A2(n_656), .B(n_1339), .Y(n_1338) );
CKINVDCx5p33_ASAP7_75t_R g1388 ( .A(n_344), .Y(n_1388) );
INVx1_ASAP7_75t_L g1809 ( .A(n_345), .Y(n_1809) );
INVxp67_ASAP7_75t_SL g1071 ( .A(n_346), .Y(n_1071) );
CKINVDCx5p33_ASAP7_75t_R g1130 ( .A(n_347), .Y(n_1130) );
OAI211xp5_ASAP7_75t_L g1490 ( .A1(n_348), .A2(n_1014), .B(n_1060), .C(n_1491), .Y(n_1490) );
INVx1_ASAP7_75t_L g1533 ( .A(n_348), .Y(n_1533) );
CKINVDCx5p33_ASAP7_75t_R g448 ( .A(n_349), .Y(n_448) );
AOI221xp5_ASAP7_75t_L g1498 ( .A1(n_350), .A2(n_367), .B1(n_612), .B2(n_644), .C(n_716), .Y(n_1498) );
INVx1_ASAP7_75t_L g1510 ( .A(n_350), .Y(n_1510) );
BUFx6f_ASAP7_75t_L g397 ( .A(n_351), .Y(n_397) );
INVx1_ASAP7_75t_L g742 ( .A(n_353), .Y(n_742) );
INVxp67_ASAP7_75t_SL g1544 ( .A(n_354), .Y(n_1544) );
NOR2xp33_ASAP7_75t_R g892 ( .A(n_355), .B(n_893), .Y(n_892) );
INVx1_ASAP7_75t_L g827 ( .A(n_356), .Y(n_827) );
INVx1_ASAP7_75t_L g578 ( .A(n_357), .Y(n_578) );
OAI221xp5_ASAP7_75t_SL g620 ( .A1(n_357), .A2(n_374), .B1(n_621), .B2(n_624), .C(n_629), .Y(n_620) );
INVx1_ASAP7_75t_L g748 ( .A(n_359), .Y(n_748) );
XNOR2xp5_ASAP7_75t_L g1850 ( .A(n_361), .B(n_1851), .Y(n_1850) );
INVx1_ASAP7_75t_L g428 ( .A(n_364), .Y(n_428) );
INVx1_ASAP7_75t_L g442 ( .A(n_364), .Y(n_442) );
INVx2_ASAP7_75t_L g461 ( .A(n_364), .Y(n_461) );
CKINVDCx5p33_ASAP7_75t_R g1262 ( .A(n_366), .Y(n_1262) );
INVxp67_ASAP7_75t_SL g1522 ( .A(n_367), .Y(n_1522) );
CKINVDCx5p33_ASAP7_75t_R g1800 ( .A(n_368), .Y(n_1800) );
OAI22xp33_ASAP7_75t_SL g681 ( .A1(n_369), .A2(n_371), .B1(n_490), .B2(n_682), .Y(n_681) );
OAI221xp5_ASAP7_75t_L g696 ( .A1(n_369), .A2(n_371), .B1(n_621), .B2(n_625), .C(n_697), .Y(n_696) );
XNOR2xp5_ASAP7_75t_L g651 ( .A(n_370), .B(n_652), .Y(n_651) );
INVx1_ASAP7_75t_L g1171 ( .A(n_372), .Y(n_1171) );
INVx1_ASAP7_75t_L g580 ( .A(n_374), .Y(n_580) );
AOI21xp5_ASAP7_75t_L g375 ( .A1(n_376), .A2(n_402), .B(n_1574), .Y(n_375) );
INVx2_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
INVx1_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
BUFx4f_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
INVx3_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
OR2x2_ASAP7_75t_L g380 ( .A(n_381), .B(n_387), .Y(n_380) );
NOR2xp33_ASAP7_75t_L g1844 ( .A(n_381), .B(n_390), .Y(n_1844) );
INVx1_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
NOR2xp33_ASAP7_75t_L g382 ( .A(n_383), .B(n_385), .Y(n_382) );
NOR2xp33_ASAP7_75t_L g1848 ( .A(n_383), .B(n_386), .Y(n_1848) );
INVx1_ASAP7_75t_L g1894 ( .A(n_383), .Y(n_1894) );
HB1xp67_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
INVx1_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
NOR2xp33_ASAP7_75t_L g1896 ( .A(n_386), .B(n_1894), .Y(n_1896) );
INVx1_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
NAND2xp5_ASAP7_75t_L g388 ( .A(n_389), .B(n_392), .Y(n_388) );
INVx1_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
AND2x4_ASAP7_75t_L g1449 ( .A(n_390), .B(n_1450), .Y(n_1449) );
INVx1_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
AND2x4_ASAP7_75t_L g525 ( .A(n_391), .B(n_401), .Y(n_525) );
AND2x4_ASAP7_75t_L g547 ( .A(n_391), .B(n_400), .Y(n_547) );
INVx1_ASAP7_75t_L g1445 ( .A(n_392), .Y(n_1445) );
AND2x4_ASAP7_75t_SL g1843 ( .A(n_392), .B(n_1844), .Y(n_1843) );
INVx3_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
OR2x6_ASAP7_75t_L g393 ( .A(n_394), .B(n_399), .Y(n_393) );
INVxp67_ASAP7_75t_L g1070 ( .A(n_394), .Y(n_1070) );
OR2x6_ASAP7_75t_L g1437 ( .A(n_394), .B(n_1438), .Y(n_1437) );
INVx2_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
BUFx4f_ASAP7_75t_L g632 ( .A(n_395), .Y(n_632) );
INVx3_ASAP7_75t_L g1208 ( .A(n_395), .Y(n_1208) );
INVx3_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
OR2x2_ASAP7_75t_L g396 ( .A(n_397), .B(n_398), .Y(n_396) );
INVx2_ASAP7_75t_L g446 ( .A(n_397), .Y(n_446) );
AND2x2_ASAP7_75t_L g511 ( .A(n_397), .B(n_512), .Y(n_511) );
INVx2_ASAP7_75t_L g517 ( .A(n_397), .Y(n_517) );
AND2x2_ASAP7_75t_L g521 ( .A(n_397), .B(n_398), .Y(n_521) );
INVx1_ASAP7_75t_L g562 ( .A(n_397), .Y(n_562) );
NAND2x1_ASAP7_75t_L g701 ( .A(n_397), .B(n_398), .Y(n_701) );
INVx1_ASAP7_75t_L g447 ( .A(n_398), .Y(n_447) );
INVx2_ASAP7_75t_L g512 ( .A(n_398), .Y(n_512) );
AND2x2_ASAP7_75t_L g516 ( .A(n_398), .B(n_517), .Y(n_516) );
BUFx2_ASAP7_75t_L g552 ( .A(n_398), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g637 ( .A(n_398), .B(n_517), .Y(n_637) );
OR2x2_ASAP7_75t_L g901 ( .A(n_398), .B(n_446), .Y(n_901) );
INVxp67_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
INVx1_ASAP7_75t_L g1425 ( .A(n_400), .Y(n_1425) );
INVx2_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
BUFx2_ASAP7_75t_L g1429 ( .A(n_401), .Y(n_1429) );
AND2x4_ASAP7_75t_L g1433 ( .A(n_401), .B(n_561), .Y(n_1433) );
XNOR2xp5_ASAP7_75t_L g402 ( .A(n_403), .B(n_1079), .Y(n_402) );
AO22x2_ASAP7_75t_L g403 ( .A1(n_404), .A2(n_405), .B1(n_1031), .B2(n_1078), .Y(n_403) );
INVx1_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
AO22x2_ASAP7_75t_L g405 ( .A1(n_406), .A2(n_752), .B1(n_753), .B2(n_1030), .Y(n_405) );
INVx1_ASAP7_75t_L g1030 ( .A(n_406), .Y(n_1030) );
XNOR2xp5_ASAP7_75t_L g406 ( .A(n_407), .B(n_649), .Y(n_406) );
XOR2xp5_ASAP7_75t_L g407 ( .A(n_408), .B(n_573), .Y(n_407) );
XNOR2xp5_ASAP7_75t_L g408 ( .A(n_409), .B(n_572), .Y(n_408) );
AND2x2_ASAP7_75t_L g409 ( .A(n_410), .B(n_498), .Y(n_409) );
AOI221xp5_ASAP7_75t_L g410 ( .A1(n_411), .A2(n_429), .B1(n_430), .B2(n_448), .C(n_449), .Y(n_410) );
NAND2xp5_ASAP7_75t_L g1099 ( .A(n_411), .B(n_1100), .Y(n_1099) );
AOI22xp5_ASAP7_75t_L g1269 ( .A1(n_411), .A2(n_1270), .B1(n_1271), .B2(n_1272), .Y(n_1269) );
AOI221xp5_ASAP7_75t_L g1313 ( .A1(n_411), .A2(n_430), .B1(n_1314), .B2(n_1315), .C(n_1316), .Y(n_1313) );
AOI221xp5_ASAP7_75t_L g1835 ( .A1(n_411), .A2(n_430), .B1(n_1817), .B2(n_1836), .C(n_1837), .Y(n_1835) );
NAND2xp5_ASAP7_75t_L g1856 ( .A(n_411), .B(n_1857), .Y(n_1856) );
INVx3_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
INVx5_ASAP7_75t_L g970 ( .A(n_412), .Y(n_970) );
OR2x6_ASAP7_75t_L g412 ( .A(n_413), .B(n_425), .Y(n_412) );
OR2x2_ASAP7_75t_L g604 ( .A(n_413), .B(n_425), .Y(n_604) );
NAND2x1p5_ASAP7_75t_L g413 ( .A(n_414), .B(n_420), .Y(n_413) );
INVx8_ASAP7_75t_L g464 ( .A(n_414), .Y(n_464) );
BUFx3_ASAP7_75t_L g862 ( .A(n_414), .Y(n_862) );
BUFx3_ASAP7_75t_L g956 ( .A(n_414), .Y(n_956) );
HB1xp67_ASAP7_75t_L g963 ( .A(n_414), .Y(n_963) );
AND2x4_ASAP7_75t_L g414 ( .A(n_415), .B(n_417), .Y(n_414) );
AND2x4_ASAP7_75t_L g470 ( .A(n_415), .B(n_471), .Y(n_470) );
INVx2_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
NAND2xp5_ASAP7_75t_L g435 ( .A(n_416), .B(n_436), .Y(n_435) );
AND2x4_ASAP7_75t_L g453 ( .A(n_416), .B(n_454), .Y(n_453) );
BUFx6f_ASAP7_75t_L g475 ( .A(n_416), .Y(n_475) );
OR2x2_ASAP7_75t_L g596 ( .A(n_416), .B(n_418), .Y(n_596) );
INVx1_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
INVx1_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
INVxp67_ASAP7_75t_L g471 ( .A(n_419), .Y(n_471) );
AND2x4_ASAP7_75t_L g455 ( .A(n_420), .B(n_441), .Y(n_455) );
INVx1_ASAP7_75t_L g864 ( .A(n_420), .Y(n_864) );
AND2x6_ASAP7_75t_L g871 ( .A(n_420), .B(n_491), .Y(n_871) );
AND2x2_ASAP7_75t_L g873 ( .A(n_420), .B(n_497), .Y(n_873) );
AND2x4_ASAP7_75t_L g420 ( .A(n_421), .B(n_423), .Y(n_420) );
NAND3x1_ASAP7_75t_L g482 ( .A(n_421), .B(n_483), .C(n_484), .Y(n_482) );
NAND2x1p5_ASAP7_75t_L g799 ( .A(n_421), .B(n_484), .Y(n_799) );
OR2x4_ASAP7_75t_L g1455 ( .A(n_421), .B(n_596), .Y(n_1455) );
INVx1_ASAP7_75t_L g1458 ( .A(n_421), .Y(n_1458) );
AND2x4_ASAP7_75t_L g1463 ( .A(n_421), .B(n_453), .Y(n_1463) );
OR2x6_ASAP7_75t_L g1478 ( .A(n_421), .B(n_668), .Y(n_1478) );
INVx3_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
BUFx3_ASAP7_75t_L g459 ( .A(n_422), .Y(n_459) );
NAND2xp33_ASAP7_75t_SL g662 ( .A(n_422), .B(n_424), .Y(n_662) );
INVx1_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
AND3x4_ASAP7_75t_L g458 ( .A(n_424), .B(n_459), .C(n_460), .Y(n_458) );
AND2x2_ASAP7_75t_L g851 ( .A(n_424), .B(n_459), .Y(n_851) );
HB1xp67_ASAP7_75t_L g1481 ( .A(n_424), .Y(n_1481) );
INVxp67_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
OR2x2_ASAP7_75t_L g559 ( .A(n_426), .B(n_560), .Y(n_559) );
INVx1_ASAP7_75t_L g810 ( .A(n_426), .Y(n_810) );
OR2x2_ASAP7_75t_L g884 ( .A(n_426), .B(n_560), .Y(n_884) );
INVx1_ASAP7_75t_L g1450 ( .A(n_426), .Y(n_1450) );
BUFx2_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
INVx2_ASAP7_75t_L g438 ( .A(n_427), .Y(n_438) );
INVx1_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
AOI221xp5_ASAP7_75t_L g513 ( .A1(n_429), .A2(n_514), .B1(n_518), .B2(n_526), .C(n_531), .Y(n_513) );
AOI21xp5_ASAP7_75t_L g601 ( .A1(n_430), .A2(n_602), .B(n_603), .Y(n_601) );
AOI21xp5_ASAP7_75t_L g653 ( .A1(n_430), .A2(n_654), .B(n_655), .Y(n_653) );
AOI21xp5_ASAP7_75t_L g747 ( .A1(n_430), .A2(n_748), .B(n_749), .Y(n_747) );
AOI211x1_ASAP7_75t_L g973 ( .A1(n_430), .A2(n_974), .B(n_975), .C(n_997), .Y(n_973) );
NAND2xp5_ASAP7_75t_L g1075 ( .A(n_430), .B(n_1076), .Y(n_1075) );
NAND2xp5_ASAP7_75t_L g1129 ( .A(n_430), .B(n_1130), .Y(n_1129) );
AOI21xp5_ASAP7_75t_L g1148 ( .A1(n_430), .A2(n_1149), .B(n_1150), .Y(n_1148) );
NAND2xp5_ASAP7_75t_L g1216 ( .A(n_430), .B(n_1217), .Y(n_1216) );
AOI21xp33_ASAP7_75t_L g1261 ( .A1(n_430), .A2(n_1262), .B(n_1263), .Y(n_1261) );
AOI21xp33_ASAP7_75t_L g1365 ( .A1(n_430), .A2(n_1366), .B(n_1367), .Y(n_1365) );
AOI21xp5_ASAP7_75t_L g1555 ( .A1(n_430), .A2(n_1556), .B(n_1557), .Y(n_1555) );
INVx8_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
AND2x4_ASAP7_75t_L g431 ( .A(n_432), .B(n_440), .Y(n_431) );
INVx1_ASAP7_75t_L g817 ( .A(n_432), .Y(n_817) );
OR2x2_ASAP7_75t_L g432 ( .A(n_433), .B(n_437), .Y(n_432) );
BUFx3_ASAP7_75t_L g960 ( .A(n_433), .Y(n_960) );
INVx1_ASAP7_75t_L g1514 ( .A(n_433), .Y(n_1514) );
INVx1_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
BUFx6f_ASAP7_75t_L g678 ( .A(n_434), .Y(n_678) );
INVx1_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
BUFx2_ASAP7_75t_L g668 ( .A(n_435), .Y(n_668) );
INVx2_ASAP7_75t_L g454 ( .A(n_436), .Y(n_454) );
INVx1_ASAP7_75t_L g566 ( .A(n_436), .Y(n_566) );
OR2x2_ASAP7_75t_L g563 ( .A(n_437), .B(n_564), .Y(n_563) );
INVx1_ASAP7_75t_L g570 ( .A(n_437), .Y(n_570) );
INVx1_ASAP7_75t_L g598 ( .A(n_437), .Y(n_598) );
OR2x2_ASAP7_75t_L g437 ( .A(n_438), .B(n_439), .Y(n_437) );
OR2x2_ASAP7_75t_L g661 ( .A(n_438), .B(n_662), .Y(n_661) );
AND2x2_ASAP7_75t_SL g897 ( .A(n_438), .B(n_525), .Y(n_897) );
INVx1_ASAP7_75t_L g1420 ( .A(n_438), .Y(n_1420) );
HB1xp67_ASAP7_75t_L g1483 ( .A(n_438), .Y(n_1483) );
INVx1_ASAP7_75t_L g838 ( .A(n_439), .Y(n_838) );
NAND2xp5_ASAP7_75t_L g914 ( .A(n_440), .B(n_915), .Y(n_914) );
OR2x2_ASAP7_75t_L g440 ( .A(n_441), .B(n_443), .Y(n_440) );
INVx1_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
INVx1_ASAP7_75t_L g483 ( .A(n_442), .Y(n_483) );
NAND2xp5_ASAP7_75t_L g894 ( .A(n_442), .B(n_505), .Y(n_894) );
NAND2xp5_ASAP7_75t_L g443 ( .A(n_444), .B(n_445), .Y(n_443) );
AND2x6_ASAP7_75t_L g531 ( .A(n_444), .B(n_520), .Y(n_531) );
AND2x2_ASAP7_75t_L g550 ( .A(n_444), .B(n_551), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g560 ( .A(n_444), .B(n_561), .Y(n_560) );
INVx1_ASAP7_75t_L g628 ( .A(n_444), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g889 ( .A(n_444), .B(n_461), .Y(n_889) );
AND2x2_ASAP7_75t_L g504 ( .A(n_445), .B(n_505), .Y(n_504) );
INVx3_ASAP7_75t_L g528 ( .A(n_445), .Y(n_528) );
BUFx6f_ASAP7_75t_L g692 ( .A(n_445), .Y(n_692) );
AND2x2_ASAP7_75t_L g445 ( .A(n_446), .B(n_447), .Y(n_445) );
HB1xp67_ASAP7_75t_L g781 ( .A(n_446), .Y(n_781) );
NAND3xp33_ASAP7_75t_SL g449 ( .A(n_450), .B(n_456), .C(n_487), .Y(n_449) );
INVx2_ASAP7_75t_SL g600 ( .A(n_450), .Y(n_600) );
AND5x1_ASAP7_75t_L g920 ( .A(n_450), .B(n_921), .C(n_948), .D(n_964), .E(n_968), .Y(n_920) );
AND4x1_ASAP7_75t_L g1169 ( .A(n_450), .B(n_1170), .C(n_1174), .D(n_1176), .Y(n_1169) );
NAND3xp33_ASAP7_75t_SL g1316 ( .A(n_450), .B(n_1317), .C(n_1320), .Y(n_1316) );
NAND5xp2_ASAP7_75t_L g1852 ( .A(n_450), .B(n_1853), .C(n_1856), .D(n_1858), .E(n_1859), .Y(n_1852) );
INVx3_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
HB1xp67_ASAP7_75t_L g658 ( .A(n_451), .Y(n_658) );
NOR3xp33_ASAP7_75t_L g733 ( .A(n_451), .B(n_734), .C(n_746), .Y(n_733) );
AOI221xp5_ASAP7_75t_L g800 ( .A1(n_451), .A2(n_683), .B1(n_779), .B2(n_801), .C(n_802), .Y(n_800) );
INVx3_ASAP7_75t_L g983 ( .A(n_451), .Y(n_983) );
NOR3xp33_ASAP7_75t_SL g1273 ( .A(n_451), .B(n_1274), .C(n_1287), .Y(n_1273) );
NOR3xp33_ASAP7_75t_L g1558 ( .A(n_451), .B(n_1559), .C(n_1568), .Y(n_1558) );
AND2x4_ASAP7_75t_L g451 ( .A(n_452), .B(n_455), .Y(n_451) );
BUFx2_ASAP7_75t_L g583 ( .A(n_452), .Y(n_583) );
BUFx2_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
BUFx2_ASAP7_75t_L g465 ( .A(n_453), .Y(n_465) );
BUFx3_ASAP7_75t_L g486 ( .A(n_453), .Y(n_486) );
BUFx2_ASAP7_75t_L g671 ( .A(n_453), .Y(n_671) );
INVx2_ASAP7_75t_L g745 ( .A(n_453), .Y(n_745) );
BUFx2_ASAP7_75t_L g1834 ( .A(n_453), .Y(n_1834) );
INVx1_ASAP7_75t_L g476 ( .A(n_454), .Y(n_476) );
NAND2x1_ASAP7_75t_L g490 ( .A(n_455), .B(n_491), .Y(n_490) );
AND2x4_ASAP7_75t_L g494 ( .A(n_455), .B(n_495), .Y(n_494) );
AND2x2_ASAP7_75t_L g579 ( .A(n_455), .B(n_491), .Y(n_579) );
AND2x4_ASAP7_75t_SL g683 ( .A(n_455), .B(n_495), .Y(n_683) );
AND2x4_ASAP7_75t_SL g801 ( .A(n_455), .B(n_491), .Y(n_801) );
AND2x2_ASAP7_75t_L g1289 ( .A(n_455), .B(n_491), .Y(n_1289) );
AOI33xp33_ASAP7_75t_L g456 ( .A1(n_457), .A2(n_462), .A3(n_466), .B1(n_477), .B2(n_479), .B3(n_485), .Y(n_456) );
AOI33xp33_ASAP7_75t_L g581 ( .A1(n_457), .A2(n_479), .A3(n_582), .B1(n_584), .B2(n_590), .B3(n_591), .Y(n_581) );
AOI33xp33_ASAP7_75t_L g984 ( .A1(n_457), .A2(n_985), .A3(n_988), .B1(n_990), .B2(n_991), .B3(n_993), .Y(n_984) );
NAND2xp5_ASAP7_75t_L g1092 ( .A(n_457), .B(n_1093), .Y(n_1092) );
AOI33xp33_ASAP7_75t_L g1138 ( .A1(n_457), .A2(n_1139), .A3(n_1140), .B1(n_1143), .B2(n_1145), .B3(n_1146), .Y(n_1138) );
AOI33xp33_ASAP7_75t_L g1176 ( .A1(n_457), .A2(n_1177), .A3(n_1178), .B1(n_1182), .B2(n_1183), .B3(n_1185), .Y(n_1176) );
BUFx3_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
AOI33xp33_ASAP7_75t_L g789 ( .A1(n_458), .A2(n_790), .A3(n_791), .B1(n_793), .B2(n_795), .B3(n_797), .Y(n_789) );
AOI33xp33_ASAP7_75t_L g1040 ( .A1(n_458), .A2(n_1041), .A3(n_1043), .B1(n_1046), .B2(n_1047), .B3(n_1048), .Y(n_1040) );
INVx1_ASAP7_75t_L g1325 ( .A(n_458), .Y(n_1325) );
AOI33xp33_ASAP7_75t_L g1372 ( .A1(n_458), .A2(n_1373), .A3(n_1374), .B1(n_1375), .B2(n_1376), .B3(n_1377), .Y(n_1372) );
AOI33xp33_ASAP7_75t_L g1562 ( .A1(n_458), .A2(n_1376), .A3(n_1563), .B1(n_1565), .B2(n_1566), .B3(n_1567), .Y(n_1562) );
INVx3_ASAP7_75t_L g1467 ( .A(n_459), .Y(n_1467) );
INVx1_ASAP7_75t_L g648 ( .A(n_460), .Y(n_648) );
OAI31xp33_ASAP7_75t_L g834 ( .A1(n_460), .A2(n_835), .A3(n_839), .B(n_865), .Y(n_834) );
INVx2_ASAP7_75t_SL g1126 ( .A(n_460), .Y(n_1126) );
INVx2_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
BUFx2_ASAP7_75t_L g556 ( .A(n_461), .Y(n_556) );
BUFx2_ASAP7_75t_L g1184 ( .A(n_463), .Y(n_1184) );
INVx8_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
INVx2_ASAP7_75t_L g569 ( .A(n_464), .Y(n_569) );
INVx3_ASAP7_75t_L g994 ( .A(n_464), .Y(n_994) );
INVx2_ASAP7_75t_L g1286 ( .A(n_464), .Y(n_1286) );
INVx1_ASAP7_75t_L g996 ( .A(n_465), .Y(n_996) );
INVx1_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
OAI22xp5_ASAP7_75t_L g1241 ( .A1(n_468), .A2(n_855), .B1(n_1242), .B2(n_1243), .Y(n_1241) );
INVx2_ASAP7_75t_SL g468 ( .A(n_469), .Y(n_468) );
AND2x4_ASAP7_75t_L g571 ( .A(n_469), .B(n_570), .Y(n_571) );
INVx2_ASAP7_75t_SL g737 ( .A(n_469), .Y(n_737) );
HB1xp67_ASAP7_75t_L g1090 ( .A(n_469), .Y(n_1090) );
INVx3_ASAP7_75t_L g1511 ( .A(n_469), .Y(n_1511) );
BUFx8_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
INVx2_ASAP7_75t_L g587 ( .A(n_470), .Y(n_587) );
BUFx6f_ASAP7_75t_L g675 ( .A(n_470), .Y(n_675) );
BUFx6f_ASAP7_75t_L g849 ( .A(n_470), .Y(n_849) );
INVx1_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
INVx2_ASAP7_75t_L g989 ( .A(n_473), .Y(n_989) );
INVx2_ASAP7_75t_R g1045 ( .A(n_473), .Y(n_1045) );
INVx5_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
BUFx3_ASAP7_75t_L g478 ( .A(n_474), .Y(n_478) );
BUFx12f_ASAP7_75t_L g589 ( .A(n_474), .Y(n_589) );
AND2x4_ASAP7_75t_L g916 ( .A(n_474), .B(n_838), .Y(n_916) );
BUFx3_ASAP7_75t_L g1091 ( .A(n_474), .Y(n_1091) );
AND2x4_ASAP7_75t_L g474 ( .A(n_475), .B(n_476), .Y(n_474) );
INVx2_ASAP7_75t_L g492 ( .A(n_475), .Y(n_492) );
NAND2x1p5_ASAP7_75t_L g565 ( .A(n_475), .B(n_566), .Y(n_565) );
BUFx2_ASAP7_75t_L g1468 ( .A(n_475), .Y(n_1468) );
INVx1_ASAP7_75t_L g497 ( .A(n_476), .Y(n_497) );
INVx1_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
OAI22xp5_ASAP7_75t_SL g734 ( .A1(n_480), .A2(n_735), .B1(n_736), .B2(n_741), .Y(n_734) );
CKINVDCx5p33_ASAP7_75t_R g480 ( .A(n_481), .Y(n_480) );
INVx2_ASAP7_75t_L g672 ( .A(n_481), .Y(n_672) );
INVx2_ASAP7_75t_L g957 ( .A(n_481), .Y(n_957) );
INVx3_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
INVx3_ASAP7_75t_L g992 ( .A(n_482), .Y(n_992) );
AOI22xp33_ASAP7_75t_L g487 ( .A1(n_488), .A2(n_489), .B1(n_493), .B2(n_494), .Y(n_487) );
AOI222xp33_ASAP7_75t_L g532 ( .A1(n_488), .A2(n_493), .B1(n_533), .B2(n_535), .C1(n_537), .C2(n_548), .Y(n_532) );
AOI221x1_ASAP7_75t_L g948 ( .A1(n_489), .A2(n_494), .B1(n_924), .B2(n_930), .C(n_949), .Y(n_948) );
AOI22xp33_ASAP7_75t_L g1170 ( .A1(n_489), .A2(n_1171), .B1(n_1172), .B2(n_1173), .Y(n_1170) );
AOI22xp33_ASAP7_75t_L g1532 ( .A1(n_489), .A2(n_494), .B1(n_1499), .B2(n_1533), .Y(n_1532) );
AOI22xp33_ASAP7_75t_L g1838 ( .A1(n_489), .A2(n_494), .B1(n_1806), .B2(n_1809), .Y(n_1838) );
INVx2_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
INVx3_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
AOI22xp33_ASAP7_75t_L g577 ( .A1(n_494), .A2(n_578), .B1(n_579), .B2(n_580), .Y(n_577) );
AO22x1_ASAP7_75t_L g977 ( .A1(n_494), .A2(n_579), .B1(n_978), .B2(n_979), .Y(n_977) );
AOI22xp33_ASAP7_75t_L g1101 ( .A1(n_494), .A2(n_579), .B1(n_1102), .B2(n_1103), .Y(n_1101) );
AOI22xp33_ASAP7_75t_L g1135 ( .A1(n_494), .A2(n_579), .B1(n_1136), .B2(n_1137), .Y(n_1135) );
HB1xp67_ASAP7_75t_L g1173 ( .A(n_494), .Y(n_1173) );
AOI22xp33_ASAP7_75t_L g1853 ( .A1(n_494), .A2(n_579), .B1(n_1854), .B2(n_1855), .Y(n_1853) );
INVx2_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
INVx1_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
AOI21xp5_ASAP7_75t_L g498 ( .A1(n_499), .A2(n_553), .B(n_557), .Y(n_498) );
NAND3xp33_ASAP7_75t_L g499 ( .A(n_500), .B(n_513), .C(n_532), .Y(n_499) );
AOI22xp33_ASAP7_75t_L g500 ( .A1(n_501), .A2(n_502), .B1(n_507), .B2(n_508), .Y(n_500) );
AOI22xp33_ASAP7_75t_L g567 ( .A1(n_501), .A2(n_507), .B1(n_568), .B2(n_571), .Y(n_567) );
AOI22xp33_ASAP7_75t_L g615 ( .A1(n_502), .A2(n_616), .B1(n_617), .B2(n_618), .Y(n_615) );
HB1xp67_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
AOI22xp33_ASAP7_75t_L g693 ( .A1(n_503), .A2(n_509), .B1(n_694), .B2(n_695), .Y(n_693) );
AOI22xp5_ASAP7_75t_L g1056 ( .A1(n_503), .A2(n_509), .B1(n_1057), .B2(n_1058), .Y(n_1056) );
AOI22xp33_ASAP7_75t_L g1106 ( .A1(n_503), .A2(n_509), .B1(n_1107), .B2(n_1108), .Y(n_1106) );
AOI22xp5_ASAP7_75t_L g1296 ( .A1(n_503), .A2(n_509), .B1(n_1297), .B2(n_1298), .Y(n_1296) );
AOI22xp5_ASAP7_75t_L g1329 ( .A1(n_503), .A2(n_509), .B1(n_1330), .B2(n_1331), .Y(n_1329) );
AOI22xp33_ASAP7_75t_L g1362 ( .A1(n_503), .A2(n_508), .B1(n_1363), .B2(n_1364), .Y(n_1362) );
NAND2xp5_ASAP7_75t_L g1503 ( .A(n_503), .B(n_1504), .Y(n_1503) );
INVx1_ASAP7_75t_L g1878 ( .A(n_503), .Y(n_1878) );
BUFx6f_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
AOI22xp33_ASAP7_75t_L g720 ( .A1(n_504), .A2(n_509), .B1(n_721), .B2(n_722), .Y(n_720) );
AND2x4_ASAP7_75t_L g832 ( .A(n_504), .B(n_810), .Y(n_832) );
INVx1_ASAP7_75t_L g1005 ( .A(n_504), .Y(n_1005) );
AND2x4_ASAP7_75t_L g509 ( .A(n_505), .B(n_510), .Y(n_509) );
AND2x4_ASAP7_75t_L g514 ( .A(n_505), .B(n_515), .Y(n_514) );
AND2x4_ASAP7_75t_SL g534 ( .A(n_505), .B(n_520), .Y(n_534) );
AND2x2_ASAP7_75t_L g761 ( .A(n_505), .B(n_762), .Y(n_761) );
BUFx2_ASAP7_75t_L g784 ( .A(n_505), .Y(n_784) );
AND2x2_ASAP7_75t_L g811 ( .A(n_505), .B(n_510), .Y(n_811) );
HB1xp67_ASAP7_75t_L g1438 ( .A(n_506), .Y(n_1438) );
AOI22xp33_ASAP7_75t_L g1552 ( .A1(n_508), .A2(n_1004), .B1(n_1553), .B2(n_1554), .Y(n_1552) );
AOI22xp33_ASAP7_75t_SL g1815 ( .A1(n_508), .A2(n_514), .B1(n_1816), .B2(n_1817), .Y(n_1815) );
INVxp67_ASAP7_75t_SL g1871 ( .A(n_508), .Y(n_1871) );
BUFx6f_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
INVx1_ASAP7_75t_L g619 ( .A(n_509), .Y(n_619) );
AOI22xp33_ASAP7_75t_L g1003 ( .A1(n_509), .A2(n_999), .B1(n_1000), .B2(n_1004), .Y(n_1003) );
HB1xp67_ASAP7_75t_L g1198 ( .A(n_509), .Y(n_1198) );
AOI22xp33_ASAP7_75t_L g1500 ( .A1(n_509), .A2(n_761), .B1(n_1501), .B2(n_1502), .Y(n_1500) );
INVx2_ASAP7_75t_L g545 ( .A(n_510), .Y(n_545) );
BUFx6f_ASAP7_75t_L g643 ( .A(n_510), .Y(n_643) );
INVx1_ASAP7_75t_L g717 ( .A(n_510), .Y(n_717) );
BUFx6f_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
BUFx3_ASAP7_75t_L g523 ( .A(n_511), .Y(n_523) );
INVx2_ASAP7_75t_L g767 ( .A(n_511), .Y(n_767) );
AND2x4_ASAP7_75t_L g1447 ( .A(n_511), .B(n_1438), .Y(n_1447) );
INVx3_ASAP7_75t_L g607 ( .A(n_514), .Y(n_607) );
INVx2_ASAP7_75t_SL g686 ( .A(n_514), .Y(n_686) );
NAND2xp5_ASAP7_75t_R g1012 ( .A(n_514), .B(n_982), .Y(n_1012) );
NAND2xp5_ASAP7_75t_L g1059 ( .A(n_514), .B(n_1039), .Y(n_1059) );
AOI221xp5_ASAP7_75t_SL g1109 ( .A1(n_514), .A2(n_531), .B1(n_1100), .B2(n_1110), .C(n_1114), .Y(n_1109) );
BUFx2_ASAP7_75t_L g1115 ( .A(n_515), .Y(n_1115) );
INVx1_ASAP7_75t_L g1195 ( .A(n_515), .Y(n_1195) );
BUFx6f_ASAP7_75t_L g515 ( .A(n_516), .Y(n_515) );
BUFx3_ASAP7_75t_L g530 ( .A(n_516), .Y(n_530) );
INVx2_ASAP7_75t_L g706 ( .A(n_516), .Y(n_706) );
BUFx3_ASAP7_75t_L g719 ( .A(n_516), .Y(n_719) );
BUFx3_ASAP7_75t_L g519 ( .A(n_520), .Y(n_519) );
BUFx6f_ASAP7_75t_L g612 ( .A(n_520), .Y(n_612) );
BUFx3_ASAP7_75t_L g715 ( .A(n_520), .Y(n_715) );
INVx1_ASAP7_75t_L g1123 ( .A(n_520), .Y(n_1123) );
BUFx3_ASAP7_75t_L g1190 ( .A(n_520), .Y(n_1190) );
AND2x2_ASAP7_75t_L g1424 ( .A(n_520), .B(n_1425), .Y(n_1424) );
BUFx6f_ASAP7_75t_L g520 ( .A(n_521), .Y(n_520) );
INVx1_ASAP7_75t_L g541 ( .A(n_521), .Y(n_541) );
BUFx2_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
INVx1_ASAP7_75t_L g1359 ( .A(n_523), .Y(n_1359) );
HB1xp67_ASAP7_75t_L g1550 ( .A(n_523), .Y(n_1550) );
HB1xp67_ASAP7_75t_SL g1255 ( .A(n_524), .Y(n_1255) );
INVx4_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
INVx1_ASAP7_75t_SL g613 ( .A(n_525), .Y(n_613) );
INVx4_ASAP7_75t_L g773 ( .A(n_525), .Y(n_773) );
NAND4xp25_ASAP7_75t_L g935 ( .A(n_525), .B(n_936), .C(n_937), .D(n_939), .Y(n_935) );
NAND2xp5_ASAP7_75t_L g1418 ( .A(n_525), .B(n_1419), .Y(n_1418) );
INVx2_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
INVx2_ASAP7_75t_SL g536 ( .A(n_528), .Y(n_536) );
INVx2_ASAP7_75t_L g770 ( .A(n_528), .Y(n_770) );
INVx1_ASAP7_75t_L g938 ( .A(n_528), .Y(n_938) );
INVx2_ASAP7_75t_L g1009 ( .A(n_528), .Y(n_1009) );
INVx1_ASAP7_75t_L g1257 ( .A(n_528), .Y(n_1257) );
BUFx3_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
INVx1_ASAP7_75t_SL g1011 ( .A(n_530), .Y(n_1011) );
HB1xp67_ASAP7_75t_L g1805 ( .A(n_530), .Y(n_1805) );
HB1xp67_ASAP7_75t_L g1814 ( .A(n_530), .Y(n_1814) );
AOI21xp5_ASAP7_75t_L g608 ( .A1(n_531), .A2(n_609), .B(n_614), .Y(n_608) );
AOI21xp5_ASAP7_75t_L g687 ( .A1(n_531), .A2(n_688), .B(n_689), .Y(n_687) );
AOI21xp5_ASAP7_75t_L g713 ( .A1(n_531), .A2(n_714), .B(n_718), .Y(n_713) );
AOI21xp5_ASAP7_75t_L g1006 ( .A1(n_531), .A2(n_1007), .B(n_1008), .Y(n_1006) );
INVx1_ASAP7_75t_L g1060 ( .A(n_531), .Y(n_1060) );
AOI21xp5_ASAP7_75t_L g1153 ( .A1(n_531), .A2(n_1154), .B(n_1156), .Y(n_1153) );
AOI21xp5_ASAP7_75t_L g1188 ( .A1(n_531), .A2(n_1189), .B(n_1191), .Y(n_1188) );
AOI21xp5_ASAP7_75t_L g1253 ( .A1(n_531), .A2(n_1254), .B(n_1256), .Y(n_1253) );
AOI221xp5_ASAP7_75t_L g1292 ( .A1(n_531), .A2(n_761), .B1(n_1272), .B2(n_1293), .C(n_1294), .Y(n_1292) );
AOI221xp5_ASAP7_75t_L g1332 ( .A1(n_531), .A2(n_761), .B1(n_1314), .B2(n_1333), .C(n_1334), .Y(n_1332) );
AOI21xp5_ASAP7_75t_L g1356 ( .A1(n_531), .A2(n_1357), .B(n_1360), .Y(n_1356) );
AOI21xp5_ASAP7_75t_L g1548 ( .A1(n_531), .A2(n_1549), .B(n_1551), .Y(n_1548) );
AOI221xp5_ASAP7_75t_L g1808 ( .A1(n_531), .A2(n_533), .B1(n_1809), .B2(n_1810), .C(n_1813), .Y(n_1808) );
NAND2xp5_ASAP7_75t_L g923 ( .A(n_533), .B(n_924), .Y(n_923) );
INVx1_ASAP7_75t_L g1125 ( .A(n_533), .Y(n_1125) );
AOI222xp33_ASAP7_75t_L g1335 ( .A1(n_533), .A2(n_550), .B1(n_1318), .B2(n_1319), .C1(n_1336), .C2(n_1337), .Y(n_1335) );
BUFx3_ASAP7_75t_L g533 ( .A(n_534), .Y(n_533) );
INVx2_ASAP7_75t_L g623 ( .A(n_534), .Y(n_623) );
INVx2_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
INVx1_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
INVx1_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
BUFx2_ASAP7_75t_L g641 ( .A(n_541), .Y(n_641) );
INVx1_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
INVx1_ASAP7_75t_L g543 ( .A(n_544), .Y(n_543) );
INVx2_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
INVx2_ASAP7_75t_L g1119 ( .A(n_545), .Y(n_1119) );
INVx1_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
INVx2_ASAP7_75t_L g644 ( .A(n_547), .Y(n_644) );
INVx2_ASAP7_75t_L g703 ( .A(n_547), .Y(n_703) );
INVx3_ASAP7_75t_L g768 ( .A(n_547), .Y(n_768) );
OAI221xp5_ASAP7_75t_L g1015 ( .A1(n_547), .A2(n_1016), .B1(n_1017), .B2(n_1018), .C(n_1021), .Y(n_1015) );
INVx1_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
INVx1_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g1349 ( .A(n_550), .B(n_1350), .Y(n_1349) );
AOI22xp33_ASAP7_75t_L g1496 ( .A1(n_550), .A2(n_1497), .B1(n_1498), .B2(n_1499), .Y(n_1496) );
NAND2xp5_ASAP7_75t_L g1541 ( .A(n_550), .B(n_1542), .Y(n_1541) );
AOI222xp33_ASAP7_75t_L g1802 ( .A1(n_550), .A2(n_1004), .B1(n_1803), .B2(n_1804), .C1(n_1806), .C2(n_1807), .Y(n_1802) );
AOI22xp5_ASAP7_75t_L g778 ( .A1(n_551), .A2(n_779), .B1(n_780), .B2(n_782), .Y(n_778) );
AOI22xp33_ASAP7_75t_L g929 ( .A1(n_551), .A2(n_780), .B1(n_930), .B2(n_931), .Y(n_929) );
BUFx2_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
INVx1_ASAP7_75t_L g627 ( .A(n_552), .Y(n_627) );
INVx1_ASAP7_75t_L g891 ( .A(n_552), .Y(n_891) );
AND2x4_ASAP7_75t_L g1428 ( .A(n_552), .B(n_1429), .Y(n_1428) );
OAI21xp5_ASAP7_75t_L g684 ( .A1(n_553), .A2(n_685), .B(n_696), .Y(n_684) );
OAI21xp5_ASAP7_75t_L g1001 ( .A1(n_553), .A2(n_1002), .B(n_1013), .Y(n_1001) );
AOI21xp5_ASAP7_75t_L g1327 ( .A1(n_553), .A2(n_1328), .B(n_1338), .Y(n_1327) );
OAI21xp5_ASAP7_75t_SL g1347 ( .A1(n_553), .A2(n_1348), .B(n_1355), .Y(n_1347) );
OAI21xp5_ASAP7_75t_L g1489 ( .A1(n_553), .A2(n_1490), .B(n_1495), .Y(n_1489) );
OAI21xp5_ASAP7_75t_SL g1539 ( .A1(n_553), .A2(n_1540), .B(n_1547), .Y(n_1539) );
INVx2_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
INVx1_ASAP7_75t_L g1308 ( .A(n_554), .Y(n_1308) );
BUFx2_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
NAND2xp5_ASAP7_75t_L g915 ( .A(n_555), .B(n_916), .Y(n_915) );
INVx1_ASAP7_75t_L g1879 ( .A(n_555), .Y(n_1879) );
INVx1_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
OR2x6_ASAP7_75t_L g798 ( .A(n_556), .B(n_799), .Y(n_798) );
AND2x4_ASAP7_75t_L g878 ( .A(n_556), .B(n_879), .Y(n_878) );
OR2x2_ASAP7_75t_L g1322 ( .A(n_556), .B(n_799), .Y(n_1322) );
HB1xp67_ASAP7_75t_L g1214 ( .A(n_558), .Y(n_1214) );
INVx2_ASAP7_75t_L g1506 ( .A(n_558), .Y(n_1506) );
AND2x4_ASAP7_75t_L g558 ( .A(n_559), .B(n_563), .Y(n_558) );
AND2x4_ASAP7_75t_L g656 ( .A(n_559), .B(n_563), .Y(n_656) );
INVx1_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
INVx2_ASAP7_75t_L g814 ( .A(n_563), .Y(n_814) );
INVx3_ASAP7_75t_L g859 ( .A(n_564), .Y(n_859) );
INVx4_ASAP7_75t_L g1520 ( .A(n_564), .Y(n_1520) );
BUFx6f_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
BUFx2_ASAP7_75t_L g846 ( .A(n_565), .Y(n_846) );
BUFx3_ASAP7_75t_L g1398 ( .A(n_565), .Y(n_1398) );
BUFx2_ASAP7_75t_L g1471 ( .A(n_566), .Y(n_1471) );
AOI22xp33_ASAP7_75t_L g707 ( .A1(n_568), .A2(n_571), .B1(n_694), .B2(n_695), .Y(n_707) );
AOI22xp33_ASAP7_75t_L g750 ( .A1(n_568), .A2(n_571), .B1(n_721), .B2(n_722), .Y(n_750) );
AOI22xp33_ASAP7_75t_L g998 ( .A1(n_568), .A2(n_571), .B1(n_999), .B2(n_1000), .Y(n_998) );
AOI22xp33_ASAP7_75t_L g1128 ( .A1(n_568), .A2(n_571), .B1(n_1107), .B2(n_1108), .Y(n_1128) );
AOI22xp33_ASAP7_75t_L g1215 ( .A1(n_568), .A2(n_571), .B1(n_1197), .B2(n_1199), .Y(n_1215) );
AOI22xp5_ASAP7_75t_L g1309 ( .A1(n_568), .A2(n_1297), .B1(n_1298), .B2(n_1310), .Y(n_1309) );
NAND2xp5_ASAP7_75t_L g1859 ( .A(n_568), .B(n_1860), .Y(n_1859) );
AND2x4_ASAP7_75t_L g568 ( .A(n_569), .B(n_570), .Y(n_568) );
AND2x4_ASAP7_75t_L g815 ( .A(n_569), .B(n_570), .Y(n_815) );
AOI22xp5_ASAP7_75t_L g866 ( .A1(n_569), .A2(n_796), .B1(n_831), .B2(n_867), .Y(n_866) );
INVx2_ASAP7_75t_L g599 ( .A(n_571), .Y(n_599) );
INVx2_ASAP7_75t_L g1230 ( .A(n_571), .Y(n_1230) );
NAND2xp5_ASAP7_75t_L g1535 ( .A(n_571), .B(n_1501), .Y(n_1535) );
NAND3xp33_ASAP7_75t_L g574 ( .A(n_575), .B(n_601), .C(n_605), .Y(n_574) );
NOR3xp33_ASAP7_75t_L g575 ( .A(n_576), .B(n_592), .C(n_600), .Y(n_575) );
NAND2xp5_ASAP7_75t_L g576 ( .A(n_577), .B(n_581), .Y(n_576) );
INVx1_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
BUFx2_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
OAI221xp5_ASAP7_75t_L g663 ( .A1(n_587), .A2(n_664), .B1(n_665), .B2(n_669), .C(n_670), .Y(n_663) );
INVx3_ASAP7_75t_L g807 ( .A(n_587), .Y(n_807) );
OR2x6_ASAP7_75t_SL g836 ( .A(n_587), .B(n_837), .Y(n_836) );
BUFx2_ASAP7_75t_L g1142 ( .A(n_587), .Y(n_1142) );
INVx1_ASAP7_75t_L g1822 ( .A(n_587), .Y(n_1822) );
BUFx2_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g966 ( .A(n_593), .B(n_967), .Y(n_966) );
OR2x6_ASAP7_75t_L g593 ( .A(n_594), .B(n_597), .Y(n_593) );
INVx2_ASAP7_75t_SL g1238 ( .A(n_594), .Y(n_1238) );
OR2x2_ASAP7_75t_L g1379 ( .A(n_594), .B(n_597), .Y(n_1379) );
INVx2_ASAP7_75t_SL g594 ( .A(n_595), .Y(n_594) );
INVx2_ASAP7_75t_L g595 ( .A(n_596), .Y(n_595) );
BUFx4f_ASAP7_75t_L g841 ( .A(n_596), .Y(n_841) );
OR2x4_ASAP7_75t_L g1476 ( .A(n_596), .B(n_1458), .Y(n_1476) );
BUFx3_ASAP7_75t_L g1516 ( .A(n_596), .Y(n_1516) );
BUFx3_ASAP7_75t_L g1527 ( .A(n_596), .Y(n_1527) );
INVxp67_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
AND2x2_ASAP7_75t_L g806 ( .A(n_598), .B(n_807), .Y(n_806) );
INVxp67_ASAP7_75t_L g1310 ( .A(n_599), .Y(n_1310) );
NOR4xp25_ASAP7_75t_L g1226 ( .A(n_600), .B(n_1227), .C(n_1229), .D(n_1231), .Y(n_1226) );
NAND2xp5_ASAP7_75t_L g908 ( .A(n_604), .B(n_909), .Y(n_908) );
OAI21xp5_ASAP7_75t_L g605 ( .A1(n_606), .A2(n_620), .B(n_645), .Y(n_605) );
INVx1_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
INVx1_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
BUFx2_ASAP7_75t_L g1155 ( .A(n_612), .Y(n_1155) );
AOI22xp33_ASAP7_75t_L g1157 ( .A1(n_618), .A2(n_1004), .B1(n_1158), .B2(n_1159), .Y(n_1157) );
INVx1_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
INVx2_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
INVx2_ASAP7_75t_L g724 ( .A(n_622), .Y(n_724) );
INVx1_ASAP7_75t_L g1014 ( .A(n_622), .Y(n_1014) );
AOI22xp33_ASAP7_75t_L g1165 ( .A1(n_622), .A2(n_626), .B1(n_1136), .B2(n_1137), .Y(n_1165) );
INVx4_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
BUFx2_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
INVx2_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
INVx2_ASAP7_75t_L g1300 ( .A(n_626), .Y(n_1300) );
NOR2x1_ASAP7_75t_L g626 ( .A(n_627), .B(n_628), .Y(n_626) );
INVx1_ASAP7_75t_L g783 ( .A(n_628), .Y(n_783) );
OAI221xp5_ASAP7_75t_L g629 ( .A1(n_630), .A2(n_633), .B1(n_634), .B2(n_638), .C(n_639), .Y(n_629) );
OAI22xp5_ASAP7_75t_L g1022 ( .A1(n_630), .A2(n_1023), .B1(n_1024), .B2(n_1025), .Y(n_1022) );
INVx2_ASAP7_75t_L g630 ( .A(n_631), .Y(n_630) );
BUFx6f_ASAP7_75t_L g631 ( .A(n_632), .Y(n_631) );
INVx3_ASAP7_75t_L g776 ( .A(n_632), .Y(n_776) );
INVx4_ASAP7_75t_L g927 ( .A(n_632), .Y(n_927) );
INVx1_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
INVx4_ASAP7_75t_L g934 ( .A(n_635), .Y(n_934) );
BUFx6f_ASAP7_75t_L g1026 ( .A(n_635), .Y(n_1026) );
INVx2_ASAP7_75t_L g1072 ( .A(n_635), .Y(n_1072) );
INVx2_ASAP7_75t_L g1211 ( .A(n_635), .Y(n_1211) );
INVx1_ASAP7_75t_L g1305 ( .A(n_635), .Y(n_1305) );
INVx2_ASAP7_75t_SL g1867 ( .A(n_635), .Y(n_1867) );
INVx8_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
OR2x2_ASAP7_75t_L g1443 ( .A(n_636), .B(n_1429), .Y(n_1443) );
BUFx2_ASAP7_75t_L g1874 ( .A(n_636), .Y(n_1874) );
BUFx6f_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
INVx1_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
INVx2_ASAP7_75t_L g1113 ( .A(n_641), .Y(n_1113) );
BUFx3_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
OAI21xp5_ASAP7_75t_L g1151 ( .A1(n_645), .A2(n_1152), .B(n_1160), .Y(n_1151) );
OAI21xp5_ASAP7_75t_L g1248 ( .A1(n_645), .A2(n_1249), .B(n_1252), .Y(n_1248) );
AOI221xp5_ASAP7_75t_L g1799 ( .A1(n_645), .A2(n_1506), .B1(n_1800), .B2(n_1801), .C(n_1818), .Y(n_1799) );
INVx2_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
INVx1_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
HB1xp67_ASAP7_75t_L g944 ( .A(n_647), .Y(n_944) );
BUFx2_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
BUFx2_ASAP7_75t_L g732 ( .A(n_648), .Y(n_732) );
AOI21x1_ASAP7_75t_L g758 ( .A1(n_648), .A2(n_759), .B(n_787), .Y(n_758) );
BUFx3_ASAP7_75t_L g649 ( .A(n_650), .Y(n_649) );
AO22x2_ASAP7_75t_L g650 ( .A1(n_651), .A2(n_708), .B1(n_709), .B2(n_751), .Y(n_650) );
INVx1_ASAP7_75t_L g751 ( .A(n_651), .Y(n_751) );
AND4x1_ASAP7_75t_L g652 ( .A(n_653), .B(n_657), .C(n_684), .D(n_707), .Y(n_652) );
INVx1_ASAP7_75t_SL g1271 ( .A(n_656), .Y(n_1271) );
NOR3xp33_ASAP7_75t_L g657 ( .A(n_658), .B(n_659), .C(n_681), .Y(n_657) );
NOR3xp33_ASAP7_75t_L g1133 ( .A(n_658), .B(n_1134), .C(n_1147), .Y(n_1133) );
NOR3xp33_ASAP7_75t_L g1368 ( .A(n_658), .B(n_1369), .C(n_1378), .Y(n_1368) );
OAI22xp5_ASAP7_75t_SL g659 ( .A1(n_660), .A2(n_663), .B1(n_672), .B2(n_673), .Y(n_659) );
BUFx3_ASAP7_75t_L g1384 ( .A(n_660), .Y(n_1384) );
BUFx4f_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
BUFx8_ASAP7_75t_L g735 ( .A(n_661), .Y(n_735) );
BUFx2_ASAP7_75t_L g950 ( .A(n_661), .Y(n_950) );
BUFx4f_ASAP7_75t_L g1275 ( .A(n_661), .Y(n_1275) );
OAI221xp5_ASAP7_75t_L g736 ( .A1(n_665), .A2(n_737), .B1(n_738), .B2(n_739), .C(n_740), .Y(n_736) );
INVx3_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
BUFx2_ASAP7_75t_L g666 ( .A(n_667), .Y(n_666) );
INVx1_ASAP7_75t_L g667 ( .A(n_668), .Y(n_667) );
BUFx3_ASAP7_75t_L g1283 ( .A(n_668), .Y(n_1283) );
OAI221xp5_ASAP7_75t_L g673 ( .A1(n_674), .A2(n_676), .B1(n_677), .B2(n_679), .C(n_680), .Y(n_673) );
INVx1_ASAP7_75t_L g1044 ( .A(n_674), .Y(n_1044) );
INVx2_ASAP7_75t_L g674 ( .A(n_675), .Y(n_674) );
BUFx6f_ASAP7_75t_L g792 ( .A(n_675), .Y(n_792) );
BUFx6f_ASAP7_75t_L g794 ( .A(n_675), .Y(n_794) );
INVx2_ASAP7_75t_L g1392 ( .A(n_675), .Y(n_1392) );
AND2x4_ASAP7_75t_L g1457 ( .A(n_675), .B(n_1458), .Y(n_1457) );
INVx2_ASAP7_75t_L g1885 ( .A(n_675), .Y(n_1885) );
OAI211xp5_ASAP7_75t_L g697 ( .A1(n_676), .A2(n_698), .B(n_702), .C(n_704), .Y(n_697) );
OAI221xp5_ASAP7_75t_L g741 ( .A1(n_677), .A2(n_726), .B1(n_737), .B2(n_742), .C(n_743), .Y(n_741) );
CKINVDCx8_ASAP7_75t_R g677 ( .A(n_678), .Y(n_677) );
INVx3_ASAP7_75t_L g843 ( .A(n_678), .Y(n_843) );
INVx3_ASAP7_75t_L g855 ( .A(n_678), .Y(n_855) );
INVx3_ASAP7_75t_L g953 ( .A(n_678), .Y(n_953) );
INVx1_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
AOI22xp5_ASAP7_75t_L g1035 ( .A1(n_683), .A2(n_801), .B1(n_1036), .B2(n_1037), .Y(n_1035) );
AOI22xp5_ASAP7_75t_L g1317 ( .A1(n_683), .A2(n_801), .B1(n_1318), .B2(n_1319), .Y(n_1317) );
AOI22xp33_ASAP7_75t_L g1370 ( .A1(n_683), .A2(n_801), .B1(n_1350), .B2(n_1371), .Y(n_1370) );
AOI22xp33_ASAP7_75t_L g1560 ( .A1(n_683), .A2(n_801), .B1(n_1542), .B2(n_1561), .Y(n_1560) );
INVx2_ASAP7_75t_SL g690 ( .A(n_691), .Y(n_690) );
INVx1_ASAP7_75t_L g1295 ( .A(n_691), .Y(n_1295) );
INVx2_ASAP7_75t_L g1361 ( .A(n_691), .Y(n_1361) );
INVx3_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
BUFx6f_ASAP7_75t_L g1193 ( .A(n_692), .Y(n_1193) );
INVx1_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
INVx2_ASAP7_75t_L g777 ( .A(n_699), .Y(n_777) );
INVx2_ASAP7_75t_L g928 ( .A(n_699), .Y(n_928) );
INVx4_ASAP7_75t_L g699 ( .A(n_700), .Y(n_699) );
BUFx4f_ASAP7_75t_L g786 ( .A(n_700), .Y(n_786) );
OR2x6_ASAP7_75t_L g904 ( .A(n_700), .B(n_905), .Y(n_904) );
BUFx4f_ASAP7_75t_L g1016 ( .A(n_700), .Y(n_1016) );
BUFx4f_ASAP7_75t_L g1053 ( .A(n_700), .Y(n_1053) );
BUFx6f_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
BUFx3_ASAP7_75t_L g729 ( .A(n_701), .Y(n_729) );
INVx1_ASAP7_75t_L g1066 ( .A(n_703), .Y(n_1066) );
INVx1_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
INVx3_ASAP7_75t_L g762 ( .A(n_706), .Y(n_762) );
INVx1_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
AND4x1_ASAP7_75t_L g710 ( .A(n_711), .B(n_733), .C(n_747), .D(n_750), .Y(n_710) );
OAI21xp5_ASAP7_75t_L g711 ( .A1(n_712), .A2(n_723), .B(n_732), .Y(n_711) );
INVx2_ASAP7_75t_SL g716 ( .A(n_717), .Y(n_716) );
OAI211xp5_ASAP7_75t_L g725 ( .A1(n_726), .A2(n_727), .B(n_730), .C(n_731), .Y(n_725) );
OAI211xp5_ASAP7_75t_L g940 ( .A1(n_727), .A2(n_941), .B(n_942), .C(n_943), .Y(n_940) );
OAI22xp5_ASAP7_75t_L g1411 ( .A1(n_727), .A2(n_933), .B1(n_1391), .B2(n_1396), .Y(n_1411) );
INVx5_ASAP7_75t_L g727 ( .A(n_728), .Y(n_727) );
INVx2_ASAP7_75t_SL g728 ( .A(n_729), .Y(n_728) );
OR2x2_ASAP7_75t_L g893 ( .A(n_729), .B(n_894), .Y(n_893) );
BUFx2_ASAP7_75t_SL g1202 ( .A(n_729), .Y(n_1202) );
O2A1O1Ixp5_ASAP7_75t_SL g1049 ( .A1(n_732), .A2(n_1050), .B(n_1061), .C(n_1073), .Y(n_1049) );
OAI33xp33_ASAP7_75t_L g1231 ( .A1(n_735), .A2(n_1232), .A3(n_1236), .B1(n_1241), .B2(n_1244), .B3(n_1247), .Y(n_1231) );
INVx2_ASAP7_75t_L g744 ( .A(n_745), .Y(n_744) );
INVx2_ASAP7_75t_L g796 ( .A(n_745), .Y(n_796) );
INVx1_ASAP7_75t_L g1042 ( .A(n_745), .Y(n_1042) );
INVx1_ASAP7_75t_L g1181 ( .A(n_745), .Y(n_1181) );
INVx1_ASAP7_75t_L g752 ( .A(n_753), .Y(n_752) );
AO22x2_ASAP7_75t_L g753 ( .A1(n_754), .A2(n_971), .B1(n_1028), .B2(n_1029), .Y(n_753) );
INVx1_ASAP7_75t_L g1028 ( .A(n_754), .Y(n_1028) );
XNOR2xp5_ASAP7_75t_L g754 ( .A(n_755), .B(n_919), .Y(n_754) );
OAI22xp5_ASAP7_75t_L g755 ( .A1(n_756), .A2(n_826), .B1(n_917), .B2(n_918), .Y(n_755) );
INVx1_ASAP7_75t_L g918 ( .A(n_756), .Y(n_918) );
NAND3xp33_ASAP7_75t_L g756 ( .A(n_757), .B(n_819), .C(n_823), .Y(n_756) );
INVx1_ASAP7_75t_L g820 ( .A(n_758), .Y(n_820) );
INVx2_ASAP7_75t_L g760 ( .A(n_761), .Y(n_760) );
AND2x4_ASAP7_75t_L g910 ( .A(n_762), .B(n_911), .Y(n_910) );
AOI22xp5_ASAP7_75t_L g763 ( .A1(n_764), .A2(n_765), .B1(n_769), .B2(n_771), .Y(n_763) );
INVx2_ASAP7_75t_L g766 ( .A(n_767), .Y(n_766) );
INVx2_ASAP7_75t_L g772 ( .A(n_767), .Y(n_772) );
INVx2_ASAP7_75t_L g1112 ( .A(n_772), .Y(n_1112) );
HB1xp67_ASAP7_75t_L g1163 ( .A(n_772), .Y(n_1163) );
INVx1_ASAP7_75t_L g1812 ( .A(n_772), .Y(n_1812) );
AOI22xp5_ASAP7_75t_L g774 ( .A1(n_775), .A2(n_783), .B1(n_784), .B2(n_785), .Y(n_774) );
INVx2_ASAP7_75t_SL g1408 ( .A(n_776), .Y(n_1408) );
INVx1_ASAP7_75t_L g780 ( .A(n_781), .Y(n_780) );
AOI222xp33_ASAP7_75t_L g813 ( .A1(n_782), .A2(n_814), .B1(n_815), .B2(n_816), .C1(n_817), .C2(n_818), .Y(n_813) );
AOI22xp5_ASAP7_75t_L g925 ( .A1(n_783), .A2(n_784), .B1(n_926), .B2(n_932), .Y(n_925) );
OAI211xp5_ASAP7_75t_L g1351 ( .A1(n_786), .A2(n_1352), .B(n_1353), .C(n_1354), .Y(n_1351) );
OAI211xp5_ASAP7_75t_L g1543 ( .A1(n_786), .A2(n_1544), .B(n_1545), .C(n_1546), .Y(n_1543) );
INVx1_ASAP7_75t_L g821 ( .A(n_788), .Y(n_821) );
AND2x2_ASAP7_75t_L g788 ( .A(n_789), .B(n_800), .Y(n_788) );
INVx2_ASAP7_75t_L g1523 ( .A(n_792), .Y(n_1523) );
INVx1_ASAP7_75t_L g1830 ( .A(n_794), .Y(n_1830) );
INVx1_ASAP7_75t_L g797 ( .A(n_798), .Y(n_797) );
INVx1_ASAP7_75t_L g1048 ( .A(n_798), .Y(n_1048) );
INVx1_ASAP7_75t_SL g1376 ( .A(n_798), .Y(n_1376) );
INVx1_ASAP7_75t_L g825 ( .A(n_803), .Y(n_825) );
NAND2xp5_ASAP7_75t_L g803 ( .A(n_804), .B(n_812), .Y(n_803) );
NAND2x1_ASAP7_75t_L g804 ( .A(n_805), .B(n_808), .Y(n_804) );
INVx2_ASAP7_75t_SL g805 ( .A(n_806), .Y(n_805) );
AOI22xp33_ASAP7_75t_L g1074 ( .A1(n_806), .A2(n_815), .B1(n_1057), .B2(n_1058), .Y(n_1074) );
AOI22xp33_ASAP7_75t_L g1339 ( .A1(n_806), .A2(n_815), .B1(n_1330), .B2(n_1331), .Y(n_1339) );
INVx2_ASAP7_75t_L g1281 ( .A(n_807), .Y(n_1281) );
INVx2_ASAP7_75t_L g808 ( .A(n_809), .Y(n_808) );
AOI22xp33_ASAP7_75t_L g830 ( .A1(n_809), .A2(n_831), .B1(n_832), .B2(n_833), .Y(n_830) );
AND2x4_ASAP7_75t_L g809 ( .A(n_810), .B(n_811), .Y(n_809) );
INVx1_ASAP7_75t_L g824 ( .A(n_813), .Y(n_824) );
AOI22xp5_ASAP7_75t_L g946 ( .A1(n_814), .A2(n_817), .B1(n_931), .B2(n_947), .Y(n_946) );
OAI21xp5_ASAP7_75t_L g819 ( .A1(n_820), .A2(n_821), .B(n_822), .Y(n_819) );
OAI21xp33_ASAP7_75t_L g823 ( .A1(n_822), .A2(n_824), .B(n_825), .Y(n_823) );
INVx1_ASAP7_75t_L g917 ( .A(n_826), .Y(n_917) );
XNOR2xp5_ASAP7_75t_L g826 ( .A(n_827), .B(n_828), .Y(n_826) );
NOR2x1_ASAP7_75t_L g828 ( .A(n_829), .B(n_874), .Y(n_828) );
NAND2xp5_ASAP7_75t_L g829 ( .A(n_830), .B(n_834), .Y(n_829) );
INVx3_ASAP7_75t_L g967 ( .A(n_832), .Y(n_967) );
INVx2_ASAP7_75t_L g837 ( .A(n_838), .Y(n_837) );
HB1xp67_ASAP7_75t_L g869 ( .A(n_838), .Y(n_869) );
OAI221xp5_ASAP7_75t_L g839 ( .A1(n_840), .A2(n_845), .B1(n_852), .B2(n_857), .C(n_863), .Y(n_839) );
OAI22xp5_ASAP7_75t_L g840 ( .A1(n_841), .A2(n_842), .B1(n_843), .B2(n_844), .Y(n_840) );
HB1xp67_ASAP7_75t_L g1387 ( .A(n_841), .Y(n_1387) );
INVx1_ASAP7_75t_L g1827 ( .A(n_841), .Y(n_1827) );
OAI22xp33_ASAP7_75t_L g1401 ( .A1(n_843), .A2(n_1387), .B1(n_1402), .B2(n_1403), .Y(n_1401) );
OAI221xp5_ASAP7_75t_L g845 ( .A1(n_846), .A2(n_847), .B1(n_848), .B2(n_850), .C(n_851), .Y(n_845) );
OR2x6_ASAP7_75t_L g863 ( .A(n_846), .B(n_864), .Y(n_863) );
INVx1_ASAP7_75t_L g1529 ( .A(n_846), .Y(n_1529) );
OAI211xp5_ASAP7_75t_L g898 ( .A1(n_847), .A2(n_899), .B(n_902), .C(n_903), .Y(n_898) );
INVx3_ASAP7_75t_L g848 ( .A(n_849), .Y(n_848) );
INVx2_ASAP7_75t_SL g853 ( .A(n_849), .Y(n_853) );
INVx5_ASAP7_75t_L g959 ( .A(n_849), .Y(n_959) );
OAI22xp5_ASAP7_75t_L g852 ( .A1(n_853), .A2(n_854), .B1(n_855), .B2(n_856), .Y(n_852) );
OAI221xp5_ASAP7_75t_L g951 ( .A1(n_853), .A2(n_952), .B1(n_953), .B2(n_954), .C(n_955), .Y(n_951) );
OAI211xp5_ASAP7_75t_L g1276 ( .A1(n_853), .A2(n_1277), .B(n_1278), .C(n_1279), .Y(n_1276) );
OAI22xp33_ASAP7_75t_L g1232 ( .A1(n_855), .A2(n_1233), .B1(n_1234), .B2(n_1235), .Y(n_1232) );
OAI22xp5_ASAP7_75t_L g1390 ( .A1(n_855), .A2(n_1391), .B1(n_1392), .B2(n_1393), .Y(n_1390) );
OAI21xp5_ASAP7_75t_SL g857 ( .A1(n_858), .A2(n_860), .B(n_861), .Y(n_857) );
INVx3_ASAP7_75t_L g858 ( .A(n_859), .Y(n_858) );
INVx2_ASAP7_75t_L g1234 ( .A(n_859), .Y(n_1234) );
INVx2_ASAP7_75t_L g1389 ( .A(n_859), .Y(n_1389) );
AOI22xp5_ASAP7_75t_L g882 ( .A1(n_867), .A2(n_883), .B1(n_885), .B2(n_886), .Y(n_882) );
INVx1_ASAP7_75t_L g868 ( .A(n_869), .Y(n_868) );
INVx4_ASAP7_75t_L g870 ( .A(n_871), .Y(n_870) );
INVx2_ASAP7_75t_L g872 ( .A(n_873), .Y(n_872) );
NAND3xp33_ASAP7_75t_L g874 ( .A(n_875), .B(n_906), .C(n_912), .Y(n_874) );
NOR3xp33_ASAP7_75t_SL g875 ( .A(n_876), .B(n_892), .C(n_895), .Y(n_875) );
OAI21xp5_ASAP7_75t_SL g876 ( .A1(n_877), .A2(n_881), .B(n_882), .Y(n_876) );
NAND2xp5_ASAP7_75t_L g877 ( .A(n_878), .B(n_880), .Y(n_877) );
INVx4_ASAP7_75t_L g1405 ( .A(n_878), .Y(n_1405) );
INVx1_ASAP7_75t_SL g883 ( .A(n_884), .Y(n_883) );
INVx2_ASAP7_75t_SL g886 ( .A(n_887), .Y(n_886) );
NAND2x2_ASAP7_75t_L g887 ( .A(n_888), .B(n_890), .Y(n_887) );
INVx1_ASAP7_75t_L g905 ( .A(n_888), .Y(n_905) );
INVx2_ASAP7_75t_L g888 ( .A(n_889), .Y(n_888) );
INVx2_ASAP7_75t_SL g890 ( .A(n_891), .Y(n_890) );
INVx1_ASAP7_75t_L g911 ( .A(n_894), .Y(n_911) );
OAI21xp5_ASAP7_75t_L g895 ( .A1(n_896), .A2(n_898), .B(n_904), .Y(n_895) );
INVx2_ASAP7_75t_L g896 ( .A(n_897), .Y(n_896) );
INVx2_ASAP7_75t_L g899 ( .A(n_900), .Y(n_899) );
INVx1_ASAP7_75t_L g900 ( .A(n_901), .Y(n_900) );
BUFx2_ASAP7_75t_L g933 ( .A(n_901), .Y(n_933) );
BUFx2_ASAP7_75t_L g1020 ( .A(n_901), .Y(n_1020) );
BUFx3_ASAP7_75t_L g1064 ( .A(n_901), .Y(n_1064) );
NAND2xp5_ASAP7_75t_L g906 ( .A(n_907), .B(n_908), .Y(n_906) );
INVx1_ASAP7_75t_L g909 ( .A(n_910), .Y(n_909) );
NAND2xp5_ASAP7_75t_L g912 ( .A(n_913), .B(n_914), .Y(n_912) );
AOI21xp5_ASAP7_75t_L g921 ( .A1(n_922), .A2(n_944), .B(n_945), .Y(n_921) );
NAND4xp25_ASAP7_75t_L g922 ( .A(n_923), .B(n_925), .C(n_935), .D(n_940), .Y(n_922) );
OAI221xp5_ASAP7_75t_L g1062 ( .A1(n_928), .A2(n_1063), .B1(n_1064), .B2(n_1065), .C(n_1066), .Y(n_1062) );
OAI22xp5_ASAP7_75t_L g1412 ( .A1(n_933), .A2(n_1388), .B1(n_1403), .B2(n_1409), .Y(n_1412) );
INVx2_ASAP7_75t_L g1410 ( .A(n_934), .Y(n_1410) );
OAI221xp5_ASAP7_75t_L g958 ( .A1(n_941), .A2(n_959), .B1(n_960), .B2(n_961), .C(n_962), .Y(n_958) );
OAI22xp5_ASAP7_75t_SL g949 ( .A1(n_950), .A2(n_951), .B1(n_957), .B2(n_958), .Y(n_949) );
OAI22xp5_ASAP7_75t_L g1883 ( .A1(n_953), .A2(n_1865), .B1(n_1884), .B2(n_1885), .Y(n_1883) );
INVx2_ASAP7_75t_SL g987 ( .A(n_956), .Y(n_987) );
BUFx3_ASAP7_75t_L g1564 ( .A(n_956), .Y(n_1564) );
OAI22xp5_ASAP7_75t_L g1274 ( .A1(n_957), .A2(n_1275), .B1(n_1276), .B2(n_1280), .Y(n_1274) );
INVx8_ASAP7_75t_L g1144 ( .A(n_959), .Y(n_1144) );
BUFx3_ASAP7_75t_L g1180 ( .A(n_959), .Y(n_1180) );
OAI22xp5_ASAP7_75t_L g1521 ( .A1(n_960), .A2(n_1522), .B1(n_1523), .B2(n_1524), .Y(n_1521) );
OAI22xp5_ASAP7_75t_L g1819 ( .A1(n_960), .A2(n_1820), .B1(n_1821), .B2(n_1823), .Y(n_1819) );
NAND2xp5_ASAP7_75t_L g964 ( .A(n_965), .B(n_966), .Y(n_964) );
NAND2xp5_ASAP7_75t_L g968 ( .A(n_969), .B(n_970), .Y(n_968) );
NAND2xp5_ASAP7_75t_L g981 ( .A(n_970), .B(n_982), .Y(n_981) );
NAND2xp5_ASAP7_75t_L g1038 ( .A(n_970), .B(n_1039), .Y(n_1038) );
NAND2xp5_ASAP7_75t_L g1174 ( .A(n_970), .B(n_1175), .Y(n_1174) );
NAND2xp5_ASAP7_75t_L g1534 ( .A(n_970), .B(n_1502), .Y(n_1534) );
INVx2_ASAP7_75t_L g1029 ( .A(n_971), .Y(n_1029) );
XOR2x2_ASAP7_75t_L g971 ( .A(n_972), .B(n_1027), .Y(n_971) );
NAND2xp5_ASAP7_75t_SL g972 ( .A(n_973), .B(n_1001), .Y(n_972) );
NAND2xp5_ASAP7_75t_L g975 ( .A(n_976), .B(n_984), .Y(n_975) );
NOR2xp33_ASAP7_75t_L g976 ( .A(n_977), .B(n_980), .Y(n_976) );
NAND2xp5_ASAP7_75t_SL g980 ( .A(n_981), .B(n_983), .Y(n_980) );
AND4x1_ASAP7_75t_L g1034 ( .A(n_983), .B(n_1035), .C(n_1038), .D(n_1040), .Y(n_1034) );
NAND3xp33_ASAP7_75t_L g1098 ( .A(n_983), .B(n_1099), .C(n_1101), .Y(n_1098) );
NAND4xp25_ASAP7_75t_L g1531 ( .A(n_983), .B(n_1532), .C(n_1534), .D(n_1535), .Y(n_1531) );
INVx2_ASAP7_75t_L g986 ( .A(n_987), .Y(n_986) );
BUFx2_ASAP7_75t_L g991 ( .A(n_992), .Y(n_991) );
BUFx2_ASAP7_75t_L g1095 ( .A(n_992), .Y(n_1095) );
BUFx2_ASAP7_75t_L g1145 ( .A(n_992), .Y(n_1145) );
BUFx2_ASAP7_75t_L g1185 ( .A(n_992), .Y(n_1185) );
INVx1_ASAP7_75t_L g995 ( .A(n_996), .Y(n_995) );
NAND3xp33_ASAP7_75t_SL g1002 ( .A(n_1003), .B(n_1006), .C(n_1012), .Y(n_1002) );
AOI22xp33_ASAP7_75t_L g1196 ( .A1(n_1004), .A2(n_1197), .B1(n_1198), .B2(n_1199), .Y(n_1196) );
AOI22xp33_ASAP7_75t_L g1258 ( .A1(n_1004), .A2(n_1198), .B1(n_1259), .B2(n_1260), .Y(n_1258) );
INVx2_ASAP7_75t_L g1004 ( .A(n_1005), .Y(n_1004) );
INVx1_ASAP7_75t_SL g1010 ( .A(n_1011), .Y(n_1010) );
OAI221xp5_ASAP7_75t_L g1201 ( .A1(n_1018), .A2(n_1066), .B1(n_1202), .B2(n_1203), .C(n_1204), .Y(n_1201) );
INVx2_ASAP7_75t_L g1018 ( .A(n_1019), .Y(n_1018) );
INVx4_ASAP7_75t_L g1019 ( .A(n_1020), .Y(n_1019) );
INVx5_ASAP7_75t_L g1025 ( .A(n_1026), .Y(n_1025) );
INVx1_ASAP7_75t_L g1078 ( .A(n_1031), .Y(n_1078) );
HB1xp67_ASAP7_75t_L g1031 ( .A(n_1032), .Y(n_1031) );
XOR2xp5_ASAP7_75t_L g1032 ( .A(n_1033), .B(n_1077), .Y(n_1032) );
NAND3xp33_ASAP7_75t_L g1033 ( .A(n_1034), .B(n_1049), .C(n_1075), .Y(n_1033) );
NAND4xp25_ASAP7_75t_L g1050 ( .A(n_1051), .B(n_1056), .C(n_1059), .D(n_1060), .Y(n_1050) );
OAI211xp5_ASAP7_75t_L g1051 ( .A1(n_1052), .A2(n_1053), .B(n_1054), .C(n_1055), .Y(n_1051) );
OAI22xp5_ASAP7_75t_L g1067 ( .A1(n_1068), .A2(n_1069), .B1(n_1071), .B2(n_1072), .Y(n_1067) );
INVx1_ASAP7_75t_L g1069 ( .A(n_1070), .Y(n_1069) );
XNOR2xp5_ASAP7_75t_L g1079 ( .A(n_1080), .B(n_1219), .Y(n_1079) );
HB1xp67_ASAP7_75t_L g1080 ( .A(n_1081), .Y(n_1080) );
XNOR2xp5_ASAP7_75t_L g1081 ( .A(n_1082), .B(n_1167), .Y(n_1081) );
OAI22x1_ASAP7_75t_L g1082 ( .A1(n_1083), .A2(n_1084), .B1(n_1131), .B2(n_1166), .Y(n_1082) );
INVx2_ASAP7_75t_L g1083 ( .A(n_1084), .Y(n_1083) );
XNOR2x1_ASAP7_75t_L g1084 ( .A(n_1085), .B(n_1086), .Y(n_1084) );
AND3x2_ASAP7_75t_L g1086 ( .A(n_1087), .B(n_1104), .C(n_1129), .Y(n_1086) );
NOR2xp33_ASAP7_75t_SL g1087 ( .A(n_1088), .B(n_1098), .Y(n_1087) );
OAI21xp5_ASAP7_75t_SL g1088 ( .A1(n_1089), .A2(n_1092), .B(n_1094), .Y(n_1088) );
NAND3xp33_ASAP7_75t_L g1094 ( .A(n_1095), .B(n_1096), .C(n_1097), .Y(n_1094) );
INVx1_ASAP7_75t_L g1247 ( .A(n_1095), .Y(n_1247) );
AOI21xp5_ASAP7_75t_SL g1104 ( .A1(n_1105), .A2(n_1126), .B(n_1127), .Y(n_1104) );
NAND3xp33_ASAP7_75t_L g1105 ( .A(n_1106), .B(n_1109), .C(n_1116), .Y(n_1105) );
INVx2_ASAP7_75t_L g1111 ( .A(n_1112), .Y(n_1111) );
AOI31xp33_ASAP7_75t_L g1116 ( .A1(n_1117), .A2(n_1120), .A3(n_1121), .B(n_1124), .Y(n_1116) );
BUFx2_ASAP7_75t_L g1118 ( .A(n_1119), .Y(n_1118) );
INVx1_ASAP7_75t_L g1122 ( .A(n_1123), .Y(n_1122) );
INVx1_ASAP7_75t_L g1493 ( .A(n_1123), .Y(n_1493) );
O2A1O1Ixp5_ASAP7_75t_L g1186 ( .A1(n_1126), .A2(n_1187), .B(n_1200), .C(n_1213), .Y(n_1186) );
INVx1_ASAP7_75t_L g1166 ( .A(n_1131), .Y(n_1166) );
NAND3xp33_ASAP7_75t_L g1132 ( .A(n_1133), .B(n_1148), .C(n_1151), .Y(n_1132) );
NAND2xp5_ASAP7_75t_L g1134 ( .A(n_1135), .B(n_1138), .Y(n_1134) );
INVx2_ASAP7_75t_L g1141 ( .A(n_1142), .Y(n_1141) );
INVx2_ASAP7_75t_L g1395 ( .A(n_1144), .Y(n_1395) );
NAND2xp5_ASAP7_75t_L g1161 ( .A(n_1162), .B(n_1164), .Y(n_1161) );
XOR2x2_ASAP7_75t_L g1167 ( .A(n_1168), .B(n_1218), .Y(n_1167) );
NAND3x1_ASAP7_75t_SL g1168 ( .A(n_1169), .B(n_1186), .C(n_1216), .Y(n_1168) );
INVx1_ASAP7_75t_L g1228 ( .A(n_1173), .Y(n_1228) );
INVx1_ASAP7_75t_L g1179 ( .A(n_1180), .Y(n_1179) );
OAI22xp5_ASAP7_75t_L g1236 ( .A1(n_1180), .A2(n_1237), .B1(n_1239), .B2(n_1240), .Y(n_1236) );
OAI221xp5_ASAP7_75t_L g1888 ( .A1(n_1180), .A2(n_1283), .B1(n_1868), .B2(n_1889), .C(n_1890), .Y(n_1888) );
INVx1_ASAP7_75t_L g1400 ( .A(n_1185), .Y(n_1400) );
HB1xp67_ASAP7_75t_L g1192 ( .A(n_1193), .Y(n_1192) );
INVx1_ASAP7_75t_L g1194 ( .A(n_1195), .Y(n_1194) );
OAI22xp33_ASAP7_75t_L g1413 ( .A1(n_1202), .A2(n_1393), .B1(n_1399), .B2(n_1414), .Y(n_1413) );
OAI22xp5_ASAP7_75t_L g1205 ( .A1(n_1206), .A2(n_1207), .B1(n_1209), .B2(n_1212), .Y(n_1205) );
OAI221xp5_ASAP7_75t_SL g1250 ( .A1(n_1207), .A2(n_1209), .B1(n_1239), .B2(n_1245), .C(n_1251), .Y(n_1250) );
OAI221xp5_ASAP7_75t_L g1864 ( .A1(n_1207), .A2(n_1865), .B1(n_1866), .B2(n_1868), .C(n_1869), .Y(n_1864) );
OAI221xp5_ASAP7_75t_L g1872 ( .A1(n_1207), .A2(n_1873), .B1(n_1874), .B2(n_1875), .C(n_1876), .Y(n_1872) );
BUFx6f_ASAP7_75t_L g1207 ( .A(n_1208), .Y(n_1207) );
BUFx3_ASAP7_75t_L g1302 ( .A(n_1208), .Y(n_1302) );
INVx2_ASAP7_75t_SL g1415 ( .A(n_1208), .Y(n_1415) );
BUFx2_ASAP7_75t_L g1209 ( .A(n_1210), .Y(n_1209) );
BUFx6f_ASAP7_75t_L g1210 ( .A(n_1211), .Y(n_1210) );
AOI22xp5_ASAP7_75t_L g1219 ( .A1(n_1220), .A2(n_1221), .B1(n_1341), .B2(n_1342), .Y(n_1219) );
INVx1_ASAP7_75t_L g1220 ( .A(n_1221), .Y(n_1220) );
AOI22xp5_ASAP7_75t_L g1221 ( .A1(n_1222), .A2(n_1223), .B1(n_1264), .B2(n_1340), .Y(n_1221) );
INVx1_ASAP7_75t_L g1222 ( .A(n_1223), .Y(n_1222) );
XNOR2xp5_ASAP7_75t_SL g1223 ( .A(n_1224), .B(n_1225), .Y(n_1223) );
AND3x2_ASAP7_75t_L g1225 ( .A(n_1226), .B(n_1248), .C(n_1261), .Y(n_1225) );
OAI22xp33_ASAP7_75t_L g1244 ( .A1(n_1234), .A2(n_1237), .B1(n_1245), .B2(n_1246), .Y(n_1244) );
OAI22xp33_ASAP7_75t_L g1824 ( .A1(n_1234), .A2(n_1825), .B1(n_1826), .B2(n_1828), .Y(n_1824) );
OAI22xp33_ASAP7_75t_L g1886 ( .A1(n_1234), .A2(n_1826), .B1(n_1873), .B2(n_1887), .Y(n_1886) );
INVx1_ASAP7_75t_L g1237 ( .A(n_1238), .Y(n_1237) );
INVx1_ASAP7_75t_L g1340 ( .A(n_1264), .Y(n_1340) );
HB1xp67_ASAP7_75t_L g1264 ( .A(n_1265), .Y(n_1264) );
XNOR2x1_ASAP7_75t_L g1265 ( .A(n_1266), .B(n_1311), .Y(n_1265) );
NAND4xp75_ASAP7_75t_L g1267 ( .A(n_1268), .B(n_1273), .C(n_1290), .D(n_1309), .Y(n_1267) );
OAI221xp5_ASAP7_75t_L g1280 ( .A1(n_1281), .A2(n_1282), .B1(n_1283), .B2(n_1284), .C(n_1285), .Y(n_1280) );
OAI221xp5_ASAP7_75t_L g1829 ( .A1(n_1283), .A2(n_1830), .B1(n_1831), .B2(n_1832), .C(n_1833), .Y(n_1829) );
INVx1_ASAP7_75t_L g1288 ( .A(n_1289), .Y(n_1288) );
OAI21xp5_ASAP7_75t_L g1290 ( .A1(n_1291), .A2(n_1299), .B(n_1308), .Y(n_1290) );
NAND2xp5_ASAP7_75t_L g1291 ( .A(n_1292), .B(n_1296), .Y(n_1291) );
OAI221xp5_ASAP7_75t_L g1301 ( .A1(n_1302), .A2(n_1303), .B1(n_1304), .B2(n_1306), .C(n_1307), .Y(n_1301) );
BUFx3_ASAP7_75t_L g1304 ( .A(n_1305), .Y(n_1304) );
AND2x2_ASAP7_75t_L g1312 ( .A(n_1313), .B(n_1327), .Y(n_1312) );
AOI22xp5_ASAP7_75t_L g1320 ( .A1(n_1321), .A2(n_1323), .B1(n_1324), .B2(n_1326), .Y(n_1320) );
NAND3xp33_ASAP7_75t_L g1328 ( .A(n_1329), .B(n_1332), .C(n_1335), .Y(n_1328) );
INVx1_ASAP7_75t_L g1341 ( .A(n_1342), .Y(n_1341) );
AO22x2_ASAP7_75t_L g1342 ( .A1(n_1343), .A2(n_1484), .B1(n_1572), .B2(n_1573), .Y(n_1342) );
INVx1_ASAP7_75t_L g1572 ( .A(n_1343), .Y(n_1572) );
XNOR2xp5_ASAP7_75t_L g1343 ( .A(n_1344), .B(n_1380), .Y(n_1343) );
INVx1_ASAP7_75t_L g1344 ( .A(n_1345), .Y(n_1344) );
NAND3xp33_ASAP7_75t_L g1346 ( .A(n_1347), .B(n_1365), .C(n_1368), .Y(n_1346) );
INVx1_ASAP7_75t_L g1358 ( .A(n_1359), .Y(n_1358) );
NAND2xp5_ASAP7_75t_L g1369 ( .A(n_1370), .B(n_1372), .Y(n_1369) );
NAND3xp33_ASAP7_75t_L g1381 ( .A(n_1382), .B(n_1421), .C(n_1451), .Y(n_1381) );
NOR2xp33_ASAP7_75t_L g1382 ( .A(n_1383), .B(n_1404), .Y(n_1382) );
OAI33xp33_ASAP7_75t_L g1383 ( .A1(n_1384), .A2(n_1385), .A3(n_1390), .B1(n_1394), .B2(n_1400), .B3(n_1401), .Y(n_1383) );
OAI22xp33_ASAP7_75t_L g1385 ( .A1(n_1386), .A2(n_1387), .B1(n_1388), .B2(n_1389), .Y(n_1385) );
OAI22xp5_ASAP7_75t_L g1406 ( .A1(n_1386), .A2(n_1402), .B1(n_1407), .B2(n_1409), .Y(n_1406) );
OAI22xp5_ASAP7_75t_L g1394 ( .A1(n_1395), .A2(n_1396), .B1(n_1397), .B2(n_1399), .Y(n_1394) );
BUFx6f_ASAP7_75t_L g1397 ( .A(n_1398), .Y(n_1397) );
INVx2_ASAP7_75t_L g1461 ( .A(n_1398), .Y(n_1461) );
OAI33xp33_ASAP7_75t_L g1404 ( .A1(n_1405), .A2(n_1406), .A3(n_1411), .B1(n_1412), .B2(n_1413), .B3(n_1416), .Y(n_1404) );
INVx2_ASAP7_75t_L g1407 ( .A(n_1408), .Y(n_1407) );
INVx2_ASAP7_75t_L g1409 ( .A(n_1410), .Y(n_1409) );
INVx2_ASAP7_75t_L g1414 ( .A(n_1415), .Y(n_1414) );
INVx2_ASAP7_75t_L g1416 ( .A(n_1417), .Y(n_1416) );
INVx1_ASAP7_75t_L g1417 ( .A(n_1418), .Y(n_1417) );
INVx1_ASAP7_75t_L g1419 ( .A(n_1420), .Y(n_1419) );
OAI31xp33_ASAP7_75t_SL g1421 ( .A1(n_1422), .A2(n_1434), .A3(n_1444), .B(n_1448), .Y(n_1421) );
INVx1_ASAP7_75t_L g1423 ( .A(n_1424), .Y(n_1423) );
AOI22xp33_ASAP7_75t_L g1426 ( .A1(n_1427), .A2(n_1430), .B1(n_1431), .B2(n_1432), .Y(n_1426) );
BUFx3_ASAP7_75t_L g1427 ( .A(n_1428), .Y(n_1427) );
AOI22xp33_ASAP7_75t_L g1464 ( .A1(n_1430), .A2(n_1465), .B1(n_1469), .B2(n_1472), .Y(n_1464) );
BUFx3_ASAP7_75t_L g1432 ( .A(n_1433), .Y(n_1432) );
INVx1_ASAP7_75t_L g1435 ( .A(n_1436), .Y(n_1435) );
INVx1_ASAP7_75t_L g1436 ( .A(n_1437), .Y(n_1436) );
INVx2_ASAP7_75t_L g1439 ( .A(n_1440), .Y(n_1439) );
INVx2_ASAP7_75t_L g1440 ( .A(n_1441), .Y(n_1440) );
INVx2_ASAP7_75t_L g1441 ( .A(n_1442), .Y(n_1441) );
INVx1_ASAP7_75t_L g1442 ( .A(n_1443), .Y(n_1442) );
INVx3_ASAP7_75t_SL g1446 ( .A(n_1447), .Y(n_1446) );
BUFx3_ASAP7_75t_L g1448 ( .A(n_1449), .Y(n_1448) );
OAI31xp33_ASAP7_75t_SL g1451 ( .A1(n_1452), .A2(n_1459), .A3(n_1473), .B(n_1479), .Y(n_1451) );
INVx1_ASAP7_75t_L g1453 ( .A(n_1454), .Y(n_1453) );
INVx1_ASAP7_75t_L g1454 ( .A(n_1455), .Y(n_1454) );
INVx1_ASAP7_75t_L g1456 ( .A(n_1457), .Y(n_1456) );
INVx2_ASAP7_75t_L g1460 ( .A(n_1461), .Y(n_1460) );
CKINVDCx8_ASAP7_75t_R g1462 ( .A(n_1463), .Y(n_1462) );
BUFx3_ASAP7_75t_L g1465 ( .A(n_1466), .Y(n_1465) );
AND2x2_ASAP7_75t_L g1466 ( .A(n_1467), .B(n_1468), .Y(n_1466) );
AND2x4_ASAP7_75t_L g1470 ( .A(n_1467), .B(n_1471), .Y(n_1470) );
BUFx6f_ASAP7_75t_L g1469 ( .A(n_1470), .Y(n_1469) );
INVx1_ASAP7_75t_L g1474 ( .A(n_1475), .Y(n_1474) );
INVx2_ASAP7_75t_SL g1475 ( .A(n_1476), .Y(n_1475) );
BUFx3_ASAP7_75t_L g1477 ( .A(n_1478), .Y(n_1477) );
AND2x2_ASAP7_75t_L g1479 ( .A(n_1480), .B(n_1482), .Y(n_1479) );
INVx1_ASAP7_75t_SL g1480 ( .A(n_1481), .Y(n_1480) );
INVx1_ASAP7_75t_L g1482 ( .A(n_1483), .Y(n_1482) );
INVx1_ASAP7_75t_L g1573 ( .A(n_1484), .Y(n_1573) );
AOI22xp5_ASAP7_75t_L g1484 ( .A1(n_1485), .A2(n_1486), .B1(n_1537), .B2(n_1571), .Y(n_1484) );
INVx1_ASAP7_75t_L g1485 ( .A(n_1486), .Y(n_1485) );
NOR3xp33_ASAP7_75t_L g1487 ( .A(n_1488), .B(n_1531), .C(n_1536), .Y(n_1487) );
NAND2xp5_ASAP7_75t_L g1488 ( .A(n_1489), .B(n_1505), .Y(n_1488) );
NAND2xp5_ASAP7_75t_L g1491 ( .A(n_1492), .B(n_1494), .Y(n_1491) );
NAND3xp33_ASAP7_75t_L g1495 ( .A(n_1496), .B(n_1500), .C(n_1503), .Y(n_1495) );
AOI21xp5_ASAP7_75t_L g1505 ( .A1(n_1506), .A2(n_1507), .B(n_1508), .Y(n_1505) );
AOI21xp5_ASAP7_75t_SL g1880 ( .A1(n_1506), .A2(n_1881), .B(n_1882), .Y(n_1880) );
OAI22xp5_ASAP7_75t_L g1509 ( .A1(n_1510), .A2(n_1511), .B1(n_1512), .B2(n_1513), .Y(n_1509) );
INVx1_ASAP7_75t_L g1513 ( .A(n_1514), .Y(n_1513) );
OAI22xp33_ASAP7_75t_L g1515 ( .A1(n_1516), .A2(n_1517), .B1(n_1518), .B2(n_1519), .Y(n_1515) );
INVx1_ASAP7_75t_L g1519 ( .A(n_1520), .Y(n_1519) );
OAI22xp5_ASAP7_75t_L g1525 ( .A1(n_1526), .A2(n_1527), .B1(n_1528), .B2(n_1530), .Y(n_1525) );
INVx1_ASAP7_75t_L g1528 ( .A(n_1529), .Y(n_1528) );
INVx1_ASAP7_75t_L g1571 ( .A(n_1537), .Y(n_1571) );
INVx1_ASAP7_75t_L g1570 ( .A(n_1538), .Y(n_1570) );
NAND3xp33_ASAP7_75t_L g1538 ( .A(n_1539), .B(n_1555), .C(n_1558), .Y(n_1538) );
NAND2xp5_ASAP7_75t_L g1559 ( .A(n_1560), .B(n_1562), .Y(n_1559) );
OAI221xp5_ASAP7_75t_SL g1574 ( .A1(n_1575), .A2(n_1792), .B1(n_1795), .B2(n_1839), .C(n_1845), .Y(n_1574) );
AOI211xp5_ASAP7_75t_L g1575 ( .A1(n_1576), .A2(n_1592), .B(n_1674), .C(n_1786), .Y(n_1575) );
NAND2xp5_ASAP7_75t_L g1726 ( .A(n_1576), .B(n_1727), .Y(n_1726) );
INVx1_ASAP7_75t_L g1777 ( .A(n_1576), .Y(n_1777) );
INVx1_ASAP7_75t_L g1576 ( .A(n_1577), .Y(n_1576) );
NAND3xp33_ASAP7_75t_L g1768 ( .A(n_1577), .B(n_1630), .C(n_1712), .Y(n_1768) );
AND2x2_ASAP7_75t_L g1785 ( .A(n_1577), .B(n_1728), .Y(n_1785) );
INVx1_ASAP7_75t_L g1577 ( .A(n_1578), .Y(n_1577) );
AOI32xp33_ASAP7_75t_L g1694 ( .A1(n_1578), .A2(n_1622), .A3(n_1664), .B1(n_1695), .B2(n_1697), .Y(n_1694) );
INVx1_ASAP7_75t_L g1698 ( .A(n_1578), .Y(n_1698) );
NOR2xp33_ASAP7_75t_L g1709 ( .A(n_1578), .B(n_1604), .Y(n_1709) );
AOI211xp5_ASAP7_75t_L g1710 ( .A1(n_1578), .A2(n_1711), .B(n_1712), .C(n_1716), .Y(n_1710) );
AND2x2_ASAP7_75t_L g1578 ( .A(n_1579), .B(n_1586), .Y(n_1578) );
AND2x6_ASAP7_75t_L g1580 ( .A(n_1581), .B(n_1582), .Y(n_1580) );
AND2x2_ASAP7_75t_L g1584 ( .A(n_1581), .B(n_1585), .Y(n_1584) );
AND2x4_ASAP7_75t_L g1587 ( .A(n_1581), .B(n_1588), .Y(n_1587) );
AND2x6_ASAP7_75t_L g1590 ( .A(n_1581), .B(n_1591), .Y(n_1590) );
AND2x2_ASAP7_75t_L g1606 ( .A(n_1581), .B(n_1585), .Y(n_1606) );
AND2x2_ASAP7_75t_L g1620 ( .A(n_1581), .B(n_1585), .Y(n_1620) );
AND2x2_ASAP7_75t_L g1588 ( .A(n_1583), .B(n_1589), .Y(n_1588) );
INVx2_ASAP7_75t_L g1794 ( .A(n_1590), .Y(n_1794) );
HB1xp67_ASAP7_75t_L g1893 ( .A(n_1591), .Y(n_1893) );
NAND5xp2_ASAP7_75t_L g1592 ( .A(n_1593), .B(n_1652), .C(n_1662), .D(n_1667), .E(n_1670), .Y(n_1592) );
AOI221xp5_ASAP7_75t_SL g1593 ( .A1(n_1594), .A2(n_1608), .B1(n_1615), .B2(n_1630), .C(n_1632), .Y(n_1593) );
O2A1O1Ixp33_ASAP7_75t_L g1753 ( .A1(n_1594), .A2(n_1696), .B(n_1754), .C(n_1756), .Y(n_1753) );
INVx1_ASAP7_75t_L g1594 ( .A(n_1595), .Y(n_1594) );
OR2x2_ASAP7_75t_L g1595 ( .A(n_1596), .B(n_1600), .Y(n_1595) );
NOR3xp33_ASAP7_75t_L g1737 ( .A(n_1596), .B(n_1704), .C(n_1738), .Y(n_1737) );
AND2x2_ASAP7_75t_L g1741 ( .A(n_1596), .B(n_1604), .Y(n_1741) );
OAI31xp33_ASAP7_75t_L g1772 ( .A1(n_1596), .A2(n_1651), .A3(n_1773), .B(n_1775), .Y(n_1772) );
INVx3_ASAP7_75t_L g1596 ( .A(n_1597), .Y(n_1596) );
NAND2xp5_ASAP7_75t_L g1631 ( .A(n_1597), .B(n_1604), .Y(n_1631) );
AND2x2_ASAP7_75t_L g1634 ( .A(n_1597), .B(n_1635), .Y(n_1634) );
AND2x2_ASAP7_75t_L g1641 ( .A(n_1597), .B(n_1642), .Y(n_1641) );
AND2x2_ASAP7_75t_L g1653 ( .A(n_1597), .B(n_1654), .Y(n_1653) );
INVx3_ASAP7_75t_L g1728 ( .A(n_1597), .Y(n_1728) );
AND2x2_ASAP7_75t_L g1734 ( .A(n_1597), .B(n_1716), .Y(n_1734) );
OR2x2_ASAP7_75t_L g1746 ( .A(n_1597), .B(n_1604), .Y(n_1746) );
AND2x2_ASAP7_75t_L g1749 ( .A(n_1597), .B(n_1698), .Y(n_1749) );
AND2x2_ASAP7_75t_L g1771 ( .A(n_1597), .B(n_1759), .Y(n_1771) );
AND2x4_ASAP7_75t_SL g1597 ( .A(n_1598), .B(n_1599), .Y(n_1597) );
INVx1_ASAP7_75t_L g1686 ( .A(n_1600), .Y(n_1686) );
OR2x2_ASAP7_75t_L g1600 ( .A(n_1601), .B(n_1604), .Y(n_1600) );
INVx1_ASAP7_75t_L g1635 ( .A(n_1601), .Y(n_1635) );
AND2x2_ASAP7_75t_L g1642 ( .A(n_1601), .B(n_1604), .Y(n_1642) );
INVx1_ASAP7_75t_L g1656 ( .A(n_1601), .Y(n_1656) );
INVx1_ASAP7_75t_L g1711 ( .A(n_1601), .Y(n_1711) );
NAND2xp5_ASAP7_75t_L g1601 ( .A(n_1602), .B(n_1603), .Y(n_1601) );
OR2x2_ASAP7_75t_L g1655 ( .A(n_1604), .B(n_1656), .Y(n_1655) );
AND2x2_ASAP7_75t_L g1604 ( .A(n_1605), .B(n_1607), .Y(n_1604) );
AND2x4_ASAP7_75t_L g1664 ( .A(n_1605), .B(n_1607), .Y(n_1664) );
AND2x2_ASAP7_75t_L g1650 ( .A(n_1608), .B(n_1618), .Y(n_1650) );
AND2x2_ASAP7_75t_L g1668 ( .A(n_1608), .B(n_1669), .Y(n_1668) );
AND2x2_ASAP7_75t_L g1682 ( .A(n_1608), .B(n_1617), .Y(n_1682) );
INVx1_ASAP7_75t_L g1774 ( .A(n_1608), .Y(n_1774) );
AND2x2_ASAP7_75t_L g1608 ( .A(n_1609), .B(n_1612), .Y(n_1608) );
INVx1_ASAP7_75t_L g1625 ( .A(n_1609), .Y(n_1625) );
INVx1_ASAP7_75t_L g1765 ( .A(n_1609), .Y(n_1765) );
NAND2xp5_ASAP7_75t_L g1609 ( .A(n_1610), .B(n_1611), .Y(n_1609) );
OR2x2_ASAP7_75t_L g1624 ( .A(n_1612), .B(n_1625), .Y(n_1624) );
INVx1_ASAP7_75t_L g1639 ( .A(n_1612), .Y(n_1639) );
INVx1_ASAP7_75t_L g1648 ( .A(n_1612), .Y(n_1648) );
AND2x2_ASAP7_75t_L g1660 ( .A(n_1612), .B(n_1625), .Y(n_1660) );
NAND2xp5_ASAP7_75t_L g1612 ( .A(n_1613), .B(n_1614), .Y(n_1612) );
INVx1_ASAP7_75t_L g1615 ( .A(n_1616), .Y(n_1615) );
AOI221xp5_ASAP7_75t_SL g1786 ( .A1(n_1616), .A2(n_1663), .B1(n_1686), .B2(n_1787), .C(n_1791), .Y(n_1786) );
OR2x2_ASAP7_75t_L g1616 ( .A(n_1617), .B(n_1622), .Y(n_1616) );
AND2x2_ASAP7_75t_L g1696 ( .A(n_1617), .B(n_1623), .Y(n_1696) );
AND2x2_ASAP7_75t_L g1701 ( .A(n_1617), .B(n_1657), .Y(n_1701) );
AND2x2_ASAP7_75t_L g1714 ( .A(n_1617), .B(n_1715), .Y(n_1714) );
AND2x2_ASAP7_75t_L g1720 ( .A(n_1617), .B(n_1647), .Y(n_1720) );
AND2x2_ASAP7_75t_L g1781 ( .A(n_1617), .B(n_1765), .Y(n_1781) );
CKINVDCx5p33_ASAP7_75t_R g1617 ( .A(n_1618), .Y(n_1617) );
AND2x2_ASAP7_75t_L g1637 ( .A(n_1618), .B(n_1638), .Y(n_1637) );
NOR2xp33_ASAP7_75t_L g1666 ( .A(n_1618), .B(n_1627), .Y(n_1666) );
AND2x2_ASAP7_75t_L g1669 ( .A(n_1618), .B(n_1627), .Y(n_1669) );
AND2x2_ASAP7_75t_L g1671 ( .A(n_1618), .B(n_1648), .Y(n_1671) );
OR2x2_ASAP7_75t_L g1755 ( .A(n_1618), .B(n_1639), .Y(n_1755) );
NAND2xp5_ASAP7_75t_L g1764 ( .A(n_1618), .B(n_1765), .Y(n_1764) );
AND2x2_ASAP7_75t_L g1618 ( .A(n_1619), .B(n_1621), .Y(n_1618) );
AND2x2_ASAP7_75t_L g1685 ( .A(n_1619), .B(n_1621), .Y(n_1685) );
NAND2xp5_ASAP7_75t_SL g1622 ( .A(n_1623), .B(n_1626), .Y(n_1622) );
AND2x2_ASAP7_75t_L g1684 ( .A(n_1623), .B(n_1685), .Y(n_1684) );
INVx1_ASAP7_75t_L g1623 ( .A(n_1624), .Y(n_1623) );
NOR2xp33_ASAP7_75t_L g1657 ( .A(n_1624), .B(n_1646), .Y(n_1657) );
AND2x2_ASAP7_75t_L g1647 ( .A(n_1625), .B(n_1648), .Y(n_1647) );
INVx1_ASAP7_75t_L g1715 ( .A(n_1625), .Y(n_1715) );
OAI322xp33_ASAP7_75t_L g1632 ( .A1(n_1626), .A2(n_1633), .A3(n_1636), .B1(n_1640), .B2(n_1643), .C1(n_1649), .C2(n_1651), .Y(n_1632) );
NAND2xp5_ASAP7_75t_L g1649 ( .A(n_1626), .B(n_1650), .Y(n_1649) );
OR2x2_ASAP7_75t_L g1680 ( .A(n_1626), .B(n_1681), .Y(n_1680) );
INVx2_ASAP7_75t_L g1725 ( .A(n_1626), .Y(n_1725) );
NAND2xp5_ASAP7_75t_L g1736 ( .A(n_1626), .B(n_1671), .Y(n_1736) );
INVx2_ASAP7_75t_L g1626 ( .A(n_1627), .Y(n_1626) );
INVx3_ASAP7_75t_L g1646 ( .A(n_1627), .Y(n_1646) );
OR2x2_ASAP7_75t_L g1704 ( .A(n_1627), .B(n_1656), .Y(n_1704) );
AND2x2_ASAP7_75t_L g1627 ( .A(n_1628), .B(n_1629), .Y(n_1627) );
INVx1_ASAP7_75t_L g1630 ( .A(n_1631), .Y(n_1630) );
NOR2xp33_ASAP7_75t_L g1756 ( .A(n_1631), .B(n_1757), .Y(n_1756) );
A2O1A1Ixp33_ASAP7_75t_SL g1729 ( .A1(n_1633), .A2(n_1730), .B(n_1731), .C(n_1733), .Y(n_1729) );
OAI221xp5_ASAP7_75t_L g1769 ( .A1(n_1633), .A2(n_1665), .B1(n_1751), .B2(n_1770), .C(n_1772), .Y(n_1769) );
INVx1_ASAP7_75t_L g1633 ( .A(n_1634), .Y(n_1633) );
INVx1_ASAP7_75t_L g1678 ( .A(n_1635), .Y(n_1678) );
NAND2xp5_ASAP7_75t_L g1688 ( .A(n_1635), .B(n_1665), .Y(n_1688) );
NAND2xp5_ASAP7_75t_L g1700 ( .A(n_1635), .B(n_1701), .Y(n_1700) );
INVx1_ASAP7_75t_L g1723 ( .A(n_1635), .Y(n_1723) );
INVx1_ASAP7_75t_L g1636 ( .A(n_1637), .Y(n_1636) );
OAI22xp5_ASAP7_75t_SL g1747 ( .A1(n_1638), .A2(n_1748), .B1(n_1750), .B2(n_1752), .Y(n_1747) );
INVx1_ASAP7_75t_L g1638 ( .A(n_1639), .Y(n_1638) );
INVx1_ASAP7_75t_L g1640 ( .A(n_1641), .Y(n_1640) );
CKINVDCx14_ASAP7_75t_R g1651 ( .A(n_1642), .Y(n_1651) );
AOI22xp5_ASAP7_75t_L g1717 ( .A1(n_1642), .A2(n_1718), .B1(n_1723), .B2(n_1724), .Y(n_1717) );
INVx1_ASAP7_75t_L g1643 ( .A(n_1644), .Y(n_1643) );
AOI321xp33_ASAP7_75t_L g1776 ( .A1(n_1644), .A2(n_1650), .A3(n_1745), .B1(n_1777), .B2(n_1778), .C(n_1779), .Y(n_1776) );
AND2x2_ASAP7_75t_L g1644 ( .A(n_1645), .B(n_1647), .Y(n_1644) );
NAND2xp5_ASAP7_75t_L g1707 ( .A(n_1645), .B(n_1660), .Y(n_1707) );
AOI21xp33_ASAP7_75t_L g1778 ( .A1(n_1645), .A2(n_1655), .B(n_1727), .Y(n_1778) );
AND2x2_ASAP7_75t_L g1783 ( .A(n_1645), .B(n_1678), .Y(n_1783) );
INVx1_ASAP7_75t_L g1645 ( .A(n_1646), .Y(n_1645) );
NAND2xp5_ASAP7_75t_L g1661 ( .A(n_1646), .B(n_1654), .Y(n_1661) );
NAND2xp5_ASAP7_75t_L g1673 ( .A(n_1646), .B(n_1656), .Y(n_1673) );
NAND2xp5_ASAP7_75t_L g1713 ( .A(n_1646), .B(n_1714), .Y(n_1713) );
AND2x2_ASAP7_75t_L g1722 ( .A(n_1646), .B(n_1660), .Y(n_1722) );
NOR2xp33_ASAP7_75t_L g1754 ( .A(n_1646), .B(n_1755), .Y(n_1754) );
AND2x2_ASAP7_75t_L g1693 ( .A(n_1647), .B(n_1685), .Y(n_1693) );
INVx1_ASAP7_75t_L g1738 ( .A(n_1647), .Y(n_1738) );
AND2x2_ASAP7_75t_L g1751 ( .A(n_1647), .B(n_1666), .Y(n_1751) );
AOI211xp5_ASAP7_75t_L g1702 ( .A1(n_1650), .A2(n_1703), .B(n_1705), .C(n_1708), .Y(n_1702) );
NAND2xp5_ASAP7_75t_L g1791 ( .A(n_1650), .B(n_1785), .Y(n_1791) );
AOI21xp5_ASAP7_75t_L g1652 ( .A1(n_1653), .A2(n_1657), .B(n_1658), .Y(n_1652) );
INVx2_ASAP7_75t_SL g1654 ( .A(n_1655), .Y(n_1654) );
OAI22xp5_ASAP7_75t_L g1787 ( .A1(n_1655), .A2(n_1716), .B1(n_1788), .B2(n_1790), .Y(n_1787) );
AND2x2_ASAP7_75t_L g1663 ( .A(n_1656), .B(n_1664), .Y(n_1663) );
INVx1_ASAP7_75t_L g1730 ( .A(n_1657), .Y(n_1730) );
NOR2xp33_ASAP7_75t_L g1658 ( .A(n_1659), .B(n_1661), .Y(n_1658) );
OR2x2_ASAP7_75t_L g1691 ( .A(n_1659), .B(n_1685), .Y(n_1691) );
INVx1_ASAP7_75t_L g1659 ( .A(n_1660), .Y(n_1659) );
AND2x2_ASAP7_75t_L g1665 ( .A(n_1660), .B(n_1666), .Y(n_1665) );
AND2x2_ASAP7_75t_L g1744 ( .A(n_1660), .B(n_1669), .Y(n_1744) );
AOI211xp5_ASAP7_75t_L g1763 ( .A1(n_1661), .A2(n_1727), .B(n_1764), .C(n_1766), .Y(n_1763) );
NAND2xp5_ASAP7_75t_L g1662 ( .A(n_1663), .B(n_1665), .Y(n_1662) );
NAND2xp5_ASAP7_75t_L g1667 ( .A(n_1663), .B(n_1668), .Y(n_1667) );
AOI21xp5_ASAP7_75t_L g1689 ( .A1(n_1663), .A2(n_1690), .B(n_1694), .Y(n_1689) );
NAND3xp33_ASAP7_75t_L g1748 ( .A(n_1663), .B(n_1725), .C(n_1749), .Y(n_1748) );
NOR2xp33_ASAP7_75t_L g1697 ( .A(n_1664), .B(n_1698), .Y(n_1697) );
INVx2_ASAP7_75t_L g1716 ( .A(n_1664), .Y(n_1716) );
NAND2xp5_ASAP7_75t_L g1757 ( .A(n_1668), .B(n_1758), .Y(n_1757) );
CKINVDCx14_ASAP7_75t_R g1775 ( .A(n_1669), .Y(n_1775) );
NAND2xp5_ASAP7_75t_L g1670 ( .A(n_1671), .B(n_1672), .Y(n_1670) );
INVx1_ASAP7_75t_L g1672 ( .A(n_1673), .Y(n_1672) );
NAND5xp2_ASAP7_75t_L g1674 ( .A(n_1675), .B(n_1753), .C(n_1760), .D(n_1769), .E(n_1776), .Y(n_1674) );
AOI321xp33_ASAP7_75t_SL g1675 ( .A1(n_1676), .A2(n_1698), .A3(n_1699), .B1(n_1726), .B2(n_1729), .C(n_1739), .Y(n_1675) );
NAND3xp33_ASAP7_75t_SL g1676 ( .A(n_1677), .B(n_1683), .C(n_1689), .Y(n_1676) );
INVxp67_ASAP7_75t_L g1790 ( .A(n_1677), .Y(n_1790) );
NAND2xp5_ASAP7_75t_L g1677 ( .A(n_1678), .B(n_1679), .Y(n_1677) );
NAND2xp5_ASAP7_75t_L g1789 ( .A(n_1678), .B(n_1705), .Y(n_1789) );
INVx1_ASAP7_75t_L g1679 ( .A(n_1680), .Y(n_1679) );
A2O1A1Ixp33_ASAP7_75t_L g1739 ( .A1(n_1680), .A2(n_1688), .B(n_1740), .C(n_1742), .Y(n_1739) );
INVx1_ASAP7_75t_L g1681 ( .A(n_1682), .Y(n_1681) );
AOI21xp5_ASAP7_75t_L g1683 ( .A1(n_1684), .A2(n_1686), .B(n_1687), .Y(n_1683) );
OR2x2_ASAP7_75t_L g1706 ( .A(n_1685), .B(n_1707), .Y(n_1706) );
AND2x2_ASAP7_75t_L g1732 ( .A(n_1685), .B(n_1722), .Y(n_1732) );
INVx1_ASAP7_75t_L g1687 ( .A(n_1688), .Y(n_1687) );
NAND2xp5_ASAP7_75t_L g1690 ( .A(n_1691), .B(n_1692), .Y(n_1690) );
INVx1_ASAP7_75t_L g1761 ( .A(n_1691), .Y(n_1761) );
INVx1_ASAP7_75t_L g1692 ( .A(n_1693), .Y(n_1692) );
INVx1_ASAP7_75t_L g1695 ( .A(n_1696), .Y(n_1695) );
A2O1A1Ixp33_ASAP7_75t_L g1699 ( .A1(n_1700), .A2(n_1702), .B(n_1710), .C(n_1717), .Y(n_1699) );
CKINVDCx14_ASAP7_75t_R g1703 ( .A(n_1704), .Y(n_1703) );
INVx1_ASAP7_75t_L g1705 ( .A(n_1706), .Y(n_1705) );
INVx1_ASAP7_75t_L g1708 ( .A(n_1709), .Y(n_1708) );
AND2x2_ASAP7_75t_L g1743 ( .A(n_1711), .B(n_1744), .Y(n_1743) );
INVx1_ASAP7_75t_L g1759 ( .A(n_1711), .Y(n_1759) );
INVx1_ASAP7_75t_L g1712 ( .A(n_1713), .Y(n_1712) );
INVx1_ASAP7_75t_L g1766 ( .A(n_1714), .Y(n_1766) );
NAND2xp5_ASAP7_75t_L g1718 ( .A(n_1719), .B(n_1721), .Y(n_1718) );
INVx1_ASAP7_75t_L g1719 ( .A(n_1720), .Y(n_1719) );
AND2x2_ASAP7_75t_L g1724 ( .A(n_1720), .B(n_1725), .Y(n_1724) );
INVx1_ASAP7_75t_L g1721 ( .A(n_1722), .Y(n_1721) );
AOI311xp33_ASAP7_75t_L g1760 ( .A1(n_1723), .A2(n_1761), .A3(n_1762), .B(n_1763), .C(n_1767), .Y(n_1760) );
INVxp67_ASAP7_75t_SL g1762 ( .A(n_1726), .Y(n_1762) );
INVx2_ASAP7_75t_L g1727 ( .A(n_1728), .Y(n_1727) );
CKINVDCx14_ASAP7_75t_R g1731 ( .A(n_1732), .Y(n_1731) );
AOI21xp5_ASAP7_75t_L g1733 ( .A1(n_1734), .A2(n_1735), .B(n_1737), .Y(n_1733) );
INVx1_ASAP7_75t_L g1752 ( .A(n_1734), .Y(n_1752) );
INVx1_ASAP7_75t_L g1735 ( .A(n_1736), .Y(n_1735) );
NAND2xp5_ASAP7_75t_L g1773 ( .A(n_1738), .B(n_1774), .Y(n_1773) );
AOI211xp5_ASAP7_75t_L g1779 ( .A1(n_1738), .A2(n_1780), .B(n_1782), .C(n_1784), .Y(n_1779) );
INVx1_ASAP7_75t_L g1740 ( .A(n_1741), .Y(n_1740) );
AOI21xp5_ASAP7_75t_L g1742 ( .A1(n_1743), .A2(n_1745), .B(n_1747), .Y(n_1742) );
INVx1_ASAP7_75t_L g1745 ( .A(n_1746), .Y(n_1745) );
INVx1_ASAP7_75t_L g1750 ( .A(n_1751), .Y(n_1750) );
INVx1_ASAP7_75t_L g1758 ( .A(n_1759), .Y(n_1758) );
INVxp67_ASAP7_75t_SL g1767 ( .A(n_1768), .Y(n_1767) );
INVx1_ASAP7_75t_L g1770 ( .A(n_1771), .Y(n_1770) );
INVx1_ASAP7_75t_L g1780 ( .A(n_1781), .Y(n_1780) );
INVxp67_ASAP7_75t_L g1782 ( .A(n_1783), .Y(n_1782) );
INVx1_ASAP7_75t_L g1784 ( .A(n_1785), .Y(n_1784) );
INVxp67_ASAP7_75t_L g1788 ( .A(n_1789), .Y(n_1788) );
CKINVDCx20_ASAP7_75t_R g1792 ( .A(n_1793), .Y(n_1792) );
CKINVDCx20_ASAP7_75t_R g1793 ( .A(n_1794), .Y(n_1793) );
INVx1_ASAP7_75t_L g1795 ( .A(n_1796), .Y(n_1795) );
XNOR2x1_ASAP7_75t_L g1796 ( .A(n_1797), .B(n_1798), .Y(n_1796) );
AND2x2_ASAP7_75t_L g1798 ( .A(n_1799), .B(n_1835), .Y(n_1798) );
NAND3xp33_ASAP7_75t_L g1801 ( .A(n_1802), .B(n_1808), .C(n_1815), .Y(n_1801) );
INVx1_ASAP7_75t_L g1811 ( .A(n_1812), .Y(n_1811) );
INVx1_ASAP7_75t_L g1821 ( .A(n_1822), .Y(n_1821) );
INVx2_ASAP7_75t_L g1826 ( .A(n_1827), .Y(n_1826) );
CKINVDCx20_ASAP7_75t_R g1839 ( .A(n_1840), .Y(n_1839) );
CKINVDCx20_ASAP7_75t_R g1840 ( .A(n_1841), .Y(n_1840) );
INVx3_ASAP7_75t_L g1841 ( .A(n_1842), .Y(n_1841) );
BUFx3_ASAP7_75t_L g1842 ( .A(n_1843), .Y(n_1842) );
BUFx3_ASAP7_75t_L g1846 ( .A(n_1847), .Y(n_1846) );
BUFx3_ASAP7_75t_L g1847 ( .A(n_1848), .Y(n_1847) );
INVxp33_ASAP7_75t_SL g1849 ( .A(n_1850), .Y(n_1849) );
NOR2x1_ASAP7_75t_L g1851 ( .A(n_1852), .B(n_1861), .Y(n_1851) );
NAND2xp5_ASAP7_75t_L g1861 ( .A(n_1862), .B(n_1880), .Y(n_1861) );
OAI31xp33_ASAP7_75t_L g1862 ( .A1(n_1863), .A2(n_1870), .A3(n_1877), .B(n_1879), .Y(n_1862) );
HB1xp67_ASAP7_75t_L g1866 ( .A(n_1867), .Y(n_1866) );
HB1xp67_ASAP7_75t_L g1891 ( .A(n_1892), .Y(n_1891) );
OAI21xp5_ASAP7_75t_L g1892 ( .A1(n_1893), .A2(n_1894), .B(n_1895), .Y(n_1892) );
INVx1_ASAP7_75t_L g1895 ( .A(n_1896), .Y(n_1895) );
endmodule