module fake_netlist_1_9068_n_857 (n_44, n_81, n_69, n_22, n_57, n_88, n_52, n_26, n_50, n_33, n_102, n_73, n_49, n_97, n_80, n_107, n_60, n_41, n_35, n_94, n_65, n_9, n_10, n_103, n_19, n_87, n_104, n_98, n_74, n_7, n_29, n_45, n_85, n_101, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_91, n_108, n_16, n_13, n_95, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_84, n_55, n_12, n_86, n_75, n_105, n_72, n_43, n_76, n_89, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_83, n_28, n_48, n_100, n_92, n_11, n_25, n_30, n_59, n_3, n_18, n_110, n_66, n_1, n_82, n_106, n_15, n_61, n_21, n_99, n_109, n_93, n_51, n_96, n_39, n_857);
input n_44;
input n_81;
input n_69;
input n_22;
input n_57;
input n_88;
input n_52;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_97;
input n_80;
input n_107;
input n_60;
input n_41;
input n_35;
input n_94;
input n_65;
input n_9;
input n_10;
input n_103;
input n_19;
input n_87;
input n_104;
input n_98;
input n_74;
input n_7;
input n_29;
input n_45;
input n_85;
input n_101;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_108;
input n_16;
input n_13;
input n_95;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_84;
input n_55;
input n_12;
input n_86;
input n_75;
input n_105;
input n_72;
input n_43;
input n_76;
input n_89;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_83;
input n_28;
input n_48;
input n_100;
input n_92;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_110;
input n_66;
input n_1;
input n_82;
input n_106;
input n_15;
input n_61;
input n_21;
input n_99;
input n_109;
input n_93;
input n_51;
input n_96;
input n_39;
output n_857;
wire n_117;
wire n_663;
wire n_707;
wire n_791;
wire n_361;
wire n_513;
wire n_838;
wire n_185;
wire n_705;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_755;
wire n_646;
wire n_792;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_848;
wire n_607;
wire n_808;
wire n_829;
wire n_125;
wire n_431;
wire n_484;
wire n_852;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_801;
wire n_292;
wire n_309;
wire n_160;
wire n_701;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_743;
wire n_523;
wire n_229;
wire n_757;
wire n_750;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_770;
wire n_252;
wire n_152;
wire n_113;
wire n_814;
wire n_637;
wire n_817;
wire n_802;
wire n_856;
wire n_353;
wire n_564;
wire n_779;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_850;
wire n_762;
wire n_672;
wire n_532;
wire n_627;
wire n_758;
wire n_544;
wire n_400;
wire n_787;
wire n_853;
wire n_296;
wire n_157;
wire n_765;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_807;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_783;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_715;
wire n_463;
wire n_131;
wire n_112;
wire n_789;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_812;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_777;
wire n_732;
wire n_752;
wire n_199;
wire n_351;
wire n_401;
wire n_461;
wire n_305;
wire n_599;
wire n_228;
wire n_724;
wire n_786;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_796;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_773;
wire n_847;
wire n_840;
wire n_392;
wire n_668;
wire n_846;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_830;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_167;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_726;
wire n_780;
wire n_712;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_809;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_854;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_764;
wire n_314;
wire n_237;
wire n_181;
wire n_255;
wire n_426;
wire n_624;
wire n_725;
wire n_769;
wire n_818;
wire n_844;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_738;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_798;
wire n_241;
wire n_575;
wire n_238;
wire n_711;
wire n_318;
wire n_471;
wire n_632;
wire n_767;
wire n_828;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_490;
wire n_247;
wire n_648;
wire n_613;
wire n_381;
wire n_550;
wire n_826;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_708;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_730;
wire n_735;
wire n_696;
wire n_771;
wire n_784;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_813;
wire n_352;
wire n_746;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_803;
wire n_299;
wire n_338;
wire n_519;
wire n_729;
wire n_699;
wire n_805;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_849;
wire n_810;
wire n_172;
wire n_329;
wire n_251;
wire n_747;
wire n_635;
wire n_731;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_719;
wire n_611;
wire n_704;
wire n_633;
wire n_271;
wire n_760;
wire n_751;
wire n_800;
wire n_626;
wire n_302;
wire n_466;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_412;
wire n_664;
wire n_827;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_788;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_839;
wire n_450;
wire n_579;
wire n_776;
wire n_403;
wire n_557;
wire n_516;
wire n_842;
wire n_254;
wire n_549;
wire n_622;
wire n_832;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_768;
wire n_797;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_666;
wire n_799;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_706;
wire n_823;
wire n_822;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_720;
wire n_568;
wire n_245;
wire n_357;
wire n_653;
wire n_716;
wire n_260;
wire n_806;
wire n_539;
wire n_201;
wire n_197;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_718;
wire n_111;
wire n_536;
wire n_816;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_754;
wire n_775;
wire n_616;
wire n_118;
wire n_365;
wire n_717;
wire n_541;
wire n_179;
wire n_363;
wire n_409;
wire n_315;
wire n_733;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_428;
wire n_364;
wire n_566;
wire n_794;
wire n_376;
wire n_639;
wire n_552;
wire n_744;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_756;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_790;
wire n_761;
wire n_615;
wire n_212;
wire n_472;
wire n_419;
wire n_851;
wire n_825;
wire n_396;
wire n_168;
wire n_804;
wire n_477;
wire n_815;
wire n_570;
wire n_508;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_721;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_821;
wire n_745;
wire n_684;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_723;
wire n_811;
wire n_749;
wire n_835;
wire n_225;
wire n_535;
wire n_530;
wire n_737;
wire n_778;
wire n_220;
wire n_358;
wire n_795;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_782;
wire n_449;
wire n_115;
wire n_300;
wire n_158;
wire n_734;
wire n_524;
wire n_121;
wire n_584;
wire n_763;
wire n_497;
wire n_728;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_841;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_180;
wire n_441;
wire n_836;
wire n_561;
wire n_335;
wire n_272;
wire n_741;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_766;
wire n_602;
wire n_831;
wire n_198;
wire n_169;
wire n_424;
wire n_714;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_837;
wire n_128;
wire n_129;
wire n_410;
wire n_774;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_855;
wire n_722;
wire n_618;
wire n_834;
wire n_727;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_785;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_748;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_820;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_843;
wire n_266;
wire n_683;
wire n_213;
wire n_824;
wire n_538;
wire n_793;
wire n_182;
wire n_492;
wire n_592;
wire n_753;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_695;
wire n_469;
wire n_742;
wire n_585;
wire n_845;
wire n_713;
wire n_123;
wire n_457;
wire n_595;
wire n_759;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_833;
wire n_736;
wire n_194;
wire n_287;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_781;
wire n_421;
wire n_175;
wire n_709;
wire n_739;
wire n_145;
wire n_740;
wire n_483;
wire n_408;
wire n_772;
wire n_290;
wire n_405;
wire n_819;
wire n_280;
wire n_132;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
CKINVDCx5p33_ASAP7_75t_R g111 ( .A(n_95), .Y(n_111) );
CKINVDCx16_ASAP7_75t_R g112 ( .A(n_57), .Y(n_112) );
CKINVDCx5p33_ASAP7_75t_R g113 ( .A(n_61), .Y(n_113) );
CKINVDCx5p33_ASAP7_75t_R g114 ( .A(n_45), .Y(n_114) );
CKINVDCx5p33_ASAP7_75t_R g115 ( .A(n_14), .Y(n_115) );
BUFx8_ASAP7_75t_SL g116 ( .A(n_105), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_69), .Y(n_117) );
CKINVDCx5p33_ASAP7_75t_R g118 ( .A(n_71), .Y(n_118) );
CKINVDCx5p33_ASAP7_75t_R g119 ( .A(n_26), .Y(n_119) );
INVx1_ASAP7_75t_SL g120 ( .A(n_26), .Y(n_120) );
CKINVDCx5p33_ASAP7_75t_R g121 ( .A(n_3), .Y(n_121) );
CKINVDCx5p33_ASAP7_75t_R g122 ( .A(n_63), .Y(n_122) );
CKINVDCx5p33_ASAP7_75t_R g123 ( .A(n_2), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_38), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_87), .Y(n_125) );
INVx1_ASAP7_75t_SL g126 ( .A(n_72), .Y(n_126) );
INVx1_ASAP7_75t_SL g127 ( .A(n_30), .Y(n_127) );
CKINVDCx5p33_ASAP7_75t_R g128 ( .A(n_33), .Y(n_128) );
CKINVDCx5p33_ASAP7_75t_R g129 ( .A(n_76), .Y(n_129) );
CKINVDCx5p33_ASAP7_75t_R g130 ( .A(n_59), .Y(n_130) );
CKINVDCx5p33_ASAP7_75t_R g131 ( .A(n_103), .Y(n_131) );
INVx1_ASAP7_75t_L g132 ( .A(n_101), .Y(n_132) );
CKINVDCx5p33_ASAP7_75t_R g133 ( .A(n_35), .Y(n_133) );
INVx1_ASAP7_75t_L g134 ( .A(n_104), .Y(n_134) );
INVx1_ASAP7_75t_L g135 ( .A(n_99), .Y(n_135) );
CKINVDCx14_ASAP7_75t_R g136 ( .A(n_93), .Y(n_136) );
CKINVDCx5p33_ASAP7_75t_R g137 ( .A(n_65), .Y(n_137) );
INVx1_ASAP7_75t_L g138 ( .A(n_15), .Y(n_138) );
INVx1_ASAP7_75t_L g139 ( .A(n_81), .Y(n_139) );
CKINVDCx20_ASAP7_75t_R g140 ( .A(n_9), .Y(n_140) );
CKINVDCx5p33_ASAP7_75t_R g141 ( .A(n_92), .Y(n_141) );
INVx2_ASAP7_75t_L g142 ( .A(n_84), .Y(n_142) );
BUFx6f_ASAP7_75t_L g143 ( .A(n_32), .Y(n_143) );
CKINVDCx14_ASAP7_75t_R g144 ( .A(n_98), .Y(n_144) );
CKINVDCx5p33_ASAP7_75t_R g145 ( .A(n_97), .Y(n_145) );
INVx1_ASAP7_75t_L g146 ( .A(n_66), .Y(n_146) );
INVx1_ASAP7_75t_L g147 ( .A(n_23), .Y(n_147) );
INVx2_ASAP7_75t_L g148 ( .A(n_21), .Y(n_148) );
BUFx3_ASAP7_75t_L g149 ( .A(n_24), .Y(n_149) );
INVx1_ASAP7_75t_L g150 ( .A(n_51), .Y(n_150) );
INVx1_ASAP7_75t_L g151 ( .A(n_96), .Y(n_151) );
INVx2_ASAP7_75t_L g152 ( .A(n_142), .Y(n_152) );
INVx1_ASAP7_75t_L g153 ( .A(n_117), .Y(n_153) );
INVx5_ASAP7_75t_L g154 ( .A(n_142), .Y(n_154) );
INVx5_ASAP7_75t_L g155 ( .A(n_142), .Y(n_155) );
NAND2xp5_ASAP7_75t_L g156 ( .A(n_124), .B(n_0), .Y(n_156) );
AND2x2_ASAP7_75t_L g157 ( .A(n_112), .B(n_0), .Y(n_157) );
HB1xp67_ASAP7_75t_L g158 ( .A(n_149), .Y(n_158) );
AND2x2_ASAP7_75t_L g159 ( .A(n_112), .B(n_1), .Y(n_159) );
AND2x4_ASAP7_75t_L g160 ( .A(n_149), .B(n_1), .Y(n_160) );
INVx1_ASAP7_75t_L g161 ( .A(n_117), .Y(n_161) );
HB1xp67_ASAP7_75t_L g162 ( .A(n_149), .Y(n_162) );
BUFx6f_ASAP7_75t_L g163 ( .A(n_143), .Y(n_163) );
INVx2_ASAP7_75t_L g164 ( .A(n_143), .Y(n_164) );
BUFx8_ASAP7_75t_L g165 ( .A(n_125), .Y(n_165) );
BUFx6f_ASAP7_75t_L g166 ( .A(n_143), .Y(n_166) );
NOR2xp33_ASAP7_75t_L g167 ( .A(n_125), .B(n_132), .Y(n_167) );
INVx5_ASAP7_75t_L g168 ( .A(n_143), .Y(n_168) );
INVx2_ASAP7_75t_SL g169 ( .A(n_132), .Y(n_169) );
INVx2_ASAP7_75t_SL g170 ( .A(n_134), .Y(n_170) );
NOR2xp33_ASAP7_75t_L g171 ( .A(n_134), .B(n_2), .Y(n_171) );
INVx5_ASAP7_75t_L g172 ( .A(n_143), .Y(n_172) );
CKINVDCx6p67_ASAP7_75t_R g173 ( .A(n_126), .Y(n_173) );
AND2x4_ASAP7_75t_L g174 ( .A(n_148), .B(n_3), .Y(n_174) );
OAI22xp33_ASAP7_75t_SL g175 ( .A1(n_156), .A2(n_119), .B1(n_120), .B2(n_127), .Y(n_175) );
INVx3_ASAP7_75t_L g176 ( .A(n_174), .Y(n_176) );
NAND2xp33_ASAP7_75t_SL g177 ( .A(n_157), .B(n_119), .Y(n_177) );
INVx2_ASAP7_75t_L g178 ( .A(n_152), .Y(n_178) );
AOI22xp5_ASAP7_75t_L g179 ( .A1(n_157), .A2(n_121), .B1(n_123), .B2(n_128), .Y(n_179) );
AOI22xp5_ASAP7_75t_L g180 ( .A1(n_157), .A2(n_114), .B1(n_115), .B2(n_133), .Y(n_180) );
INVx2_ASAP7_75t_L g181 ( .A(n_152), .Y(n_181) );
NAND2xp5_ASAP7_75t_L g182 ( .A(n_158), .B(n_118), .Y(n_182) );
INVx2_ASAP7_75t_L g183 ( .A(n_152), .Y(n_183) );
OAI22xp33_ASAP7_75t_L g184 ( .A1(n_156), .A2(n_140), .B1(n_147), .B2(n_138), .Y(n_184) );
OAI22xp33_ASAP7_75t_L g185 ( .A1(n_156), .A2(n_140), .B1(n_147), .B2(n_138), .Y(n_185) );
AND2x2_ASAP7_75t_L g186 ( .A(n_158), .B(n_136), .Y(n_186) );
OAI22xp33_ASAP7_75t_L g187 ( .A1(n_157), .A2(n_124), .B1(n_127), .B2(n_120), .Y(n_187) );
AOI22xp5_ASAP7_75t_L g188 ( .A1(n_159), .A2(n_136), .B1(n_144), .B2(n_148), .Y(n_188) );
OAI22xp33_ASAP7_75t_L g189 ( .A1(n_159), .A2(n_162), .B1(n_158), .B2(n_148), .Y(n_189) );
INVx1_ASAP7_75t_L g190 ( .A(n_162), .Y(n_190) );
AND2x2_ASAP7_75t_L g191 ( .A(n_162), .B(n_144), .Y(n_191) );
OR2x2_ASAP7_75t_L g192 ( .A(n_159), .B(n_143), .Y(n_192) );
AOI22xp5_ASAP7_75t_L g193 ( .A1(n_159), .A2(n_118), .B1(n_145), .B2(n_143), .Y(n_193) );
OAI22xp5_ASAP7_75t_L g194 ( .A1(n_173), .A2(n_145), .B1(n_126), .B2(n_151), .Y(n_194) );
AND2x4_ASAP7_75t_L g195 ( .A(n_159), .B(n_135), .Y(n_195) );
OAI22xp33_ASAP7_75t_L g196 ( .A1(n_153), .A2(n_151), .B1(n_150), .B2(n_146), .Y(n_196) );
AND2x2_ASAP7_75t_L g197 ( .A(n_173), .B(n_111), .Y(n_197) );
AOI22xp5_ASAP7_75t_L g198 ( .A1(n_173), .A2(n_150), .B1(n_146), .B2(n_135), .Y(n_198) );
NOR2xp33_ASAP7_75t_L g199 ( .A(n_167), .B(n_139), .Y(n_199) );
OA22x2_ASAP7_75t_L g200 ( .A1(n_174), .A2(n_139), .B1(n_141), .B2(n_137), .Y(n_200) );
CKINVDCx20_ASAP7_75t_R g201 ( .A(n_173), .Y(n_201) );
INVx5_ASAP7_75t_L g202 ( .A(n_160), .Y(n_202) );
AOI22xp5_ASAP7_75t_L g203 ( .A1(n_173), .A2(n_131), .B1(n_130), .B2(n_129), .Y(n_203) );
INVx2_ASAP7_75t_L g204 ( .A(n_152), .Y(n_204) );
OAI22xp33_ASAP7_75t_L g205 ( .A1(n_153), .A2(n_122), .B1(n_113), .B2(n_116), .Y(n_205) );
AND2x2_ASAP7_75t_L g206 ( .A(n_160), .B(n_4), .Y(n_206) );
AND2x2_ASAP7_75t_L g207 ( .A(n_160), .B(n_4), .Y(n_207) );
AO22x2_ASAP7_75t_L g208 ( .A1(n_160), .A2(n_116), .B1(n_6), .B2(n_7), .Y(n_208) );
OR2x6_ASAP7_75t_L g209 ( .A(n_174), .B(n_5), .Y(n_209) );
OA22x2_ASAP7_75t_L g210 ( .A1(n_174), .A2(n_5), .B1(n_6), .B2(n_7), .Y(n_210) );
OAI22xp33_ASAP7_75t_L g211 ( .A1(n_153), .A2(n_8), .B1(n_9), .B2(n_10), .Y(n_211) );
BUFx10_ASAP7_75t_L g212 ( .A(n_160), .Y(n_212) );
OA22x2_ASAP7_75t_L g213 ( .A1(n_174), .A2(n_8), .B1(n_10), .B2(n_11), .Y(n_213) );
AOI22xp5_ASAP7_75t_L g214 ( .A1(n_160), .A2(n_12), .B1(n_13), .B2(n_14), .Y(n_214) );
OAI22xp33_ASAP7_75t_L g215 ( .A1(n_153), .A2(n_12), .B1(n_13), .B2(n_15), .Y(n_215) );
OAI22xp33_ASAP7_75t_SL g216 ( .A1(n_174), .A2(n_16), .B1(n_17), .B2(n_18), .Y(n_216) );
AOI22xp5_ASAP7_75t_L g217 ( .A1(n_160), .A2(n_16), .B1(n_17), .B2(n_18), .Y(n_217) );
OAI22xp33_ASAP7_75t_L g218 ( .A1(n_161), .A2(n_19), .B1(n_20), .B2(n_21), .Y(n_218) );
AND2x2_ASAP7_75t_L g219 ( .A(n_160), .B(n_19), .Y(n_219) );
OAI22xp5_ASAP7_75t_SL g220 ( .A1(n_171), .A2(n_20), .B1(n_22), .B2(n_23), .Y(n_220) );
CKINVDCx5p33_ASAP7_75t_R g221 ( .A(n_201), .Y(n_221) );
NAND2xp5_ASAP7_75t_L g222 ( .A(n_186), .B(n_165), .Y(n_222) );
INVx1_ASAP7_75t_L g223 ( .A(n_176), .Y(n_223) );
INVx2_ASAP7_75t_L g224 ( .A(n_178), .Y(n_224) );
INVx1_ASAP7_75t_L g225 ( .A(n_176), .Y(n_225) );
AND2x2_ASAP7_75t_L g226 ( .A(n_195), .B(n_174), .Y(n_226) );
INVx1_ASAP7_75t_L g227 ( .A(n_181), .Y(n_227) );
INVx1_ASAP7_75t_L g228 ( .A(n_183), .Y(n_228) );
NOR2xp67_ASAP7_75t_L g229 ( .A(n_202), .B(n_169), .Y(n_229) );
NOR2xp33_ASAP7_75t_L g230 ( .A(n_190), .B(n_167), .Y(n_230) );
AND2x2_ASAP7_75t_L g231 ( .A(n_195), .B(n_174), .Y(n_231) );
INVx1_ASAP7_75t_L g232 ( .A(n_204), .Y(n_232) );
NOR2xp33_ASAP7_75t_L g233 ( .A(n_182), .B(n_167), .Y(n_233) );
INVx1_ASAP7_75t_L g234 ( .A(n_212), .Y(n_234) );
INVx1_ASAP7_75t_L g235 ( .A(n_212), .Y(n_235) );
INVx1_ASAP7_75t_L g236 ( .A(n_206), .Y(n_236) );
AND2x2_ASAP7_75t_L g237 ( .A(n_191), .B(n_161), .Y(n_237) );
INVx1_ASAP7_75t_L g238 ( .A(n_207), .Y(n_238) );
NOR2xp33_ASAP7_75t_L g239 ( .A(n_179), .B(n_165), .Y(n_239) );
INVx2_ASAP7_75t_L g240 ( .A(n_202), .Y(n_240) );
AND2x2_ASAP7_75t_SL g241 ( .A(n_219), .B(n_161), .Y(n_241) );
BUFx3_ASAP7_75t_L g242 ( .A(n_209), .Y(n_242) );
INVx1_ASAP7_75t_L g243 ( .A(n_210), .Y(n_243) );
NAND2xp5_ASAP7_75t_L g244 ( .A(n_199), .B(n_165), .Y(n_244) );
BUFx8_ASAP7_75t_L g245 ( .A(n_197), .Y(n_245) );
OAI21xp5_ASAP7_75t_L g246 ( .A1(n_200), .A2(n_170), .B(n_169), .Y(n_246) );
NOR2xp67_ASAP7_75t_L g247 ( .A(n_202), .B(n_169), .Y(n_247) );
AND2x2_ASAP7_75t_L g248 ( .A(n_209), .B(n_161), .Y(n_248) );
OR2x6_ASAP7_75t_L g249 ( .A(n_209), .B(n_169), .Y(n_249) );
AND2x2_ASAP7_75t_L g250 ( .A(n_192), .B(n_171), .Y(n_250) );
XOR2xp5_ASAP7_75t_L g251 ( .A(n_208), .B(n_22), .Y(n_251) );
INVx2_ASAP7_75t_SL g252 ( .A(n_202), .Y(n_252) );
NAND2xp5_ASAP7_75t_L g253 ( .A(n_189), .B(n_165), .Y(n_253) );
NOR2xp33_ASAP7_75t_L g254 ( .A(n_180), .B(n_165), .Y(n_254) );
INVx2_ASAP7_75t_L g255 ( .A(n_200), .Y(n_255) );
INVx1_ASAP7_75t_L g256 ( .A(n_210), .Y(n_256) );
INVx1_ASAP7_75t_L g257 ( .A(n_213), .Y(n_257) );
INVx1_ASAP7_75t_L g258 ( .A(n_213), .Y(n_258) );
NAND2xp5_ASAP7_75t_L g259 ( .A(n_189), .B(n_165), .Y(n_259) );
BUFx3_ASAP7_75t_L g260 ( .A(n_198), .Y(n_260) );
XNOR2x1_ASAP7_75t_L g261 ( .A(n_208), .B(n_24), .Y(n_261) );
INVx1_ASAP7_75t_L g262 ( .A(n_214), .Y(n_262) );
INVx1_ASAP7_75t_L g263 ( .A(n_217), .Y(n_263) );
INVx1_ASAP7_75t_L g264 ( .A(n_216), .Y(n_264) );
INVx1_ASAP7_75t_L g265 ( .A(n_196), .Y(n_265) );
INVx1_ASAP7_75t_L g266 ( .A(n_196), .Y(n_266) );
INVx1_ASAP7_75t_L g267 ( .A(n_208), .Y(n_267) );
NAND2xp5_ASAP7_75t_L g268 ( .A(n_193), .B(n_165), .Y(n_268) );
AND2x2_ASAP7_75t_L g269 ( .A(n_188), .B(n_171), .Y(n_269) );
AND2x4_ASAP7_75t_L g270 ( .A(n_203), .B(n_169), .Y(n_270) );
AOI21x1_ASAP7_75t_L g271 ( .A1(n_194), .A2(n_152), .B(n_164), .Y(n_271) );
INVx3_ASAP7_75t_L g272 ( .A(n_175), .Y(n_272) );
XOR2xp5_ASAP7_75t_L g273 ( .A(n_205), .B(n_25), .Y(n_273) );
INVx1_ASAP7_75t_L g274 ( .A(n_220), .Y(n_274) );
OR2x2_ASAP7_75t_L g275 ( .A(n_184), .B(n_170), .Y(n_275) );
XOR2xp5_ASAP7_75t_L g276 ( .A(n_205), .B(n_25), .Y(n_276) );
NOR2xp33_ASAP7_75t_L g277 ( .A(n_177), .B(n_170), .Y(n_277) );
INVx1_ASAP7_75t_L g278 ( .A(n_211), .Y(n_278) );
INVx1_ASAP7_75t_L g279 ( .A(n_211), .Y(n_279) );
INVxp33_ASAP7_75t_L g280 ( .A(n_184), .Y(n_280) );
NOR2xp33_ASAP7_75t_SL g281 ( .A(n_185), .B(n_152), .Y(n_281) );
HB1xp67_ASAP7_75t_L g282 ( .A(n_249), .Y(n_282) );
AND2x2_ASAP7_75t_L g283 ( .A(n_249), .B(n_170), .Y(n_283) );
AND2x2_ASAP7_75t_SL g284 ( .A(n_248), .B(n_163), .Y(n_284) );
CKINVDCx12_ASAP7_75t_R g285 ( .A(n_249), .Y(n_285) );
AND2x2_ASAP7_75t_L g286 ( .A(n_249), .B(n_170), .Y(n_286) );
INVx1_ASAP7_75t_L g287 ( .A(n_223), .Y(n_287) );
INVx2_ASAP7_75t_L g288 ( .A(n_224), .Y(n_288) );
INVx2_ASAP7_75t_L g289 ( .A(n_224), .Y(n_289) );
INVx4_ASAP7_75t_L g290 ( .A(n_249), .Y(n_290) );
AND2x2_ASAP7_75t_L g291 ( .A(n_237), .B(n_154), .Y(n_291) );
BUFx5_ASAP7_75t_L g292 ( .A(n_241), .Y(n_292) );
INVxp67_ASAP7_75t_L g293 ( .A(n_242), .Y(n_293) );
NAND2xp5_ASAP7_75t_L g294 ( .A(n_241), .B(n_185), .Y(n_294) );
INVx1_ASAP7_75t_L g295 ( .A(n_223), .Y(n_295) );
AND2x2_ASAP7_75t_L g296 ( .A(n_237), .B(n_154), .Y(n_296) );
BUFx6f_ASAP7_75t_L g297 ( .A(n_224), .Y(n_297) );
INVx1_ASAP7_75t_L g298 ( .A(n_225), .Y(n_298) );
HB1xp67_ASAP7_75t_L g299 ( .A(n_242), .Y(n_299) );
INVx1_ASAP7_75t_SL g300 ( .A(n_242), .Y(n_300) );
INVx3_ASAP7_75t_L g301 ( .A(n_240), .Y(n_301) );
INVx2_ASAP7_75t_L g302 ( .A(n_227), .Y(n_302) );
INVx2_ASAP7_75t_SL g303 ( .A(n_248), .Y(n_303) );
AND2x6_ASAP7_75t_L g304 ( .A(n_267), .B(n_215), .Y(n_304) );
INVx4_ASAP7_75t_L g305 ( .A(n_241), .Y(n_305) );
INVxp67_ASAP7_75t_L g306 ( .A(n_234), .Y(n_306) );
CKINVDCx5p33_ASAP7_75t_R g307 ( .A(n_245), .Y(n_307) );
INVx2_ASAP7_75t_L g308 ( .A(n_227), .Y(n_308) );
INVx2_ASAP7_75t_L g309 ( .A(n_228), .Y(n_309) );
BUFx3_ASAP7_75t_L g310 ( .A(n_245), .Y(n_310) );
BUFx4f_ASAP7_75t_L g311 ( .A(n_234), .Y(n_311) );
NAND2xp5_ASAP7_75t_L g312 ( .A(n_264), .B(n_187), .Y(n_312) );
INVx2_ASAP7_75t_L g313 ( .A(n_228), .Y(n_313) );
NOR2xp33_ASAP7_75t_L g314 ( .A(n_233), .B(n_187), .Y(n_314) );
AND2x2_ASAP7_75t_L g315 ( .A(n_253), .B(n_154), .Y(n_315) );
NAND2xp5_ASAP7_75t_L g316 ( .A(n_264), .B(n_154), .Y(n_316) );
AND2x2_ASAP7_75t_L g317 ( .A(n_253), .B(n_154), .Y(n_317) );
NAND2x1p5_ASAP7_75t_L g318 ( .A(n_267), .B(n_154), .Y(n_318) );
AND2x4_ASAP7_75t_L g319 ( .A(n_226), .B(n_154), .Y(n_319) );
HB1xp67_ASAP7_75t_L g320 ( .A(n_235), .Y(n_320) );
AND2x2_ASAP7_75t_L g321 ( .A(n_259), .B(n_154), .Y(n_321) );
BUFx3_ASAP7_75t_L g322 ( .A(n_245), .Y(n_322) );
NAND2xp5_ASAP7_75t_L g323 ( .A(n_269), .B(n_154), .Y(n_323) );
NAND2xp5_ASAP7_75t_L g324 ( .A(n_269), .B(n_154), .Y(n_324) );
INVx1_ASAP7_75t_L g325 ( .A(n_225), .Y(n_325) );
AND2x2_ASAP7_75t_L g326 ( .A(n_259), .B(n_154), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g327 ( .A(n_262), .B(n_154), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g328 ( .A(n_262), .B(n_154), .Y(n_328) );
OAI21x1_ASAP7_75t_L g329 ( .A1(n_271), .A2(n_164), .B(n_155), .Y(n_329) );
INVx2_ASAP7_75t_L g330 ( .A(n_232), .Y(n_330) );
INVx1_ASAP7_75t_L g331 ( .A(n_232), .Y(n_331) );
HB1xp67_ASAP7_75t_L g332 ( .A(n_235), .Y(n_332) );
INVx2_ASAP7_75t_L g333 ( .A(n_240), .Y(n_333) );
AND2x4_ASAP7_75t_L g334 ( .A(n_290), .B(n_226), .Y(n_334) );
INVx2_ASAP7_75t_L g335 ( .A(n_288), .Y(n_335) );
NAND2xp5_ASAP7_75t_L g336 ( .A(n_314), .B(n_263), .Y(n_336) );
NAND2xp5_ASAP7_75t_L g337 ( .A(n_314), .B(n_263), .Y(n_337) );
NOR2xp33_ASAP7_75t_L g338 ( .A(n_314), .B(n_260), .Y(n_338) );
OR2x6_ASAP7_75t_L g339 ( .A(n_290), .B(n_243), .Y(n_339) );
INVx2_ASAP7_75t_L g340 ( .A(n_288), .Y(n_340) );
INVx3_ASAP7_75t_L g341 ( .A(n_290), .Y(n_341) );
BUFx3_ASAP7_75t_L g342 ( .A(n_310), .Y(n_342) );
NAND2xp5_ASAP7_75t_L g343 ( .A(n_294), .B(n_265), .Y(n_343) );
AND2x4_ASAP7_75t_L g344 ( .A(n_290), .B(n_231), .Y(n_344) );
OR2x2_ASAP7_75t_SL g345 ( .A(n_282), .B(n_261), .Y(n_345) );
NAND2xp5_ASAP7_75t_L g346 ( .A(n_294), .B(n_265), .Y(n_346) );
INVx2_ASAP7_75t_L g347 ( .A(n_288), .Y(n_347) );
OR2x2_ASAP7_75t_L g348 ( .A(n_292), .B(n_261), .Y(n_348) );
OR2x6_ASAP7_75t_L g349 ( .A(n_290), .B(n_243), .Y(n_349) );
AND2x4_ASAP7_75t_L g350 ( .A(n_290), .B(n_231), .Y(n_350) );
INVx8_ASAP7_75t_L g351 ( .A(n_283), .Y(n_351) );
CKINVDCx5p33_ASAP7_75t_R g352 ( .A(n_307), .Y(n_352) );
NOR2xp33_ASAP7_75t_SL g353 ( .A(n_290), .B(n_305), .Y(n_353) );
INVx1_ASAP7_75t_L g354 ( .A(n_302), .Y(n_354) );
AND2x4_ASAP7_75t_L g355 ( .A(n_305), .B(n_236), .Y(n_355) );
INVx1_ASAP7_75t_L g356 ( .A(n_302), .Y(n_356) );
INVx4_ASAP7_75t_L g357 ( .A(n_310), .Y(n_357) );
BUFx2_ASAP7_75t_L g358 ( .A(n_292), .Y(n_358) );
INVx2_ASAP7_75t_L g359 ( .A(n_288), .Y(n_359) );
BUFx2_ASAP7_75t_SL g360 ( .A(n_292), .Y(n_360) );
INVx3_ASAP7_75t_L g361 ( .A(n_302), .Y(n_361) );
AND2x2_ASAP7_75t_SL g362 ( .A(n_305), .B(n_275), .Y(n_362) );
NOR2xp33_ASAP7_75t_L g363 ( .A(n_305), .B(n_260), .Y(n_363) );
NAND2x1p5_ASAP7_75t_L g364 ( .A(n_305), .B(n_256), .Y(n_364) );
NAND2x1p5_ASAP7_75t_L g365 ( .A(n_305), .B(n_256), .Y(n_365) );
INVx2_ASAP7_75t_L g366 ( .A(n_288), .Y(n_366) );
BUFx8_ASAP7_75t_L g367 ( .A(n_342), .Y(n_367) );
AND2x2_ASAP7_75t_L g368 ( .A(n_354), .B(n_292), .Y(n_368) );
NAND2x1p5_ASAP7_75t_L g369 ( .A(n_361), .B(n_305), .Y(n_369) );
NAND2x1p5_ASAP7_75t_L g370 ( .A(n_361), .B(n_310), .Y(n_370) );
BUFx10_ASAP7_75t_L g371 ( .A(n_355), .Y(n_371) );
BUFx3_ASAP7_75t_L g372 ( .A(n_342), .Y(n_372) );
OAI22xp5_ASAP7_75t_L g373 ( .A1(n_345), .A2(n_294), .B1(n_261), .B2(n_251), .Y(n_373) );
NOR2xp33_ASAP7_75t_L g374 ( .A(n_338), .B(n_280), .Y(n_374) );
BUFx2_ASAP7_75t_L g375 ( .A(n_354), .Y(n_375) );
BUFx4_ASAP7_75t_SL g376 ( .A(n_352), .Y(n_376) );
NAND2x1p5_ASAP7_75t_L g377 ( .A(n_361), .B(n_310), .Y(n_377) );
NAND2xp5_ASAP7_75t_L g378 ( .A(n_336), .B(n_266), .Y(n_378) );
CKINVDCx14_ASAP7_75t_R g379 ( .A(n_352), .Y(n_379) );
AOI22xp33_ASAP7_75t_L g380 ( .A1(n_338), .A2(n_304), .B1(n_251), .B2(n_292), .Y(n_380) );
INVx4_ASAP7_75t_L g381 ( .A(n_357), .Y(n_381) );
INVx5_ASAP7_75t_L g382 ( .A(n_357), .Y(n_382) );
OR2x6_ASAP7_75t_L g383 ( .A(n_360), .B(n_310), .Y(n_383) );
INVx2_ASAP7_75t_SL g384 ( .A(n_342), .Y(n_384) );
INVx1_ASAP7_75t_L g385 ( .A(n_354), .Y(n_385) );
BUFx3_ASAP7_75t_L g386 ( .A(n_342), .Y(n_386) );
INVx2_ASAP7_75t_L g387 ( .A(n_366), .Y(n_387) );
AND2x2_ASAP7_75t_L g388 ( .A(n_356), .B(n_292), .Y(n_388) );
AND2x4_ASAP7_75t_L g389 ( .A(n_357), .B(n_322), .Y(n_389) );
BUFx2_ASAP7_75t_L g390 ( .A(n_356), .Y(n_390) );
INVx1_ASAP7_75t_L g391 ( .A(n_356), .Y(n_391) );
BUFx2_ASAP7_75t_SL g392 ( .A(n_357), .Y(n_392) );
BUFx6f_ASAP7_75t_L g393 ( .A(n_361), .Y(n_393) );
BUFx12f_ASAP7_75t_L g394 ( .A(n_357), .Y(n_394) );
CKINVDCx5p33_ASAP7_75t_R g395 ( .A(n_351), .Y(n_395) );
CKINVDCx20_ASAP7_75t_R g396 ( .A(n_379), .Y(n_396) );
INVx1_ASAP7_75t_L g397 ( .A(n_385), .Y(n_397) );
BUFx4f_ASAP7_75t_SL g398 ( .A(n_394), .Y(n_398) );
AND2x2_ASAP7_75t_L g399 ( .A(n_375), .B(n_335), .Y(n_399) );
INVx3_ASAP7_75t_L g400 ( .A(n_394), .Y(n_400) );
AOI22xp33_ASAP7_75t_L g401 ( .A1(n_373), .A2(n_304), .B1(n_348), .B2(n_362), .Y(n_401) );
AOI22xp33_ASAP7_75t_SL g402 ( .A1(n_373), .A2(n_362), .B1(n_292), .B2(n_348), .Y(n_402) );
OAI22xp5_ASAP7_75t_L g403 ( .A1(n_380), .A2(n_345), .B1(n_362), .B2(n_348), .Y(n_403) );
INVx2_ASAP7_75t_L g404 ( .A(n_387), .Y(n_404) );
BUFx12f_ASAP7_75t_L g405 ( .A(n_394), .Y(n_405) );
INVxp67_ASAP7_75t_L g406 ( .A(n_375), .Y(n_406) );
AND2x2_ASAP7_75t_L g407 ( .A(n_375), .B(n_366), .Y(n_407) );
AOI22xp33_ASAP7_75t_L g408 ( .A1(n_380), .A2(n_304), .B1(n_362), .B2(n_363), .Y(n_408) );
NAND2xp5_ASAP7_75t_L g409 ( .A(n_385), .B(n_343), .Y(n_409) );
AOI22xp33_ASAP7_75t_SL g410 ( .A1(n_392), .A2(n_292), .B1(n_360), .B2(n_353), .Y(n_410) );
BUFx8_ASAP7_75t_L g411 ( .A(n_394), .Y(n_411) );
CKINVDCx5p33_ASAP7_75t_R g412 ( .A(n_376), .Y(n_412) );
INVx6_ASAP7_75t_SL g413 ( .A(n_371), .Y(n_413) );
CKINVDCx5p33_ASAP7_75t_R g414 ( .A(n_379), .Y(n_414) );
AOI22xp33_ASAP7_75t_L g415 ( .A1(n_374), .A2(n_304), .B1(n_363), .B2(n_292), .Y(n_415) );
INVx6_ASAP7_75t_L g416 ( .A(n_367), .Y(n_416) );
OAI22xp5_ASAP7_75t_SL g417 ( .A1(n_381), .A2(n_345), .B1(n_273), .B2(n_276), .Y(n_417) );
AOI22xp33_ASAP7_75t_L g418 ( .A1(n_374), .A2(n_304), .B1(n_292), .B2(n_360), .Y(n_418) );
CKINVDCx5p33_ASAP7_75t_R g419 ( .A(n_367), .Y(n_419) );
INVx2_ASAP7_75t_L g420 ( .A(n_387), .Y(n_420) );
INVx1_ASAP7_75t_L g421 ( .A(n_385), .Y(n_421) );
INVx2_ASAP7_75t_L g422 ( .A(n_387), .Y(n_422) );
BUFx6f_ASAP7_75t_L g423 ( .A(n_393), .Y(n_423) );
INVx1_ASAP7_75t_L g424 ( .A(n_391), .Y(n_424) );
AOI22xp33_ASAP7_75t_L g425 ( .A1(n_392), .A2(n_304), .B1(n_292), .B2(n_355), .Y(n_425) );
AOI22xp33_ASAP7_75t_SL g426 ( .A1(n_392), .A2(n_292), .B1(n_353), .B2(n_304), .Y(n_426) );
BUFx3_ASAP7_75t_L g427 ( .A(n_367), .Y(n_427) );
BUFx2_ASAP7_75t_R g428 ( .A(n_395), .Y(n_428) );
INVx3_ASAP7_75t_SL g429 ( .A(n_382), .Y(n_429) );
CKINVDCx20_ASAP7_75t_R g430 ( .A(n_367), .Y(n_430) );
INVx4_ASAP7_75t_L g431 ( .A(n_382), .Y(n_431) );
NAND2xp5_ASAP7_75t_L g432 ( .A(n_391), .B(n_343), .Y(n_432) );
INVx4_ASAP7_75t_L g433 ( .A(n_382), .Y(n_433) );
INVx4_ASAP7_75t_L g434 ( .A(n_382), .Y(n_434) );
AOI22xp33_ASAP7_75t_L g435 ( .A1(n_381), .A2(n_304), .B1(n_292), .B2(n_355), .Y(n_435) );
AOI22xp33_ASAP7_75t_L g436 ( .A1(n_381), .A2(n_304), .B1(n_292), .B2(n_355), .Y(n_436) );
INVx1_ASAP7_75t_L g437 ( .A(n_391), .Y(n_437) );
INVx2_ASAP7_75t_L g438 ( .A(n_387), .Y(n_438) );
OAI22xp5_ASAP7_75t_L g439 ( .A1(n_401), .A2(n_382), .B1(n_381), .B2(n_390), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_397), .Y(n_440) );
AOI22xp33_ASAP7_75t_L g441 ( .A1(n_403), .A2(n_304), .B1(n_381), .B2(n_292), .Y(n_441) );
INVx1_ASAP7_75t_SL g442 ( .A(n_398), .Y(n_442) );
BUFx4f_ASAP7_75t_L g443 ( .A(n_429), .Y(n_443) );
INVx1_ASAP7_75t_L g444 ( .A(n_397), .Y(n_444) );
INVx1_ASAP7_75t_L g445 ( .A(n_421), .Y(n_445) );
INVx2_ASAP7_75t_L g446 ( .A(n_404), .Y(n_446) );
AOI22xp33_ASAP7_75t_L g447 ( .A1(n_403), .A2(n_417), .B1(n_402), .B2(n_401), .Y(n_447) );
OAI22xp5_ASAP7_75t_L g448 ( .A1(n_417), .A2(n_382), .B1(n_381), .B2(n_390), .Y(n_448) );
OAI22xp5_ASAP7_75t_L g449 ( .A1(n_402), .A2(n_382), .B1(n_390), .B2(n_383), .Y(n_449) );
AOI22xp33_ASAP7_75t_L g450 ( .A1(n_408), .A2(n_304), .B1(n_292), .B2(n_322), .Y(n_450) );
OAI22xp5_ASAP7_75t_L g451 ( .A1(n_426), .A2(n_382), .B1(n_383), .B2(n_273), .Y(n_451) );
OAI21xp5_ASAP7_75t_SL g452 ( .A1(n_400), .A2(n_276), .B(n_389), .Y(n_452) );
BUFx2_ASAP7_75t_L g453 ( .A(n_433), .Y(n_453) );
INVx1_ASAP7_75t_L g454 ( .A(n_424), .Y(n_454) );
OAI22xp5_ASAP7_75t_SL g455 ( .A1(n_430), .A2(n_285), .B1(n_307), .B2(n_221), .Y(n_455) );
AOI22xp33_ASAP7_75t_L g456 ( .A1(n_408), .A2(n_304), .B1(n_292), .B2(n_322), .Y(n_456) );
OAI22xp33_ASAP7_75t_L g457 ( .A1(n_398), .A2(n_382), .B1(n_322), .B2(n_383), .Y(n_457) );
INVx1_ASAP7_75t_L g458 ( .A(n_424), .Y(n_458) );
INVx2_ASAP7_75t_L g459 ( .A(n_404), .Y(n_459) );
AOI22xp33_ASAP7_75t_SL g460 ( .A1(n_416), .A2(n_367), .B1(n_322), .B2(n_389), .Y(n_460) );
CKINVDCx5p33_ASAP7_75t_R g461 ( .A(n_412), .Y(n_461) );
HB1xp67_ASAP7_75t_L g462 ( .A(n_399), .Y(n_462) );
AOI22xp33_ASAP7_75t_L g463 ( .A1(n_415), .A2(n_304), .B1(n_292), .B2(n_367), .Y(n_463) );
AOI22xp33_ASAP7_75t_SL g464 ( .A1(n_416), .A2(n_389), .B1(n_371), .B2(n_304), .Y(n_464) );
OAI21xp33_ASAP7_75t_L g465 ( .A1(n_426), .A2(n_281), .B(n_279), .Y(n_465) );
AND2x4_ASAP7_75t_L g466 ( .A(n_427), .B(n_389), .Y(n_466) );
AOI22xp33_ASAP7_75t_SL g467 ( .A1(n_416), .A2(n_389), .B1(n_371), .B2(n_372), .Y(n_467) );
OAI22xp5_ASAP7_75t_L g468 ( .A1(n_425), .A2(n_383), .B1(n_369), .B2(n_389), .Y(n_468) );
AOI22xp33_ASAP7_75t_L g469 ( .A1(n_415), .A2(n_358), .B1(n_371), .B2(n_355), .Y(n_469) );
INVx2_ASAP7_75t_L g470 ( .A(n_404), .Y(n_470) );
OR2x2_ASAP7_75t_L g471 ( .A(n_406), .B(n_369), .Y(n_471) );
AOI22xp33_ASAP7_75t_L g472 ( .A1(n_435), .A2(n_358), .B1(n_371), .B2(n_355), .Y(n_472) );
INVx1_ASAP7_75t_L g473 ( .A(n_437), .Y(n_473) );
NAND2xp5_ASAP7_75t_L g474 ( .A(n_437), .B(n_278), .Y(n_474) );
NAND2xp5_ASAP7_75t_L g475 ( .A(n_399), .B(n_278), .Y(n_475) );
AOI22xp33_ASAP7_75t_SL g476 ( .A1(n_416), .A2(n_371), .B1(n_372), .B2(n_386), .Y(n_476) );
OAI22xp5_ASAP7_75t_L g477 ( .A1(n_435), .A2(n_383), .B1(n_369), .B2(n_370), .Y(n_477) );
AOI22xp33_ASAP7_75t_L g478 ( .A1(n_436), .A2(n_358), .B1(n_383), .B2(n_337), .Y(n_478) );
NOR2xp33_ASAP7_75t_L g479 ( .A(n_414), .B(n_274), .Y(n_479) );
AOI22xp33_ASAP7_75t_L g480 ( .A1(n_436), .A2(n_336), .B1(n_337), .B2(n_350), .Y(n_480) );
NAND3xp33_ASAP7_75t_L g481 ( .A(n_411), .B(n_246), .C(n_281), .Y(n_481) );
OAI21xp5_ASAP7_75t_L g482 ( .A1(n_418), .A2(n_254), .B(n_239), .Y(n_482) );
NAND2xp5_ASAP7_75t_L g483 ( .A(n_399), .B(n_279), .Y(n_483) );
AOI22xp33_ASAP7_75t_L g484 ( .A1(n_418), .A2(n_350), .B1(n_334), .B2(n_344), .Y(n_484) );
INVx1_ASAP7_75t_L g485 ( .A(n_420), .Y(n_485) );
BUFx2_ASAP7_75t_L g486 ( .A(n_433), .Y(n_486) );
AOI22xp33_ASAP7_75t_SL g487 ( .A1(n_416), .A2(n_427), .B1(n_405), .B2(n_411), .Y(n_487) );
AND2x2_ASAP7_75t_L g488 ( .A(n_407), .B(n_368), .Y(n_488) );
OAI22xp5_ASAP7_75t_L g489 ( .A1(n_427), .A2(n_369), .B1(n_377), .B2(n_370), .Y(n_489) );
AOI22xp33_ASAP7_75t_SL g490 ( .A1(n_405), .A2(n_372), .B1(n_386), .B2(n_351), .Y(n_490) );
INVx1_ASAP7_75t_L g491 ( .A(n_420), .Y(n_491) );
OAI22xp5_ASAP7_75t_L g492 ( .A1(n_410), .A2(n_370), .B1(n_377), .B2(n_282), .Y(n_492) );
NAND2xp5_ASAP7_75t_L g493 ( .A(n_407), .B(n_368), .Y(n_493) );
AOI22xp33_ASAP7_75t_L g494 ( .A1(n_411), .A2(n_350), .B1(n_334), .B2(n_344), .Y(n_494) );
AOI22xp33_ASAP7_75t_SL g495 ( .A1(n_411), .A2(n_372), .B1(n_386), .B2(n_351), .Y(n_495) );
OAI22xp5_ASAP7_75t_L g496 ( .A1(n_410), .A2(n_370), .B1(n_377), .B2(n_282), .Y(n_496) );
INVx2_ASAP7_75t_L g497 ( .A(n_420), .Y(n_497) );
AOI22xp33_ASAP7_75t_SL g498 ( .A1(n_411), .A2(n_386), .B1(n_351), .B2(n_384), .Y(n_498) );
AOI22xp33_ASAP7_75t_L g499 ( .A1(n_433), .A2(n_344), .B1(n_334), .B2(n_350), .Y(n_499) );
AOI22xp33_ASAP7_75t_SL g500 ( .A1(n_400), .A2(n_351), .B1(n_384), .B2(n_377), .Y(n_500) );
INVx2_ASAP7_75t_L g501 ( .A(n_422), .Y(n_501) );
OAI22xp5_ASAP7_75t_L g502 ( .A1(n_400), .A2(n_377), .B1(n_341), .B2(n_339), .Y(n_502) );
AOI22xp33_ASAP7_75t_SL g503 ( .A1(n_400), .A2(n_351), .B1(n_384), .B2(n_341), .Y(n_503) );
INVx2_ASAP7_75t_L g504 ( .A(n_422), .Y(n_504) );
AOI22xp33_ASAP7_75t_L g505 ( .A1(n_433), .A2(n_344), .B1(n_334), .B2(n_350), .Y(n_505) );
INVx1_ASAP7_75t_L g506 ( .A(n_422), .Y(n_506) );
INVx1_ASAP7_75t_SL g507 ( .A(n_396), .Y(n_507) );
AOI22xp33_ASAP7_75t_SL g508 ( .A1(n_451), .A2(n_433), .B1(n_434), .B2(n_431), .Y(n_508) );
AOI22xp33_ASAP7_75t_L g509 ( .A1(n_447), .A2(n_434), .B1(n_431), .B2(n_413), .Y(n_509) );
OAI221xp5_ASAP7_75t_L g510 ( .A1(n_452), .A2(n_272), .B1(n_274), .B2(n_312), .C(n_378), .Y(n_510) );
OAI22xp5_ASAP7_75t_L g511 ( .A1(n_441), .A2(n_406), .B1(n_434), .B2(n_431), .Y(n_511) );
AOI22xp5_ASAP7_75t_L g512 ( .A1(n_448), .A2(n_419), .B1(n_215), .B2(n_218), .Y(n_512) );
AOI22xp33_ASAP7_75t_SL g513 ( .A1(n_453), .A2(n_434), .B1(n_431), .B2(n_407), .Y(n_513) );
AOI22xp33_ASAP7_75t_SL g514 ( .A1(n_453), .A2(n_351), .B1(n_432), .B2(n_409), .Y(n_514) );
AOI22xp33_ASAP7_75t_L g515 ( .A1(n_463), .A2(n_413), .B1(n_429), .B2(n_341), .Y(n_515) );
AOI22xp33_ASAP7_75t_L g516 ( .A1(n_450), .A2(n_413), .B1(n_429), .B2(n_341), .Y(n_516) );
AOI22xp33_ASAP7_75t_SL g517 ( .A1(n_486), .A2(n_351), .B1(n_432), .B2(n_409), .Y(n_517) );
AOI22xp33_ASAP7_75t_L g518 ( .A1(n_456), .A2(n_413), .B1(n_341), .B2(n_388), .Y(n_518) );
OAI221xp5_ASAP7_75t_SL g519 ( .A1(n_480), .A2(n_218), .B1(n_312), .B2(n_378), .C(n_272), .Y(n_519) );
AOI22xp33_ASAP7_75t_L g520 ( .A1(n_449), .A2(n_413), .B1(n_341), .B2(n_368), .Y(n_520) );
OAI221xp5_ASAP7_75t_L g521 ( .A1(n_487), .A2(n_272), .B1(n_312), .B2(n_246), .C(n_266), .Y(n_521) );
AOI22xp33_ASAP7_75t_L g522 ( .A1(n_464), .A2(n_468), .B1(n_478), .B2(n_482), .Y(n_522) );
HB1xp67_ASAP7_75t_L g523 ( .A(n_486), .Y(n_523) );
AND2x2_ASAP7_75t_L g524 ( .A(n_462), .B(n_438), .Y(n_524) );
INVx1_ASAP7_75t_L g525 ( .A(n_440), .Y(n_525) );
AOI22xp33_ASAP7_75t_L g526 ( .A1(n_465), .A2(n_388), .B1(n_339), .B2(n_349), .Y(n_526) );
HB1xp67_ASAP7_75t_L g527 ( .A(n_471), .Y(n_527) );
AOI22xp33_ASAP7_75t_L g528 ( .A1(n_465), .A2(n_388), .B1(n_339), .B2(n_349), .Y(n_528) );
INVx1_ASAP7_75t_L g529 ( .A(n_440), .Y(n_529) );
OAI22xp5_ASAP7_75t_L g530 ( .A1(n_443), .A2(n_438), .B1(n_428), .B2(n_361), .Y(n_530) );
AOI22xp33_ASAP7_75t_L g531 ( .A1(n_439), .A2(n_339), .B1(n_349), .B2(n_344), .Y(n_531) );
AOI22xp33_ASAP7_75t_L g532 ( .A1(n_484), .A2(n_339), .B1(n_349), .B2(n_344), .Y(n_532) );
AOI22xp33_ASAP7_75t_SL g533 ( .A1(n_443), .A2(n_245), .B1(n_438), .B2(n_423), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_488), .B(n_255), .Y(n_534) );
OAI22xp5_ASAP7_75t_L g535 ( .A1(n_443), .A2(n_428), .B1(n_349), .B2(n_339), .Y(n_535) );
AOI22xp33_ASAP7_75t_L g536 ( .A1(n_469), .A2(n_339), .B1(n_349), .B2(n_334), .Y(n_536) );
AOI22xp5_ASAP7_75t_L g537 ( .A1(n_460), .A2(n_285), .B1(n_346), .B2(n_334), .Y(n_537) );
AOI22xp33_ASAP7_75t_L g538 ( .A1(n_477), .A2(n_349), .B1(n_350), .B2(n_255), .Y(n_538) );
AOI22xp33_ASAP7_75t_L g539 ( .A1(n_472), .A2(n_255), .B1(n_258), .B2(n_257), .Y(n_539) );
OAI22xp5_ASAP7_75t_L g540 ( .A1(n_499), .A2(n_364), .B1(n_365), .B2(n_366), .Y(n_540) );
AOI22xp33_ASAP7_75t_L g541 ( .A1(n_466), .A2(n_364), .B1(n_365), .B2(n_326), .Y(n_541) );
AOI22xp33_ASAP7_75t_SL g542 ( .A1(n_466), .A2(n_423), .B1(n_393), .B2(n_270), .Y(n_542) );
AOI22xp33_ASAP7_75t_L g543 ( .A1(n_466), .A2(n_364), .B1(n_365), .B2(n_326), .Y(n_543) );
OAI222xp33_ASAP7_75t_L g544 ( .A1(n_467), .A2(n_365), .B1(n_364), .B2(n_275), .C1(n_300), .C2(n_293), .Y(n_544) );
OAI22xp5_ASAP7_75t_L g545 ( .A1(n_505), .A2(n_365), .B1(n_366), .B2(n_347), .Y(n_545) );
AOI22xp33_ASAP7_75t_L g546 ( .A1(n_492), .A2(n_326), .B1(n_321), .B2(n_317), .Y(n_546) );
OAI22xp33_ASAP7_75t_L g547 ( .A1(n_496), .A2(n_300), .B1(n_393), .B2(n_293), .Y(n_547) );
AOI22xp5_ASAP7_75t_L g548 ( .A1(n_495), .A2(n_303), .B1(n_283), .B2(n_286), .Y(n_548) );
AOI22xp5_ASAP7_75t_L g549 ( .A1(n_498), .A2(n_303), .B1(n_283), .B2(n_286), .Y(n_549) );
OAI22xp5_ASAP7_75t_L g550 ( .A1(n_500), .A2(n_340), .B1(n_359), .B2(n_347), .Y(n_550) );
AOI22xp33_ASAP7_75t_L g551 ( .A1(n_481), .A2(n_326), .B1(n_321), .B2(n_317), .Y(n_551) );
OAI222xp33_ASAP7_75t_L g552 ( .A1(n_489), .A2(n_300), .B1(n_293), .B2(n_340), .C1(n_347), .C2(n_359), .Y(n_552) );
AOI22xp5_ASAP7_75t_L g553 ( .A1(n_457), .A2(n_303), .B1(n_283), .B2(n_286), .Y(n_553) );
OAI22xp5_ASAP7_75t_SL g554 ( .A1(n_455), .A2(n_423), .B1(n_284), .B2(n_299), .Y(n_554) );
AOI22xp33_ASAP7_75t_L g555 ( .A1(n_490), .A2(n_317), .B1(n_315), .B2(n_321), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g556 ( .A(n_488), .B(n_335), .Y(n_556) );
AOI22xp5_ASAP7_75t_SL g557 ( .A1(n_442), .A2(n_423), .B1(n_393), .B2(n_299), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g558 ( .A(n_475), .B(n_335), .Y(n_558) );
AOI22xp5_ASAP7_75t_L g559 ( .A1(n_494), .A2(n_303), .B1(n_286), .B2(n_270), .Y(n_559) );
AOI22xp33_ASAP7_75t_SL g560 ( .A1(n_502), .A2(n_423), .B1(n_393), .B2(n_270), .Y(n_560) );
AOI22xp33_ASAP7_75t_L g561 ( .A1(n_471), .A2(n_315), .B1(n_393), .B2(n_303), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g562 ( .A(n_483), .B(n_335), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g563 ( .A(n_444), .B(n_340), .Y(n_563) );
AOI22xp33_ASAP7_75t_L g564 ( .A1(n_476), .A2(n_393), .B1(n_260), .B2(n_299), .Y(n_564) );
OAI22xp5_ASAP7_75t_L g565 ( .A1(n_503), .A2(n_359), .B1(n_347), .B2(n_340), .Y(n_565) );
AND2x2_ASAP7_75t_L g566 ( .A(n_445), .B(n_423), .Y(n_566) );
OAI22xp5_ASAP7_75t_L g567 ( .A1(n_493), .A2(n_359), .B1(n_393), .B2(n_284), .Y(n_567) );
AOI22xp33_ASAP7_75t_SL g568 ( .A1(n_455), .A2(n_423), .B1(n_284), .B2(n_291), .Y(n_568) );
OAI22xp5_ASAP7_75t_L g569 ( .A1(n_445), .A2(n_284), .B1(n_306), .B2(n_302), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g570 ( .A(n_454), .B(n_316), .Y(n_570) );
AOI22xp33_ASAP7_75t_L g571 ( .A1(n_454), .A2(n_284), .B1(n_331), .B2(n_316), .Y(n_571) );
AOI22xp33_ASAP7_75t_L g572 ( .A1(n_458), .A2(n_284), .B1(n_331), .B2(n_316), .Y(n_572) );
OAI22xp5_ASAP7_75t_L g573 ( .A1(n_507), .A2(n_306), .B1(n_320), .B2(n_332), .Y(n_573) );
AOI22xp33_ASAP7_75t_L g574 ( .A1(n_458), .A2(n_331), .B1(n_328), .B2(n_327), .Y(n_574) );
NOR2xp33_ASAP7_75t_L g575 ( .A(n_479), .B(n_461), .Y(n_575) );
AOI22xp33_ASAP7_75t_L g576 ( .A1(n_473), .A2(n_327), .B1(n_328), .B2(n_324), .Y(n_576) );
AOI222xp33_ASAP7_75t_L g577 ( .A1(n_474), .A2(n_327), .B1(n_328), .B2(n_323), .C1(n_324), .C2(n_250), .Y(n_577) );
AOI22xp33_ASAP7_75t_L g578 ( .A1(n_473), .A2(n_323), .B1(n_324), .B2(n_318), .Y(n_578) );
AOI22xp33_ASAP7_75t_L g579 ( .A1(n_485), .A2(n_323), .B1(n_318), .B2(n_330), .Y(n_579) );
AOI22xp33_ASAP7_75t_L g580 ( .A1(n_485), .A2(n_318), .B1(n_330), .B2(n_302), .Y(n_580) );
AOI22xp33_ASAP7_75t_L g581 ( .A1(n_491), .A2(n_506), .B1(n_504), .B2(n_501), .Y(n_581) );
NAND2xp33_ASAP7_75t_SL g582 ( .A(n_491), .B(n_320), .Y(n_582) );
AOI22xp33_ASAP7_75t_L g583 ( .A1(n_506), .A2(n_318), .B1(n_330), .B2(n_308), .Y(n_583) );
AOI22xp33_ASAP7_75t_L g584 ( .A1(n_446), .A2(n_318), .B1(n_330), .B2(n_308), .Y(n_584) );
CKINVDCx11_ASAP7_75t_R g585 ( .A(n_446), .Y(n_585) );
AOI22xp33_ASAP7_75t_L g586 ( .A1(n_459), .A2(n_318), .B1(n_330), .B2(n_308), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g587 ( .A(n_459), .B(n_308), .Y(n_587) );
AND2x2_ASAP7_75t_L g588 ( .A(n_470), .B(n_164), .Y(n_588) );
AOI22xp33_ASAP7_75t_L g589 ( .A1(n_470), .A2(n_308), .B1(n_309), .B2(n_313), .Y(n_589) );
AOI22xp33_ASAP7_75t_L g590 ( .A1(n_504), .A2(n_309), .B1(n_313), .B2(n_295), .Y(n_590) );
AOI22xp33_ASAP7_75t_L g591 ( .A1(n_497), .A2(n_309), .B1(n_313), .B2(n_295), .Y(n_591) );
AOI22xp33_ASAP7_75t_L g592 ( .A1(n_497), .A2(n_309), .B1(n_313), .B2(n_295), .Y(n_592) );
AOI22xp33_ASAP7_75t_SL g593 ( .A1(n_501), .A2(n_296), .B1(n_291), .B2(n_311), .Y(n_593) );
OAI22xp33_ASAP7_75t_L g594 ( .A1(n_452), .A2(n_311), .B1(n_332), .B2(n_313), .Y(n_594) );
AOI222xp33_ASAP7_75t_L g595 ( .A1(n_452), .A2(n_250), .B1(n_230), .B2(n_296), .C1(n_291), .C2(n_236), .Y(n_595) );
NAND3xp33_ASAP7_75t_SL g596 ( .A(n_452), .B(n_164), .C(n_222), .Y(n_596) );
AOI22xp33_ASAP7_75t_L g597 ( .A1(n_447), .A2(n_309), .B1(n_295), .B2(n_287), .Y(n_597) );
AOI22xp33_ASAP7_75t_L g598 ( .A1(n_447), .A2(n_287), .B1(n_298), .B2(n_325), .Y(n_598) );
AOI22xp5_ASAP7_75t_L g599 ( .A1(n_452), .A2(n_332), .B1(n_277), .B2(n_291), .Y(n_599) );
AOI22xp33_ASAP7_75t_L g600 ( .A1(n_447), .A2(n_287), .B1(n_325), .B2(n_298), .Y(n_600) );
AOI22xp33_ASAP7_75t_L g601 ( .A1(n_447), .A2(n_325), .B1(n_298), .B2(n_296), .Y(n_601) );
OAI222xp33_ASAP7_75t_L g602 ( .A1(n_448), .A2(n_296), .B1(n_155), .B2(n_271), .C1(n_222), .C2(n_289), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g603 ( .A(n_527), .B(n_27), .Y(n_603) );
AND2x2_ASAP7_75t_L g604 ( .A(n_566), .B(n_164), .Y(n_604) );
AND2x2_ASAP7_75t_L g605 ( .A(n_566), .B(n_163), .Y(n_605) );
AOI21xp5_ASAP7_75t_SL g606 ( .A1(n_535), .A2(n_289), .B(n_319), .Y(n_606) );
AOI22xp33_ASAP7_75t_SL g607 ( .A1(n_554), .A2(n_311), .B1(n_319), .B2(n_155), .Y(n_607) );
AND2x2_ASAP7_75t_L g608 ( .A(n_524), .B(n_163), .Y(n_608) );
AND2x2_ASAP7_75t_L g609 ( .A(n_524), .B(n_163), .Y(n_609) );
AOI221xp5_ASAP7_75t_L g610 ( .A1(n_519), .A2(n_163), .B1(n_166), .B2(n_155), .C(n_319), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g611 ( .A(n_525), .B(n_27), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g612 ( .A(n_525), .B(n_28), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g613 ( .A(n_529), .B(n_28), .Y(n_613) );
OAI221xp5_ASAP7_75t_SL g614 ( .A1(n_599), .A2(n_238), .B1(n_268), .B2(n_244), .C(n_333), .Y(n_614) );
AOI22xp5_ASAP7_75t_L g615 ( .A1(n_596), .A2(n_238), .B1(n_319), .B2(n_311), .Y(n_615) );
NAND2x1_ASAP7_75t_L g616 ( .A(n_530), .B(n_163), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g617 ( .A(n_585), .B(n_29), .Y(n_617) );
AND2x2_ASAP7_75t_L g618 ( .A(n_581), .B(n_163), .Y(n_618) );
NAND3xp33_ASAP7_75t_L g619 ( .A(n_595), .B(n_163), .C(n_166), .Y(n_619) );
NAND2xp5_ASAP7_75t_L g620 ( .A(n_523), .B(n_556), .Y(n_620) );
NAND3xp33_ASAP7_75t_L g621 ( .A(n_595), .B(n_163), .C(n_166), .Y(n_621) );
AND2x2_ASAP7_75t_L g622 ( .A(n_520), .B(n_163), .Y(n_622) );
AND2x2_ASAP7_75t_L g623 ( .A(n_513), .B(n_163), .Y(n_623) );
NAND2xp5_ASAP7_75t_L g624 ( .A(n_514), .B(n_29), .Y(n_624) );
OAI22xp5_ASAP7_75t_L g625 ( .A1(n_599), .A2(n_311), .B1(n_289), .B2(n_333), .Y(n_625) );
NOR3xp33_ASAP7_75t_L g626 ( .A(n_521), .B(n_301), .C(n_244), .Y(n_626) );
AND2x2_ASAP7_75t_L g627 ( .A(n_557), .B(n_166), .Y(n_627) );
OAI22xp5_ASAP7_75t_L g628 ( .A1(n_537), .A2(n_311), .B1(n_289), .B2(n_333), .Y(n_628) );
OAI221xp5_ASAP7_75t_SL g629 ( .A1(n_512), .A2(n_268), .B1(n_333), .B2(n_289), .C(n_301), .Y(n_629) );
OAI21xp5_ASAP7_75t_SL g630 ( .A1(n_533), .A2(n_319), .B(n_166), .Y(n_630) );
NAND2xp5_ASAP7_75t_L g631 ( .A(n_517), .B(n_30), .Y(n_631) );
NAND2xp5_ASAP7_75t_L g632 ( .A(n_570), .B(n_31), .Y(n_632) );
NAND3xp33_ASAP7_75t_L g633 ( .A(n_568), .B(n_560), .C(n_582), .Y(n_633) );
OAI22xp5_ASAP7_75t_L g634 ( .A1(n_537), .A2(n_333), .B1(n_155), .B2(n_301), .Y(n_634) );
NAND2xp5_ASAP7_75t_L g635 ( .A(n_567), .B(n_31), .Y(n_635) );
NAND2xp5_ASAP7_75t_L g636 ( .A(n_567), .B(n_32), .Y(n_636) );
OAI22xp5_ASAP7_75t_L g637 ( .A1(n_594), .A2(n_155), .B1(n_301), .B2(n_319), .Y(n_637) );
NAND2xp5_ASAP7_75t_SL g638 ( .A(n_557), .B(n_155), .Y(n_638) );
NAND2xp5_ASAP7_75t_L g639 ( .A(n_522), .B(n_33), .Y(n_639) );
NAND2xp5_ASAP7_75t_SL g640 ( .A(n_530), .B(n_155), .Y(n_640) );
OA211x2_ASAP7_75t_L g641 ( .A1(n_509), .A2(n_34), .B(n_36), .C(n_37), .Y(n_641) );
AND2x2_ASAP7_75t_L g642 ( .A(n_588), .B(n_166), .Y(n_642) );
NAND2xp5_ASAP7_75t_SL g643 ( .A(n_554), .B(n_155), .Y(n_643) );
OAI221xp5_ASAP7_75t_SL g644 ( .A1(n_601), .A2(n_301), .B1(n_36), .B2(n_37), .C(n_38), .Y(n_644) );
NAND2xp5_ASAP7_75t_L g645 ( .A(n_534), .B(n_34), .Y(n_645) );
NAND2xp5_ASAP7_75t_L g646 ( .A(n_558), .B(n_39), .Y(n_646) );
NAND2xp5_ASAP7_75t_L g647 ( .A(n_562), .B(n_39), .Y(n_647) );
NAND2xp5_ASAP7_75t_L g648 ( .A(n_508), .B(n_40), .Y(n_648) );
NAND2xp5_ASAP7_75t_L g649 ( .A(n_538), .B(n_40), .Y(n_649) );
NAND2xp5_ASAP7_75t_L g650 ( .A(n_563), .B(n_41), .Y(n_650) );
NAND3xp33_ASAP7_75t_L g651 ( .A(n_542), .B(n_166), .C(n_168), .Y(n_651) );
OAI22xp5_ASAP7_75t_L g652 ( .A1(n_548), .A2(n_155), .B1(n_301), .B2(n_319), .Y(n_652) );
NAND2xp5_ASAP7_75t_L g653 ( .A(n_577), .B(n_41), .Y(n_653) );
OAI221xp5_ASAP7_75t_SL g654 ( .A1(n_598), .A2(n_301), .B1(n_43), .B2(n_44), .C(n_45), .Y(n_654) );
AND2x4_ASAP7_75t_SL g655 ( .A(n_548), .B(n_553), .Y(n_655) );
NAND2xp5_ASAP7_75t_SL g656 ( .A(n_550), .B(n_155), .Y(n_656) );
NAND3xp33_ASAP7_75t_L g657 ( .A(n_600), .B(n_166), .C(n_168), .Y(n_657) );
NAND2xp5_ASAP7_75t_L g658 ( .A(n_577), .B(n_42), .Y(n_658) );
NAND2xp5_ASAP7_75t_L g659 ( .A(n_576), .B(n_43), .Y(n_659) );
AND2x2_ASAP7_75t_L g660 ( .A(n_540), .B(n_172), .Y(n_660) );
OAI21xp33_ASAP7_75t_SL g661 ( .A1(n_531), .A2(n_329), .B(n_46), .Y(n_661) );
AOI221xp5_ASAP7_75t_L g662 ( .A1(n_510), .A2(n_155), .B1(n_319), .B2(n_172), .C(n_168), .Y(n_662) );
NAND2xp5_ASAP7_75t_L g663 ( .A(n_574), .B(n_44), .Y(n_663) );
NAND3xp33_ASAP7_75t_L g664 ( .A(n_550), .B(n_168), .C(n_172), .Y(n_664) );
NAND2xp5_ASAP7_75t_L g665 ( .A(n_569), .B(n_46), .Y(n_665) );
NAND2xp5_ASAP7_75t_L g666 ( .A(n_545), .B(n_47), .Y(n_666) );
BUFx2_ASAP7_75t_L g667 ( .A(n_587), .Y(n_667) );
OAI22xp5_ASAP7_75t_L g668 ( .A1(n_549), .A2(n_155), .B1(n_297), .B2(n_168), .Y(n_668) );
NAND2xp5_ASAP7_75t_L g669 ( .A(n_597), .B(n_47), .Y(n_669) );
OAI22xp5_ASAP7_75t_L g670 ( .A1(n_549), .A2(n_297), .B1(n_168), .B2(n_172), .Y(n_670) );
AOI221xp5_ASAP7_75t_L g671 ( .A1(n_573), .A2(n_172), .B1(n_168), .B2(n_240), .C(n_252), .Y(n_671) );
AND2x2_ASAP7_75t_L g672 ( .A(n_526), .B(n_172), .Y(n_672) );
NAND2xp5_ASAP7_75t_L g673 ( .A(n_528), .B(n_172), .Y(n_673) );
NAND2xp5_ASAP7_75t_L g674 ( .A(n_546), .B(n_172), .Y(n_674) );
NAND2xp5_ASAP7_75t_L g675 ( .A(n_511), .B(n_172), .Y(n_675) );
AND2x2_ASAP7_75t_L g676 ( .A(n_511), .B(n_172), .Y(n_676) );
NAND2xp5_ASAP7_75t_L g677 ( .A(n_551), .B(n_571), .Y(n_677) );
NAND2xp5_ASAP7_75t_L g678 ( .A(n_572), .B(n_168), .Y(n_678) );
AOI22x1_ASAP7_75t_L g679 ( .A1(n_544), .A2(n_297), .B1(n_252), .B2(n_50), .Y(n_679) );
NAND2xp5_ASAP7_75t_SL g680 ( .A(n_547), .B(n_297), .Y(n_680) );
AOI22xp33_ASAP7_75t_L g681 ( .A1(n_532), .A2(n_329), .B1(n_297), .B2(n_168), .Y(n_681) );
AND2x2_ASAP7_75t_L g682 ( .A(n_565), .B(n_168), .Y(n_682) );
NOR2xp33_ASAP7_75t_L g683 ( .A(n_575), .B(n_48), .Y(n_683) );
NAND2xp5_ASAP7_75t_L g684 ( .A(n_589), .B(n_329), .Y(n_684) );
AOI21xp5_ASAP7_75t_SL g685 ( .A1(n_559), .A2(n_297), .B(n_247), .Y(n_685) );
OAI21xp33_ASAP7_75t_L g686 ( .A1(n_593), .A2(n_297), .B(n_252), .Y(n_686) );
AND2x2_ASAP7_75t_L g687 ( .A(n_541), .B(n_49), .Y(n_687) );
AND2x2_ASAP7_75t_L g688 ( .A(n_543), .B(n_52), .Y(n_688) );
NAND3xp33_ASAP7_75t_L g689 ( .A(n_515), .B(n_297), .C(n_229), .Y(n_689) );
AND2x2_ASAP7_75t_L g690 ( .A(n_578), .B(n_53), .Y(n_690) );
NAND2xp5_ASAP7_75t_SL g691 ( .A(n_564), .B(n_297), .Y(n_691) );
OAI21xp5_ASAP7_75t_L g692 ( .A1(n_552), .A2(n_229), .B(n_55), .Y(n_692) );
NOR2xp33_ASAP7_75t_R g693 ( .A(n_536), .B(n_54), .Y(n_693) );
NAND2xp5_ASAP7_75t_L g694 ( .A(n_561), .B(n_56), .Y(n_694) );
NAND3xp33_ASAP7_75t_L g695 ( .A(n_638), .B(n_516), .C(n_518), .Y(n_695) );
NAND3xp33_ASAP7_75t_L g696 ( .A(n_638), .B(n_555), .C(n_579), .Y(n_696) );
NOR2xp33_ASAP7_75t_L g697 ( .A(n_617), .B(n_559), .Y(n_697) );
BUFx2_ASAP7_75t_L g698 ( .A(n_608), .Y(n_698) );
NAND4xp75_ASAP7_75t_L g699 ( .A(n_643), .B(n_602), .C(n_580), .D(n_583), .Y(n_699) );
AND2x2_ASAP7_75t_SL g700 ( .A(n_627), .B(n_586), .Y(n_700) );
NAND3xp33_ASAP7_75t_L g701 ( .A(n_643), .B(n_584), .C(n_591), .Y(n_701) );
NOR3xp33_ASAP7_75t_L g702 ( .A(n_639), .B(n_539), .C(n_592), .Y(n_702) );
AOI22xp33_ASAP7_75t_L g703 ( .A1(n_633), .A2(n_590), .B1(n_60), .B2(n_62), .Y(n_703) );
OR2x2_ASAP7_75t_L g704 ( .A(n_620), .B(n_58), .Y(n_704) );
AOI22xp33_ASAP7_75t_L g705 ( .A1(n_655), .A2(n_64), .B1(n_67), .B2(n_68), .Y(n_705) );
NOR2xp33_ASAP7_75t_L g706 ( .A(n_603), .B(n_70), .Y(n_706) );
AND2x2_ASAP7_75t_L g707 ( .A(n_604), .B(n_73), .Y(n_707) );
XOR2x2_ASAP7_75t_L g708 ( .A(n_619), .B(n_74), .Y(n_708) );
AND2x2_ASAP7_75t_L g709 ( .A(n_604), .B(n_75), .Y(n_709) );
NAND2xp5_ASAP7_75t_L g710 ( .A(n_667), .B(n_77), .Y(n_710) );
AOI22xp5_ASAP7_75t_SL g711 ( .A1(n_627), .A2(n_78), .B1(n_79), .B2(n_80), .Y(n_711) );
NAND3xp33_ASAP7_75t_L g712 ( .A(n_607), .B(n_82), .C(n_83), .Y(n_712) );
NAND2xp5_ASAP7_75t_L g713 ( .A(n_609), .B(n_605), .Y(n_713) );
INVx2_ASAP7_75t_SL g714 ( .A(n_609), .Y(n_714) );
NOR3xp33_ASAP7_75t_L g715 ( .A(n_644), .B(n_654), .C(n_658), .Y(n_715) );
AOI22xp33_ASAP7_75t_L g716 ( .A1(n_655), .A2(n_85), .B1(n_86), .B2(n_88), .Y(n_716) );
OR2x2_ASAP7_75t_L g717 ( .A(n_611), .B(n_89), .Y(n_717) );
NOR3xp33_ASAP7_75t_L g718 ( .A(n_653), .B(n_90), .C(n_91), .Y(n_718) );
OA211x2_ASAP7_75t_L g719 ( .A1(n_640), .A2(n_94), .B(n_100), .C(n_102), .Y(n_719) );
AND2x2_ASAP7_75t_L g720 ( .A(n_642), .B(n_106), .Y(n_720) );
NOR3xp33_ASAP7_75t_L g721 ( .A(n_648), .B(n_107), .C(n_108), .Y(n_721) );
NAND3xp33_ASAP7_75t_L g722 ( .A(n_679), .B(n_689), .C(n_640), .Y(n_722) );
AND2x2_ASAP7_75t_L g723 ( .A(n_642), .B(n_109), .Y(n_723) );
NAND2xp5_ASAP7_75t_L g724 ( .A(n_635), .B(n_110), .Y(n_724) );
NOR3xp33_ASAP7_75t_SL g725 ( .A(n_630), .B(n_621), .C(n_614), .Y(n_725) );
NOR2xp33_ASAP7_75t_L g726 ( .A(n_683), .B(n_624), .Y(n_726) );
NOR2x1_ASAP7_75t_L g727 ( .A(n_606), .B(n_685), .Y(n_727) );
NAND2xp5_ASAP7_75t_L g728 ( .A(n_636), .B(n_612), .Y(n_728) );
NAND2xp5_ASAP7_75t_L g729 ( .A(n_613), .B(n_666), .Y(n_729) );
AOI22xp33_ASAP7_75t_SL g730 ( .A1(n_693), .A2(n_625), .B1(n_628), .B2(n_692), .Y(n_730) );
NAND2xp5_ASAP7_75t_L g731 ( .A(n_665), .B(n_618), .Y(n_731) );
INVx1_ASAP7_75t_L g732 ( .A(n_618), .Y(n_732) );
NAND4xp75_ASAP7_75t_L g733 ( .A(n_641), .B(n_661), .C(n_631), .D(n_676), .Y(n_733) );
NAND3xp33_ASAP7_75t_L g734 ( .A(n_623), .B(n_610), .C(n_626), .Y(n_734) );
NAND3xp33_ASAP7_75t_L g735 ( .A(n_623), .B(n_664), .C(n_647), .Y(n_735) );
AOI22xp5_ASAP7_75t_L g736 ( .A1(n_677), .A2(n_634), .B1(n_637), .B2(n_662), .Y(n_736) );
AOI22xp33_ASAP7_75t_L g737 ( .A1(n_693), .A2(n_660), .B1(n_657), .B2(n_656), .Y(n_737) );
OR2x2_ASAP7_75t_L g738 ( .A(n_680), .B(n_646), .Y(n_738) );
NOR3xp33_ASAP7_75t_L g739 ( .A(n_632), .B(n_659), .C(n_663), .Y(n_739) );
NOR3xp33_ASAP7_75t_L g740 ( .A(n_650), .B(n_645), .C(n_649), .Y(n_740) );
OR2x2_ASAP7_75t_L g741 ( .A(n_680), .B(n_675), .Y(n_741) );
NOR2xp33_ASAP7_75t_L g742 ( .A(n_669), .B(n_673), .Y(n_742) );
AND2x2_ASAP7_75t_L g743 ( .A(n_622), .B(n_672), .Y(n_743) );
NAND3xp33_ASAP7_75t_L g744 ( .A(n_616), .B(n_651), .C(n_671), .Y(n_744) );
NAND3xp33_ASAP7_75t_L g745 ( .A(n_629), .B(n_682), .C(n_672), .Y(n_745) );
NOR3xp33_ASAP7_75t_SL g746 ( .A(n_686), .B(n_652), .C(n_691), .Y(n_746) );
NAND3xp33_ASAP7_75t_L g747 ( .A(n_682), .B(n_691), .C(n_615), .Y(n_747) );
OR2x2_ASAP7_75t_L g748 ( .A(n_684), .B(n_678), .Y(n_748) );
NOR3xp33_ASAP7_75t_L g749 ( .A(n_694), .B(n_668), .C(n_688), .Y(n_749) );
NAND3xp33_ASAP7_75t_L g750 ( .A(n_681), .B(n_690), .C(n_688), .Y(n_750) );
INVx1_ASAP7_75t_L g751 ( .A(n_687), .Y(n_751) );
NOR2xp33_ASAP7_75t_L g752 ( .A(n_674), .B(n_690), .Y(n_752) );
OR2x2_ASAP7_75t_L g753 ( .A(n_687), .B(n_670), .Y(n_753) );
NOR3xp33_ASAP7_75t_L g754 ( .A(n_639), .B(n_644), .C(n_654), .Y(n_754) );
INVxp33_ASAP7_75t_SL g755 ( .A(n_617), .Y(n_755) );
NOR3xp33_ASAP7_75t_L g756 ( .A(n_639), .B(n_644), .C(n_654), .Y(n_756) );
OR2x2_ASAP7_75t_L g757 ( .A(n_620), .B(n_527), .Y(n_757) );
AOI22xp33_ASAP7_75t_SL g758 ( .A1(n_627), .A2(n_655), .B1(n_633), .B2(n_417), .Y(n_758) );
INVx3_ASAP7_75t_L g759 ( .A(n_627), .Y(n_759) );
NAND2xp5_ASAP7_75t_L g760 ( .A(n_620), .B(n_604), .Y(n_760) );
AOI22xp33_ASAP7_75t_SL g761 ( .A1(n_627), .A2(n_655), .B1(n_633), .B2(n_417), .Y(n_761) );
NAND3xp33_ASAP7_75t_L g762 ( .A(n_638), .B(n_643), .C(n_627), .Y(n_762) );
NAND3xp33_ASAP7_75t_L g763 ( .A(n_638), .B(n_643), .C(n_627), .Y(n_763) );
NAND4xp75_ASAP7_75t_L g764 ( .A(n_727), .B(n_700), .C(n_725), .D(n_726), .Y(n_764) );
OR2x2_ASAP7_75t_L g765 ( .A(n_757), .B(n_760), .Y(n_765) );
XOR2x2_ASAP7_75t_L g766 ( .A(n_755), .B(n_762), .Y(n_766) );
XOR2x2_ASAP7_75t_L g767 ( .A(n_763), .B(n_708), .Y(n_767) );
XNOR2x2_ASAP7_75t_L g768 ( .A(n_722), .B(n_733), .Y(n_768) );
XOR2x2_ASAP7_75t_L g769 ( .A(n_711), .B(n_697), .Y(n_769) );
AOI22xp5_ASAP7_75t_L g770 ( .A1(n_758), .A2(n_761), .B1(n_715), .B2(n_754), .Y(n_770) );
XOR2xp5_ASAP7_75t_L g771 ( .A(n_758), .B(n_761), .Y(n_771) );
NOR3xp33_ASAP7_75t_SL g772 ( .A(n_734), .B(n_695), .C(n_744), .Y(n_772) );
INVx1_ASAP7_75t_L g773 ( .A(n_713), .Y(n_773) );
HB1xp67_ASAP7_75t_L g774 ( .A(n_714), .Y(n_774) );
NAND2xp5_ASAP7_75t_L g775 ( .A(n_732), .B(n_728), .Y(n_775) );
NAND4xp75_ASAP7_75t_SL g776 ( .A(n_742), .B(n_730), .C(n_706), .D(n_752), .Y(n_776) );
NAND4xp75_ASAP7_75t_L g777 ( .A(n_725), .B(n_746), .C(n_729), .D(n_719), .Y(n_777) );
INVx2_ASAP7_75t_L g778 ( .A(n_759), .Y(n_778) );
INVx4_ASAP7_75t_L g779 ( .A(n_759), .Y(n_779) );
INVx2_ASAP7_75t_L g780 ( .A(n_741), .Y(n_780) );
NAND2xp5_ASAP7_75t_L g781 ( .A(n_751), .B(n_731), .Y(n_781) );
NOR4xp25_ASAP7_75t_L g782 ( .A(n_735), .B(n_696), .C(n_738), .D(n_745), .Y(n_782) );
NAND4xp75_ASAP7_75t_L g783 ( .A(n_746), .B(n_736), .C(n_710), .D(n_720), .Y(n_783) );
AND2x4_ASAP7_75t_L g784 ( .A(n_748), .B(n_743), .Y(n_784) );
NAND2xp5_ASAP7_75t_L g785 ( .A(n_739), .B(n_740), .Y(n_785) );
XOR2x2_ASAP7_75t_L g786 ( .A(n_715), .B(n_699), .Y(n_786) );
XOR2x2_ASAP7_75t_L g787 ( .A(n_754), .B(n_756), .Y(n_787) );
INVx5_ASAP7_75t_L g788 ( .A(n_723), .Y(n_788) );
XNOR2xp5_ASAP7_75t_L g789 ( .A(n_730), .B(n_750), .Y(n_789) );
XOR2x2_ASAP7_75t_L g790 ( .A(n_756), .B(n_718), .Y(n_790) );
XOR2x2_ASAP7_75t_L g791 ( .A(n_718), .B(n_739), .Y(n_791) );
NAND4xp75_ASAP7_75t_L g792 ( .A(n_707), .B(n_709), .C(n_724), .D(n_737), .Y(n_792) );
INVx2_ASAP7_75t_L g793 ( .A(n_704), .Y(n_793) );
NAND4xp75_ASAP7_75t_L g794 ( .A(n_749), .B(n_747), .C(n_716), .D(n_705), .Y(n_794) );
NAND2xp5_ASAP7_75t_L g795 ( .A(n_753), .B(n_749), .Y(n_795) );
INVxp33_ASAP7_75t_SL g796 ( .A(n_701), .Y(n_796) );
XOR2x2_ASAP7_75t_L g797 ( .A(n_721), .B(n_712), .Y(n_797) );
AND2x6_ASAP7_75t_L g798 ( .A(n_703), .B(n_702), .Y(n_798) );
INVx2_ASAP7_75t_L g799 ( .A(n_717), .Y(n_799) );
INVx1_ASAP7_75t_L g800 ( .A(n_702), .Y(n_800) );
NAND4xp75_ASAP7_75t_L g801 ( .A(n_727), .B(n_700), .C(n_638), .D(n_643), .Y(n_801) );
INVx2_ASAP7_75t_L g802 ( .A(n_698), .Y(n_802) );
AO22x2_ASAP7_75t_L g803 ( .A1(n_771), .A2(n_800), .B1(n_764), .B2(n_776), .Y(n_803) );
INVx2_ASAP7_75t_L g804 ( .A(n_780), .Y(n_804) );
INVxp33_ASAP7_75t_L g805 ( .A(n_766), .Y(n_805) );
INVxp67_ASAP7_75t_L g806 ( .A(n_768), .Y(n_806) );
INVxp67_ASAP7_75t_L g807 ( .A(n_768), .Y(n_807) );
NOR2xp33_ASAP7_75t_L g808 ( .A(n_796), .B(n_770), .Y(n_808) );
XNOR2xp5_ASAP7_75t_L g809 ( .A(n_786), .B(n_787), .Y(n_809) );
XOR2x2_ASAP7_75t_L g810 ( .A(n_786), .B(n_787), .Y(n_810) );
OAI22xp5_ASAP7_75t_SL g811 ( .A1(n_789), .A2(n_782), .B1(n_785), .B2(n_788), .Y(n_811) );
XNOR2x1_ASAP7_75t_L g812 ( .A(n_790), .B(n_769), .Y(n_812) );
AO22x2_ASAP7_75t_L g813 ( .A1(n_783), .A2(n_801), .B1(n_795), .B2(n_794), .Y(n_813) );
NAND2xp5_ASAP7_75t_L g814 ( .A(n_784), .B(n_773), .Y(n_814) );
XNOR2xp5_ASAP7_75t_L g815 ( .A(n_769), .B(n_790), .Y(n_815) );
INVxp33_ASAP7_75t_L g816 ( .A(n_777), .Y(n_816) );
XNOR2x1_ASAP7_75t_SL g817 ( .A(n_791), .B(n_772), .Y(n_817) );
OAI22x1_ASAP7_75t_L g818 ( .A1(n_815), .A2(n_779), .B1(n_788), .B2(n_772), .Y(n_818) );
XOR2xp5_ASAP7_75t_L g819 ( .A(n_809), .B(n_791), .Y(n_819) );
AO22x2_ASAP7_75t_L g820 ( .A1(n_812), .A2(n_792), .B1(n_775), .B2(n_765), .Y(n_820) );
INVxp67_ASAP7_75t_L g821 ( .A(n_808), .Y(n_821) );
INVx1_ASAP7_75t_L g822 ( .A(n_814), .Y(n_822) );
NAND2xp5_ASAP7_75t_L g823 ( .A(n_806), .B(n_781), .Y(n_823) );
AOI22x1_ASAP7_75t_L g824 ( .A1(n_817), .A2(n_774), .B1(n_802), .B2(n_767), .Y(n_824) );
AOI22xp5_ASAP7_75t_L g825 ( .A1(n_813), .A2(n_798), .B1(n_767), .B2(n_797), .Y(n_825) );
INVx2_ASAP7_75t_L g826 ( .A(n_804), .Y(n_826) );
OA22x2_ASAP7_75t_L g827 ( .A1(n_815), .A2(n_778), .B1(n_799), .B2(n_793), .Y(n_827) );
BUFx2_ASAP7_75t_L g828 ( .A(n_818), .Y(n_828) );
INVx1_ASAP7_75t_SL g829 ( .A(n_823), .Y(n_829) );
INVx2_ASAP7_75t_L g830 ( .A(n_826), .Y(n_830) );
NAND2xp5_ASAP7_75t_L g831 ( .A(n_821), .B(n_807), .Y(n_831) );
INVx1_ASAP7_75t_SL g832 ( .A(n_823), .Y(n_832) );
INVx1_ASAP7_75t_L g833 ( .A(n_822), .Y(n_833) );
INVx1_ASAP7_75t_L g834 ( .A(n_831), .Y(n_834) );
INVx1_ASAP7_75t_L g835 ( .A(n_833), .Y(n_835) );
AOI22xp5_ASAP7_75t_L g836 ( .A1(n_829), .A2(n_825), .B1(n_812), .B2(n_813), .Y(n_836) );
AOI22xp5_ASAP7_75t_L g837 ( .A1(n_832), .A2(n_813), .B1(n_803), .B2(n_820), .Y(n_837) );
INVx2_ASAP7_75t_L g838 ( .A(n_830), .Y(n_838) );
OAI22xp5_ASAP7_75t_L g839 ( .A1(n_837), .A2(n_820), .B1(n_805), .B2(n_824), .Y(n_839) );
NAND2xp5_ASAP7_75t_L g840 ( .A(n_836), .B(n_809), .Y(n_840) );
AOI22x1_ASAP7_75t_L g841 ( .A1(n_834), .A2(n_817), .B1(n_828), .B2(n_820), .Y(n_841) );
AOI22xp5_ASAP7_75t_L g842 ( .A1(n_839), .A2(n_810), .B1(n_803), .B2(n_819), .Y(n_842) );
INVx2_ASAP7_75t_L g843 ( .A(n_841), .Y(n_843) );
NAND2xp5_ASAP7_75t_L g844 ( .A(n_842), .B(n_810), .Y(n_844) );
CKINVDCx20_ASAP7_75t_R g845 ( .A(n_843), .Y(n_845) );
INVxp67_ASAP7_75t_SL g846 ( .A(n_845), .Y(n_846) );
INVx2_ASAP7_75t_L g847 ( .A(n_844), .Y(n_847) );
INVx1_ASAP7_75t_L g848 ( .A(n_846), .Y(n_848) );
INVx2_ASAP7_75t_L g849 ( .A(n_847), .Y(n_849) );
INVx1_ASAP7_75t_L g850 ( .A(n_848), .Y(n_850) );
INVx1_ASAP7_75t_L g851 ( .A(n_850), .Y(n_851) );
AO22x2_ASAP7_75t_L g852 ( .A1(n_851), .A2(n_849), .B1(n_840), .B2(n_821), .Y(n_852) );
INVx1_ASAP7_75t_L g853 ( .A(n_852), .Y(n_853) );
OAI22xp5_ASAP7_75t_L g854 ( .A1(n_853), .A2(n_849), .B1(n_828), .B2(n_816), .Y(n_854) );
INVx1_ASAP7_75t_L g855 ( .A(n_854), .Y(n_855) );
AOI221xp5_ASAP7_75t_L g856 ( .A1(n_855), .A2(n_835), .B1(n_833), .B2(n_838), .C(n_811), .Y(n_856) );
AOI22xp33_ASAP7_75t_L g857 ( .A1(n_856), .A2(n_811), .B1(n_827), .B2(n_830), .Y(n_857) );
endmodule