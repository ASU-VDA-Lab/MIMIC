module fake_jpeg_30384_n_101 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_101);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_101;

wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

BUFx12_ASAP7_75t_L g11 ( 
.A(n_9),
.Y(n_11)
);

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_6),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_9),
.Y(n_13)
);

BUFx3_ASAP7_75t_L g14 ( 
.A(n_2),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_0),
.Y(n_15)
);

INVx2_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

BUFx8_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_3),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_10),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_1),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_4),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_6),
.Y(n_22)
);

AOI21xp33_ASAP7_75t_L g23 ( 
.A1(n_15),
.A2(n_0),
.B(n_1),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_23),
.B(n_29),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_24),
.Y(n_32)
);

INVx5_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_25),
.Y(n_41)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_27),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_16),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_SL g30 ( 
.A(n_15),
.B(n_0),
.Y(n_30)
);

XNOR2xp5_ASAP7_75t_L g35 ( 
.A(n_30),
.B(n_20),
.Y(n_35)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_31),
.B(n_17),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_35),
.B(n_17),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_36),
.B(n_17),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_L g38 ( 
.A1(n_24),
.A2(n_20),
.B1(n_22),
.B2(n_21),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_38),
.A2(n_27),
.B1(n_24),
.B2(n_29),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g39 ( 
.A1(n_30),
.A2(n_14),
.B1(n_22),
.B2(n_13),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g46 ( 
.A1(n_39),
.A2(n_18),
.B1(n_21),
.B2(n_19),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_42),
.B(n_50),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g43 ( 
.A1(n_37),
.A2(n_26),
.B1(n_25),
.B2(n_28),
.Y(n_43)
);

INVxp67_ASAP7_75t_L g59 ( 
.A(n_43),
.Y(n_59)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_37),
.Y(n_44)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_44),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_34),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_45),
.B(n_49),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g61 ( 
.A1(n_46),
.A2(n_47),
.B1(n_52),
.B2(n_32),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g47 ( 
.A1(n_33),
.A2(n_31),
.B1(n_28),
.B2(n_27),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_40),
.Y(n_48)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_48),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_35),
.B(n_29),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_51),
.Y(n_63)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_32),
.Y(n_53)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_53),
.Y(n_64)
);

AND2x6_ASAP7_75t_L g54 ( 
.A(n_50),
.B(n_13),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_54),
.B(n_2),
.Y(n_70)
);

XOR2xp5_ASAP7_75t_L g60 ( 
.A(n_52),
.B(n_26),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_60),
.B(n_34),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_61),
.A2(n_53),
.B1(n_41),
.B2(n_17),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_48),
.A2(n_19),
.B1(n_18),
.B2(n_34),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_62),
.A2(n_41),
.B1(n_44),
.B2(n_51),
.Y(n_65)
);

OAI21xp5_ASAP7_75t_L g75 ( 
.A1(n_65),
.A2(n_59),
.B(n_17),
.Y(n_75)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_57),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_66),
.B(n_71),
.Y(n_76)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_64),
.Y(n_67)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_67),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_68),
.B(n_56),
.Y(n_80)
);

BUFx5_ASAP7_75t_L g69 ( 
.A(n_58),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_69),
.B(n_70),
.Y(n_79)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_63),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_72),
.B(n_73),
.Y(n_78)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_55),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_75),
.A2(n_11),
.B1(n_5),
.B2(n_7),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_SL g77 ( 
.A1(n_68),
.A2(n_59),
.B(n_54),
.Y(n_77)
);

OAI21xp5_ASAP7_75t_SL g86 ( 
.A1(n_77),
.A2(n_81),
.B(n_11),
.Y(n_86)
);

OAI21xp33_ASAP7_75t_L g82 ( 
.A1(n_80),
.A2(n_65),
.B(n_67),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_SL g81 ( 
.A1(n_69),
.A2(n_60),
.B(n_61),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_82),
.B(n_83),
.Y(n_89)
);

XOR2x1_ASAP7_75t_SL g83 ( 
.A(n_80),
.B(n_79),
.Y(n_83)
);

INVxp33_ASAP7_75t_L g84 ( 
.A(n_76),
.Y(n_84)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_84),
.Y(n_91)
);

HB1xp67_ASAP7_75t_L g85 ( 
.A(n_74),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_85),
.A2(n_87),
.B1(n_4),
.B2(n_5),
.Y(n_88)
);

O2A1O1Ixp33_ASAP7_75t_SL g90 ( 
.A1(n_86),
.A2(n_78),
.B(n_11),
.C(n_10),
.Y(n_90)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_88),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_90),
.B(n_7),
.Y(n_92)
);

NAND2xp33_ASAP7_75t_SL g97 ( 
.A(n_92),
.B(n_8),
.Y(n_97)
);

XOR2xp5_ASAP7_75t_L g94 ( 
.A(n_89),
.B(n_82),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_94),
.B(n_89),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_95),
.B(n_96),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_L g96 ( 
.A1(n_93),
.A2(n_91),
.B(n_8),
.Y(n_96)
);

NAND2x1_ASAP7_75t_L g99 ( 
.A(n_97),
.B(n_11),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_99),
.A2(n_11),
.B1(n_94),
.B2(n_98),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_100),
.B(n_99),
.Y(n_101)
);


endmodule