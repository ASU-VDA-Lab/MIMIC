module fake_jpeg_3410_n_210 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_210);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_210;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_207;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_202;
wire n_75;
wire n_122;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_91;
wire n_93;
wire n_54;
wire n_161;
wire n_209;
wire n_208;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx11_ASAP7_75t_SL g51 ( 
.A(n_29),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_45),
.B(n_42),
.Y(n_52)
);

BUFx4f_ASAP7_75t_SL g53 ( 
.A(n_23),
.Y(n_53)
);

BUFx5_ASAP7_75t_L g54 ( 
.A(n_12),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_20),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_22),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_6),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_36),
.Y(n_58)
);

INVx6_ASAP7_75t_SL g59 ( 
.A(n_34),
.Y(n_59)
);

BUFx5_ASAP7_75t_L g60 ( 
.A(n_1),
.Y(n_60)
);

BUFx5_ASAP7_75t_L g61 ( 
.A(n_6),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_2),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_19),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_7),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_3),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_0),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_2),
.Y(n_67)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_24),
.Y(n_68)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_25),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_26),
.Y(n_70)
);

BUFx5_ASAP7_75t_L g71 ( 
.A(n_11),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_43),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_28),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_50),
.Y(n_74)
);

BUFx12f_ASAP7_75t_L g75 ( 
.A(n_59),
.Y(n_75)
);

INVx8_ASAP7_75t_L g90 ( 
.A(n_75),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_55),
.Y(n_76)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_76),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_55),
.Y(n_77)
);

INVx6_ASAP7_75t_L g95 ( 
.A(n_77),
.Y(n_95)
);

INVx3_ASAP7_75t_SL g78 ( 
.A(n_51),
.Y(n_78)
);

BUFx2_ASAP7_75t_L g89 ( 
.A(n_78),
.Y(n_89)
);

INVx6_ASAP7_75t_L g79 ( 
.A(n_67),
.Y(n_79)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_79),
.Y(n_96)
);

CKINVDCx16_ASAP7_75t_R g80 ( 
.A(n_53),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_80),
.B(n_78),
.Y(n_93)
);

INVx5_ASAP7_75t_L g81 ( 
.A(n_59),
.Y(n_81)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_81),
.Y(n_85)
);

INVx11_ASAP7_75t_L g82 ( 
.A(n_51),
.Y(n_82)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_82),
.Y(n_92)
);

BUFx16f_ASAP7_75t_L g84 ( 
.A(n_78),
.Y(n_84)
);

INVxp67_ASAP7_75t_SL g105 ( 
.A(n_84),
.Y(n_105)
);

OAI21xp33_ASAP7_75t_L g86 ( 
.A1(n_80),
.A2(n_68),
.B(n_69),
.Y(n_86)
);

INVx1_ASAP7_75t_SL g113 ( 
.A(n_86),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_75),
.B(n_62),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_87),
.B(n_75),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_79),
.A2(n_69),
.B1(n_67),
.B2(n_68),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_88),
.A2(n_53),
.B1(n_77),
.B2(n_76),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_82),
.A2(n_64),
.B1(n_57),
.B2(n_65),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_91),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_93),
.B(n_94),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_82),
.A2(n_64),
.B1(n_66),
.B2(n_61),
.Y(n_94)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_96),
.Y(n_97)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_97),
.Y(n_116)
);

OAI32xp33_ASAP7_75t_L g98 ( 
.A1(n_86),
.A2(n_70),
.A3(n_52),
.B1(n_79),
.B2(n_60),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g133 ( 
.A(n_98),
.B(n_103),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_85),
.B(n_70),
.C(n_63),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_101),
.B(n_53),
.C(n_90),
.Y(n_120)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_84),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_102),
.Y(n_115)
);

AO22x1_ASAP7_75t_SL g104 ( 
.A1(n_96),
.A2(n_77),
.B1(n_76),
.B2(n_75),
.Y(n_104)
);

AND2x2_ASAP7_75t_L g135 ( 
.A(n_104),
.B(n_27),
.Y(n_135)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_83),
.Y(n_106)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_106),
.Y(n_123)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_84),
.Y(n_107)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_107),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_108),
.A2(n_95),
.B1(n_83),
.B2(n_81),
.Y(n_121)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_92),
.Y(n_109)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_109),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_85),
.B(n_73),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_110),
.B(n_111),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_90),
.B(n_74),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_89),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_112),
.B(n_92),
.Y(n_119)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_89),
.Y(n_114)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_114),
.Y(n_132)
);

AOI32xp33_ASAP7_75t_L g117 ( 
.A1(n_100),
.A2(n_56),
.A3(n_58),
.B1(n_72),
.B2(n_54),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_117),
.B(n_120),
.Y(n_154)
);

CKINVDCx14_ASAP7_75t_R g118 ( 
.A(n_113),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_118),
.B(n_129),
.Y(n_144)
);

CKINVDCx16_ASAP7_75t_R g152 ( 
.A(n_119),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_L g159 ( 
.A1(n_121),
.A2(n_31),
.B1(n_47),
.B2(n_46),
.Y(n_159)
);

BUFx24_ASAP7_75t_L g122 ( 
.A(n_105),
.Y(n_122)
);

INVx2_ASAP7_75t_SL g140 ( 
.A(n_122),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_102),
.B(n_107),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g145 ( 
.A(n_125),
.B(n_127),
.Y(n_145)
);

NOR2x1_ASAP7_75t_L g127 ( 
.A(n_113),
.B(n_81),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_105),
.B(n_0),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_99),
.A2(n_95),
.B1(n_71),
.B2(n_61),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_130),
.A2(n_135),
.B1(n_3),
.B2(n_4),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_99),
.A2(n_71),
.B1(n_60),
.B2(n_54),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_131),
.A2(n_5),
.B1(n_7),
.B2(n_8),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_109),
.B(n_1),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_134),
.B(n_8),
.Y(n_147)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_128),
.Y(n_136)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_136),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_133),
.A2(n_104),
.B1(n_4),
.B2(n_5),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_137),
.A2(n_14),
.B1(n_15),
.B2(n_16),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_115),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_138),
.B(n_139),
.Y(n_170)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_132),
.Y(n_139)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_123),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_141),
.B(n_146),
.Y(n_175)
);

INVxp67_ASAP7_75t_L g168 ( 
.A(n_142),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_143),
.A2(n_156),
.B1(n_159),
.B2(n_13),
.Y(n_169)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_116),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_147),
.B(n_148),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_133),
.B(n_32),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_124),
.Y(n_149)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_149),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_115),
.Y(n_150)
);

AOI322xp5_ASAP7_75t_SL g165 ( 
.A1(n_150),
.A2(n_151),
.A3(n_157),
.B1(n_158),
.B2(n_9),
.C1(n_10),
.C2(n_12),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_126),
.Y(n_151)
);

INVx3_ASAP7_75t_L g153 ( 
.A(n_122),
.Y(n_153)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_153),
.Y(n_167)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_127),
.Y(n_155)
);

INVxp33_ASAP7_75t_L g176 ( 
.A(n_155),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_135),
.B(n_49),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_122),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_130),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_152),
.A2(n_120),
.B1(n_10),
.B2(n_11),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_160),
.A2(n_166),
.B1(n_174),
.B2(n_140),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_148),
.B(n_30),
.C(n_44),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_161),
.B(n_164),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_SL g164 ( 
.A1(n_144),
.A2(n_21),
.B(n_41),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_165),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_142),
.A2(n_9),
.B1(n_13),
.B2(n_14),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_169),
.B(n_171),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_136),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_172),
.A2(n_177),
.B1(n_159),
.B2(n_156),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_145),
.A2(n_48),
.B1(n_35),
.B2(n_37),
.Y(n_173)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_173),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_L g174 ( 
.A1(n_154),
.A2(n_15),
.B(n_16),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_137),
.A2(n_17),
.B1(n_18),
.B2(n_33),
.Y(n_177)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_179),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_SL g180 ( 
.A(n_178),
.B(n_147),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_180),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_182),
.B(n_186),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_175),
.Y(n_185)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_185),
.Y(n_194)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_170),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_162),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_187),
.B(n_174),
.C(n_163),
.Y(n_189)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_189),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_188),
.B(n_161),
.C(n_160),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_190),
.B(n_192),
.Y(n_200)
);

AOI322xp5_ASAP7_75t_L g192 ( 
.A1(n_181),
.A2(n_168),
.A3(n_176),
.B1(n_172),
.B2(n_167),
.C1(n_177),
.C2(n_173),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_182),
.B(n_176),
.Y(n_195)
);

AND2x2_ASAP7_75t_L g198 ( 
.A(n_195),
.B(n_140),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_198),
.B(n_191),
.Y(n_204)
);

AOI31xp67_ASAP7_75t_L g199 ( 
.A1(n_194),
.A2(n_183),
.A3(n_168),
.B(n_184),
.Y(n_199)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_199),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_193),
.A2(n_183),
.B1(n_153),
.B2(n_184),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_201),
.B(n_195),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_202),
.B(n_204),
.Y(n_206)
);

AOI21xp5_ASAP7_75t_L g205 ( 
.A1(n_203),
.A2(n_200),
.B(n_197),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_SL g207 ( 
.A(n_205),
.B(n_196),
.Y(n_207)
);

NOR4xp25_ASAP7_75t_L g208 ( 
.A(n_207),
.B(n_206),
.C(n_192),
.D(n_17),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_208),
.B(n_40),
.Y(n_209)
);

AOI21xp5_ASAP7_75t_L g210 ( 
.A1(n_209),
.A2(n_38),
.B(n_39),
.Y(n_210)
);


endmodule