module fake_jpeg_31258_n_5 (n_0, n_1, n_5);

input n_0;
input n_1;

output n_5;

wire n_3;
wire n_2;
wire n_4;

INVx2_ASAP7_75t_L g2 ( 
.A(n_0),
.Y(n_2)
);

HB1xp67_ASAP7_75t_L g3 ( 
.A(n_2),
.Y(n_3)
);

NAND2xp5_ASAP7_75t_L g4 ( 
.A(n_3),
.B(n_1),
.Y(n_4)
);

BUFx24_ASAP7_75t_SL g5 ( 
.A(n_4),
.Y(n_5)
);


endmodule