module fake_netlist_5_2225_n_1983 (n_137, n_168, n_164, n_191, n_91, n_82, n_122, n_194, n_142, n_176, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_182, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_180, n_184, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_189, n_165, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_177, n_60, n_155, n_152, n_197, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_195, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_203, n_205, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_179, n_125, n_35, n_167, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_202, n_130, n_157, n_29, n_79, n_193, n_131, n_151, n_47, n_173, n_192, n_25, n_53, n_160, n_198, n_188, n_190, n_8, n_201, n_158, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_159, n_163, n_95, n_119, n_183, n_185, n_175, n_169, n_59, n_26, n_133, n_55, n_196, n_99, n_2, n_181, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_178, n_12, n_67, n_121, n_36, n_76, n_200, n_87, n_150, n_162, n_27, n_170, n_64, n_77, n_102, n_106, n_161, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_174, n_186, n_199, n_134, n_187, n_32, n_41, n_104, n_172, n_103, n_56, n_51, n_63, n_97, n_141, n_166, n_11, n_171, n_153, n_7, n_15, n_145, n_48, n_204, n_50, n_52, n_88, n_110, n_1983);

input n_137;
input n_168;
input n_164;
input n_191;
input n_91;
input n_82;
input n_122;
input n_194;
input n_142;
input n_176;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_182;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_180;
input n_184;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_189;
input n_165;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_177;
input n_60;
input n_155;
input n_152;
input n_197;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_195;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_203;
input n_205;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_179;
input n_125;
input n_35;
input n_167;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_202;
input n_130;
input n_157;
input n_29;
input n_79;
input n_193;
input n_131;
input n_151;
input n_47;
input n_173;
input n_192;
input n_25;
input n_53;
input n_160;
input n_198;
input n_188;
input n_190;
input n_8;
input n_201;
input n_158;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_159;
input n_163;
input n_95;
input n_119;
input n_183;
input n_185;
input n_175;
input n_169;
input n_59;
input n_26;
input n_133;
input n_55;
input n_196;
input n_99;
input n_2;
input n_181;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_178;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_200;
input n_87;
input n_150;
input n_162;
input n_27;
input n_170;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_174;
input n_186;
input n_199;
input n_134;
input n_187;
input n_32;
input n_41;
input n_104;
input n_172;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_166;
input n_11;
input n_171;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_204;
input n_50;
input n_52;
input n_88;
input n_110;

output n_1983;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1729;
wire n_1166;
wire n_1751;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1859;
wire n_1677;
wire n_1150;
wire n_226;
wire n_1780;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1738;
wire n_1021;
wire n_1960;
wire n_551;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1695;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_1789;
wire n_1666;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_1545;
wire n_864;
wire n_859;
wire n_951;
wire n_1947;
wire n_1264;
wire n_447;
wire n_247;
wire n_1494;
wire n_292;
wire n_625;
wire n_854;
wire n_1462;
wire n_1799;
wire n_1580;
wire n_674;
wire n_417;
wire n_1939;
wire n_1806;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_1869;
wire n_1607;
wire n_1563;
wire n_606;
wire n_275;
wire n_877;
wire n_1696;
wire n_755;
wire n_1118;
wire n_1686;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1860;
wire n_1359;
wire n_530;
wire n_1107;
wire n_1728;
wire n_556;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_1896;
wire n_929;
wire n_1124;
wire n_1818;
wire n_902;
wire n_1576;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1705;
wire n_1257;
wire n_1182;
wire n_579;
wire n_1698;
wire n_1261;
wire n_938;
wire n_1098;
wire n_320;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_519;
wire n_406;
wire n_1016;
wire n_1243;
wire n_546;
wire n_1280;
wire n_1845;
wire n_281;
wire n_240;
wire n_291;
wire n_231;
wire n_257;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_317;
wire n_1236;
wire n_1633;
wire n_569;
wire n_1778;
wire n_227;
wire n_920;
wire n_1289;
wire n_1517;
wire n_335;
wire n_1669;
wire n_370;
wire n_976;
wire n_1949;
wire n_343;
wire n_1449;
wire n_308;
wire n_1946;
wire n_1566;
wire n_297;
wire n_1078;
wire n_1670;
wire n_775;
wire n_219;
wire n_600;
wire n_1484;
wire n_1374;
wire n_1328;
wire n_223;
wire n_1948;
wire n_264;
wire n_1877;
wire n_1831;
wire n_1598;
wire n_1723;
wire n_955;
wire n_1850;
wire n_339;
wire n_1146;
wire n_882;
wire n_243;
wire n_1036;
wire n_1097;
wire n_1749;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_215;
wire n_350;
wire n_798;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_290;
wire n_580;
wire n_1040;
wire n_1872;
wire n_1852;
wire n_578;
wire n_926;
wire n_344;
wire n_1218;
wire n_1931;
wire n_422;
wire n_475;
wire n_777;
wire n_1070;
wire n_1547;
wire n_1030;
wire n_1755;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1801;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_845;
wire n_663;
wire n_1862;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_1796;
wire n_680;
wire n_1473;
wire n_1587;
wire n_395;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_214;
wire n_1748;
wire n_1672;
wire n_675;
wire n_888;
wire n_1880;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1384;
wire n_1556;
wire n_446;
wire n_1863;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_1706;
wire n_468;
wire n_213;
wire n_342;
wire n_464;
wire n_363;
wire n_1582;
wire n_1069;
wire n_1784;
wire n_1075;
wire n_1836;
wire n_1450;
wire n_1322;
wire n_1471;
wire n_1750;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_1700;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1971;
wire n_1599;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_1950;
wire n_907;
wire n_1447;
wire n_1377;
wire n_989;
wire n_1039;
wire n_228;
wire n_283;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_310;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_1667;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1926;
wire n_1248;
wire n_230;
wire n_1331;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_1819;
wire n_476;
wire n_1527;
wire n_534;
wire n_1882;
wire n_884;
wire n_345;
wire n_944;
wire n_1754;
wire n_1623;
wire n_1854;
wire n_1565;
wire n_1809;
wire n_1856;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_857;
wire n_832;
wire n_207;
wire n_561;
wire n_1319;
wire n_1825;
wire n_1951;
wire n_1883;
wire n_1906;
wire n_1712;
wire n_1387;
wire n_1532;
wire n_1027;
wire n_971;
wire n_1156;
wire n_326;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1775;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_1709;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1538;
wire n_1838;
wire n_1199;
wire n_1847;
wire n_1779;
wire n_352;
wire n_1884;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_1841;
wire n_1660;
wire n_887;
wire n_1905;
wire n_300;
wire n_809;
wire n_870;
wire n_931;
wire n_599;
wire n_1891;
wire n_1662;
wire n_1711;
wire n_1481;
wire n_1942;
wire n_434;
wire n_1978;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1629;
wire n_1293;
wire n_965;
wire n_1876;
wire n_1743;
wire n_935;
wire n_1175;
wire n_817;
wire n_360;
wire n_1479;
wire n_1810;
wire n_1888;
wire n_759;
wire n_1892;
wire n_806;
wire n_1766;
wire n_1477;
wire n_324;
wire n_1635;
wire n_1963;
wire n_1571;
wire n_1189;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_784;
wire n_1733;
wire n_1244;
wire n_431;
wire n_1194;
wire n_1925;
wire n_1815;
wire n_615;
wire n_851;
wire n_1759;
wire n_843;
wire n_1788;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_1679;
wire n_776;
wire n_1798;
wire n_1790;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1746;
wire n_1647;
wire n_1829;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_1674;
wire n_1833;
wire n_1830;
wire n_1710;
wire n_284;
wire n_1128;
wire n_1734;
wire n_744;
wire n_590;
wire n_629;
wire n_1308;
wire n_1767;
wire n_254;
wire n_1680;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_526;
wire n_1916;
wire n_372;
wire n_293;
wire n_677;
wire n_244;
wire n_1333;
wire n_1121;
wire n_433;
wire n_314;
wire n_604;
wire n_368;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_498;
wire n_1468;
wire n_1559;
wire n_1765;
wire n_1866;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_252;
wire n_624;
wire n_1380;
wire n_1744;
wire n_1617;
wire n_295;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_1839;
wire n_1837;
wire n_610;
wire n_1760;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_1832;
wire n_259;
wire n_448;
wire n_1851;
wire n_758;
wire n_999;
wire n_1933;
wire n_1656;
wire n_1158;
wire n_1509;
wire n_1874;
wire n_563;
wire n_1145;
wire n_878;
wire n_524;
wire n_394;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_1871;
wire n_1964;
wire n_331;
wire n_906;
wire n_1163;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_1781;
wire n_658;
wire n_1740;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_1923;
wire n_1773;
wire n_592;
wire n_1169;
wire n_1596;
wire n_1692;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_1095;
wire n_1828;
wire n_1614;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_1431;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1640;
wire n_1732;
wire n_1009;
wire n_1148;
wire n_742;
wire n_750;
wire n_995;
wire n_454;
wire n_1609;
wire n_374;
wire n_396;
wire n_1887;
wire n_1383;
wire n_1073;
wire n_255;
wire n_662;
wire n_459;
wire n_218;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1920;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1721;
wire n_1959;
wire n_1758;
wire n_1574;
wire n_473;
wire n_1921;
wire n_1309;
wire n_1878;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_1800;
wire n_1548;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_208;
wire n_743;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_1240;
wire n_1820;
wire n_829;
wire n_1612;
wire n_1416;
wire n_1724;
wire n_361;
wire n_700;
wire n_1237;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1785;
wire n_1568;
wire n_1006;
wire n_329;
wire n_274;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_1870;
wire n_309;
wire n_512;
wire n_1591;
wire n_322;
wire n_1682;
wire n_1980;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1927;
wire n_1349;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_1909;
wire n_224;
wire n_1562;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_1965;
wire n_239;
wire n_630;
wire n_1902;
wire n_1941;
wire n_1913;
wire n_504;
wire n_1823;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_1875;
wire n_1982;
wire n_1304;
wire n_1324;
wire n_987;
wire n_1846;
wire n_261;
wire n_1885;
wire n_1455;
wire n_767;
wire n_993;
wire n_1903;
wire n_1407;
wire n_1551;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_1805;
wire n_1816;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_1849;
wire n_729;
wire n_1131;
wire n_1084;
wire n_1961;
wire n_970;
wire n_1935;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_340;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_1645;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_1684;
wire n_233;
wire n_1717;
wire n_572;
wire n_366;
wire n_815;
wire n_1795;
wire n_1821;
wire n_327;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_1708;
wire n_426;
wire n_1438;
wire n_1082;
wire n_1840;
wire n_589;
wire n_716;
wire n_1630;
wire n_562;
wire n_1436;
wire n_1691;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_1776;
wire n_531;
wire n_1757;
wire n_890;
wire n_1897;
wire n_764;
wire n_1919;
wire n_1056;
wire n_1424;
wire n_960;
wire n_1893;
wire n_222;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_634;
wire n_1958;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_1519;
wire n_256;
wire n_950;
wire n_1553;
wire n_1811;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1808;
wire n_1060;
wire n_1141;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_912;
wire n_315;
wire n_968;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_1699;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_1954;
wire n_1608;
wire n_983;
wire n_1844;
wire n_280;
wire n_1305;
wire n_873;
wire n_1826;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_1644;
wire n_690;
wire n_1974;
wire n_583;
wire n_302;
wire n_1343;
wire n_1203;
wire n_1631;
wire n_821;
wire n_1763;
wire n_1966;
wire n_1768;
wire n_321;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1719;
wire n_1288;
wire n_385;
wire n_212;
wire n_507;
wire n_1560;
wire n_1605;
wire n_330;
wire n_1228;
wire n_972;
wire n_692;
wire n_1953;
wire n_1938;
wire n_820;
wire n_1200;
wire n_1911;
wire n_1301;
wire n_1363;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_1967;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_1688;
wire n_945;
wire n_492;
wire n_1504;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_1932;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_286;
wire n_1643;
wire n_883;
wire n_470;
wire n_325;
wire n_449;
wire n_1594;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_856;
wire n_1793;
wire n_1976;
wire n_918;
wire n_942;
wire n_1804;
wire n_1147;
wire n_1557;
wire n_1977;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_356;
wire n_894;
wire n_1636;
wire n_1730;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1865;
wire n_1470;
wire n_1096;
wire n_234;
wire n_1575;
wire n_1697;
wire n_1735;
wire n_833;
wire n_1646;
wire n_225;
wire n_1307;
wire n_1881;
wire n_988;
wire n_1940;
wire n_814;
wire n_1549;
wire n_1934;
wire n_1201;
wire n_1114;
wire n_655;
wire n_1616;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_1807;
wire n_387;
wire n_1149;
wire n_398;
wire n_1671;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_211;
wire n_1824;
wire n_1917;
wire n_1219;
wire n_1204;
wire n_1814;
wire n_1035;
wire n_287;
wire n_555;
wire n_783;
wire n_1848;
wire n_1928;
wire n_1188;
wire n_1722;
wire n_661;
wire n_1802;
wire n_849;
wire n_584;
wire n_336;
wire n_681;
wire n_1638;
wire n_1786;
wire n_430;
wire n_510;
wire n_216;
wire n_311;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_1655;
wire n_445;
wire n_749;
wire n_1895;
wire n_1134;
wire n_1358;
wire n_717;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_249;
wire n_304;
wire n_1338;
wire n_577;
wire n_1522;
wire n_1687;
wire n_1637;
wire n_1419;
wire n_338;
wire n_1653;
wire n_693;
wire n_1506;
wire n_836;
wire n_990;
wire n_1886;
wire n_1389;
wire n_1894;
wire n_975;
wire n_1908;
wire n_1256;
wire n_1702;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_306;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_1843;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1929;
wire n_1164;
wire n_1659;
wire n_1834;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_1572;
wire n_1968;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1736;
wire n_1685;
wire n_601;
wire n_917;
wire n_1714;
wire n_966;
wire n_253;
wire n_1116;
wire n_1661;
wire n_1212;
wire n_1541;
wire n_206;
wire n_217;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_1731;
wire n_818;
wire n_1970;
wire n_861;
wire n_1713;
wire n_1183;
wire n_1658;
wire n_899;
wire n_1253;
wire n_210;
wire n_1737;
wire n_1904;
wire n_774;
wire n_1628;
wire n_1335;
wire n_1514;
wire n_1777;
wire n_1957;
wire n_1059;
wire n_1345;
wire n_1133;
wire n_1771;
wire n_1912;
wire n_1899;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_1168;
wire n_707;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_1584;
wire n_665;
wire n_1726;
wire n_1835;
wire n_1440;
wire n_421;
wire n_1853;
wire n_1356;
wire n_1787;
wire n_910;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1774;
wire n_1725;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_1812;
wire n_735;
wire n_232;
wire n_1915;
wire n_1109;
wire n_895;
wire n_1310;
wire n_1803;
wire n_427;
wire n_1399;
wire n_1543;
wire n_1979;
wire n_791;
wire n_732;
wire n_1533;
wire n_808;
wire n_797;
wire n_1025;
wire n_1930;
wire n_1955;
wire n_500;
wire n_1067;
wire n_1720;
wire n_435;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1742;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_594;
wire n_1291;
wire n_1297;
wire n_1753;
wire n_1782;
wire n_1155;
wire n_1418;
wire n_1972;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_985;
wire n_1855;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1703;
wire n_1352;
wire n_626;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_305;
wire n_676;
wire n_294;
wire n_318;
wire n_653;
wire n_642;
wire n_1602;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_268;
wire n_664;
wire n_503;
wire n_235;
wire n_1372;
wire n_605;
wire n_1273;
wire n_1822;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_1783;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_1907;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_1898;
wire n_581;
wire n_382;
wire n_554;
wire n_1625;
wire n_898;
wire n_1762;
wire n_1013;
wire n_1452;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_1791;
wire n_1890;
wire n_1747;
wire n_714;
wire n_1683;
wire n_1817;
wire n_909;
wire n_1944;
wire n_1530;
wire n_1497;
wire n_997;
wire n_932;
wire n_612;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_1981;
wire n_508;
wire n_506;
wire n_1320;
wire n_1663;
wire n_737;
wire n_1718;
wire n_986;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1715;
wire n_1281;
wire n_1952;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_1889;
wire n_209;
wire n_1792;
wire n_1564;
wire n_1868;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1922;
wire n_1376;
wire n_941;
wire n_981;
wire n_1569;
wire n_867;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_518;
wire n_505;
wire n_1772;
wire n_282;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1861;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1901;
wire n_1900;
wire n_1620;
wire n_381;
wire n_220;
wire n_390;
wire n_1330;
wire n_1867;
wire n_1945;
wire n_481;
wire n_1675;
wire n_1924;
wire n_1727;
wire n_1554;
wire n_1745;
wire n_769;
wire n_1046;
wire n_271;
wire n_934;
wire n_1618;
wire n_826;
wire n_1813;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_428;
wire n_379;
wire n_1341;
wire n_570;
wire n_1641;
wire n_1361;
wire n_1707;
wire n_853;
wire n_377;
wire n_751;
wire n_1973;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_704;
wire n_787;
wire n_1770;
wire n_961;
wire n_1756;
wire n_771;
wire n_276;
wire n_1716;
wire n_1225;
wire n_1520;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_1873;
wire n_1411;
wire n_221;
wire n_622;
wire n_1962;
wire n_1577;
wire n_1087;
wire n_386;
wire n_994;
wire n_1701;
wire n_848;
wire n_1550;
wire n_1498;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1857;
wire n_1344;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_1797;
wire n_432;
wire n_1769;
wire n_839;
wire n_1210;
wire n_1364;
wire n_328;
wire n_1250;
wire n_369;
wire n_1842;
wire n_871;
wire n_685;
wire n_598;
wire n_928;
wire n_608;
wire n_1367;
wire n_1943;
wire n_1460;
wire n_772;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_413;
wire n_402;
wire n_1086;
wire n_796;
wire n_1858;
wire n_1619;
wire n_236;
wire n_1502;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_903;
wire n_1525;
wire n_1752;
wire n_740;
wire n_384;
wire n_1404;
wire n_1794;
wire n_1315;
wire n_277;
wire n_1061;
wire n_1910;
wire n_333;
wire n_1298;
wire n_1652;
wire n_462;
wire n_1193;
wire n_1676;
wire n_1255;
wire n_258;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_844;
wire n_471;
wire n_852;
wire n_1487;
wire n_1864;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_1673;
wire n_465;
wire n_362;
wire n_1321;
wire n_1975;
wire n_273;
wire n_1937;
wire n_585;
wire n_1739;
wire n_270;
wire n_616;
wire n_1914;
wire n_745;
wire n_1654;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_1761;
wire n_641;
wire n_730;
wire n_1325;
wire n_1595;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_229;
wire n_1936;
wire n_1956;
wire n_437;
wire n_1642;
wire n_453;
wire n_403;
wire n_1130;
wire n_720;
wire n_1918;
wire n_1526;
wire n_863;
wire n_805;
wire n_1604;
wire n_1275;
wire n_1764;
wire n_712;
wire n_246;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_269;
wire n_285;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1741;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_1621;
wire n_251;
wire n_566;
wire n_565;
wire n_1448;
wire n_1507;
wire n_1398;
wire n_1879;
wire n_597;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_651;
wire n_1340;
wire n_334;
wire n_811;
wire n_1558;
wire n_807;
wire n_835;
wire n_666;
wire n_262;
wire n_1433;
wire n_1704;
wire n_1254;
wire n_1026;
wire n_1969;
wire n_1234;
wire n_319;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_242;
wire n_1681;
wire n_1018;
wire n_1693;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_1180;
wire n_1827;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;
wire n_278;

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_187),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_141),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_23),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_176),
.Y(n_209)
);

INVx1_ASAP7_75t_SL g210 ( 
.A(n_191),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_79),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_12),
.Y(n_212)
);

INVx3_ASAP7_75t_L g213 ( 
.A(n_101),
.Y(n_213)
);

CKINVDCx16_ASAP7_75t_R g214 ( 
.A(n_19),
.Y(n_214)
);

BUFx3_ASAP7_75t_L g215 ( 
.A(n_86),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_22),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_90),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_71),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_55),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_120),
.Y(n_220)
);

BUFx6f_ASAP7_75t_L g221 ( 
.A(n_173),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_148),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_47),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_134),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_24),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_106),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_41),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_61),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_23),
.Y(n_229)
);

HB1xp67_ASAP7_75t_L g230 ( 
.A(n_117),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_159),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_59),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_123),
.Y(n_233)
);

CKINVDCx16_ASAP7_75t_R g234 ( 
.A(n_24),
.Y(n_234)
);

BUFx10_ASAP7_75t_L g235 ( 
.A(n_161),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_169),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_64),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_20),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_143),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_105),
.Y(n_240)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_131),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_93),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_55),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_183),
.Y(n_244)
);

BUFx6f_ASAP7_75t_L g245 ( 
.A(n_132),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_7),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_188),
.Y(n_247)
);

BUFx2_ASAP7_75t_L g248 ( 
.A(n_66),
.Y(n_248)
);

INVx1_ASAP7_75t_SL g249 ( 
.A(n_153),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_94),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_56),
.Y(n_251)
);

BUFx3_ASAP7_75t_L g252 ( 
.A(n_170),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_51),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_158),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_195),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_78),
.Y(n_256)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_139),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_20),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_128),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_172),
.Y(n_260)
);

INVx2_ASAP7_75t_SL g261 ( 
.A(n_180),
.Y(n_261)
);

BUFx6f_ASAP7_75t_L g262 ( 
.A(n_177),
.Y(n_262)
);

BUFx5_ASAP7_75t_L g263 ( 
.A(n_89),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_103),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_11),
.Y(n_265)
);

BUFx3_ASAP7_75t_L g266 ( 
.A(n_10),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_174),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_202),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_185),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_107),
.Y(n_270)
);

INVx2_ASAP7_75t_SL g271 ( 
.A(n_127),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_74),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_114),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_178),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_160),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_5),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_190),
.Y(n_277)
);

BUFx10_ASAP7_75t_L g278 ( 
.A(n_34),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_29),
.Y(n_279)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_167),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_49),
.Y(n_281)
);

INVx1_ASAP7_75t_SL g282 ( 
.A(n_137),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_0),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_164),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_66),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_44),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_77),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_21),
.Y(n_288)
);

CKINVDCx16_ASAP7_75t_R g289 ( 
.A(n_3),
.Y(n_289)
);

INVx2_ASAP7_75t_SL g290 ( 
.A(n_16),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_201),
.Y(n_291)
);

BUFx10_ASAP7_75t_L g292 ( 
.A(n_75),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_196),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_133),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_73),
.Y(n_295)
);

CKINVDCx14_ASAP7_75t_R g296 ( 
.A(n_13),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_150),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_108),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_163),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_154),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_43),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_113),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_88),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_49),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_96),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_166),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_192),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_126),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_81),
.Y(n_309)
);

BUFx10_ASAP7_75t_L g310 ( 
.A(n_41),
.Y(n_310)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_186),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_122),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_142),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_12),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_72),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_44),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_5),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_82),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_109),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_175),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_9),
.Y(n_321)
);

INVx1_ASAP7_75t_SL g322 ( 
.A(n_43),
.Y(n_322)
);

BUFx10_ASAP7_75t_L g323 ( 
.A(n_28),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_1),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_121),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_46),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_10),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_48),
.Y(n_328)
);

CKINVDCx16_ASAP7_75t_R g329 ( 
.A(n_69),
.Y(n_329)
);

BUFx6f_ASAP7_75t_L g330 ( 
.A(n_27),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_145),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_84),
.Y(n_332)
);

BUFx6f_ASAP7_75t_L g333 ( 
.A(n_45),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_4),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_50),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_146),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_85),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_3),
.Y(n_338)
);

INVx2_ASAP7_75t_L g339 ( 
.A(n_60),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_70),
.Y(n_340)
);

BUFx2_ASAP7_75t_SL g341 ( 
.A(n_26),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_184),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_14),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_48),
.Y(n_344)
);

BUFx10_ASAP7_75t_L g345 ( 
.A(n_182),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_29),
.Y(n_346)
);

BUFx3_ASAP7_75t_L g347 ( 
.A(n_168),
.Y(n_347)
);

INVx1_ASAP7_75t_SL g348 ( 
.A(n_47),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_45),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_13),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_198),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_87),
.Y(n_352)
);

INVx2_ASAP7_75t_SL g353 ( 
.A(n_67),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_136),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_9),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_203),
.Y(n_356)
);

INVx1_ASAP7_75t_SL g357 ( 
.A(n_165),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_147),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_1),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_193),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_155),
.Y(n_361)
);

INVx2_ASAP7_75t_SL g362 ( 
.A(n_32),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_25),
.Y(n_363)
);

BUFx10_ASAP7_75t_L g364 ( 
.A(n_116),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_68),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_34),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_100),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_56),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_35),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_28),
.Y(n_370)
);

CKINVDCx20_ASAP7_75t_R g371 ( 
.A(n_189),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_50),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_61),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_197),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_19),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_17),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_91),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_30),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_16),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_111),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_157),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_37),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_33),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_194),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_17),
.Y(n_385)
);

INVx1_ASAP7_75t_SL g386 ( 
.A(n_95),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_144),
.Y(n_387)
);

INVx2_ASAP7_75t_SL g388 ( 
.A(n_130),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_102),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_25),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_138),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_51),
.Y(n_392)
);

INVx2_ASAP7_75t_L g393 ( 
.A(n_39),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_204),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_151),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_135),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_92),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_156),
.Y(n_398)
);

INVx1_ASAP7_75t_SL g399 ( 
.A(n_15),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_26),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_15),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_39),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_4),
.Y(n_403)
);

BUFx6f_ASAP7_75t_L g404 ( 
.A(n_52),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_129),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_31),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_38),
.Y(n_407)
);

CKINVDCx20_ASAP7_75t_R g408 ( 
.A(n_217),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_207),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_211),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_L g411 ( 
.A(n_230),
.B(n_0),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_330),
.Y(n_412)
);

CKINVDCx20_ASAP7_75t_R g413 ( 
.A(n_217),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_330),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_254),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_255),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_330),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_330),
.Y(n_418)
);

INVx2_ASAP7_75t_L g419 ( 
.A(n_330),
.Y(n_419)
);

NOR2xp33_ASAP7_75t_L g420 ( 
.A(n_296),
.B(n_2),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_259),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_333),
.Y(n_422)
);

CKINVDCx20_ASAP7_75t_R g423 ( 
.A(n_247),
.Y(n_423)
);

NOR2xp67_ASAP7_75t_L g424 ( 
.A(n_213),
.B(n_2),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_260),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_333),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_333),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_333),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_333),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_404),
.Y(n_430)
);

INVxp67_ASAP7_75t_SL g431 ( 
.A(n_215),
.Y(n_431)
);

HB1xp67_ASAP7_75t_L g432 ( 
.A(n_214),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_404),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_404),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_264),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_268),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_404),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_404),
.Y(n_438)
);

INVxp33_ASAP7_75t_SL g439 ( 
.A(n_223),
.Y(n_439)
);

BUFx6f_ASAP7_75t_SL g440 ( 
.A(n_235),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_339),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_273),
.Y(n_442)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_263),
.Y(n_443)
);

CKINVDCx20_ASAP7_75t_R g444 ( 
.A(n_247),
.Y(n_444)
);

INVxp33_ASAP7_75t_SL g445 ( 
.A(n_223),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_274),
.Y(n_446)
);

CKINVDCx20_ASAP7_75t_R g447 ( 
.A(n_275),
.Y(n_447)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_263),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_339),
.Y(n_449)
);

CKINVDCx20_ASAP7_75t_R g450 ( 
.A(n_275),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_393),
.Y(n_451)
);

CKINVDCx20_ASAP7_75t_R g452 ( 
.A(n_297),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_277),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_284),
.Y(n_454)
);

HB1xp67_ASAP7_75t_L g455 ( 
.A(n_234),
.Y(n_455)
);

INVx2_ASAP7_75t_L g456 ( 
.A(n_263),
.Y(n_456)
);

CKINVDCx20_ASAP7_75t_R g457 ( 
.A(n_297),
.Y(n_457)
);

CKINVDCx20_ASAP7_75t_R g458 ( 
.A(n_371),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_294),
.Y(n_459)
);

INVxp67_ASAP7_75t_SL g460 ( 
.A(n_215),
.Y(n_460)
);

INVxp67_ASAP7_75t_SL g461 ( 
.A(n_252),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_393),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_295),
.Y(n_463)
);

CKINVDCx20_ASAP7_75t_R g464 ( 
.A(n_371),
.Y(n_464)
);

CKINVDCx5p33_ASAP7_75t_R g465 ( 
.A(n_298),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_266),
.Y(n_466)
);

INVxp67_ASAP7_75t_L g467 ( 
.A(n_248),
.Y(n_467)
);

CKINVDCx5p33_ASAP7_75t_R g468 ( 
.A(n_299),
.Y(n_468)
);

CKINVDCx20_ASAP7_75t_R g469 ( 
.A(n_329),
.Y(n_469)
);

CKINVDCx5p33_ASAP7_75t_R g470 ( 
.A(n_302),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_266),
.Y(n_471)
);

CKINVDCx5p33_ASAP7_75t_R g472 ( 
.A(n_303),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_407),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_216),
.Y(n_474)
);

BUFx2_ASAP7_75t_L g475 ( 
.A(n_227),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_219),
.Y(n_476)
);

CKINVDCx5p33_ASAP7_75t_R g477 ( 
.A(n_305),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_225),
.Y(n_478)
);

NOR2xp67_ASAP7_75t_L g479 ( 
.A(n_213),
.B(n_6),
.Y(n_479)
);

CKINVDCx5p33_ASAP7_75t_R g480 ( 
.A(n_306),
.Y(n_480)
);

CKINVDCx14_ASAP7_75t_R g481 ( 
.A(n_278),
.Y(n_481)
);

INVxp67_ASAP7_75t_L g482 ( 
.A(n_278),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_232),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_237),
.Y(n_484)
);

INVxp67_ASAP7_75t_SL g485 ( 
.A(n_252),
.Y(n_485)
);

CKINVDCx5p33_ASAP7_75t_R g486 ( 
.A(n_307),
.Y(n_486)
);

CKINVDCx5p33_ASAP7_75t_R g487 ( 
.A(n_308),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_243),
.Y(n_488)
);

CKINVDCx5p33_ASAP7_75t_R g489 ( 
.A(n_309),
.Y(n_489)
);

NOR2xp33_ASAP7_75t_L g490 ( 
.A(n_261),
.B(n_6),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_246),
.Y(n_491)
);

AND2x2_ASAP7_75t_L g492 ( 
.A(n_290),
.B(n_7),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_265),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_276),
.Y(n_494)
);

BUFx3_ASAP7_75t_L g495 ( 
.A(n_347),
.Y(n_495)
);

CKINVDCx5p33_ASAP7_75t_R g496 ( 
.A(n_313),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_283),
.Y(n_497)
);

CKINVDCx5p33_ASAP7_75t_R g498 ( 
.A(n_318),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_285),
.Y(n_499)
);

CKINVDCx5p33_ASAP7_75t_R g500 ( 
.A(n_319),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_288),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_304),
.Y(n_502)
);

BUFx3_ASAP7_75t_L g503 ( 
.A(n_347),
.Y(n_503)
);

CKINVDCx20_ASAP7_75t_R g504 ( 
.A(n_320),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_261),
.B(n_8),
.Y(n_505)
);

CKINVDCx5p33_ASAP7_75t_R g506 ( 
.A(n_325),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_316),
.Y(n_507)
);

NOR2xp67_ASAP7_75t_L g508 ( 
.A(n_213),
.B(n_8),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_317),
.Y(n_509)
);

BUFx3_ASAP7_75t_L g510 ( 
.A(n_235),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_327),
.Y(n_511)
);

CKINVDCx5p33_ASAP7_75t_R g512 ( 
.A(n_337),
.Y(n_512)
);

INVxp33_ASAP7_75t_SL g513 ( 
.A(n_227),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_328),
.Y(n_514)
);

AOI22xp5_ASAP7_75t_L g515 ( 
.A1(n_420),
.A2(n_289),
.B1(n_379),
.B2(n_378),
.Y(n_515)
);

CKINVDCx5p33_ASAP7_75t_R g516 ( 
.A(n_504),
.Y(n_516)
);

INVxp67_ASAP7_75t_L g517 ( 
.A(n_432),
.Y(n_517)
);

AND2x4_ASAP7_75t_L g518 ( 
.A(n_492),
.B(n_271),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_SL g519 ( 
.A(n_510),
.B(n_439),
.Y(n_519)
);

INVx3_ASAP7_75t_L g520 ( 
.A(n_419),
.Y(n_520)
);

AND2x4_ASAP7_75t_L g521 ( 
.A(n_492),
.B(n_424),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_409),
.B(n_271),
.Y(n_522)
);

INVx3_ASAP7_75t_L g523 ( 
.A(n_419),
.Y(n_523)
);

CKINVDCx5p33_ASAP7_75t_R g524 ( 
.A(n_410),
.Y(n_524)
);

CKINVDCx20_ASAP7_75t_R g525 ( 
.A(n_408),
.Y(n_525)
);

BUFx6f_ASAP7_75t_L g526 ( 
.A(n_412),
.Y(n_526)
);

BUFx2_ASAP7_75t_L g527 ( 
.A(n_469),
.Y(n_527)
);

AND2x4_ASAP7_75t_L g528 ( 
.A(n_479),
.B(n_388),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_415),
.B(n_416),
.Y(n_529)
);

CKINVDCx20_ASAP7_75t_R g530 ( 
.A(n_413),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_L g531 ( 
.A(n_421),
.B(n_388),
.Y(n_531)
);

BUFx6f_ASAP7_75t_L g532 ( 
.A(n_412),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_414),
.Y(n_533)
);

CKINVDCx20_ASAP7_75t_R g534 ( 
.A(n_423),
.Y(n_534)
);

BUFx3_ASAP7_75t_L g535 ( 
.A(n_495),
.Y(n_535)
);

INVx2_ASAP7_75t_L g536 ( 
.A(n_414),
.Y(n_536)
);

CKINVDCx11_ASAP7_75t_R g537 ( 
.A(n_444),
.Y(n_537)
);

CKINVDCx20_ASAP7_75t_R g538 ( 
.A(n_447),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_SL g539 ( 
.A(n_510),
.B(n_235),
.Y(n_539)
);

CKINVDCx20_ASAP7_75t_R g540 ( 
.A(n_450),
.Y(n_540)
);

CKINVDCx5p33_ASAP7_75t_R g541 ( 
.A(n_425),
.Y(n_541)
);

AND2x6_ASAP7_75t_L g542 ( 
.A(n_443),
.B(n_221),
.Y(n_542)
);

INVx2_ASAP7_75t_L g543 ( 
.A(n_417),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_417),
.Y(n_544)
);

CKINVDCx5p33_ASAP7_75t_R g545 ( 
.A(n_435),
.Y(n_545)
);

CKINVDCx5p33_ASAP7_75t_R g546 ( 
.A(n_436),
.Y(n_546)
);

CKINVDCx16_ASAP7_75t_R g547 ( 
.A(n_481),
.Y(n_547)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_418),
.Y(n_548)
);

AND2x6_ASAP7_75t_L g549 ( 
.A(n_443),
.B(n_221),
.Y(n_549)
);

CKINVDCx11_ASAP7_75t_R g550 ( 
.A(n_452),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_418),
.Y(n_551)
);

NOR2xp33_ASAP7_75t_L g552 ( 
.A(n_442),
.B(n_210),
.Y(n_552)
);

BUFx2_ASAP7_75t_L g553 ( 
.A(n_455),
.Y(n_553)
);

BUFx3_ASAP7_75t_L g554 ( 
.A(n_495),
.Y(n_554)
);

OA21x2_ASAP7_75t_L g555 ( 
.A1(n_422),
.A2(n_257),
.B(n_241),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_422),
.Y(n_556)
);

INVx2_ASAP7_75t_L g557 ( 
.A(n_426),
.Y(n_557)
);

INVx2_ASAP7_75t_L g558 ( 
.A(n_427),
.Y(n_558)
);

CKINVDCx5p33_ASAP7_75t_R g559 ( 
.A(n_446),
.Y(n_559)
);

INVx3_ASAP7_75t_L g560 ( 
.A(n_427),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_428),
.Y(n_561)
);

CKINVDCx20_ASAP7_75t_R g562 ( 
.A(n_457),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_428),
.Y(n_563)
);

BUFx8_ASAP7_75t_L g564 ( 
.A(n_440),
.Y(n_564)
);

CKINVDCx5p33_ASAP7_75t_R g565 ( 
.A(n_453),
.Y(n_565)
);

AND2x6_ASAP7_75t_L g566 ( 
.A(n_448),
.B(n_221),
.Y(n_566)
);

BUFx6f_ASAP7_75t_L g567 ( 
.A(n_429),
.Y(n_567)
);

AND2x6_ASAP7_75t_L g568 ( 
.A(n_448),
.B(n_221),
.Y(n_568)
);

INVx5_ASAP7_75t_L g569 ( 
.A(n_456),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_430),
.Y(n_570)
);

BUFx6f_ASAP7_75t_L g571 ( 
.A(n_430),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_433),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_433),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_434),
.Y(n_574)
);

BUFx6f_ASAP7_75t_L g575 ( 
.A(n_434),
.Y(n_575)
);

CKINVDCx20_ASAP7_75t_R g576 ( 
.A(n_458),
.Y(n_576)
);

INVx3_ASAP7_75t_L g577 ( 
.A(n_437),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_437),
.Y(n_578)
);

CKINVDCx5p33_ASAP7_75t_R g579 ( 
.A(n_454),
.Y(n_579)
);

HB1xp67_ASAP7_75t_L g580 ( 
.A(n_459),
.Y(n_580)
);

CKINVDCx5p33_ASAP7_75t_R g581 ( 
.A(n_463),
.Y(n_581)
);

CKINVDCx20_ASAP7_75t_R g582 ( 
.A(n_464),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_438),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_438),
.Y(n_584)
);

CKINVDCx5p33_ASAP7_75t_R g585 ( 
.A(n_465),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_488),
.Y(n_586)
);

CKINVDCx5p33_ASAP7_75t_R g587 ( 
.A(n_468),
.Y(n_587)
);

INVx3_ASAP7_75t_L g588 ( 
.A(n_456),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_466),
.Y(n_589)
);

INVx2_ASAP7_75t_L g590 ( 
.A(n_441),
.Y(n_590)
);

CKINVDCx5p33_ASAP7_75t_R g591 ( 
.A(n_470),
.Y(n_591)
);

NOR2xp33_ASAP7_75t_R g592 ( 
.A(n_472),
.B(n_351),
.Y(n_592)
);

BUFx6f_ASAP7_75t_L g593 ( 
.A(n_441),
.Y(n_593)
);

NOR2xp67_ASAP7_75t_L g594 ( 
.A(n_477),
.B(n_209),
.Y(n_594)
);

AND2x4_ASAP7_75t_L g595 ( 
.A(n_508),
.B(n_241),
.Y(n_595)
);

INVx3_ASAP7_75t_L g596 ( 
.A(n_588),
.Y(n_596)
);

BUFx3_ASAP7_75t_L g597 ( 
.A(n_535),
.Y(n_597)
);

OR2x2_ASAP7_75t_L g598 ( 
.A(n_553),
.B(n_475),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_SL g599 ( 
.A(n_521),
.B(n_257),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_L g600 ( 
.A(n_521),
.B(n_480),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_L g601 ( 
.A(n_521),
.B(n_486),
.Y(n_601)
);

INVxp67_ASAP7_75t_SL g602 ( 
.A(n_588),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_589),
.Y(n_603)
);

AND2x4_ASAP7_75t_L g604 ( 
.A(n_535),
.B(n_503),
.Y(n_604)
);

INVx5_ASAP7_75t_L g605 ( 
.A(n_542),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_586),
.Y(n_606)
);

INVx2_ASAP7_75t_L g607 ( 
.A(n_526),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_533),
.Y(n_608)
);

INVx5_ASAP7_75t_L g609 ( 
.A(n_542),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_544),
.Y(n_610)
);

OAI22xp33_ASAP7_75t_L g611 ( 
.A1(n_515),
.A2(n_251),
.B1(n_353),
.B2(n_290),
.Y(n_611)
);

NOR2xp33_ASAP7_75t_L g612 ( 
.A(n_522),
.B(n_445),
.Y(n_612)
);

NOR2xp33_ASAP7_75t_L g613 ( 
.A(n_531),
.B(n_513),
.Y(n_613)
);

BUFx3_ASAP7_75t_L g614 ( 
.A(n_554),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_551),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_SL g616 ( 
.A(n_528),
.B(n_280),
.Y(n_616)
);

INVx2_ASAP7_75t_SL g617 ( 
.A(n_554),
.Y(n_617)
);

AOI22xp33_ASAP7_75t_L g618 ( 
.A1(n_518),
.A2(n_490),
.B1(n_505),
.B2(n_411),
.Y(n_618)
);

INVx1_ASAP7_75t_SL g619 ( 
.A(n_525),
.Y(n_619)
);

AND2x6_ASAP7_75t_L g620 ( 
.A(n_518),
.B(n_280),
.Y(n_620)
);

NOR2xp33_ASAP7_75t_L g621 ( 
.A(n_552),
.B(n_487),
.Y(n_621)
);

CKINVDCx6p67_ASAP7_75t_R g622 ( 
.A(n_547),
.Y(n_622)
);

AOI22xp33_ASAP7_75t_L g623 ( 
.A1(n_518),
.A2(n_353),
.B1(n_362),
.B2(n_311),
.Y(n_623)
);

NAND2xp33_ASAP7_75t_L g624 ( 
.A(n_592),
.B(n_489),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_SL g625 ( 
.A(n_528),
.B(n_311),
.Y(n_625)
);

BUFx10_ASAP7_75t_L g626 ( 
.A(n_524),
.Y(n_626)
);

INVx1_ASAP7_75t_SL g627 ( 
.A(n_525),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_556),
.Y(n_628)
);

BUFx3_ASAP7_75t_L g629 ( 
.A(n_526),
.Y(n_629)
);

BUFx3_ASAP7_75t_L g630 ( 
.A(n_526),
.Y(n_630)
);

AOI22xp5_ASAP7_75t_L g631 ( 
.A1(n_519),
.A2(n_498),
.B1(n_500),
.B2(n_496),
.Y(n_631)
);

INVx3_ASAP7_75t_L g632 ( 
.A(n_588),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_561),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_SL g634 ( 
.A(n_528),
.B(n_221),
.Y(n_634)
);

BUFx3_ASAP7_75t_L g635 ( 
.A(n_595),
.Y(n_635)
);

INVx2_ASAP7_75t_L g636 ( 
.A(n_526),
.Y(n_636)
);

INVx4_ASAP7_75t_L g637 ( 
.A(n_532),
.Y(n_637)
);

INVxp67_ASAP7_75t_SL g638 ( 
.A(n_555),
.Y(n_638)
);

INVx5_ASAP7_75t_L g639 ( 
.A(n_542),
.Y(n_639)
);

INVx8_ASAP7_75t_L g640 ( 
.A(n_524),
.Y(n_640)
);

CKINVDCx20_ASAP7_75t_R g641 ( 
.A(n_530),
.Y(n_641)
);

NAND2xp33_ASAP7_75t_SL g642 ( 
.A(n_595),
.B(n_362),
.Y(n_642)
);

NOR2xp33_ASAP7_75t_L g643 ( 
.A(n_529),
.B(n_506),
.Y(n_643)
);

BUFx3_ASAP7_75t_L g644 ( 
.A(n_532),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_570),
.Y(n_645)
);

INVx4_ASAP7_75t_L g646 ( 
.A(n_532),
.Y(n_646)
);

INVx5_ASAP7_75t_L g647 ( 
.A(n_542),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_SL g648 ( 
.A(n_595),
.B(n_245),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_SL g649 ( 
.A(n_594),
.B(n_245),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_572),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_573),
.Y(n_651)
);

AND2x4_ASAP7_75t_L g652 ( 
.A(n_539),
.B(n_503),
.Y(n_652)
);

INVx3_ASAP7_75t_L g653 ( 
.A(n_532),
.Y(n_653)
);

NOR2x1p5_ASAP7_75t_L g654 ( 
.A(n_541),
.B(n_228),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_578),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_584),
.Y(n_656)
);

BUFx10_ASAP7_75t_L g657 ( 
.A(n_541),
.Y(n_657)
);

AO22x2_ASAP7_75t_L g658 ( 
.A1(n_517),
.A2(n_341),
.B1(n_467),
.B2(n_348),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_560),
.Y(n_659)
);

OAI22xp33_ASAP7_75t_L g660 ( 
.A1(n_545),
.A2(n_251),
.B1(n_399),
.B2(n_322),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_L g661 ( 
.A(n_560),
.B(n_512),
.Y(n_661)
);

AOI22xp33_ASAP7_75t_L g662 ( 
.A1(n_555),
.A2(n_343),
.B1(n_344),
.B2(n_334),
.Y(n_662)
);

INVx2_ASAP7_75t_L g663 ( 
.A(n_532),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_577),
.B(n_431),
.Y(n_664)
);

INVx2_ASAP7_75t_L g665 ( 
.A(n_567),
.Y(n_665)
);

BUFx2_ASAP7_75t_L g666 ( 
.A(n_530),
.Y(n_666)
);

INVx2_ASAP7_75t_L g667 ( 
.A(n_567),
.Y(n_667)
);

BUFx3_ASAP7_75t_L g668 ( 
.A(n_527),
.Y(n_668)
);

NAND2xp33_ASAP7_75t_R g669 ( 
.A(n_545),
.B(n_475),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_SL g670 ( 
.A(n_546),
.B(n_245),
.Y(n_670)
);

OR2x2_ASAP7_75t_L g671 ( 
.A(n_580),
.B(n_460),
.Y(n_671)
);

INVx4_ASAP7_75t_L g672 ( 
.A(n_567),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_SL g673 ( 
.A(n_546),
.B(n_245),
.Y(n_673)
);

NOR2xp33_ASAP7_75t_L g674 ( 
.A(n_559),
.B(n_461),
.Y(n_674)
);

OR2x6_ASAP7_75t_L g675 ( 
.A(n_564),
.B(n_482),
.Y(n_675)
);

INVx3_ASAP7_75t_L g676 ( 
.A(n_567),
.Y(n_676)
);

INVx1_ASAP7_75t_SL g677 ( 
.A(n_534),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_577),
.Y(n_678)
);

AOI22xp33_ASAP7_75t_L g679 ( 
.A1(n_555),
.A2(n_359),
.B1(n_369),
.B2(n_372),
.Y(n_679)
);

INVx4_ASAP7_75t_SL g680 ( 
.A(n_542),
.Y(n_680)
);

AO22x2_ASAP7_75t_L g681 ( 
.A1(n_536),
.A2(n_349),
.B1(n_383),
.B2(n_390),
.Y(n_681)
);

AO22x2_ASAP7_75t_L g682 ( 
.A1(n_536),
.A2(n_291),
.B1(n_222),
.B2(n_231),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_567),
.Y(n_683)
);

INVx1_ASAP7_75t_SL g684 ( 
.A(n_534),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_L g685 ( 
.A(n_571),
.B(n_485),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_L g686 ( 
.A(n_571),
.B(n_249),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_571),
.B(n_282),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_571),
.Y(n_688)
);

INVx1_ASAP7_75t_SL g689 ( 
.A(n_538),
.Y(n_689)
);

CKINVDCx20_ASAP7_75t_R g690 ( 
.A(n_538),
.Y(n_690)
);

INVx6_ASAP7_75t_L g691 ( 
.A(n_564),
.Y(n_691)
);

AOI22xp5_ASAP7_75t_L g692 ( 
.A1(n_559),
.A2(n_440),
.B1(n_244),
.B2(n_315),
.Y(n_692)
);

BUFx6f_ASAP7_75t_L g693 ( 
.A(n_571),
.Y(n_693)
);

OR2x2_ASAP7_75t_L g694 ( 
.A(n_565),
.B(n_471),
.Y(n_694)
);

INVx4_ASAP7_75t_SL g695 ( 
.A(n_542),
.Y(n_695)
);

OAI22xp33_ASAP7_75t_L g696 ( 
.A1(n_565),
.A2(n_228),
.B1(n_229),
.B2(n_238),
.Y(n_696)
);

INVx2_ASAP7_75t_L g697 ( 
.A(n_575),
.Y(n_697)
);

AND2x4_ASAP7_75t_L g698 ( 
.A(n_590),
.B(n_473),
.Y(n_698)
);

BUFx2_ASAP7_75t_L g699 ( 
.A(n_540),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_575),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_SL g701 ( 
.A(n_579),
.B(n_245),
.Y(n_701)
);

NOR2xp33_ASAP7_75t_L g702 ( 
.A(n_579),
.B(n_440),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_575),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_575),
.Y(n_704)
);

BUFx10_ASAP7_75t_L g705 ( 
.A(n_581),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_L g706 ( 
.A(n_575),
.B(n_357),
.Y(n_706)
);

OR2x2_ASAP7_75t_L g707 ( 
.A(n_581),
.B(n_473),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_543),
.Y(n_708)
);

INVx4_ASAP7_75t_L g709 ( 
.A(n_549),
.Y(n_709)
);

AND2x6_ASAP7_75t_L g710 ( 
.A(n_543),
.B(n_262),
.Y(n_710)
);

INVx2_ASAP7_75t_L g711 ( 
.A(n_520),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_L g712 ( 
.A(n_548),
.B(n_557),
.Y(n_712)
);

AND2x2_ASAP7_75t_SL g713 ( 
.A(n_590),
.B(n_262),
.Y(n_713)
);

INVx2_ASAP7_75t_L g714 ( 
.A(n_520),
.Y(n_714)
);

CKINVDCx20_ASAP7_75t_R g715 ( 
.A(n_540),
.Y(n_715)
);

INVx1_ASAP7_75t_SL g716 ( 
.A(n_562),
.Y(n_716)
);

INVx2_ASAP7_75t_L g717 ( 
.A(n_520),
.Y(n_717)
);

AOI22xp33_ASAP7_75t_L g718 ( 
.A1(n_549),
.A2(n_494),
.B1(n_511),
.B2(n_509),
.Y(n_718)
);

INVx2_ASAP7_75t_L g719 ( 
.A(n_523),
.Y(n_719)
);

BUFx6f_ASAP7_75t_L g720 ( 
.A(n_593),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_557),
.Y(n_721)
);

INVxp67_ASAP7_75t_L g722 ( 
.A(n_593),
.Y(n_722)
);

INVx4_ASAP7_75t_SL g723 ( 
.A(n_549),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_L g724 ( 
.A(n_558),
.B(n_563),
.Y(n_724)
);

INVx2_ASAP7_75t_L g725 ( 
.A(n_523),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_SL g726 ( 
.A(n_585),
.B(n_262),
.Y(n_726)
);

OR2x6_ASAP7_75t_L g727 ( 
.A(n_564),
.B(n_474),
.Y(n_727)
);

BUFx6f_ASAP7_75t_L g728 ( 
.A(n_593),
.Y(n_728)
);

NOR2x1p5_ASAP7_75t_L g729 ( 
.A(n_585),
.B(n_229),
.Y(n_729)
);

CKINVDCx5p33_ASAP7_75t_R g730 ( 
.A(n_587),
.Y(n_730)
);

INVx2_ASAP7_75t_L g731 ( 
.A(n_523),
.Y(n_731)
);

AO21x2_ASAP7_75t_L g732 ( 
.A1(n_563),
.A2(n_242),
.B(n_236),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_SL g733 ( 
.A(n_587),
.B(n_262),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_L g734 ( 
.A(n_574),
.B(n_583),
.Y(n_734)
);

INVx3_ASAP7_75t_L g735 ( 
.A(n_593),
.Y(n_735)
);

AND2x4_ASAP7_75t_L g736 ( 
.A(n_574),
.B(n_474),
.Y(n_736)
);

OAI22xp5_ASAP7_75t_L g737 ( 
.A1(n_591),
.A2(n_314),
.B1(n_338),
.B2(n_335),
.Y(n_737)
);

BUFx6f_ASAP7_75t_L g738 ( 
.A(n_635),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_643),
.B(n_591),
.Y(n_739)
);

BUFx6f_ASAP7_75t_L g740 ( 
.A(n_614),
.Y(n_740)
);

BUFx3_ASAP7_75t_L g741 ( 
.A(n_597),
.Y(n_741)
);

NOR2xp33_ASAP7_75t_L g742 ( 
.A(n_621),
.B(n_386),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_L g743 ( 
.A(n_643),
.B(n_583),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_L g744 ( 
.A(n_621),
.B(n_549),
.Y(n_744)
);

INVx2_ASAP7_75t_SL g745 ( 
.A(n_604),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_L g746 ( 
.A(n_602),
.B(n_549),
.Y(n_746)
);

AND2x2_ASAP7_75t_L g747 ( 
.A(n_674),
.B(n_516),
.Y(n_747)
);

OAI22xp33_ASAP7_75t_L g748 ( 
.A1(n_611),
.A2(n_392),
.B1(n_385),
.B2(n_382),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_602),
.B(n_549),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_L g750 ( 
.A(n_664),
.B(n_566),
.Y(n_750)
);

AND2x4_ASAP7_75t_L g751 ( 
.A(n_614),
.B(n_617),
.Y(n_751)
);

NOR2xp33_ASAP7_75t_L g752 ( 
.A(n_612),
.B(n_206),
.Y(n_752)
);

INVx2_ASAP7_75t_SL g753 ( 
.A(n_604),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_L g754 ( 
.A(n_638),
.B(n_685),
.Y(n_754)
);

A2O1A1Ixp33_ASAP7_75t_L g755 ( 
.A1(n_618),
.A2(n_391),
.B(n_256),
.C(n_267),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_606),
.Y(n_756)
);

AOI22xp5_ASAP7_75t_L g757 ( 
.A1(n_612),
.A2(n_356),
.B1(n_374),
.B2(n_361),
.Y(n_757)
);

OR2x6_ASAP7_75t_L g758 ( 
.A(n_640),
.B(n_476),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_638),
.B(n_566),
.Y(n_759)
);

INVx2_ASAP7_75t_L g760 ( 
.A(n_596),
.Y(n_760)
);

INVx4_ASAP7_75t_L g761 ( 
.A(n_720),
.Y(n_761)
);

NOR3xp33_ASAP7_75t_L g762 ( 
.A(n_611),
.B(n_550),
.C(n_537),
.Y(n_762)
);

NOR2x1p5_ASAP7_75t_L g763 ( 
.A(n_622),
.B(n_516),
.Y(n_763)
);

NOR2xp33_ASAP7_75t_L g764 ( 
.A(n_613),
.B(n_707),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_603),
.Y(n_765)
);

AOI22xp33_ASAP7_75t_L g766 ( 
.A1(n_662),
.A2(n_262),
.B1(n_300),
.B2(n_384),
.Y(n_766)
);

INVx2_ASAP7_75t_L g767 ( 
.A(n_632),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_L g768 ( 
.A(n_613),
.B(n_566),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_L g769 ( 
.A(n_713),
.B(n_566),
.Y(n_769)
);

AND2x2_ASAP7_75t_L g770 ( 
.A(n_674),
.B(n_278),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_713),
.B(n_566),
.Y(n_771)
);

NOR2x2_ASAP7_75t_L g772 ( 
.A(n_727),
.B(n_562),
.Y(n_772)
);

NOR3xp33_ASAP7_75t_L g773 ( 
.A(n_660),
.B(n_478),
.C(n_476),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_L g774 ( 
.A(n_599),
.B(n_566),
.Y(n_774)
);

INVx2_ASAP7_75t_L g775 ( 
.A(n_632),
.Y(n_775)
);

AOI22xp5_ASAP7_75t_L g776 ( 
.A1(n_600),
.A2(n_601),
.B1(n_599),
.B2(n_618),
.Y(n_776)
);

AND2x2_ASAP7_75t_L g777 ( 
.A(n_694),
.B(n_310),
.Y(n_777)
);

INVx2_ASAP7_75t_L g778 ( 
.A(n_711),
.Y(n_778)
);

OAI221xp5_ASAP7_75t_L g779 ( 
.A1(n_623),
.A2(n_342),
.B1(n_340),
.B2(n_367),
.C(n_250),
.Y(n_779)
);

AOI22xp33_ASAP7_75t_L g780 ( 
.A1(n_679),
.A2(n_336),
.B1(n_332),
.B2(n_331),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_661),
.B(n_568),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_698),
.Y(n_782)
);

NOR2xp33_ASAP7_75t_L g783 ( 
.A(n_671),
.B(n_206),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_SL g784 ( 
.A(n_605),
.B(n_263),
.Y(n_784)
);

INVxp67_ASAP7_75t_L g785 ( 
.A(n_598),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_L g786 ( 
.A(n_608),
.B(n_568),
.Y(n_786)
);

OR2x6_ASAP7_75t_L g787 ( 
.A(n_640),
.B(n_691),
.Y(n_787)
);

AND2x2_ASAP7_75t_L g788 ( 
.A(n_652),
.B(n_310),
.Y(n_788)
);

INVx2_ASAP7_75t_L g789 ( 
.A(n_714),
.Y(n_789)
);

AOI22xp5_ASAP7_75t_L g790 ( 
.A1(n_620),
.A2(n_360),
.B1(n_358),
.B2(n_354),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_SL g791 ( 
.A(n_605),
.B(n_263),
.Y(n_791)
);

OAI221xp5_ASAP7_75t_L g792 ( 
.A1(n_623),
.A2(n_270),
.B1(n_312),
.B2(n_397),
.C(n_396),
.Y(n_792)
);

INVx2_ASAP7_75t_SL g793 ( 
.A(n_652),
.Y(n_793)
);

AOI22xp33_ASAP7_75t_L g794 ( 
.A1(n_679),
.A2(n_398),
.B1(n_293),
.B2(n_272),
.Y(n_794)
);

INVx2_ASAP7_75t_L g795 ( 
.A(n_717),
.Y(n_795)
);

AOI21xp5_ASAP7_75t_L g796 ( 
.A1(n_686),
.A2(n_569),
.B(n_287),
.Y(n_796)
);

NOR2xp67_ASAP7_75t_L g797 ( 
.A(n_702),
.B(n_631),
.Y(n_797)
);

OAI22xp33_ASAP7_75t_L g798 ( 
.A1(n_660),
.A2(n_382),
.B1(n_385),
.B2(n_392),
.Y(n_798)
);

BUFx2_ASAP7_75t_L g799 ( 
.A(n_641),
.Y(n_799)
);

AOI22xp33_ASAP7_75t_L g800 ( 
.A1(n_620),
.A2(n_269),
.B1(n_381),
.B2(n_263),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_L g801 ( 
.A(n_610),
.B(n_568),
.Y(n_801)
);

NOR2xp33_ASAP7_75t_L g802 ( 
.A(n_670),
.B(n_218),
.Y(n_802)
);

NOR2xp33_ASAP7_75t_L g803 ( 
.A(n_670),
.B(n_218),
.Y(n_803)
);

AOI21xp5_ASAP7_75t_L g804 ( 
.A1(n_687),
.A2(n_706),
.B(n_722),
.Y(n_804)
);

INVx2_ASAP7_75t_L g805 ( 
.A(n_719),
.Y(n_805)
);

INVx1_ASAP7_75t_SL g806 ( 
.A(n_690),
.Y(n_806)
);

NOR2xp33_ASAP7_75t_L g807 ( 
.A(n_673),
.B(n_220),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_L g808 ( 
.A(n_615),
.B(n_568),
.Y(n_808)
);

NOR2xp33_ASAP7_75t_L g809 ( 
.A(n_673),
.B(n_220),
.Y(n_809)
);

AOI22xp5_ASAP7_75t_L g810 ( 
.A1(n_620),
.A2(n_352),
.B1(n_380),
.B2(n_377),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_698),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_SL g812 ( 
.A(n_605),
.B(n_263),
.Y(n_812)
);

NOR2xp33_ASAP7_75t_L g813 ( 
.A(n_701),
.B(n_224),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_SL g814 ( 
.A(n_605),
.B(n_224),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_L g815 ( 
.A(n_628),
.B(n_568),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_736),
.Y(n_816)
);

INVx2_ASAP7_75t_L g817 ( 
.A(n_725),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_SL g818 ( 
.A(n_609),
.B(n_226),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_L g819 ( 
.A(n_633),
.B(n_568),
.Y(n_819)
);

AOI21xp5_ASAP7_75t_L g820 ( 
.A1(n_722),
.A2(n_569),
.B(n_483),
.Y(n_820)
);

INVx2_ASAP7_75t_L g821 ( 
.A(n_731),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_SL g822 ( 
.A(n_701),
.B(n_226),
.Y(n_822)
);

INVx8_ASAP7_75t_L g823 ( 
.A(n_640),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_SL g824 ( 
.A(n_609),
.B(n_233),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_736),
.Y(n_825)
);

HB1xp67_ASAP7_75t_L g826 ( 
.A(n_681),
.Y(n_826)
);

NAND2xp33_ASAP7_75t_SL g827 ( 
.A(n_654),
.B(n_238),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_L g828 ( 
.A(n_645),
.B(n_569),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_L g829 ( 
.A(n_650),
.B(n_569),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_L g830 ( 
.A(n_651),
.B(n_233),
.Y(n_830)
);

INVx2_ASAP7_75t_L g831 ( 
.A(n_708),
.Y(n_831)
);

AOI22xp5_ASAP7_75t_L g832 ( 
.A1(n_620),
.A2(n_240),
.B1(n_244),
.B2(n_315),
.Y(n_832)
);

NOR3xp33_ASAP7_75t_L g833 ( 
.A(n_737),
.B(n_478),
.C(n_514),
.Y(n_833)
);

INVx4_ASAP7_75t_L g834 ( 
.A(n_720),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_SL g835 ( 
.A(n_609),
.B(n_239),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_SL g836 ( 
.A(n_726),
.B(n_239),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_L g837 ( 
.A(n_655),
.B(n_240),
.Y(n_837)
);

AO221x1_ASAP7_75t_L g838 ( 
.A1(n_696),
.A2(n_514),
.B1(n_483),
.B2(n_484),
.C(n_491),
.Y(n_838)
);

BUFx6f_ASAP7_75t_L g839 ( 
.A(n_620),
.Y(n_839)
);

AOI22xp5_ASAP7_75t_L g840 ( 
.A1(n_726),
.A2(n_395),
.B1(n_405),
.B2(n_394),
.Y(n_840)
);

NAND2xp33_ASAP7_75t_L g841 ( 
.A(n_718),
.B(n_387),
.Y(n_841)
);

AND2x2_ASAP7_75t_L g842 ( 
.A(n_626),
.B(n_323),
.Y(n_842)
);

AOI21xp5_ASAP7_75t_L g843 ( 
.A1(n_712),
.A2(n_491),
.B(n_509),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_656),
.Y(n_844)
);

INVx3_ASAP7_75t_L g845 ( 
.A(n_629),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_L g846 ( 
.A(n_659),
.B(n_387),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_678),
.Y(n_847)
);

OR2x2_ASAP7_75t_L g848 ( 
.A(n_619),
.B(n_484),
.Y(n_848)
);

NOR2xp33_ASAP7_75t_SL g849 ( 
.A(n_730),
.B(n_576),
.Y(n_849)
);

AOI221xp5_ASAP7_75t_L g850 ( 
.A1(n_696),
.A2(n_400),
.B1(n_401),
.B2(n_402),
.C(n_403),
.Y(n_850)
);

AOI22xp5_ASAP7_75t_L g851 ( 
.A1(n_733),
.A2(n_405),
.B1(n_395),
.B2(n_394),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_721),
.Y(n_852)
);

CKINVDCx5p33_ASAP7_75t_R g853 ( 
.A(n_626),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_735),
.B(n_389),
.Y(n_854)
);

OR2x2_ASAP7_75t_L g855 ( 
.A(n_627),
.B(n_493),
.Y(n_855)
);

NOR2xp33_ASAP7_75t_L g856 ( 
.A(n_733),
.B(n_389),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_735),
.B(n_494),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_L g858 ( 
.A(n_653),
.B(n_497),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_L g859 ( 
.A(n_653),
.B(n_497),
.Y(n_859)
);

AOI22xp33_ASAP7_75t_L g860 ( 
.A1(n_681),
.A2(n_406),
.B1(n_400),
.B2(n_403),
.Y(n_860)
);

AOI22xp33_ASAP7_75t_L g861 ( 
.A1(n_681),
.A2(n_406),
.B1(n_401),
.B2(n_402),
.Y(n_861)
);

NOR2xp33_ASAP7_75t_L g862 ( 
.A(n_692),
.B(n_208),
.Y(n_862)
);

CKINVDCx5p33_ASAP7_75t_R g863 ( 
.A(n_657),
.Y(n_863)
);

AOI22xp5_ASAP7_75t_L g864 ( 
.A1(n_624),
.A2(n_364),
.B1(n_292),
.B2(n_345),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_676),
.B(n_499),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_L g866 ( 
.A(n_676),
.B(n_499),
.Y(n_866)
);

AOI22xp33_ASAP7_75t_L g867 ( 
.A1(n_682),
.A2(n_323),
.B1(n_501),
.B2(n_507),
.Y(n_867)
);

NOR2xp33_ASAP7_75t_L g868 ( 
.A(n_702),
.B(n_212),
.Y(n_868)
);

AND2x2_ASAP7_75t_L g869 ( 
.A(n_657),
.B(n_705),
.Y(n_869)
);

INVx3_ASAP7_75t_L g870 ( 
.A(n_629),
.Y(n_870)
);

AND2x2_ASAP7_75t_L g871 ( 
.A(n_705),
.B(n_323),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_630),
.B(n_501),
.Y(n_872)
);

OAI22xp5_ASAP7_75t_SL g873 ( 
.A1(n_715),
.A2(n_582),
.B1(n_576),
.B2(n_253),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_SL g874 ( 
.A(n_609),
.B(n_292),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_SL g875 ( 
.A(n_639),
.B(n_647),
.Y(n_875)
);

NOR2xp33_ASAP7_75t_L g876 ( 
.A(n_616),
.B(n_258),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_SL g877 ( 
.A(n_639),
.B(n_292),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_630),
.B(n_502),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_SL g879 ( 
.A(n_642),
.B(n_345),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_L g880 ( 
.A(n_644),
.B(n_502),
.Y(n_880)
);

AND2x4_ASAP7_75t_L g881 ( 
.A(n_616),
.B(n_507),
.Y(n_881)
);

INVx3_ASAP7_75t_L g882 ( 
.A(n_644),
.Y(n_882)
);

O2A1O1Ixp33_ASAP7_75t_L g883 ( 
.A1(n_625),
.A2(n_462),
.B(n_451),
.C(n_449),
.Y(n_883)
);

AND2x2_ASAP7_75t_SL g884 ( 
.A(n_718),
.B(n_449),
.Y(n_884)
);

INVx2_ASAP7_75t_L g885 ( 
.A(n_724),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_L g886 ( 
.A(n_634),
.B(n_279),
.Y(n_886)
);

AND2x6_ASAP7_75t_SL g887 ( 
.A(n_675),
.B(n_451),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_734),
.Y(n_888)
);

AND2x6_ASAP7_75t_SL g889 ( 
.A(n_675),
.B(n_727),
.Y(n_889)
);

AND2x6_ASAP7_75t_SL g890 ( 
.A(n_675),
.B(n_462),
.Y(n_890)
);

NOR2xp33_ASAP7_75t_L g891 ( 
.A(n_625),
.B(n_281),
.Y(n_891)
);

O2A1O1Ixp5_ASAP7_75t_L g892 ( 
.A1(n_648),
.A2(n_364),
.B(n_345),
.C(n_375),
.Y(n_892)
);

NOR2xp33_ASAP7_75t_L g893 ( 
.A(n_642),
.B(n_286),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_SL g894 ( 
.A(n_639),
.B(n_364),
.Y(n_894)
);

NOR3xp33_ASAP7_75t_L g895 ( 
.A(n_677),
.B(n_363),
.C(n_376),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_L g896 ( 
.A(n_634),
.B(n_301),
.Y(n_896)
);

OR2x6_ASAP7_75t_L g897 ( 
.A(n_691),
.B(n_582),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_L g898 ( 
.A(n_683),
.B(n_321),
.Y(n_898)
);

NOR2xp33_ASAP7_75t_L g899 ( 
.A(n_742),
.B(n_684),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_L g900 ( 
.A(n_888),
.B(n_732),
.Y(n_900)
);

O2A1O1Ixp33_ASAP7_75t_L g901 ( 
.A1(n_755),
.A2(n_648),
.B(n_649),
.C(n_732),
.Y(n_901)
);

AOI21xp5_ASAP7_75t_L g902 ( 
.A1(n_754),
.A2(n_709),
.B(n_637),
.Y(n_902)
);

AOI21xp5_ASAP7_75t_L g903 ( 
.A1(n_804),
.A2(n_709),
.B(n_637),
.Y(n_903)
);

BUFx2_ASAP7_75t_L g904 ( 
.A(n_799),
.Y(n_904)
);

AOI21xp5_ASAP7_75t_L g905 ( 
.A1(n_759),
.A2(n_646),
.B(n_672),
.Y(n_905)
);

INVx3_ASAP7_75t_L g906 ( 
.A(n_845),
.Y(n_906)
);

AOI21xp5_ASAP7_75t_L g907 ( 
.A1(n_743),
.A2(n_781),
.B(n_750),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_L g908 ( 
.A(n_742),
.B(n_688),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_885),
.B(n_700),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_782),
.Y(n_910)
);

BUFx6f_ASAP7_75t_L g911 ( 
.A(n_740),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_776),
.B(n_703),
.Y(n_912)
);

BUFx2_ASAP7_75t_L g913 ( 
.A(n_785),
.Y(n_913)
);

A2O1A1Ixp33_ASAP7_75t_L g914 ( 
.A1(n_752),
.A2(n_729),
.B(n_649),
.C(n_704),
.Y(n_914)
);

AOI21x1_ASAP7_75t_L g915 ( 
.A1(n_744),
.A2(n_749),
.B(n_746),
.Y(n_915)
);

AOI21xp5_ASAP7_75t_L g916 ( 
.A1(n_870),
.A2(n_639),
.B(n_647),
.Y(n_916)
);

AOI21xp5_ASAP7_75t_L g917 ( 
.A1(n_870),
.A2(n_647),
.B(n_728),
.Y(n_917)
);

A2O1A1Ixp33_ASAP7_75t_L g918 ( 
.A1(n_752),
.A2(n_663),
.B(n_665),
.C(n_636),
.Y(n_918)
);

OAI21xp5_ASAP7_75t_L g919 ( 
.A1(n_766),
.A2(n_667),
.B(n_607),
.Y(n_919)
);

AOI21xp5_ASAP7_75t_L g920 ( 
.A1(n_882),
.A2(n_647),
.B(n_728),
.Y(n_920)
);

AOI21xp5_ASAP7_75t_L g921 ( 
.A1(n_882),
.A2(n_834),
.B(n_761),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_L g922 ( 
.A(n_764),
.B(n_697),
.Y(n_922)
);

AND2x6_ASAP7_75t_L g923 ( 
.A(n_839),
.B(n_668),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_L g924 ( 
.A(n_764),
.B(n_682),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_811),
.Y(n_925)
);

INVxp67_ASAP7_75t_L g926 ( 
.A(n_848),
.Y(n_926)
);

AOI21x1_ASAP7_75t_L g927 ( 
.A1(n_768),
.A2(n_682),
.B(n_693),
.Y(n_927)
);

OAI321xp33_ASAP7_75t_L g928 ( 
.A1(n_748),
.A2(n_658),
.A3(n_727),
.B1(n_669),
.B2(n_666),
.C(n_699),
.Y(n_928)
);

O2A1O1Ixp33_ASAP7_75t_L g929 ( 
.A1(n_826),
.A2(n_716),
.B(n_689),
.C(n_658),
.Y(n_929)
);

AND2x2_ASAP7_75t_L g930 ( 
.A(n_770),
.B(n_658),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_816),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_825),
.Y(n_932)
);

AND2x2_ASAP7_75t_L g933 ( 
.A(n_747),
.B(n_691),
.Y(n_933)
);

OAI21xp33_ASAP7_75t_L g934 ( 
.A1(n_783),
.A2(n_368),
.B(n_326),
.Y(n_934)
);

NAND3xp33_ASAP7_75t_L g935 ( 
.A(n_783),
.B(n_669),
.C(n_324),
.Y(n_935)
);

INVx2_ASAP7_75t_SL g936 ( 
.A(n_855),
.Y(n_936)
);

NOR2xp33_ASAP7_75t_L g937 ( 
.A(n_739),
.B(n_346),
.Y(n_937)
);

A2O1A1Ixp33_ASAP7_75t_L g938 ( 
.A1(n_802),
.A2(n_373),
.B(n_355),
.C(n_365),
.Y(n_938)
);

AOI21x1_ASAP7_75t_L g939 ( 
.A1(n_786),
.A2(n_693),
.B(n_695),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_L g940 ( 
.A(n_766),
.B(n_693),
.Y(n_940)
);

HB1xp67_ASAP7_75t_L g941 ( 
.A(n_826),
.Y(n_941)
);

BUFx6f_ASAP7_75t_L g942 ( 
.A(n_740),
.Y(n_942)
);

AOI21xp5_ASAP7_75t_L g943 ( 
.A1(n_774),
.A2(n_723),
.B(n_695),
.Y(n_943)
);

AOI21xp5_ASAP7_75t_L g944 ( 
.A1(n_875),
.A2(n_723),
.B(n_695),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_SL g945 ( 
.A(n_797),
.B(n_723),
.Y(n_945)
);

AOI21xp5_ASAP7_75t_L g946 ( 
.A1(n_875),
.A2(n_808),
.B(n_801),
.Y(n_946)
);

AOI21xp5_ASAP7_75t_L g947 ( 
.A1(n_815),
.A2(n_680),
.B(n_710),
.Y(n_947)
);

NAND3xp33_ASAP7_75t_L g948 ( 
.A(n_868),
.B(n_350),
.C(n_366),
.Y(n_948)
);

AO21x2_ASAP7_75t_L g949 ( 
.A1(n_769),
.A2(n_771),
.B(n_847),
.Y(n_949)
);

AOI21x1_ASAP7_75t_L g950 ( 
.A1(n_819),
.A2(n_710),
.B(n_125),
.Y(n_950)
);

NAND3xp33_ASAP7_75t_L g951 ( 
.A(n_868),
.B(n_862),
.C(n_850),
.Y(n_951)
);

INVxp67_ASAP7_75t_L g952 ( 
.A(n_777),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_SL g953 ( 
.A(n_738),
.B(n_370),
.Y(n_953)
);

AOI21x1_ASAP7_75t_L g954 ( 
.A1(n_828),
.A2(n_710),
.B(n_205),
.Y(n_954)
);

BUFx6f_ASAP7_75t_L g955 ( 
.A(n_740),
.Y(n_955)
);

AOI21xp5_ASAP7_75t_L g956 ( 
.A1(n_829),
.A2(n_710),
.B(n_200),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_765),
.Y(n_957)
);

NAND2xp33_ASAP7_75t_L g958 ( 
.A(n_839),
.B(n_780),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_L g959 ( 
.A(n_780),
.B(n_11),
.Y(n_959)
);

BUFx3_ASAP7_75t_L g960 ( 
.A(n_741),
.Y(n_960)
);

AND2x4_ASAP7_75t_L g961 ( 
.A(n_751),
.B(n_199),
.Y(n_961)
);

A2O1A1Ixp33_ASAP7_75t_L g962 ( 
.A1(n_802),
.A2(n_18),
.B(n_21),
.C(n_22),
.Y(n_962)
);

AOI21xp5_ASAP7_75t_L g963 ( 
.A1(n_760),
.A2(n_181),
.B(n_179),
.Y(n_963)
);

AOI21x1_ASAP7_75t_L g964 ( 
.A1(n_796),
.A2(n_171),
.B(n_162),
.Y(n_964)
);

CKINVDCx5p33_ASAP7_75t_R g965 ( 
.A(n_853),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_L g966 ( 
.A(n_794),
.B(n_112),
.Y(n_966)
);

BUFx4f_ASAP7_75t_L g967 ( 
.A(n_823),
.Y(n_967)
);

A2O1A1Ixp33_ASAP7_75t_L g968 ( 
.A1(n_803),
.A2(n_18),
.B(n_27),
.C(n_30),
.Y(n_968)
);

OAI22xp5_ASAP7_75t_L g969 ( 
.A1(n_794),
.A2(n_32),
.B1(n_33),
.B2(n_35),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_L g970 ( 
.A(n_884),
.B(n_110),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_L g971 ( 
.A(n_884),
.B(n_152),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_L g972 ( 
.A(n_881),
.B(n_104),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_L g973 ( 
.A(n_881),
.B(n_149),
.Y(n_973)
);

AND2x6_ASAP7_75t_L g974 ( 
.A(n_839),
.B(n_140),
.Y(n_974)
);

BUFx2_ASAP7_75t_L g975 ( 
.A(n_897),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_844),
.Y(n_976)
);

AOI22x1_ASAP7_75t_L g977 ( 
.A1(n_767),
.A2(n_124),
.B1(n_119),
.B2(n_118),
.Y(n_977)
);

INVxp67_ASAP7_75t_L g978 ( 
.A(n_788),
.Y(n_978)
);

AOI21xp5_ASAP7_75t_L g979 ( 
.A1(n_775),
.A2(n_115),
.B(n_99),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_SL g980 ( 
.A(n_738),
.B(n_740),
.Y(n_980)
);

OAI21xp5_ASAP7_75t_L g981 ( 
.A1(n_800),
.A2(n_98),
.B(n_97),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_L g982 ( 
.A(n_803),
.B(n_36),
.Y(n_982)
);

AOI21xp5_ASAP7_75t_L g983 ( 
.A1(n_854),
.A2(n_83),
.B(n_80),
.Y(n_983)
);

CKINVDCx5p33_ASAP7_75t_R g984 ( 
.A(n_863),
.Y(n_984)
);

AOI21xp5_ASAP7_75t_L g985 ( 
.A1(n_898),
.A2(n_76),
.B(n_37),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_L g986 ( 
.A(n_807),
.B(n_36),
.Y(n_986)
);

AOI21xp5_ASAP7_75t_L g987 ( 
.A1(n_872),
.A2(n_38),
.B(n_40),
.Y(n_987)
);

AOI21xp5_ASAP7_75t_L g988 ( 
.A1(n_878),
.A2(n_880),
.B(n_846),
.Y(n_988)
);

INVx2_ASAP7_75t_L g989 ( 
.A(n_852),
.Y(n_989)
);

OAI22xp5_ASAP7_75t_L g990 ( 
.A1(n_860),
.A2(n_40),
.B1(n_42),
.B2(n_46),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_L g991 ( 
.A(n_807),
.B(n_42),
.Y(n_991)
);

AND2x4_ASAP7_75t_L g992 ( 
.A(n_751),
.B(n_52),
.Y(n_992)
);

NOR2xp33_ASAP7_75t_SL g993 ( 
.A(n_849),
.B(n_53),
.Y(n_993)
);

OAI22xp5_ASAP7_75t_L g994 ( 
.A1(n_860),
.A2(n_53),
.B1(n_54),
.B2(n_57),
.Y(n_994)
);

BUFx12f_ASAP7_75t_L g995 ( 
.A(n_887),
.Y(n_995)
);

AOI22xp33_ASAP7_75t_L g996 ( 
.A1(n_838),
.A2(n_58),
.B1(n_59),
.B2(n_60),
.Y(n_996)
);

AO22x1_ASAP7_75t_L g997 ( 
.A1(n_862),
.A2(n_58),
.B1(n_62),
.B2(n_63),
.Y(n_997)
);

AND2x2_ASAP7_75t_L g998 ( 
.A(n_842),
.B(n_62),
.Y(n_998)
);

A2O1A1Ixp33_ASAP7_75t_L g999 ( 
.A1(n_809),
.A2(n_68),
.B(n_64),
.C(n_65),
.Y(n_999)
);

INVx4_ASAP7_75t_L g1000 ( 
.A(n_823),
.Y(n_1000)
);

NAND3xp33_ASAP7_75t_L g1001 ( 
.A(n_809),
.B(n_63),
.C(n_65),
.Y(n_1001)
);

O2A1O1Ixp33_ASAP7_75t_L g1002 ( 
.A1(n_779),
.A2(n_67),
.B(n_792),
.C(n_841),
.Y(n_1002)
);

BUFx8_ASAP7_75t_SL g1003 ( 
.A(n_897),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_L g1004 ( 
.A(n_813),
.B(n_856),
.Y(n_1004)
);

AOI21xp33_ASAP7_75t_L g1005 ( 
.A1(n_813),
.A2(n_856),
.B(n_891),
.Y(n_1005)
);

A2O1A1Ixp33_ASAP7_75t_L g1006 ( 
.A1(n_876),
.A2(n_891),
.B(n_893),
.C(n_756),
.Y(n_1006)
);

AOI21xp5_ASAP7_75t_L g1007 ( 
.A1(n_784),
.A2(n_812),
.B(n_791),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_L g1008 ( 
.A(n_876),
.B(n_857),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_858),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_L g1010 ( 
.A(n_859),
.B(n_866),
.Y(n_1010)
);

AOI21xp5_ASAP7_75t_L g1011 ( 
.A1(n_745),
.A2(n_753),
.B(n_795),
.Y(n_1011)
);

AO21x1_ASAP7_75t_L g1012 ( 
.A1(n_822),
.A2(n_836),
.B(n_893),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_L g1013 ( 
.A(n_865),
.B(n_793),
.Y(n_1013)
);

O2A1O1Ixp33_ASAP7_75t_L g1014 ( 
.A1(n_748),
.A2(n_798),
.B(n_886),
.C(n_896),
.Y(n_1014)
);

AOI21xp5_ASAP7_75t_L g1015 ( 
.A1(n_778),
.A2(n_821),
.B(n_817),
.Y(n_1015)
);

AOI22xp5_ASAP7_75t_L g1016 ( 
.A1(n_738),
.A2(n_789),
.B1(n_805),
.B2(n_832),
.Y(n_1016)
);

OA22x2_ASAP7_75t_L g1017 ( 
.A1(n_864),
.A2(n_758),
.B1(n_871),
.B2(n_873),
.Y(n_1017)
);

NOR3xp33_ASAP7_75t_L g1018 ( 
.A(n_798),
.B(n_827),
.C(n_806),
.Y(n_1018)
);

NOR2xp33_ASAP7_75t_L g1019 ( 
.A(n_757),
.B(n_837),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_L g1020 ( 
.A(n_830),
.B(n_851),
.Y(n_1020)
);

NAND2xp5_ASAP7_75t_L g1021 ( 
.A(n_840),
.B(n_833),
.Y(n_1021)
);

AOI21xp5_ASAP7_75t_L g1022 ( 
.A1(n_800),
.A2(n_835),
.B(n_818),
.Y(n_1022)
);

BUFx3_ASAP7_75t_L g1023 ( 
.A(n_823),
.Y(n_1023)
);

OAI21xp5_ASAP7_75t_L g1024 ( 
.A1(n_892),
.A2(n_810),
.B(n_790),
.Y(n_1024)
);

AOI21xp5_ASAP7_75t_L g1025 ( 
.A1(n_814),
.A2(n_835),
.B(n_824),
.Y(n_1025)
);

AND2x2_ASAP7_75t_L g1026 ( 
.A(n_758),
.B(n_861),
.Y(n_1026)
);

AOI21xp5_ASAP7_75t_L g1027 ( 
.A1(n_814),
.A2(n_824),
.B(n_818),
.Y(n_1027)
);

NOR2x1p5_ASAP7_75t_L g1028 ( 
.A(n_772),
.B(n_787),
.Y(n_1028)
);

INVx2_ASAP7_75t_L g1029 ( 
.A(n_874),
.Y(n_1029)
);

AOI21xp5_ASAP7_75t_L g1030 ( 
.A1(n_820),
.A2(n_874),
.B(n_894),
.Y(n_1030)
);

NAND2xp5_ASAP7_75t_L g1031 ( 
.A(n_867),
.B(n_843),
.Y(n_1031)
);

AOI21xp5_ASAP7_75t_L g1032 ( 
.A1(n_877),
.A2(n_894),
.B(n_879),
.Y(n_1032)
);

NAND2xp5_ASAP7_75t_L g1033 ( 
.A(n_877),
.B(n_861),
.Y(n_1033)
);

AOI21xp5_ASAP7_75t_L g1034 ( 
.A1(n_883),
.A2(n_895),
.B(n_787),
.Y(n_1034)
);

NAND2xp5_ASAP7_75t_L g1035 ( 
.A(n_773),
.B(n_787),
.Y(n_1035)
);

INVx3_ASAP7_75t_SL g1036 ( 
.A(n_763),
.Y(n_1036)
);

NAND2xp5_ASAP7_75t_L g1037 ( 
.A(n_762),
.B(n_890),
.Y(n_1037)
);

OAI321xp33_ASAP7_75t_L g1038 ( 
.A1(n_889),
.A2(n_748),
.A3(n_742),
.B1(n_611),
.B2(n_798),
.C(n_752),
.Y(n_1038)
);

INVx5_ASAP7_75t_L g1039 ( 
.A(n_839),
.Y(n_1039)
);

INVx2_ASAP7_75t_L g1040 ( 
.A(n_831),
.Y(n_1040)
);

AOI21xp5_ASAP7_75t_L g1041 ( 
.A1(n_754),
.A2(n_638),
.B(n_804),
.Y(n_1041)
);

INVx5_ASAP7_75t_L g1042 ( 
.A(n_839),
.Y(n_1042)
);

NAND3xp33_ASAP7_75t_L g1043 ( 
.A(n_742),
.B(n_752),
.C(n_764),
.Y(n_1043)
);

INVx1_ASAP7_75t_L g1044 ( 
.A(n_782),
.Y(n_1044)
);

INVx1_ASAP7_75t_SL g1045 ( 
.A(n_848),
.Y(n_1045)
);

INVx1_ASAP7_75t_L g1046 ( 
.A(n_782),
.Y(n_1046)
);

INVx1_ASAP7_75t_SL g1047 ( 
.A(n_848),
.Y(n_1047)
);

OAI21xp5_ASAP7_75t_L g1048 ( 
.A1(n_754),
.A2(n_638),
.B(n_759),
.Y(n_1048)
);

NOR2xp33_ASAP7_75t_L g1049 ( 
.A(n_742),
.B(n_764),
.Y(n_1049)
);

NAND2xp5_ASAP7_75t_L g1050 ( 
.A(n_888),
.B(n_742),
.Y(n_1050)
);

AND2x2_ASAP7_75t_L g1051 ( 
.A(n_764),
.B(n_770),
.Y(n_1051)
);

NOR2xp33_ASAP7_75t_L g1052 ( 
.A(n_742),
.B(n_764),
.Y(n_1052)
);

AOI21xp5_ASAP7_75t_L g1053 ( 
.A1(n_754),
.A2(n_638),
.B(n_804),
.Y(n_1053)
);

O2A1O1Ixp33_ASAP7_75t_L g1054 ( 
.A1(n_755),
.A2(n_742),
.B(n_826),
.C(n_752),
.Y(n_1054)
);

BUFx2_ASAP7_75t_SL g1055 ( 
.A(n_869),
.Y(n_1055)
);

AOI21xp5_ASAP7_75t_L g1056 ( 
.A1(n_754),
.A2(n_638),
.B(n_804),
.Y(n_1056)
);

O2A1O1Ixp33_ASAP7_75t_L g1057 ( 
.A1(n_755),
.A2(n_742),
.B(n_826),
.C(n_752),
.Y(n_1057)
);

AOI21xp5_ASAP7_75t_L g1058 ( 
.A1(n_754),
.A2(n_638),
.B(n_804),
.Y(n_1058)
);

NAND2xp5_ASAP7_75t_SL g1059 ( 
.A(n_742),
.B(n_739),
.Y(n_1059)
);

A2O1A1Ixp33_ASAP7_75t_L g1060 ( 
.A1(n_742),
.A2(n_752),
.B(n_764),
.C(n_776),
.Y(n_1060)
);

AOI21xp5_ASAP7_75t_L g1061 ( 
.A1(n_754),
.A2(n_638),
.B(n_804),
.Y(n_1061)
);

AO21x1_ASAP7_75t_L g1062 ( 
.A1(n_742),
.A2(n_752),
.B(n_802),
.Y(n_1062)
);

AND2x2_ASAP7_75t_L g1063 ( 
.A(n_764),
.B(n_770),
.Y(n_1063)
);

INVx5_ASAP7_75t_L g1064 ( 
.A(n_839),
.Y(n_1064)
);

OAI21xp5_ASAP7_75t_L g1065 ( 
.A1(n_754),
.A2(n_638),
.B(n_759),
.Y(n_1065)
);

NAND2xp5_ASAP7_75t_L g1066 ( 
.A(n_888),
.B(n_742),
.Y(n_1066)
);

AOI21xp5_ASAP7_75t_L g1067 ( 
.A1(n_958),
.A2(n_1053),
.B(n_1041),
.Y(n_1067)
);

OAI21x1_ASAP7_75t_L g1068 ( 
.A1(n_946),
.A2(n_939),
.B(n_903),
.Y(n_1068)
);

INVx2_ASAP7_75t_L g1069 ( 
.A(n_989),
.Y(n_1069)
);

AOI21xp5_ASAP7_75t_L g1070 ( 
.A1(n_1056),
.A2(n_1061),
.B(n_1058),
.Y(n_1070)
);

BUFx2_ASAP7_75t_L g1071 ( 
.A(n_904),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_L g1072 ( 
.A(n_1049),
.B(n_1052),
.Y(n_1072)
);

OAI21x1_ASAP7_75t_L g1073 ( 
.A1(n_915),
.A2(n_905),
.B(n_907),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_L g1074 ( 
.A(n_1060),
.B(n_1051),
.Y(n_1074)
);

AOI21xp5_ASAP7_75t_L g1075 ( 
.A1(n_1004),
.A2(n_1008),
.B(n_1048),
.Y(n_1075)
);

AOI21xp5_ASAP7_75t_L g1076 ( 
.A1(n_1065),
.A2(n_1005),
.B(n_1006),
.Y(n_1076)
);

BUFx6f_ASAP7_75t_L g1077 ( 
.A(n_911),
.Y(n_1077)
);

BUFx6f_ASAP7_75t_L g1078 ( 
.A(n_911),
.Y(n_1078)
);

NAND2x1p5_ASAP7_75t_L g1079 ( 
.A(n_1039),
.B(n_1042),
.Y(n_1079)
);

OAI22xp5_ASAP7_75t_L g1080 ( 
.A1(n_1043),
.A2(n_951),
.B1(n_1066),
.B2(n_1050),
.Y(n_1080)
);

BUFx2_ASAP7_75t_L g1081 ( 
.A(n_913),
.Y(n_1081)
);

AND2x2_ASAP7_75t_L g1082 ( 
.A(n_1063),
.B(n_1045),
.Y(n_1082)
);

HB1xp67_ASAP7_75t_L g1083 ( 
.A(n_941),
.Y(n_1083)
);

AOI21xp5_ASAP7_75t_L g1084 ( 
.A1(n_1005),
.A2(n_902),
.B(n_1022),
.Y(n_1084)
);

NAND2xp5_ASAP7_75t_L g1085 ( 
.A(n_1050),
.B(n_1066),
.Y(n_1085)
);

AOI21xp5_ASAP7_75t_L g1086 ( 
.A1(n_912),
.A2(n_988),
.B(n_1010),
.Y(n_1086)
);

NAND2x1p5_ASAP7_75t_L g1087 ( 
.A(n_1039),
.B(n_1042),
.Y(n_1087)
);

BUFx2_ASAP7_75t_L g1088 ( 
.A(n_975),
.Y(n_1088)
);

BUFx2_ASAP7_75t_L g1089 ( 
.A(n_936),
.Y(n_1089)
);

OAI21x1_ASAP7_75t_L g1090 ( 
.A1(n_921),
.A2(n_927),
.B(n_1007),
.Y(n_1090)
);

AO31x2_ASAP7_75t_L g1091 ( 
.A1(n_1062),
.A2(n_918),
.A3(n_914),
.B(n_1012),
.Y(n_1091)
);

INVx3_ASAP7_75t_L g1092 ( 
.A(n_942),
.Y(n_1092)
);

INVx1_ASAP7_75t_L g1093 ( 
.A(n_957),
.Y(n_1093)
);

NAND2xp5_ASAP7_75t_L g1094 ( 
.A(n_1059),
.B(n_922),
.Y(n_1094)
);

OAI21x1_ASAP7_75t_L g1095 ( 
.A1(n_919),
.A2(n_1030),
.B(n_920),
.Y(n_1095)
);

NAND2xp5_ASAP7_75t_SL g1096 ( 
.A(n_1019),
.B(n_899),
.Y(n_1096)
);

OAI21x1_ASAP7_75t_L g1097 ( 
.A1(n_919),
.A2(n_917),
.B(n_1025),
.Y(n_1097)
);

INVx2_ASAP7_75t_SL g1098 ( 
.A(n_1047),
.Y(n_1098)
);

CKINVDCx20_ASAP7_75t_R g1099 ( 
.A(n_965),
.Y(n_1099)
);

A2O1A1Ixp33_ASAP7_75t_L g1100 ( 
.A1(n_1054),
.A2(n_1057),
.B(n_1014),
.C(n_937),
.Y(n_1100)
);

INVx3_ASAP7_75t_L g1101 ( 
.A(n_942),
.Y(n_1101)
);

AOI21xp5_ASAP7_75t_L g1102 ( 
.A1(n_900),
.A2(n_901),
.B(n_940),
.Y(n_1102)
);

A2O1A1Ixp33_ASAP7_75t_L g1103 ( 
.A1(n_1021),
.A2(n_986),
.B(n_982),
.C(n_991),
.Y(n_1103)
);

AOI21xp33_ASAP7_75t_L g1104 ( 
.A1(n_1002),
.A2(n_1033),
.B(n_924),
.Y(n_1104)
);

NOR2xp33_ASAP7_75t_L g1105 ( 
.A(n_926),
.B(n_1038),
.Y(n_1105)
);

OAI21xp5_ASAP7_75t_L g1106 ( 
.A1(n_970),
.A2(n_971),
.B(n_1027),
.Y(n_1106)
);

NAND2xp5_ASAP7_75t_SL g1107 ( 
.A(n_952),
.B(n_933),
.Y(n_1107)
);

O2A1O1Ixp5_ASAP7_75t_L g1108 ( 
.A1(n_1024),
.A2(n_908),
.B(n_1032),
.C(n_1034),
.Y(n_1108)
);

OAI21x1_ASAP7_75t_L g1109 ( 
.A1(n_1015),
.A2(n_950),
.B(n_909),
.Y(n_1109)
);

AOI21xp5_ASAP7_75t_L g1110 ( 
.A1(n_900),
.A2(n_970),
.B(n_971),
.Y(n_1110)
);

OAI21x1_ASAP7_75t_SL g1111 ( 
.A1(n_981),
.A2(n_973),
.B(n_972),
.Y(n_1111)
);

NAND2xp5_ASAP7_75t_L g1112 ( 
.A(n_1009),
.B(n_908),
.Y(n_1112)
);

NAND2x1p5_ASAP7_75t_L g1113 ( 
.A(n_1039),
.B(n_1042),
.Y(n_1113)
);

OAI21x1_ASAP7_75t_L g1114 ( 
.A1(n_909),
.A2(n_947),
.B(n_943),
.Y(n_1114)
);

AND2x2_ASAP7_75t_L g1115 ( 
.A(n_930),
.B(n_998),
.Y(n_1115)
);

AND2x4_ASAP7_75t_L g1116 ( 
.A(n_1023),
.B(n_1000),
.Y(n_1116)
);

OAI22xp33_ASAP7_75t_L g1117 ( 
.A1(n_1038),
.A2(n_993),
.B1(n_1017),
.B2(n_928),
.Y(n_1117)
);

NAND2xp5_ASAP7_75t_SL g1118 ( 
.A(n_1020),
.B(n_961),
.Y(n_1118)
);

NOR2xp33_ASAP7_75t_SL g1119 ( 
.A(n_984),
.B(n_967),
.Y(n_1119)
);

OAI21x1_ASAP7_75t_L g1120 ( 
.A1(n_916),
.A2(n_964),
.B(n_954),
.Y(n_1120)
);

AOI21xp5_ASAP7_75t_L g1121 ( 
.A1(n_1031),
.A2(n_981),
.B(n_972),
.Y(n_1121)
);

OAI21x1_ASAP7_75t_L g1122 ( 
.A1(n_906),
.A2(n_973),
.B(n_945),
.Y(n_1122)
);

OAI22xp5_ASAP7_75t_L g1123 ( 
.A1(n_966),
.A2(n_959),
.B1(n_994),
.B2(n_990),
.Y(n_1123)
);

OAI21xp5_ASAP7_75t_L g1124 ( 
.A1(n_1024),
.A2(n_966),
.B(n_948),
.Y(n_1124)
);

BUFx2_ASAP7_75t_L g1125 ( 
.A(n_992),
.Y(n_1125)
);

OAI22xp5_ASAP7_75t_L g1126 ( 
.A1(n_990),
.A2(n_994),
.B1(n_969),
.B2(n_961),
.Y(n_1126)
);

A2O1A1Ixp33_ASAP7_75t_L g1127 ( 
.A1(n_935),
.A2(n_934),
.B(n_1029),
.C(n_938),
.Y(n_1127)
);

AND2x4_ASAP7_75t_L g1128 ( 
.A(n_1000),
.B(n_960),
.Y(n_1128)
);

BUFx6f_ASAP7_75t_L g1129 ( 
.A(n_942),
.Y(n_1129)
);

AOI21xp5_ASAP7_75t_L g1130 ( 
.A1(n_1013),
.A2(n_980),
.B(n_949),
.Y(n_1130)
);

OAI21x1_ASAP7_75t_L g1131 ( 
.A1(n_1011),
.A2(n_944),
.B(n_1016),
.Y(n_1131)
);

BUFx2_ASAP7_75t_SL g1132 ( 
.A(n_923),
.Y(n_1132)
);

AOI21xp5_ASAP7_75t_L g1133 ( 
.A1(n_949),
.A2(n_953),
.B(n_1035),
.Y(n_1133)
);

INVx2_ASAP7_75t_L g1134 ( 
.A(n_910),
.Y(n_1134)
);

NAND2xp5_ASAP7_75t_L g1135 ( 
.A(n_976),
.B(n_931),
.Y(n_1135)
);

NAND2xp5_ASAP7_75t_SL g1136 ( 
.A(n_978),
.B(n_955),
.Y(n_1136)
);

O2A1O1Ixp5_ASAP7_75t_L g1137 ( 
.A1(n_985),
.A2(n_983),
.B(n_956),
.C(n_1040),
.Y(n_1137)
);

OAI21x1_ASAP7_75t_L g1138 ( 
.A1(n_963),
.A2(n_979),
.B(n_977),
.Y(n_1138)
);

CKINVDCx5p33_ASAP7_75t_R g1139 ( 
.A(n_1003),
.Y(n_1139)
);

AO21x1_ASAP7_75t_L g1140 ( 
.A1(n_969),
.A2(n_929),
.B(n_987),
.Y(n_1140)
);

INVx2_ASAP7_75t_L g1141 ( 
.A(n_925),
.Y(n_1141)
);

OAI222xp33_ASAP7_75t_L g1142 ( 
.A1(n_1017),
.A2(n_996),
.B1(n_1026),
.B2(n_1046),
.C1(n_932),
.C2(n_1044),
.Y(n_1142)
);

INVx5_ASAP7_75t_L g1143 ( 
.A(n_974),
.Y(n_1143)
);

AOI21xp33_ASAP7_75t_L g1144 ( 
.A1(n_1001),
.A2(n_928),
.B(n_968),
.Y(n_1144)
);

OAI21xp5_ASAP7_75t_L g1145 ( 
.A1(n_962),
.A2(n_999),
.B(n_1018),
.Y(n_1145)
);

AOI21xp5_ASAP7_75t_L g1146 ( 
.A1(n_1039),
.A2(n_1064),
.B(n_1042),
.Y(n_1146)
);

NAND2xp5_ASAP7_75t_L g1147 ( 
.A(n_955),
.B(n_1064),
.Y(n_1147)
);

INVx1_ASAP7_75t_L g1148 ( 
.A(n_992),
.Y(n_1148)
);

OAI21x1_ASAP7_75t_L g1149 ( 
.A1(n_1064),
.A2(n_1028),
.B(n_1037),
.Y(n_1149)
);

AOI21x1_ASAP7_75t_L g1150 ( 
.A1(n_997),
.A2(n_955),
.B(n_974),
.Y(n_1150)
);

OAI21x1_ASAP7_75t_L g1151 ( 
.A1(n_1064),
.A2(n_974),
.B(n_967),
.Y(n_1151)
);

AO31x2_ASAP7_75t_L g1152 ( 
.A1(n_974),
.A2(n_923),
.A3(n_1055),
.B(n_1036),
.Y(n_1152)
);

AND2x4_ASAP7_75t_L g1153 ( 
.A(n_923),
.B(n_995),
.Y(n_1153)
);

OAI21x1_ASAP7_75t_L g1154 ( 
.A1(n_923),
.A2(n_946),
.B(n_939),
.Y(n_1154)
);

OAI21x1_ASAP7_75t_L g1155 ( 
.A1(n_946),
.A2(n_939),
.B(n_903),
.Y(n_1155)
);

NAND2xp5_ASAP7_75t_L g1156 ( 
.A(n_1049),
.B(n_1052),
.Y(n_1156)
);

AND2x2_ASAP7_75t_L g1157 ( 
.A(n_1051),
.B(n_1063),
.Y(n_1157)
);

OAI21x1_ASAP7_75t_L g1158 ( 
.A1(n_946),
.A2(n_939),
.B(n_903),
.Y(n_1158)
);

AOI21xp5_ASAP7_75t_L g1159 ( 
.A1(n_958),
.A2(n_1053),
.B(n_1041),
.Y(n_1159)
);

AOI21xp5_ASAP7_75t_SL g1160 ( 
.A1(n_1060),
.A2(n_981),
.B(n_839),
.Y(n_1160)
);

INVx2_ASAP7_75t_SL g1161 ( 
.A(n_936),
.Y(n_1161)
);

OAI21x1_ASAP7_75t_L g1162 ( 
.A1(n_946),
.A2(n_939),
.B(n_903),
.Y(n_1162)
);

BUFx6f_ASAP7_75t_L g1163 ( 
.A(n_911),
.Y(n_1163)
);

NAND2xp5_ASAP7_75t_L g1164 ( 
.A(n_1049),
.B(n_1052),
.Y(n_1164)
);

AOI21xp5_ASAP7_75t_L g1165 ( 
.A1(n_958),
.A2(n_1053),
.B(n_1041),
.Y(n_1165)
);

OAI21xp5_ASAP7_75t_SL g1166 ( 
.A1(n_1049),
.A2(n_1052),
.B(n_951),
.Y(n_1166)
);

NAND2xp5_ASAP7_75t_L g1167 ( 
.A(n_1049),
.B(n_1052),
.Y(n_1167)
);

OAI21xp5_ASAP7_75t_L g1168 ( 
.A1(n_1060),
.A2(n_1043),
.B(n_1004),
.Y(n_1168)
);

BUFx12f_ASAP7_75t_L g1169 ( 
.A(n_904),
.Y(n_1169)
);

OAI21x1_ASAP7_75t_L g1170 ( 
.A1(n_946),
.A2(n_939),
.B(n_903),
.Y(n_1170)
);

NOR2xp33_ASAP7_75t_L g1171 ( 
.A(n_1049),
.B(n_1052),
.Y(n_1171)
);

AO31x2_ASAP7_75t_L g1172 ( 
.A1(n_1062),
.A2(n_1060),
.A3(n_918),
.B(n_914),
.Y(n_1172)
);

AOI21xp5_ASAP7_75t_L g1173 ( 
.A1(n_958),
.A2(n_1053),
.B(n_1041),
.Y(n_1173)
);

AOI21xp5_ASAP7_75t_L g1174 ( 
.A1(n_958),
.A2(n_1053),
.B(n_1041),
.Y(n_1174)
);

NAND2xp5_ASAP7_75t_L g1175 ( 
.A(n_1049),
.B(n_1052),
.Y(n_1175)
);

OAI21x1_ASAP7_75t_L g1176 ( 
.A1(n_946),
.A2(n_939),
.B(n_903),
.Y(n_1176)
);

INVx2_ASAP7_75t_SL g1177 ( 
.A(n_936),
.Y(n_1177)
);

NAND2xp5_ASAP7_75t_L g1178 ( 
.A(n_1049),
.B(n_1052),
.Y(n_1178)
);

AO31x2_ASAP7_75t_L g1179 ( 
.A1(n_1062),
.A2(n_1060),
.A3(n_918),
.B(n_914),
.Y(n_1179)
);

A2O1A1Ixp33_ASAP7_75t_L g1180 ( 
.A1(n_1049),
.A2(n_1052),
.B(n_951),
.C(n_1043),
.Y(n_1180)
);

AOI21x1_ASAP7_75t_L g1181 ( 
.A1(n_915),
.A2(n_927),
.B(n_900),
.Y(n_1181)
);

NAND2xp5_ASAP7_75t_L g1182 ( 
.A(n_1049),
.B(n_1052),
.Y(n_1182)
);

NAND2xp5_ASAP7_75t_L g1183 ( 
.A(n_1049),
.B(n_1052),
.Y(n_1183)
);

OAI21x1_ASAP7_75t_SL g1184 ( 
.A1(n_981),
.A2(n_973),
.B(n_972),
.Y(n_1184)
);

AND2x2_ASAP7_75t_L g1185 ( 
.A(n_1051),
.B(n_1063),
.Y(n_1185)
);

AO31x2_ASAP7_75t_L g1186 ( 
.A1(n_1062),
.A2(n_1060),
.A3(n_918),
.B(n_914),
.Y(n_1186)
);

NOR2xp33_ASAP7_75t_L g1187 ( 
.A(n_1049),
.B(n_1052),
.Y(n_1187)
);

INVx3_ASAP7_75t_L g1188 ( 
.A(n_911),
.Y(n_1188)
);

AO31x2_ASAP7_75t_L g1189 ( 
.A1(n_1062),
.A2(n_1060),
.A3(n_918),
.B(n_914),
.Y(n_1189)
);

OAI21x1_ASAP7_75t_L g1190 ( 
.A1(n_946),
.A2(n_939),
.B(n_903),
.Y(n_1190)
);

OAI21x1_ASAP7_75t_L g1191 ( 
.A1(n_946),
.A2(n_939),
.B(n_903),
.Y(n_1191)
);

BUFx2_ASAP7_75t_L g1192 ( 
.A(n_904),
.Y(n_1192)
);

AOI21xp5_ASAP7_75t_L g1193 ( 
.A1(n_958),
.A2(n_1053),
.B(n_1041),
.Y(n_1193)
);

NAND2x1_ASAP7_75t_L g1194 ( 
.A(n_906),
.B(n_761),
.Y(n_1194)
);

OAI21x1_ASAP7_75t_L g1195 ( 
.A1(n_946),
.A2(n_939),
.B(n_903),
.Y(n_1195)
);

AOI21xp5_ASAP7_75t_L g1196 ( 
.A1(n_958),
.A2(n_1053),
.B(n_1041),
.Y(n_1196)
);

AOI21xp5_ASAP7_75t_L g1197 ( 
.A1(n_958),
.A2(n_1053),
.B(n_1041),
.Y(n_1197)
);

OAI22x1_ASAP7_75t_L g1198 ( 
.A1(n_1049),
.A2(n_1052),
.B1(n_951),
.B2(n_1043),
.Y(n_1198)
);

AND2x4_ASAP7_75t_L g1199 ( 
.A(n_1023),
.B(n_1000),
.Y(n_1199)
);

OAI21x1_ASAP7_75t_L g1200 ( 
.A1(n_946),
.A2(n_939),
.B(n_903),
.Y(n_1200)
);

INVx2_ASAP7_75t_SL g1201 ( 
.A(n_936),
.Y(n_1201)
);

BUFx6f_ASAP7_75t_L g1202 ( 
.A(n_911),
.Y(n_1202)
);

AOI21xp5_ASAP7_75t_L g1203 ( 
.A1(n_958),
.A2(n_1053),
.B(n_1041),
.Y(n_1203)
);

OAI21x1_ASAP7_75t_L g1204 ( 
.A1(n_946),
.A2(n_939),
.B(n_903),
.Y(n_1204)
);

NAND2xp5_ASAP7_75t_L g1205 ( 
.A(n_1049),
.B(n_1052),
.Y(n_1205)
);

OAI21x1_ASAP7_75t_L g1206 ( 
.A1(n_946),
.A2(n_939),
.B(n_903),
.Y(n_1206)
);

AOI21xp5_ASAP7_75t_L g1207 ( 
.A1(n_958),
.A2(n_1053),
.B(n_1041),
.Y(n_1207)
);

NAND2xp5_ASAP7_75t_L g1208 ( 
.A(n_1049),
.B(n_1052),
.Y(n_1208)
);

NAND2xp5_ASAP7_75t_L g1209 ( 
.A(n_1049),
.B(n_1052),
.Y(n_1209)
);

INVx5_ASAP7_75t_L g1210 ( 
.A(n_974),
.Y(n_1210)
);

OAI21x1_ASAP7_75t_L g1211 ( 
.A1(n_946),
.A2(n_939),
.B(n_903),
.Y(n_1211)
);

INVx3_ASAP7_75t_L g1212 ( 
.A(n_1143),
.Y(n_1212)
);

HB1xp67_ASAP7_75t_L g1213 ( 
.A(n_1081),
.Y(n_1213)
);

NOR2xp33_ASAP7_75t_SL g1214 ( 
.A(n_1099),
.B(n_1119),
.Y(n_1214)
);

OR2x2_ASAP7_75t_L g1215 ( 
.A(n_1166),
.B(n_1072),
.Y(n_1215)
);

AOI22xp5_ASAP7_75t_L g1216 ( 
.A1(n_1171),
.A2(n_1187),
.B1(n_1096),
.B2(n_1164),
.Y(n_1216)
);

NAND2xp5_ASAP7_75t_L g1217 ( 
.A(n_1072),
.B(n_1156),
.Y(n_1217)
);

AND2x2_ASAP7_75t_SL g1218 ( 
.A(n_1156),
.B(n_1164),
.Y(n_1218)
);

AOI21xp5_ASAP7_75t_L g1219 ( 
.A1(n_1067),
.A2(n_1165),
.B(n_1159),
.Y(n_1219)
);

AND2x4_ASAP7_75t_L g1220 ( 
.A(n_1128),
.B(n_1116),
.Y(n_1220)
);

AND2x4_ASAP7_75t_L g1221 ( 
.A(n_1128),
.B(n_1116),
.Y(n_1221)
);

NAND3xp33_ASAP7_75t_L g1222 ( 
.A(n_1180),
.B(n_1175),
.C(n_1167),
.Y(n_1222)
);

O2A1O1Ixp33_ASAP7_75t_L g1223 ( 
.A1(n_1167),
.A2(n_1209),
.B(n_1178),
.C(n_1205),
.Y(n_1223)
);

AND2x4_ASAP7_75t_L g1224 ( 
.A(n_1199),
.B(n_1148),
.Y(n_1224)
);

AND2x4_ASAP7_75t_L g1225 ( 
.A(n_1199),
.B(n_1125),
.Y(n_1225)
);

NAND2xp5_ASAP7_75t_L g1226 ( 
.A(n_1175),
.B(n_1178),
.Y(n_1226)
);

AOI22xp5_ASAP7_75t_L g1227 ( 
.A1(n_1182),
.A2(n_1205),
.B1(n_1183),
.B2(n_1208),
.Y(n_1227)
);

INVx5_ASAP7_75t_L g1228 ( 
.A(n_1143),
.Y(n_1228)
);

A2O1A1Ixp33_ASAP7_75t_L g1229 ( 
.A1(n_1100),
.A2(n_1121),
.B(n_1103),
.C(n_1182),
.Y(n_1229)
);

AND2x4_ASAP7_75t_L g1230 ( 
.A(n_1153),
.B(n_1141),
.Y(n_1230)
);

NAND2xp5_ASAP7_75t_L g1231 ( 
.A(n_1183),
.B(n_1208),
.Y(n_1231)
);

INVxp33_ASAP7_75t_L g1232 ( 
.A(n_1071),
.Y(n_1232)
);

OAI22xp5_ASAP7_75t_L g1233 ( 
.A1(n_1209),
.A2(n_1085),
.B1(n_1126),
.B2(n_1112),
.Y(n_1233)
);

CKINVDCx5p33_ASAP7_75t_R g1234 ( 
.A(n_1169),
.Y(n_1234)
);

INVxp67_ASAP7_75t_SL g1235 ( 
.A(n_1098),
.Y(n_1235)
);

CKINVDCx11_ASAP7_75t_R g1236 ( 
.A(n_1192),
.Y(n_1236)
);

INVx1_ASAP7_75t_SL g1237 ( 
.A(n_1089),
.Y(n_1237)
);

INVx1_ASAP7_75t_L g1238 ( 
.A(n_1135),
.Y(n_1238)
);

AOI21xp5_ASAP7_75t_L g1239 ( 
.A1(n_1067),
.A2(n_1207),
.B(n_1203),
.Y(n_1239)
);

NAND2xp5_ASAP7_75t_L g1240 ( 
.A(n_1085),
.B(n_1112),
.Y(n_1240)
);

NAND2xp5_ASAP7_75t_L g1241 ( 
.A(n_1080),
.B(n_1094),
.Y(n_1241)
);

AND2x4_ASAP7_75t_L g1242 ( 
.A(n_1153),
.B(n_1069),
.Y(n_1242)
);

OAI22xp5_ASAP7_75t_L g1243 ( 
.A1(n_1126),
.A2(n_1123),
.B1(n_1117),
.B2(n_1105),
.Y(n_1243)
);

AND2x2_ASAP7_75t_L g1244 ( 
.A(n_1082),
.B(n_1115),
.Y(n_1244)
);

OAI21xp5_ASAP7_75t_L g1245 ( 
.A1(n_1076),
.A2(n_1075),
.B(n_1124),
.Y(n_1245)
);

NAND2xp5_ASAP7_75t_SL g1246 ( 
.A(n_1080),
.B(n_1198),
.Y(n_1246)
);

NAND2xp5_ASAP7_75t_L g1247 ( 
.A(n_1094),
.B(n_1074),
.Y(n_1247)
);

AOI21xp5_ASAP7_75t_L g1248 ( 
.A1(n_1159),
.A2(n_1207),
.B(n_1197),
.Y(n_1248)
);

NAND2xp5_ASAP7_75t_L g1249 ( 
.A(n_1074),
.B(n_1168),
.Y(n_1249)
);

O2A1O1Ixp33_ASAP7_75t_SL g1250 ( 
.A1(n_1127),
.A2(n_1144),
.B(n_1118),
.C(n_1123),
.Y(n_1250)
);

CKINVDCx5p33_ASAP7_75t_R g1251 ( 
.A(n_1139),
.Y(n_1251)
);

OAI22xp5_ASAP7_75t_L g1252 ( 
.A1(n_1143),
.A2(n_1210),
.B1(n_1160),
.B2(n_1076),
.Y(n_1252)
);

OAI21x1_ASAP7_75t_L g1253 ( 
.A1(n_1154),
.A2(n_1114),
.B(n_1211),
.Y(n_1253)
);

NOR2xp33_ASAP7_75t_L g1254 ( 
.A(n_1107),
.B(n_1161),
.Y(n_1254)
);

BUFx2_ASAP7_75t_L g1255 ( 
.A(n_1088),
.Y(n_1255)
);

INVx2_ASAP7_75t_SL g1256 ( 
.A(n_1177),
.Y(n_1256)
);

BUFx6f_ASAP7_75t_L g1257 ( 
.A(n_1077),
.Y(n_1257)
);

HB1xp67_ASAP7_75t_L g1258 ( 
.A(n_1083),
.Y(n_1258)
);

INVxp67_ASAP7_75t_L g1259 ( 
.A(n_1201),
.Y(n_1259)
);

NOR4xp25_ASAP7_75t_L g1260 ( 
.A(n_1144),
.B(n_1145),
.C(n_1142),
.D(n_1106),
.Y(n_1260)
);

BUFx3_ASAP7_75t_L g1261 ( 
.A(n_1077),
.Y(n_1261)
);

OAI21xp5_ASAP7_75t_L g1262 ( 
.A1(n_1075),
.A2(n_1121),
.B(n_1108),
.Y(n_1262)
);

CKINVDCx11_ASAP7_75t_R g1263 ( 
.A(n_1077),
.Y(n_1263)
);

AOI21xp5_ASAP7_75t_L g1264 ( 
.A1(n_1086),
.A2(n_1173),
.B(n_1196),
.Y(n_1264)
);

AOI21xp5_ASAP7_75t_L g1265 ( 
.A1(n_1086),
.A2(n_1173),
.B(n_1196),
.Y(n_1265)
);

A2O1A1Ixp33_ASAP7_75t_L g1266 ( 
.A1(n_1133),
.A2(n_1104),
.B(n_1110),
.C(n_1084),
.Y(n_1266)
);

A2O1A1Ixp33_ASAP7_75t_L g1267 ( 
.A1(n_1133),
.A2(n_1104),
.B(n_1110),
.C(n_1084),
.Y(n_1267)
);

INVx2_ASAP7_75t_L g1268 ( 
.A(n_1092),
.Y(n_1268)
);

HB1xp67_ASAP7_75t_L g1269 ( 
.A(n_1078),
.Y(n_1269)
);

INVx2_ASAP7_75t_L g1270 ( 
.A(n_1092),
.Y(n_1270)
);

INVx1_ASAP7_75t_L g1271 ( 
.A(n_1136),
.Y(n_1271)
);

NOR2xp33_ASAP7_75t_L g1272 ( 
.A(n_1140),
.B(n_1150),
.Y(n_1272)
);

AND2x4_ASAP7_75t_L g1273 ( 
.A(n_1149),
.B(n_1210),
.Y(n_1273)
);

OA21x2_ASAP7_75t_L g1274 ( 
.A1(n_1070),
.A2(n_1102),
.B(n_1165),
.Y(n_1274)
);

AOI221xp5_ASAP7_75t_L g1275 ( 
.A1(n_1111),
.A2(n_1184),
.B1(n_1174),
.B2(n_1193),
.C(n_1130),
.Y(n_1275)
);

OAI22xp5_ASAP7_75t_L g1276 ( 
.A1(n_1143),
.A2(n_1210),
.B1(n_1132),
.B2(n_1174),
.Y(n_1276)
);

BUFx6f_ASAP7_75t_L g1277 ( 
.A(n_1078),
.Y(n_1277)
);

AOI21xp5_ASAP7_75t_L g1278 ( 
.A1(n_1070),
.A2(n_1073),
.B(n_1137),
.Y(n_1278)
);

CKINVDCx16_ASAP7_75t_R g1279 ( 
.A(n_1078),
.Y(n_1279)
);

INVx1_ASAP7_75t_L g1280 ( 
.A(n_1101),
.Y(n_1280)
);

INVxp67_ASAP7_75t_L g1281 ( 
.A(n_1129),
.Y(n_1281)
);

INVx1_ASAP7_75t_L g1282 ( 
.A(n_1101),
.Y(n_1282)
);

BUFx12f_ASAP7_75t_L g1283 ( 
.A(n_1129),
.Y(n_1283)
);

AOI22xp33_ASAP7_75t_L g1284 ( 
.A1(n_1210),
.A2(n_1188),
.B1(n_1130),
.B2(n_1202),
.Y(n_1284)
);

CKINVDCx8_ASAP7_75t_R g1285 ( 
.A(n_1129),
.Y(n_1285)
);

INVx1_ASAP7_75t_SL g1286 ( 
.A(n_1163),
.Y(n_1286)
);

AOI21xp5_ASAP7_75t_L g1287 ( 
.A1(n_1146),
.A2(n_1095),
.B(n_1158),
.Y(n_1287)
);

AOI21xp5_ASAP7_75t_L g1288 ( 
.A1(n_1146),
.A2(n_1068),
.B(n_1206),
.Y(n_1288)
);

NOR2x1_ASAP7_75t_L g1289 ( 
.A(n_1188),
.B(n_1147),
.Y(n_1289)
);

INVx2_ASAP7_75t_SL g1290 ( 
.A(n_1163),
.Y(n_1290)
);

AND2x4_ASAP7_75t_L g1291 ( 
.A(n_1152),
.B(n_1151),
.Y(n_1291)
);

NAND2x1_ASAP7_75t_L g1292 ( 
.A(n_1163),
.B(n_1202),
.Y(n_1292)
);

OR2x6_ASAP7_75t_SL g1293 ( 
.A(n_1147),
.B(n_1152),
.Y(n_1293)
);

AND2x2_ASAP7_75t_L g1294 ( 
.A(n_1152),
.B(n_1091),
.Y(n_1294)
);

CKINVDCx5p33_ASAP7_75t_R g1295 ( 
.A(n_1194),
.Y(n_1295)
);

BUFx6f_ASAP7_75t_L g1296 ( 
.A(n_1079),
.Y(n_1296)
);

AND2x2_ASAP7_75t_L g1297 ( 
.A(n_1091),
.B(n_1186),
.Y(n_1297)
);

AOI21xp5_ASAP7_75t_L g1298 ( 
.A1(n_1155),
.A2(n_1204),
.B(n_1162),
.Y(n_1298)
);

AOI21xp5_ASAP7_75t_SL g1299 ( 
.A1(n_1079),
.A2(n_1113),
.B(n_1087),
.Y(n_1299)
);

BUFx2_ASAP7_75t_L g1300 ( 
.A(n_1091),
.Y(n_1300)
);

BUFx2_ASAP7_75t_L g1301 ( 
.A(n_1087),
.Y(n_1301)
);

AOI21xp5_ASAP7_75t_L g1302 ( 
.A1(n_1170),
.A2(n_1200),
.B(n_1195),
.Y(n_1302)
);

NAND2xp5_ASAP7_75t_SL g1303 ( 
.A(n_1113),
.B(n_1122),
.Y(n_1303)
);

INVx1_ASAP7_75t_L g1304 ( 
.A(n_1172),
.Y(n_1304)
);

AND2x2_ASAP7_75t_L g1305 ( 
.A(n_1179),
.B(n_1189),
.Y(n_1305)
);

OA21x2_ASAP7_75t_L g1306 ( 
.A1(n_1097),
.A2(n_1191),
.B(n_1190),
.Y(n_1306)
);

NAND2xp5_ASAP7_75t_SL g1307 ( 
.A(n_1181),
.B(n_1131),
.Y(n_1307)
);

AND2x2_ASAP7_75t_L g1308 ( 
.A(n_1179),
.B(n_1189),
.Y(n_1308)
);

BUFx3_ASAP7_75t_L g1309 ( 
.A(n_1090),
.Y(n_1309)
);

AOI22xp33_ASAP7_75t_L g1310 ( 
.A1(n_1138),
.A2(n_1109),
.B1(n_1176),
.B2(n_1120),
.Y(n_1310)
);

OAI22xp5_ASAP7_75t_L g1311 ( 
.A1(n_1171),
.A2(n_1187),
.B1(n_1049),
.B2(n_1052),
.Y(n_1311)
);

INVxp67_ASAP7_75t_L g1312 ( 
.A(n_1098),
.Y(n_1312)
);

BUFx2_ASAP7_75t_L g1313 ( 
.A(n_1081),
.Y(n_1313)
);

NAND2xp5_ASAP7_75t_L g1314 ( 
.A(n_1171),
.B(n_1187),
.Y(n_1314)
);

AND2x2_ASAP7_75t_L g1315 ( 
.A(n_1157),
.B(n_1185),
.Y(n_1315)
);

OAI22xp5_ASAP7_75t_L g1316 ( 
.A1(n_1171),
.A2(n_1187),
.B1(n_1049),
.B2(n_1052),
.Y(n_1316)
);

AOI21xp5_ASAP7_75t_L g1317 ( 
.A1(n_1067),
.A2(n_1165),
.B(n_1159),
.Y(n_1317)
);

OAI22xp5_ASAP7_75t_L g1318 ( 
.A1(n_1171),
.A2(n_1187),
.B1(n_1049),
.B2(n_1052),
.Y(n_1318)
);

OAI22xp5_ASAP7_75t_L g1319 ( 
.A1(n_1171),
.A2(n_1187),
.B1(n_1049),
.B2(n_1052),
.Y(n_1319)
);

BUFx6f_ASAP7_75t_L g1320 ( 
.A(n_1077),
.Y(n_1320)
);

NAND2xp5_ASAP7_75t_L g1321 ( 
.A(n_1171),
.B(n_1187),
.Y(n_1321)
);

OR2x6_ASAP7_75t_L g1322 ( 
.A(n_1132),
.B(n_823),
.Y(n_1322)
);

OR2x2_ASAP7_75t_L g1323 ( 
.A(n_1166),
.B(n_1045),
.Y(n_1323)
);

INVx3_ASAP7_75t_L g1324 ( 
.A(n_1143),
.Y(n_1324)
);

NOR2xp33_ASAP7_75t_L g1325 ( 
.A(n_1171),
.B(n_1049),
.Y(n_1325)
);

INVx1_ASAP7_75t_L g1326 ( 
.A(n_1093),
.Y(n_1326)
);

AND2x2_ASAP7_75t_L g1327 ( 
.A(n_1157),
.B(n_1185),
.Y(n_1327)
);

INVx5_ASAP7_75t_L g1328 ( 
.A(n_1143),
.Y(n_1328)
);

OAI221xp5_ASAP7_75t_L g1329 ( 
.A1(n_1171),
.A2(n_1049),
.B1(n_1052),
.B2(n_1187),
.C(n_1166),
.Y(n_1329)
);

INVx2_ASAP7_75t_L g1330 ( 
.A(n_1134),
.Y(n_1330)
);

OAI22xp5_ASAP7_75t_L g1331 ( 
.A1(n_1171),
.A2(n_1187),
.B1(n_1049),
.B2(n_1052),
.Y(n_1331)
);

NAND2xp5_ASAP7_75t_L g1332 ( 
.A(n_1171),
.B(n_1187),
.Y(n_1332)
);

INVx1_ASAP7_75t_L g1333 ( 
.A(n_1093),
.Y(n_1333)
);

NAND2xp5_ASAP7_75t_L g1334 ( 
.A(n_1171),
.B(n_1187),
.Y(n_1334)
);

AOI21xp5_ASAP7_75t_L g1335 ( 
.A1(n_1067),
.A2(n_1165),
.B(n_1159),
.Y(n_1335)
);

AND2x4_ASAP7_75t_L g1336 ( 
.A(n_1128),
.B(n_1116),
.Y(n_1336)
);

NAND2xp5_ASAP7_75t_L g1337 ( 
.A(n_1171),
.B(n_1187),
.Y(n_1337)
);

INVx3_ASAP7_75t_SL g1338 ( 
.A(n_1139),
.Y(n_1338)
);

NAND2xp5_ASAP7_75t_L g1339 ( 
.A(n_1171),
.B(n_1187),
.Y(n_1339)
);

INVx5_ASAP7_75t_L g1340 ( 
.A(n_1143),
.Y(n_1340)
);

INVx2_ASAP7_75t_L g1341 ( 
.A(n_1134),
.Y(n_1341)
);

INVx2_ASAP7_75t_L g1342 ( 
.A(n_1134),
.Y(n_1342)
);

INVx2_ASAP7_75t_L g1343 ( 
.A(n_1134),
.Y(n_1343)
);

AND2x2_ASAP7_75t_L g1344 ( 
.A(n_1157),
.B(n_1185),
.Y(n_1344)
);

AND2x2_ASAP7_75t_L g1345 ( 
.A(n_1157),
.B(n_1185),
.Y(n_1345)
);

AND2x2_ASAP7_75t_L g1346 ( 
.A(n_1157),
.B(n_1185),
.Y(n_1346)
);

INVx1_ASAP7_75t_L g1347 ( 
.A(n_1093),
.Y(n_1347)
);

INVx3_ASAP7_75t_L g1348 ( 
.A(n_1143),
.Y(n_1348)
);

NOR2xp33_ASAP7_75t_L g1349 ( 
.A(n_1171),
.B(n_1049),
.Y(n_1349)
);

NAND2xp5_ASAP7_75t_L g1350 ( 
.A(n_1171),
.B(n_1187),
.Y(n_1350)
);

NOR2xp33_ASAP7_75t_L g1351 ( 
.A(n_1171),
.B(n_1049),
.Y(n_1351)
);

INVx1_ASAP7_75t_L g1352 ( 
.A(n_1093),
.Y(n_1352)
);

NAND2xp5_ASAP7_75t_L g1353 ( 
.A(n_1171),
.B(n_1187),
.Y(n_1353)
);

INVx2_ASAP7_75t_L g1354 ( 
.A(n_1134),
.Y(n_1354)
);

INVx2_ASAP7_75t_SL g1355 ( 
.A(n_1169),
.Y(n_1355)
);

AND2x2_ASAP7_75t_L g1356 ( 
.A(n_1157),
.B(n_1185),
.Y(n_1356)
);

NAND2xp5_ASAP7_75t_L g1357 ( 
.A(n_1171),
.B(n_1187),
.Y(n_1357)
);

BUFx2_ASAP7_75t_L g1358 ( 
.A(n_1293),
.Y(n_1358)
);

BUFx6f_ASAP7_75t_L g1359 ( 
.A(n_1228),
.Y(n_1359)
);

CKINVDCx14_ASAP7_75t_R g1360 ( 
.A(n_1236),
.Y(n_1360)
);

OR2x6_ASAP7_75t_L g1361 ( 
.A(n_1252),
.B(n_1219),
.Y(n_1361)
);

AOI22xp33_ASAP7_75t_L g1362 ( 
.A1(n_1325),
.A2(n_1349),
.B1(n_1351),
.B2(n_1329),
.Y(n_1362)
);

INVx1_ASAP7_75t_L g1363 ( 
.A(n_1304),
.Y(n_1363)
);

BUFx8_ASAP7_75t_SL g1364 ( 
.A(n_1251),
.Y(n_1364)
);

AOI22xp33_ASAP7_75t_L g1365 ( 
.A1(n_1329),
.A2(n_1319),
.B1(n_1318),
.B2(n_1311),
.Y(n_1365)
);

HB1xp67_ASAP7_75t_L g1366 ( 
.A(n_1213),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_1305),
.Y(n_1367)
);

AND2x2_ASAP7_75t_L g1368 ( 
.A(n_1215),
.B(n_1218),
.Y(n_1368)
);

INVx1_ASAP7_75t_L g1369 ( 
.A(n_1308),
.Y(n_1369)
);

CKINVDCx11_ASAP7_75t_R g1370 ( 
.A(n_1338),
.Y(n_1370)
);

INVx6_ASAP7_75t_L g1371 ( 
.A(n_1228),
.Y(n_1371)
);

HB1xp67_ASAP7_75t_L g1372 ( 
.A(n_1258),
.Y(n_1372)
);

NAND2x1p5_ASAP7_75t_L g1373 ( 
.A(n_1228),
.B(n_1328),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_1300),
.Y(n_1374)
);

OAI21x1_ASAP7_75t_L g1375 ( 
.A1(n_1288),
.A2(n_1253),
.B(n_1298),
.Y(n_1375)
);

INVxp67_ASAP7_75t_L g1376 ( 
.A(n_1313),
.Y(n_1376)
);

INVx1_ASAP7_75t_L g1377 ( 
.A(n_1297),
.Y(n_1377)
);

INVx2_ASAP7_75t_SL g1378 ( 
.A(n_1328),
.Y(n_1378)
);

AOI21x1_ASAP7_75t_L g1379 ( 
.A1(n_1287),
.A2(n_1302),
.B(n_1298),
.Y(n_1379)
);

HB1xp67_ASAP7_75t_L g1380 ( 
.A(n_1237),
.Y(n_1380)
);

HB1xp67_ASAP7_75t_L g1381 ( 
.A(n_1312),
.Y(n_1381)
);

AND2x4_ASAP7_75t_L g1382 ( 
.A(n_1273),
.B(n_1291),
.Y(n_1382)
);

INVx3_ASAP7_75t_L g1383 ( 
.A(n_1309),
.Y(n_1383)
);

BUFx2_ASAP7_75t_L g1384 ( 
.A(n_1294),
.Y(n_1384)
);

HB1xp67_ASAP7_75t_L g1385 ( 
.A(n_1244),
.Y(n_1385)
);

AOI22xp33_ASAP7_75t_L g1386 ( 
.A1(n_1311),
.A2(n_1331),
.B1(n_1319),
.B2(n_1316),
.Y(n_1386)
);

BUFx4f_ASAP7_75t_L g1387 ( 
.A(n_1220),
.Y(n_1387)
);

HB1xp67_ASAP7_75t_L g1388 ( 
.A(n_1255),
.Y(n_1388)
);

INVx2_ASAP7_75t_L g1389 ( 
.A(n_1326),
.Y(n_1389)
);

AOI22xp33_ASAP7_75t_L g1390 ( 
.A1(n_1316),
.A2(n_1331),
.B1(n_1318),
.B2(n_1243),
.Y(n_1390)
);

AND2x2_ASAP7_75t_L g1391 ( 
.A(n_1240),
.B(n_1238),
.Y(n_1391)
);

INVx2_ASAP7_75t_L g1392 ( 
.A(n_1333),
.Y(n_1392)
);

INVx5_ASAP7_75t_L g1393 ( 
.A(n_1340),
.Y(n_1393)
);

NAND2xp5_ASAP7_75t_L g1394 ( 
.A(n_1314),
.B(n_1321),
.Y(n_1394)
);

AOI22xp33_ASAP7_75t_L g1395 ( 
.A1(n_1243),
.A2(n_1222),
.B1(n_1246),
.B2(n_1314),
.Y(n_1395)
);

AOI21x1_ASAP7_75t_L g1396 ( 
.A1(n_1302),
.A2(n_1307),
.B(n_1278),
.Y(n_1396)
);

INVx2_ASAP7_75t_L g1397 ( 
.A(n_1347),
.Y(n_1397)
);

BUFx2_ASAP7_75t_L g1398 ( 
.A(n_1241),
.Y(n_1398)
);

BUFx2_ASAP7_75t_L g1399 ( 
.A(n_1241),
.Y(n_1399)
);

AOI21x1_ASAP7_75t_L g1400 ( 
.A1(n_1239),
.A2(n_1335),
.B(n_1317),
.Y(n_1400)
);

OA21x2_ASAP7_75t_L g1401 ( 
.A1(n_1266),
.A2(n_1267),
.B(n_1262),
.Y(n_1401)
);

HB1xp67_ASAP7_75t_L g1402 ( 
.A(n_1315),
.Y(n_1402)
);

BUFx2_ASAP7_75t_SL g1403 ( 
.A(n_1340),
.Y(n_1403)
);

INVx2_ASAP7_75t_L g1404 ( 
.A(n_1352),
.Y(n_1404)
);

HB1xp67_ASAP7_75t_L g1405 ( 
.A(n_1327),
.Y(n_1405)
);

INVx1_ASAP7_75t_L g1406 ( 
.A(n_1272),
.Y(n_1406)
);

AOI22xp33_ASAP7_75t_L g1407 ( 
.A1(n_1321),
.A2(n_1357),
.B1(n_1332),
.B2(n_1334),
.Y(n_1407)
);

BUFx3_ASAP7_75t_L g1408 ( 
.A(n_1220),
.Y(n_1408)
);

NOR2xp33_ASAP7_75t_L g1409 ( 
.A(n_1332),
.B(n_1334),
.Y(n_1409)
);

OAI22xp5_ASAP7_75t_L g1410 ( 
.A1(n_1216),
.A2(n_1357),
.B1(n_1353),
.B2(n_1350),
.Y(n_1410)
);

INVx1_ASAP7_75t_L g1411 ( 
.A(n_1249),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_1249),
.Y(n_1412)
);

INVx2_ASAP7_75t_L g1413 ( 
.A(n_1330),
.Y(n_1413)
);

AND2x2_ASAP7_75t_L g1414 ( 
.A(n_1240),
.B(n_1233),
.Y(n_1414)
);

INVx1_ASAP7_75t_L g1415 ( 
.A(n_1250),
.Y(n_1415)
);

INVx1_ASAP7_75t_L g1416 ( 
.A(n_1247),
.Y(n_1416)
);

INVx1_ASAP7_75t_L g1417 ( 
.A(n_1247),
.Y(n_1417)
);

INVx2_ASAP7_75t_L g1418 ( 
.A(n_1341),
.Y(n_1418)
);

INVx1_ASAP7_75t_L g1419 ( 
.A(n_1274),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_1274),
.Y(n_1420)
);

BUFx3_ASAP7_75t_L g1421 ( 
.A(n_1221),
.Y(n_1421)
);

INVx2_ASAP7_75t_L g1422 ( 
.A(n_1342),
.Y(n_1422)
);

INVx1_ASAP7_75t_L g1423 ( 
.A(n_1229),
.Y(n_1423)
);

CKINVDCx11_ASAP7_75t_R g1424 ( 
.A(n_1263),
.Y(n_1424)
);

CKINVDCx5p33_ASAP7_75t_R g1425 ( 
.A(n_1234),
.Y(n_1425)
);

INVx3_ASAP7_75t_L g1426 ( 
.A(n_1273),
.Y(n_1426)
);

INVx2_ASAP7_75t_L g1427 ( 
.A(n_1343),
.Y(n_1427)
);

AOI22xp5_ASAP7_75t_L g1428 ( 
.A1(n_1337),
.A2(n_1350),
.B1(n_1339),
.B2(n_1353),
.Y(n_1428)
);

BUFx3_ASAP7_75t_L g1429 ( 
.A(n_1221),
.Y(n_1429)
);

INVx1_ASAP7_75t_L g1430 ( 
.A(n_1245),
.Y(n_1430)
);

CKINVDCx11_ASAP7_75t_R g1431 ( 
.A(n_1285),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_1233),
.Y(n_1432)
);

INVx2_ASAP7_75t_L g1433 ( 
.A(n_1354),
.Y(n_1433)
);

BUFx6f_ASAP7_75t_L g1434 ( 
.A(n_1340),
.Y(n_1434)
);

BUFx2_ASAP7_75t_L g1435 ( 
.A(n_1235),
.Y(n_1435)
);

AND2x2_ASAP7_75t_L g1436 ( 
.A(n_1227),
.B(n_1217),
.Y(n_1436)
);

OAI22xp33_ASAP7_75t_L g1437 ( 
.A1(n_1337),
.A2(n_1339),
.B1(n_1323),
.B2(n_1217),
.Y(n_1437)
);

AO21x1_ASAP7_75t_SL g1438 ( 
.A1(n_1284),
.A2(n_1260),
.B(n_1310),
.Y(n_1438)
);

HB1xp67_ASAP7_75t_L g1439 ( 
.A(n_1344),
.Y(n_1439)
);

AOI22xp33_ASAP7_75t_L g1440 ( 
.A1(n_1345),
.A2(n_1356),
.B1(n_1346),
.B2(n_1231),
.Y(n_1440)
);

OAI21xp5_ASAP7_75t_L g1441 ( 
.A1(n_1223),
.A2(n_1231),
.B(n_1226),
.Y(n_1441)
);

INVx5_ASAP7_75t_L g1442 ( 
.A(n_1340),
.Y(n_1442)
);

INVx1_ASAP7_75t_L g1443 ( 
.A(n_1303),
.Y(n_1443)
);

OAI21x1_ASAP7_75t_L g1444 ( 
.A1(n_1264),
.A2(n_1265),
.B(n_1248),
.Y(n_1444)
);

AND2x2_ASAP7_75t_L g1445 ( 
.A(n_1226),
.B(n_1271),
.Y(n_1445)
);

CKINVDCx11_ASAP7_75t_R g1446 ( 
.A(n_1279),
.Y(n_1446)
);

AOI22xp5_ASAP7_75t_L g1447 ( 
.A1(n_1254),
.A2(n_1214),
.B1(n_1230),
.B2(n_1242),
.Y(n_1447)
);

INVx2_ASAP7_75t_L g1448 ( 
.A(n_1306),
.Y(n_1448)
);

CKINVDCx5p33_ASAP7_75t_R g1449 ( 
.A(n_1283),
.Y(n_1449)
);

INVx1_ASAP7_75t_L g1450 ( 
.A(n_1275),
.Y(n_1450)
);

OAI21xp5_ASAP7_75t_L g1451 ( 
.A1(n_1275),
.A2(n_1276),
.B(n_1289),
.Y(n_1451)
);

HB1xp67_ASAP7_75t_L g1452 ( 
.A(n_1259),
.Y(n_1452)
);

OAI21x1_ASAP7_75t_L g1453 ( 
.A1(n_1276),
.A2(n_1212),
.B(n_1348),
.Y(n_1453)
);

INVx1_ASAP7_75t_L g1454 ( 
.A(n_1280),
.Y(n_1454)
);

AOI22xp33_ASAP7_75t_SL g1455 ( 
.A1(n_1230),
.A2(n_1242),
.B1(n_1224),
.B2(n_1225),
.Y(n_1455)
);

INVx1_ASAP7_75t_L g1456 ( 
.A(n_1282),
.Y(n_1456)
);

CKINVDCx5p33_ASAP7_75t_R g1457 ( 
.A(n_1355),
.Y(n_1457)
);

INVx2_ASAP7_75t_SL g1458 ( 
.A(n_1336),
.Y(n_1458)
);

INVx1_ASAP7_75t_L g1459 ( 
.A(n_1348),
.Y(n_1459)
);

AOI22xp33_ASAP7_75t_SL g1460 ( 
.A1(n_1224),
.A2(n_1225),
.B1(n_1336),
.B2(n_1212),
.Y(n_1460)
);

INVx2_ASAP7_75t_L g1461 ( 
.A(n_1324),
.Y(n_1461)
);

INVx2_ASAP7_75t_L g1462 ( 
.A(n_1324),
.Y(n_1462)
);

AOI22xp33_ASAP7_75t_L g1463 ( 
.A1(n_1232),
.A2(n_1270),
.B1(n_1268),
.B2(n_1256),
.Y(n_1463)
);

BUFx2_ASAP7_75t_L g1464 ( 
.A(n_1269),
.Y(n_1464)
);

CKINVDCx5p33_ASAP7_75t_R g1465 ( 
.A(n_1261),
.Y(n_1465)
);

OAI22xp33_ASAP7_75t_L g1466 ( 
.A1(n_1322),
.A2(n_1295),
.B1(n_1281),
.B2(n_1286),
.Y(n_1466)
);

INVx2_ASAP7_75t_L g1467 ( 
.A(n_1296),
.Y(n_1467)
);

INVx2_ASAP7_75t_L g1468 ( 
.A(n_1296),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_1296),
.Y(n_1469)
);

INVx2_ASAP7_75t_L g1470 ( 
.A(n_1301),
.Y(n_1470)
);

NAND2xp5_ASAP7_75t_L g1471 ( 
.A(n_1290),
.B(n_1257),
.Y(n_1471)
);

AOI22xp33_ASAP7_75t_L g1472 ( 
.A1(n_1322),
.A2(n_1257),
.B1(n_1277),
.B2(n_1320),
.Y(n_1472)
);

OAI22xp33_ASAP7_75t_L g1473 ( 
.A1(n_1322),
.A2(n_1277),
.B1(n_1320),
.B2(n_1292),
.Y(n_1473)
);

INVxp67_ASAP7_75t_L g1474 ( 
.A(n_1277),
.Y(n_1474)
);

AOI22xp33_ASAP7_75t_L g1475 ( 
.A1(n_1320),
.A2(n_1049),
.B1(n_1052),
.B2(n_951),
.Y(n_1475)
);

INVx2_ASAP7_75t_L g1476 ( 
.A(n_1299),
.Y(n_1476)
);

AND2x2_ASAP7_75t_L g1477 ( 
.A(n_1215),
.B(n_1218),
.Y(n_1477)
);

BUFx3_ASAP7_75t_L g1478 ( 
.A(n_1220),
.Y(n_1478)
);

INVx1_ASAP7_75t_SL g1479 ( 
.A(n_1237),
.Y(n_1479)
);

CKINVDCx20_ASAP7_75t_R g1480 ( 
.A(n_1236),
.Y(n_1480)
);

NOR2xp33_ASAP7_75t_L g1481 ( 
.A(n_1325),
.B(n_1349),
.Y(n_1481)
);

INVxp33_ASAP7_75t_L g1482 ( 
.A(n_1213),
.Y(n_1482)
);

CKINVDCx5p33_ASAP7_75t_R g1483 ( 
.A(n_1251),
.Y(n_1483)
);

INVx1_ASAP7_75t_L g1484 ( 
.A(n_1304),
.Y(n_1484)
);

OA21x2_ASAP7_75t_L g1485 ( 
.A1(n_1266),
.A2(n_1267),
.B(n_1278),
.Y(n_1485)
);

AOI22xp33_ASAP7_75t_L g1486 ( 
.A1(n_1325),
.A2(n_1049),
.B1(n_1052),
.B2(n_951),
.Y(n_1486)
);

AOI22xp33_ASAP7_75t_SL g1487 ( 
.A1(n_1311),
.A2(n_1052),
.B1(n_1049),
.B2(n_1171),
.Y(n_1487)
);

NAND2xp5_ASAP7_75t_L g1488 ( 
.A(n_1325),
.B(n_1171),
.Y(n_1488)
);

INVx1_ASAP7_75t_L g1489 ( 
.A(n_1363),
.Y(n_1489)
);

OAI21xp5_ASAP7_75t_L g1490 ( 
.A1(n_1487),
.A2(n_1486),
.B(n_1362),
.Y(n_1490)
);

AND2x4_ASAP7_75t_SL g1491 ( 
.A(n_1359),
.B(n_1434),
.Y(n_1491)
);

AND2x4_ASAP7_75t_L g1492 ( 
.A(n_1382),
.B(n_1426),
.Y(n_1492)
);

NAND2xp5_ASAP7_75t_L g1493 ( 
.A(n_1410),
.B(n_1437),
.Y(n_1493)
);

AOI21x1_ASAP7_75t_L g1494 ( 
.A1(n_1379),
.A2(n_1396),
.B(n_1400),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_1484),
.Y(n_1495)
);

OAI21x1_ASAP7_75t_L g1496 ( 
.A1(n_1379),
.A2(n_1375),
.B(n_1396),
.Y(n_1496)
);

AND2x2_ASAP7_75t_L g1497 ( 
.A(n_1377),
.B(n_1367),
.Y(n_1497)
);

NAND2xp5_ASAP7_75t_L g1498 ( 
.A(n_1428),
.B(n_1409),
.Y(n_1498)
);

AND2x2_ASAP7_75t_L g1499 ( 
.A(n_1377),
.B(n_1367),
.Y(n_1499)
);

BUFx12f_ASAP7_75t_L g1500 ( 
.A(n_1424),
.Y(n_1500)
);

INVx3_ASAP7_75t_SL g1501 ( 
.A(n_1465),
.Y(n_1501)
);

BUFx2_ASAP7_75t_L g1502 ( 
.A(n_1374),
.Y(n_1502)
);

AND2x2_ASAP7_75t_L g1503 ( 
.A(n_1369),
.B(n_1414),
.Y(n_1503)
);

CKINVDCx11_ASAP7_75t_R g1504 ( 
.A(n_1480),
.Y(n_1504)
);

INVxp33_ASAP7_75t_L g1505 ( 
.A(n_1385),
.Y(n_1505)
);

OA21x2_ASAP7_75t_L g1506 ( 
.A1(n_1444),
.A2(n_1451),
.B(n_1420),
.Y(n_1506)
);

AND2x2_ASAP7_75t_L g1507 ( 
.A(n_1369),
.B(n_1414),
.Y(n_1507)
);

OAI21x1_ASAP7_75t_L g1508 ( 
.A1(n_1375),
.A2(n_1444),
.B(n_1400),
.Y(n_1508)
);

OAI21x1_ASAP7_75t_L g1509 ( 
.A1(n_1453),
.A2(n_1420),
.B(n_1419),
.Y(n_1509)
);

BUFx2_ASAP7_75t_L g1510 ( 
.A(n_1374),
.Y(n_1510)
);

OR2x6_ASAP7_75t_L g1511 ( 
.A(n_1361),
.B(n_1401),
.Y(n_1511)
);

NAND2xp5_ASAP7_75t_L g1512 ( 
.A(n_1428),
.B(n_1436),
.Y(n_1512)
);

HB1xp67_ASAP7_75t_L g1513 ( 
.A(n_1435),
.Y(n_1513)
);

CKINVDCx5p33_ASAP7_75t_R g1514 ( 
.A(n_1364),
.Y(n_1514)
);

HB1xp67_ASAP7_75t_L g1515 ( 
.A(n_1435),
.Y(n_1515)
);

OR2x6_ASAP7_75t_L g1516 ( 
.A(n_1361),
.B(n_1401),
.Y(n_1516)
);

AND2x2_ASAP7_75t_L g1517 ( 
.A(n_1384),
.B(n_1368),
.Y(n_1517)
);

INVxp67_ASAP7_75t_L g1518 ( 
.A(n_1366),
.Y(n_1518)
);

AND2x2_ASAP7_75t_L g1519 ( 
.A(n_1384),
.B(n_1368),
.Y(n_1519)
);

INVx3_ASAP7_75t_L g1520 ( 
.A(n_1382),
.Y(n_1520)
);

BUFx2_ASAP7_75t_L g1521 ( 
.A(n_1443),
.Y(n_1521)
);

INVx3_ASAP7_75t_L g1522 ( 
.A(n_1382),
.Y(n_1522)
);

AND2x4_ASAP7_75t_L g1523 ( 
.A(n_1382),
.B(n_1426),
.Y(n_1523)
);

BUFx2_ASAP7_75t_SL g1524 ( 
.A(n_1393),
.Y(n_1524)
);

HB1xp67_ASAP7_75t_L g1525 ( 
.A(n_1372),
.Y(n_1525)
);

OR2x2_ASAP7_75t_L g1526 ( 
.A(n_1430),
.B(n_1450),
.Y(n_1526)
);

NAND2x1p5_ASAP7_75t_L g1527 ( 
.A(n_1393),
.B(n_1442),
.Y(n_1527)
);

HB1xp67_ASAP7_75t_L g1528 ( 
.A(n_1464),
.Y(n_1528)
);

CKINVDCx14_ASAP7_75t_R g1529 ( 
.A(n_1360),
.Y(n_1529)
);

HB1xp67_ASAP7_75t_L g1530 ( 
.A(n_1464),
.Y(n_1530)
);

AND2x4_ASAP7_75t_L g1531 ( 
.A(n_1426),
.B(n_1383),
.Y(n_1531)
);

OR2x2_ASAP7_75t_L g1532 ( 
.A(n_1430),
.B(n_1450),
.Y(n_1532)
);

AND2x4_ASAP7_75t_L g1533 ( 
.A(n_1426),
.B(n_1383),
.Y(n_1533)
);

OR2x2_ASAP7_75t_L g1534 ( 
.A(n_1406),
.B(n_1398),
.Y(n_1534)
);

BUFx2_ASAP7_75t_L g1535 ( 
.A(n_1443),
.Y(n_1535)
);

NAND2xp5_ASAP7_75t_L g1536 ( 
.A(n_1436),
.B(n_1407),
.Y(n_1536)
);

HB1xp67_ASAP7_75t_L g1537 ( 
.A(n_1445),
.Y(n_1537)
);

HB1xp67_ASAP7_75t_L g1538 ( 
.A(n_1445),
.Y(n_1538)
);

BUFx2_ASAP7_75t_L g1539 ( 
.A(n_1358),
.Y(n_1539)
);

AOI21xp33_ASAP7_75t_L g1540 ( 
.A1(n_1395),
.A2(n_1365),
.B(n_1481),
.Y(n_1540)
);

OA21x2_ASAP7_75t_L g1541 ( 
.A1(n_1448),
.A2(n_1432),
.B(n_1406),
.Y(n_1541)
);

BUFx4f_ASAP7_75t_SL g1542 ( 
.A(n_1479),
.Y(n_1542)
);

INVxp67_ASAP7_75t_L g1543 ( 
.A(n_1381),
.Y(n_1543)
);

INVx1_ASAP7_75t_L g1544 ( 
.A(n_1398),
.Y(n_1544)
);

OR2x2_ASAP7_75t_L g1545 ( 
.A(n_1399),
.B(n_1358),
.Y(n_1545)
);

INVx1_ASAP7_75t_L g1546 ( 
.A(n_1432),
.Y(n_1546)
);

BUFx2_ASAP7_75t_L g1547 ( 
.A(n_1361),
.Y(n_1547)
);

OAI21xp5_ASAP7_75t_L g1548 ( 
.A1(n_1488),
.A2(n_1475),
.B(n_1390),
.Y(n_1548)
);

BUFx3_ASAP7_75t_L g1549 ( 
.A(n_1371),
.Y(n_1549)
);

AOI21x1_ASAP7_75t_L g1550 ( 
.A1(n_1361),
.A2(n_1476),
.B(n_1415),
.Y(n_1550)
);

INVx3_ASAP7_75t_L g1551 ( 
.A(n_1485),
.Y(n_1551)
);

INVx1_ASAP7_75t_L g1552 ( 
.A(n_1401),
.Y(n_1552)
);

INVx1_ASAP7_75t_L g1553 ( 
.A(n_1401),
.Y(n_1553)
);

AND2x2_ASAP7_75t_L g1554 ( 
.A(n_1477),
.B(n_1391),
.Y(n_1554)
);

AO21x2_ASAP7_75t_L g1555 ( 
.A1(n_1441),
.A2(n_1415),
.B(n_1423),
.Y(n_1555)
);

INVx1_ASAP7_75t_L g1556 ( 
.A(n_1389),
.Y(n_1556)
);

INVx1_ASAP7_75t_L g1557 ( 
.A(n_1392),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_1397),
.Y(n_1558)
);

INVx1_ASAP7_75t_L g1559 ( 
.A(n_1404),
.Y(n_1559)
);

INVx1_ASAP7_75t_L g1560 ( 
.A(n_1416),
.Y(n_1560)
);

NOR2xp33_ASAP7_75t_L g1561 ( 
.A(n_1394),
.B(n_1482),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1416),
.Y(n_1562)
);

INVx1_ASAP7_75t_L g1563 ( 
.A(n_1417),
.Y(n_1563)
);

INVx1_ASAP7_75t_L g1564 ( 
.A(n_1417),
.Y(n_1564)
);

AO21x1_ASAP7_75t_SL g1565 ( 
.A1(n_1386),
.A2(n_1447),
.B(n_1411),
.Y(n_1565)
);

AO21x2_ASAP7_75t_L g1566 ( 
.A1(n_1459),
.A2(n_1411),
.B(n_1412),
.Y(n_1566)
);

OAI21x1_ASAP7_75t_L g1567 ( 
.A1(n_1494),
.A2(n_1373),
.B(n_1412),
.Y(n_1567)
);

OR2x2_ASAP7_75t_L g1568 ( 
.A(n_1545),
.B(n_1544),
.Y(n_1568)
);

AO31x2_ASAP7_75t_L g1569 ( 
.A1(n_1552),
.A2(n_1459),
.A3(n_1456),
.B(n_1454),
.Y(n_1569)
);

AND2x2_ASAP7_75t_L g1570 ( 
.A(n_1503),
.B(n_1507),
.Y(n_1570)
);

INVxp67_ASAP7_75t_L g1571 ( 
.A(n_1528),
.Y(n_1571)
);

INVxp67_ASAP7_75t_L g1572 ( 
.A(n_1530),
.Y(n_1572)
);

NAND2xp5_ASAP7_75t_L g1573 ( 
.A(n_1512),
.B(n_1391),
.Y(n_1573)
);

INVxp67_ASAP7_75t_L g1574 ( 
.A(n_1513),
.Y(n_1574)
);

NAND2xp5_ASAP7_75t_L g1575 ( 
.A(n_1526),
.B(n_1477),
.Y(n_1575)
);

INVx1_ASAP7_75t_L g1576 ( 
.A(n_1489),
.Y(n_1576)
);

AND2x2_ASAP7_75t_L g1577 ( 
.A(n_1503),
.B(n_1438),
.Y(n_1577)
);

OR2x2_ASAP7_75t_L g1578 ( 
.A(n_1545),
.B(n_1402),
.Y(n_1578)
);

INVx3_ASAP7_75t_L g1579 ( 
.A(n_1509),
.Y(n_1579)
);

NAND2xp5_ASAP7_75t_L g1580 ( 
.A(n_1526),
.B(n_1405),
.Y(n_1580)
);

OR2x2_ASAP7_75t_L g1581 ( 
.A(n_1544),
.B(n_1439),
.Y(n_1581)
);

NOR2xp33_ASAP7_75t_L g1582 ( 
.A(n_1542),
.B(n_1483),
.Y(n_1582)
);

AND2x4_ASAP7_75t_L g1583 ( 
.A(n_1520),
.B(n_1393),
.Y(n_1583)
);

AND2x2_ASAP7_75t_L g1584 ( 
.A(n_1507),
.B(n_1438),
.Y(n_1584)
);

INVx2_ASAP7_75t_L g1585 ( 
.A(n_1495),
.Y(n_1585)
);

OR2x6_ASAP7_75t_L g1586 ( 
.A(n_1511),
.B(n_1403),
.Y(n_1586)
);

INVx2_ASAP7_75t_L g1587 ( 
.A(n_1495),
.Y(n_1587)
);

OAI21xp5_ASAP7_75t_L g1588 ( 
.A1(n_1490),
.A2(n_1447),
.B(n_1440),
.Y(n_1588)
);

AND2x2_ASAP7_75t_L g1589 ( 
.A(n_1517),
.B(n_1456),
.Y(n_1589)
);

AND2x2_ASAP7_75t_L g1590 ( 
.A(n_1517),
.B(n_1462),
.Y(n_1590)
);

HB1xp67_ASAP7_75t_L g1591 ( 
.A(n_1515),
.Y(n_1591)
);

INVx2_ASAP7_75t_SL g1592 ( 
.A(n_1531),
.Y(n_1592)
);

AND2x2_ASAP7_75t_L g1593 ( 
.A(n_1519),
.B(n_1462),
.Y(n_1593)
);

AND2x2_ASAP7_75t_L g1594 ( 
.A(n_1519),
.B(n_1461),
.Y(n_1594)
);

NAND2xp5_ASAP7_75t_L g1595 ( 
.A(n_1532),
.B(n_1413),
.Y(n_1595)
);

AND2x4_ASAP7_75t_L g1596 ( 
.A(n_1520),
.B(n_1522),
.Y(n_1596)
);

OR2x2_ASAP7_75t_L g1597 ( 
.A(n_1552),
.B(n_1388),
.Y(n_1597)
);

AND2x2_ASAP7_75t_L g1598 ( 
.A(n_1554),
.B(n_1497),
.Y(n_1598)
);

NOR2x1_ASAP7_75t_SL g1599 ( 
.A(n_1511),
.B(n_1403),
.Y(n_1599)
);

INVxp67_ASAP7_75t_SL g1600 ( 
.A(n_1553),
.Y(n_1600)
);

AO21x2_ASAP7_75t_L g1601 ( 
.A1(n_1494),
.A2(n_1473),
.B(n_1466),
.Y(n_1601)
);

NAND2xp5_ASAP7_75t_L g1602 ( 
.A(n_1532),
.B(n_1422),
.Y(n_1602)
);

INVx3_ASAP7_75t_L g1603 ( 
.A(n_1531),
.Y(n_1603)
);

AOI21xp33_ASAP7_75t_SL g1604 ( 
.A1(n_1540),
.A2(n_1483),
.B(n_1425),
.Y(n_1604)
);

INVx1_ASAP7_75t_L g1605 ( 
.A(n_1566),
.Y(n_1605)
);

INVx1_ASAP7_75t_L g1606 ( 
.A(n_1566),
.Y(n_1606)
);

NAND2xp5_ASAP7_75t_L g1607 ( 
.A(n_1498),
.B(n_1433),
.Y(n_1607)
);

INVx3_ASAP7_75t_L g1608 ( 
.A(n_1531),
.Y(n_1608)
);

AND2x2_ASAP7_75t_L g1609 ( 
.A(n_1499),
.B(n_1427),
.Y(n_1609)
);

HB1xp67_ASAP7_75t_L g1610 ( 
.A(n_1502),
.Y(n_1610)
);

CKINVDCx20_ASAP7_75t_R g1611 ( 
.A(n_1504),
.Y(n_1611)
);

AND2x2_ASAP7_75t_L g1612 ( 
.A(n_1537),
.B(n_1427),
.Y(n_1612)
);

AND2x2_ASAP7_75t_L g1613 ( 
.A(n_1538),
.B(n_1433),
.Y(n_1613)
);

BUFx3_ASAP7_75t_L g1614 ( 
.A(n_1549),
.Y(n_1614)
);

INVx2_ASAP7_75t_SL g1615 ( 
.A(n_1531),
.Y(n_1615)
);

AND2x2_ASAP7_75t_L g1616 ( 
.A(n_1547),
.B(n_1522),
.Y(n_1616)
);

INVx1_ASAP7_75t_L g1617 ( 
.A(n_1566),
.Y(n_1617)
);

HB1xp67_ASAP7_75t_L g1618 ( 
.A(n_1502),
.Y(n_1618)
);

AND2x2_ASAP7_75t_L g1619 ( 
.A(n_1547),
.B(n_1418),
.Y(n_1619)
);

HB1xp67_ASAP7_75t_L g1620 ( 
.A(n_1510),
.Y(n_1620)
);

AOI22xp33_ASAP7_75t_L g1621 ( 
.A1(n_1548),
.A2(n_1455),
.B1(n_1478),
.B2(n_1421),
.Y(n_1621)
);

AND2x2_ASAP7_75t_L g1622 ( 
.A(n_1511),
.B(n_1413),
.Y(n_1622)
);

OAI22xp33_ASAP7_75t_L g1623 ( 
.A1(n_1493),
.A2(n_1387),
.B1(n_1408),
.B2(n_1429),
.Y(n_1623)
);

NAND2xp5_ASAP7_75t_L g1624 ( 
.A(n_1573),
.B(n_1525),
.Y(n_1624)
);

NAND3xp33_ASAP7_75t_L g1625 ( 
.A(n_1588),
.B(n_1536),
.C(n_1463),
.Y(n_1625)
);

OAI22xp5_ASAP7_75t_L g1626 ( 
.A1(n_1621),
.A2(n_1501),
.B1(n_1460),
.B2(n_1472),
.Y(n_1626)
);

NAND3xp33_ASAP7_75t_L g1627 ( 
.A(n_1588),
.B(n_1534),
.C(n_1561),
.Y(n_1627)
);

NAND3xp33_ASAP7_75t_L g1628 ( 
.A(n_1604),
.B(n_1534),
.C(n_1543),
.Y(n_1628)
);

NOR2xp33_ASAP7_75t_L g1629 ( 
.A(n_1604),
.B(n_1505),
.Y(n_1629)
);

NAND2xp5_ASAP7_75t_L g1630 ( 
.A(n_1575),
.B(n_1518),
.Y(n_1630)
);

NAND2xp5_ASAP7_75t_L g1631 ( 
.A(n_1580),
.B(n_1539),
.Y(n_1631)
);

NAND2xp5_ASAP7_75t_SL g1632 ( 
.A(n_1623),
.B(n_1492),
.Y(n_1632)
);

OAI21xp5_ASAP7_75t_SL g1633 ( 
.A1(n_1577),
.A2(n_1529),
.B(n_1491),
.Y(n_1633)
);

NAND3xp33_ASAP7_75t_L g1634 ( 
.A(n_1607),
.B(n_1574),
.C(n_1572),
.Y(n_1634)
);

NOR2xp33_ASAP7_75t_L g1635 ( 
.A(n_1578),
.B(n_1501),
.Y(n_1635)
);

NAND2xp5_ASAP7_75t_L g1636 ( 
.A(n_1591),
.B(n_1510),
.Y(n_1636)
);

OAI21xp5_ASAP7_75t_SL g1637 ( 
.A1(n_1577),
.A2(n_1491),
.B(n_1527),
.Y(n_1637)
);

AND2x2_ASAP7_75t_L g1638 ( 
.A(n_1570),
.B(n_1511),
.Y(n_1638)
);

NAND2xp5_ASAP7_75t_L g1639 ( 
.A(n_1571),
.B(n_1521),
.Y(n_1639)
);

NAND2xp5_ASAP7_75t_L g1640 ( 
.A(n_1571),
.B(n_1521),
.Y(n_1640)
);

NAND3xp33_ASAP7_75t_L g1641 ( 
.A(n_1607),
.B(n_1574),
.C(n_1572),
.Y(n_1641)
);

NAND2xp5_ASAP7_75t_L g1642 ( 
.A(n_1578),
.B(n_1535),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1576),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_1585),
.Y(n_1644)
);

NAND4xp25_ASAP7_75t_SL g1645 ( 
.A(n_1584),
.B(n_1471),
.C(n_1469),
.D(n_1563),
.Y(n_1645)
);

NAND2xp5_ASAP7_75t_L g1646 ( 
.A(n_1612),
.B(n_1535),
.Y(n_1646)
);

NAND2xp5_ASAP7_75t_L g1647 ( 
.A(n_1612),
.B(n_1613),
.Y(n_1647)
);

NAND3xp33_ASAP7_75t_L g1648 ( 
.A(n_1597),
.B(n_1380),
.C(n_1376),
.Y(n_1648)
);

AND2x2_ASAP7_75t_L g1649 ( 
.A(n_1570),
.B(n_1511),
.Y(n_1649)
);

NOR2xp33_ASAP7_75t_L g1650 ( 
.A(n_1611),
.B(n_1501),
.Y(n_1650)
);

NAND2xp5_ASAP7_75t_L g1651 ( 
.A(n_1613),
.B(n_1560),
.Y(n_1651)
);

AND2x2_ASAP7_75t_L g1652 ( 
.A(n_1616),
.B(n_1516),
.Y(n_1652)
);

AOI22xp33_ASAP7_75t_L g1653 ( 
.A1(n_1584),
.A2(n_1565),
.B1(n_1523),
.B2(n_1492),
.Y(n_1653)
);

AOI21xp33_ASAP7_75t_L g1654 ( 
.A1(n_1601),
.A2(n_1555),
.B(n_1516),
.Y(n_1654)
);

OA21x2_ASAP7_75t_L g1655 ( 
.A1(n_1605),
.A2(n_1496),
.B(n_1508),
.Y(n_1655)
);

AND2x2_ASAP7_75t_L g1656 ( 
.A(n_1616),
.B(n_1516),
.Y(n_1656)
);

NAND2xp5_ASAP7_75t_L g1657 ( 
.A(n_1598),
.B(n_1562),
.Y(n_1657)
);

AND2x2_ASAP7_75t_L g1658 ( 
.A(n_1603),
.B(n_1516),
.Y(n_1658)
);

OAI21xp5_ASAP7_75t_SL g1659 ( 
.A1(n_1582),
.A2(n_1527),
.B(n_1523),
.Y(n_1659)
);

NAND2xp5_ASAP7_75t_SL g1660 ( 
.A(n_1595),
.B(n_1492),
.Y(n_1660)
);

OAI22xp5_ASAP7_75t_L g1661 ( 
.A1(n_1581),
.A2(n_1387),
.B1(n_1478),
.B2(n_1429),
.Y(n_1661)
);

AND2x2_ASAP7_75t_L g1662 ( 
.A(n_1603),
.B(n_1608),
.Y(n_1662)
);

AND2x2_ASAP7_75t_L g1663 ( 
.A(n_1603),
.B(n_1516),
.Y(n_1663)
);

OAI21xp5_ASAP7_75t_L g1664 ( 
.A1(n_1567),
.A2(n_1469),
.B(n_1533),
.Y(n_1664)
);

NAND3xp33_ASAP7_75t_L g1665 ( 
.A(n_1597),
.B(n_1546),
.C(n_1558),
.Y(n_1665)
);

OA211x2_ASAP7_75t_L g1666 ( 
.A1(n_1595),
.A2(n_1602),
.B(n_1599),
.C(n_1474),
.Y(n_1666)
);

AND2x2_ASAP7_75t_L g1667 ( 
.A(n_1603),
.B(n_1541),
.Y(n_1667)
);

OAI221xp5_ASAP7_75t_SL g1668 ( 
.A1(n_1586),
.A2(n_1452),
.B1(n_1470),
.B2(n_1564),
.C(n_1563),
.Y(n_1668)
);

AND2x2_ASAP7_75t_L g1669 ( 
.A(n_1608),
.B(n_1541),
.Y(n_1669)
);

AND2x2_ASAP7_75t_SL g1670 ( 
.A(n_1583),
.B(n_1506),
.Y(n_1670)
);

AOI22xp33_ASAP7_75t_L g1671 ( 
.A1(n_1622),
.A2(n_1565),
.B1(n_1523),
.B2(n_1492),
.Y(n_1671)
);

NOR2xp33_ASAP7_75t_R g1672 ( 
.A(n_1614),
.B(n_1514),
.Y(n_1672)
);

AND2x4_ASAP7_75t_L g1673 ( 
.A(n_1592),
.B(n_1533),
.Y(n_1673)
);

NAND2xp5_ASAP7_75t_L g1674 ( 
.A(n_1590),
.B(n_1562),
.Y(n_1674)
);

AND2x2_ASAP7_75t_L g1675 ( 
.A(n_1608),
.B(n_1541),
.Y(n_1675)
);

INVxp67_ASAP7_75t_SL g1676 ( 
.A(n_1610),
.Y(n_1676)
);

NAND2xp5_ASAP7_75t_L g1677 ( 
.A(n_1590),
.B(n_1564),
.Y(n_1677)
);

NAND2xp5_ASAP7_75t_L g1678 ( 
.A(n_1593),
.B(n_1594),
.Y(n_1678)
);

AND2x2_ASAP7_75t_L g1679 ( 
.A(n_1608),
.B(n_1541),
.Y(n_1679)
);

NAND4xp25_ASAP7_75t_L g1680 ( 
.A(n_1581),
.B(n_1559),
.C(n_1556),
.D(n_1558),
.Y(n_1680)
);

AOI22xp33_ASAP7_75t_SL g1681 ( 
.A1(n_1601),
.A2(n_1524),
.B1(n_1500),
.B2(n_1555),
.Y(n_1681)
);

HB1xp67_ASAP7_75t_L g1682 ( 
.A(n_1618),
.Y(n_1682)
);

AND2x2_ASAP7_75t_L g1683 ( 
.A(n_1592),
.B(n_1551),
.Y(n_1683)
);

NAND2xp5_ASAP7_75t_L g1684 ( 
.A(n_1593),
.B(n_1556),
.Y(n_1684)
);

AND2x2_ASAP7_75t_L g1685 ( 
.A(n_1592),
.B(n_1551),
.Y(n_1685)
);

AOI22xp5_ASAP7_75t_L g1686 ( 
.A1(n_1622),
.A2(n_1523),
.B1(n_1458),
.B2(n_1555),
.Y(n_1686)
);

NAND3xp33_ASAP7_75t_L g1687 ( 
.A(n_1605),
.B(n_1617),
.C(n_1606),
.Y(n_1687)
);

NAND2xp5_ASAP7_75t_L g1688 ( 
.A(n_1594),
.B(n_1557),
.Y(n_1688)
);

INVx2_ASAP7_75t_L g1689 ( 
.A(n_1667),
.Y(n_1689)
);

NAND2xp5_ASAP7_75t_L g1690 ( 
.A(n_1624),
.B(n_1619),
.Y(n_1690)
);

AND2x4_ASAP7_75t_L g1691 ( 
.A(n_1658),
.B(n_1586),
.Y(n_1691)
);

HB1xp67_ASAP7_75t_L g1692 ( 
.A(n_1682),
.Y(n_1692)
);

AND2x4_ASAP7_75t_L g1693 ( 
.A(n_1658),
.B(n_1586),
.Y(n_1693)
);

AND2x2_ASAP7_75t_L g1694 ( 
.A(n_1638),
.B(n_1615),
.Y(n_1694)
);

AND2x2_ASAP7_75t_L g1695 ( 
.A(n_1638),
.B(n_1615),
.Y(n_1695)
);

INVx2_ASAP7_75t_L g1696 ( 
.A(n_1667),
.Y(n_1696)
);

INVx1_ASAP7_75t_L g1697 ( 
.A(n_1644),
.Y(n_1697)
);

AND2x2_ASAP7_75t_L g1698 ( 
.A(n_1649),
.B(n_1586),
.Y(n_1698)
);

AND2x2_ASAP7_75t_L g1699 ( 
.A(n_1662),
.B(n_1586),
.Y(n_1699)
);

INVx1_ASAP7_75t_L g1700 ( 
.A(n_1644),
.Y(n_1700)
);

OR2x2_ASAP7_75t_L g1701 ( 
.A(n_1642),
.B(n_1568),
.Y(n_1701)
);

AND2x2_ASAP7_75t_L g1702 ( 
.A(n_1652),
.B(n_1596),
.Y(n_1702)
);

NOR2x1_ASAP7_75t_L g1703 ( 
.A(n_1687),
.B(n_1606),
.Y(n_1703)
);

AOI211xp5_ASAP7_75t_L g1704 ( 
.A1(n_1627),
.A2(n_1457),
.B(n_1465),
.C(n_1568),
.Y(n_1704)
);

INVx1_ASAP7_75t_L g1705 ( 
.A(n_1643),
.Y(n_1705)
);

AND2x2_ASAP7_75t_L g1706 ( 
.A(n_1652),
.B(n_1596),
.Y(n_1706)
);

INVx3_ASAP7_75t_L g1707 ( 
.A(n_1669),
.Y(n_1707)
);

INVx1_ASAP7_75t_L g1708 ( 
.A(n_1669),
.Y(n_1708)
);

OR2x2_ASAP7_75t_L g1709 ( 
.A(n_1631),
.B(n_1620),
.Y(n_1709)
);

AND2x4_ASAP7_75t_L g1710 ( 
.A(n_1663),
.B(n_1599),
.Y(n_1710)
);

INVx2_ASAP7_75t_L g1711 ( 
.A(n_1675),
.Y(n_1711)
);

INVxp67_ASAP7_75t_L g1712 ( 
.A(n_1636),
.Y(n_1712)
);

INVx1_ASAP7_75t_L g1713 ( 
.A(n_1675),
.Y(n_1713)
);

INVx1_ASAP7_75t_L g1714 ( 
.A(n_1679),
.Y(n_1714)
);

INVxp67_ASAP7_75t_L g1715 ( 
.A(n_1639),
.Y(n_1715)
);

AND2x2_ASAP7_75t_L g1716 ( 
.A(n_1656),
.B(n_1589),
.Y(n_1716)
);

NOR2xp33_ASAP7_75t_L g1717 ( 
.A(n_1650),
.B(n_1500),
.Y(n_1717)
);

INVx1_ASAP7_75t_L g1718 ( 
.A(n_1679),
.Y(n_1718)
);

INVx6_ASAP7_75t_L g1719 ( 
.A(n_1673),
.Y(n_1719)
);

AND2x2_ASAP7_75t_L g1720 ( 
.A(n_1663),
.B(n_1673),
.Y(n_1720)
);

INVx2_ASAP7_75t_L g1721 ( 
.A(n_1683),
.Y(n_1721)
);

AND2x4_ASAP7_75t_L g1722 ( 
.A(n_1683),
.B(n_1583),
.Y(n_1722)
);

INVx1_ASAP7_75t_L g1723 ( 
.A(n_1665),
.Y(n_1723)
);

BUFx3_ASAP7_75t_L g1724 ( 
.A(n_1673),
.Y(n_1724)
);

AND2x2_ASAP7_75t_L g1725 ( 
.A(n_1670),
.B(n_1600),
.Y(n_1725)
);

OR2x2_ASAP7_75t_L g1726 ( 
.A(n_1646),
.B(n_1676),
.Y(n_1726)
);

NAND2x1_ASAP7_75t_L g1727 ( 
.A(n_1686),
.B(n_1585),
.Y(n_1727)
);

AND2x2_ASAP7_75t_L g1728 ( 
.A(n_1670),
.B(n_1600),
.Y(n_1728)
);

INVx1_ASAP7_75t_L g1729 ( 
.A(n_1685),
.Y(n_1729)
);

OR2x2_ASAP7_75t_L g1730 ( 
.A(n_1640),
.B(n_1647),
.Y(n_1730)
);

INVx1_ASAP7_75t_L g1731 ( 
.A(n_1651),
.Y(n_1731)
);

AND2x2_ASAP7_75t_L g1732 ( 
.A(n_1678),
.B(n_1587),
.Y(n_1732)
);

INVx2_ASAP7_75t_L g1733 ( 
.A(n_1655),
.Y(n_1733)
);

INVx1_ASAP7_75t_L g1734 ( 
.A(n_1684),
.Y(n_1734)
);

INVx1_ASAP7_75t_L g1735 ( 
.A(n_1688),
.Y(n_1735)
);

NOR2xp33_ASAP7_75t_L g1736 ( 
.A(n_1630),
.B(n_1370),
.Y(n_1736)
);

AND2x2_ASAP7_75t_L g1737 ( 
.A(n_1660),
.B(n_1587),
.Y(n_1737)
);

OR2x2_ASAP7_75t_L g1738 ( 
.A(n_1657),
.B(n_1617),
.Y(n_1738)
);

INVx2_ASAP7_75t_L g1739 ( 
.A(n_1689),
.Y(n_1739)
);

NOR2xp33_ASAP7_75t_L g1740 ( 
.A(n_1717),
.B(n_1736),
.Y(n_1740)
);

INVx1_ASAP7_75t_L g1741 ( 
.A(n_1697),
.Y(n_1741)
);

NOR2xp33_ASAP7_75t_SL g1742 ( 
.A(n_1703),
.B(n_1668),
.Y(n_1742)
);

INVx1_ASAP7_75t_L g1743 ( 
.A(n_1697),
.Y(n_1743)
);

NOR2x1_ASAP7_75t_L g1744 ( 
.A(n_1703),
.B(n_1628),
.Y(n_1744)
);

BUFx2_ASAP7_75t_L g1745 ( 
.A(n_1724),
.Y(n_1745)
);

INVx1_ASAP7_75t_SL g1746 ( 
.A(n_1692),
.Y(n_1746)
);

NAND2xp5_ASAP7_75t_L g1747 ( 
.A(n_1723),
.B(n_1634),
.Y(n_1747)
);

AND2x2_ASAP7_75t_L g1748 ( 
.A(n_1722),
.B(n_1681),
.Y(n_1748)
);

AND2x2_ASAP7_75t_L g1749 ( 
.A(n_1722),
.B(n_1635),
.Y(n_1749)
);

AND2x2_ASAP7_75t_L g1750 ( 
.A(n_1722),
.B(n_1659),
.Y(n_1750)
);

OR2x2_ASAP7_75t_L g1751 ( 
.A(n_1723),
.B(n_1641),
.Y(n_1751)
);

INVx1_ASAP7_75t_L g1752 ( 
.A(n_1700),
.Y(n_1752)
);

NAND2xp5_ASAP7_75t_L g1753 ( 
.A(n_1715),
.B(n_1660),
.Y(n_1753)
);

NAND2xp5_ASAP7_75t_L g1754 ( 
.A(n_1712),
.B(n_1648),
.Y(n_1754)
);

NAND2x1p5_ASAP7_75t_L g1755 ( 
.A(n_1727),
.B(n_1550),
.Y(n_1755)
);

NOR2xp33_ASAP7_75t_SL g1756 ( 
.A(n_1725),
.B(n_1633),
.Y(n_1756)
);

AND2x2_ASAP7_75t_L g1757 ( 
.A(n_1722),
.B(n_1637),
.Y(n_1757)
);

AND2x2_ASAP7_75t_L g1758 ( 
.A(n_1720),
.B(n_1664),
.Y(n_1758)
);

NOR2x1_ASAP7_75t_R g1759 ( 
.A(n_1704),
.B(n_1431),
.Y(n_1759)
);

AND2x4_ASAP7_75t_L g1760 ( 
.A(n_1691),
.B(n_1579),
.Y(n_1760)
);

AND2x2_ASAP7_75t_L g1761 ( 
.A(n_1720),
.B(n_1654),
.Y(n_1761)
);

NOR2xp33_ASAP7_75t_SL g1762 ( 
.A(n_1725),
.B(n_1625),
.Y(n_1762)
);

NOR3xp33_ASAP7_75t_L g1763 ( 
.A(n_1704),
.B(n_1629),
.C(n_1626),
.Y(n_1763)
);

INVx1_ASAP7_75t_L g1764 ( 
.A(n_1700),
.Y(n_1764)
);

NAND2xp5_ASAP7_75t_L g1765 ( 
.A(n_1731),
.B(n_1674),
.Y(n_1765)
);

NAND2xp5_ASAP7_75t_L g1766 ( 
.A(n_1731),
.B(n_1677),
.Y(n_1766)
);

INVx1_ASAP7_75t_L g1767 ( 
.A(n_1705),
.Y(n_1767)
);

INVx2_ASAP7_75t_SL g1768 ( 
.A(n_1719),
.Y(n_1768)
);

AND2x2_ASAP7_75t_L g1769 ( 
.A(n_1699),
.B(n_1671),
.Y(n_1769)
);

OR2x2_ASAP7_75t_L g1770 ( 
.A(n_1727),
.B(n_1680),
.Y(n_1770)
);

INVx1_ASAP7_75t_L g1771 ( 
.A(n_1705),
.Y(n_1771)
);

AND2x2_ASAP7_75t_L g1772 ( 
.A(n_1699),
.B(n_1632),
.Y(n_1772)
);

INVxp67_ASAP7_75t_L g1773 ( 
.A(n_1726),
.Y(n_1773)
);

INVx1_ASAP7_75t_L g1774 ( 
.A(n_1737),
.Y(n_1774)
);

NAND2xp5_ASAP7_75t_L g1775 ( 
.A(n_1734),
.B(n_1609),
.Y(n_1775)
);

INVx2_ASAP7_75t_L g1776 ( 
.A(n_1689),
.Y(n_1776)
);

OR2x2_ASAP7_75t_L g1777 ( 
.A(n_1708),
.B(n_1569),
.Y(n_1777)
);

AND2x4_ASAP7_75t_L g1778 ( 
.A(n_1691),
.B(n_1579),
.Y(n_1778)
);

INVx1_ASAP7_75t_L g1779 ( 
.A(n_1737),
.Y(n_1779)
);

NOR2xp33_ASAP7_75t_L g1780 ( 
.A(n_1730),
.B(n_1457),
.Y(n_1780)
);

AND2x2_ASAP7_75t_L g1781 ( 
.A(n_1724),
.B(n_1632),
.Y(n_1781)
);

AND2x2_ASAP7_75t_L g1782 ( 
.A(n_1724),
.B(n_1583),
.Y(n_1782)
);

INVxp33_ASAP7_75t_L g1783 ( 
.A(n_1690),
.Y(n_1783)
);

INVx2_ASAP7_75t_L g1784 ( 
.A(n_1689),
.Y(n_1784)
);

INVx1_ASAP7_75t_L g1785 ( 
.A(n_1767),
.Y(n_1785)
);

INVx2_ASAP7_75t_L g1786 ( 
.A(n_1739),
.Y(n_1786)
);

AND2x2_ASAP7_75t_L g1787 ( 
.A(n_1748),
.B(n_1710),
.Y(n_1787)
);

AND2x2_ASAP7_75t_L g1788 ( 
.A(n_1748),
.B(n_1710),
.Y(n_1788)
);

INVx1_ASAP7_75t_L g1789 ( 
.A(n_1767),
.Y(n_1789)
);

AND2x2_ASAP7_75t_L g1790 ( 
.A(n_1757),
.B(n_1750),
.Y(n_1790)
);

AND2x2_ASAP7_75t_L g1791 ( 
.A(n_1757),
.B(n_1710),
.Y(n_1791)
);

INVx1_ASAP7_75t_L g1792 ( 
.A(n_1771),
.Y(n_1792)
);

AND2x2_ASAP7_75t_L g1793 ( 
.A(n_1750),
.B(n_1710),
.Y(n_1793)
);

INVx2_ASAP7_75t_L g1794 ( 
.A(n_1739),
.Y(n_1794)
);

HB1xp67_ASAP7_75t_L g1795 ( 
.A(n_1746),
.Y(n_1795)
);

NAND2xp5_ASAP7_75t_L g1796 ( 
.A(n_1747),
.B(n_1734),
.Y(n_1796)
);

OAI22xp5_ASAP7_75t_L g1797 ( 
.A1(n_1763),
.A2(n_1653),
.B1(n_1719),
.B2(n_1666),
.Y(n_1797)
);

NAND2xp5_ASAP7_75t_L g1798 ( 
.A(n_1751),
.B(n_1735),
.Y(n_1798)
);

HB1xp67_ASAP7_75t_L g1799 ( 
.A(n_1773),
.Y(n_1799)
);

AOI211xp5_ASAP7_75t_SL g1800 ( 
.A1(n_1742),
.A2(n_1661),
.B(n_1728),
.C(n_1693),
.Y(n_1800)
);

NOR2x1p5_ASAP7_75t_L g1801 ( 
.A(n_1754),
.B(n_1691),
.Y(n_1801)
);

OAI21xp33_ASAP7_75t_L g1802 ( 
.A1(n_1742),
.A2(n_1728),
.B(n_1645),
.Y(n_1802)
);

OAI21xp33_ASAP7_75t_L g1803 ( 
.A1(n_1762),
.A2(n_1726),
.B(n_1735),
.Y(n_1803)
);

OR2x2_ASAP7_75t_L g1804 ( 
.A(n_1751),
.B(n_1738),
.Y(n_1804)
);

INVx1_ASAP7_75t_L g1805 ( 
.A(n_1771),
.Y(n_1805)
);

INVx1_ASAP7_75t_L g1806 ( 
.A(n_1741),
.Y(n_1806)
);

OR2x2_ASAP7_75t_L g1807 ( 
.A(n_1774),
.B(n_1738),
.Y(n_1807)
);

INVx1_ASAP7_75t_L g1808 ( 
.A(n_1741),
.Y(n_1808)
);

AOI211xp5_ASAP7_75t_SL g1809 ( 
.A1(n_1762),
.A2(n_1691),
.B(n_1693),
.C(n_1698),
.Y(n_1809)
);

OR2x2_ASAP7_75t_L g1810 ( 
.A(n_1774),
.B(n_1696),
.Y(n_1810)
);

INVx1_ASAP7_75t_L g1811 ( 
.A(n_1743),
.Y(n_1811)
);

INVx2_ASAP7_75t_L g1812 ( 
.A(n_1776),
.Y(n_1812)
);

NAND2xp5_ASAP7_75t_L g1813 ( 
.A(n_1753),
.B(n_1716),
.Y(n_1813)
);

HB1xp67_ASAP7_75t_L g1814 ( 
.A(n_1744),
.Y(n_1814)
);

INVx1_ASAP7_75t_L g1815 ( 
.A(n_1743),
.Y(n_1815)
);

OR2x2_ASAP7_75t_L g1816 ( 
.A(n_1779),
.B(n_1696),
.Y(n_1816)
);

INVx1_ASAP7_75t_L g1817 ( 
.A(n_1752),
.Y(n_1817)
);

INVxp67_ASAP7_75t_SL g1818 ( 
.A(n_1744),
.Y(n_1818)
);

NAND2x2_ASAP7_75t_L g1819 ( 
.A(n_1759),
.B(n_1614),
.Y(n_1819)
);

INVx2_ASAP7_75t_L g1820 ( 
.A(n_1776),
.Y(n_1820)
);

OR2x2_ASAP7_75t_L g1821 ( 
.A(n_1779),
.B(n_1696),
.Y(n_1821)
);

AOI211xp5_ASAP7_75t_L g1822 ( 
.A1(n_1759),
.A2(n_1672),
.B(n_1698),
.C(n_1693),
.Y(n_1822)
);

NAND2xp5_ASAP7_75t_L g1823 ( 
.A(n_1783),
.B(n_1716),
.Y(n_1823)
);

INVx1_ASAP7_75t_L g1824 ( 
.A(n_1752),
.Y(n_1824)
);

INVx1_ASAP7_75t_L g1825 ( 
.A(n_1764),
.Y(n_1825)
);

INVx1_ASAP7_75t_L g1826 ( 
.A(n_1764),
.Y(n_1826)
);

OAI21xp33_ASAP7_75t_SL g1827 ( 
.A1(n_1772),
.A2(n_1706),
.B(n_1702),
.Y(n_1827)
);

NAND2xp5_ASAP7_75t_L g1828 ( 
.A(n_1765),
.B(n_1732),
.Y(n_1828)
);

CKINVDCx16_ASAP7_75t_R g1829 ( 
.A(n_1756),
.Y(n_1829)
);

INVx1_ASAP7_75t_L g1830 ( 
.A(n_1777),
.Y(n_1830)
);

INVx1_ASAP7_75t_L g1831 ( 
.A(n_1785),
.Y(n_1831)
);

INVx1_ASAP7_75t_SL g1832 ( 
.A(n_1829),
.Y(n_1832)
);

INVx1_ASAP7_75t_L g1833 ( 
.A(n_1785),
.Y(n_1833)
);

HB1xp67_ASAP7_75t_L g1834 ( 
.A(n_1795),
.Y(n_1834)
);

INVx1_ASAP7_75t_L g1835 ( 
.A(n_1808),
.Y(n_1835)
);

HB1xp67_ASAP7_75t_L g1836 ( 
.A(n_1814),
.Y(n_1836)
);

NOR2x1_ASAP7_75t_L g1837 ( 
.A(n_1801),
.B(n_1770),
.Y(n_1837)
);

NAND2xp5_ASAP7_75t_L g1838 ( 
.A(n_1799),
.B(n_1772),
.Y(n_1838)
);

AOI21xp5_ASAP7_75t_L g1839 ( 
.A1(n_1818),
.A2(n_1802),
.B(n_1800),
.Y(n_1839)
);

INVx1_ASAP7_75t_L g1840 ( 
.A(n_1808),
.Y(n_1840)
);

INVx1_ASAP7_75t_L g1841 ( 
.A(n_1811),
.Y(n_1841)
);

CKINVDCx6p67_ASAP7_75t_R g1842 ( 
.A(n_1819),
.Y(n_1842)
);

INVx1_ASAP7_75t_L g1843 ( 
.A(n_1811),
.Y(n_1843)
);

INVx2_ASAP7_75t_L g1844 ( 
.A(n_1786),
.Y(n_1844)
);

INVx1_ASAP7_75t_L g1845 ( 
.A(n_1815),
.Y(n_1845)
);

AOI21xp5_ASAP7_75t_L g1846 ( 
.A1(n_1822),
.A2(n_1770),
.B(n_1740),
.Y(n_1846)
);

NOR2x1_ASAP7_75t_L g1847 ( 
.A(n_1797),
.B(n_1745),
.Y(n_1847)
);

INVx2_ASAP7_75t_L g1848 ( 
.A(n_1786),
.Y(n_1848)
);

NAND2xp5_ASAP7_75t_L g1849 ( 
.A(n_1796),
.B(n_1798),
.Y(n_1849)
);

INVx1_ASAP7_75t_L g1850 ( 
.A(n_1815),
.Y(n_1850)
);

OR2x2_ASAP7_75t_L g1851 ( 
.A(n_1804),
.B(n_1784),
.Y(n_1851)
);

BUFx3_ASAP7_75t_L g1852 ( 
.A(n_1790),
.Y(n_1852)
);

INVx1_ASAP7_75t_L g1853 ( 
.A(n_1817),
.Y(n_1853)
);

NAND2xp5_ASAP7_75t_L g1854 ( 
.A(n_1790),
.B(n_1803),
.Y(n_1854)
);

AND2x2_ASAP7_75t_L g1855 ( 
.A(n_1809),
.B(n_1781),
.Y(n_1855)
);

OAI22xp5_ASAP7_75t_L g1856 ( 
.A1(n_1819),
.A2(n_1781),
.B1(n_1755),
.B2(n_1719),
.Y(n_1856)
);

AND2x4_ASAP7_75t_L g1857 ( 
.A(n_1787),
.B(n_1745),
.Y(n_1857)
);

AND2x2_ASAP7_75t_L g1858 ( 
.A(n_1787),
.B(n_1758),
.Y(n_1858)
);

AND2x2_ASAP7_75t_L g1859 ( 
.A(n_1788),
.B(n_1758),
.Y(n_1859)
);

INVx1_ASAP7_75t_L g1860 ( 
.A(n_1817),
.Y(n_1860)
);

NAND2xp5_ASAP7_75t_L g1861 ( 
.A(n_1813),
.B(n_1780),
.Y(n_1861)
);

INVxp67_ASAP7_75t_L g1862 ( 
.A(n_1804),
.Y(n_1862)
);

OR2x2_ASAP7_75t_L g1863 ( 
.A(n_1807),
.B(n_1784),
.Y(n_1863)
);

NAND2xp5_ASAP7_75t_L g1864 ( 
.A(n_1823),
.B(n_1769),
.Y(n_1864)
);

AOI21xp33_ASAP7_75t_SL g1865 ( 
.A1(n_1788),
.A2(n_1768),
.B(n_1755),
.Y(n_1865)
);

INVx2_ASAP7_75t_L g1866 ( 
.A(n_1794),
.Y(n_1866)
);

OR2x2_ASAP7_75t_L g1867 ( 
.A(n_1807),
.B(n_1777),
.Y(n_1867)
);

NAND2xp5_ASAP7_75t_L g1868 ( 
.A(n_1828),
.B(n_1769),
.Y(n_1868)
);

INVx1_ASAP7_75t_L g1869 ( 
.A(n_1824),
.Y(n_1869)
);

AOI22xp5_ASAP7_75t_L g1870 ( 
.A1(n_1847),
.A2(n_1791),
.B1(n_1793),
.B2(n_1827),
.Y(n_1870)
);

NAND2xp5_ASAP7_75t_L g1871 ( 
.A(n_1834),
.B(n_1791),
.Y(n_1871)
);

AOI21xp33_ASAP7_75t_SL g1872 ( 
.A1(n_1854),
.A2(n_1425),
.B(n_1755),
.Y(n_1872)
);

AO22x1_ASAP7_75t_L g1873 ( 
.A1(n_1832),
.A2(n_1768),
.B1(n_1793),
.B2(n_1792),
.Y(n_1873)
);

OAI221xp5_ASAP7_75t_L g1874 ( 
.A1(n_1839),
.A2(n_1805),
.B1(n_1789),
.B2(n_1825),
.C(n_1806),
.Y(n_1874)
);

AOI221xp5_ASAP7_75t_L g1875 ( 
.A1(n_1855),
.A2(n_1846),
.B1(n_1862),
.B2(n_1836),
.C(n_1852),
.Y(n_1875)
);

NAND2xp5_ASAP7_75t_L g1876 ( 
.A(n_1852),
.B(n_1761),
.Y(n_1876)
);

NAND2xp5_ASAP7_75t_L g1877 ( 
.A(n_1838),
.B(n_1761),
.Y(n_1877)
);

NAND2xp5_ASAP7_75t_L g1878 ( 
.A(n_1861),
.B(n_1855),
.Y(n_1878)
);

NOR2xp67_ASAP7_75t_L g1879 ( 
.A(n_1865),
.B(n_1826),
.Y(n_1879)
);

INVx1_ASAP7_75t_L g1880 ( 
.A(n_1835),
.Y(n_1880)
);

OAI222xp33_ASAP7_75t_L g1881 ( 
.A1(n_1837),
.A2(n_1821),
.B1(n_1810),
.B2(n_1816),
.C1(n_1824),
.C2(n_1830),
.Y(n_1881)
);

NAND2xp5_ASAP7_75t_L g1882 ( 
.A(n_1864),
.B(n_1749),
.Y(n_1882)
);

INVx1_ASAP7_75t_L g1883 ( 
.A(n_1835),
.Y(n_1883)
);

OAI22xp5_ASAP7_75t_L g1884 ( 
.A1(n_1842),
.A2(n_1719),
.B1(n_1693),
.B2(n_1749),
.Y(n_1884)
);

AOI211xp5_ASAP7_75t_L g1885 ( 
.A1(n_1856),
.A2(n_1672),
.B(n_1830),
.C(n_1812),
.Y(n_1885)
);

NAND2xp5_ASAP7_75t_SL g1886 ( 
.A(n_1857),
.B(n_1794),
.Y(n_1886)
);

OAI221xp5_ASAP7_75t_L g1887 ( 
.A1(n_1849),
.A2(n_1821),
.B1(n_1810),
.B2(n_1816),
.C(n_1812),
.Y(n_1887)
);

OAI22xp5_ASAP7_75t_L g1888 ( 
.A1(n_1842),
.A2(n_1719),
.B1(n_1778),
.B2(n_1760),
.Y(n_1888)
);

INVx1_ASAP7_75t_L g1889 ( 
.A(n_1840),
.Y(n_1889)
);

INVx1_ASAP7_75t_L g1890 ( 
.A(n_1840),
.Y(n_1890)
);

OAI22xp5_ASAP7_75t_L g1891 ( 
.A1(n_1857),
.A2(n_1778),
.B1(n_1760),
.B2(n_1782),
.Y(n_1891)
);

INVx1_ASAP7_75t_L g1892 ( 
.A(n_1841),
.Y(n_1892)
);

AOI22xp5_ASAP7_75t_L g1893 ( 
.A1(n_1857),
.A2(n_1868),
.B1(n_1859),
.B2(n_1858),
.Y(n_1893)
);

INVx1_ASAP7_75t_L g1894 ( 
.A(n_1841),
.Y(n_1894)
);

INVx1_ASAP7_75t_L g1895 ( 
.A(n_1850),
.Y(n_1895)
);

AND2x2_ASAP7_75t_L g1896 ( 
.A(n_1858),
.B(n_1760),
.Y(n_1896)
);

INVx1_ASAP7_75t_SL g1897 ( 
.A(n_1859),
.Y(n_1897)
);

NOR2x1_ASAP7_75t_L g1898 ( 
.A(n_1850),
.B(n_1820),
.Y(n_1898)
);

INVx1_ASAP7_75t_L g1899 ( 
.A(n_1898),
.Y(n_1899)
);

HB1xp67_ASAP7_75t_L g1900 ( 
.A(n_1897),
.Y(n_1900)
);

INVx3_ASAP7_75t_SL g1901 ( 
.A(n_1886),
.Y(n_1901)
);

NOR2xp33_ASAP7_75t_SL g1902 ( 
.A(n_1874),
.B(n_1449),
.Y(n_1902)
);

INVxp67_ASAP7_75t_SL g1903 ( 
.A(n_1886),
.Y(n_1903)
);

INVxp67_ASAP7_75t_SL g1904 ( 
.A(n_1873),
.Y(n_1904)
);

AND2x2_ASAP7_75t_L g1905 ( 
.A(n_1893),
.B(n_1844),
.Y(n_1905)
);

INVx1_ASAP7_75t_L g1906 ( 
.A(n_1880),
.Y(n_1906)
);

AND2x2_ASAP7_75t_L g1907 ( 
.A(n_1870),
.B(n_1844),
.Y(n_1907)
);

NAND2xp5_ASAP7_75t_L g1908 ( 
.A(n_1875),
.B(n_1831),
.Y(n_1908)
);

NAND2xp5_ASAP7_75t_L g1909 ( 
.A(n_1878),
.B(n_1833),
.Y(n_1909)
);

NAND2xp5_ASAP7_75t_L g1910 ( 
.A(n_1871),
.B(n_1882),
.Y(n_1910)
);

OR2x2_ASAP7_75t_L g1911 ( 
.A(n_1877),
.B(n_1876),
.Y(n_1911)
);

INVx2_ASAP7_75t_L g1912 ( 
.A(n_1896),
.Y(n_1912)
);

INVx1_ASAP7_75t_SL g1913 ( 
.A(n_1896),
.Y(n_1913)
);

OR2x2_ASAP7_75t_L g1914 ( 
.A(n_1887),
.B(n_1851),
.Y(n_1914)
);

INVx1_ASAP7_75t_L g1915 ( 
.A(n_1883),
.Y(n_1915)
);

INVxp67_ASAP7_75t_L g1916 ( 
.A(n_1879),
.Y(n_1916)
);

NAND2xp5_ASAP7_75t_L g1917 ( 
.A(n_1889),
.B(n_1843),
.Y(n_1917)
);

AND2x2_ASAP7_75t_L g1918 ( 
.A(n_1885),
.B(n_1848),
.Y(n_1918)
);

NAND2xp5_ASAP7_75t_L g1919 ( 
.A(n_1890),
.B(n_1845),
.Y(n_1919)
);

OA22x2_ASAP7_75t_L g1920 ( 
.A1(n_1892),
.A2(n_1860),
.B1(n_1853),
.B2(n_1869),
.Y(n_1920)
);

INVx2_ASAP7_75t_L g1921 ( 
.A(n_1894),
.Y(n_1921)
);

AOI22xp5_ASAP7_75t_L g1922 ( 
.A1(n_1904),
.A2(n_1884),
.B1(n_1888),
.B2(n_1891),
.Y(n_1922)
);

NAND3xp33_ASAP7_75t_L g1923 ( 
.A(n_1908),
.B(n_1872),
.C(n_1895),
.Y(n_1923)
);

AOI321xp33_ASAP7_75t_L g1924 ( 
.A1(n_1903),
.A2(n_1881),
.A3(n_1869),
.B1(n_1848),
.B2(n_1866),
.C(n_1851),
.Y(n_1924)
);

OAI221xp5_ASAP7_75t_L g1925 ( 
.A1(n_1902),
.A2(n_1901),
.B1(n_1916),
.B2(n_1914),
.C(n_1900),
.Y(n_1925)
);

HB1xp67_ASAP7_75t_L g1926 ( 
.A(n_1899),
.Y(n_1926)
);

NAND2xp5_ASAP7_75t_L g1927 ( 
.A(n_1901),
.B(n_1866),
.Y(n_1927)
);

AOI222xp33_ASAP7_75t_L g1928 ( 
.A1(n_1905),
.A2(n_1881),
.B1(n_1820),
.B2(n_1733),
.C1(n_1446),
.C2(n_1766),
.Y(n_1928)
);

AOI32xp33_ASAP7_75t_L g1929 ( 
.A1(n_1907),
.A2(n_1863),
.A3(n_1867),
.B1(n_1782),
.B2(n_1778),
.Y(n_1929)
);

INVx1_ASAP7_75t_L g1930 ( 
.A(n_1920),
.Y(n_1930)
);

INVx1_ASAP7_75t_L g1931 ( 
.A(n_1920),
.Y(n_1931)
);

AOI221xp5_ASAP7_75t_L g1932 ( 
.A1(n_1905),
.A2(n_1863),
.B1(n_1867),
.B2(n_1733),
.C(n_1760),
.Y(n_1932)
);

AOI21xp5_ASAP7_75t_L g1933 ( 
.A1(n_1914),
.A2(n_1778),
.B(n_1775),
.Y(n_1933)
);

OAI221xp5_ASAP7_75t_L g1934 ( 
.A1(n_1910),
.A2(n_1709),
.B1(n_1730),
.B2(n_1449),
.C(n_1707),
.Y(n_1934)
);

AOI22xp5_ASAP7_75t_L g1935 ( 
.A1(n_1913),
.A2(n_1614),
.B1(n_1601),
.B2(n_1707),
.Y(n_1935)
);

NOR3xp33_ASAP7_75t_L g1936 ( 
.A(n_1918),
.B(n_1458),
.C(n_1467),
.Y(n_1936)
);

OR2x2_ASAP7_75t_L g1937 ( 
.A(n_1927),
.B(n_1911),
.Y(n_1937)
);

HB1xp67_ASAP7_75t_L g1938 ( 
.A(n_1926),
.Y(n_1938)
);

NOR2xp33_ASAP7_75t_L g1939 ( 
.A(n_1925),
.B(n_1911),
.Y(n_1939)
);

AOI22xp5_ASAP7_75t_L g1940 ( 
.A1(n_1922),
.A2(n_1912),
.B1(n_1907),
.B2(n_1918),
.Y(n_1940)
);

NOR2x1_ASAP7_75t_L g1941 ( 
.A(n_1930),
.B(n_1899),
.Y(n_1941)
);

NOR3xp33_ASAP7_75t_L g1942 ( 
.A(n_1923),
.B(n_1909),
.C(n_1915),
.Y(n_1942)
);

NOR2x1_ASAP7_75t_L g1943 ( 
.A(n_1931),
.B(n_1921),
.Y(n_1943)
);

NOR2xp33_ASAP7_75t_L g1944 ( 
.A(n_1934),
.B(n_1912),
.Y(n_1944)
);

AOI211xp5_ASAP7_75t_L g1945 ( 
.A1(n_1924),
.A2(n_1919),
.B(n_1917),
.C(n_1906),
.Y(n_1945)
);

NAND3xp33_ASAP7_75t_L g1946 ( 
.A(n_1928),
.B(n_1921),
.C(n_1906),
.Y(n_1946)
);

NOR2xp33_ASAP7_75t_L g1947 ( 
.A(n_1933),
.B(n_1920),
.Y(n_1947)
);

NOR2xp33_ASAP7_75t_L g1948 ( 
.A(n_1937),
.B(n_1936),
.Y(n_1948)
);

NOR2xp33_ASAP7_75t_SL g1949 ( 
.A(n_1938),
.B(n_1929),
.Y(n_1949)
);

NOR2x1_ASAP7_75t_L g1950 ( 
.A(n_1943),
.B(n_1932),
.Y(n_1950)
);

NAND4xp25_ASAP7_75t_SL g1951 ( 
.A(n_1945),
.B(n_1935),
.C(n_1709),
.D(n_1718),
.Y(n_1951)
);

NAND3xp33_ASAP7_75t_L g1952 ( 
.A(n_1942),
.B(n_1468),
.C(n_1467),
.Y(n_1952)
);

NAND4xp25_ASAP7_75t_L g1953 ( 
.A(n_1940),
.B(n_1421),
.C(n_1408),
.D(n_1429),
.Y(n_1953)
);

AOI221xp5_ASAP7_75t_L g1954 ( 
.A1(n_1947),
.A2(n_1733),
.B1(n_1707),
.B2(n_1714),
.C(n_1713),
.Y(n_1954)
);

INVx1_ASAP7_75t_L g1955 ( 
.A(n_1950),
.Y(n_1955)
);

INVx2_ASAP7_75t_L g1956 ( 
.A(n_1952),
.Y(n_1956)
);

AOI22xp5_ASAP7_75t_L g1957 ( 
.A1(n_1949),
.A2(n_1939),
.B1(n_1944),
.B2(n_1946),
.Y(n_1957)
);

INVx1_ASAP7_75t_L g1958 ( 
.A(n_1948),
.Y(n_1958)
);

AOI22xp5_ASAP7_75t_L g1959 ( 
.A1(n_1951),
.A2(n_1941),
.B1(n_1707),
.B2(n_1713),
.Y(n_1959)
);

INVx1_ASAP7_75t_L g1960 ( 
.A(n_1953),
.Y(n_1960)
);

INVx1_ASAP7_75t_L g1961 ( 
.A(n_1954),
.Y(n_1961)
);

NAND3xp33_ASAP7_75t_SL g1962 ( 
.A(n_1955),
.B(n_1957),
.C(n_1958),
.Y(n_1962)
);

AND2x4_ASAP7_75t_L g1963 ( 
.A(n_1956),
.B(n_1694),
.Y(n_1963)
);

NOR2xp33_ASAP7_75t_L g1964 ( 
.A(n_1961),
.B(n_1701),
.Y(n_1964)
);

NOR3xp33_ASAP7_75t_L g1965 ( 
.A(n_1960),
.B(n_1959),
.C(n_1468),
.Y(n_1965)
);

NOR2x1_ASAP7_75t_L g1966 ( 
.A(n_1955),
.B(n_1359),
.Y(n_1966)
);

NOR2xp33_ASAP7_75t_L g1967 ( 
.A(n_1955),
.B(n_1701),
.Y(n_1967)
);

AOI22xp5_ASAP7_75t_SL g1968 ( 
.A1(n_1967),
.A2(n_1524),
.B1(n_1434),
.B2(n_1359),
.Y(n_1968)
);

XNOR2xp5_ASAP7_75t_L g1969 ( 
.A(n_1962),
.B(n_1373),
.Y(n_1969)
);

AND2x4_ASAP7_75t_L g1970 ( 
.A(n_1963),
.B(n_1694),
.Y(n_1970)
);

OAI22xp5_ASAP7_75t_SL g1971 ( 
.A1(n_1966),
.A2(n_1442),
.B1(n_1371),
.B2(n_1373),
.Y(n_1971)
);

INVx1_ASAP7_75t_L g1972 ( 
.A(n_1969),
.Y(n_1972)
);

INVx1_ASAP7_75t_L g1973 ( 
.A(n_1972),
.Y(n_1973)
);

NAND2xp5_ASAP7_75t_L g1974 ( 
.A(n_1973),
.B(n_1964),
.Y(n_1974)
);

INVx2_ASAP7_75t_L g1975 ( 
.A(n_1973),
.Y(n_1975)
);

NAND2xp5_ASAP7_75t_L g1976 ( 
.A(n_1975),
.B(n_1965),
.Y(n_1976)
);

OR2x6_ASAP7_75t_L g1977 ( 
.A(n_1974),
.B(n_1970),
.Y(n_1977)
);

INVxp33_ASAP7_75t_L g1978 ( 
.A(n_1976),
.Y(n_1978)
);

AND2x2_ASAP7_75t_L g1979 ( 
.A(n_1977),
.B(n_1968),
.Y(n_1979)
);

AO21x2_ASAP7_75t_L g1980 ( 
.A1(n_1979),
.A2(n_1971),
.B(n_1714),
.Y(n_1980)
);

AOI322xp5_ASAP7_75t_L g1981 ( 
.A1(n_1980),
.A2(n_1978),
.A3(n_1708),
.B1(n_1718),
.B2(n_1711),
.C1(n_1729),
.C2(n_1695),
.Y(n_1981)
);

OAI221xp5_ASAP7_75t_R g1982 ( 
.A1(n_1981),
.A2(n_1711),
.B1(n_1371),
.B2(n_1442),
.C(n_1721),
.Y(n_1982)
);

AOI211xp5_ASAP7_75t_L g1983 ( 
.A1(n_1982),
.A2(n_1359),
.B(n_1434),
.C(n_1378),
.Y(n_1983)
);


endmodule