module fake_netlist_6_548_n_2159 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_193, n_147, n_154, n_191, n_88, n_3, n_209, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_199, n_138, n_22, n_161, n_208, n_68, n_166, n_28, n_184, n_50, n_158, n_49, n_7, n_210, n_83, n_206, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_188, n_102, n_186, n_204, n_0, n_87, n_195, n_189, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_197, n_11, n_137, n_17, n_23, n_203, n_142, n_20, n_143, n_207, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_205, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_202, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_196, n_200, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_198, n_104, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_190, n_14, n_123, n_136, n_72, n_187, n_89, n_173, n_201, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_194, n_171, n_31, n_192, n_57, n_169, n_53, n_51, n_44, n_56, n_2159);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_193;
input n_147;
input n_154;
input n_191;
input n_88;
input n_3;
input n_209;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_199;
input n_138;
input n_22;
input n_161;
input n_208;
input n_68;
input n_166;
input n_28;
input n_184;
input n_50;
input n_158;
input n_49;
input n_7;
input n_210;
input n_83;
input n_206;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_188;
input n_102;
input n_186;
input n_204;
input n_0;
input n_87;
input n_195;
input n_189;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_197;
input n_11;
input n_137;
input n_17;
input n_23;
input n_203;
input n_142;
input n_20;
input n_143;
input n_207;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_205;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_202;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_196;
input n_200;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_190;
input n_14;
input n_123;
input n_136;
input n_72;
input n_187;
input n_89;
input n_173;
input n_201;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_194;
input n_171;
input n_31;
input n_192;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_2159;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_726;
wire n_2157;
wire n_212;
wire n_700;
wire n_1307;
wire n_2003;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_1853;
wire n_783;
wire n_1738;
wire n_798;
wire n_1575;
wire n_1854;
wire n_1923;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_2051;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1691;
wire n_1688;
wire n_1975;
wire n_1009;
wire n_1743;
wire n_1930;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1991;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_1844;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_1985;
wire n_447;
wire n_1803;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1867;
wire n_1704;
wire n_1078;
wire n_544;
wire n_250;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_2019;
wire n_836;
wire n_375;
wire n_2074;
wire n_522;
wire n_2129;
wire n_1261;
wire n_945;
wire n_1649;
wire n_2018;
wire n_2094;
wire n_1903;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_616;
wire n_658;
wire n_1874;
wire n_1119;
wire n_2013;
wire n_428;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_2044;
wire n_1954;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_1971;
wire n_2058;
wire n_2090;
wire n_405;
wire n_213;
wire n_538;
wire n_2004;
wire n_1106;
wire n_886;
wire n_1471;
wire n_953;
wire n_343;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_494;
wire n_539;
wire n_493;
wire n_2108;
wire n_454;
wire n_1421;
wire n_1936;
wire n_638;
wire n_1404;
wire n_1211;
wire n_2124;
wire n_381;
wire n_887;
wire n_1660;
wire n_1961;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_2155;
wire n_224;
wire n_1445;
wire n_1560;
wire n_1526;
wire n_734;
wire n_1088;
wire n_1894;
wire n_1231;
wire n_1978;
wire n_2085;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_1815;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1967;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1911;
wire n_1956;
wire n_1644;
wire n_2011;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_1986;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_2113;
wire n_1918;
wire n_577;
wire n_1843;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1909;
wire n_2080;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_2104;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_2093;
wire n_483;
wire n_1970;
wire n_608;
wire n_261;
wire n_2101;
wire n_630;
wire n_2059;
wire n_541;
wire n_512;
wire n_2073;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_1957;
wire n_219;
wire n_1907;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1876;
wire n_1895;
wire n_2123;
wire n_1697;
wire n_2143;
wire n_243;
wire n_979;
wire n_1873;
wire n_905;
wire n_1866;
wire n_1680;
wire n_322;
wire n_993;
wire n_689;
wire n_2031;
wire n_354;
wire n_2130;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1988;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_2009;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_2068;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_2072;
wire n_1354;
wire n_586;
wire n_423;
wire n_1875;
wire n_1865;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_1950;
wire n_530;
wire n_1563;
wire n_1912;
wire n_277;
wire n_1982;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_1927;
wire n_2028;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_2008;
wire n_1926;
wire n_1175;
wire n_328;
wire n_1386;
wire n_1896;
wire n_429;
wire n_1747;
wire n_1012;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1977;
wire n_1802;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_835;
wire n_242;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1801;
wire n_1886;
wire n_2092;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_2096;
wire n_1965;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_484;
wire n_2036;
wire n_2152;
wire n_1709;
wire n_1825;
wire n_1757;
wire n_1796;
wire n_1792;
wire n_891;
wire n_2067;
wire n_2136;
wire n_2082;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_2075;
wire n_1987;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_1052;
wire n_462;
wire n_1033;
wire n_1296;
wire n_1990;
wire n_304;
wire n_694;
wire n_2150;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_2078;
wire n_297;
wire n_595;
wire n_627;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1858;
wire n_1044;
wire n_2133;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_382;
wire n_673;
wire n_1969;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_2145;
wire n_1968;
wire n_898;
wire n_255;
wire n_284;
wire n_1952;
wire n_865;
wire n_925;
wire n_1932;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_2151;
wire n_1451;
wire n_963;
wire n_639;
wire n_320;
wire n_794;
wire n_727;
wire n_894;
wire n_1839;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_1863;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_1308;
wire n_2089;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_1913;
wire n_510;
wire n_837;
wire n_2097;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_2148;
wire n_977;
wire n_1005;
wire n_1947;
wire n_536;
wire n_1788;
wire n_1999;
wire n_622;
wire n_1469;
wire n_2060;
wire n_1838;
wire n_1835;
wire n_1776;
wire n_1766;
wire n_1959;
wire n_2002;
wire n_581;
wire n_2138;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_1878;
wire n_899;
wire n_738;
wire n_2012;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_2134;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_2069;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_1181;
wire n_2119;
wire n_1822;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_1992;
wire n_648;
wire n_657;
wire n_1049;
wire n_2057;
wire n_2103;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_1817;
wire n_927;
wire n_1849;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_2127;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_2137;
wire n_1626;
wire n_1507;
wire n_552;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_216;
wire n_912;
wire n_1857;
wire n_1519;
wire n_2144;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_2110;
wire n_731;
wire n_1502;
wire n_1659;
wire n_1955;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_683;
wire n_811;
wire n_1207;
wire n_527;
wire n_312;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_1897;
wire n_2064;
wire n_880;
wire n_2053;
wire n_2121;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_1966;
wire n_1942;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_1837;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_2132;
wire n_2063;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_211;
wire n_1483;
wire n_1834;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1993;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1919;
wire n_1080;
wire n_723;
wire n_1877;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1939;
wire n_2030;
wire n_1769;
wire n_1220;
wire n_1893;
wire n_556;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_2025;
wire n_1125;
wire n_970;
wire n_1980;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_1951;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_1286;
wire n_1773;
wire n_1775;
wire n_2115;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_1745;
wire n_914;
wire n_759;
wire n_1831;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_2146;
wire n_2131;
wire n_488;
wire n_497;
wire n_773;
wire n_1901;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1892;
wire n_1933;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_2000;
wire n_1917;
wire n_1580;
wire n_1425;
wire n_1881;
wire n_1267;
wire n_1281;
wire n_1806;
wire n_983;
wire n_2023;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_2158;
wire n_2087;
wire n_1855;
wire n_1636;
wire n_1437;
wire n_2135;
wire n_1645;
wire n_1832;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_2049;
wire n_1331;
wire n_736;
wire n_613;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_2100;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1995;
wire n_1594;
wire n_664;
wire n_1869;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_1889;
wire n_435;
wire n_1905;
wire n_2016;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_1937;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_2139;
wire n_2142;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1934;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_1871;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_1859;
wire n_2102;
wire n_238;
wire n_1095;
wire n_2024;
wire n_1595;
wire n_2156;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_1916;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_2153;
wire n_1847;
wire n_2052;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1841;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_1997;
wire n_340;
wire n_710;
wire n_1108;
wire n_1818;
wire n_1182;
wire n_1298;
wire n_2088;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1960;
wire n_2061;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1943;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1983;
wire n_1938;
wire n_1262;
wire n_218;
wire n_1891;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_239;
wire n_2037;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_2120;
wire n_1472;
wire n_2050;
wire n_1081;
wire n_402;
wire n_1870;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_2006;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_2017;
wire n_370;
wire n_1695;
wire n_1828;
wire n_2046;
wire n_650;
wire n_1046;
wire n_1940;
wire n_1979;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_1963;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1883;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_2084;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_1823;
wire n_227;
wire n_1974;
wire n_1720;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_1964;
wire n_1920;
wire n_2099;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_2007;
wire n_2039;
wire n_1946;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_1846;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_2141;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_1676;
wire n_833;
wire n_1830;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_1900;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_2021;
wire n_2114;
wire n_1086;
wire n_1066;
wire n_1948;
wire n_2125;
wire n_2026;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_2154;
wire n_560;
wire n_1906;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_1758;
wire n_1925;
wire n_737;
wire n_1318;
wire n_1914;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_2056;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1984;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_1931;
wire n_2083;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_1941;
wire n_2128;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1962;
wire n_1559;
wire n_1725;
wire n_1928;
wire n_1872;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1741;
wire n_1325;
wire n_1002;
wire n_1746;
wire n_1949;
wire n_545;
wire n_489;
wire n_1804;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_2054;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_2062;
wire n_2041;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1860;
wire n_1904;
wire n_1200;
wire n_2070;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1908;
wire n_1454;
wire n_2126;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_2045;
wire n_817;
wire n_262;
wire n_897;
wire n_846;
wire n_2066;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1800;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1882;
wire n_1076;
wire n_1118;
wire n_1007;
wire n_1807;
wire n_1929;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_1879;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_680;
wire n_367;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_1953;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1976;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_2122;
wire n_2109;
wire n_1435;
wire n_969;
wire n_988;
wire n_2140;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_2029;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_1810;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_2020;
wire n_1729;
wire n_669;
wire n_2048;
wire n_300;
wire n_222;
wire n_2005;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_2076;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1785;
wire n_763;
wire n_1147;
wire n_1848;
wire n_360;
wire n_1754;
wire n_2149;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_1994;
wire n_895;
wire n_866;
wire n_1227;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_1924;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_1174;
wire n_1944;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_844;
wire n_448;
wire n_1017;
wire n_2117;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_2081;
wire n_234;
wire n_2022;
wire n_1945;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_2112;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_2034;
wire n_576;
wire n_1028;
wire n_2106;
wire n_472;
wire n_270;
wire n_414;
wire n_1922;
wire n_563;
wire n_2032;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_1973;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_2015;
wire n_2118;
wire n_2111;
wire n_390;
wire n_1148;
wire n_334;
wire n_1989;
wire n_1161;
wire n_1085;
wire n_232;
wire n_2014;
wire n_2042;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1972;
wire n_1525;
wire n_455;
wire n_1585;
wire n_1851;
wire n_363;
wire n_1799;
wire n_1090;
wire n_2147;
wire n_592;
wire n_1816;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_1829;
wire n_503;
wire n_2035;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_2033;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_2071;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_2010;
wire n_1651;
wire n_1198;
wire n_2047;
wire n_2095;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1998;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1981;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_1996;
wire n_249;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_2043;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1921;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_2065;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_271;
wire n_404;
wire n_2001;
wire n_2107;
wire n_1884;
wire n_2040;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1819;
wire n_2055;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_2038;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_373;
wire n_1632;
wire n_1890;
wire n_1805;
wire n_257;
wire n_1557;
wire n_1888;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_1850;
wire n_1898;
wire n_1868;
wire n_2079;
wire n_1089;
wire n_1887;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_1242;
wire n_2086;
wire n_1836;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1899;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1856;
wire n_1862;
wire n_1958;
wire n_2077;
wire n_339;
wire n_784;
wire n_434;
wire n_315;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_2105;
wire n_2098;
wire n_540;
wire n_1423;
wire n_1935;
wire n_2027;
wire n_457;
wire n_2091;
wire n_364;
wire n_1915;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_2116;
wire n_336;
wire n_1885;
wire n_1013;
wire n_1259;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_157),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_145),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_62),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_147),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_16),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_79),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_206),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_156),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_59),
.Y(n_219)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_111),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_53),
.Y(n_221)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_59),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_170),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_96),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_152),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_140),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_207),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_204),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_198),
.Y(n_229)
);

CKINVDCx16_ASAP7_75t_R g230 ( 
.A(n_27),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_33),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_117),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_42),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_62),
.Y(n_234)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_188),
.Y(n_235)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_112),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_75),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_44),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_104),
.Y(n_239)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_82),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_86),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_15),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_14),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_179),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_175),
.Y(n_245)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_84),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_16),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_201),
.Y(n_248)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_186),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_139),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_133),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_172),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_122),
.Y(n_253)
);

BUFx3_ASAP7_75t_L g254 ( 
.A(n_108),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_9),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_116),
.Y(n_256)
);

INVx2_ASAP7_75t_SL g257 ( 
.A(n_200),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_56),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_103),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_25),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_185),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_88),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_202),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_126),
.Y(n_264)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_183),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_89),
.Y(n_266)
);

INVx1_ASAP7_75t_SL g267 ( 
.A(n_0),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_44),
.Y(n_268)
);

INVx1_ASAP7_75t_SL g269 ( 
.A(n_49),
.Y(n_269)
);

CKINVDCx16_ASAP7_75t_R g270 ( 
.A(n_38),
.Y(n_270)
);

BUFx2_ASAP7_75t_SL g271 ( 
.A(n_13),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_41),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_171),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_73),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_43),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_191),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_36),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_168),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_107),
.Y(n_279)
);

INVx1_ASAP7_75t_SL g280 ( 
.A(n_41),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_197),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_77),
.Y(n_282)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_165),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_160),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_78),
.Y(n_285)
);

INVx2_ASAP7_75t_SL g286 ( 
.A(n_72),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_124),
.Y(n_287)
);

BUFx3_ASAP7_75t_L g288 ( 
.A(n_80),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_159),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_129),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_73),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_28),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_187),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_6),
.Y(n_294)
);

CKINVDCx16_ASAP7_75t_R g295 ( 
.A(n_24),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_74),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_97),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_82),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_98),
.Y(n_299)
);

BUFx8_ASAP7_75t_SL g300 ( 
.A(n_65),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_130),
.Y(n_301)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_192),
.Y(n_302)
);

BUFx10_ASAP7_75t_L g303 ( 
.A(n_195),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_46),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_177),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_203),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_56),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_146),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_127),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_35),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_138),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_79),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_189),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_99),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_13),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_27),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_0),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_55),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_45),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_46),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_178),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_23),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_109),
.Y(n_323)
);

HB1xp67_ASAP7_75t_L g324 ( 
.A(n_182),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_135),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_7),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_153),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_33),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_12),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_15),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_72),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_29),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_21),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_53),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_83),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_184),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_2),
.Y(n_337)
);

BUFx10_ASAP7_75t_L g338 ( 
.A(n_106),
.Y(n_338)
);

INVx2_ASAP7_75t_L g339 ( 
.A(n_50),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_81),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_199),
.Y(n_341)
);

INVx2_ASAP7_75t_L g342 ( 
.A(n_162),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_36),
.Y(n_343)
);

BUFx8_ASAP7_75t_SL g344 ( 
.A(n_173),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_113),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_205),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_74),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_196),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_180),
.Y(n_349)
);

BUFx10_ASAP7_75t_L g350 ( 
.A(n_174),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_52),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_71),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_63),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_93),
.Y(n_354)
);

BUFx10_ASAP7_75t_L g355 ( 
.A(n_83),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_120),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_141),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_17),
.Y(n_358)
);

INVx2_ASAP7_75t_L g359 ( 
.A(n_125),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_63),
.Y(n_360)
);

BUFx10_ASAP7_75t_L g361 ( 
.A(n_22),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_194),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_176),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_17),
.Y(n_364)
);

BUFx6f_ASAP7_75t_L g365 ( 
.A(n_5),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_136),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_64),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_69),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_22),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_210),
.Y(n_370)
);

INVx1_ASAP7_75t_SL g371 ( 
.A(n_11),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_6),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_48),
.Y(n_373)
);

BUFx3_ASAP7_75t_L g374 ( 
.A(n_60),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_31),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_69),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_5),
.Y(n_377)
);

CKINVDCx20_ASAP7_75t_R g378 ( 
.A(n_42),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_87),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_57),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_149),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_102),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_26),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_32),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_84),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_3),
.Y(n_386)
);

INVx2_ASAP7_75t_SL g387 ( 
.A(n_86),
.Y(n_387)
);

BUFx10_ASAP7_75t_L g388 ( 
.A(n_14),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_94),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_123),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_91),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_181),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_54),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_155),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_3),
.Y(n_395)
);

BUFx3_ASAP7_75t_L g396 ( 
.A(n_164),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_34),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_11),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_134),
.Y(n_399)
);

CKINVDCx16_ASAP7_75t_R g400 ( 
.A(n_40),
.Y(n_400)
);

BUFx6f_ASAP7_75t_L g401 ( 
.A(n_101),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_45),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_7),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_54),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_208),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_25),
.Y(n_406)
);

CKINVDCx20_ASAP7_75t_R g407 ( 
.A(n_190),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_52),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_8),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_92),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_67),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_71),
.Y(n_412)
);

BUFx10_ASAP7_75t_L g413 ( 
.A(n_2),
.Y(n_413)
);

CKINVDCx20_ASAP7_75t_R g414 ( 
.A(n_218),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_344),
.Y(n_415)
);

NOR2xp67_ASAP7_75t_L g416 ( 
.A(n_286),
.B(n_1),
.Y(n_416)
);

HB1xp67_ASAP7_75t_L g417 ( 
.A(n_230),
.Y(n_417)
);

HB1xp67_ASAP7_75t_L g418 ( 
.A(n_230),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_365),
.Y(n_419)
);

INVxp67_ASAP7_75t_SL g420 ( 
.A(n_324),
.Y(n_420)
);

BUFx6f_ASAP7_75t_L g421 ( 
.A(n_401),
.Y(n_421)
);

CKINVDCx20_ASAP7_75t_R g422 ( 
.A(n_226),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_365),
.Y(n_423)
);

INVxp67_ASAP7_75t_SL g424 ( 
.A(n_254),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_365),
.Y(n_425)
);

INVx2_ASAP7_75t_L g426 ( 
.A(n_249),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_365),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_365),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_300),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_211),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_365),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_222),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_222),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_212),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_240),
.Y(n_435)
);

CKINVDCx16_ASAP7_75t_R g436 ( 
.A(n_270),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_214),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_217),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_228),
.Y(n_439)
);

CKINVDCx20_ASAP7_75t_R g440 ( 
.A(n_297),
.Y(n_440)
);

BUFx2_ASAP7_75t_SL g441 ( 
.A(n_257),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_232),
.Y(n_442)
);

HB1xp67_ASAP7_75t_L g443 ( 
.A(n_270),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_244),
.Y(n_444)
);

CKINVDCx20_ASAP7_75t_R g445 ( 
.A(n_407),
.Y(n_445)
);

NOR2xp33_ASAP7_75t_L g446 ( 
.A(n_257),
.B(n_1),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_240),
.Y(n_447)
);

INVxp67_ASAP7_75t_SL g448 ( 
.A(n_237),
.Y(n_448)
);

NOR2xp33_ASAP7_75t_L g449 ( 
.A(n_223),
.B(n_4),
.Y(n_449)
);

HB1xp67_ASAP7_75t_L g450 ( 
.A(n_295),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_245),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_246),
.Y(n_452)
);

AND2x2_ASAP7_75t_L g453 ( 
.A(n_288),
.B(n_4),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_248),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_246),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_339),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_251),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_339),
.Y(n_458)
);

HB1xp67_ASAP7_75t_L g459 ( 
.A(n_295),
.Y(n_459)
);

INVxp67_ASAP7_75t_L g460 ( 
.A(n_286),
.Y(n_460)
);

CKINVDCx20_ASAP7_75t_R g461 ( 
.A(n_259),
.Y(n_461)
);

CKINVDCx5p33_ASAP7_75t_R g462 ( 
.A(n_263),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_266),
.Y(n_463)
);

CKINVDCx20_ASAP7_75t_R g464 ( 
.A(n_276),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_288),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_288),
.Y(n_466)
);

NAND2xp33_ASAP7_75t_R g467 ( 
.A(n_279),
.B(n_8),
.Y(n_467)
);

CKINVDCx20_ASAP7_75t_R g468 ( 
.A(n_284),
.Y(n_468)
);

CKINVDCx20_ASAP7_75t_R g469 ( 
.A(n_287),
.Y(n_469)
);

INVxp67_ASAP7_75t_L g470 ( 
.A(n_387),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_374),
.Y(n_471)
);

CKINVDCx5p33_ASAP7_75t_R g472 ( 
.A(n_290),
.Y(n_472)
);

CKINVDCx5p33_ASAP7_75t_R g473 ( 
.A(n_293),
.Y(n_473)
);

INVx2_ASAP7_75t_L g474 ( 
.A(n_249),
.Y(n_474)
);

INVxp67_ASAP7_75t_SL g475 ( 
.A(n_237),
.Y(n_475)
);

CKINVDCx20_ASAP7_75t_R g476 ( 
.A(n_301),
.Y(n_476)
);

NOR2xp67_ASAP7_75t_L g477 ( 
.A(n_387),
.B(n_9),
.Y(n_477)
);

INVxp67_ASAP7_75t_L g478 ( 
.A(n_255),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_374),
.Y(n_479)
);

HB1xp67_ASAP7_75t_L g480 ( 
.A(n_400),
.Y(n_480)
);

INVxp67_ASAP7_75t_L g481 ( 
.A(n_255),
.Y(n_481)
);

INVxp67_ASAP7_75t_SL g482 ( 
.A(n_254),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_374),
.Y(n_483)
);

CKINVDCx20_ASAP7_75t_R g484 ( 
.A(n_305),
.Y(n_484)
);

HB1xp67_ASAP7_75t_L g485 ( 
.A(n_400),
.Y(n_485)
);

NOR2xp33_ASAP7_75t_L g486 ( 
.A(n_223),
.B(n_10),
.Y(n_486)
);

CKINVDCx5p33_ASAP7_75t_R g487 ( 
.A(n_306),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_272),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_272),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_277),
.Y(n_490)
);

INVx2_ASAP7_75t_L g491 ( 
.A(n_249),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_277),
.Y(n_492)
);

CKINVDCx5p33_ASAP7_75t_R g493 ( 
.A(n_308),
.Y(n_493)
);

AND2x2_ASAP7_75t_L g494 ( 
.A(n_254),
.B(n_12),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_285),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_285),
.Y(n_496)
);

CKINVDCx5p33_ASAP7_75t_R g497 ( 
.A(n_311),
.Y(n_497)
);

CKINVDCx20_ASAP7_75t_R g498 ( 
.A(n_314),
.Y(n_498)
);

AND2x2_ASAP7_75t_L g499 ( 
.A(n_396),
.B(n_294),
.Y(n_499)
);

NOR2xp33_ASAP7_75t_L g500 ( 
.A(n_224),
.B(n_18),
.Y(n_500)
);

CKINVDCx5p33_ASAP7_75t_R g501 ( 
.A(n_321),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_294),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_298),
.Y(n_503)
);

CKINVDCx5p33_ASAP7_75t_R g504 ( 
.A(n_323),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_298),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_329),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_329),
.Y(n_507)
);

CKINVDCx5p33_ASAP7_75t_R g508 ( 
.A(n_325),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_334),
.Y(n_509)
);

INVxp67_ASAP7_75t_L g510 ( 
.A(n_334),
.Y(n_510)
);

CKINVDCx20_ASAP7_75t_R g511 ( 
.A(n_327),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_347),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_347),
.Y(n_513)
);

CKINVDCx5p33_ASAP7_75t_R g514 ( 
.A(n_336),
.Y(n_514)
);

CKINVDCx5p33_ASAP7_75t_R g515 ( 
.A(n_362),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_351),
.Y(n_516)
);

NOR2xp33_ASAP7_75t_R g517 ( 
.A(n_370),
.B(n_90),
.Y(n_517)
);

CKINVDCx5p33_ASAP7_75t_R g518 ( 
.A(n_379),
.Y(n_518)
);

CKINVDCx5p33_ASAP7_75t_R g519 ( 
.A(n_381),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_351),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_360),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_360),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_419),
.Y(n_523)
);

INVx2_ASAP7_75t_L g524 ( 
.A(n_421),
.Y(n_524)
);

OAI21x1_ASAP7_75t_L g525 ( 
.A1(n_426),
.A2(n_235),
.B(n_220),
.Y(n_525)
);

INVx2_ASAP7_75t_L g526 ( 
.A(n_421),
.Y(n_526)
);

INVx2_ASAP7_75t_L g527 ( 
.A(n_421),
.Y(n_527)
);

INVx2_ASAP7_75t_L g528 ( 
.A(n_421),
.Y(n_528)
);

AND2x4_ASAP7_75t_L g529 ( 
.A(n_494),
.B(n_396),
.Y(n_529)
);

BUFx6f_ASAP7_75t_L g530 ( 
.A(n_421),
.Y(n_530)
);

AND2x2_ASAP7_75t_L g531 ( 
.A(n_499),
.B(n_396),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_419),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_423),
.Y(n_533)
);

OAI21x1_ASAP7_75t_L g534 ( 
.A1(n_426),
.A2(n_235),
.B(n_220),
.Y(n_534)
);

INVx3_ASAP7_75t_L g535 ( 
.A(n_421),
.Y(n_535)
);

NOR2xp33_ASAP7_75t_SL g536 ( 
.A(n_436),
.B(n_355),
.Y(n_536)
);

AND2x4_ASAP7_75t_L g537 ( 
.A(n_494),
.B(n_236),
.Y(n_537)
);

INVx2_ASAP7_75t_L g538 ( 
.A(n_426),
.Y(n_538)
);

BUFx6f_ASAP7_75t_L g539 ( 
.A(n_474),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_423),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_L g541 ( 
.A(n_424),
.B(n_382),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_SL g542 ( 
.A(n_416),
.B(n_303),
.Y(n_542)
);

CKINVDCx5p33_ASAP7_75t_R g543 ( 
.A(n_461),
.Y(n_543)
);

BUFx6f_ASAP7_75t_L g544 ( 
.A(n_474),
.Y(n_544)
);

BUFx6f_ASAP7_75t_L g545 ( 
.A(n_474),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_425),
.Y(n_546)
);

BUFx6f_ASAP7_75t_L g547 ( 
.A(n_491),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_L g548 ( 
.A(n_482),
.B(n_389),
.Y(n_548)
);

BUFx6f_ASAP7_75t_L g549 ( 
.A(n_491),
.Y(n_549)
);

NAND2xp33_ASAP7_75t_SL g550 ( 
.A(n_453),
.B(n_238),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_425),
.Y(n_551)
);

OA21x2_ASAP7_75t_L g552 ( 
.A1(n_491),
.A2(n_368),
.B(n_364),
.Y(n_552)
);

BUFx2_ASAP7_75t_L g553 ( 
.A(n_417),
.Y(n_553)
);

INVx3_ASAP7_75t_L g554 ( 
.A(n_427),
.Y(n_554)
);

BUFx2_ASAP7_75t_L g555 ( 
.A(n_418),
.Y(n_555)
);

OA21x2_ASAP7_75t_L g556 ( 
.A1(n_427),
.A2(n_368),
.B(n_364),
.Y(n_556)
);

BUFx6f_ASAP7_75t_L g557 ( 
.A(n_428),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_428),
.Y(n_558)
);

INVx4_ASAP7_75t_L g559 ( 
.A(n_499),
.Y(n_559)
);

INVx3_ASAP7_75t_L g560 ( 
.A(n_431),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_431),
.Y(n_561)
);

BUFx2_ASAP7_75t_L g562 ( 
.A(n_443),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_L g563 ( 
.A(n_446),
.B(n_392),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_488),
.Y(n_564)
);

BUFx6f_ASAP7_75t_L g565 ( 
.A(n_432),
.Y(n_565)
);

CKINVDCx14_ASAP7_75t_R g566 ( 
.A(n_415),
.Y(n_566)
);

AND2x2_ASAP7_75t_L g567 ( 
.A(n_453),
.B(n_342),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_L g568 ( 
.A(n_441),
.B(n_465),
.Y(n_568)
);

AND2x2_ASAP7_75t_L g569 ( 
.A(n_465),
.B(n_342),
.Y(n_569)
);

CKINVDCx5p33_ASAP7_75t_R g570 ( 
.A(n_464),
.Y(n_570)
);

INVx2_ASAP7_75t_L g571 ( 
.A(n_432),
.Y(n_571)
);

INVx2_ASAP7_75t_L g572 ( 
.A(n_433),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_488),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_433),
.Y(n_574)
);

INVx2_ASAP7_75t_L g575 ( 
.A(n_435),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_489),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_489),
.Y(n_577)
);

INVx3_ASAP7_75t_L g578 ( 
.A(n_435),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_490),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_490),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_492),
.Y(n_581)
);

BUFx6f_ASAP7_75t_L g582 ( 
.A(n_447),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_492),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_L g584 ( 
.A(n_441),
.B(n_466),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_L g585 ( 
.A(n_466),
.B(n_399),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_L g586 ( 
.A(n_471),
.B(n_405),
.Y(n_586)
);

BUFx6f_ASAP7_75t_L g587 ( 
.A(n_447),
.Y(n_587)
);

INVx2_ASAP7_75t_L g588 ( 
.A(n_452),
.Y(n_588)
);

BUFx2_ASAP7_75t_L g589 ( 
.A(n_450),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_495),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_495),
.Y(n_591)
);

AND2x2_ASAP7_75t_L g592 ( 
.A(n_471),
.B(n_342),
.Y(n_592)
);

AND2x4_ASAP7_75t_L g593 ( 
.A(n_479),
.B(n_236),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_496),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_L g595 ( 
.A(n_479),
.B(n_265),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_L g596 ( 
.A(n_483),
.B(n_265),
.Y(n_596)
);

OAI22xp5_ASAP7_75t_L g597 ( 
.A1(n_436),
.A2(n_268),
.B1(n_307),
.B2(n_241),
.Y(n_597)
);

INVx3_ASAP7_75t_L g598 ( 
.A(n_452),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_496),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_502),
.Y(n_600)
);

INVx2_ASAP7_75t_L g601 ( 
.A(n_455),
.Y(n_601)
);

OAI22xp5_ASAP7_75t_SL g602 ( 
.A1(n_414),
.A2(n_378),
.B1(n_326),
.B2(n_333),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_502),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_503),
.Y(n_604)
);

HB1xp67_ASAP7_75t_L g605 ( 
.A(n_459),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_503),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_505),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_505),
.Y(n_608)
);

BUFx6f_ASAP7_75t_L g609 ( 
.A(n_455),
.Y(n_609)
);

INVxp67_ASAP7_75t_SL g610 ( 
.A(n_568),
.Y(n_610)
);

INVx2_ASAP7_75t_L g611 ( 
.A(n_538),
.Y(n_611)
);

NAND3xp33_ASAP7_75t_L g612 ( 
.A(n_550),
.B(n_420),
.C(n_430),
.Y(n_612)
);

INVx2_ASAP7_75t_L g613 ( 
.A(n_538),
.Y(n_613)
);

AND2x2_ASAP7_75t_L g614 ( 
.A(n_559),
.B(n_483),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_552),
.Y(n_615)
);

INVx4_ASAP7_75t_L g616 ( 
.A(n_559),
.Y(n_616)
);

BUFx10_ASAP7_75t_L g617 ( 
.A(n_529),
.Y(n_617)
);

INVx2_ASAP7_75t_L g618 ( 
.A(n_538),
.Y(n_618)
);

AND2x6_ASAP7_75t_L g619 ( 
.A(n_567),
.B(n_359),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_L g620 ( 
.A(n_559),
.B(n_434),
.Y(n_620)
);

OR2x6_ASAP7_75t_L g621 ( 
.A(n_542),
.B(n_271),
.Y(n_621)
);

AND2x2_ASAP7_75t_SL g622 ( 
.A(n_567),
.B(n_359),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_552),
.Y(n_623)
);

CKINVDCx5p33_ASAP7_75t_R g624 ( 
.A(n_543),
.Y(n_624)
);

INVx2_ASAP7_75t_L g625 ( 
.A(n_538),
.Y(n_625)
);

BUFx6f_ASAP7_75t_L g626 ( 
.A(n_530),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_552),
.Y(n_627)
);

INVx2_ASAP7_75t_SL g628 ( 
.A(n_531),
.Y(n_628)
);

INVx2_ASAP7_75t_L g629 ( 
.A(n_532),
.Y(n_629)
);

BUFx4f_ASAP7_75t_L g630 ( 
.A(n_556),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_552),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_552),
.Y(n_632)
);

NOR2xp33_ASAP7_75t_L g633 ( 
.A(n_541),
.B(n_437),
.Y(n_633)
);

INVx2_ASAP7_75t_L g634 ( 
.A(n_532),
.Y(n_634)
);

BUFx6f_ASAP7_75t_L g635 ( 
.A(n_530),
.Y(n_635)
);

OR2x2_ASAP7_75t_L g636 ( 
.A(n_605),
.B(n_553),
.Y(n_636)
);

NOR2x1p5_ASAP7_75t_L g637 ( 
.A(n_568),
.B(n_429),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_552),
.Y(n_638)
);

INVx2_ASAP7_75t_L g639 ( 
.A(n_533),
.Y(n_639)
);

INVx2_ASAP7_75t_L g640 ( 
.A(n_533),
.Y(n_640)
);

INVx2_ASAP7_75t_L g641 ( 
.A(n_540),
.Y(n_641)
);

AND2x4_ASAP7_75t_L g642 ( 
.A(n_559),
.B(n_224),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_556),
.Y(n_643)
);

BUFx6f_ASAP7_75t_L g644 ( 
.A(n_530),
.Y(n_644)
);

NAND2xp33_ASAP7_75t_L g645 ( 
.A(n_563),
.B(n_438),
.Y(n_645)
);

OAI22xp5_ASAP7_75t_L g646 ( 
.A1(n_563),
.A2(n_469),
.B1(n_476),
.B2(n_468),
.Y(n_646)
);

INVx3_ASAP7_75t_L g647 ( 
.A(n_530),
.Y(n_647)
);

INVx2_ASAP7_75t_L g648 ( 
.A(n_540),
.Y(n_648)
);

OR2x2_ASAP7_75t_L g649 ( 
.A(n_605),
.B(n_480),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_556),
.Y(n_650)
);

OR2x6_ASAP7_75t_L g651 ( 
.A(n_542),
.B(n_271),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_SL g652 ( 
.A(n_559),
.B(n_439),
.Y(n_652)
);

CKINVDCx20_ASAP7_75t_R g653 ( 
.A(n_543),
.Y(n_653)
);

INVx2_ASAP7_75t_L g654 ( 
.A(n_546),
.Y(n_654)
);

INVx3_ASAP7_75t_L g655 ( 
.A(n_530),
.Y(n_655)
);

INVx2_ASAP7_75t_L g656 ( 
.A(n_546),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_L g657 ( 
.A(n_541),
.B(n_442),
.Y(n_657)
);

BUFx10_ASAP7_75t_L g658 ( 
.A(n_529),
.Y(n_658)
);

INVxp67_ASAP7_75t_L g659 ( 
.A(n_553),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_556),
.Y(n_660)
);

OAI22xp5_ASAP7_75t_L g661 ( 
.A1(n_548),
.A2(n_498),
.B1(n_511),
.B2(n_484),
.Y(n_661)
);

INVxp67_ASAP7_75t_L g662 ( 
.A(n_553),
.Y(n_662)
);

NOR2xp33_ASAP7_75t_L g663 ( 
.A(n_548),
.B(n_444),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_529),
.B(n_567),
.Y(n_664)
);

INVx2_ASAP7_75t_L g665 ( 
.A(n_551),
.Y(n_665)
);

BUFx2_ASAP7_75t_L g666 ( 
.A(n_550),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_556),
.Y(n_667)
);

INVx2_ASAP7_75t_L g668 ( 
.A(n_551),
.Y(n_668)
);

INVx2_ASAP7_75t_L g669 ( 
.A(n_561),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_SL g670 ( 
.A(n_536),
.B(n_451),
.Y(n_670)
);

NOR2xp33_ASAP7_75t_L g671 ( 
.A(n_585),
.B(n_454),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_529),
.B(n_457),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_556),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_561),
.Y(n_674)
);

INVx2_ASAP7_75t_L g675 ( 
.A(n_523),
.Y(n_675)
);

OAI22xp5_ASAP7_75t_L g676 ( 
.A1(n_529),
.A2(n_463),
.B1(n_472),
.B2(n_462),
.Y(n_676)
);

AND2x6_ASAP7_75t_L g677 ( 
.A(n_537),
.B(n_359),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_SL g678 ( 
.A(n_536),
.B(n_473),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_523),
.Y(n_679)
);

AOI21x1_ASAP7_75t_L g680 ( 
.A1(n_523),
.A2(n_227),
.B(n_225),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_558),
.Y(n_681)
);

INVx2_ASAP7_75t_L g682 ( 
.A(n_558),
.Y(n_682)
);

CKINVDCx5p33_ASAP7_75t_R g683 ( 
.A(n_570),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_558),
.Y(n_684)
);

NAND2xp33_ASAP7_75t_L g685 ( 
.A(n_585),
.B(n_487),
.Y(n_685)
);

OR2x6_ASAP7_75t_L g686 ( 
.A(n_584),
.B(n_225),
.Y(n_686)
);

NOR2xp33_ASAP7_75t_L g687 ( 
.A(n_586),
.B(n_493),
.Y(n_687)
);

INVx2_ASAP7_75t_SL g688 ( 
.A(n_531),
.Y(n_688)
);

BUFx3_ASAP7_75t_L g689 ( 
.A(n_531),
.Y(n_689)
);

INVx2_ASAP7_75t_L g690 ( 
.A(n_539),
.Y(n_690)
);

AOI22xp5_ASAP7_75t_L g691 ( 
.A1(n_555),
.A2(n_322),
.B1(n_486),
.B2(n_449),
.Y(n_691)
);

HB1xp67_ASAP7_75t_L g692 ( 
.A(n_555),
.Y(n_692)
);

AND2x2_ASAP7_75t_L g693 ( 
.A(n_569),
.B(n_448),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_564),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_564),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_573),
.Y(n_696)
);

INVx1_ASAP7_75t_SL g697 ( 
.A(n_570),
.Y(n_697)
);

INVx2_ASAP7_75t_SL g698 ( 
.A(n_537),
.Y(n_698)
);

NAND3xp33_ASAP7_75t_L g699 ( 
.A(n_586),
.B(n_501),
.C(n_497),
.Y(n_699)
);

INVx2_ASAP7_75t_SL g700 ( 
.A(n_537),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_573),
.Y(n_701)
);

INVx2_ASAP7_75t_L g702 ( 
.A(n_539),
.Y(n_702)
);

INVx2_ASAP7_75t_L g703 ( 
.A(n_539),
.Y(n_703)
);

INVx2_ASAP7_75t_L g704 ( 
.A(n_539),
.Y(n_704)
);

INVx2_ASAP7_75t_L g705 ( 
.A(n_539),
.Y(n_705)
);

NOR2xp33_ASAP7_75t_L g706 ( 
.A(n_584),
.B(n_504),
.Y(n_706)
);

AND2x2_ASAP7_75t_L g707 ( 
.A(n_569),
.B(n_448),
.Y(n_707)
);

INVx2_ASAP7_75t_L g708 ( 
.A(n_539),
.Y(n_708)
);

INVx3_ASAP7_75t_L g709 ( 
.A(n_530),
.Y(n_709)
);

AND2x2_ASAP7_75t_L g710 ( 
.A(n_569),
.B(n_475),
.Y(n_710)
);

INVx4_ASAP7_75t_L g711 ( 
.A(n_530),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_576),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_L g713 ( 
.A(n_537),
.B(n_508),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_L g714 ( 
.A(n_537),
.B(n_514),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_576),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_577),
.Y(n_716)
);

OR2x2_ASAP7_75t_L g717 ( 
.A(n_555),
.B(n_485),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_577),
.Y(n_718)
);

NOR2xp33_ASAP7_75t_L g719 ( 
.A(n_562),
.B(n_515),
.Y(n_719)
);

AND2x2_ASAP7_75t_L g720 ( 
.A(n_592),
.B(n_475),
.Y(n_720)
);

INVx2_ASAP7_75t_L g721 ( 
.A(n_539),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_579),
.Y(n_722)
);

INVx2_ASAP7_75t_L g723 ( 
.A(n_539),
.Y(n_723)
);

AND2x2_ASAP7_75t_L g724 ( 
.A(n_592),
.B(n_456),
.Y(n_724)
);

NOR2xp33_ASAP7_75t_L g725 ( 
.A(n_562),
.B(n_518),
.Y(n_725)
);

BUFx3_ASAP7_75t_L g726 ( 
.A(n_593),
.Y(n_726)
);

BUFx6f_ASAP7_75t_L g727 ( 
.A(n_530),
.Y(n_727)
);

XOR2xp5_ASAP7_75t_L g728 ( 
.A(n_602),
.B(n_422),
.Y(n_728)
);

AND2x2_ASAP7_75t_L g729 ( 
.A(n_592),
.B(n_456),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_579),
.Y(n_730)
);

AND2x4_ASAP7_75t_L g731 ( 
.A(n_593),
.B(n_227),
.Y(n_731)
);

AND2x6_ASAP7_75t_L g732 ( 
.A(n_593),
.B(n_401),
.Y(n_732)
);

AND2x6_ASAP7_75t_L g733 ( 
.A(n_593),
.B(n_401),
.Y(n_733)
);

INVx5_ASAP7_75t_L g734 ( 
.A(n_544),
.Y(n_734)
);

INVx2_ASAP7_75t_L g735 ( 
.A(n_544),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_SL g736 ( 
.A(n_562),
.B(n_519),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_L g737 ( 
.A(n_535),
.B(n_554),
.Y(n_737)
);

OR2x6_ASAP7_75t_L g738 ( 
.A(n_589),
.B(n_416),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_580),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_580),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_SL g741 ( 
.A(n_589),
.B(n_517),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_L g742 ( 
.A(n_535),
.B(n_229),
.Y(n_742)
);

BUFx3_ASAP7_75t_L g743 ( 
.A(n_593),
.Y(n_743)
);

INVx1_ASAP7_75t_SL g744 ( 
.A(n_589),
.Y(n_744)
);

INVx2_ASAP7_75t_SL g745 ( 
.A(n_581),
.Y(n_745)
);

OR2x6_ASAP7_75t_L g746 ( 
.A(n_595),
.B(n_477),
.Y(n_746)
);

AOI22xp33_ASAP7_75t_L g747 ( 
.A1(n_595),
.A2(n_500),
.B1(n_477),
.B2(n_380),
.Y(n_747)
);

CKINVDCx16_ASAP7_75t_R g748 ( 
.A(n_597),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_SL g749 ( 
.A(n_597),
.B(n_303),
.Y(n_749)
);

INVx2_ASAP7_75t_L g750 ( 
.A(n_544),
.Y(n_750)
);

INVx6_ASAP7_75t_L g751 ( 
.A(n_557),
.Y(n_751)
);

AOI22xp33_ASAP7_75t_L g752 ( 
.A1(n_596),
.A2(n_380),
.B1(n_386),
.B2(n_372),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_581),
.Y(n_753)
);

INVx2_ASAP7_75t_L g754 ( 
.A(n_544),
.Y(n_754)
);

INVx2_ASAP7_75t_L g755 ( 
.A(n_544),
.Y(n_755)
);

INVx4_ASAP7_75t_L g756 ( 
.A(n_557),
.Y(n_756)
);

BUFx3_ASAP7_75t_L g757 ( 
.A(n_583),
.Y(n_757)
);

INVx2_ASAP7_75t_SL g758 ( 
.A(n_583),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_535),
.B(n_229),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_590),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_535),
.B(n_239),
.Y(n_761)
);

INVx2_ASAP7_75t_L g762 ( 
.A(n_544),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_SL g763 ( 
.A(n_706),
.B(n_440),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_L g764 ( 
.A(n_610),
.B(n_622),
.Y(n_764)
);

INVx4_ASAP7_75t_L g765 ( 
.A(n_616),
.Y(n_765)
);

INVx2_ASAP7_75t_L g766 ( 
.A(n_629),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_L g767 ( 
.A(n_622),
.B(n_578),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_698),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_698),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_L g770 ( 
.A(n_622),
.B(n_578),
.Y(n_770)
);

INVx2_ASAP7_75t_SL g771 ( 
.A(n_636),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_SL g772 ( 
.A(n_700),
.B(n_401),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_633),
.B(n_578),
.Y(n_773)
);

INVx2_ASAP7_75t_L g774 ( 
.A(n_629),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_663),
.B(n_578),
.Y(n_775)
);

BUFx6f_ASAP7_75t_L g776 ( 
.A(n_617),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_L g777 ( 
.A(n_671),
.B(n_578),
.Y(n_777)
);

AOI22xp5_ASAP7_75t_L g778 ( 
.A1(n_687),
.A2(n_445),
.B1(n_467),
.B2(n_566),
.Y(n_778)
);

NOR2xp33_ASAP7_75t_L g779 ( 
.A(n_657),
.B(n_566),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_700),
.B(n_598),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_628),
.B(n_598),
.Y(n_781)
);

NOR2xp33_ASAP7_75t_L g782 ( 
.A(n_719),
.B(n_725),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_SL g783 ( 
.A(n_630),
.B(n_401),
.Y(n_783)
);

NAND2x1p5_ASAP7_75t_L g784 ( 
.A(n_616),
.B(n_525),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_689),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_L g786 ( 
.A(n_628),
.B(n_598),
.Y(n_786)
);

INVx2_ASAP7_75t_L g787 ( 
.A(n_634),
.Y(n_787)
);

NAND2x1_ASAP7_75t_L g788 ( 
.A(n_615),
.B(n_535),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_689),
.Y(n_789)
);

INVx2_ASAP7_75t_L g790 ( 
.A(n_634),
.Y(n_790)
);

NOR2xp67_ASAP7_75t_L g791 ( 
.A(n_699),
.B(n_590),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_SL g792 ( 
.A(n_630),
.B(n_401),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_L g793 ( 
.A(n_688),
.B(n_598),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_726),
.Y(n_794)
);

NOR2xp33_ASAP7_75t_L g795 ( 
.A(n_713),
.B(n_602),
.Y(n_795)
);

AND2x2_ASAP7_75t_L g796 ( 
.A(n_693),
.B(n_460),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_SL g797 ( 
.A(n_630),
.B(n_283),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_688),
.B(n_598),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_SL g799 ( 
.A(n_616),
.B(n_283),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_L g800 ( 
.A(n_614),
.B(n_554),
.Y(n_800)
);

BUFx6f_ASAP7_75t_L g801 ( 
.A(n_617),
.Y(n_801)
);

INVx3_ASAP7_75t_L g802 ( 
.A(n_617),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_SL g803 ( 
.A(n_664),
.B(n_302),
.Y(n_803)
);

AND2x4_ASAP7_75t_SL g804 ( 
.A(n_738),
.B(n_692),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_SL g805 ( 
.A(n_642),
.B(n_302),
.Y(n_805)
);

INVx2_ASAP7_75t_L g806 ( 
.A(n_639),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_L g807 ( 
.A(n_614),
.B(n_554),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_SL g808 ( 
.A(n_693),
.B(n_707),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_L g809 ( 
.A(n_745),
.B(n_554),
.Y(n_809)
);

NOR2xp33_ASAP7_75t_L g810 ( 
.A(n_714),
.B(n_267),
.Y(n_810)
);

INVx2_ASAP7_75t_L g811 ( 
.A(n_639),
.Y(n_811)
);

INVx2_ASAP7_75t_SL g812 ( 
.A(n_636),
.Y(n_812)
);

AND2x4_ASAP7_75t_SL g813 ( 
.A(n_738),
.B(n_303),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_726),
.Y(n_814)
);

INVx2_ASAP7_75t_L g815 ( 
.A(n_640),
.Y(n_815)
);

OR2x2_ASAP7_75t_L g816 ( 
.A(n_717),
.B(n_269),
.Y(n_816)
);

NAND2x1_ASAP7_75t_L g817 ( 
.A(n_615),
.B(n_554),
.Y(n_817)
);

AND2x2_ASAP7_75t_L g818 ( 
.A(n_707),
.B(n_460),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_743),
.Y(n_819)
);

INVxp33_ASAP7_75t_L g820 ( 
.A(n_717),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_L g821 ( 
.A(n_745),
.B(n_560),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_743),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_L g823 ( 
.A(n_758),
.B(n_560),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_SL g824 ( 
.A(n_710),
.B(n_303),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_SL g825 ( 
.A(n_642),
.B(n_658),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_L g826 ( 
.A(n_758),
.B(n_560),
.Y(n_826)
);

AOI22xp5_ASAP7_75t_L g827 ( 
.A1(n_746),
.A2(n_250),
.B1(n_252),
.B2(n_239),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_757),
.Y(n_828)
);

NOR2xp33_ASAP7_75t_L g829 ( 
.A(n_672),
.B(n_280),
.Y(n_829)
);

BUFx3_ASAP7_75t_L g830 ( 
.A(n_724),
.Y(n_830)
);

INVx2_ASAP7_75t_L g831 ( 
.A(n_640),
.Y(n_831)
);

BUFx2_ASAP7_75t_L g832 ( 
.A(n_649),
.Y(n_832)
);

AND2x2_ASAP7_75t_L g833 ( 
.A(n_710),
.B(n_470),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_720),
.B(n_560),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_SL g835 ( 
.A(n_642),
.B(n_565),
.Y(n_835)
);

NOR2xp33_ASAP7_75t_L g836 ( 
.A(n_659),
.B(n_371),
.Y(n_836)
);

O2A1O1Ixp33_ASAP7_75t_L g837 ( 
.A1(n_643),
.A2(n_596),
.B(n_594),
.C(n_591),
.Y(n_837)
);

INVx2_ASAP7_75t_L g838 ( 
.A(n_641),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_L g839 ( 
.A(n_720),
.B(n_560),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_SL g840 ( 
.A(n_642),
.B(n_609),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_724),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_729),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_SL g843 ( 
.A(n_658),
.B(n_609),
.Y(n_843)
);

AND2x2_ASAP7_75t_L g844 ( 
.A(n_744),
.B(n_470),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_SL g845 ( 
.A(n_658),
.B(n_565),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_L g846 ( 
.A(n_694),
.B(n_565),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_L g847 ( 
.A(n_694),
.B(n_565),
.Y(n_847)
);

NOR2xp33_ASAP7_75t_L g848 ( 
.A(n_662),
.B(n_676),
.Y(n_848)
);

AOI22xp5_ASAP7_75t_L g849 ( 
.A1(n_746),
.A2(n_252),
.B1(n_253),
.B2(n_250),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_695),
.B(n_565),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_SL g851 ( 
.A(n_623),
.B(n_565),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_SL g852 ( 
.A(n_623),
.B(n_565),
.Y(n_852)
);

AND2x6_ASAP7_75t_L g853 ( 
.A(n_627),
.B(n_253),
.Y(n_853)
);

OAI22xp5_ASAP7_75t_L g854 ( 
.A1(n_620),
.A2(n_261),
.B1(n_262),
.B2(n_256),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_L g855 ( 
.A(n_695),
.B(n_565),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_SL g856 ( 
.A(n_627),
.B(n_582),
.Y(n_856)
);

INVx2_ASAP7_75t_L g857 ( 
.A(n_641),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_L g858 ( 
.A(n_696),
.B(n_582),
.Y(n_858)
);

OR2x6_ASAP7_75t_L g859 ( 
.A(n_738),
.B(n_478),
.Y(n_859)
);

NOR2xp33_ASAP7_75t_L g860 ( 
.A(n_741),
.B(n_213),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_L g861 ( 
.A(n_696),
.B(n_582),
.Y(n_861)
);

NOR2xp67_ASAP7_75t_L g862 ( 
.A(n_646),
.B(n_591),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_L g863 ( 
.A(n_701),
.B(n_582),
.Y(n_863)
);

INVxp67_ASAP7_75t_SL g864 ( 
.A(n_631),
.Y(n_864)
);

INVx2_ASAP7_75t_L g865 ( 
.A(n_648),
.Y(n_865)
);

NOR2xp33_ASAP7_75t_L g866 ( 
.A(n_612),
.B(n_736),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_SL g867 ( 
.A(n_631),
.B(n_582),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_SL g868 ( 
.A(n_632),
.B(n_582),
.Y(n_868)
);

OAI221xp5_ASAP7_75t_L g869 ( 
.A1(n_747),
.A2(n_478),
.B1(n_481),
.B2(n_510),
.C(n_372),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_SL g870 ( 
.A(n_632),
.B(n_582),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_L g871 ( 
.A(n_701),
.B(n_582),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_SL g872 ( 
.A(n_638),
.B(n_609),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_SL g873 ( 
.A(n_638),
.B(n_609),
.Y(n_873)
);

INVx2_ASAP7_75t_L g874 ( 
.A(n_648),
.Y(n_874)
);

A2O1A1Ixp33_ASAP7_75t_L g875 ( 
.A1(n_643),
.A2(n_534),
.B(n_525),
.C(n_261),
.Y(n_875)
);

NOR2xp33_ASAP7_75t_L g876 ( 
.A(n_661),
.B(n_670),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_L g877 ( 
.A(n_712),
.B(n_587),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_712),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_715),
.B(n_587),
.Y(n_879)
);

NAND2xp33_ASAP7_75t_L g880 ( 
.A(n_619),
.B(n_256),
.Y(n_880)
);

INVx1_ASAP7_75t_SL g881 ( 
.A(n_697),
.Y(n_881)
);

BUFx4_ASAP7_75t_L g882 ( 
.A(n_653),
.Y(n_882)
);

INVx5_ASAP7_75t_L g883 ( 
.A(n_677),
.Y(n_883)
);

HB1xp67_ASAP7_75t_L g884 ( 
.A(n_649),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_SL g885 ( 
.A(n_650),
.B(n_660),
.Y(n_885)
);

INVx2_ASAP7_75t_L g886 ( 
.A(n_654),
.Y(n_886)
);

NAND2xp33_ASAP7_75t_SL g887 ( 
.A(n_749),
.B(n_215),
.Y(n_887)
);

AND2x2_ASAP7_75t_L g888 ( 
.A(n_738),
.B(n_481),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_L g889 ( 
.A(n_715),
.B(n_587),
.Y(n_889)
);

AND2x4_ASAP7_75t_L g890 ( 
.A(n_731),
.B(n_594),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_SL g891 ( 
.A(n_666),
.B(n_338),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_716),
.Y(n_892)
);

INVxp67_ASAP7_75t_L g893 ( 
.A(n_666),
.Y(n_893)
);

INVx2_ASAP7_75t_L g894 ( 
.A(n_654),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_SL g895 ( 
.A(n_650),
.B(n_587),
.Y(n_895)
);

NOR2xp33_ASAP7_75t_SL g896 ( 
.A(n_624),
.B(n_338),
.Y(n_896)
);

NAND2x1_ASAP7_75t_L g897 ( 
.A(n_677),
.B(n_524),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_SL g898 ( 
.A(n_660),
.B(n_587),
.Y(n_898)
);

NOR2xp33_ASAP7_75t_L g899 ( 
.A(n_678),
.B(n_216),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_SL g900 ( 
.A(n_667),
.B(n_673),
.Y(n_900)
);

NOR2x1_ASAP7_75t_L g901 ( 
.A(n_637),
.B(n_262),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_L g902 ( 
.A(n_716),
.B(n_587),
.Y(n_902)
);

NOR2xp33_ASAP7_75t_L g903 ( 
.A(n_645),
.B(n_219),
.Y(n_903)
);

BUFx6f_ASAP7_75t_L g904 ( 
.A(n_677),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_718),
.Y(n_905)
);

INVxp33_ASAP7_75t_L g906 ( 
.A(n_728),
.Y(n_906)
);

BUFx8_ASAP7_75t_L g907 ( 
.A(n_731),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_L g908 ( 
.A(n_718),
.B(n_587),
.Y(n_908)
);

NOR2xp33_ASAP7_75t_L g909 ( 
.A(n_652),
.B(n_685),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_L g910 ( 
.A(n_722),
.B(n_587),
.Y(n_910)
);

BUFx3_ASAP7_75t_L g911 ( 
.A(n_677),
.Y(n_911)
);

NOR2xp33_ASAP7_75t_L g912 ( 
.A(n_621),
.B(n_221),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_SL g913 ( 
.A(n_667),
.B(n_673),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_SL g914 ( 
.A(n_731),
.B(n_609),
.Y(n_914)
);

OR2x2_ASAP7_75t_L g915 ( 
.A(n_748),
.B(n_510),
.Y(n_915)
);

BUFx3_ASAP7_75t_L g916 ( 
.A(n_677),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_L g917 ( 
.A(n_722),
.B(n_609),
.Y(n_917)
);

AND2x2_ASAP7_75t_L g918 ( 
.A(n_691),
.B(n_599),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_SL g919 ( 
.A(n_691),
.B(n_338),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_SL g920 ( 
.A(n_731),
.B(n_609),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_L g921 ( 
.A(n_730),
.B(n_609),
.Y(n_921)
);

INVx2_ASAP7_75t_L g922 ( 
.A(n_656),
.Y(n_922)
);

AOI22xp5_ASAP7_75t_L g923 ( 
.A1(n_746),
.A2(n_363),
.B1(n_273),
.B2(n_278),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_SL g924 ( 
.A(n_730),
.B(n_264),
.Y(n_924)
);

NOR2xp33_ASAP7_75t_L g925 ( 
.A(n_621),
.B(n_231),
.Y(n_925)
);

AOI22xp33_ASAP7_75t_L g926 ( 
.A1(n_619),
.A2(n_394),
.B1(n_273),
.B2(n_278),
.Y(n_926)
);

OAI22xp33_ASAP7_75t_L g927 ( 
.A1(n_621),
.A2(n_651),
.B1(n_746),
.B2(n_686),
.Y(n_927)
);

AOI22xp5_ASAP7_75t_L g928 ( 
.A1(n_619),
.A2(n_313),
.B1(n_410),
.B2(n_394),
.Y(n_928)
);

AOI22xp5_ASAP7_75t_L g929 ( 
.A1(n_619),
.A2(n_363),
.B1(n_281),
.B2(n_289),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_739),
.B(n_740),
.Y(n_930)
);

OAI22xp5_ASAP7_75t_SL g931 ( 
.A1(n_728),
.A2(n_312),
.B1(n_296),
.B2(n_292),
.Y(n_931)
);

NOR2xp67_ASAP7_75t_L g932 ( 
.A(n_624),
.B(n_599),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_L g933 ( 
.A(n_764),
.B(n_739),
.Y(n_933)
);

AOI22xp5_ASAP7_75t_L g934 ( 
.A1(n_782),
.A2(n_619),
.B1(n_677),
.B2(n_651),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_SL g935 ( 
.A(n_927),
.B(n_740),
.Y(n_935)
);

CKINVDCx5p33_ASAP7_75t_R g936 ( 
.A(n_881),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_L g937 ( 
.A(n_808),
.B(n_753),
.Y(n_937)
);

AOI21xp5_ASAP7_75t_L g938 ( 
.A1(n_825),
.A2(n_711),
.B(n_635),
.Y(n_938)
);

HB1xp67_ASAP7_75t_L g939 ( 
.A(n_771),
.Y(n_939)
);

AOI21xp5_ASAP7_75t_L g940 ( 
.A1(n_825),
.A2(n_711),
.B(n_635),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_L g941 ( 
.A(n_864),
.B(n_753),
.Y(n_941)
);

AOI21xp5_ASAP7_75t_L g942 ( 
.A1(n_883),
.A2(n_711),
.B(n_635),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_L g943 ( 
.A(n_810),
.B(n_760),
.Y(n_943)
);

AOI22xp5_ASAP7_75t_L g944 ( 
.A1(n_876),
.A2(n_619),
.B1(n_677),
.B2(n_651),
.Y(n_944)
);

AOI21xp5_ASAP7_75t_L g945 ( 
.A1(n_883),
.A2(n_635),
.B(n_626),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_L g946 ( 
.A(n_829),
.B(n_760),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_L g947 ( 
.A(n_796),
.B(n_686),
.Y(n_947)
);

AOI21xp5_ASAP7_75t_L g948 ( 
.A1(n_883),
.A2(n_635),
.B(n_626),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_L g949 ( 
.A(n_818),
.B(n_686),
.Y(n_949)
);

AND2x2_ASAP7_75t_L g950 ( 
.A(n_833),
.B(n_683),
.Y(n_950)
);

INVxp67_ASAP7_75t_L g951 ( 
.A(n_844),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_SL g952 ( 
.A(n_883),
.B(n_674),
.Y(n_952)
);

AOI21xp5_ASAP7_75t_L g953 ( 
.A1(n_767),
.A2(n_644),
.B(n_626),
.Y(n_953)
);

AND2x4_ASAP7_75t_L g954 ( 
.A(n_830),
.B(n_637),
.Y(n_954)
);

AO21x1_ASAP7_75t_L g955 ( 
.A1(n_797),
.A2(n_680),
.B(n_679),
.Y(n_955)
);

NOR2xp33_ASAP7_75t_L g956 ( 
.A(n_893),
.B(n_621),
.Y(n_956)
);

O2A1O1Ixp33_ASAP7_75t_L g957 ( 
.A1(n_803),
.A2(n_686),
.B(n_651),
.C(n_742),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_L g958 ( 
.A(n_878),
.B(n_892),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_SL g959 ( 
.A(n_904),
.B(n_674),
.Y(n_959)
);

INVx3_ASAP7_75t_L g960 ( 
.A(n_890),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_L g961 ( 
.A(n_905),
.B(n_686),
.Y(n_961)
);

INVx2_ASAP7_75t_L g962 ( 
.A(n_766),
.Y(n_962)
);

AOI21xp5_ASAP7_75t_L g963 ( 
.A1(n_770),
.A2(n_644),
.B(n_626),
.Y(n_963)
);

O2A1O1Ixp33_ASAP7_75t_L g964 ( 
.A1(n_803),
.A2(n_761),
.B(n_759),
.C(n_681),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_L g965 ( 
.A(n_830),
.B(n_619),
.Y(n_965)
);

AND2x4_ASAP7_75t_L g966 ( 
.A(n_785),
.B(n_656),
.Y(n_966)
);

AOI22xp5_ASAP7_75t_L g967 ( 
.A1(n_795),
.A2(n_681),
.B1(n_684),
.B2(n_679),
.Y(n_967)
);

INVx2_ASAP7_75t_L g968 ( 
.A(n_766),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_774),
.Y(n_969)
);

O2A1O1Ixp33_ASAP7_75t_L g970 ( 
.A1(n_924),
.A2(n_684),
.B(n_668),
.C(n_669),
.Y(n_970)
);

INVx3_ASAP7_75t_L g971 ( 
.A(n_890),
.Y(n_971)
);

OAI22xp5_ASAP7_75t_L g972 ( 
.A1(n_909),
.A2(n_752),
.B1(n_668),
.B2(n_669),
.Y(n_972)
);

BUFx2_ASAP7_75t_L g973 ( 
.A(n_832),
.Y(n_973)
);

NOR3xp33_ASAP7_75t_L g974 ( 
.A(n_763),
.B(n_683),
.C(n_603),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_L g975 ( 
.A(n_777),
.B(n_665),
.Y(n_975)
);

AO21x1_ASAP7_75t_L g976 ( 
.A1(n_797),
.A2(n_680),
.B(n_281),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_L g977 ( 
.A(n_834),
.B(n_665),
.Y(n_977)
);

OR2x2_ASAP7_75t_SL g978 ( 
.A(n_915),
.B(n_386),
.Y(n_978)
);

OAI21xp5_ASAP7_75t_L g979 ( 
.A1(n_783),
.A2(n_737),
.B(n_534),
.Y(n_979)
);

AOI21xp5_ASAP7_75t_L g980 ( 
.A1(n_773),
.A2(n_644),
.B(n_626),
.Y(n_980)
);

AOI21x1_ASAP7_75t_L g981 ( 
.A1(n_783),
.A2(n_682),
.B(n_675),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_L g982 ( 
.A(n_839),
.B(n_930),
.Y(n_982)
);

NOR2xp33_ASAP7_75t_L g983 ( 
.A(n_812),
.B(n_675),
.Y(n_983)
);

INVx2_ASAP7_75t_L g984 ( 
.A(n_774),
.Y(n_984)
);

AND2x2_ASAP7_75t_L g985 ( 
.A(n_836),
.B(n_888),
.Y(n_985)
);

AOI21xp5_ASAP7_75t_L g986 ( 
.A1(n_775),
.A2(n_727),
.B(n_644),
.Y(n_986)
);

OAI22xp5_ASAP7_75t_L g987 ( 
.A1(n_911),
.A2(n_682),
.B1(n_289),
.B2(n_299),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_SL g988 ( 
.A(n_904),
.B(n_644),
.Y(n_988)
);

AOI21xp5_ASAP7_75t_L g989 ( 
.A1(n_843),
.A2(n_727),
.B(n_756),
.Y(n_989)
);

INVx2_ASAP7_75t_L g990 ( 
.A(n_787),
.Y(n_990)
);

AND2x2_ASAP7_75t_L g991 ( 
.A(n_816),
.B(n_600),
.Y(n_991)
);

INVxp67_ASAP7_75t_L g992 ( 
.A(n_884),
.Y(n_992)
);

AOI21xp5_ASAP7_75t_L g993 ( 
.A1(n_843),
.A2(n_727),
.B(n_756),
.Y(n_993)
);

AOI21xp5_ASAP7_75t_L g994 ( 
.A1(n_845),
.A2(n_727),
.B(n_756),
.Y(n_994)
);

AOI22xp33_ASAP7_75t_L g995 ( 
.A1(n_853),
.A2(n_900),
.B1(n_913),
.B2(n_885),
.Y(n_995)
);

AND2x2_ASAP7_75t_L g996 ( 
.A(n_820),
.B(n_600),
.Y(n_996)
);

BUFx6f_ASAP7_75t_L g997 ( 
.A(n_904),
.Y(n_997)
);

AND2x2_ASAP7_75t_L g998 ( 
.A(n_918),
.B(n_603),
.Y(n_998)
);

A2O1A1Ixp33_ASAP7_75t_L g999 ( 
.A1(n_866),
.A2(n_395),
.B(n_397),
.C(n_393),
.Y(n_999)
);

AOI21xp5_ASAP7_75t_L g1000 ( 
.A1(n_845),
.A2(n_727),
.B(n_702),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_L g1001 ( 
.A(n_768),
.B(n_769),
.Y(n_1001)
);

BUFx2_ASAP7_75t_L g1002 ( 
.A(n_859),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_L g1003 ( 
.A(n_841),
.B(n_647),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_L g1004 ( 
.A(n_842),
.B(n_647),
.Y(n_1004)
);

HB1xp67_ASAP7_75t_L g1005 ( 
.A(n_789),
.Y(n_1005)
);

OAI22xp5_ASAP7_75t_L g1006 ( 
.A1(n_911),
.A2(n_299),
.B1(n_309),
.B2(n_264),
.Y(n_1006)
);

NAND2xp33_ASAP7_75t_L g1007 ( 
.A(n_776),
.B(n_732),
.Y(n_1007)
);

INVx3_ASAP7_75t_L g1008 ( 
.A(n_890),
.Y(n_1008)
);

BUFx6f_ASAP7_75t_L g1009 ( 
.A(n_904),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_SL g1010 ( 
.A(n_776),
.B(n_801),
.Y(n_1010)
);

OAI21x1_ASAP7_75t_L g1011 ( 
.A1(n_817),
.A2(n_655),
.B(n_647),
.Y(n_1011)
);

NAND2x1_ASAP7_75t_L g1012 ( 
.A(n_776),
.B(n_751),
.Y(n_1012)
);

AOI21xp5_ASAP7_75t_L g1013 ( 
.A1(n_792),
.A2(n_702),
.B(n_690),
.Y(n_1013)
);

OAI21xp5_ASAP7_75t_L g1014 ( 
.A1(n_792),
.A2(n_534),
.B(n_525),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_SL g1015 ( 
.A(n_776),
.B(n_655),
.Y(n_1015)
);

A2O1A1Ixp33_ASAP7_75t_L g1016 ( 
.A1(n_912),
.A2(n_395),
.B(n_397),
.C(n_393),
.Y(n_1016)
);

AOI21xp33_ASAP7_75t_L g1017 ( 
.A1(n_903),
.A2(n_313),
.B(n_309),
.Y(n_1017)
);

OAI21xp5_ASAP7_75t_L g1018 ( 
.A1(n_885),
.A2(n_709),
.B(n_655),
.Y(n_1018)
);

AND2x2_ASAP7_75t_L g1019 ( 
.A(n_932),
.B(n_604),
.Y(n_1019)
);

AOI21xp5_ASAP7_75t_L g1020 ( 
.A1(n_835),
.A2(n_703),
.B(n_690),
.Y(n_1020)
);

NOR2x1_ASAP7_75t_R g1021 ( 
.A(n_919),
.B(n_233),
.Y(n_1021)
);

OAI21xp5_ASAP7_75t_L g1022 ( 
.A1(n_900),
.A2(n_709),
.B(n_704),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_SL g1023 ( 
.A(n_801),
.B(n_703),
.Y(n_1023)
);

A2O1A1Ixp33_ASAP7_75t_L g1024 ( 
.A1(n_925),
.A2(n_404),
.B(n_406),
.C(n_409),
.Y(n_1024)
);

OAI21xp33_ASAP7_75t_L g1025 ( 
.A1(n_896),
.A2(n_242),
.B(n_234),
.Y(n_1025)
);

INVx1_ASAP7_75t_L g1026 ( 
.A(n_790),
.Y(n_1026)
);

INVx2_ASAP7_75t_L g1027 ( 
.A(n_790),
.Y(n_1027)
);

OAI21xp33_ASAP7_75t_L g1028 ( 
.A1(n_860),
.A2(n_247),
.B(n_243),
.Y(n_1028)
);

AOI21x1_ASAP7_75t_L g1029 ( 
.A1(n_895),
.A2(n_708),
.B(n_705),
.Y(n_1029)
);

AOI33xp33_ASAP7_75t_L g1030 ( 
.A1(n_804),
.A2(n_506),
.A3(n_513),
.B1(n_516),
.B2(n_520),
.B3(n_521),
.Y(n_1030)
);

NOR2xp33_ASAP7_75t_L g1031 ( 
.A(n_848),
.B(n_258),
.Y(n_1031)
);

INVx1_ASAP7_75t_L g1032 ( 
.A(n_806),
.Y(n_1032)
);

AO21x1_ASAP7_75t_L g1033 ( 
.A1(n_799),
.A2(n_345),
.B(n_341),
.Y(n_1033)
);

OAI21xp5_ASAP7_75t_L g1034 ( 
.A1(n_913),
.A2(n_852),
.B(n_851),
.Y(n_1034)
);

OAI21xp33_ASAP7_75t_L g1035 ( 
.A1(n_899),
.A2(n_274),
.B(n_260),
.Y(n_1035)
);

BUFx4f_ASAP7_75t_L g1036 ( 
.A(n_859),
.Y(n_1036)
);

AOI21xp5_ASAP7_75t_L g1037 ( 
.A1(n_835),
.A2(n_708),
.B(n_705),
.Y(n_1037)
);

O2A1O1Ixp5_ASAP7_75t_L g1038 ( 
.A1(n_799),
.A2(n_805),
.B(n_772),
.C(n_924),
.Y(n_1038)
);

NOR2xp67_ASAP7_75t_L g1039 ( 
.A(n_778),
.B(n_604),
.Y(n_1039)
);

INVx2_ASAP7_75t_L g1040 ( 
.A(n_806),
.Y(n_1040)
);

AOI21xp5_ASAP7_75t_L g1041 ( 
.A1(n_840),
.A2(n_723),
.B(n_721),
.Y(n_1041)
);

AOI21xp5_ASAP7_75t_L g1042 ( 
.A1(n_840),
.A2(n_723),
.B(n_721),
.Y(n_1042)
);

NAND2xp5_ASAP7_75t_L g1043 ( 
.A(n_828),
.B(n_735),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_L g1044 ( 
.A(n_781),
.B(n_735),
.Y(n_1044)
);

O2A1O1Ixp33_ASAP7_75t_L g1045 ( 
.A1(n_854),
.A2(n_346),
.B(n_391),
.C(n_390),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_L g1046 ( 
.A(n_786),
.B(n_750),
.Y(n_1046)
);

AOI21xp5_ASAP7_75t_L g1047 ( 
.A1(n_851),
.A2(n_754),
.B(n_750),
.Y(n_1047)
);

AOI21xp5_ASAP7_75t_L g1048 ( 
.A1(n_852),
.A2(n_755),
.B(n_754),
.Y(n_1048)
);

NAND2xp5_ASAP7_75t_L g1049 ( 
.A(n_793),
.B(n_755),
.Y(n_1049)
);

A2O1A1Ixp33_ASAP7_75t_L g1050 ( 
.A1(n_869),
.A2(n_404),
.B(n_406),
.C(n_409),
.Y(n_1050)
);

AND2x2_ASAP7_75t_L g1051 ( 
.A(n_859),
.B(n_606),
.Y(n_1051)
);

BUFx6f_ASAP7_75t_L g1052 ( 
.A(n_801),
.Y(n_1052)
);

AOI21xp5_ASAP7_75t_L g1053 ( 
.A1(n_856),
.A2(n_762),
.B(n_734),
.Y(n_1053)
);

O2A1O1Ixp33_ASAP7_75t_L g1054 ( 
.A1(n_805),
.A2(n_346),
.B(n_341),
.C(n_345),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_L g1055 ( 
.A(n_798),
.B(n_611),
.Y(n_1055)
);

NAND2xp5_ASAP7_75t_L g1056 ( 
.A(n_862),
.B(n_611),
.Y(n_1056)
);

BUFx6f_ASAP7_75t_L g1057 ( 
.A(n_801),
.Y(n_1057)
);

O2A1O1Ixp33_ASAP7_75t_L g1058 ( 
.A1(n_824),
.A2(n_366),
.B(n_357),
.C(n_390),
.Y(n_1058)
);

AND2x4_ASAP7_75t_L g1059 ( 
.A(n_791),
.B(n_606),
.Y(n_1059)
);

BUFx4f_ASAP7_75t_L g1060 ( 
.A(n_853),
.Y(n_1060)
);

AOI21xp5_ASAP7_75t_L g1061 ( 
.A1(n_867),
.A2(n_734),
.B(n_618),
.Y(n_1061)
);

AOI21xp5_ASAP7_75t_L g1062 ( 
.A1(n_867),
.A2(n_734),
.B(n_618),
.Y(n_1062)
);

NOR2xp33_ASAP7_75t_L g1063 ( 
.A(n_891),
.B(n_275),
.Y(n_1063)
);

AOI21xp5_ASAP7_75t_L g1064 ( 
.A1(n_868),
.A2(n_734),
.B(n_625),
.Y(n_1064)
);

INVxp67_ASAP7_75t_L g1065 ( 
.A(n_901),
.Y(n_1065)
);

AOI21xp5_ASAP7_75t_L g1066 ( 
.A1(n_868),
.A2(n_734),
.B(n_625),
.Y(n_1066)
);

NAND2xp5_ASAP7_75t_L g1067 ( 
.A(n_794),
.B(n_814),
.Y(n_1067)
);

AOI21xp5_ASAP7_75t_L g1068 ( 
.A1(n_870),
.A2(n_613),
.B(n_545),
.Y(n_1068)
);

AOI22xp33_ASAP7_75t_L g1069 ( 
.A1(n_853),
.A2(n_410),
.B1(n_356),
.B2(n_354),
.Y(n_1069)
);

INVx4_ASAP7_75t_L g1070 ( 
.A(n_765),
.Y(n_1070)
);

CKINVDCx20_ASAP7_75t_R g1071 ( 
.A(n_779),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_L g1072 ( 
.A(n_819),
.B(n_613),
.Y(n_1072)
);

OAI22xp5_ASAP7_75t_L g1073 ( 
.A1(n_916),
.A2(n_357),
.B1(n_349),
.B2(n_354),
.Y(n_1073)
);

INVx2_ASAP7_75t_L g1074 ( 
.A(n_811),
.Y(n_1074)
);

NAND2xp5_ASAP7_75t_L g1075 ( 
.A(n_822),
.B(n_348),
.Y(n_1075)
);

NAND2xp5_ASAP7_75t_L g1076 ( 
.A(n_815),
.B(n_348),
.Y(n_1076)
);

INVx4_ASAP7_75t_L g1077 ( 
.A(n_765),
.Y(n_1077)
);

NOR2xp33_ASAP7_75t_L g1078 ( 
.A(n_813),
.B(n_282),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_L g1079 ( 
.A(n_815),
.B(n_349),
.Y(n_1079)
);

NAND2xp5_ASAP7_75t_L g1080 ( 
.A(n_831),
.B(n_356),
.Y(n_1080)
);

BUFx6f_ASAP7_75t_L g1081 ( 
.A(n_916),
.Y(n_1081)
);

NAND2xp5_ASAP7_75t_L g1082 ( 
.A(n_831),
.B(n_838),
.Y(n_1082)
);

NAND2xp5_ASAP7_75t_L g1083 ( 
.A(n_838),
.B(n_366),
.Y(n_1083)
);

INVx1_ASAP7_75t_L g1084 ( 
.A(n_857),
.Y(n_1084)
);

OAI21xp5_ASAP7_75t_L g1085 ( 
.A1(n_872),
.A2(n_733),
.B(n_732),
.Y(n_1085)
);

NAND2xp5_ASAP7_75t_SL g1086 ( 
.A(n_802),
.B(n_391),
.Y(n_1086)
);

NAND2xp5_ASAP7_75t_L g1087 ( 
.A(n_857),
.B(n_732),
.Y(n_1087)
);

INVx2_ASAP7_75t_L g1088 ( 
.A(n_865),
.Y(n_1088)
);

NAND2xp5_ASAP7_75t_L g1089 ( 
.A(n_865),
.B(n_732),
.Y(n_1089)
);

NAND2xp5_ASAP7_75t_L g1090 ( 
.A(n_874),
.B(n_732),
.Y(n_1090)
);

AOI21x1_ASAP7_75t_L g1091 ( 
.A1(n_895),
.A2(n_526),
.B(n_524),
.Y(n_1091)
);

AOI21xp5_ASAP7_75t_L g1092 ( 
.A1(n_872),
.A2(n_545),
.B(n_544),
.Y(n_1092)
);

AOI21xp5_ASAP7_75t_L g1093 ( 
.A1(n_873),
.A2(n_545),
.B(n_544),
.Y(n_1093)
);

AOI21x1_ASAP7_75t_L g1094 ( 
.A1(n_898),
.A2(n_526),
.B(n_524),
.Y(n_1094)
);

NOR2xp33_ASAP7_75t_L g1095 ( 
.A(n_813),
.B(n_291),
.Y(n_1095)
);

AOI21xp5_ASAP7_75t_L g1096 ( 
.A1(n_873),
.A2(n_547),
.B(n_545),
.Y(n_1096)
);

INVx3_ASAP7_75t_L g1097 ( 
.A(n_874),
.Y(n_1097)
);

BUFx4f_ASAP7_75t_L g1098 ( 
.A(n_853),
.Y(n_1098)
);

NAND2xp5_ASAP7_75t_L g1099 ( 
.A(n_886),
.B(n_733),
.Y(n_1099)
);

NAND2xp5_ASAP7_75t_L g1100 ( 
.A(n_886),
.B(n_733),
.Y(n_1100)
);

NAND2xp5_ASAP7_75t_L g1101 ( 
.A(n_894),
.B(n_733),
.Y(n_1101)
);

OAI321xp33_ASAP7_75t_L g1102 ( 
.A1(n_931),
.A2(n_516),
.A3(n_520),
.B1(n_521),
.B2(n_522),
.C(n_506),
.Y(n_1102)
);

INVx2_ASAP7_75t_L g1103 ( 
.A(n_894),
.Y(n_1103)
);

CKINVDCx10_ASAP7_75t_R g1104 ( 
.A(n_882),
.Y(n_1104)
);

NAND2xp5_ASAP7_75t_L g1105 ( 
.A(n_922),
.B(n_802),
.Y(n_1105)
);

AOI21x1_ASAP7_75t_L g1106 ( 
.A1(n_788),
.A2(n_526),
.B(n_524),
.Y(n_1106)
);

NAND2xp5_ASAP7_75t_L g1107 ( 
.A(n_922),
.B(n_733),
.Y(n_1107)
);

O2A1O1Ixp33_ASAP7_75t_L g1108 ( 
.A1(n_837),
.A2(n_608),
.B(n_607),
.C(n_513),
.Y(n_1108)
);

INVx1_ASAP7_75t_L g1109 ( 
.A(n_846),
.Y(n_1109)
);

BUFx3_ASAP7_75t_L g1110 ( 
.A(n_907),
.Y(n_1110)
);

OAI21x1_ASAP7_75t_L g1111 ( 
.A1(n_784),
.A2(n_527),
.B(n_526),
.Y(n_1111)
);

A2O1A1Ixp33_ASAP7_75t_L g1112 ( 
.A1(n_827),
.A2(n_607),
.B(n_608),
.C(n_512),
.Y(n_1112)
);

OAI21xp5_ASAP7_75t_L g1113 ( 
.A1(n_800),
.A2(n_528),
.B(n_527),
.Y(n_1113)
);

AOI21xp5_ASAP7_75t_L g1114 ( 
.A1(n_807),
.A2(n_547),
.B(n_545),
.Y(n_1114)
);

INVx4_ASAP7_75t_L g1115 ( 
.A(n_853),
.Y(n_1115)
);

NAND2xp5_ASAP7_75t_L g1116 ( 
.A(n_849),
.B(n_751),
.Y(n_1116)
);

NOR2xp33_ASAP7_75t_L g1117 ( 
.A(n_923),
.B(n_304),
.Y(n_1117)
);

NAND2xp33_ASAP7_75t_SL g1118 ( 
.A(n_950),
.B(n_906),
.Y(n_1118)
);

NAND2xp5_ASAP7_75t_SL g1119 ( 
.A(n_944),
.B(n_780),
.Y(n_1119)
);

NAND2xp5_ASAP7_75t_SL g1120 ( 
.A(n_934),
.B(n_784),
.Y(n_1120)
);

OAI22xp5_ASAP7_75t_L g1121 ( 
.A1(n_995),
.A2(n_926),
.B1(n_929),
.B2(n_928),
.Y(n_1121)
);

CKINVDCx6p67_ASAP7_75t_R g1122 ( 
.A(n_1104),
.Y(n_1122)
);

NAND2xp5_ASAP7_75t_L g1123 ( 
.A(n_943),
.B(n_809),
.Y(n_1123)
);

INVx3_ASAP7_75t_L g1124 ( 
.A(n_1052),
.Y(n_1124)
);

A2O1A1Ixp33_ASAP7_75t_L g1125 ( 
.A1(n_1031),
.A2(n_887),
.B(n_880),
.C(n_875),
.Y(n_1125)
);

INVxp67_ASAP7_75t_SL g1126 ( 
.A(n_1052),
.Y(n_1126)
);

CKINVDCx10_ASAP7_75t_R g1127 ( 
.A(n_936),
.Y(n_1127)
);

AOI21xp5_ASAP7_75t_L g1128 ( 
.A1(n_982),
.A2(n_920),
.B(n_914),
.Y(n_1128)
);

OR2x2_ASAP7_75t_L g1129 ( 
.A(n_951),
.B(n_772),
.Y(n_1129)
);

AND2x2_ASAP7_75t_L g1130 ( 
.A(n_985),
.B(n_355),
.Y(n_1130)
);

AOI22xp5_ASAP7_75t_L g1131 ( 
.A1(n_1071),
.A2(n_907),
.B1(n_920),
.B2(n_914),
.Y(n_1131)
);

AOI21xp5_ASAP7_75t_L g1132 ( 
.A1(n_975),
.A2(n_897),
.B(n_823),
.Y(n_1132)
);

OAI22xp5_ASAP7_75t_L g1133 ( 
.A1(n_995),
.A2(n_821),
.B1(n_826),
.B2(n_910),
.Y(n_1133)
);

INVx1_ASAP7_75t_L g1134 ( 
.A(n_1005),
.Y(n_1134)
);

BUFx12f_ASAP7_75t_L g1135 ( 
.A(n_973),
.Y(n_1135)
);

HB1xp67_ASAP7_75t_L g1136 ( 
.A(n_939),
.Y(n_1136)
);

AOI21xp5_ASAP7_75t_L g1137 ( 
.A1(n_933),
.A2(n_850),
.B(n_847),
.Y(n_1137)
);

O2A1O1Ixp33_ASAP7_75t_SL g1138 ( 
.A1(n_1017),
.A2(n_921),
.B(n_917),
.C(n_908),
.Y(n_1138)
);

INVx2_ASAP7_75t_L g1139 ( 
.A(n_1097),
.Y(n_1139)
);

NAND2xp5_ASAP7_75t_SL g1140 ( 
.A(n_960),
.B(n_855),
.Y(n_1140)
);

NAND2xp5_ASAP7_75t_L g1141 ( 
.A(n_946),
.B(n_858),
.Y(n_1141)
);

AOI21xp5_ASAP7_75t_L g1142 ( 
.A1(n_977),
.A2(n_863),
.B(n_861),
.Y(n_1142)
);

INVx1_ASAP7_75t_L g1143 ( 
.A(n_1005),
.Y(n_1143)
);

INVx2_ASAP7_75t_L g1144 ( 
.A(n_1097),
.Y(n_1144)
);

INVx1_ASAP7_75t_L g1145 ( 
.A(n_969),
.Y(n_1145)
);

BUFx6f_ASAP7_75t_L g1146 ( 
.A(n_1052),
.Y(n_1146)
);

NAND2xp5_ASAP7_75t_L g1147 ( 
.A(n_998),
.B(n_1019),
.Y(n_1147)
);

AND2x2_ASAP7_75t_L g1148 ( 
.A(n_991),
.B(n_355),
.Y(n_1148)
);

A2O1A1Ixp33_ASAP7_75t_L g1149 ( 
.A1(n_1117),
.A2(n_871),
.B(n_902),
.C(n_889),
.Y(n_1149)
);

BUFx12f_ASAP7_75t_L g1150 ( 
.A(n_1110),
.Y(n_1150)
);

AOI33xp33_ASAP7_75t_L g1151 ( 
.A1(n_996),
.A2(n_522),
.A3(n_512),
.B1(n_509),
.B2(n_507),
.B3(n_458),
.Y(n_1151)
);

OAI22xp5_ASAP7_75t_L g1152 ( 
.A1(n_1081),
.A2(n_879),
.B1(n_877),
.B2(n_751),
.Y(n_1152)
);

NAND2xp5_ASAP7_75t_L g1153 ( 
.A(n_947),
.B(n_907),
.Y(n_1153)
);

OR2x2_ASAP7_75t_L g1154 ( 
.A(n_992),
.B(n_507),
.Y(n_1154)
);

OAI22xp5_ASAP7_75t_L g1155 ( 
.A1(n_1081),
.A2(n_751),
.B1(n_376),
.B2(n_375),
.Y(n_1155)
);

NAND3xp33_ASAP7_75t_SL g1156 ( 
.A(n_1028),
.B(n_369),
.C(n_315),
.Y(n_1156)
);

INVx1_ASAP7_75t_L g1157 ( 
.A(n_1026),
.Y(n_1157)
);

NAND2xp5_ASAP7_75t_L g1158 ( 
.A(n_949),
.B(n_958),
.Y(n_1158)
);

AOI21xp5_ASAP7_75t_L g1159 ( 
.A1(n_953),
.A2(n_963),
.B(n_980),
.Y(n_1159)
);

INVx5_ASAP7_75t_L g1160 ( 
.A(n_1052),
.Y(n_1160)
);

INVx1_ASAP7_75t_L g1161 ( 
.A(n_1032),
.Y(n_1161)
);

BUFx3_ASAP7_75t_L g1162 ( 
.A(n_939),
.Y(n_1162)
);

AOI21xp5_ASAP7_75t_L g1163 ( 
.A1(n_986),
.A2(n_549),
.B(n_545),
.Y(n_1163)
);

A2O1A1Ixp33_ASAP7_75t_L g1164 ( 
.A1(n_1050),
.A2(n_509),
.B(n_310),
.C(n_367),
.Y(n_1164)
);

INVx1_ASAP7_75t_L g1165 ( 
.A(n_1084),
.Y(n_1165)
);

INVx1_ASAP7_75t_L g1166 ( 
.A(n_962),
.Y(n_1166)
);

AND2x2_ASAP7_75t_L g1167 ( 
.A(n_1051),
.B(n_355),
.Y(n_1167)
);

A2O1A1Ixp33_ASAP7_75t_L g1168 ( 
.A1(n_1050),
.A2(n_377),
.B(n_317),
.C(n_318),
.Y(n_1168)
);

OAI22xp5_ASAP7_75t_L g1169 ( 
.A1(n_1081),
.A2(n_385),
.B1(n_319),
.B2(n_320),
.Y(n_1169)
);

INVx2_ASAP7_75t_L g1170 ( 
.A(n_968),
.Y(n_1170)
);

NAND2xp5_ASAP7_75t_SL g1171 ( 
.A(n_960),
.B(n_338),
.Y(n_1171)
);

O2A1O1Ixp33_ASAP7_75t_L g1172 ( 
.A1(n_1102),
.A2(n_458),
.B(n_588),
.C(n_575),
.Y(n_1172)
);

BUFx4f_ASAP7_75t_L g1173 ( 
.A(n_954),
.Y(n_1173)
);

INVxp67_ASAP7_75t_L g1174 ( 
.A(n_983),
.Y(n_1174)
);

OAI22xp5_ASAP7_75t_L g1175 ( 
.A1(n_1081),
.A2(n_398),
.B1(n_328),
.B2(n_330),
.Y(n_1175)
);

O2A1O1Ixp33_ASAP7_75t_L g1176 ( 
.A1(n_1016),
.A2(n_588),
.B(n_575),
.C(n_574),
.Y(n_1176)
);

CKINVDCx5p33_ASAP7_75t_R g1177 ( 
.A(n_1002),
.Y(n_1177)
);

AND2x2_ASAP7_75t_L g1178 ( 
.A(n_1063),
.B(n_1117),
.Y(n_1178)
);

AOI21x1_ASAP7_75t_L g1179 ( 
.A1(n_1023),
.A2(n_528),
.B(n_527),
.Y(n_1179)
);

AOI21xp5_ASAP7_75t_L g1180 ( 
.A1(n_965),
.A2(n_545),
.B(n_547),
.Y(n_1180)
);

CKINVDCx14_ASAP7_75t_R g1181 ( 
.A(n_1036),
.Y(n_1181)
);

INVx2_ASAP7_75t_L g1182 ( 
.A(n_984),
.Y(n_1182)
);

NAND2xp5_ASAP7_75t_L g1183 ( 
.A(n_983),
.B(n_571),
.Y(n_1183)
);

NAND2xp5_ASAP7_75t_SL g1184 ( 
.A(n_971),
.B(n_350),
.Y(n_1184)
);

NAND2xp5_ASAP7_75t_L g1185 ( 
.A(n_937),
.B(n_571),
.Y(n_1185)
);

CKINVDCx8_ASAP7_75t_R g1186 ( 
.A(n_954),
.Y(n_1186)
);

AOI21xp5_ASAP7_75t_L g1187 ( 
.A1(n_942),
.A2(n_988),
.B(n_1105),
.Y(n_1187)
);

BUFx4f_ASAP7_75t_L g1188 ( 
.A(n_1057),
.Y(n_1188)
);

INVx1_ASAP7_75t_L g1189 ( 
.A(n_990),
.Y(n_1189)
);

NAND2xp5_ASAP7_75t_SL g1190 ( 
.A(n_971),
.B(n_350),
.Y(n_1190)
);

CKINVDCx8_ASAP7_75t_R g1191 ( 
.A(n_1057),
.Y(n_1191)
);

AOI21xp5_ASAP7_75t_L g1192 ( 
.A1(n_988),
.A2(n_979),
.B(n_940),
.Y(n_1192)
);

A2O1A1Ixp33_ASAP7_75t_L g1193 ( 
.A1(n_1016),
.A2(n_384),
.B(n_331),
.C(n_332),
.Y(n_1193)
);

AOI21xp5_ASAP7_75t_L g1194 ( 
.A1(n_938),
.A2(n_545),
.B(n_547),
.Y(n_1194)
);

A2O1A1Ixp33_ASAP7_75t_L g1195 ( 
.A1(n_1024),
.A2(n_402),
.B(n_335),
.C(n_337),
.Y(n_1195)
);

INVx4_ASAP7_75t_L g1196 ( 
.A(n_1057),
.Y(n_1196)
);

OAI22x1_ASAP7_75t_L g1197 ( 
.A1(n_1063),
.A2(n_316),
.B1(n_340),
.B2(n_343),
.Y(n_1197)
);

AOI22xp33_ASAP7_75t_L g1198 ( 
.A1(n_1069),
.A2(n_361),
.B1(n_388),
.B2(n_413),
.Y(n_1198)
);

OAI22xp5_ASAP7_75t_L g1199 ( 
.A1(n_967),
.A2(n_373),
.B1(n_383),
.B2(n_403),
.Y(n_1199)
);

HB1xp67_ASAP7_75t_L g1200 ( 
.A(n_1008),
.Y(n_1200)
);

NAND2xp5_ASAP7_75t_SL g1201 ( 
.A(n_1008),
.B(n_350),
.Y(n_1201)
);

NOR2xp33_ASAP7_75t_L g1202 ( 
.A(n_978),
.B(n_352),
.Y(n_1202)
);

AOI21xp5_ASAP7_75t_L g1203 ( 
.A1(n_941),
.A2(n_547),
.B(n_549),
.Y(n_1203)
);

BUFx2_ASAP7_75t_SL g1204 ( 
.A(n_1057),
.Y(n_1204)
);

A2O1A1Ixp33_ASAP7_75t_L g1205 ( 
.A1(n_1024),
.A2(n_358),
.B(n_408),
.C(n_411),
.Y(n_1205)
);

AO32x1_ASAP7_75t_L g1206 ( 
.A1(n_972),
.A2(n_601),
.A3(n_588),
.B1(n_575),
.B2(n_574),
.Y(n_1206)
);

AND2x2_ASAP7_75t_L g1207 ( 
.A(n_974),
.B(n_361),
.Y(n_1207)
);

INVx2_ASAP7_75t_L g1208 ( 
.A(n_990),
.Y(n_1208)
);

AOI21xp5_ASAP7_75t_L g1209 ( 
.A1(n_989),
.A2(n_547),
.B(n_549),
.Y(n_1209)
);

NAND2xp5_ASAP7_75t_L g1210 ( 
.A(n_1109),
.B(n_571),
.Y(n_1210)
);

AOI21xp5_ASAP7_75t_L g1211 ( 
.A1(n_993),
.A2(n_547),
.B(n_549),
.Y(n_1211)
);

INVx3_ASAP7_75t_L g1212 ( 
.A(n_997),
.Y(n_1212)
);

NAND2xp5_ASAP7_75t_L g1213 ( 
.A(n_1059),
.B(n_571),
.Y(n_1213)
);

INVx4_ASAP7_75t_L g1214 ( 
.A(n_997),
.Y(n_1214)
);

BUFx6f_ASAP7_75t_L g1215 ( 
.A(n_997),
.Y(n_1215)
);

A2O1A1Ixp33_ASAP7_75t_L g1216 ( 
.A1(n_999),
.A2(n_353),
.B(n_412),
.C(n_575),
.Y(n_1216)
);

NAND3xp33_ASAP7_75t_SL g1217 ( 
.A(n_1035),
.B(n_1025),
.C(n_1078),
.Y(n_1217)
);

NAND2xp5_ASAP7_75t_L g1218 ( 
.A(n_1059),
.B(n_572),
.Y(n_1218)
);

NAND2xp5_ASAP7_75t_L g1219 ( 
.A(n_1001),
.B(n_572),
.Y(n_1219)
);

OAI22xp5_ASAP7_75t_L g1220 ( 
.A1(n_935),
.A2(n_601),
.B1(n_588),
.B2(n_574),
.Y(n_1220)
);

A2O1A1Ixp33_ASAP7_75t_L g1221 ( 
.A1(n_999),
.A2(n_601),
.B(n_574),
.C(n_572),
.Y(n_1221)
);

BUFx2_ASAP7_75t_L g1222 ( 
.A(n_1065),
.Y(n_1222)
);

NAND2xp5_ASAP7_75t_L g1223 ( 
.A(n_966),
.B(n_1039),
.Y(n_1223)
);

INVx2_ASAP7_75t_L g1224 ( 
.A(n_1027),
.Y(n_1224)
);

AOI21xp5_ASAP7_75t_L g1225 ( 
.A1(n_994),
.A2(n_549),
.B(n_547),
.Y(n_1225)
);

INVx1_ASAP7_75t_L g1226 ( 
.A(n_1040),
.Y(n_1226)
);

HB1xp67_ASAP7_75t_L g1227 ( 
.A(n_997),
.Y(n_1227)
);

BUFx2_ASAP7_75t_L g1228 ( 
.A(n_1036),
.Y(n_1228)
);

NAND2xp5_ASAP7_75t_L g1229 ( 
.A(n_966),
.B(n_572),
.Y(n_1229)
);

BUFx2_ASAP7_75t_L g1230 ( 
.A(n_1021),
.Y(n_1230)
);

AND2x2_ASAP7_75t_L g1231 ( 
.A(n_1078),
.B(n_361),
.Y(n_1231)
);

CKINVDCx5p33_ASAP7_75t_R g1232 ( 
.A(n_1095),
.Y(n_1232)
);

INVx2_ASAP7_75t_L g1233 ( 
.A(n_1040),
.Y(n_1233)
);

HB1xp67_ASAP7_75t_L g1234 ( 
.A(n_1009),
.Y(n_1234)
);

OA21x2_ASAP7_75t_L g1235 ( 
.A1(n_1014),
.A2(n_528),
.B(n_601),
.Y(n_1235)
);

AO32x1_ASAP7_75t_L g1236 ( 
.A1(n_1006),
.A2(n_528),
.A3(n_350),
.B1(n_388),
.B2(n_413),
.Y(n_1236)
);

INVx2_ASAP7_75t_L g1237 ( 
.A(n_1074),
.Y(n_1237)
);

AOI21xp5_ASAP7_75t_L g1238 ( 
.A1(n_1034),
.A2(n_549),
.B(n_557),
.Y(n_1238)
);

A2O1A1Ixp33_ASAP7_75t_L g1239 ( 
.A1(n_956),
.A2(n_413),
.B(n_388),
.C(n_361),
.Y(n_1239)
);

NAND2xp5_ASAP7_75t_L g1240 ( 
.A(n_961),
.B(n_557),
.Y(n_1240)
);

AOI22xp33_ASAP7_75t_L g1241 ( 
.A1(n_1069),
.A2(n_413),
.B1(n_388),
.B2(n_557),
.Y(n_1241)
);

AOI21xp5_ASAP7_75t_L g1242 ( 
.A1(n_1007),
.A2(n_549),
.B(n_557),
.Y(n_1242)
);

AOI21xp5_ASAP7_75t_L g1243 ( 
.A1(n_945),
.A2(n_549),
.B(n_557),
.Y(n_1243)
);

BUFx3_ASAP7_75t_L g1244 ( 
.A(n_1009),
.Y(n_1244)
);

BUFx3_ASAP7_75t_L g1245 ( 
.A(n_1009),
.Y(n_1245)
);

NAND2xp5_ASAP7_75t_L g1246 ( 
.A(n_956),
.B(n_557),
.Y(n_1246)
);

INVx3_ASAP7_75t_L g1247 ( 
.A(n_1070),
.Y(n_1247)
);

O2A1O1Ixp33_ASAP7_75t_L g1248 ( 
.A1(n_935),
.A2(n_18),
.B(n_19),
.C(n_20),
.Y(n_1248)
);

INVx3_ASAP7_75t_L g1249 ( 
.A(n_1070),
.Y(n_1249)
);

INVx1_ASAP7_75t_SL g1250 ( 
.A(n_1075),
.Y(n_1250)
);

INVx1_ASAP7_75t_SL g1251 ( 
.A(n_1067),
.Y(n_1251)
);

AOI21xp5_ASAP7_75t_L g1252 ( 
.A1(n_948),
.A2(n_1046),
.B(n_1044),
.Y(n_1252)
);

INVx8_ASAP7_75t_L g1253 ( 
.A(n_1030),
.Y(n_1253)
);

OR2x6_ASAP7_75t_L g1254 ( 
.A(n_1077),
.B(n_95),
.Y(n_1254)
);

NOR2xp33_ASAP7_75t_L g1255 ( 
.A(n_1095),
.B(n_24),
.Y(n_1255)
);

AOI21xp5_ASAP7_75t_L g1256 ( 
.A1(n_1049),
.A2(n_209),
.B(n_193),
.Y(n_1256)
);

HB1xp67_ASAP7_75t_L g1257 ( 
.A(n_1074),
.Y(n_1257)
);

NOR2xp33_ASAP7_75t_L g1258 ( 
.A(n_1003),
.B(n_30),
.Y(n_1258)
);

OAI21xp5_ASAP7_75t_L g1259 ( 
.A1(n_1038),
.A2(n_169),
.B(n_167),
.Y(n_1259)
);

AOI21xp5_ASAP7_75t_L g1260 ( 
.A1(n_1023),
.A2(n_957),
.B(n_1010),
.Y(n_1260)
);

INVx1_ASAP7_75t_L g1261 ( 
.A(n_1088),
.Y(n_1261)
);

NAND2xp5_ASAP7_75t_L g1262 ( 
.A(n_1030),
.B(n_31),
.Y(n_1262)
);

BUFx3_ASAP7_75t_L g1263 ( 
.A(n_1012),
.Y(n_1263)
);

OAI21xp33_ASAP7_75t_L g1264 ( 
.A1(n_1112),
.A2(n_32),
.B(n_34),
.Y(n_1264)
);

NAND2xp5_ASAP7_75t_L g1265 ( 
.A(n_1088),
.B(n_35),
.Y(n_1265)
);

NAND2x1p5_ASAP7_75t_L g1266 ( 
.A(n_1077),
.B(n_166),
.Y(n_1266)
);

NOR2xp33_ASAP7_75t_R g1267 ( 
.A(n_1060),
.B(n_132),
.Y(n_1267)
);

AOI21xp5_ASAP7_75t_L g1268 ( 
.A1(n_1010),
.A2(n_163),
.B(n_161),
.Y(n_1268)
);

INVxp67_ASAP7_75t_L g1269 ( 
.A(n_1086),
.Y(n_1269)
);

INVx1_ASAP7_75t_L g1270 ( 
.A(n_1103),
.Y(n_1270)
);

OAI21xp5_ASAP7_75t_L g1271 ( 
.A1(n_1047),
.A2(n_158),
.B(n_154),
.Y(n_1271)
);

OAI21xp5_ASAP7_75t_L g1272 ( 
.A1(n_1260),
.A2(n_1116),
.B(n_1056),
.Y(n_1272)
);

AO31x2_ASAP7_75t_L g1273 ( 
.A1(n_1125),
.A2(n_955),
.A3(n_1033),
.B(n_987),
.Y(n_1273)
);

BUFx2_ASAP7_75t_L g1274 ( 
.A(n_1135),
.Y(n_1274)
);

O2A1O1Ixp33_ASAP7_75t_L g1275 ( 
.A1(n_1255),
.A2(n_1045),
.B(n_1058),
.C(n_1073),
.Y(n_1275)
);

OAI21x1_ASAP7_75t_L g1276 ( 
.A1(n_1187),
.A2(n_981),
.B(n_1029),
.Y(n_1276)
);

NOR2xp33_ASAP7_75t_L g1277 ( 
.A(n_1178),
.B(n_1251),
.Y(n_1277)
);

NAND2xp5_ASAP7_75t_L g1278 ( 
.A(n_1147),
.B(n_1004),
.Y(n_1278)
);

BUFx6f_ASAP7_75t_L g1279 ( 
.A(n_1191),
.Y(n_1279)
);

NAND2x1_ASAP7_75t_L g1280 ( 
.A(n_1214),
.B(n_1115),
.Y(n_1280)
);

NAND2x1p5_ASAP7_75t_L g1281 ( 
.A(n_1160),
.B(n_1115),
.Y(n_1281)
);

OAI22xp5_ASAP7_75t_L g1282 ( 
.A1(n_1131),
.A2(n_1060),
.B1(n_1098),
.B2(n_959),
.Y(n_1282)
);

AOI21xp5_ASAP7_75t_L g1283 ( 
.A1(n_1252),
.A2(n_1098),
.B(n_964),
.Y(n_1283)
);

AOI21xp5_ASAP7_75t_L g1284 ( 
.A1(n_1120),
.A2(n_1055),
.B(n_1113),
.Y(n_1284)
);

INVxp67_ASAP7_75t_L g1285 ( 
.A(n_1136),
.Y(n_1285)
);

INVx1_ASAP7_75t_L g1286 ( 
.A(n_1257),
.Y(n_1286)
);

OAI21x1_ASAP7_75t_L g1287 ( 
.A1(n_1194),
.A2(n_1011),
.B(n_1013),
.Y(n_1287)
);

OAI21x1_ASAP7_75t_L g1288 ( 
.A1(n_1209),
.A2(n_1094),
.B(n_1091),
.Y(n_1288)
);

INVx1_ASAP7_75t_L g1289 ( 
.A(n_1257),
.Y(n_1289)
);

INVx5_ASAP7_75t_L g1290 ( 
.A(n_1146),
.Y(n_1290)
);

OAI21xp5_ASAP7_75t_L g1291 ( 
.A1(n_1119),
.A2(n_1114),
.B(n_970),
.Y(n_1291)
);

OAI22xp33_ASAP7_75t_L g1292 ( 
.A1(n_1232),
.A2(n_1255),
.B1(n_1250),
.B2(n_1223),
.Y(n_1292)
);

A2O1A1Ixp33_ASAP7_75t_L g1293 ( 
.A1(n_1125),
.A2(n_1217),
.B(n_1259),
.C(n_1158),
.Y(n_1293)
);

OAI21x1_ASAP7_75t_L g1294 ( 
.A1(n_1211),
.A2(n_1048),
.B(n_1000),
.Y(n_1294)
);

OAI21x1_ASAP7_75t_L g1295 ( 
.A1(n_1225),
.A2(n_1106),
.B(n_1041),
.Y(n_1295)
);

OAI22xp5_ASAP7_75t_L g1296 ( 
.A1(n_1269),
.A2(n_952),
.B1(n_1015),
.B2(n_1082),
.Y(n_1296)
);

INVxp67_ASAP7_75t_L g1297 ( 
.A(n_1136),
.Y(n_1297)
);

OAI21x1_ASAP7_75t_L g1298 ( 
.A1(n_1163),
.A2(n_1020),
.B(n_1037),
.Y(n_1298)
);

NAND2xp5_ASAP7_75t_L g1299 ( 
.A(n_1174),
.B(n_1043),
.Y(n_1299)
);

AOI221x1_ASAP7_75t_L g1300 ( 
.A1(n_1264),
.A2(n_1079),
.B1(n_1076),
.B2(n_1080),
.C(n_1083),
.Y(n_1300)
);

NOR4xp25_ASAP7_75t_L g1301 ( 
.A(n_1248),
.B(n_1108),
.C(n_1054),
.D(n_1072),
.Y(n_1301)
);

BUFx6f_ASAP7_75t_L g1302 ( 
.A(n_1188),
.Y(n_1302)
);

OAI21x1_ASAP7_75t_L g1303 ( 
.A1(n_1238),
.A2(n_1042),
.B(n_1068),
.Y(n_1303)
);

INVx1_ASAP7_75t_L g1304 ( 
.A(n_1145),
.Y(n_1304)
);

INVx5_ASAP7_75t_SL g1305 ( 
.A(n_1122),
.Y(n_1305)
);

OAI22xp5_ASAP7_75t_L g1306 ( 
.A1(n_1269),
.A2(n_952),
.B1(n_1015),
.B2(n_1085),
.Y(n_1306)
);

AO31x2_ASAP7_75t_L g1307 ( 
.A1(n_1192),
.A2(n_1092),
.A3(n_1093),
.B(n_1096),
.Y(n_1307)
);

AO21x1_ASAP7_75t_L g1308 ( 
.A1(n_1271),
.A2(n_1053),
.B(n_1022),
.Y(n_1308)
);

BUFx2_ASAP7_75t_L g1309 ( 
.A(n_1162),
.Y(n_1309)
);

NAND2xp5_ASAP7_75t_L g1310 ( 
.A(n_1174),
.B(n_1123),
.Y(n_1310)
);

AOI21xp5_ASAP7_75t_L g1311 ( 
.A1(n_1120),
.A2(n_1018),
.B(n_1061),
.Y(n_1311)
);

OR2x6_ASAP7_75t_L g1312 ( 
.A(n_1254),
.B(n_1107),
.Y(n_1312)
);

OAI22x1_ASAP7_75t_L g1313 ( 
.A1(n_1207),
.A2(n_1101),
.B1(n_1100),
.B2(n_1099),
.Y(n_1313)
);

BUFx2_ASAP7_75t_L g1314 ( 
.A(n_1222),
.Y(n_1314)
);

OAI21xp5_ASAP7_75t_L g1315 ( 
.A1(n_1119),
.A2(n_1066),
.B(n_1064),
.Y(n_1315)
);

AND2x2_ASAP7_75t_L g1316 ( 
.A(n_1148),
.B(n_1090),
.Y(n_1316)
);

OAI21xp5_ASAP7_75t_L g1317 ( 
.A1(n_1149),
.A2(n_1062),
.B(n_1089),
.Y(n_1317)
);

AOI21xp5_ASAP7_75t_L g1318 ( 
.A1(n_1128),
.A2(n_1087),
.B(n_151),
.Y(n_1318)
);

CKINVDCx5p33_ASAP7_75t_R g1319 ( 
.A(n_1127),
.Y(n_1319)
);

AOI22xp5_ASAP7_75t_L g1320 ( 
.A1(n_1118),
.A2(n_37),
.B1(n_38),
.B2(n_39),
.Y(n_1320)
);

OAI21xp5_ASAP7_75t_L g1321 ( 
.A1(n_1137),
.A2(n_150),
.B(n_148),
.Y(n_1321)
);

OAI21x1_ASAP7_75t_L g1322 ( 
.A1(n_1180),
.A2(n_144),
.B(n_143),
.Y(n_1322)
);

HB1xp67_ASAP7_75t_L g1323 ( 
.A(n_1134),
.Y(n_1323)
);

INVx1_ASAP7_75t_SL g1324 ( 
.A(n_1154),
.Y(n_1324)
);

INVx2_ASAP7_75t_SL g1325 ( 
.A(n_1177),
.Y(n_1325)
);

AOI21xp5_ASAP7_75t_L g1326 ( 
.A1(n_1141),
.A2(n_142),
.B(n_137),
.Y(n_1326)
);

NAND2xp5_ASAP7_75t_L g1327 ( 
.A(n_1130),
.B(n_37),
.Y(n_1327)
);

AOI21xp5_ASAP7_75t_L g1328 ( 
.A1(n_1142),
.A2(n_131),
.B(n_128),
.Y(n_1328)
);

NAND2xp5_ASAP7_75t_L g1329 ( 
.A(n_1231),
.B(n_39),
.Y(n_1329)
);

NAND2xp5_ASAP7_75t_L g1330 ( 
.A(n_1258),
.B(n_40),
.Y(n_1330)
);

NAND2xp5_ASAP7_75t_L g1331 ( 
.A(n_1258),
.B(n_1129),
.Y(n_1331)
);

NAND2xp5_ASAP7_75t_L g1332 ( 
.A(n_1167),
.B(n_47),
.Y(n_1332)
);

AOI22xp5_ASAP7_75t_L g1333 ( 
.A1(n_1202),
.A2(n_47),
.B1(n_48),
.B2(n_49),
.Y(n_1333)
);

AO21x1_ASAP7_75t_L g1334 ( 
.A1(n_1246),
.A2(n_50),
.B(n_51),
.Y(n_1334)
);

NAND3xp33_ASAP7_75t_L g1335 ( 
.A(n_1239),
.B(n_1202),
.C(n_1195),
.Y(n_1335)
);

AOI21xp5_ASAP7_75t_L g1336 ( 
.A1(n_1138),
.A2(n_121),
.B(n_119),
.Y(n_1336)
);

NAND2xp5_ASAP7_75t_L g1337 ( 
.A(n_1151),
.B(n_51),
.Y(n_1337)
);

O2A1O1Ixp33_ASAP7_75t_L g1338 ( 
.A1(n_1239),
.A2(n_57),
.B(n_58),
.C(n_60),
.Y(n_1338)
);

AOI21xp5_ASAP7_75t_L g1339 ( 
.A1(n_1138),
.A2(n_118),
.B(n_115),
.Y(n_1339)
);

AOI221x1_ASAP7_75t_L g1340 ( 
.A1(n_1216),
.A2(n_58),
.B1(n_61),
.B2(n_64),
.C(n_65),
.Y(n_1340)
);

BUFx6f_ASAP7_75t_L g1341 ( 
.A(n_1188),
.Y(n_1341)
);

INVx1_ASAP7_75t_L g1342 ( 
.A(n_1157),
.Y(n_1342)
);

NAND2xp5_ASAP7_75t_L g1343 ( 
.A(n_1143),
.B(n_61),
.Y(n_1343)
);

O2A1O1Ixp33_ASAP7_75t_SL g1344 ( 
.A1(n_1216),
.A2(n_114),
.B(n_110),
.C(n_105),
.Y(n_1344)
);

NAND3xp33_ASAP7_75t_L g1345 ( 
.A(n_1193),
.B(n_1205),
.C(n_1195),
.Y(n_1345)
);

NAND2xp5_ASAP7_75t_L g1346 ( 
.A(n_1253),
.B(n_66),
.Y(n_1346)
);

INVx4_ASAP7_75t_L g1347 ( 
.A(n_1160),
.Y(n_1347)
);

AOI22xp5_ASAP7_75t_L g1348 ( 
.A1(n_1253),
.A2(n_66),
.B1(n_67),
.B2(n_68),
.Y(n_1348)
);

NOR2xp33_ASAP7_75t_SL g1349 ( 
.A(n_1186),
.B(n_68),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_1161),
.Y(n_1350)
);

OAI21x1_ASAP7_75t_L g1351 ( 
.A1(n_1132),
.A2(n_100),
.B(n_75),
.Y(n_1351)
);

NAND2xp33_ASAP7_75t_L g1352 ( 
.A(n_1200),
.B(n_1160),
.Y(n_1352)
);

AOI21xp5_ASAP7_75t_L g1353 ( 
.A1(n_1133),
.A2(n_70),
.B(n_76),
.Y(n_1353)
);

NAND2xp5_ASAP7_75t_L g1354 ( 
.A(n_1253),
.B(n_70),
.Y(n_1354)
);

AOI21xp5_ASAP7_75t_L g1355 ( 
.A1(n_1183),
.A2(n_76),
.B(n_77),
.Y(n_1355)
);

NOR2xp33_ASAP7_75t_L g1356 ( 
.A(n_1153),
.B(n_80),
.Y(n_1356)
);

AOI21xp5_ASAP7_75t_L g1357 ( 
.A1(n_1219),
.A2(n_81),
.B(n_85),
.Y(n_1357)
);

NOR2xp67_ASAP7_75t_L g1358 ( 
.A(n_1160),
.B(n_85),
.Y(n_1358)
);

AO31x2_ASAP7_75t_L g1359 ( 
.A1(n_1221),
.A2(n_1164),
.A3(n_1220),
.B(n_1205),
.Y(n_1359)
);

INVx2_ASAP7_75t_L g1360 ( 
.A(n_1170),
.Y(n_1360)
);

A2O1A1Ixp33_ASAP7_75t_L g1361 ( 
.A1(n_1156),
.A2(n_1164),
.B(n_1193),
.C(n_1168),
.Y(n_1361)
);

NAND3xp33_ASAP7_75t_L g1362 ( 
.A(n_1199),
.B(n_1198),
.C(n_1168),
.Y(n_1362)
);

AOI21xp5_ASAP7_75t_L g1363 ( 
.A1(n_1240),
.A2(n_1152),
.B(n_1185),
.Y(n_1363)
);

INVx3_ASAP7_75t_L g1364 ( 
.A(n_1214),
.Y(n_1364)
);

INVx1_ASAP7_75t_L g1365 ( 
.A(n_1165),
.Y(n_1365)
);

AOI21xp5_ASAP7_75t_L g1366 ( 
.A1(n_1210),
.A2(n_1126),
.B(n_1140),
.Y(n_1366)
);

AND2x2_ASAP7_75t_L g1367 ( 
.A(n_1173),
.B(n_1228),
.Y(n_1367)
);

AOI21xp5_ASAP7_75t_L g1368 ( 
.A1(n_1126),
.A2(n_1140),
.B(n_1203),
.Y(n_1368)
);

BUFx3_ASAP7_75t_L g1369 ( 
.A(n_1150),
.Y(n_1369)
);

BUFx10_ASAP7_75t_L g1370 ( 
.A(n_1254),
.Y(n_1370)
);

OAI21x1_ASAP7_75t_L g1371 ( 
.A1(n_1243),
.A2(n_1242),
.B(n_1235),
.Y(n_1371)
);

BUFx3_ASAP7_75t_L g1372 ( 
.A(n_1173),
.Y(n_1372)
);

O2A1O1Ixp33_ASAP7_75t_L g1373 ( 
.A1(n_1171),
.A2(n_1201),
.B(n_1184),
.C(n_1190),
.Y(n_1373)
);

CKINVDCx6p67_ASAP7_75t_R g1374 ( 
.A(n_1254),
.Y(n_1374)
);

AO31x2_ASAP7_75t_L g1375 ( 
.A1(n_1221),
.A2(n_1265),
.A3(n_1206),
.B(n_1197),
.Y(n_1375)
);

AO31x2_ASAP7_75t_L g1376 ( 
.A1(n_1206),
.A2(n_1262),
.A3(n_1256),
.B(n_1261),
.Y(n_1376)
);

AO21x2_ASAP7_75t_L g1377 ( 
.A1(n_1213),
.A2(n_1218),
.B(n_1270),
.Y(n_1377)
);

OR2x2_ASAP7_75t_L g1378 ( 
.A(n_1229),
.B(n_1175),
.Y(n_1378)
);

CKINVDCx16_ASAP7_75t_R g1379 ( 
.A(n_1181),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_1182),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_1208),
.Y(n_1381)
);

AND2x4_ASAP7_75t_L g1382 ( 
.A(n_1263),
.B(n_1247),
.Y(n_1382)
);

NOR2xp67_ASAP7_75t_L g1383 ( 
.A(n_1247),
.B(n_1249),
.Y(n_1383)
);

AOI21xp5_ASAP7_75t_SL g1384 ( 
.A1(n_1215),
.A2(n_1266),
.B(n_1146),
.Y(n_1384)
);

OA21x2_ASAP7_75t_L g1385 ( 
.A1(n_1166),
.A2(n_1226),
.B(n_1189),
.Y(n_1385)
);

AOI22xp33_ASAP7_75t_L g1386 ( 
.A1(n_1198),
.A2(n_1200),
.B1(n_1230),
.B2(n_1241),
.Y(n_1386)
);

AOI21xp5_ASAP7_75t_L g1387 ( 
.A1(n_1235),
.A2(n_1249),
.B(n_1206),
.Y(n_1387)
);

INVx5_ASAP7_75t_L g1388 ( 
.A(n_1146),
.Y(n_1388)
);

AOI21xp5_ASAP7_75t_L g1389 ( 
.A1(n_1235),
.A2(n_1268),
.B(n_1215),
.Y(n_1389)
);

INVx4_ASAP7_75t_L g1390 ( 
.A(n_1146),
.Y(n_1390)
);

CKINVDCx5p33_ASAP7_75t_R g1391 ( 
.A(n_1267),
.Y(n_1391)
);

NAND2xp5_ASAP7_75t_SL g1392 ( 
.A(n_1169),
.B(n_1215),
.Y(n_1392)
);

CKINVDCx5p33_ASAP7_75t_R g1393 ( 
.A(n_1267),
.Y(n_1393)
);

OAI21x1_ASAP7_75t_L g1394 ( 
.A1(n_1176),
.A2(n_1237),
.B(n_1224),
.Y(n_1394)
);

NAND2xp5_ASAP7_75t_L g1395 ( 
.A(n_1233),
.B(n_1139),
.Y(n_1395)
);

INVx2_ASAP7_75t_L g1396 ( 
.A(n_1144),
.Y(n_1396)
);

O2A1O1Ixp33_ASAP7_75t_L g1397 ( 
.A1(n_1155),
.A2(n_1172),
.B(n_1266),
.C(n_1234),
.Y(n_1397)
);

AO21x2_ASAP7_75t_L g1398 ( 
.A1(n_1227),
.A2(n_1234),
.B(n_1236),
.Y(n_1398)
);

HB1xp67_ASAP7_75t_L g1399 ( 
.A(n_1227),
.Y(n_1399)
);

AO31x2_ASAP7_75t_L g1400 ( 
.A1(n_1236),
.A2(n_1196),
.A3(n_1241),
.B(n_1212),
.Y(n_1400)
);

AOI21xp5_ASAP7_75t_L g1401 ( 
.A1(n_1215),
.A2(n_1196),
.B(n_1124),
.Y(n_1401)
);

NOR2xp33_ASAP7_75t_L g1402 ( 
.A(n_1244),
.B(n_1245),
.Y(n_1402)
);

BUFx2_ASAP7_75t_R g1403 ( 
.A(n_1204),
.Y(n_1403)
);

NAND2x1p5_ASAP7_75t_L g1404 ( 
.A(n_1236),
.B(n_1160),
.Y(n_1404)
);

BUFx6f_ASAP7_75t_SL g1405 ( 
.A(n_1162),
.Y(n_1405)
);

OAI22xp5_ASAP7_75t_L g1406 ( 
.A1(n_1178),
.A2(n_782),
.B1(n_764),
.B2(n_1147),
.Y(n_1406)
);

AOI21xp5_ASAP7_75t_L g1407 ( 
.A1(n_1252),
.A2(n_883),
.B(n_982),
.Y(n_1407)
);

CKINVDCx20_ASAP7_75t_R g1408 ( 
.A(n_1122),
.Y(n_1408)
);

OAI22xp5_ASAP7_75t_L g1409 ( 
.A1(n_1178),
.A2(n_782),
.B1(n_764),
.B2(n_1147),
.Y(n_1409)
);

AOI22xp5_ASAP7_75t_L g1410 ( 
.A1(n_1178),
.A2(n_782),
.B1(n_1031),
.B2(n_1255),
.Y(n_1410)
);

INVx1_ASAP7_75t_L g1411 ( 
.A(n_1257),
.Y(n_1411)
);

AO31x2_ASAP7_75t_L g1412 ( 
.A1(n_1260),
.A2(n_955),
.A3(n_976),
.B(n_1159),
.Y(n_1412)
);

OA21x2_ASAP7_75t_L g1413 ( 
.A1(n_1260),
.A2(n_1192),
.B(n_1259),
.Y(n_1413)
);

INVx1_ASAP7_75t_L g1414 ( 
.A(n_1257),
.Y(n_1414)
);

NOR2xp67_ASAP7_75t_SL g1415 ( 
.A(n_1191),
.B(n_936),
.Y(n_1415)
);

O2A1O1Ixp33_ASAP7_75t_L g1416 ( 
.A1(n_1255),
.A2(n_782),
.B(n_1031),
.C(n_1178),
.Y(n_1416)
);

AO32x2_ASAP7_75t_L g1417 ( 
.A1(n_1133),
.A2(n_972),
.A3(n_1073),
.B1(n_1006),
.B2(n_1121),
.Y(n_1417)
);

AOI21xp5_ASAP7_75t_L g1418 ( 
.A1(n_1252),
.A2(n_883),
.B(n_982),
.Y(n_1418)
);

AOI21xp5_ASAP7_75t_L g1419 ( 
.A1(n_1252),
.A2(n_883),
.B(n_982),
.Y(n_1419)
);

OAI22x1_ASAP7_75t_L g1420 ( 
.A1(n_1178),
.A2(n_1255),
.B1(n_782),
.B2(n_876),
.Y(n_1420)
);

AOI22xp5_ASAP7_75t_L g1421 ( 
.A1(n_1178),
.A2(n_782),
.B1(n_1031),
.B2(n_1255),
.Y(n_1421)
);

O2A1O1Ixp33_ASAP7_75t_L g1422 ( 
.A1(n_1255),
.A2(n_782),
.B(n_1031),
.C(n_1178),
.Y(n_1422)
);

AOI21xp5_ASAP7_75t_L g1423 ( 
.A1(n_1252),
.A2(n_883),
.B(n_982),
.Y(n_1423)
);

NAND2xp5_ASAP7_75t_L g1424 ( 
.A(n_1147),
.B(n_782),
.Y(n_1424)
);

AND2x2_ASAP7_75t_L g1425 ( 
.A(n_1178),
.B(n_950),
.Y(n_1425)
);

BUFx6f_ASAP7_75t_L g1426 ( 
.A(n_1191),
.Y(n_1426)
);

AO31x2_ASAP7_75t_L g1427 ( 
.A1(n_1260),
.A2(n_955),
.A3(n_976),
.B(n_1159),
.Y(n_1427)
);

INVx1_ASAP7_75t_L g1428 ( 
.A(n_1257),
.Y(n_1428)
);

OAI21x1_ASAP7_75t_L g1429 ( 
.A1(n_1179),
.A2(n_1111),
.B(n_1159),
.Y(n_1429)
);

AND2x2_ASAP7_75t_L g1430 ( 
.A(n_1178),
.B(n_950),
.Y(n_1430)
);

NOR2xp67_ASAP7_75t_SL g1431 ( 
.A(n_1191),
.B(n_936),
.Y(n_1431)
);

OR2x2_ASAP7_75t_L g1432 ( 
.A(n_1178),
.B(n_915),
.Y(n_1432)
);

AOI21xp5_ASAP7_75t_L g1433 ( 
.A1(n_1252),
.A2(n_883),
.B(n_982),
.Y(n_1433)
);

BUFx3_ASAP7_75t_L g1434 ( 
.A(n_1135),
.Y(n_1434)
);

OAI21x1_ASAP7_75t_SL g1435 ( 
.A1(n_1158),
.A2(n_1262),
.B(n_1259),
.Y(n_1435)
);

NAND2xp5_ASAP7_75t_L g1436 ( 
.A(n_1147),
.B(n_782),
.Y(n_1436)
);

NAND2xp5_ASAP7_75t_L g1437 ( 
.A(n_1147),
.B(n_782),
.Y(n_1437)
);

INVx2_ASAP7_75t_L g1438 ( 
.A(n_1170),
.Y(n_1438)
);

INVx4_ASAP7_75t_L g1439 ( 
.A(n_1302),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_1304),
.Y(n_1440)
);

INVx2_ASAP7_75t_SL g1441 ( 
.A(n_1279),
.Y(n_1441)
);

INVx2_ASAP7_75t_L g1442 ( 
.A(n_1385),
.Y(n_1442)
);

AOI22xp33_ASAP7_75t_L g1443 ( 
.A1(n_1410),
.A2(n_1421),
.B1(n_1420),
.B2(n_1362),
.Y(n_1443)
);

INVx2_ASAP7_75t_L g1444 ( 
.A(n_1385),
.Y(n_1444)
);

INVx2_ASAP7_75t_L g1445 ( 
.A(n_1360),
.Y(n_1445)
);

AOI22xp33_ASAP7_75t_L g1446 ( 
.A1(n_1410),
.A2(n_1421),
.B1(n_1362),
.B2(n_1330),
.Y(n_1446)
);

INVx2_ASAP7_75t_L g1447 ( 
.A(n_1438),
.Y(n_1447)
);

INVx1_ASAP7_75t_L g1448 ( 
.A(n_1342),
.Y(n_1448)
);

CKINVDCx20_ASAP7_75t_R g1449 ( 
.A(n_1408),
.Y(n_1449)
);

INVx6_ASAP7_75t_L g1450 ( 
.A(n_1279),
.Y(n_1450)
);

BUFx2_ASAP7_75t_L g1451 ( 
.A(n_1314),
.Y(n_1451)
);

BUFx4f_ASAP7_75t_SL g1452 ( 
.A(n_1279),
.Y(n_1452)
);

OAI22xp33_ASAP7_75t_L g1453 ( 
.A1(n_1349),
.A2(n_1333),
.B1(n_1320),
.B2(n_1348),
.Y(n_1453)
);

OAI22xp5_ASAP7_75t_L g1454 ( 
.A1(n_1416),
.A2(n_1422),
.B1(n_1277),
.B2(n_1292),
.Y(n_1454)
);

BUFx3_ASAP7_75t_L g1455 ( 
.A(n_1426),
.Y(n_1455)
);

AOI22xp33_ASAP7_75t_SL g1456 ( 
.A1(n_1349),
.A2(n_1335),
.B1(n_1356),
.B2(n_1329),
.Y(n_1456)
);

INVx6_ASAP7_75t_L g1457 ( 
.A(n_1426),
.Y(n_1457)
);

AOI22xp33_ASAP7_75t_L g1458 ( 
.A1(n_1333),
.A2(n_1335),
.B1(n_1348),
.B2(n_1320),
.Y(n_1458)
);

AOI22xp5_ASAP7_75t_L g1459 ( 
.A1(n_1425),
.A2(n_1430),
.B1(n_1436),
.B2(n_1424),
.Y(n_1459)
);

BUFx2_ASAP7_75t_L g1460 ( 
.A(n_1309),
.Y(n_1460)
);

INVx6_ASAP7_75t_L g1461 ( 
.A(n_1426),
.Y(n_1461)
);

INVx1_ASAP7_75t_L g1462 ( 
.A(n_1350),
.Y(n_1462)
);

INVx2_ASAP7_75t_L g1463 ( 
.A(n_1380),
.Y(n_1463)
);

CKINVDCx11_ASAP7_75t_R g1464 ( 
.A(n_1379),
.Y(n_1464)
);

AOI22xp33_ASAP7_75t_L g1465 ( 
.A1(n_1437),
.A2(n_1409),
.B1(n_1406),
.B2(n_1331),
.Y(n_1465)
);

BUFx10_ASAP7_75t_L g1466 ( 
.A(n_1405),
.Y(n_1466)
);

BUFx4f_ASAP7_75t_SL g1467 ( 
.A(n_1434),
.Y(n_1467)
);

NAND2x1p5_ASAP7_75t_L g1468 ( 
.A(n_1290),
.B(n_1388),
.Y(n_1468)
);

INVxp67_ASAP7_75t_L g1469 ( 
.A(n_1323),
.Y(n_1469)
);

INVx2_ASAP7_75t_L g1470 ( 
.A(n_1381),
.Y(n_1470)
);

AOI22xp33_ASAP7_75t_L g1471 ( 
.A1(n_1345),
.A2(n_1334),
.B1(n_1353),
.B2(n_1432),
.Y(n_1471)
);

OAI22xp33_ASAP7_75t_L g1472 ( 
.A1(n_1374),
.A2(n_1324),
.B1(n_1393),
.B2(n_1391),
.Y(n_1472)
);

CKINVDCx11_ASAP7_75t_R g1473 ( 
.A(n_1274),
.Y(n_1473)
);

AOI22xp33_ASAP7_75t_L g1474 ( 
.A1(n_1345),
.A2(n_1435),
.B1(n_1337),
.B2(n_1386),
.Y(n_1474)
);

INVx2_ASAP7_75t_SL g1475 ( 
.A(n_1325),
.Y(n_1475)
);

NAND2xp5_ASAP7_75t_L g1476 ( 
.A(n_1310),
.B(n_1324),
.Y(n_1476)
);

CKINVDCx20_ASAP7_75t_R g1477 ( 
.A(n_1319),
.Y(n_1477)
);

AND2x2_ASAP7_75t_L g1478 ( 
.A(n_1367),
.B(n_1399),
.Y(n_1478)
);

BUFx12f_ASAP7_75t_L g1479 ( 
.A(n_1370),
.Y(n_1479)
);

INVx8_ASAP7_75t_L g1480 ( 
.A(n_1290),
.Y(n_1480)
);

HB1xp67_ASAP7_75t_L g1481 ( 
.A(n_1285),
.Y(n_1481)
);

AOI22xp33_ASAP7_75t_L g1482 ( 
.A1(n_1355),
.A2(n_1321),
.B1(n_1357),
.B2(n_1354),
.Y(n_1482)
);

AOI22xp33_ASAP7_75t_SL g1483 ( 
.A1(n_1321),
.A2(n_1332),
.B1(n_1346),
.B2(n_1327),
.Y(n_1483)
);

INVx2_ASAP7_75t_L g1484 ( 
.A(n_1394),
.Y(n_1484)
);

AND2x2_ASAP7_75t_L g1485 ( 
.A(n_1286),
.B(n_1289),
.Y(n_1485)
);

OAI21xp5_ASAP7_75t_SL g1486 ( 
.A1(n_1338),
.A2(n_1340),
.B(n_1361),
.Y(n_1486)
);

INVx2_ASAP7_75t_SL g1487 ( 
.A(n_1369),
.Y(n_1487)
);

OAI22xp5_ASAP7_75t_L g1488 ( 
.A1(n_1293),
.A2(n_1372),
.B1(n_1299),
.B2(n_1297),
.Y(n_1488)
);

AOI22xp33_ASAP7_75t_L g1489 ( 
.A1(n_1316),
.A2(n_1278),
.B1(n_1378),
.B2(n_1343),
.Y(n_1489)
);

INVx6_ASAP7_75t_L g1490 ( 
.A(n_1302),
.Y(n_1490)
);

OAI22xp33_ASAP7_75t_SL g1491 ( 
.A1(n_1392),
.A2(n_1312),
.B1(n_1428),
.B2(n_1411),
.Y(n_1491)
);

AOI22xp33_ASAP7_75t_L g1492 ( 
.A1(n_1414),
.A2(n_1365),
.B1(n_1413),
.B2(n_1370),
.Y(n_1492)
);

INVx1_ASAP7_75t_SL g1493 ( 
.A(n_1403),
.Y(n_1493)
);

CKINVDCx11_ASAP7_75t_R g1494 ( 
.A(n_1302),
.Y(n_1494)
);

AOI22xp33_ASAP7_75t_L g1495 ( 
.A1(n_1413),
.A2(n_1272),
.B1(n_1313),
.B2(n_1326),
.Y(n_1495)
);

AOI22xp33_ASAP7_75t_L g1496 ( 
.A1(n_1308),
.A2(n_1396),
.B1(n_1282),
.B2(n_1312),
.Y(n_1496)
);

CKINVDCx16_ASAP7_75t_R g1497 ( 
.A(n_1405),
.Y(n_1497)
);

AOI22xp5_ASAP7_75t_L g1498 ( 
.A1(n_1415),
.A2(n_1431),
.B1(n_1312),
.B2(n_1382),
.Y(n_1498)
);

INVx3_ASAP7_75t_L g1499 ( 
.A(n_1347),
.Y(n_1499)
);

INVxp67_ASAP7_75t_SL g1500 ( 
.A(n_1352),
.Y(n_1500)
);

AND2x2_ASAP7_75t_L g1501 ( 
.A(n_1402),
.B(n_1382),
.Y(n_1501)
);

INVx3_ASAP7_75t_L g1502 ( 
.A(n_1341),
.Y(n_1502)
);

AOI22xp5_ASAP7_75t_L g1503 ( 
.A1(n_1358),
.A2(n_1306),
.B1(n_1296),
.B2(n_1383),
.Y(n_1503)
);

AOI22xp33_ASAP7_75t_L g1504 ( 
.A1(n_1377),
.A2(n_1328),
.B1(n_1358),
.B2(n_1291),
.Y(n_1504)
);

AOI22xp33_ASAP7_75t_SL g1505 ( 
.A1(n_1336),
.A2(n_1339),
.B1(n_1305),
.B2(n_1341),
.Y(n_1505)
);

AOI22xp33_ASAP7_75t_L g1506 ( 
.A1(n_1377),
.A2(n_1291),
.B1(n_1284),
.B2(n_1395),
.Y(n_1506)
);

AOI22xp33_ASAP7_75t_L g1507 ( 
.A1(n_1363),
.A2(n_1366),
.B1(n_1317),
.B2(n_1311),
.Y(n_1507)
);

OAI22xp33_ASAP7_75t_L g1508 ( 
.A1(n_1341),
.A2(n_1300),
.B1(n_1383),
.B2(n_1364),
.Y(n_1508)
);

BUFx2_ASAP7_75t_SL g1509 ( 
.A(n_1388),
.Y(n_1509)
);

INVx6_ASAP7_75t_L g1510 ( 
.A(n_1390),
.Y(n_1510)
);

CKINVDCx11_ASAP7_75t_R g1511 ( 
.A(n_1305),
.Y(n_1511)
);

AOI22xp33_ASAP7_75t_SL g1512 ( 
.A1(n_1351),
.A2(n_1283),
.B1(n_1404),
.B2(n_1322),
.Y(n_1512)
);

OAI21xp33_ASAP7_75t_L g1513 ( 
.A1(n_1275),
.A2(n_1373),
.B(n_1301),
.Y(n_1513)
);

AOI22xp33_ASAP7_75t_SL g1514 ( 
.A1(n_1417),
.A2(n_1318),
.B1(n_1364),
.B2(n_1281),
.Y(n_1514)
);

AOI22xp33_ASAP7_75t_SL g1515 ( 
.A1(n_1417),
.A2(n_1317),
.B1(n_1315),
.B2(n_1344),
.Y(n_1515)
);

BUFx12f_ASAP7_75t_L g1516 ( 
.A(n_1390),
.Y(n_1516)
);

CKINVDCx5p33_ASAP7_75t_R g1517 ( 
.A(n_1384),
.Y(n_1517)
);

AOI22xp33_ASAP7_75t_L g1518 ( 
.A1(n_1417),
.A2(n_1315),
.B1(n_1398),
.B2(n_1368),
.Y(n_1518)
);

INVx5_ASAP7_75t_L g1519 ( 
.A(n_1280),
.Y(n_1519)
);

INVx1_ASAP7_75t_L g1520 ( 
.A(n_1398),
.Y(n_1520)
);

OAI21xp5_ASAP7_75t_L g1521 ( 
.A1(n_1397),
.A2(n_1433),
.B(n_1423),
.Y(n_1521)
);

INVx1_ASAP7_75t_L g1522 ( 
.A(n_1376),
.Y(n_1522)
);

CKINVDCx11_ASAP7_75t_R g1523 ( 
.A(n_1401),
.Y(n_1523)
);

OAI22xp5_ASAP7_75t_SL g1524 ( 
.A1(n_1301),
.A2(n_1359),
.B1(n_1400),
.B2(n_1375),
.Y(n_1524)
);

INVx1_ASAP7_75t_L g1525 ( 
.A(n_1359),
.Y(n_1525)
);

BUFx6f_ASAP7_75t_L g1526 ( 
.A(n_1371),
.Y(n_1526)
);

AOI22xp33_ASAP7_75t_L g1527 ( 
.A1(n_1407),
.A2(n_1419),
.B1(n_1418),
.B2(n_1387),
.Y(n_1527)
);

AOI22xp33_ASAP7_75t_L g1528 ( 
.A1(n_1389),
.A2(n_1276),
.B1(n_1303),
.B2(n_1298),
.Y(n_1528)
);

NAND2xp5_ASAP7_75t_L g1529 ( 
.A(n_1359),
.B(n_1427),
.Y(n_1529)
);

CKINVDCx6p67_ASAP7_75t_R g1530 ( 
.A(n_1400),
.Y(n_1530)
);

INVx1_ASAP7_75t_L g1531 ( 
.A(n_1375),
.Y(n_1531)
);

OAI22xp33_ASAP7_75t_L g1532 ( 
.A1(n_1375),
.A2(n_1273),
.B1(n_1400),
.B2(n_1412),
.Y(n_1532)
);

INVxp67_ASAP7_75t_L g1533 ( 
.A(n_1288),
.Y(n_1533)
);

INVx1_ASAP7_75t_L g1534 ( 
.A(n_1412),
.Y(n_1534)
);

INVx1_ASAP7_75t_L g1535 ( 
.A(n_1427),
.Y(n_1535)
);

AOI22xp33_ASAP7_75t_L g1536 ( 
.A1(n_1294),
.A2(n_1295),
.B1(n_1429),
.B2(n_1287),
.Y(n_1536)
);

AOI22xp33_ASAP7_75t_L g1537 ( 
.A1(n_1273),
.A2(n_1178),
.B1(n_1421),
.B2(n_1410),
.Y(n_1537)
);

INVx1_ASAP7_75t_L g1538 ( 
.A(n_1427),
.Y(n_1538)
);

BUFx3_ASAP7_75t_L g1539 ( 
.A(n_1307),
.Y(n_1539)
);

AOI22xp33_ASAP7_75t_L g1540 ( 
.A1(n_1273),
.A2(n_1178),
.B1(n_1421),
.B2(n_1410),
.Y(n_1540)
);

INVx8_ASAP7_75t_L g1541 ( 
.A(n_1307),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_1307),
.Y(n_1542)
);

BUFx3_ASAP7_75t_L g1543 ( 
.A(n_1279),
.Y(n_1543)
);

AOI22xp33_ASAP7_75t_SL g1544 ( 
.A1(n_1349),
.A2(n_1178),
.B1(n_782),
.B2(n_536),
.Y(n_1544)
);

AOI22xp33_ASAP7_75t_L g1545 ( 
.A1(n_1410),
.A2(n_1178),
.B1(n_1421),
.B2(n_782),
.Y(n_1545)
);

INVx6_ASAP7_75t_L g1546 ( 
.A(n_1279),
.Y(n_1546)
);

BUFx4f_ASAP7_75t_SL g1547 ( 
.A(n_1408),
.Y(n_1547)
);

AND2x2_ASAP7_75t_L g1548 ( 
.A(n_1425),
.B(n_1430),
.Y(n_1548)
);

AOI22xp33_ASAP7_75t_SL g1549 ( 
.A1(n_1349),
.A2(n_1178),
.B1(n_782),
.B2(n_536),
.Y(n_1549)
);

INVx4_ASAP7_75t_L g1550 ( 
.A(n_1302),
.Y(n_1550)
);

INVx2_ASAP7_75t_L g1551 ( 
.A(n_1385),
.Y(n_1551)
);

OAI21xp5_ASAP7_75t_SL g1552 ( 
.A1(n_1410),
.A2(n_1178),
.B(n_782),
.Y(n_1552)
);

AOI22xp33_ASAP7_75t_L g1553 ( 
.A1(n_1410),
.A2(n_1178),
.B1(n_1421),
.B2(n_782),
.Y(n_1553)
);

INVx8_ASAP7_75t_L g1554 ( 
.A(n_1290),
.Y(n_1554)
);

INVx2_ASAP7_75t_L g1555 ( 
.A(n_1385),
.Y(n_1555)
);

INVx1_ASAP7_75t_L g1556 ( 
.A(n_1304),
.Y(n_1556)
);

INVx1_ASAP7_75t_L g1557 ( 
.A(n_1304),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_1304),
.Y(n_1558)
);

HB1xp67_ASAP7_75t_L g1559 ( 
.A(n_1324),
.Y(n_1559)
);

OAI22xp33_ASAP7_75t_L g1560 ( 
.A1(n_1410),
.A2(n_1421),
.B1(n_896),
.B2(n_782),
.Y(n_1560)
);

INVx1_ASAP7_75t_SL g1561 ( 
.A(n_1314),
.Y(n_1561)
);

AOI22xp33_ASAP7_75t_L g1562 ( 
.A1(n_1410),
.A2(n_1178),
.B1(n_1421),
.B2(n_782),
.Y(n_1562)
);

INVx3_ASAP7_75t_L g1563 ( 
.A(n_1347),
.Y(n_1563)
);

CKINVDCx5p33_ASAP7_75t_R g1564 ( 
.A(n_1319),
.Y(n_1564)
);

OAI22xp33_ASAP7_75t_L g1565 ( 
.A1(n_1410),
.A2(n_1421),
.B1(n_896),
.B2(n_782),
.Y(n_1565)
);

INVx2_ASAP7_75t_L g1566 ( 
.A(n_1385),
.Y(n_1566)
);

AOI22xp33_ASAP7_75t_L g1567 ( 
.A1(n_1410),
.A2(n_1178),
.B1(n_1421),
.B2(n_782),
.Y(n_1567)
);

INVx1_ASAP7_75t_L g1568 ( 
.A(n_1304),
.Y(n_1568)
);

AOI22xp33_ASAP7_75t_L g1569 ( 
.A1(n_1410),
.A2(n_1178),
.B1(n_1421),
.B2(n_782),
.Y(n_1569)
);

AOI22xp33_ASAP7_75t_SL g1570 ( 
.A1(n_1349),
.A2(n_1178),
.B1(n_782),
.B2(n_536),
.Y(n_1570)
);

AOI22xp33_ASAP7_75t_SL g1571 ( 
.A1(n_1349),
.A2(n_1178),
.B1(n_782),
.B2(n_536),
.Y(n_1571)
);

NAND2xp5_ASAP7_75t_L g1572 ( 
.A(n_1424),
.B(n_1436),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_1304),
.Y(n_1573)
);

OAI22xp33_ASAP7_75t_L g1574 ( 
.A1(n_1410),
.A2(n_1421),
.B1(n_896),
.B2(n_782),
.Y(n_1574)
);

NAND2xp5_ASAP7_75t_L g1575 ( 
.A(n_1424),
.B(n_1436),
.Y(n_1575)
);

AOI22xp33_ASAP7_75t_SL g1576 ( 
.A1(n_1349),
.A2(n_1178),
.B1(n_782),
.B2(n_536),
.Y(n_1576)
);

NAND2xp5_ASAP7_75t_L g1577 ( 
.A(n_1424),
.B(n_1436),
.Y(n_1577)
);

INVx2_ASAP7_75t_SL g1578 ( 
.A(n_1279),
.Y(n_1578)
);

BUFx4_ASAP7_75t_SL g1579 ( 
.A(n_1408),
.Y(n_1579)
);

AOI22xp33_ASAP7_75t_SL g1580 ( 
.A1(n_1349),
.A2(n_1178),
.B1(n_782),
.B2(n_536),
.Y(n_1580)
);

INVx1_ASAP7_75t_L g1581 ( 
.A(n_1304),
.Y(n_1581)
);

OAI22xp33_ASAP7_75t_L g1582 ( 
.A1(n_1410),
.A2(n_1421),
.B1(n_896),
.B2(n_782),
.Y(n_1582)
);

INVx1_ASAP7_75t_L g1583 ( 
.A(n_1304),
.Y(n_1583)
);

AOI22xp33_ASAP7_75t_L g1584 ( 
.A1(n_1410),
.A2(n_1178),
.B1(n_1421),
.B2(n_782),
.Y(n_1584)
);

INVx1_ASAP7_75t_SL g1585 ( 
.A(n_1314),
.Y(n_1585)
);

BUFx12f_ASAP7_75t_L g1586 ( 
.A(n_1319),
.Y(n_1586)
);

AOI22xp33_ASAP7_75t_SL g1587 ( 
.A1(n_1349),
.A2(n_1178),
.B1(n_782),
.B2(n_536),
.Y(n_1587)
);

BUFx6f_ASAP7_75t_L g1588 ( 
.A(n_1290),
.Y(n_1588)
);

AOI22xp33_ASAP7_75t_L g1589 ( 
.A1(n_1410),
.A2(n_1178),
.B1(n_1421),
.B2(n_782),
.Y(n_1589)
);

INVx1_ASAP7_75t_SL g1590 ( 
.A(n_1314),
.Y(n_1590)
);

AOI22xp33_ASAP7_75t_L g1591 ( 
.A1(n_1410),
.A2(n_1178),
.B1(n_1421),
.B2(n_782),
.Y(n_1591)
);

INVx4_ASAP7_75t_L g1592 ( 
.A(n_1302),
.Y(n_1592)
);

AND2x2_ASAP7_75t_L g1593 ( 
.A(n_1425),
.B(n_1430),
.Y(n_1593)
);

OAI22xp5_ASAP7_75t_L g1594 ( 
.A1(n_1410),
.A2(n_1421),
.B1(n_782),
.B2(n_1178),
.Y(n_1594)
);

AOI22xp33_ASAP7_75t_L g1595 ( 
.A1(n_1410),
.A2(n_1178),
.B1(n_1421),
.B2(n_782),
.Y(n_1595)
);

AND2x2_ASAP7_75t_L g1596 ( 
.A(n_1425),
.B(n_1430),
.Y(n_1596)
);

NAND2xp5_ASAP7_75t_L g1597 ( 
.A(n_1424),
.B(n_1436),
.Y(n_1597)
);

INVx8_ASAP7_75t_L g1598 ( 
.A(n_1290),
.Y(n_1598)
);

BUFx2_ASAP7_75t_SL g1599 ( 
.A(n_1405),
.Y(n_1599)
);

INVx2_ASAP7_75t_L g1600 ( 
.A(n_1442),
.Y(n_1600)
);

INVx2_ASAP7_75t_L g1601 ( 
.A(n_1442),
.Y(n_1601)
);

INVx2_ASAP7_75t_SL g1602 ( 
.A(n_1480),
.Y(n_1602)
);

INVx2_ASAP7_75t_L g1603 ( 
.A(n_1444),
.Y(n_1603)
);

HB1xp67_ASAP7_75t_L g1604 ( 
.A(n_1559),
.Y(n_1604)
);

INVx1_ASAP7_75t_L g1605 ( 
.A(n_1444),
.Y(n_1605)
);

INVx1_ASAP7_75t_SL g1606 ( 
.A(n_1548),
.Y(n_1606)
);

OAI21xp5_ASAP7_75t_L g1607 ( 
.A1(n_1483),
.A2(n_1594),
.B(n_1552),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_1551),
.Y(n_1608)
);

HB1xp67_ASAP7_75t_L g1609 ( 
.A(n_1485),
.Y(n_1609)
);

INVxp67_ASAP7_75t_L g1610 ( 
.A(n_1593),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_1555),
.Y(n_1611)
);

OA21x2_ASAP7_75t_L g1612 ( 
.A1(n_1520),
.A2(n_1521),
.B(n_1513),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1566),
.Y(n_1613)
);

OAI21xp5_ASAP7_75t_L g1614 ( 
.A1(n_1482),
.A2(n_1565),
.B(n_1560),
.Y(n_1614)
);

OR2x6_ASAP7_75t_L g1615 ( 
.A(n_1541),
.B(n_1486),
.Y(n_1615)
);

AND2x2_ASAP7_75t_L g1616 ( 
.A(n_1443),
.B(n_1537),
.Y(n_1616)
);

BUFx3_ASAP7_75t_L g1617 ( 
.A(n_1523),
.Y(n_1617)
);

HB1xp67_ASAP7_75t_L g1618 ( 
.A(n_1469),
.Y(n_1618)
);

AND2x4_ASAP7_75t_L g1619 ( 
.A(n_1539),
.B(n_1525),
.Y(n_1619)
);

HB1xp67_ASAP7_75t_L g1620 ( 
.A(n_1481),
.Y(n_1620)
);

AND2x4_ASAP7_75t_L g1621 ( 
.A(n_1539),
.B(n_1533),
.Y(n_1621)
);

INVx3_ASAP7_75t_L g1622 ( 
.A(n_1526),
.Y(n_1622)
);

NAND2xp5_ASAP7_75t_L g1623 ( 
.A(n_1572),
.B(n_1575),
.Y(n_1623)
);

INVx2_ASAP7_75t_L g1624 ( 
.A(n_1463),
.Y(n_1624)
);

AND2x2_ASAP7_75t_L g1625 ( 
.A(n_1443),
.B(n_1537),
.Y(n_1625)
);

AND2x4_ASAP7_75t_L g1626 ( 
.A(n_1463),
.B(n_1470),
.Y(n_1626)
);

INVx2_ASAP7_75t_L g1627 ( 
.A(n_1470),
.Y(n_1627)
);

HB1xp67_ASAP7_75t_L g1628 ( 
.A(n_1478),
.Y(n_1628)
);

INVx1_ASAP7_75t_L g1629 ( 
.A(n_1534),
.Y(n_1629)
);

OAI21x1_ASAP7_75t_L g1630 ( 
.A1(n_1536),
.A2(n_1528),
.B(n_1527),
.Y(n_1630)
);

OAI21x1_ASAP7_75t_L g1631 ( 
.A1(n_1536),
.A2(n_1528),
.B(n_1527),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_1535),
.Y(n_1632)
);

INVx1_ASAP7_75t_L g1633 ( 
.A(n_1538),
.Y(n_1633)
);

OAI21x1_ASAP7_75t_L g1634 ( 
.A1(n_1484),
.A2(n_1507),
.B(n_1495),
.Y(n_1634)
);

INVx3_ASAP7_75t_L g1635 ( 
.A(n_1526),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_1531),
.Y(n_1636)
);

NAND2xp5_ASAP7_75t_L g1637 ( 
.A(n_1577),
.B(n_1597),
.Y(n_1637)
);

OAI21x1_ASAP7_75t_L g1638 ( 
.A1(n_1484),
.A2(n_1507),
.B(n_1495),
.Y(n_1638)
);

OAI21x1_ASAP7_75t_L g1639 ( 
.A1(n_1504),
.A2(n_1542),
.B(n_1518),
.Y(n_1639)
);

AND2x2_ASAP7_75t_L g1640 ( 
.A(n_1540),
.B(n_1446),
.Y(n_1640)
);

OAI21x1_ASAP7_75t_L g1641 ( 
.A1(n_1504),
.A2(n_1518),
.B(n_1506),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_1522),
.Y(n_1642)
);

NAND2xp5_ASAP7_75t_L g1643 ( 
.A(n_1476),
.B(n_1459),
.Y(n_1643)
);

INVx2_ASAP7_75t_SL g1644 ( 
.A(n_1480),
.Y(n_1644)
);

HB1xp67_ASAP7_75t_L g1645 ( 
.A(n_1451),
.Y(n_1645)
);

INVx1_ASAP7_75t_L g1646 ( 
.A(n_1529),
.Y(n_1646)
);

INVx1_ASAP7_75t_L g1647 ( 
.A(n_1524),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_1541),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_1541),
.Y(n_1649)
);

OAI21x1_ASAP7_75t_L g1650 ( 
.A1(n_1506),
.A2(n_1496),
.B(n_1492),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_1440),
.Y(n_1651)
);

OR2x2_ASAP7_75t_L g1652 ( 
.A(n_1540),
.B(n_1446),
.Y(n_1652)
);

INVx2_ASAP7_75t_L g1653 ( 
.A(n_1448),
.Y(n_1653)
);

HB1xp67_ASAP7_75t_L g1654 ( 
.A(n_1488),
.Y(n_1654)
);

NAND2xp5_ASAP7_75t_L g1655 ( 
.A(n_1465),
.B(n_1545),
.Y(n_1655)
);

INVx1_ASAP7_75t_L g1656 ( 
.A(n_1462),
.Y(n_1656)
);

AO21x2_ASAP7_75t_L g1657 ( 
.A1(n_1532),
.A2(n_1503),
.B(n_1508),
.Y(n_1657)
);

OR2x2_ASAP7_75t_L g1658 ( 
.A(n_1489),
.B(n_1492),
.Y(n_1658)
);

INVx2_ASAP7_75t_L g1659 ( 
.A(n_1556),
.Y(n_1659)
);

NOR2xp33_ASAP7_75t_L g1660 ( 
.A(n_1596),
.B(n_1501),
.Y(n_1660)
);

NAND2xp5_ASAP7_75t_L g1661 ( 
.A(n_1465),
.B(n_1545),
.Y(n_1661)
);

OAI21x1_ASAP7_75t_L g1662 ( 
.A1(n_1496),
.A2(n_1482),
.B(n_1474),
.Y(n_1662)
);

BUFx6f_ASAP7_75t_L g1663 ( 
.A(n_1523),
.Y(n_1663)
);

OA21x2_ASAP7_75t_L g1664 ( 
.A1(n_1474),
.A2(n_1471),
.B(n_1458),
.Y(n_1664)
);

INVx11_ASAP7_75t_L g1665 ( 
.A(n_1586),
.Y(n_1665)
);

OAI21xp5_ASAP7_75t_L g1666 ( 
.A1(n_1574),
.A2(n_1582),
.B(n_1456),
.Y(n_1666)
);

AND2x2_ASAP7_75t_L g1667 ( 
.A(n_1515),
.B(n_1557),
.Y(n_1667)
);

INVx1_ASAP7_75t_L g1668 ( 
.A(n_1558),
.Y(n_1668)
);

AND2x2_ASAP7_75t_L g1669 ( 
.A(n_1568),
.B(n_1573),
.Y(n_1669)
);

AND2x4_ASAP7_75t_L g1670 ( 
.A(n_1498),
.B(n_1445),
.Y(n_1670)
);

INVx1_ASAP7_75t_L g1671 ( 
.A(n_1581),
.Y(n_1671)
);

INVx6_ASAP7_75t_L g1672 ( 
.A(n_1439),
.Y(n_1672)
);

INVx2_ASAP7_75t_L g1673 ( 
.A(n_1583),
.Y(n_1673)
);

INVxp67_ASAP7_75t_L g1674 ( 
.A(n_1460),
.Y(n_1674)
);

BUFx2_ASAP7_75t_L g1675 ( 
.A(n_1500),
.Y(n_1675)
);

BUFx2_ASAP7_75t_L g1676 ( 
.A(n_1530),
.Y(n_1676)
);

INVx2_ASAP7_75t_L g1677 ( 
.A(n_1445),
.Y(n_1677)
);

OA21x2_ASAP7_75t_L g1678 ( 
.A1(n_1471),
.A2(n_1458),
.B(n_1489),
.Y(n_1678)
);

HB1xp67_ASAP7_75t_L g1679 ( 
.A(n_1561),
.Y(n_1679)
);

INVx1_ASAP7_75t_L g1680 ( 
.A(n_1447),
.Y(n_1680)
);

OA21x2_ASAP7_75t_L g1681 ( 
.A1(n_1553),
.A2(n_1562),
.B(n_1569),
.Y(n_1681)
);

INVx1_ASAP7_75t_L g1682 ( 
.A(n_1447),
.Y(n_1682)
);

OAI21xp33_ASAP7_75t_SL g1683 ( 
.A1(n_1553),
.A2(n_1569),
.B(n_1595),
.Y(n_1683)
);

HB1xp67_ASAP7_75t_L g1684 ( 
.A(n_1585),
.Y(n_1684)
);

HB1xp67_ASAP7_75t_L g1685 ( 
.A(n_1590),
.Y(n_1685)
);

INVx1_ASAP7_75t_L g1686 ( 
.A(n_1491),
.Y(n_1686)
);

O2A1O1Ixp33_ASAP7_75t_L g1687 ( 
.A1(n_1453),
.A2(n_1454),
.B(n_1589),
.C(n_1562),
.Y(n_1687)
);

INVx1_ASAP7_75t_L g1688 ( 
.A(n_1512),
.Y(n_1688)
);

NAND2xp5_ASAP7_75t_L g1689 ( 
.A(n_1567),
.B(n_1589),
.Y(n_1689)
);

INVx1_ASAP7_75t_L g1690 ( 
.A(n_1514),
.Y(n_1690)
);

CKINVDCx6p67_ASAP7_75t_R g1691 ( 
.A(n_1511),
.Y(n_1691)
);

BUFx6f_ASAP7_75t_L g1692 ( 
.A(n_1588),
.Y(n_1692)
);

INVx3_ASAP7_75t_L g1693 ( 
.A(n_1519),
.Y(n_1693)
);

INVx1_ASAP7_75t_L g1694 ( 
.A(n_1519),
.Y(n_1694)
);

AND2x2_ASAP7_75t_L g1695 ( 
.A(n_1567),
.B(n_1584),
.Y(n_1695)
);

AND2x4_ASAP7_75t_SL g1696 ( 
.A(n_1466),
.B(n_1588),
.Y(n_1696)
);

INVx1_ASAP7_75t_L g1697 ( 
.A(n_1499),
.Y(n_1697)
);

INVx1_ASAP7_75t_L g1698 ( 
.A(n_1563),
.Y(n_1698)
);

AND2x2_ASAP7_75t_L g1699 ( 
.A(n_1584),
.B(n_1591),
.Y(n_1699)
);

INVxp67_ASAP7_75t_L g1700 ( 
.A(n_1475),
.Y(n_1700)
);

NOR2xp33_ASAP7_75t_L g1701 ( 
.A(n_1472),
.B(n_1493),
.Y(n_1701)
);

INVx2_ASAP7_75t_SL g1702 ( 
.A(n_1480),
.Y(n_1702)
);

NAND2xp5_ASAP7_75t_L g1703 ( 
.A(n_1591),
.B(n_1595),
.Y(n_1703)
);

NAND2xp5_ASAP7_75t_L g1704 ( 
.A(n_1544),
.B(n_1571),
.Y(n_1704)
);

INVx2_ASAP7_75t_L g1705 ( 
.A(n_1588),
.Y(n_1705)
);

AND2x2_ASAP7_75t_L g1706 ( 
.A(n_1549),
.B(n_1576),
.Y(n_1706)
);

INVx1_ASAP7_75t_L g1707 ( 
.A(n_1505),
.Y(n_1707)
);

INVx2_ASAP7_75t_L g1708 ( 
.A(n_1588),
.Y(n_1708)
);

OAI21xp5_ASAP7_75t_L g1709 ( 
.A1(n_1570),
.A2(n_1580),
.B(n_1587),
.Y(n_1709)
);

INVx2_ASAP7_75t_L g1710 ( 
.A(n_1468),
.Y(n_1710)
);

OA21x2_ASAP7_75t_L g1711 ( 
.A1(n_1517),
.A2(n_1441),
.B(n_1578),
.Y(n_1711)
);

BUFx2_ASAP7_75t_L g1712 ( 
.A(n_1479),
.Y(n_1712)
);

INVx3_ASAP7_75t_L g1713 ( 
.A(n_1554),
.Y(n_1713)
);

INVx2_ASAP7_75t_L g1714 ( 
.A(n_1554),
.Y(n_1714)
);

INVx1_ASAP7_75t_L g1715 ( 
.A(n_1509),
.Y(n_1715)
);

INVx1_ASAP7_75t_L g1716 ( 
.A(n_1598),
.Y(n_1716)
);

HB1xp67_ASAP7_75t_L g1717 ( 
.A(n_1510),
.Y(n_1717)
);

CKINVDCx5p33_ASAP7_75t_R g1718 ( 
.A(n_1579),
.Y(n_1718)
);

CKINVDCx5p33_ASAP7_75t_R g1719 ( 
.A(n_1564),
.Y(n_1719)
);

AOI22xp33_ASAP7_75t_L g1720 ( 
.A1(n_1473),
.A2(n_1464),
.B1(n_1479),
.B2(n_1599),
.Y(n_1720)
);

OAI21xp5_ASAP7_75t_L g1721 ( 
.A1(n_1487),
.A2(n_1502),
.B(n_1439),
.Y(n_1721)
);

AOI21x1_ASAP7_75t_L g1722 ( 
.A1(n_1598),
.A2(n_1510),
.B(n_1516),
.Y(n_1722)
);

NAND2xp5_ASAP7_75t_L g1723 ( 
.A(n_1455),
.B(n_1543),
.Y(n_1723)
);

AND2x2_ASAP7_75t_L g1724 ( 
.A(n_1502),
.B(n_1543),
.Y(n_1724)
);

HB1xp67_ASAP7_75t_L g1725 ( 
.A(n_1510),
.Y(n_1725)
);

HB1xp67_ASAP7_75t_L g1726 ( 
.A(n_1455),
.Y(n_1726)
);

INVx1_ASAP7_75t_L g1727 ( 
.A(n_1439),
.Y(n_1727)
);

BUFx3_ASAP7_75t_L g1728 ( 
.A(n_1516),
.Y(n_1728)
);

OAI211xp5_ASAP7_75t_L g1729 ( 
.A1(n_1709),
.A2(n_1494),
.B(n_1473),
.C(n_1464),
.Y(n_1729)
);

AND2x2_ASAP7_75t_L g1730 ( 
.A(n_1628),
.B(n_1461),
.Y(n_1730)
);

OAI21x1_ASAP7_75t_SL g1731 ( 
.A1(n_1687),
.A2(n_1666),
.B(n_1607),
.Y(n_1731)
);

NAND2xp5_ASAP7_75t_L g1732 ( 
.A(n_1646),
.B(n_1550),
.Y(n_1732)
);

AND2x2_ASAP7_75t_L g1733 ( 
.A(n_1660),
.B(n_1461),
.Y(n_1733)
);

AND2x2_ASAP7_75t_L g1734 ( 
.A(n_1609),
.B(n_1461),
.Y(n_1734)
);

AND2x4_ASAP7_75t_L g1735 ( 
.A(n_1626),
.B(n_1550),
.Y(n_1735)
);

AND2x4_ASAP7_75t_L g1736 ( 
.A(n_1626),
.B(n_1550),
.Y(n_1736)
);

AOI221xp5_ASAP7_75t_L g1737 ( 
.A1(n_1683),
.A2(n_1497),
.B1(n_1592),
.B2(n_1449),
.C(n_1477),
.Y(n_1737)
);

OA21x2_ASAP7_75t_L g1738 ( 
.A1(n_1641),
.A2(n_1466),
.B(n_1450),
.Y(n_1738)
);

INVx1_ASAP7_75t_L g1739 ( 
.A(n_1651),
.Y(n_1739)
);

CKINVDCx20_ASAP7_75t_R g1740 ( 
.A(n_1718),
.Y(n_1740)
);

O2A1O1Ixp5_ASAP7_75t_L g1741 ( 
.A1(n_1614),
.A2(n_1592),
.B(n_1466),
.C(n_1457),
.Y(n_1741)
);

AND2x4_ASAP7_75t_L g1742 ( 
.A(n_1626),
.B(n_1449),
.Y(n_1742)
);

INVx1_ASAP7_75t_L g1743 ( 
.A(n_1651),
.Y(n_1743)
);

OR2x6_ASAP7_75t_L g1744 ( 
.A(n_1615),
.B(n_1450),
.Y(n_1744)
);

OAI21xp5_ASAP7_75t_L g1745 ( 
.A1(n_1683),
.A2(n_1477),
.B(n_1457),
.Y(n_1745)
);

OA21x2_ASAP7_75t_L g1746 ( 
.A1(n_1641),
.A2(n_1450),
.B(n_1546),
.Y(n_1746)
);

AND2x2_ASAP7_75t_L g1747 ( 
.A(n_1606),
.B(n_1457),
.Y(n_1747)
);

AO32x2_ASAP7_75t_L g1748 ( 
.A1(n_1647),
.A2(n_1452),
.A3(n_1490),
.B1(n_1511),
.B2(n_1467),
.Y(n_1748)
);

AND2x4_ASAP7_75t_SL g1749 ( 
.A(n_1663),
.B(n_1691),
.Y(n_1749)
);

AND2x4_ASAP7_75t_L g1750 ( 
.A(n_1626),
.B(n_1490),
.Y(n_1750)
);

AND2x2_ASAP7_75t_L g1751 ( 
.A(n_1610),
.B(n_1586),
.Y(n_1751)
);

CKINVDCx5p33_ASAP7_75t_R g1752 ( 
.A(n_1719),
.Y(n_1752)
);

AOI21xp5_ASAP7_75t_L g1753 ( 
.A1(n_1664),
.A2(n_1547),
.B(n_1612),
.Y(n_1753)
);

AOI221xp5_ASAP7_75t_L g1754 ( 
.A1(n_1706),
.A2(n_1704),
.B1(n_1654),
.B2(n_1655),
.C(n_1661),
.Y(n_1754)
);

INVx2_ASAP7_75t_L g1755 ( 
.A(n_1669),
.Y(n_1755)
);

BUFx2_ASAP7_75t_L g1756 ( 
.A(n_1663),
.Y(n_1756)
);

HB1xp67_ASAP7_75t_L g1757 ( 
.A(n_1604),
.Y(n_1757)
);

OR2x6_ASAP7_75t_L g1758 ( 
.A(n_1615),
.B(n_1662),
.Y(n_1758)
);

AND2x2_ASAP7_75t_L g1759 ( 
.A(n_1686),
.B(n_1670),
.Y(n_1759)
);

AND2x2_ASAP7_75t_L g1760 ( 
.A(n_1686),
.B(n_1670),
.Y(n_1760)
);

AND2x2_ASAP7_75t_L g1761 ( 
.A(n_1670),
.B(n_1667),
.Y(n_1761)
);

OR2x6_ASAP7_75t_L g1762 ( 
.A(n_1615),
.B(n_1662),
.Y(n_1762)
);

A2O1A1Ixp33_ASAP7_75t_L g1763 ( 
.A1(n_1652),
.A2(n_1640),
.B(n_1695),
.C(n_1699),
.Y(n_1763)
);

OAI22xp5_ASAP7_75t_L g1764 ( 
.A1(n_1652),
.A2(n_1703),
.B1(n_1689),
.B2(n_1643),
.Y(n_1764)
);

AOI221xp5_ASAP7_75t_L g1765 ( 
.A1(n_1616),
.A2(n_1625),
.B1(n_1640),
.B2(n_1695),
.C(n_1699),
.Y(n_1765)
);

OAI21xp5_ASAP7_75t_L g1766 ( 
.A1(n_1650),
.A2(n_1664),
.B(n_1678),
.Y(n_1766)
);

AND2x4_ASAP7_75t_L g1767 ( 
.A(n_1648),
.B(n_1649),
.Y(n_1767)
);

A2O1A1Ixp33_ASAP7_75t_L g1768 ( 
.A1(n_1616),
.A2(n_1625),
.B(n_1650),
.C(n_1617),
.Y(n_1768)
);

AND2x4_ASAP7_75t_L g1769 ( 
.A(n_1648),
.B(n_1649),
.Y(n_1769)
);

NOR2xp33_ASAP7_75t_L g1770 ( 
.A(n_1623),
.B(n_1637),
.Y(n_1770)
);

HB1xp67_ASAP7_75t_L g1771 ( 
.A(n_1675),
.Y(n_1771)
);

NAND2xp5_ASAP7_75t_L g1772 ( 
.A(n_1659),
.B(n_1656),
.Y(n_1772)
);

AND2x4_ASAP7_75t_L g1773 ( 
.A(n_1676),
.B(n_1653),
.Y(n_1773)
);

INVxp67_ASAP7_75t_L g1774 ( 
.A(n_1679),
.Y(n_1774)
);

AND2x4_ASAP7_75t_L g1775 ( 
.A(n_1676),
.B(n_1653),
.Y(n_1775)
);

OR2x2_ASAP7_75t_L g1776 ( 
.A(n_1658),
.B(n_1673),
.Y(n_1776)
);

OAI21xp5_ASAP7_75t_L g1777 ( 
.A1(n_1664),
.A2(n_1678),
.B(n_1707),
.Y(n_1777)
);

NOR2xp33_ASAP7_75t_L g1778 ( 
.A(n_1701),
.B(n_1700),
.Y(n_1778)
);

AOI21xp5_ASAP7_75t_L g1779 ( 
.A1(n_1612),
.A2(n_1678),
.B(n_1675),
.Y(n_1779)
);

NAND2xp5_ASAP7_75t_L g1780 ( 
.A(n_1668),
.B(n_1671),
.Y(n_1780)
);

INVxp67_ASAP7_75t_L g1781 ( 
.A(n_1684),
.Y(n_1781)
);

A2O1A1Ixp33_ASAP7_75t_L g1782 ( 
.A1(n_1617),
.A2(n_1688),
.B(n_1690),
.C(n_1663),
.Y(n_1782)
);

INVx4_ASAP7_75t_L g1783 ( 
.A(n_1663),
.Y(n_1783)
);

AOI211xp5_ASAP7_75t_L g1784 ( 
.A1(n_1617),
.A2(n_1688),
.B(n_1663),
.C(n_1685),
.Y(n_1784)
);

OR2x2_ASAP7_75t_L g1785 ( 
.A(n_1620),
.B(n_1668),
.Y(n_1785)
);

AND2x2_ASAP7_75t_L g1786 ( 
.A(n_1645),
.B(n_1724),
.Y(n_1786)
);

OR2x2_ASAP7_75t_L g1787 ( 
.A(n_1671),
.B(n_1618),
.Y(n_1787)
);

AOI22xp5_ASAP7_75t_L g1788 ( 
.A1(n_1681),
.A2(n_1663),
.B1(n_1720),
.B2(n_1615),
.Y(n_1788)
);

OAI21xp5_ASAP7_75t_L g1789 ( 
.A1(n_1681),
.A2(n_1634),
.B(n_1638),
.Y(n_1789)
);

AND2x2_ASAP7_75t_L g1790 ( 
.A(n_1724),
.B(n_1726),
.Y(n_1790)
);

OAI21xp5_ASAP7_75t_L g1791 ( 
.A1(n_1681),
.A2(n_1638),
.B(n_1634),
.Y(n_1791)
);

OAI21xp5_ASAP7_75t_L g1792 ( 
.A1(n_1681),
.A2(n_1612),
.B(n_1631),
.Y(n_1792)
);

INVx1_ASAP7_75t_L g1793 ( 
.A(n_1636),
.Y(n_1793)
);

AND2x2_ASAP7_75t_L g1794 ( 
.A(n_1615),
.B(n_1674),
.Y(n_1794)
);

AND2x2_ASAP7_75t_L g1795 ( 
.A(n_1624),
.B(n_1627),
.Y(n_1795)
);

NAND2xp5_ASAP7_75t_L g1796 ( 
.A(n_1627),
.B(n_1605),
.Y(n_1796)
);

A2O1A1Ixp33_ASAP7_75t_L g1797 ( 
.A1(n_1639),
.A2(n_1631),
.B(n_1630),
.C(n_1721),
.Y(n_1797)
);

AND2x2_ASAP7_75t_L g1798 ( 
.A(n_1705),
.B(n_1708),
.Y(n_1798)
);

AOI22xp5_ASAP7_75t_L g1799 ( 
.A1(n_1691),
.A2(n_1712),
.B1(n_1657),
.B2(n_1728),
.Y(n_1799)
);

AO32x2_ASAP7_75t_L g1800 ( 
.A1(n_1602),
.A2(n_1644),
.A3(n_1702),
.B1(n_1657),
.B2(n_1642),
.Y(n_1800)
);

OA21x2_ASAP7_75t_L g1801 ( 
.A1(n_1639),
.A2(n_1630),
.B(n_1642),
.Y(n_1801)
);

OAI22xp5_ASAP7_75t_L g1802 ( 
.A1(n_1712),
.A2(n_1711),
.B1(n_1723),
.B2(n_1715),
.Y(n_1802)
);

NAND2xp5_ASAP7_75t_L g1803 ( 
.A(n_1605),
.B(n_1608),
.Y(n_1803)
);

INVx3_ASAP7_75t_L g1804 ( 
.A(n_1692),
.Y(n_1804)
);

OA21x2_ASAP7_75t_L g1805 ( 
.A1(n_1629),
.A2(n_1632),
.B(n_1633),
.Y(n_1805)
);

AND2x2_ASAP7_75t_L g1806 ( 
.A(n_1705),
.B(n_1708),
.Y(n_1806)
);

OAI21x1_ASAP7_75t_L g1807 ( 
.A1(n_1693),
.A2(n_1622),
.B(n_1635),
.Y(n_1807)
);

INVxp67_ASAP7_75t_L g1808 ( 
.A(n_1717),
.Y(n_1808)
);

AOI221xp5_ASAP7_75t_L g1809 ( 
.A1(n_1657),
.A2(n_1682),
.B1(n_1680),
.B2(n_1677),
.C(n_1629),
.Y(n_1809)
);

O2A1O1Ixp33_ASAP7_75t_SL g1810 ( 
.A1(n_1716),
.A2(n_1715),
.B(n_1602),
.C(n_1644),
.Y(n_1810)
);

OR2x6_ASAP7_75t_L g1811 ( 
.A(n_1711),
.B(n_1619),
.Y(n_1811)
);

NAND2xp5_ASAP7_75t_SL g1812 ( 
.A(n_1770),
.B(n_1714),
.Y(n_1812)
);

OR2x2_ASAP7_75t_L g1813 ( 
.A(n_1811),
.B(n_1600),
.Y(n_1813)
);

INVx1_ASAP7_75t_L g1814 ( 
.A(n_1805),
.Y(n_1814)
);

INVx1_ASAP7_75t_L g1815 ( 
.A(n_1805),
.Y(n_1815)
);

INVx2_ASAP7_75t_L g1816 ( 
.A(n_1793),
.Y(n_1816)
);

AND2x2_ASAP7_75t_L g1817 ( 
.A(n_1792),
.B(n_1600),
.Y(n_1817)
);

AND2x4_ASAP7_75t_L g1818 ( 
.A(n_1811),
.B(n_1622),
.Y(n_1818)
);

INVx2_ASAP7_75t_L g1819 ( 
.A(n_1739),
.Y(n_1819)
);

OAI22xp5_ASAP7_75t_L g1820 ( 
.A1(n_1754),
.A2(n_1763),
.B1(n_1737),
.B2(n_1745),
.Y(n_1820)
);

AND2x4_ASAP7_75t_L g1821 ( 
.A(n_1811),
.B(n_1622),
.Y(n_1821)
);

NAND2x1_ASAP7_75t_L g1822 ( 
.A(n_1744),
.B(n_1711),
.Y(n_1822)
);

OAI22xp5_ASAP7_75t_L g1823 ( 
.A1(n_1737),
.A2(n_1711),
.B1(n_1696),
.B2(n_1672),
.Y(n_1823)
);

AND2x2_ASAP7_75t_L g1824 ( 
.A(n_1792),
.B(n_1789),
.Y(n_1824)
);

BUFx2_ASAP7_75t_L g1825 ( 
.A(n_1800),
.Y(n_1825)
);

INVx2_ASAP7_75t_L g1826 ( 
.A(n_1743),
.Y(n_1826)
);

NAND2xp5_ASAP7_75t_L g1827 ( 
.A(n_1776),
.B(n_1755),
.Y(n_1827)
);

HB1xp67_ASAP7_75t_L g1828 ( 
.A(n_1771),
.Y(n_1828)
);

NOR2x1_ASAP7_75t_L g1829 ( 
.A(n_1802),
.B(n_1694),
.Y(n_1829)
);

BUFx2_ASAP7_75t_L g1830 ( 
.A(n_1800),
.Y(n_1830)
);

AND2x2_ASAP7_75t_L g1831 ( 
.A(n_1791),
.B(n_1766),
.Y(n_1831)
);

AND2x4_ASAP7_75t_L g1832 ( 
.A(n_1807),
.B(n_1622),
.Y(n_1832)
);

OR2x2_ASAP7_75t_L g1833 ( 
.A(n_1766),
.B(n_1601),
.Y(n_1833)
);

AND2x2_ASAP7_75t_L g1834 ( 
.A(n_1801),
.B(n_1601),
.Y(n_1834)
);

BUFx2_ASAP7_75t_L g1835 ( 
.A(n_1800),
.Y(n_1835)
);

NOR2xp33_ASAP7_75t_L g1836 ( 
.A(n_1729),
.B(n_1728),
.Y(n_1836)
);

AOI22xp33_ASAP7_75t_L g1837 ( 
.A1(n_1731),
.A2(n_1728),
.B1(n_1680),
.B2(n_1682),
.Y(n_1837)
);

NAND2xp5_ASAP7_75t_L g1838 ( 
.A(n_1757),
.B(n_1613),
.Y(n_1838)
);

BUFx3_ASAP7_75t_L g1839 ( 
.A(n_1749),
.Y(n_1839)
);

BUFx2_ASAP7_75t_L g1840 ( 
.A(n_1759),
.Y(n_1840)
);

NOR2x1_ASAP7_75t_L g1841 ( 
.A(n_1802),
.B(n_1694),
.Y(n_1841)
);

OR2x2_ASAP7_75t_L g1842 ( 
.A(n_1779),
.B(n_1603),
.Y(n_1842)
);

INVx1_ASAP7_75t_L g1843 ( 
.A(n_1780),
.Y(n_1843)
);

NAND2xp5_ASAP7_75t_L g1844 ( 
.A(n_1760),
.B(n_1611),
.Y(n_1844)
);

AND2x2_ASAP7_75t_L g1845 ( 
.A(n_1758),
.B(n_1762),
.Y(n_1845)
);

INVx1_ASAP7_75t_L g1846 ( 
.A(n_1780),
.Y(n_1846)
);

INVx2_ASAP7_75t_L g1847 ( 
.A(n_1795),
.Y(n_1847)
);

AND2x4_ASAP7_75t_SL g1848 ( 
.A(n_1744),
.B(n_1619),
.Y(n_1848)
);

AOI22xp33_ASAP7_75t_L g1849 ( 
.A1(n_1745),
.A2(n_1619),
.B1(n_1677),
.B2(n_1621),
.Y(n_1849)
);

INVx1_ASAP7_75t_L g1850 ( 
.A(n_1772),
.Y(n_1850)
);

BUFx3_ASAP7_75t_L g1851 ( 
.A(n_1756),
.Y(n_1851)
);

AOI22xp33_ASAP7_75t_L g1852 ( 
.A1(n_1764),
.A2(n_1621),
.B1(n_1725),
.B2(n_1710),
.Y(n_1852)
);

INVx2_ASAP7_75t_SL g1853 ( 
.A(n_1773),
.Y(n_1853)
);

OAI21xp33_ASAP7_75t_L g1854 ( 
.A1(n_1768),
.A2(n_1696),
.B(n_1727),
.Y(n_1854)
);

OAI221xp5_ASAP7_75t_L g1855 ( 
.A1(n_1820),
.A2(n_1799),
.B1(n_1788),
.B2(n_1784),
.C(n_1782),
.Y(n_1855)
);

AOI221xp5_ASAP7_75t_L g1856 ( 
.A1(n_1820),
.A2(n_1764),
.B1(n_1765),
.B2(n_1753),
.C(n_1781),
.Y(n_1856)
);

NAND4xp25_ASAP7_75t_SL g1857 ( 
.A(n_1829),
.B(n_1784),
.C(n_1809),
.D(n_1797),
.Y(n_1857)
);

OR2x2_ASAP7_75t_L g1858 ( 
.A(n_1833),
.B(n_1785),
.Y(n_1858)
);

INVx1_ASAP7_75t_L g1859 ( 
.A(n_1816),
.Y(n_1859)
);

HB1xp67_ASAP7_75t_L g1860 ( 
.A(n_1828),
.Y(n_1860)
);

AOI211xp5_ASAP7_75t_L g1861 ( 
.A1(n_1854),
.A2(n_1777),
.B(n_1778),
.C(n_1794),
.Y(n_1861)
);

INVx1_ASAP7_75t_L g1862 ( 
.A(n_1816),
.Y(n_1862)
);

AND2x2_ASAP7_75t_L g1863 ( 
.A(n_1840),
.B(n_1761),
.Y(n_1863)
);

AND2x4_ASAP7_75t_L g1864 ( 
.A(n_1818),
.B(n_1744),
.Y(n_1864)
);

INVx1_ASAP7_75t_L g1865 ( 
.A(n_1816),
.Y(n_1865)
);

NAND3xp33_ASAP7_75t_SL g1866 ( 
.A(n_1854),
.B(n_1741),
.C(n_1777),
.Y(n_1866)
);

AND2x2_ASAP7_75t_L g1867 ( 
.A(n_1845),
.B(n_1738),
.Y(n_1867)
);

AND2x4_ASAP7_75t_L g1868 ( 
.A(n_1818),
.B(n_1773),
.Y(n_1868)
);

INVx3_ASAP7_75t_L g1869 ( 
.A(n_1832),
.Y(n_1869)
);

INVx2_ASAP7_75t_L g1870 ( 
.A(n_1814),
.Y(n_1870)
);

NAND2xp5_ASAP7_75t_L g1871 ( 
.A(n_1843),
.B(n_1774),
.Y(n_1871)
);

OR2x2_ASAP7_75t_L g1872 ( 
.A(n_1833),
.B(n_1787),
.Y(n_1872)
);

HB1xp67_ASAP7_75t_L g1873 ( 
.A(n_1828),
.Y(n_1873)
);

INVx1_ASAP7_75t_L g1874 ( 
.A(n_1819),
.Y(n_1874)
);

INVx5_ASAP7_75t_L g1875 ( 
.A(n_1834),
.Y(n_1875)
);

BUFx3_ASAP7_75t_L g1876 ( 
.A(n_1839),
.Y(n_1876)
);

INVxp67_ASAP7_75t_L g1877 ( 
.A(n_1812),
.Y(n_1877)
);

AOI322xp5_ASAP7_75t_L g1878 ( 
.A1(n_1829),
.A2(n_1809),
.A3(n_1742),
.B1(n_1733),
.B2(n_1747),
.C1(n_1751),
.C2(n_1786),
.Y(n_1878)
);

OAI22xp5_ASAP7_75t_L g1879 ( 
.A1(n_1849),
.A2(n_1783),
.B1(n_1808),
.B2(n_1742),
.Y(n_1879)
);

OAI322xp33_ASAP7_75t_L g1880 ( 
.A1(n_1833),
.A2(n_1732),
.A3(n_1796),
.B1(n_1803),
.B2(n_1633),
.C1(n_1734),
.C2(n_1730),
.Y(n_1880)
);

NAND4xp25_ASAP7_75t_L g1881 ( 
.A(n_1837),
.B(n_1732),
.C(n_1775),
.D(n_1806),
.Y(n_1881)
);

OAI31xp33_ASAP7_75t_L g1882 ( 
.A1(n_1823),
.A2(n_1836),
.A3(n_1831),
.B(n_1824),
.Y(n_1882)
);

INVx2_ASAP7_75t_L g1883 ( 
.A(n_1814),
.Y(n_1883)
);

AND2x2_ASAP7_75t_L g1884 ( 
.A(n_1845),
.B(n_1738),
.Y(n_1884)
);

AND2x2_ASAP7_75t_L g1885 ( 
.A(n_1845),
.B(n_1746),
.Y(n_1885)
);

OAI22xp5_ASAP7_75t_L g1886 ( 
.A1(n_1849),
.A2(n_1769),
.B1(n_1767),
.B2(n_1672),
.Y(n_1886)
);

BUFx3_ASAP7_75t_L g1887 ( 
.A(n_1839),
.Y(n_1887)
);

BUFx6f_ASAP7_75t_L g1888 ( 
.A(n_1839),
.Y(n_1888)
);

NAND2xp5_ASAP7_75t_SL g1889 ( 
.A(n_1841),
.B(n_1775),
.Y(n_1889)
);

OR2x2_ASAP7_75t_L g1890 ( 
.A(n_1827),
.B(n_1746),
.Y(n_1890)
);

OAI221xp5_ASAP7_75t_SL g1891 ( 
.A1(n_1837),
.A2(n_1831),
.B1(n_1824),
.B2(n_1852),
.C(n_1835),
.Y(n_1891)
);

OR2x2_ASAP7_75t_L g1892 ( 
.A(n_1827),
.B(n_1803),
.Y(n_1892)
);

BUFx3_ASAP7_75t_L g1893 ( 
.A(n_1851),
.Y(n_1893)
);

AOI22xp33_ASAP7_75t_L g1894 ( 
.A1(n_1823),
.A2(n_1735),
.B1(n_1736),
.B2(n_1750),
.Y(n_1894)
);

NOR2xp33_ASAP7_75t_L g1895 ( 
.A(n_1838),
.B(n_1752),
.Y(n_1895)
);

OR2x2_ASAP7_75t_L g1896 ( 
.A(n_1847),
.B(n_1790),
.Y(n_1896)
);

INVx2_ASAP7_75t_SL g1897 ( 
.A(n_1851),
.Y(n_1897)
);

OR2x6_ASAP7_75t_SL g1898 ( 
.A(n_1813),
.B(n_1748),
.Y(n_1898)
);

NAND2xp33_ASAP7_75t_R g1899 ( 
.A(n_1831),
.B(n_1798),
.Y(n_1899)
);

AND2x4_ASAP7_75t_L g1900 ( 
.A(n_1818),
.B(n_1804),
.Y(n_1900)
);

XNOR2xp5_ASAP7_75t_L g1901 ( 
.A(n_1841),
.B(n_1740),
.Y(n_1901)
);

OAI22xp5_ASAP7_75t_L g1902 ( 
.A1(n_1848),
.A2(n_1769),
.B1(n_1767),
.B2(n_1672),
.Y(n_1902)
);

OAI211xp5_ASAP7_75t_L g1903 ( 
.A1(n_1824),
.A2(n_1810),
.B(n_1697),
.C(n_1698),
.Y(n_1903)
);

INVx1_ASAP7_75t_L g1904 ( 
.A(n_1826),
.Y(n_1904)
);

INVx3_ASAP7_75t_L g1905 ( 
.A(n_1832),
.Y(n_1905)
);

BUFx2_ASAP7_75t_L g1906 ( 
.A(n_1832),
.Y(n_1906)
);

BUFx2_ASAP7_75t_L g1907 ( 
.A(n_1832),
.Y(n_1907)
);

OAI21xp5_ASAP7_75t_SL g1908 ( 
.A1(n_1825),
.A2(n_1696),
.B(n_1722),
.Y(n_1908)
);

AND2x2_ASAP7_75t_L g1909 ( 
.A(n_1847),
.B(n_1853),
.Y(n_1909)
);

HB1xp67_ASAP7_75t_L g1910 ( 
.A(n_1870),
.Y(n_1910)
);

INVx1_ASAP7_75t_L g1911 ( 
.A(n_1870),
.Y(n_1911)
);

AND2x2_ASAP7_75t_L g1912 ( 
.A(n_1875),
.B(n_1825),
.Y(n_1912)
);

INVx2_ASAP7_75t_L g1913 ( 
.A(n_1883),
.Y(n_1913)
);

AND2x2_ASAP7_75t_L g1914 ( 
.A(n_1875),
.B(n_1830),
.Y(n_1914)
);

OAI211xp5_ASAP7_75t_SL g1915 ( 
.A1(n_1856),
.A2(n_1838),
.B(n_1844),
.C(n_1842),
.Y(n_1915)
);

AND2x4_ASAP7_75t_SL g1916 ( 
.A(n_1888),
.B(n_1864),
.Y(n_1916)
);

INVx1_ASAP7_75t_L g1917 ( 
.A(n_1883),
.Y(n_1917)
);

INVx3_ASAP7_75t_L g1918 ( 
.A(n_1875),
.Y(n_1918)
);

AND2x2_ASAP7_75t_L g1919 ( 
.A(n_1875),
.B(n_1830),
.Y(n_1919)
);

AND2x2_ASAP7_75t_L g1920 ( 
.A(n_1875),
.B(n_1906),
.Y(n_1920)
);

OA21x2_ASAP7_75t_L g1921 ( 
.A1(n_1906),
.A2(n_1835),
.B(n_1815),
.Y(n_1921)
);

INVx1_ASAP7_75t_L g1922 ( 
.A(n_1859),
.Y(n_1922)
);

NAND2xp5_ASAP7_75t_L g1923 ( 
.A(n_1860),
.B(n_1843),
.Y(n_1923)
);

INVx2_ASAP7_75t_L g1924 ( 
.A(n_1890),
.Y(n_1924)
);

NOR2xp33_ASAP7_75t_R g1925 ( 
.A(n_1901),
.B(n_1722),
.Y(n_1925)
);

INVx1_ASAP7_75t_L g1926 ( 
.A(n_1862),
.Y(n_1926)
);

INVx1_ASAP7_75t_L g1927 ( 
.A(n_1865),
.Y(n_1927)
);

AND2x2_ASAP7_75t_L g1928 ( 
.A(n_1907),
.B(n_1869),
.Y(n_1928)
);

INVx1_ASAP7_75t_L g1929 ( 
.A(n_1874),
.Y(n_1929)
);

AND2x2_ASAP7_75t_L g1930 ( 
.A(n_1907),
.B(n_1817),
.Y(n_1930)
);

NAND2xp5_ASAP7_75t_SL g1931 ( 
.A(n_1901),
.B(n_1818),
.Y(n_1931)
);

INVx3_ASAP7_75t_L g1932 ( 
.A(n_1869),
.Y(n_1932)
);

AND2x2_ASAP7_75t_L g1933 ( 
.A(n_1885),
.B(n_1818),
.Y(n_1933)
);

HB1xp67_ASAP7_75t_L g1934 ( 
.A(n_1873),
.Y(n_1934)
);

NAND2xp5_ASAP7_75t_L g1935 ( 
.A(n_1872),
.B(n_1846),
.Y(n_1935)
);

NAND2xp5_ASAP7_75t_SL g1936 ( 
.A(n_1861),
.B(n_1821),
.Y(n_1936)
);

AND2x2_ASAP7_75t_L g1937 ( 
.A(n_1885),
.B(n_1867),
.Y(n_1937)
);

AND2x2_ASAP7_75t_L g1938 ( 
.A(n_1867),
.B(n_1884),
.Y(n_1938)
);

AND2x4_ASAP7_75t_L g1939 ( 
.A(n_1905),
.B(n_1821),
.Y(n_1939)
);

NAND2xp5_ASAP7_75t_L g1940 ( 
.A(n_1872),
.B(n_1892),
.Y(n_1940)
);

NAND2xp5_ASAP7_75t_L g1941 ( 
.A(n_1892),
.B(n_1846),
.Y(n_1941)
);

NAND2x1_ASAP7_75t_L g1942 ( 
.A(n_1884),
.B(n_1821),
.Y(n_1942)
);

INVx2_ASAP7_75t_L g1943 ( 
.A(n_1890),
.Y(n_1943)
);

AND2x2_ASAP7_75t_L g1944 ( 
.A(n_1905),
.B(n_1909),
.Y(n_1944)
);

HB1xp67_ASAP7_75t_L g1945 ( 
.A(n_1904),
.Y(n_1945)
);

NAND2xp5_ASAP7_75t_L g1946 ( 
.A(n_1858),
.B(n_1850),
.Y(n_1946)
);

INVx3_ASAP7_75t_L g1947 ( 
.A(n_1905),
.Y(n_1947)
);

INVx1_ASAP7_75t_SL g1948 ( 
.A(n_1889),
.Y(n_1948)
);

OAI21xp5_ASAP7_75t_L g1949 ( 
.A1(n_1855),
.A2(n_1822),
.B(n_1842),
.Y(n_1949)
);

AND2x2_ASAP7_75t_L g1950 ( 
.A(n_1898),
.B(n_1909),
.Y(n_1950)
);

INVxp67_ASAP7_75t_L g1951 ( 
.A(n_1898),
.Y(n_1951)
);

NAND2xp5_ASAP7_75t_L g1952 ( 
.A(n_1951),
.B(n_1877),
.Y(n_1952)
);

AND2x2_ASAP7_75t_L g1953 ( 
.A(n_1916),
.B(n_1900),
.Y(n_1953)
);

NAND2x1_ASAP7_75t_L g1954 ( 
.A(n_1918),
.B(n_1888),
.Y(n_1954)
);

AND2x2_ASAP7_75t_L g1955 ( 
.A(n_1916),
.B(n_1900),
.Y(n_1955)
);

AOI22xp33_ASAP7_75t_L g1956 ( 
.A1(n_1936),
.A2(n_1857),
.B1(n_1882),
.B2(n_1866),
.Y(n_1956)
);

NAND2xp5_ASAP7_75t_L g1957 ( 
.A(n_1951),
.B(n_1878),
.Y(n_1957)
);

INVx1_ASAP7_75t_L g1958 ( 
.A(n_1945),
.Y(n_1958)
);

AND2x2_ASAP7_75t_L g1959 ( 
.A(n_1916),
.B(n_1900),
.Y(n_1959)
);

INVx1_ASAP7_75t_L g1960 ( 
.A(n_1945),
.Y(n_1960)
);

INVxp67_ASAP7_75t_L g1961 ( 
.A(n_1934),
.Y(n_1961)
);

NOR2xp67_ASAP7_75t_L g1962 ( 
.A(n_1918),
.B(n_1889),
.Y(n_1962)
);

INVx1_ASAP7_75t_L g1963 ( 
.A(n_1922),
.Y(n_1963)
);

INVx1_ASAP7_75t_L g1964 ( 
.A(n_1922),
.Y(n_1964)
);

INVx1_ASAP7_75t_L g1965 ( 
.A(n_1922),
.Y(n_1965)
);

INVx1_ASAP7_75t_SL g1966 ( 
.A(n_1948),
.Y(n_1966)
);

AND2x2_ASAP7_75t_L g1967 ( 
.A(n_1916),
.B(n_1868),
.Y(n_1967)
);

INVx1_ASAP7_75t_L g1968 ( 
.A(n_1926),
.Y(n_1968)
);

AND2x4_ASAP7_75t_L g1969 ( 
.A(n_1918),
.B(n_1864),
.Y(n_1969)
);

INVx2_ASAP7_75t_L g1970 ( 
.A(n_1921),
.Y(n_1970)
);

AND2x2_ASAP7_75t_L g1971 ( 
.A(n_1950),
.B(n_1868),
.Y(n_1971)
);

AND2x2_ASAP7_75t_L g1972 ( 
.A(n_1950),
.B(n_1868),
.Y(n_1972)
);

NAND2xp5_ASAP7_75t_L g1973 ( 
.A(n_1949),
.B(n_1871),
.Y(n_1973)
);

INVx2_ASAP7_75t_SL g1974 ( 
.A(n_1918),
.Y(n_1974)
);

BUFx2_ASAP7_75t_L g1975 ( 
.A(n_1925),
.Y(n_1975)
);

INVx2_ASAP7_75t_L g1976 ( 
.A(n_1921),
.Y(n_1976)
);

AND2x2_ASAP7_75t_L g1977 ( 
.A(n_1950),
.B(n_1888),
.Y(n_1977)
);

INVx2_ASAP7_75t_L g1978 ( 
.A(n_1921),
.Y(n_1978)
);

O2A1O1Ixp5_ASAP7_75t_SL g1979 ( 
.A1(n_1936),
.A2(n_1903),
.B(n_1815),
.C(n_1727),
.Y(n_1979)
);

INVx1_ASAP7_75t_L g1980 ( 
.A(n_1926),
.Y(n_1980)
);

OR2x2_ASAP7_75t_L g1981 ( 
.A(n_1940),
.B(n_1935),
.Y(n_1981)
);

AND2x2_ASAP7_75t_L g1982 ( 
.A(n_1933),
.B(n_1912),
.Y(n_1982)
);

INVx1_ASAP7_75t_L g1983 ( 
.A(n_1926),
.Y(n_1983)
);

OR2x2_ASAP7_75t_L g1984 ( 
.A(n_1940),
.B(n_1858),
.Y(n_1984)
);

INVxp67_ASAP7_75t_L g1985 ( 
.A(n_1934),
.Y(n_1985)
);

INVx1_ASAP7_75t_L g1986 ( 
.A(n_1927),
.Y(n_1986)
);

AND2x4_ASAP7_75t_L g1987 ( 
.A(n_1918),
.B(n_1864),
.Y(n_1987)
);

INVx2_ASAP7_75t_SL g1988 ( 
.A(n_1918),
.Y(n_1988)
);

HB1xp67_ASAP7_75t_L g1989 ( 
.A(n_1921),
.Y(n_1989)
);

INVx1_ASAP7_75t_L g1990 ( 
.A(n_1927),
.Y(n_1990)
);

INVx1_ASAP7_75t_L g1991 ( 
.A(n_1927),
.Y(n_1991)
);

OAI22xp33_ASAP7_75t_L g1992 ( 
.A1(n_1931),
.A2(n_1899),
.B1(n_1908),
.B2(n_1881),
.Y(n_1992)
);

NAND2xp5_ASAP7_75t_L g1993 ( 
.A(n_1949),
.B(n_1863),
.Y(n_1993)
);

NAND2xp5_ASAP7_75t_L g1994 ( 
.A(n_1941),
.B(n_1863),
.Y(n_1994)
);

OR2x2_ASAP7_75t_L g1995 ( 
.A(n_1935),
.B(n_1896),
.Y(n_1995)
);

INVx1_ASAP7_75t_L g1996 ( 
.A(n_1929),
.Y(n_1996)
);

AND2x2_ASAP7_75t_L g1997 ( 
.A(n_1933),
.B(n_1888),
.Y(n_1997)
);

AND2x2_ASAP7_75t_L g1998 ( 
.A(n_1933),
.B(n_1888),
.Y(n_1998)
);

XNOR2xp5_ASAP7_75t_L g1999 ( 
.A(n_1956),
.B(n_1931),
.Y(n_1999)
);

AND2x2_ASAP7_75t_L g2000 ( 
.A(n_1977),
.B(n_1948),
.Y(n_2000)
);

NAND2xp5_ASAP7_75t_L g2001 ( 
.A(n_1957),
.B(n_1924),
.Y(n_2001)
);

INVx1_ASAP7_75t_L g2002 ( 
.A(n_1963),
.Y(n_2002)
);

OR2x2_ASAP7_75t_L g2003 ( 
.A(n_1952),
.B(n_1924),
.Y(n_2003)
);

AND2x4_ASAP7_75t_L g2004 ( 
.A(n_1962),
.B(n_1920),
.Y(n_2004)
);

NAND2xp5_ASAP7_75t_L g2005 ( 
.A(n_1961),
.B(n_1924),
.Y(n_2005)
);

INVx1_ASAP7_75t_L g2006 ( 
.A(n_1963),
.Y(n_2006)
);

INVx1_ASAP7_75t_L g2007 ( 
.A(n_1964),
.Y(n_2007)
);

OR2x2_ASAP7_75t_L g2008 ( 
.A(n_1952),
.B(n_1981),
.Y(n_2008)
);

INVx1_ASAP7_75t_L g2009 ( 
.A(n_1964),
.Y(n_2009)
);

INVx1_ASAP7_75t_L g2010 ( 
.A(n_1965),
.Y(n_2010)
);

AND2x2_ASAP7_75t_L g2011 ( 
.A(n_1977),
.B(n_1920),
.Y(n_2011)
);

INVx2_ASAP7_75t_L g2012 ( 
.A(n_1970),
.Y(n_2012)
);

HB1xp67_ASAP7_75t_L g2013 ( 
.A(n_1966),
.Y(n_2013)
);

AND2x2_ASAP7_75t_L g2014 ( 
.A(n_1962),
.B(n_1920),
.Y(n_2014)
);

NOR2x1_ASAP7_75t_L g2015 ( 
.A(n_1975),
.B(n_1915),
.Y(n_2015)
);

OAI31xp33_ASAP7_75t_L g2016 ( 
.A1(n_1992),
.A2(n_1915),
.A3(n_1891),
.B(n_1879),
.Y(n_2016)
);

NAND2xp5_ASAP7_75t_L g2017 ( 
.A(n_1985),
.B(n_1966),
.Y(n_2017)
);

BUFx2_ASAP7_75t_L g2018 ( 
.A(n_1967),
.Y(n_2018)
);

NOR2xp33_ASAP7_75t_L g2019 ( 
.A(n_1973),
.B(n_1665),
.Y(n_2019)
);

AO21x1_ASAP7_75t_L g2020 ( 
.A1(n_1954),
.A2(n_1914),
.B(n_1912),
.Y(n_2020)
);

INVx3_ASAP7_75t_L g2021 ( 
.A(n_1954),
.Y(n_2021)
);

INVx1_ASAP7_75t_SL g2022 ( 
.A(n_1975),
.Y(n_2022)
);

NAND2xp5_ASAP7_75t_L g2023 ( 
.A(n_1958),
.B(n_1924),
.Y(n_2023)
);

AND2x2_ASAP7_75t_L g2024 ( 
.A(n_1971),
.B(n_1972),
.Y(n_2024)
);

NAND2xp5_ASAP7_75t_L g2025 ( 
.A(n_1958),
.B(n_1943),
.Y(n_2025)
);

INVx1_ASAP7_75t_L g2026 ( 
.A(n_1965),
.Y(n_2026)
);

AND2x2_ASAP7_75t_L g2027 ( 
.A(n_1971),
.B(n_1912),
.Y(n_2027)
);

AOI22xp33_ASAP7_75t_L g2028 ( 
.A1(n_1993),
.A2(n_1925),
.B1(n_1894),
.B2(n_1886),
.Y(n_2028)
);

INVx2_ASAP7_75t_L g2029 ( 
.A(n_1970),
.Y(n_2029)
);

INVx1_ASAP7_75t_L g2030 ( 
.A(n_1968),
.Y(n_2030)
);

INVx2_ASAP7_75t_L g2031 ( 
.A(n_1970),
.Y(n_2031)
);

INVx2_ASAP7_75t_L g2032 ( 
.A(n_1976),
.Y(n_2032)
);

AND2x2_ASAP7_75t_L g2033 ( 
.A(n_1972),
.B(n_1914),
.Y(n_2033)
);

AND2x2_ASAP7_75t_L g2034 ( 
.A(n_1982),
.B(n_1914),
.Y(n_2034)
);

INVx1_ASAP7_75t_L g2035 ( 
.A(n_1968),
.Y(n_2035)
);

OAI21xp33_ASAP7_75t_L g2036 ( 
.A1(n_1979),
.A2(n_1919),
.B(n_1943),
.Y(n_2036)
);

OR2x2_ASAP7_75t_L g2037 ( 
.A(n_1981),
.B(n_1943),
.Y(n_2037)
);

NAND2xp5_ASAP7_75t_L g2038 ( 
.A(n_2022),
.B(n_1982),
.Y(n_2038)
);

HB1xp67_ASAP7_75t_L g2039 ( 
.A(n_2013),
.Y(n_2039)
);

BUFx6f_ASAP7_75t_L g2040 ( 
.A(n_2021),
.Y(n_2040)
);

NAND2xp5_ASAP7_75t_L g2041 ( 
.A(n_2022),
.B(n_1997),
.Y(n_2041)
);

INVx1_ASAP7_75t_L g2042 ( 
.A(n_2013),
.Y(n_2042)
);

INVx1_ASAP7_75t_L g2043 ( 
.A(n_2002),
.Y(n_2043)
);

NAND2xp5_ASAP7_75t_L g2044 ( 
.A(n_1999),
.B(n_1997),
.Y(n_2044)
);

INVx2_ASAP7_75t_L g2045 ( 
.A(n_2021),
.Y(n_2045)
);

INVx1_ASAP7_75t_L g2046 ( 
.A(n_2002),
.Y(n_2046)
);

INVx1_ASAP7_75t_L g2047 ( 
.A(n_2006),
.Y(n_2047)
);

O2A1O1Ixp33_ASAP7_75t_SL g2048 ( 
.A1(n_1999),
.A2(n_1989),
.B(n_1974),
.C(n_1988),
.Y(n_2048)
);

OAI322xp33_ASAP7_75t_L g2049 ( 
.A1(n_2001),
.A2(n_1960),
.A3(n_1976),
.B1(n_1978),
.B2(n_1943),
.C1(n_1984),
.C2(n_1995),
.Y(n_2049)
);

INVx1_ASAP7_75t_L g2050 ( 
.A(n_2006),
.Y(n_2050)
);

INVx1_ASAP7_75t_L g2051 ( 
.A(n_2007),
.Y(n_2051)
);

INVx1_ASAP7_75t_L g2052 ( 
.A(n_2007),
.Y(n_2052)
);

OAI22xp5_ASAP7_75t_L g2053 ( 
.A1(n_2015),
.A2(n_1967),
.B1(n_1994),
.B2(n_1959),
.Y(n_2053)
);

NAND2xp5_ASAP7_75t_L g2054 ( 
.A(n_2015),
.B(n_2000),
.Y(n_2054)
);

NAND3xp33_ASAP7_75t_L g2055 ( 
.A(n_2016),
.B(n_1979),
.C(n_1960),
.Y(n_2055)
);

AOI332xp33_ASAP7_75t_L g2056 ( 
.A1(n_2001),
.A2(n_1978),
.A3(n_1976),
.B1(n_1980),
.B2(n_1991),
.B3(n_1990),
.C1(n_1983),
.C2(n_1996),
.Y(n_2056)
);

NAND2x1_ASAP7_75t_SL g2057 ( 
.A(n_2004),
.B(n_1953),
.Y(n_2057)
);

AOI222xp33_ASAP7_75t_L g2058 ( 
.A1(n_2017),
.A2(n_2036),
.B1(n_2028),
.B2(n_2016),
.C1(n_2000),
.C2(n_2018),
.Y(n_2058)
);

OAI221xp5_ASAP7_75t_L g2059 ( 
.A1(n_2017),
.A2(n_1942),
.B1(n_1984),
.B2(n_1974),
.C(n_1988),
.Y(n_2059)
);

INVxp33_ASAP7_75t_L g2060 ( 
.A(n_2019),
.Y(n_2060)
);

OAI21xp5_ASAP7_75t_L g2061 ( 
.A1(n_2036),
.A2(n_2004),
.B(n_2008),
.Y(n_2061)
);

XNOR2x1_ASAP7_75t_L g2062 ( 
.A(n_2008),
.B(n_1998),
.Y(n_2062)
);

NAND2xp5_ASAP7_75t_L g2063 ( 
.A(n_2018),
.B(n_1998),
.Y(n_2063)
);

INVx1_ASAP7_75t_L g2064 ( 
.A(n_2009),
.Y(n_2064)
);

AOI22xp5_ASAP7_75t_L g2065 ( 
.A1(n_2024),
.A2(n_1969),
.B1(n_1987),
.B2(n_1955),
.Y(n_2065)
);

AO22x1_ASAP7_75t_L g2066 ( 
.A1(n_2021),
.A2(n_1969),
.B1(n_1987),
.B2(n_1959),
.Y(n_2066)
);

OAI21xp5_ASAP7_75t_SL g2067 ( 
.A1(n_2058),
.A2(n_2011),
.B(n_2024),
.Y(n_2067)
);

AOI22xp33_ASAP7_75t_L g2068 ( 
.A1(n_2055),
.A2(n_2003),
.B1(n_2020),
.B2(n_2011),
.Y(n_2068)
);

OAI21xp5_ASAP7_75t_L g2069 ( 
.A1(n_2061),
.A2(n_2004),
.B(n_2003),
.Y(n_2069)
);

INVx1_ASAP7_75t_L g2070 ( 
.A(n_2039),
.Y(n_2070)
);

INVx2_ASAP7_75t_L g2071 ( 
.A(n_2040),
.Y(n_2071)
);

NAND2xp5_ASAP7_75t_L g2072 ( 
.A(n_2042),
.B(n_2024),
.Y(n_2072)
);

AOI222xp33_ASAP7_75t_L g2073 ( 
.A1(n_2054),
.A2(n_2005),
.B1(n_2014),
.B2(n_2004),
.C1(n_2034),
.C2(n_2033),
.Y(n_2073)
);

AOI31xp33_ASAP7_75t_L g2074 ( 
.A1(n_2060),
.A2(n_2044),
.A3(n_2039),
.B(n_2062),
.Y(n_2074)
);

OAI22xp5_ASAP7_75t_L g2075 ( 
.A1(n_2065),
.A2(n_2021),
.B1(n_2033),
.B2(n_2027),
.Y(n_2075)
);

OAI221xp5_ASAP7_75t_L g2076 ( 
.A1(n_2057),
.A2(n_2005),
.B1(n_2014),
.B2(n_2037),
.C(n_2023),
.Y(n_2076)
);

INVx2_ASAP7_75t_L g2077 ( 
.A(n_2040),
.Y(n_2077)
);

INVx2_ASAP7_75t_SL g2078 ( 
.A(n_2040),
.Y(n_2078)
);

AOI21xp33_ASAP7_75t_L g2079 ( 
.A1(n_2060),
.A2(n_2025),
.B(n_2023),
.Y(n_2079)
);

INVx1_ASAP7_75t_L g2080 ( 
.A(n_2043),
.Y(n_2080)
);

OAI21xp5_ASAP7_75t_L g2081 ( 
.A1(n_2048),
.A2(n_2014),
.B(n_2025),
.Y(n_2081)
);

OAI31xp33_ASAP7_75t_L g2082 ( 
.A1(n_2053),
.A2(n_2033),
.A3(n_2027),
.B(n_2034),
.Y(n_2082)
);

OR2x2_ASAP7_75t_L g2083 ( 
.A(n_2038),
.B(n_2037),
.Y(n_2083)
);

INVx1_ASAP7_75t_L g2084 ( 
.A(n_2046),
.Y(n_2084)
);

NAND2xp5_ASAP7_75t_L g2085 ( 
.A(n_2041),
.B(n_2034),
.Y(n_2085)
);

INVx1_ASAP7_75t_L g2086 ( 
.A(n_2047),
.Y(n_2086)
);

OAI22xp33_ASAP7_75t_L g2087 ( 
.A1(n_2059),
.A2(n_2063),
.B1(n_1942),
.B2(n_2040),
.Y(n_2087)
);

INVx1_ASAP7_75t_L g2088 ( 
.A(n_2050),
.Y(n_2088)
);

OAI222xp33_ASAP7_75t_L g2089 ( 
.A1(n_2056),
.A2(n_1969),
.B1(n_1987),
.B2(n_1942),
.C1(n_1978),
.C2(n_1919),
.Y(n_2089)
);

NAND2xp5_ASAP7_75t_L g2090 ( 
.A(n_2066),
.B(n_2020),
.Y(n_2090)
);

INVx1_ASAP7_75t_SL g2091 ( 
.A(n_2083),
.Y(n_2091)
);

INVx1_ASAP7_75t_L g2092 ( 
.A(n_2070),
.Y(n_2092)
);

AOI31xp33_ASAP7_75t_L g2093 ( 
.A1(n_2069),
.A2(n_2068),
.A3(n_2070),
.B(n_2090),
.Y(n_2093)
);

INVx1_ASAP7_75t_L g2094 ( 
.A(n_2072),
.Y(n_2094)
);

INVx2_ASAP7_75t_SL g2095 ( 
.A(n_2078),
.Y(n_2095)
);

INVx1_ASAP7_75t_L g2096 ( 
.A(n_2071),
.Y(n_2096)
);

AOI21xp33_ASAP7_75t_L g2097 ( 
.A1(n_2074),
.A2(n_2045),
.B(n_2051),
.Y(n_2097)
);

O2A1O1Ixp5_ASAP7_75t_L g2098 ( 
.A1(n_2089),
.A2(n_2049),
.B(n_2048),
.C(n_2064),
.Y(n_2098)
);

AND2x2_ASAP7_75t_L g2099 ( 
.A(n_2073),
.B(n_1953),
.Y(n_2099)
);

NOR2xp33_ASAP7_75t_L g2100 ( 
.A(n_2067),
.B(n_1665),
.Y(n_2100)
);

NAND2xp5_ASAP7_75t_SL g2101 ( 
.A(n_2087),
.B(n_1969),
.Y(n_2101)
);

INVx1_ASAP7_75t_L g2102 ( 
.A(n_2071),
.Y(n_2102)
);

HB1xp67_ASAP7_75t_L g2103 ( 
.A(n_2078),
.Y(n_2103)
);

INVx1_ASAP7_75t_L g2104 ( 
.A(n_2077),
.Y(n_2104)
);

NOR3xp33_ASAP7_75t_L g2105 ( 
.A(n_2093),
.B(n_2079),
.C(n_2077),
.Y(n_2105)
);

AND2x2_ASAP7_75t_L g2106 ( 
.A(n_2099),
.B(n_2085),
.Y(n_2106)
);

AOI21xp33_ASAP7_75t_SL g2107 ( 
.A1(n_2097),
.A2(n_2100),
.B(n_2082),
.Y(n_2107)
);

OAI32xp33_ASAP7_75t_L g2108 ( 
.A1(n_2091),
.A2(n_2068),
.A3(n_2081),
.B1(n_2076),
.B2(n_2075),
.Y(n_2108)
);

AND2x2_ASAP7_75t_L g2109 ( 
.A(n_2099),
.B(n_2083),
.Y(n_2109)
);

NAND2xp5_ASAP7_75t_L g2110 ( 
.A(n_2103),
.B(n_2080),
.Y(n_2110)
);

INVx1_ASAP7_75t_L g2111 ( 
.A(n_2092),
.Y(n_2111)
);

INVx1_ASAP7_75t_L g2112 ( 
.A(n_2092),
.Y(n_2112)
);

OAI21xp5_ASAP7_75t_L g2113 ( 
.A1(n_2098),
.A2(n_2086),
.B(n_2084),
.Y(n_2113)
);

NAND2xp5_ASAP7_75t_L g2114 ( 
.A(n_2095),
.B(n_2088),
.Y(n_2114)
);

OAI21xp33_ASAP7_75t_SL g2115 ( 
.A1(n_2101),
.A2(n_2052),
.B(n_2010),
.Y(n_2115)
);

OAI211xp5_ASAP7_75t_L g2116 ( 
.A1(n_2094),
.A2(n_2035),
.B(n_2009),
.C(n_2010),
.Y(n_2116)
);

AOI322xp5_ASAP7_75t_L g2117 ( 
.A1(n_2094),
.A2(n_2035),
.A3(n_2026),
.B1(n_2030),
.B2(n_2031),
.C1(n_2029),
.C2(n_2032),
.Y(n_2117)
);

OR2x2_ASAP7_75t_L g2118 ( 
.A(n_2095),
.B(n_2096),
.Y(n_2118)
);

O2A1O1Ixp33_ASAP7_75t_L g2119 ( 
.A1(n_2108),
.A2(n_2104),
.B(n_2102),
.C(n_2026),
.Y(n_2119)
);

NAND2xp5_ASAP7_75t_L g2120 ( 
.A(n_2109),
.B(n_2104),
.Y(n_2120)
);

OAI211xp5_ASAP7_75t_L g2121 ( 
.A1(n_2113),
.A2(n_2102),
.B(n_2030),
.C(n_2031),
.Y(n_2121)
);

INVx1_ASAP7_75t_L g2122 ( 
.A(n_2118),
.Y(n_2122)
);

AOI221xp5_ASAP7_75t_L g2123 ( 
.A1(n_2107),
.A2(n_2032),
.B1(n_2031),
.B2(n_2029),
.C(n_2012),
.Y(n_2123)
);

INVx1_ASAP7_75t_L g2124 ( 
.A(n_2114),
.Y(n_2124)
);

NAND4xp25_ASAP7_75t_L g2125 ( 
.A(n_2105),
.B(n_1895),
.C(n_2029),
.D(n_2012),
.Y(n_2125)
);

AOI221xp5_ASAP7_75t_L g2126 ( 
.A1(n_2115),
.A2(n_2106),
.B1(n_2110),
.B2(n_2112),
.C(n_2111),
.Y(n_2126)
);

AOI211xp5_ASAP7_75t_L g2127 ( 
.A1(n_2116),
.A2(n_1987),
.B(n_2012),
.C(n_2032),
.Y(n_2127)
);

AOI221xp5_ASAP7_75t_L g2128 ( 
.A1(n_2119),
.A2(n_2117),
.B1(n_1919),
.B2(n_1983),
.C(n_1991),
.Y(n_2128)
);

OAI221xp5_ASAP7_75t_SL g2129 ( 
.A1(n_2126),
.A2(n_2117),
.B1(n_1955),
.B2(n_1995),
.C(n_1887),
.Y(n_2129)
);

AOI22xp5_ASAP7_75t_L g2130 ( 
.A1(n_2122),
.A2(n_1996),
.B1(n_1990),
.B2(n_1986),
.Y(n_2130)
);

NOR3x1_ASAP7_75t_L g2131 ( 
.A(n_2120),
.B(n_1986),
.C(n_1980),
.Y(n_2131)
);

AOI211xp5_ASAP7_75t_L g2132 ( 
.A1(n_2125),
.A2(n_1880),
.B(n_1902),
.C(n_1928),
.Y(n_2132)
);

OAI22xp5_ASAP7_75t_L g2133 ( 
.A1(n_2124),
.A2(n_1921),
.B1(n_1947),
.B2(n_1932),
.Y(n_2133)
);

AOI222xp33_ASAP7_75t_L g2134 ( 
.A1(n_2121),
.A2(n_1930),
.B1(n_1938),
.B2(n_1937),
.C1(n_1928),
.C2(n_1910),
.Y(n_2134)
);

OAI211xp5_ASAP7_75t_L g2135 ( 
.A1(n_2123),
.A2(n_1921),
.B(n_1947),
.C(n_1932),
.Y(n_2135)
);

INVxp67_ASAP7_75t_L g2136 ( 
.A(n_2130),
.Y(n_2136)
);

NAND4xp75_ASAP7_75t_L g2137 ( 
.A(n_2131),
.B(n_2127),
.C(n_1928),
.D(n_1938),
.Y(n_2137)
);

AND2x2_ASAP7_75t_L g2138 ( 
.A(n_2132),
.B(n_1938),
.Y(n_2138)
);

AO22x1_ASAP7_75t_L g2139 ( 
.A1(n_2129),
.A2(n_1928),
.B1(n_1947),
.B2(n_1932),
.Y(n_2139)
);

NAND2xp5_ASAP7_75t_L g2140 ( 
.A(n_2128),
.B(n_1937),
.Y(n_2140)
);

NOR2xp33_ASAP7_75t_L g2141 ( 
.A(n_2135),
.B(n_1876),
.Y(n_2141)
);

OAI221xp5_ASAP7_75t_L g2142 ( 
.A1(n_2136),
.A2(n_2133),
.B1(n_2134),
.B2(n_1947),
.C(n_1932),
.Y(n_2142)
);

NAND3x1_ASAP7_75t_SL g2143 ( 
.A(n_2138),
.B(n_1748),
.C(n_1937),
.Y(n_2143)
);

NOR2x1p5_ASAP7_75t_L g2144 ( 
.A(n_2137),
.B(n_1876),
.Y(n_2144)
);

OAI221xp5_ASAP7_75t_SL g2145 ( 
.A1(n_2140),
.A2(n_1887),
.B1(n_1947),
.B2(n_1932),
.C(n_1893),
.Y(n_2145)
);

NAND2xp5_ASAP7_75t_L g2146 ( 
.A(n_2144),
.B(n_2139),
.Y(n_2146)
);

OAI21xp33_ASAP7_75t_L g2147 ( 
.A1(n_2145),
.A2(n_2141),
.B(n_1893),
.Y(n_2147)
);

AO22x2_ASAP7_75t_L g2148 ( 
.A1(n_2146),
.A2(n_2143),
.B1(n_2142),
.B2(n_1947),
.Y(n_2148)
);

OAI21x1_ASAP7_75t_L g2149 ( 
.A1(n_2148),
.A2(n_2147),
.B(n_1932),
.Y(n_2149)
);

OAI22xp5_ASAP7_75t_L g2150 ( 
.A1(n_2148),
.A2(n_1941),
.B1(n_1923),
.B2(n_1910),
.Y(n_2150)
);

AOI21xp33_ASAP7_75t_L g2151 ( 
.A1(n_2149),
.A2(n_1923),
.B(n_1913),
.Y(n_2151)
);

OAI22xp5_ASAP7_75t_L g2152 ( 
.A1(n_2150),
.A2(n_1946),
.B1(n_1913),
.B2(n_1944),
.Y(n_2152)
);

AOI22x1_ASAP7_75t_L g2153 ( 
.A1(n_2151),
.A2(n_1702),
.B1(n_1913),
.B2(n_1716),
.Y(n_2153)
);

INVx1_ASAP7_75t_L g2154 ( 
.A(n_2152),
.Y(n_2154)
);

XOR2xp5_ASAP7_75t_L g2155 ( 
.A(n_2154),
.B(n_1692),
.Y(n_2155)
);

AOI21xp33_ASAP7_75t_SL g2156 ( 
.A1(n_2155),
.A2(n_2153),
.B(n_1713),
.Y(n_2156)
);

INVx1_ASAP7_75t_L g2157 ( 
.A(n_2156),
.Y(n_2157)
);

OAI221xp5_ASAP7_75t_R g2158 ( 
.A1(n_2157),
.A2(n_1748),
.B1(n_1913),
.B2(n_1939),
.C(n_1897),
.Y(n_2158)
);

AOI211xp5_ASAP7_75t_L g2159 ( 
.A1(n_2158),
.A2(n_1692),
.B(n_1911),
.C(n_1917),
.Y(n_2159)
);


endmodule