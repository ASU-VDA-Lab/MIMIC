module fake_jpeg_28414_n_225 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_225);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_225;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_1),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

INVx1_ASAP7_75t_SL g20 ( 
.A(n_4),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_5),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_0),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_12),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_1),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_16),
.Y(n_32)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_4),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_18),
.Y(n_36)
);

OR2x2_ASAP7_75t_SL g73 ( 
.A(n_36),
.B(n_40),
.Y(n_73)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_27),
.Y(n_37)
);

BUFx4f_ASAP7_75t_SL g79 ( 
.A(n_37),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g38 ( 
.A(n_20),
.Y(n_38)
);

INVx4_ASAP7_75t_SL g55 ( 
.A(n_38),
.Y(n_55)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_18),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_28),
.B(n_16),
.Y(n_41)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_41),
.B(n_32),
.Y(n_70)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_27),
.Y(n_42)
);

CKINVDCx9p33_ASAP7_75t_R g69 ( 
.A(n_42),
.Y(n_69)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_27),
.Y(n_43)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_43),
.Y(n_64)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_31),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_44),
.B(n_48),
.Y(n_80)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_27),
.Y(n_45)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_45),
.Y(n_62)
);

INVx13_ASAP7_75t_L g46 ( 
.A(n_30),
.Y(n_46)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_46),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_30),
.Y(n_47)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_47),
.Y(n_68)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_31),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_21),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_49),
.Y(n_61)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_30),
.Y(n_50)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_50),
.Y(n_77)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_30),
.Y(n_51)
);

INVx6_ASAP7_75t_L g78 ( 
.A(n_51),
.Y(n_78)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_17),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_52),
.Y(n_54)
);

CKINVDCx12_ASAP7_75t_R g53 ( 
.A(n_37),
.Y(n_53)
);

INVxp67_ASAP7_75t_L g83 ( 
.A(n_53),
.Y(n_83)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_47),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_56),
.B(n_59),
.Y(n_89)
);

AOI21xp5_ASAP7_75t_L g58 ( 
.A1(n_38),
.A2(n_20),
.B(n_2),
.Y(n_58)
);

AOI21xp5_ASAP7_75t_L g86 ( 
.A1(n_58),
.A2(n_1),
.B(n_3),
.Y(n_86)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_47),
.Y(n_59)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_39),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_60),
.B(n_66),
.Y(n_101)
);

AO22x1_ASAP7_75t_SL g63 ( 
.A1(n_52),
.A2(n_17),
.B1(n_34),
.B2(n_24),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_63),
.A2(n_44),
.B1(n_48),
.B2(n_19),
.Y(n_85)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_43),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_36),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_67),
.B(n_75),
.Y(n_102)
);

OR2x2_ASAP7_75t_L g109 ( 
.A(n_70),
.B(n_23),
.Y(n_109)
);

OAI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_50),
.A2(n_33),
.B1(n_29),
.B2(n_26),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_71),
.A2(n_72),
.B1(n_25),
.B2(n_23),
.Y(n_100)
);

OAI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_51),
.A2(n_33),
.B1(n_29),
.B2(n_26),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_L g74 ( 
.A1(n_46),
.A2(n_17),
.B1(n_34),
.B2(n_24),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_74),
.A2(n_35),
.B1(n_19),
.B2(n_42),
.Y(n_90)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_40),
.Y(n_75)
);

INVx2_ASAP7_75t_SL g76 ( 
.A(n_46),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_76),
.B(n_55),
.Y(n_105)
);

NAND4xp25_ASAP7_75t_L g81 ( 
.A(n_61),
.B(n_49),
.C(n_32),
.D(n_28),
.Y(n_81)
);

NOR2x1_ASAP7_75t_L g116 ( 
.A(n_81),
.B(n_73),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_80),
.B(n_21),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_82),
.B(n_88),
.Y(n_111)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_77),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_84),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_85),
.A2(n_90),
.B1(n_68),
.B2(n_62),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_86),
.A2(n_100),
.B1(n_104),
.B2(n_88),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_63),
.B(n_45),
.C(n_43),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g128 ( 
.A(n_87),
.B(n_99),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_71),
.B(n_35),
.Y(n_88)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_54),
.Y(n_91)
);

INVx1_ASAP7_75t_SL g131 ( 
.A(n_91),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_72),
.B(n_34),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_92),
.B(n_98),
.Y(n_113)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_57),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_93),
.B(n_105),
.Y(n_118)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_54),
.Y(n_94)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_94),
.Y(n_117)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_62),
.Y(n_95)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_95),
.Y(n_132)
);

BUFx12_ASAP7_75t_L g96 ( 
.A(n_69),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_96),
.Y(n_114)
);

BUFx2_ASAP7_75t_L g97 ( 
.A(n_76),
.Y(n_97)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_97),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_70),
.B(n_24),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_57),
.B(n_45),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_65),
.B(n_45),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_103),
.B(n_79),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_55),
.A2(n_25),
.B1(n_23),
.B2(n_22),
.Y(n_104)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_74),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_106),
.B(n_109),
.Y(n_133)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_78),
.Y(n_107)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_107),
.Y(n_125)
);

BUFx8_ASAP7_75t_L g108 ( 
.A(n_79),
.Y(n_108)
);

INVx5_ASAP7_75t_L g112 ( 
.A(n_108),
.Y(n_112)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_78),
.Y(n_110)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_110),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_115),
.A2(n_94),
.B1(n_84),
.B2(n_83),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_116),
.B(n_120),
.Y(n_139)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_95),
.Y(n_120)
);

NOR2x1_ASAP7_75t_L g121 ( 
.A(n_100),
.B(n_65),
.Y(n_121)
);

OR2x2_ASAP7_75t_L g138 ( 
.A(n_121),
.B(n_124),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_122),
.B(n_123),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_82),
.B(n_43),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_102),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_129),
.B(n_109),
.Y(n_134)
);

A2O1A1Ixp33_ASAP7_75t_SL g130 ( 
.A1(n_87),
.A2(n_68),
.B(n_64),
.C(n_22),
.Y(n_130)
);

OAI22x1_ASAP7_75t_L g148 ( 
.A1(n_130),
.A2(n_99),
.B1(n_91),
.B2(n_107),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_134),
.B(n_141),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_115),
.A2(n_92),
.B1(n_85),
.B2(n_104),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_135),
.A2(n_149),
.B1(n_131),
.B2(n_132),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_111),
.B(n_103),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_137),
.B(n_142),
.Y(n_159)
);

XOR2xp5_ASAP7_75t_L g140 ( 
.A(n_113),
.B(n_98),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g157 ( 
.A(n_140),
.B(n_150),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_123),
.B(n_101),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_122),
.Y(n_142)
);

NAND3xp33_ASAP7_75t_L g143 ( 
.A(n_116),
.B(n_111),
.C(n_113),
.Y(n_143)
);

NOR2x1_ASAP7_75t_L g160 ( 
.A(n_143),
.B(n_12),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_126),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_144),
.B(n_145),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_126),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_121),
.A2(n_128),
.B1(n_133),
.B2(n_130),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_146),
.A2(n_125),
.B1(n_131),
.B2(n_117),
.Y(n_158)
);

A2O1A1Ixp33_ASAP7_75t_L g147 ( 
.A1(n_128),
.A2(n_86),
.B(n_99),
.C(n_89),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_L g168 ( 
.A1(n_147),
.A2(n_114),
.B(n_5),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_SL g167 ( 
.A1(n_148),
.A2(n_119),
.B(n_114),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_128),
.B(n_108),
.C(n_83),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_118),
.B(n_22),
.Y(n_151)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_151),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_L g152 ( 
.A(n_130),
.B(n_108),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_152),
.B(n_155),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_127),
.B(n_3),
.Y(n_153)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_153),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_130),
.B(n_97),
.C(n_96),
.Y(n_154)
);

INVxp67_ASAP7_75t_L g163 ( 
.A(n_154),
.Y(n_163)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_125),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g156 ( 
.A(n_137),
.B(n_127),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_SL g176 ( 
.A(n_156),
.B(n_136),
.Y(n_176)
);

AOI221xp5_ASAP7_75t_L g175 ( 
.A1(n_158),
.A2(n_160),
.B1(n_139),
.B2(n_151),
.C(n_153),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_164),
.B(n_138),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_148),
.A2(n_120),
.B1(n_119),
.B2(n_112),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_165),
.B(n_145),
.Y(n_183)
);

XNOR2x2_ASAP7_75t_SL g166 ( 
.A(n_136),
.B(n_3),
.Y(n_166)
);

A2O1A1Ixp33_ASAP7_75t_L g179 ( 
.A1(n_166),
.A2(n_138),
.B(n_154),
.C(n_142),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_L g181 ( 
.A1(n_167),
.A2(n_168),
.B(n_172),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_L g172 ( 
.A1(n_147),
.A2(n_4),
.B(n_5),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_135),
.A2(n_112),
.B1(n_7),
.B2(n_8),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_173),
.Y(n_174)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_175),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_176),
.B(n_177),
.Y(n_196)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_161),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_159),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_178),
.B(n_183),
.Y(n_194)
);

AOI21xp5_ASAP7_75t_L g192 ( 
.A1(n_179),
.A2(n_185),
.B(n_187),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_180),
.A2(n_165),
.B1(n_162),
.B2(n_166),
.Y(n_197)
);

AOI221xp5_ASAP7_75t_L g182 ( 
.A1(n_168),
.A2(n_146),
.B1(n_152),
.B2(n_140),
.C(n_150),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_182),
.B(n_157),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_156),
.B(n_155),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_SL g198 ( 
.A(n_184),
.B(n_171),
.Y(n_198)
);

AOI21xp5_ASAP7_75t_L g185 ( 
.A1(n_167),
.A2(n_144),
.B(n_8),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_157),
.B(n_96),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_186),
.B(n_164),
.Y(n_190)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_159),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_188),
.B(n_190),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_186),
.B(n_170),
.C(n_163),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_189),
.B(n_191),
.C(n_195),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_178),
.B(n_163),
.C(n_169),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_187),
.B(n_169),
.C(n_162),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_197),
.B(n_198),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_188),
.B(n_177),
.C(n_179),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_200),
.B(n_203),
.C(n_13),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g202 ( 
.A(n_190),
.B(n_181),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_202),
.B(n_189),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_193),
.B(n_181),
.C(n_172),
.Y(n_203)
);

OAI22xp33_ASAP7_75t_SL g205 ( 
.A1(n_192),
.A2(n_183),
.B1(n_185),
.B2(n_174),
.Y(n_205)
);

AOI21xp5_ASAP7_75t_L g209 ( 
.A1(n_205),
.A2(n_191),
.B(n_195),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_194),
.A2(n_174),
.B1(n_173),
.B2(n_160),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_206),
.B(n_196),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_207),
.B(n_208),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_209),
.A2(n_210),
.B1(n_201),
.B2(n_9),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_199),
.B(n_14),
.C(n_8),
.Y(n_211)
);

INVxp67_ASAP7_75t_L g213 ( 
.A(n_211),
.Y(n_213)
);

AND2x2_ASAP7_75t_L g212 ( 
.A(n_202),
.B(n_6),
.Y(n_212)
);

AOI322xp5_ASAP7_75t_L g217 ( 
.A1(n_212),
.A2(n_6),
.A3(n_9),
.B1(n_10),
.B2(n_11),
.C1(n_172),
.C2(n_139),
.Y(n_217)
);

AOI221xp5_ASAP7_75t_L g214 ( 
.A1(n_212),
.A2(n_204),
.B1(n_205),
.B2(n_201),
.C(n_14),
.Y(n_214)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_214),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_215),
.B(n_217),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_SL g218 ( 
.A(n_216),
.B(n_207),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_218),
.B(n_213),
.Y(n_222)
);

AOI21xp5_ASAP7_75t_SL g221 ( 
.A1(n_220),
.A2(n_213),
.B(n_9),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_221),
.B(n_222),
.Y(n_223)
);

NOR2xp67_ASAP7_75t_L g224 ( 
.A(n_223),
.B(n_219),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_224),
.B(n_6),
.Y(n_225)
);


endmodule