module fake_jpeg_19704_n_118 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_118);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_118;

wire n_117;
wire n_10;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_112;
wire n_95;
wire n_97;
wire n_9;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g9 ( 
.A(n_1),
.Y(n_9)
);

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_2),
.Y(n_10)
);

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_8),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_2),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_2),
.Y(n_13)
);

INVx6_ASAP7_75t_L g14 ( 
.A(n_3),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_7),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_6),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

INVx3_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_18),
.B(n_19),
.Y(n_32)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_15),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_20),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_21),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

INVx1_ASAP7_75t_SL g31 ( 
.A(n_22),
.Y(n_31)
);

BUFx2_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_23),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_12),
.Y(n_24)
);

AOI22xp33_ASAP7_75t_L g27 ( 
.A1(n_24),
.A2(n_9),
.B1(n_16),
.B2(n_13),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_SL g26 ( 
.A1(n_18),
.A2(n_14),
.B1(n_17),
.B2(n_12),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_SL g38 ( 
.A1(n_26),
.A2(n_29),
.B1(n_31),
.B2(n_24),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_27),
.B(n_11),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_L g29 ( 
.A1(n_18),
.A2(n_14),
.B1(n_17),
.B2(n_12),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_32),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_33),
.B(n_34),
.Y(n_49)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_30),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_25),
.Y(n_35)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_35),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_32),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_36),
.B(n_39),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_25),
.Y(n_37)
);

INVxp67_ASAP7_75t_L g45 ( 
.A(n_37),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_L g42 ( 
.A1(n_38),
.A2(n_41),
.B1(n_31),
.B2(n_30),
.Y(n_42)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_26),
.Y(n_39)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_40),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_42),
.B(n_23),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g44 ( 
.A1(n_33),
.A2(n_31),
.B1(n_14),
.B2(n_17),
.Y(n_44)
);

CKINVDCx14_ASAP7_75t_R g60 ( 
.A(n_44),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_39),
.A2(n_28),
.B1(n_19),
.B2(n_26),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_46),
.B(n_47),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g47 ( 
.A1(n_36),
.A2(n_38),
.B1(n_41),
.B2(n_28),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_34),
.A2(n_28),
.B1(n_19),
.B2(n_29),
.Y(n_50)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_50),
.Y(n_55)
);

AOI21xp5_ASAP7_75t_L g52 ( 
.A1(n_51),
.A2(n_0),
.B(n_40),
.Y(n_52)
);

OAI21xp5_ASAP7_75t_SL g66 ( 
.A1(n_52),
.A2(n_53),
.B(n_45),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g54 ( 
.A(n_51),
.B(n_21),
.C(n_20),
.Y(n_54)
);

XNOR2xp5_ASAP7_75t_L g70 ( 
.A(n_54),
.B(n_50),
.Y(n_70)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_49),
.Y(n_57)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_57),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_49),
.B(n_27),
.Y(n_58)
);

OAI21xp33_ASAP7_75t_L g64 ( 
.A1(n_58),
.A2(n_44),
.B(n_42),
.Y(n_64)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_48),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_59),
.B(n_48),
.Y(n_69)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_46),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_61),
.Y(n_63)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_64),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_57),
.B(n_47),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_65),
.B(n_68),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_66),
.B(n_70),
.Y(n_74)
);

NOR3xp33_ASAP7_75t_L g67 ( 
.A(n_52),
.B(n_16),
.C(n_13),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_67),
.B(n_16),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g68 ( 
.A(n_54),
.Y(n_68)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_69),
.Y(n_78)
);

AOI21xp5_ASAP7_75t_L g71 ( 
.A1(n_60),
.A2(n_0),
.B(n_13),
.Y(n_71)
);

AOI21x1_ASAP7_75t_L g76 ( 
.A1(n_71),
.A2(n_56),
.B(n_0),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g72 ( 
.A(n_62),
.B(n_58),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_72),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_L g85 ( 
.A1(n_76),
.A2(n_55),
.B(n_11),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_70),
.B(n_56),
.C(n_61),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_77),
.B(n_80),
.C(n_15),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_79),
.A2(n_11),
.B1(n_10),
.B2(n_9),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_65),
.B(n_55),
.C(n_59),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_68),
.B(n_63),
.Y(n_81)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_81),
.Y(n_89)
);

AOI322xp5_ASAP7_75t_SL g83 ( 
.A1(n_76),
.A2(n_78),
.A3(n_71),
.B1(n_74),
.B2(n_75),
.C1(n_77),
.C2(n_66),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_83),
.B(n_84),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_85),
.A2(n_10),
.B1(n_0),
.B2(n_3),
.Y(n_97)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_80),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_86),
.B(n_88),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_87),
.B(n_37),
.C(n_35),
.Y(n_92)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_73),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_80),
.A2(n_43),
.B1(n_37),
.B2(n_35),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_90),
.A2(n_43),
.B1(n_25),
.B2(n_22),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_82),
.A2(n_43),
.B1(n_10),
.B2(n_9),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_91),
.B(n_95),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_92),
.B(n_96),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_90),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_97),
.B(n_85),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_98),
.B(n_99),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_94),
.B(n_87),
.C(n_86),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g102 ( 
.A(n_92),
.B(n_89),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_102),
.B(n_100),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_93),
.B(n_88),
.C(n_96),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_103),
.B(n_23),
.Y(n_107)
);

OAI21xp33_ASAP7_75t_L g105 ( 
.A1(n_101),
.A2(n_95),
.B(n_3),
.Y(n_105)
);

XOR2xp5_ASAP7_75t_L g110 ( 
.A(n_105),
.B(n_1),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_106),
.A2(n_107),
.B1(n_1),
.B2(n_4),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_101),
.A2(n_25),
.B1(n_22),
.B2(n_20),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_108),
.A2(n_21),
.B1(n_5),
.B2(n_7),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_109),
.B(n_110),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_104),
.A2(n_23),
.B1(n_21),
.B2(n_6),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_111),
.B(n_112),
.C(n_110),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_113),
.B(n_111),
.Y(n_115)
);

O2A1O1Ixp33_ASAP7_75t_SL g117 ( 
.A1(n_115),
.A2(n_116),
.B(n_4),
.C(n_5),
.Y(n_117)
);

NOR3xp33_ASAP7_75t_L g116 ( 
.A(n_114),
.B(n_4),
.C(n_5),
.Y(n_116)
);

XOR2xp5_ASAP7_75t_L g118 ( 
.A(n_117),
.B(n_7),
.Y(n_118)
);


endmodule