module fake_netlist_1_691_n_24 (n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_24);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_24;
wire n_20;
wire n_23;
wire n_22;
wire n_11;
wire n_16;
wire n_13;
wire n_18;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_19;
wire n_21;
NAND2xp33_ASAP7_75t_R g11 ( .A(n_5), .B(n_6), .Y(n_11) );
CKINVDCx5p33_ASAP7_75t_R g12 ( .A(n_10), .Y(n_12) );
AND2x2_ASAP7_75t_L g13 ( .A(n_9), .B(n_2), .Y(n_13) );
BUFx2_ASAP7_75t_L g14 ( .A(n_4), .Y(n_14) );
CKINVDCx5p33_ASAP7_75t_R g15 ( .A(n_3), .Y(n_15) );
INVx1_ASAP7_75t_L g16 ( .A(n_14), .Y(n_16) );
BUFx4f_ASAP7_75t_L g17 ( .A(n_13), .Y(n_17) );
INVxp67_ASAP7_75t_L g18 ( .A(n_16), .Y(n_18) );
AND2x4_ASAP7_75t_L g19 ( .A(n_18), .B(n_15), .Y(n_19) );
AOI22xp5_ASAP7_75t_L g20 ( .A1(n_19), .A2(n_17), .B1(n_12), .B2(n_11), .Y(n_20) );
INVx1_ASAP7_75t_SL g21 ( .A(n_20), .Y(n_21) );
AND2x2_ASAP7_75t_L g22 ( .A(n_21), .B(n_0), .Y(n_22) );
CKINVDCx20_ASAP7_75t_R g23 ( .A(n_22), .Y(n_23) );
AOI22xp5_ASAP7_75t_SL g24 ( .A1(n_23), .A2(n_1), .B1(n_7), .B2(n_8), .Y(n_24) );
endmodule