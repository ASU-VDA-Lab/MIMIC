module fake_jpeg_12133_n_192 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_51, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_192);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_51;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_192;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_76;
wire n_127;
wire n_154;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_143;
wire n_122;
wire n_75;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_91;
wire n_93;
wire n_54;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

INVx4_ASAP7_75t_L g52 ( 
.A(n_9),
.Y(n_52)
);

CKINVDCx16_ASAP7_75t_R g53 ( 
.A(n_37),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_24),
.Y(n_54)
);

BUFx5_ASAP7_75t_L g55 ( 
.A(n_28),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_3),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_10),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_4),
.Y(n_58)
);

INVx1_ASAP7_75t_SL g59 ( 
.A(n_4),
.Y(n_59)
);

INVx1_ASAP7_75t_SL g60 ( 
.A(n_13),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_51),
.Y(n_61)
);

BUFx8_ASAP7_75t_L g62 ( 
.A(n_12),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_48),
.Y(n_63)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_2),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_43),
.Y(n_65)
);

BUFx5_ASAP7_75t_L g66 ( 
.A(n_17),
.Y(n_66)
);

INVxp67_ASAP7_75t_L g67 ( 
.A(n_21),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_50),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_14),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_23),
.Y(n_70)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_25),
.Y(n_71)
);

BUFx5_ASAP7_75t_L g72 ( 
.A(n_49),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_15),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_1),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_42),
.Y(n_75)
);

BUFx12_ASAP7_75t_L g76 ( 
.A(n_6),
.Y(n_76)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_3),
.Y(n_77)
);

BUFx12_ASAP7_75t_L g78 ( 
.A(n_31),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_47),
.Y(n_79)
);

INVx2_ASAP7_75t_SL g80 ( 
.A(n_34),
.Y(n_80)
);

AND2x2_ASAP7_75t_SL g81 ( 
.A(n_62),
.B(n_29),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_81),
.B(n_83),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_74),
.B(n_0),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_82),
.B(n_84),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_78),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_78),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_76),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_85),
.B(n_86),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_59),
.B(n_0),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_56),
.Y(n_87)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_87),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_63),
.Y(n_88)
);

INVx6_ASAP7_75t_L g91 ( 
.A(n_88),
.Y(n_91)
);

INVx8_ASAP7_75t_L g89 ( 
.A(n_55),
.Y(n_89)
);

INVx5_ASAP7_75t_L g93 ( 
.A(n_89),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_76),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_90),
.B(n_60),
.Y(n_105)
);

INVx5_ASAP7_75t_L g94 ( 
.A(n_89),
.Y(n_94)
);

BUFx2_ASAP7_75t_L g121 ( 
.A(n_94),
.Y(n_121)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_88),
.Y(n_95)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_95),
.Y(n_110)
);

BUFx5_ASAP7_75t_L g96 ( 
.A(n_81),
.Y(n_96)
);

BUFx12f_ASAP7_75t_L g107 ( 
.A(n_96),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_81),
.A2(n_57),
.B1(n_52),
.B2(n_77),
.Y(n_98)
);

AOI21xp5_ASAP7_75t_L g123 ( 
.A1(n_98),
.A2(n_101),
.B(n_80),
.Y(n_123)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_87),
.Y(n_100)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_100),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_89),
.A2(n_57),
.B1(n_64),
.B2(n_71),
.Y(n_101)
);

INVx11_ASAP7_75t_L g102 ( 
.A(n_89),
.Y(n_102)
);

INVx8_ASAP7_75t_L g113 ( 
.A(n_102),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_88),
.A2(n_69),
.B1(n_65),
.B2(n_73),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_103),
.A2(n_68),
.B1(n_58),
.B2(n_53),
.Y(n_126)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_87),
.Y(n_104)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_104),
.Y(n_116)
);

AND2x2_ASAP7_75t_L g120 ( 
.A(n_105),
.B(n_62),
.Y(n_120)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_99),
.Y(n_108)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_108),
.Y(n_133)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_91),
.Y(n_109)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_109),
.Y(n_136)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_91),
.Y(n_111)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_111),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_96),
.B(n_56),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g147 ( 
.A(n_112),
.B(n_7),
.Y(n_147)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_93),
.Y(n_114)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_114),
.Y(n_135)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_93),
.Y(n_117)
);

BUFx3_ASAP7_75t_L g137 ( 
.A(n_117),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_102),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_118),
.B(n_119),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_97),
.B(n_79),
.Y(n_119)
);

AND2x2_ASAP7_75t_L g130 ( 
.A(n_120),
.B(n_123),
.Y(n_130)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_94),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_122),
.Y(n_132)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_92),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_124),
.B(n_120),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_106),
.B(n_79),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_125),
.B(n_5),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_126),
.A2(n_127),
.B1(n_67),
.B2(n_72),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_98),
.A2(n_58),
.B1(n_61),
.B2(n_54),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_112),
.B(n_54),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_131),
.B(n_134),
.Y(n_151)
);

NOR2x1_ASAP7_75t_L g138 ( 
.A(n_107),
.B(n_61),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_138),
.B(n_141),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_107),
.A2(n_101),
.B1(n_75),
.B2(n_70),
.Y(n_139)
);

OAI22x1_ASAP7_75t_SL g165 ( 
.A1(n_139),
.A2(n_39),
.B1(n_40),
.B2(n_41),
.Y(n_165)
);

AND2x2_ASAP7_75t_L g140 ( 
.A(n_115),
.B(n_1),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g150 ( 
.A(n_140),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_116),
.B(n_2),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_142),
.A2(n_148),
.B1(n_11),
.B2(n_16),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_143),
.B(n_144),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_121),
.B(n_5),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_118),
.B(n_6),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_145),
.B(n_146),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_110),
.Y(n_146)
);

OR2x2_ASAP7_75t_L g156 ( 
.A(n_147),
.B(n_22),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_113),
.A2(n_66),
.B1(n_8),
.B2(n_9),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g149 ( 
.A(n_124),
.B(n_7),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_149),
.B(n_38),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_SL g152 ( 
.A(n_130),
.B(n_35),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_152),
.B(n_46),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_130),
.A2(n_8),
.B1(n_10),
.B2(n_11),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_153),
.A2(n_155),
.B1(n_159),
.B2(n_165),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_154),
.A2(n_160),
.B1(n_44),
.B2(n_45),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_SL g155 ( 
.A1(n_137),
.A2(n_18),
.B1(n_19),
.B2(n_20),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_156),
.B(n_157),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_129),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_140),
.A2(n_26),
.B1(n_27),
.B2(n_30),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_139),
.A2(n_32),
.B1(n_33),
.B2(n_36),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_161),
.B(n_166),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_138),
.B(n_133),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_163),
.B(n_167),
.Y(n_173)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_136),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_132),
.B(n_128),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_164),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_168),
.Y(n_180)
);

AOI22x1_ASAP7_75t_L g169 ( 
.A1(n_150),
.A2(n_135),
.B1(n_132),
.B2(n_137),
.Y(n_169)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_169),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_150),
.A2(n_158),
.B1(n_151),
.B2(n_155),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g181 ( 
.A(n_170),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_172),
.B(n_174),
.Y(n_178)
);

CKINVDCx16_ASAP7_75t_R g175 ( 
.A(n_162),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_L g182 ( 
.A1(n_175),
.A2(n_156),
.B(n_152),
.Y(n_182)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_182),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_178),
.B(n_176),
.C(n_174),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_183),
.B(n_177),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_185),
.B(n_180),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_186),
.B(n_173),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_187),
.B(n_184),
.Y(n_188)
);

MAJx2_ASAP7_75t_L g189 ( 
.A(n_188),
.B(n_170),
.C(n_171),
.Y(n_189)
);

MAJx2_ASAP7_75t_L g190 ( 
.A(n_189),
.B(n_179),
.C(n_181),
.Y(n_190)
);

BUFx24_ASAP7_75t_SL g191 ( 
.A(n_190),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_191),
.B(n_181),
.Y(n_192)
);


endmodule