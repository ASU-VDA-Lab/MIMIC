module real_jpeg_16972_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_425;
wire n_455;
wire n_50;
wire n_409;
wire n_186;
wire n_137;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_366;
wire n_456;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_432;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_411;
wire n_382;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_450;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_404;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_343;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_447;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

INVx1_ASAP7_75t_SL g82 ( 
.A(n_0),
.Y(n_82)
);

AOI21xp5_ASAP7_75t_L g18 ( 
.A1(n_1),
.A2(n_19),
.B(n_460),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g460 ( 
.A(n_1),
.B(n_461),
.Y(n_460)
);

AND2x2_ASAP7_75t_L g39 ( 
.A(n_2),
.B(n_40),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_2),
.B(n_84),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_2),
.B(n_36),
.Y(n_110)
);

AND2x2_ASAP7_75t_L g119 ( 
.A(n_2),
.B(n_120),
.Y(n_119)
);

AND2x2_ASAP7_75t_L g135 ( 
.A(n_2),
.B(n_124),
.Y(n_135)
);

AND2x2_ASAP7_75t_L g145 ( 
.A(n_2),
.B(n_146),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_2),
.B(n_302),
.Y(n_301)
);

AND2x2_ASAP7_75t_L g446 ( 
.A(n_2),
.B(n_447),
.Y(n_446)
);

AND2x2_ASAP7_75t_L g35 ( 
.A(n_3),
.B(n_36),
.Y(n_35)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_3),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_3),
.B(n_96),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g166 ( 
.A(n_3),
.B(n_167),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g306 ( 
.A(n_3),
.B(n_307),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_4),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_4),
.B(n_69),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_4),
.B(n_132),
.Y(n_131)
);

AND2x2_ASAP7_75t_L g147 ( 
.A(n_4),
.B(n_106),
.Y(n_147)
);

AND2x2_ASAP7_75t_SL g193 ( 
.A(n_4),
.B(n_194),
.Y(n_193)
);

AND2x2_ASAP7_75t_SL g338 ( 
.A(n_4),
.B(n_339),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_SL g343 ( 
.A(n_4),
.B(n_344),
.Y(n_343)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_5),
.B(n_59),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_5),
.B(n_73),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_5),
.B(n_128),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_5),
.B(n_163),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_5),
.B(n_45),
.Y(n_186)
);

CKINVDCx16_ASAP7_75t_R g297 ( 
.A(n_5),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_SL g431 ( 
.A(n_5),
.B(n_132),
.Y(n_431)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_6),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_6),
.Y(n_125)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_6),
.Y(n_192)
);

BUFx3_ASAP7_75t_L g265 ( 
.A(n_6),
.Y(n_265)
);

BUFx5_ASAP7_75t_L g75 ( 
.A(n_7),
.Y(n_75)
);

BUFx5_ASAP7_75t_L g84 ( 
.A(n_7),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_7),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g200 ( 
.A(n_7),
.Y(n_200)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_8),
.B(n_78),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_8),
.B(n_231),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_8),
.B(n_258),
.Y(n_257)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_8),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_8),
.B(n_383),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_SL g387 ( 
.A(n_8),
.B(n_388),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_SL g391 ( 
.A(n_8),
.B(n_392),
.Y(n_391)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_9),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_9),
.Y(n_47)
);

INVx2_ASAP7_75t_L g373 ( 
.A(n_9),
.Y(n_373)
);

AND2x2_ASAP7_75t_SL g49 ( 
.A(n_10),
.B(n_50),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_10),
.B(n_105),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_10),
.B(n_116),
.Y(n_115)
);

AND2x2_ASAP7_75t_SL g188 ( 
.A(n_10),
.B(n_189),
.Y(n_188)
);

AND2x2_ASAP7_75t_SL g261 ( 
.A(n_10),
.B(n_262),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_SL g331 ( 
.A(n_10),
.B(n_84),
.Y(n_331)
);

AND2x2_ASAP7_75t_SL g333 ( 
.A(n_10),
.B(n_334),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_10),
.B(n_371),
.Y(n_370)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_11),
.Y(n_81)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_11),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_11),
.Y(n_129)
);

BUFx3_ASAP7_75t_L g169 ( 
.A(n_11),
.Y(n_169)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_11),
.Y(n_197)
);

BUFx5_ASAP7_75t_L g263 ( 
.A(n_11),
.Y(n_263)
);

BUFx3_ASAP7_75t_L g324 ( 
.A(n_11),
.Y(n_324)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_12),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_12),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_12),
.Y(n_134)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_13),
.Y(n_461)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_14),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_14),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g30 ( 
.A(n_15),
.B(n_31),
.Y(n_30)
);

AND2x2_ASAP7_75t_L g55 ( 
.A(n_15),
.B(n_56),
.Y(n_55)
);

AND2x2_ASAP7_75t_SL g224 ( 
.A(n_15),
.B(n_225),
.Y(n_224)
);

AND2x2_ASAP7_75t_L g264 ( 
.A(n_15),
.B(n_265),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g320 ( 
.A(n_15),
.B(n_321),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_15),
.B(n_367),
.Y(n_366)
);

AND2x2_ASAP7_75t_SL g378 ( 
.A(n_15),
.B(n_379),
.Y(n_378)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_16),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g346 ( 
.A(n_16),
.Y(n_346)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_17),
.Y(n_33)
);

BUFx8_ASAP7_75t_L g447 ( 
.A(n_17),
.Y(n_447)
);

XOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_423),
.Y(n_19)
);

HB1xp67_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_310),
.Y(n_21)
);

A2O1A1O1Ixp25_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_211),
.B(n_267),
.C(n_268),
.D(n_309),
.Y(n_22)
);

INVx2_ASAP7_75t_SL g23 ( 
.A(n_24),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_24),
.B(n_269),
.Y(n_311)
);

AND2x2_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_174),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_25),
.B(n_174),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_100),
.Y(n_25)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_26),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_67),
.C(n_85),
.Y(n_26)
);

INVxp67_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_28),
.B(n_177),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_41),
.C(n_54),
.Y(n_28)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_29),
.B(n_233),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_34),
.Y(n_29)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_30),
.B(n_35),
.C(n_39),
.Y(n_87)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx5_ASAP7_75t_L g78 ( 
.A(n_32),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g287 ( 
.A(n_32),
.Y(n_287)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_33),
.Y(n_107)
);

XNOR2xp5_ASAP7_75t_L g34 ( 
.A(n_35),
.B(n_39),
.Y(n_34)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g337 ( 
.A(n_38),
.Y(n_337)
);

XNOR2xp5_ASAP7_75t_L g351 ( 
.A(n_39),
.B(n_154),
.Y(n_351)
);

AND2x2_ASAP7_75t_L g111 ( 
.A(n_40),
.B(n_90),
.Y(n_111)
);

INVx3_ASAP7_75t_L g340 ( 
.A(n_40),
.Y(n_340)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_41),
.A2(n_42),
.B1(n_54),
.B2(n_234),
.Y(n_233)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

AOI21xp5_ASAP7_75t_L g221 ( 
.A1(n_42),
.A2(n_43),
.B(n_49),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_43),
.B(n_49),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_SL g43 ( 
.A(n_44),
.B(n_48),
.Y(n_43)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx5_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g450 ( 
.A(n_48),
.B(n_451),
.Y(n_450)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_52),
.Y(n_146)
);

INVx3_ASAP7_75t_L g296 ( 
.A(n_52),
.Y(n_296)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_53),
.Y(n_71)
);

BUFx5_ASAP7_75t_L g260 ( 
.A(n_53),
.Y(n_260)
);

BUFx6f_ASAP7_75t_L g452 ( 
.A(n_53),
.Y(n_452)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_54),
.Y(n_234)
);

MAJx2_ASAP7_75t_L g54 ( 
.A(n_55),
.B(n_58),
.C(n_62),
.Y(n_54)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_55),
.B(n_58),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_56),
.B(n_90),
.Y(n_152)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx4_ASAP7_75t_L g304 ( 
.A(n_57),
.Y(n_304)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

AND2x2_ASAP7_75t_L g154 ( 
.A(n_61),
.B(n_90),
.Y(n_154)
);

BUFx3_ASAP7_75t_L g369 ( 
.A(n_61),
.Y(n_369)
);

XNOR2xp5_ASAP7_75t_SL g181 ( 
.A(n_62),
.B(n_182),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_63),
.B(n_64),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g352 ( 
.A(n_63),
.B(n_353),
.Y(n_352)
);

HB1xp67_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_67),
.A2(n_85),
.B1(n_86),
.B2(n_178),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_67),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g67 ( 
.A(n_68),
.B(n_72),
.C(n_76),
.Y(n_67)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_68),
.B(n_72),
.Y(n_202)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx2_ASAP7_75t_SL g353 ( 
.A(n_75),
.Y(n_353)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_76),
.B(n_202),
.Y(n_201)
);

MAJx2_ASAP7_75t_L g76 ( 
.A(n_77),
.B(n_79),
.C(n_83),
.Y(n_76)
);

XNOR2xp5_ASAP7_75t_SL g217 ( 
.A(n_77),
.B(n_218),
.Y(n_217)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_79),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g432 ( 
.A1(n_79),
.A2(n_198),
.B1(n_220),
.B2(n_253),
.Y(n_432)
);

OR2x2_ASAP7_75t_L g79 ( 
.A(n_80),
.B(n_82),
.Y(n_79)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx3_ASAP7_75t_L g384 ( 
.A(n_81),
.Y(n_384)
);

INVx1_ASAP7_75t_SL g90 ( 
.A(n_82),
.Y(n_90)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_83),
.B(n_161),
.Y(n_160)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_83),
.Y(n_219)
);

INVx1_ASAP7_75t_SL g85 ( 
.A(n_86),
.Y(n_85)
);

XNOR2xp5_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_88),
.Y(n_86)
);

MAJx2_ASAP7_75t_L g140 ( 
.A(n_87),
.B(n_89),
.C(n_95),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_89),
.A2(n_94),
.B1(n_95),
.B2(n_99),
.Y(n_88)
);

INVx1_ASAP7_75t_SL g99 ( 
.A(n_89),
.Y(n_99)
);

NAND2x1_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_91),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g123 ( 
.A(n_90),
.B(n_124),
.Y(n_123)
);

AND2x2_ASAP7_75t_L g198 ( 
.A(n_90),
.B(n_199),
.Y(n_198)
);

AND2x2_ASAP7_75t_L g285 ( 
.A(n_90),
.B(n_286),
.Y(n_285)
);

INVx6_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_93),
.Y(n_228)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx6_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_101),
.A2(n_150),
.B1(n_172),
.B2(n_173),
.Y(n_100)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_101),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_138),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_102),
.B(n_139),
.C(n_276),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_113),
.C(n_126),
.Y(n_102)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_103),
.B(n_113),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_108),
.Y(n_103)
);

OAI21xp33_ASAP7_75t_L g158 ( 
.A1(n_104),
.A2(n_110),
.B(n_111),
.Y(n_158)
);

BUFx2_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_109),
.A2(n_110),
.B1(n_111),
.B2(n_112),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_109),
.A2(n_110),
.B1(n_185),
.B2(n_186),
.Y(n_254)
);

INVx1_ASAP7_75t_SL g109 ( 
.A(n_110),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_110),
.B(n_111),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_110),
.B(n_185),
.Y(n_184)
);

INVx1_ASAP7_75t_SL g112 ( 
.A(n_111),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_111),
.A2(n_112),
.B1(n_154),
.B2(n_155),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_111),
.B(n_152),
.C(n_155),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g342 ( 
.A(n_111),
.B(n_343),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_112),
.B(n_343),
.Y(n_349)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_119),
.C(n_123),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_114),
.A2(n_115),
.B1(n_123),
.B2(n_206),
.Y(n_205)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

HB1xp67_ASAP7_75t_L g231 ( 
.A(n_118),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_119),
.A2(n_204),
.B1(n_205),
.B2(n_207),
.Y(n_203)
);

INVx1_ASAP7_75t_SL g207 ( 
.A(n_119),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_119),
.A2(n_207),
.B1(n_306),
.B2(n_308),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g435 ( 
.A(n_119),
.B(n_308),
.C(n_436),
.Y(n_435)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx1_ASAP7_75t_SL g206 ( 
.A(n_123),
.Y(n_206)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_125),
.Y(n_165)
);

XOR2x1_ASAP7_75t_L g209 ( 
.A(n_126),
.B(n_210),
.Y(n_209)
);

XNOR2x1_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_130),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_127),
.B(n_131),
.C(n_137),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_131),
.A2(n_135),
.B1(n_136),
.B2(n_137),
.Y(n_130)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_131),
.Y(n_136)
);

INVx4_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx4_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_135),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_L g449 ( 
.A(n_137),
.B(n_450),
.Y(n_449)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_139),
.A2(n_140),
.B1(n_141),
.B2(n_149),
.Y(n_138)
);

INVx1_ASAP7_75t_SL g139 ( 
.A(n_140),
.Y(n_139)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_141),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_143),
.Y(n_141)
);

MAJx2_ASAP7_75t_L g281 ( 
.A(n_142),
.B(n_144),
.C(n_148),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_144),
.A2(n_145),
.B1(n_147),
.B2(n_148),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_144),
.A2(n_145),
.B1(n_285),
.B2(n_288),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g441 ( 
.A(n_144),
.B(n_285),
.C(n_442),
.Y(n_441)
);

INVx3_ASAP7_75t_SL g144 ( 
.A(n_145),
.Y(n_144)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_147),
.Y(n_148)
);

HB1xp67_ASAP7_75t_L g276 ( 
.A(n_149),
.Y(n_276)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_150),
.Y(n_173)
);

HB1xp67_ASAP7_75t_L g273 ( 
.A(n_150),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_156),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_151),
.B(n_157),
.C(n_160),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_153),
.Y(n_151)
);

INVx1_ASAP7_75t_SL g155 ( 
.A(n_154),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_L g291 ( 
.A1(n_154),
.A2(n_155),
.B1(n_198),
.B2(n_253),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_SL g434 ( 
.A(n_155),
.B(n_198),
.C(n_292),
.Y(n_434)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_160),
.Y(n_156)
);

AND2x2_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_159),
.Y(n_157)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_159),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g408 ( 
.A1(n_159),
.A2(n_223),
.B1(n_409),
.B2(n_410),
.Y(n_408)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_162),
.A2(n_166),
.B1(n_170),
.B2(n_171),
.Y(n_161)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_162),
.Y(n_171)
);

INVx5_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

INVx5_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_166),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_166),
.B(n_171),
.C(n_219),
.Y(n_299)
);

INVx3_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

INVx5_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

HB1xp67_ASAP7_75t_L g271 ( 
.A(n_172),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_179),
.C(n_208),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g236 ( 
.A1(n_175),
.A2(n_176),
.B1(n_209),
.B2(n_237),
.Y(n_236)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_179),
.B(n_236),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_201),
.C(n_203),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_180),
.B(n_215),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_183),
.C(n_187),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_SL g246 ( 
.A(n_181),
.B(n_247),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_183),
.A2(n_184),
.B1(n_187),
.B2(n_248),
.Y(n_247)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_187),
.Y(n_248)
);

MAJx2_ASAP7_75t_L g187 ( 
.A(n_188),
.B(n_193),
.C(n_198),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_188),
.A2(n_198),
.B1(n_252),
.B2(n_253),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_188),
.Y(n_252)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

BUFx6f_ASAP7_75t_L g307 ( 
.A(n_191),
.Y(n_307)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_SL g250 ( 
.A(n_193),
.B(n_251),
.Y(n_250)
);

INVx3_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

INVx1_ASAP7_75t_SL g253 ( 
.A(n_198),
.Y(n_253)
);

BUFx6f_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVx6_ASAP7_75t_L g380 ( 
.A(n_200),
.Y(n_380)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_201),
.B(n_203),
.Y(n_215)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

HB1xp67_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_209),
.Y(n_237)
);

AOI21x1_ASAP7_75t_L g211 ( 
.A1(n_212),
.A2(n_238),
.B(n_266),
.Y(n_211)
);

OR2x2_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_235),
.Y(n_212)
);

AND2x2_ASAP7_75t_L g266 ( 
.A(n_213),
.B(n_235),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_216),
.C(n_232),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_214),
.B(n_240),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_216),
.B(n_232),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_221),
.C(n_222),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_217),
.B(n_221),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_220),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_222),
.B(n_244),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_224),
.C(n_229),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g410 ( 
.A1(n_224),
.A2(n_229),
.B1(n_230),
.B2(n_411),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_224),
.Y(n_411)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

INVx2_ASAP7_75t_SL g227 ( 
.A(n_228),
.Y(n_227)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_239),
.B(n_241),
.Y(n_238)
);

OR2x2_ASAP7_75t_L g312 ( 
.A(n_239),
.B(n_241),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_245),
.C(n_249),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g419 ( 
.A1(n_242),
.A2(n_243),
.B1(n_420),
.B2(n_421),
.Y(n_419)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g421 ( 
.A(n_246),
.B(n_249),
.Y(n_421)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_254),
.C(n_255),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g413 ( 
.A(n_250),
.B(n_414),
.Y(n_413)
);

XNOR2xp5_ASAP7_75t_L g414 ( 
.A(n_254),
.B(n_255),
.Y(n_414)
);

MAJx2_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_261),
.C(n_264),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g360 ( 
.A1(n_256),
.A2(n_257),
.B1(n_264),
.B2(n_361),
.Y(n_360)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

INVx2_ASAP7_75t_SL g259 ( 
.A(n_260),
.Y(n_259)
);

XNOR2x1_ASAP7_75t_L g359 ( 
.A(n_261),
.B(n_360),
.Y(n_359)
);

BUFx6f_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

CKINVDCx16_ASAP7_75t_R g361 ( 
.A(n_264),
.Y(n_361)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_265),
.Y(n_330)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_266),
.Y(n_313)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

AND2x2_ASAP7_75t_L g269 ( 
.A(n_270),
.B(n_274),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_270),
.B(n_274),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_271),
.B(n_272),
.C(n_273),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_275),
.B(n_277),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_R g456 ( 
.A(n_275),
.B(n_278),
.C(n_457),
.Y(n_456)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_278),
.B(n_289),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_279),
.B(n_280),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g454 ( 
.A(n_279),
.B(n_281),
.C(n_455),
.Y(n_454)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_281),
.B(n_282),
.Y(n_280)
);

HB1xp67_ASAP7_75t_L g455 ( 
.A(n_282),
.Y(n_455)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_283),
.B(n_284),
.Y(n_282)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_283),
.Y(n_442)
);

INVx1_ASAP7_75t_SL g288 ( 
.A(n_285),
.Y(n_288)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

HB1xp67_ASAP7_75t_L g457 ( 
.A(n_289),
.Y(n_457)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_290),
.B(n_298),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g453 ( 
.A(n_290),
.B(n_299),
.C(n_300),
.Y(n_453)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_291),
.B(n_292),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_293),
.B(n_297),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

BUFx3_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_299),
.B(n_300),
.Y(n_298)
);

XNOR2x1_ASAP7_75t_SL g300 ( 
.A(n_301),
.B(n_305),
.Y(n_300)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_301),
.Y(n_436)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

INVx6_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_306),
.Y(n_308)
);

NAND4xp25_ASAP7_75t_L g310 ( 
.A(n_311),
.B(n_312),
.C(n_313),
.D(n_314),
.Y(n_310)
);

OAI21xp5_ASAP7_75t_L g314 ( 
.A1(n_315),
.A2(n_417),
.B(n_422),
.Y(n_314)
);

AOI21x1_ASAP7_75t_SL g315 ( 
.A1(n_316),
.A2(n_405),
.B(n_416),
.Y(n_315)
);

OAI21x1_ASAP7_75t_L g316 ( 
.A1(n_317),
.A2(n_362),
.B(n_404),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_318),
.B(n_347),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_318),
.B(n_347),
.Y(n_404)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_319),
.B(n_332),
.C(n_341),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_L g400 ( 
.A(n_319),
.B(n_401),
.Y(n_400)
);

XOR2xp5_ASAP7_75t_L g319 ( 
.A(n_320),
.B(n_325),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g357 ( 
.A(n_320),
.B(n_331),
.C(n_358),
.Y(n_357)
);

INVx1_ASAP7_75t_SL g321 ( 
.A(n_322),
.Y(n_321)
);

BUFx2_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

INVx3_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_L g325 ( 
.A(n_326),
.B(n_331),
.Y(n_325)
);

INVxp67_ASAP7_75t_L g358 ( 
.A(n_326),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_327),
.B(n_328),
.Y(n_326)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_L g401 ( 
.A1(n_332),
.A2(n_341),
.B1(n_342),
.B2(n_402),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_332),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_333),
.B(n_338),
.Y(n_332)
);

XOR2xp5_ASAP7_75t_L g375 ( 
.A(n_333),
.B(n_338),
.Y(n_375)
);

INVx2_ASAP7_75t_L g334 ( 
.A(n_335),
.Y(n_334)
);

INVx2_ASAP7_75t_L g335 ( 
.A(n_336),
.Y(n_335)
);

INVx2_ASAP7_75t_L g336 ( 
.A(n_337),
.Y(n_336)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_340),
.Y(n_339)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_342),
.Y(n_341)
);

BUFx3_ASAP7_75t_L g344 ( 
.A(n_345),
.Y(n_344)
);

BUFx3_ASAP7_75t_L g345 ( 
.A(n_346),
.Y(n_345)
);

XNOR2xp5_ASAP7_75t_L g347 ( 
.A(n_348),
.B(n_356),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g415 ( 
.A(n_348),
.B(n_357),
.C(n_359),
.Y(n_415)
);

XNOR2xp5_ASAP7_75t_L g348 ( 
.A(n_349),
.B(n_350),
.Y(n_348)
);

MAJIxp5_ASAP7_75t_L g412 ( 
.A(n_349),
.B(n_352),
.C(n_354),
.Y(n_412)
);

AOI22xp5_ASAP7_75t_SL g350 ( 
.A1(n_351),
.A2(n_352),
.B1(n_354),
.B2(n_355),
.Y(n_350)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_351),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_352),
.Y(n_355)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_353),
.Y(n_388)
);

XNOR2xp5_ASAP7_75t_L g356 ( 
.A(n_357),
.B(n_359),
.Y(n_356)
);

AOI21xp5_ASAP7_75t_L g362 ( 
.A1(n_363),
.A2(n_398),
.B(n_403),
.Y(n_362)
);

OAI21xp5_ASAP7_75t_SL g363 ( 
.A1(n_364),
.A2(n_385),
.B(n_397),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_L g364 ( 
.A(n_365),
.B(n_374),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_SL g397 ( 
.A(n_365),
.B(n_374),
.Y(n_397)
);

NOR2xp33_ASAP7_75t_L g365 ( 
.A(n_366),
.B(n_370),
.Y(n_365)
);

XNOR2xp5_ASAP7_75t_L g389 ( 
.A(n_366),
.B(n_370),
.Y(n_389)
);

NOR2xp33_ASAP7_75t_L g390 ( 
.A(n_366),
.B(n_391),
.Y(n_390)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_368),
.Y(n_367)
);

INVx3_ASAP7_75t_L g368 ( 
.A(n_369),
.Y(n_368)
);

BUFx6f_ASAP7_75t_L g371 ( 
.A(n_372),
.Y(n_371)
);

INVx3_ASAP7_75t_L g372 ( 
.A(n_373),
.Y(n_372)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_373),
.Y(n_395)
);

XOR2xp5_ASAP7_75t_L g374 ( 
.A(n_375),
.B(n_376),
.Y(n_374)
);

MAJIxp5_ASAP7_75t_L g399 ( 
.A(n_375),
.B(n_378),
.C(n_381),
.Y(n_399)
);

OAI22xp5_ASAP7_75t_SL g376 ( 
.A1(n_377),
.A2(n_378),
.B1(n_381),
.B2(n_382),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_378),
.Y(n_377)
);

INVx4_ASAP7_75t_L g379 ( 
.A(n_380),
.Y(n_379)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_382),
.Y(n_381)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_384),
.Y(n_383)
);

AOI21xp5_ASAP7_75t_L g385 ( 
.A1(n_386),
.A2(n_390),
.B(n_396),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_387),
.B(n_389),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_L g396 ( 
.A(n_387),
.B(n_389),
.Y(n_396)
);

BUFx3_ASAP7_75t_L g392 ( 
.A(n_393),
.Y(n_392)
);

BUFx6f_ASAP7_75t_L g393 ( 
.A(n_394),
.Y(n_393)
);

BUFx6f_ASAP7_75t_L g394 ( 
.A(n_395),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_399),
.B(n_400),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_L g403 ( 
.A(n_399),
.B(n_400),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_SL g405 ( 
.A(n_406),
.B(n_415),
.Y(n_405)
);

NOR2xp67_ASAP7_75t_L g416 ( 
.A(n_406),
.B(n_415),
.Y(n_416)
);

XNOR2xp5_ASAP7_75t_L g406 ( 
.A(n_407),
.B(n_413),
.Y(n_406)
);

XNOR2xp5_ASAP7_75t_L g407 ( 
.A(n_408),
.B(n_412),
.Y(n_407)
);

MAJIxp5_ASAP7_75t_L g418 ( 
.A(n_408),
.B(n_412),
.C(n_413),
.Y(n_418)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_410),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_L g417 ( 
.A(n_418),
.B(n_419),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_418),
.B(n_419),
.Y(n_422)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_421),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_L g423 ( 
.A(n_424),
.B(n_458),
.Y(n_423)
);

INVxp33_ASAP7_75t_L g424 ( 
.A(n_425),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_SL g425 ( 
.A(n_426),
.B(n_456),
.Y(n_425)
);

OR2x2_ASAP7_75t_L g459 ( 
.A(n_426),
.B(n_456),
.Y(n_459)
);

XOR2xp5_ASAP7_75t_L g426 ( 
.A(n_427),
.B(n_454),
.Y(n_426)
);

AOI22xp5_ASAP7_75t_L g427 ( 
.A1(n_428),
.A2(n_429),
.B1(n_437),
.B2(n_438),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_429),
.Y(n_428)
);

XNOR2xp5_ASAP7_75t_L g429 ( 
.A(n_430),
.B(n_433),
.Y(n_429)
);

XNOR2xp5_ASAP7_75t_SL g430 ( 
.A(n_431),
.B(n_432),
.Y(n_430)
);

XNOR2xp5_ASAP7_75t_L g433 ( 
.A(n_434),
.B(n_435),
.Y(n_433)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_438),
.Y(n_437)
);

XOR2xp5_ASAP7_75t_L g438 ( 
.A(n_439),
.B(n_453),
.Y(n_438)
);

OAI22xp5_ASAP7_75t_SL g439 ( 
.A1(n_440),
.A2(n_441),
.B1(n_443),
.B2(n_444),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_441),
.Y(n_440)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_444),
.Y(n_443)
);

AOI22xp5_ASAP7_75t_L g444 ( 
.A1(n_445),
.A2(n_446),
.B1(n_448),
.B2(n_449),
.Y(n_444)
);

CKINVDCx20_ASAP7_75t_R g445 ( 
.A(n_446),
.Y(n_445)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_449),
.Y(n_448)
);

INVx2_ASAP7_75t_L g451 ( 
.A(n_452),
.Y(n_451)
);

INVxp33_ASAP7_75t_L g458 ( 
.A(n_459),
.Y(n_458)
);


endmodule