module fake_jpeg_28677_n_415 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_415);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_415;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_4),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_12),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_4),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_1),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

CKINVDCx16_ASAP7_75t_R g28 ( 
.A(n_9),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_10),
.Y(n_35)
);

BUFx8_ASAP7_75t_L g36 ( 
.A(n_11),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

INVx13_ASAP7_75t_L g38 ( 
.A(n_7),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_1),
.Y(n_39)
);

BUFx12_ASAP7_75t_L g40 ( 
.A(n_7),
.Y(n_40)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_3),
.Y(n_41)
);

INVx11_ASAP7_75t_L g42 ( 
.A(n_4),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_9),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_3),
.Y(n_44)
);

INVx13_ASAP7_75t_L g45 ( 
.A(n_41),
.Y(n_45)
);

INVx13_ASAP7_75t_L g90 ( 
.A(n_45),
.Y(n_90)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_24),
.Y(n_46)
);

INVx5_ASAP7_75t_L g96 ( 
.A(n_46),
.Y(n_96)
);

INVxp67_ASAP7_75t_SL g47 ( 
.A(n_36),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_47),
.B(n_50),
.Y(n_91)
);

BUFx5_ASAP7_75t_L g48 ( 
.A(n_25),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g92 ( 
.A(n_48),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_15),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_49),
.Y(n_89)
);

INVx2_ASAP7_75t_SL g50 ( 
.A(n_41),
.Y(n_50)
);

BUFx5_ASAP7_75t_L g51 ( 
.A(n_25),
.Y(n_51)
);

INVx5_ASAP7_75t_L g119 ( 
.A(n_51),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_15),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_52),
.Y(n_93)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_53),
.B(n_77),
.Y(n_104)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_54),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_15),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_55),
.Y(n_99)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_24),
.Y(n_56)
);

INVx4_ASAP7_75t_L g128 ( 
.A(n_56),
.Y(n_128)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

INVx4_ASAP7_75t_L g129 ( 
.A(n_57),
.Y(n_129)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_24),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_58),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_16),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_59),
.Y(n_133)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_19),
.Y(n_60)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_60),
.Y(n_115)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_21),
.Y(n_61)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_61),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_16),
.Y(n_62)
);

INVx6_ASAP7_75t_L g88 ( 
.A(n_62),
.Y(n_88)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_21),
.Y(n_63)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_63),
.Y(n_94)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_38),
.Y(n_64)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_64),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_16),
.Y(n_65)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_65),
.Y(n_117)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_33),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_66),
.Y(n_134)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_19),
.Y(n_67)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_67),
.Y(n_87)
);

INVx11_ASAP7_75t_L g68 ( 
.A(n_20),
.Y(n_68)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_68),
.Y(n_102)
);

INVx11_ASAP7_75t_L g69 ( 
.A(n_20),
.Y(n_69)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_69),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_20),
.Y(n_70)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_70),
.Y(n_118)
);

INVx4_ASAP7_75t_SL g71 ( 
.A(n_33),
.Y(n_71)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_71),
.Y(n_123)
);

OAI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_31),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_72),
.A2(n_17),
.B1(n_43),
.B2(n_18),
.Y(n_116)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_19),
.Y(n_73)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_73),
.Y(n_124)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_29),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g101 ( 
.A(n_74),
.B(n_76),
.Y(n_101)
);

INVx8_ASAP7_75t_L g75 ( 
.A(n_36),
.Y(n_75)
);

BUFx4f_ASAP7_75t_L g120 ( 
.A(n_75),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_31),
.Y(n_76)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_29),
.Y(n_77)
);

INVx8_ASAP7_75t_L g78 ( 
.A(n_36),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_78),
.B(n_79),
.Y(n_105)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_18),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_28),
.B(n_0),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_80),
.B(n_81),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_31),
.Y(n_81)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_29),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_82),
.B(n_83),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_28),
.B(n_0),
.Y(n_83)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_34),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_84),
.B(n_85),
.Y(n_113)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_34),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_34),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_86),
.B(n_36),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_64),
.B(n_23),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_97),
.B(n_121),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_47),
.Y(n_98)
);

CKINVDCx14_ASAP7_75t_R g143 ( 
.A(n_98),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_72),
.B(n_44),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_103),
.B(n_111),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_50),
.A2(n_23),
.B1(n_35),
.B2(n_22),
.Y(n_108)
);

AOI21xp5_ASAP7_75t_L g136 ( 
.A1(n_108),
.A2(n_39),
.B(n_46),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_71),
.A2(n_26),
.B1(n_32),
.B2(n_27),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_110),
.A2(n_112),
.B1(n_114),
.B2(n_125),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_49),
.B(n_44),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_75),
.A2(n_32),
.B1(n_26),
.B2(n_27),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_86),
.A2(n_22),
.B1(n_35),
.B2(n_17),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_116),
.A2(n_40),
.B1(n_2),
.B2(n_3),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_61),
.Y(n_121)
);

OA22x2_ASAP7_75t_L g122 ( 
.A1(n_73),
.A2(n_32),
.B1(n_26),
.B2(n_43),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g162 ( 
.A(n_122),
.B(n_130),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_52),
.A2(n_30),
.B1(n_39),
.B2(n_42),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_66),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_126),
.B(n_127),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_64),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_78),
.A2(n_27),
.B1(n_25),
.B2(n_30),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_132),
.A2(n_55),
.B1(n_42),
.B2(n_68),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_SL g219 ( 
.A1(n_136),
.A2(n_128),
.B(n_9),
.Y(n_219)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_131),
.Y(n_137)
);

INVx2_ASAP7_75t_SL g189 ( 
.A(n_137),
.Y(n_189)
);

INVx5_ASAP7_75t_L g138 ( 
.A(n_131),
.Y(n_138)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_138),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_104),
.B(n_74),
.C(n_57),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_139),
.B(n_179),
.C(n_170),
.Y(n_183)
);

OAI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_103),
.A2(n_81),
.B1(n_76),
.B2(n_70),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_142),
.A2(n_161),
.B1(n_173),
.B2(n_180),
.Y(n_190)
);

O2A1O1Ixp33_ASAP7_75t_L g144 ( 
.A1(n_122),
.A2(n_45),
.B(n_58),
.C(n_69),
.Y(n_144)
);

CKINVDCx16_ASAP7_75t_R g212 ( 
.A(n_144),
.Y(n_212)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_87),
.Y(n_146)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_146),
.Y(n_196)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_87),
.Y(n_147)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_147),
.Y(n_201)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_111),
.Y(n_148)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_148),
.Y(n_208)
);

INVxp67_ASAP7_75t_L g149 ( 
.A(n_91),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_149),
.B(n_151),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_116),
.B(n_65),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_150),
.B(n_156),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_105),
.Y(n_151)
);

CKINVDCx14_ASAP7_75t_R g152 ( 
.A(n_92),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_152),
.B(n_153),
.Y(n_199)
);

CKINVDCx16_ASAP7_75t_R g153 ( 
.A(n_123),
.Y(n_153)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_95),
.Y(n_155)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_155),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_108),
.B(n_62),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_107),
.B(n_59),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_157),
.B(n_168),
.Y(n_197)
);

AND2x4_ASAP7_75t_L g158 ( 
.A(n_122),
.B(n_38),
.Y(n_158)
);

NAND2x1_ASAP7_75t_L g221 ( 
.A(n_158),
.B(n_8),
.Y(n_221)
);

HB1xp67_ASAP7_75t_L g159 ( 
.A(n_129),
.Y(n_159)
);

INVxp67_ASAP7_75t_L g184 ( 
.A(n_159),
.Y(n_184)
);

BUFx2_ASAP7_75t_L g160 ( 
.A(n_135),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_160),
.Y(n_188)
);

AOI22xp33_ASAP7_75t_L g163 ( 
.A1(n_122),
.A2(n_27),
.B1(n_25),
.B2(n_42),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_163),
.A2(n_167),
.B1(n_119),
.B2(n_134),
.Y(n_209)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_124),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_164),
.B(n_165),
.Y(n_205)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_124),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_SL g166 ( 
.A1(n_123),
.A2(n_27),
.B1(n_25),
.B2(n_38),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_SL g215 ( 
.A1(n_166),
.A2(n_181),
.B1(n_119),
.B2(n_92),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_109),
.B(n_1),
.Y(n_168)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_95),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_169),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_101),
.A2(n_40),
.B1(n_5),
.B2(n_6),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g185 ( 
.A(n_170),
.Y(n_185)
);

BUFx2_ASAP7_75t_L g171 ( 
.A(n_135),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_171),
.Y(n_213)
);

INVx4_ASAP7_75t_L g172 ( 
.A(n_96),
.Y(n_172)
);

INVx8_ASAP7_75t_L g198 ( 
.A(n_172),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_113),
.A2(n_40),
.B1(n_5),
.B2(n_6),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_120),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_SL g222 ( 
.A(n_174),
.B(n_177),
.Y(n_222)
);

INVxp67_ASAP7_75t_L g175 ( 
.A(n_120),
.Y(n_175)
);

INVxp67_ASAP7_75t_L g186 ( 
.A(n_175),
.Y(n_186)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_115),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g204 ( 
.A(n_176),
.Y(n_204)
);

OR2x2_ASAP7_75t_L g177 ( 
.A(n_90),
.B(n_101),
.Y(n_177)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_115),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_178),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_101),
.B(n_40),
.C(n_6),
.Y(n_179)
);

OAI22xp33_ASAP7_75t_SL g180 ( 
.A1(n_88),
.A2(n_2),
.B1(n_6),
.B2(n_8),
.Y(n_180)
);

INVx5_ASAP7_75t_L g181 ( 
.A(n_96),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_118),
.Y(n_182)
);

INVxp67_ASAP7_75t_L g206 ( 
.A(n_182),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_183),
.B(n_178),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_148),
.A2(n_118),
.B1(n_88),
.B2(n_99),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_187),
.A2(n_194),
.B1(n_209),
.B2(n_210),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_162),
.A2(n_117),
.B1(n_102),
.B2(n_106),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_192),
.A2(n_218),
.B1(n_223),
.B2(n_177),
.Y(n_225)
);

OAI22xp33_ASAP7_75t_L g194 ( 
.A1(n_150),
.A2(n_89),
.B1(n_133),
.B2(n_93),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_145),
.B(n_106),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_200),
.B(n_202),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_145),
.B(n_102),
.Y(n_202)
);

A2O1A1Ixp33_ASAP7_75t_L g207 ( 
.A1(n_156),
.A2(n_98),
.B(n_120),
.C(n_90),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_SL g238 ( 
.A1(n_207),
.A2(n_219),
.B(n_179),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_162),
.A2(n_117),
.B1(n_133),
.B2(n_93),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_162),
.B(n_134),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_211),
.B(n_221),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_136),
.A2(n_99),
.B1(n_89),
.B2(n_100),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_214),
.A2(n_173),
.B1(n_176),
.B2(n_146),
.Y(n_242)
);

INVxp67_ASAP7_75t_L g227 ( 
.A(n_215),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_L g216 ( 
.A1(n_144),
.A2(n_94),
.B(n_100),
.Y(n_216)
);

AOI21xp5_ASAP7_75t_SL g226 ( 
.A1(n_216),
.A2(n_158),
.B(n_157),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_141),
.A2(n_129),
.B1(n_94),
.B2(n_128),
.Y(n_218)
);

OR2x4_ASAP7_75t_L g241 ( 
.A(n_221),
.B(n_208),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_158),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_225),
.A2(n_229),
.B1(n_242),
.B2(n_251),
.Y(n_276)
);

OAI21xp5_ASAP7_75t_SL g287 ( 
.A1(n_226),
.A2(n_240),
.B(n_243),
.Y(n_287)
);

AOI22xp33_ASAP7_75t_SL g228 ( 
.A1(n_215),
.A2(n_143),
.B1(n_171),
.B2(n_160),
.Y(n_228)
);

INVxp67_ASAP7_75t_L g285 ( 
.A(n_228),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_195),
.A2(n_158),
.B1(n_167),
.B2(n_139),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_196),
.Y(n_230)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_230),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_231),
.B(n_211),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_183),
.B(n_208),
.C(n_200),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_232),
.B(n_245),
.C(n_210),
.Y(n_281)
);

BUFx6f_ASAP7_75t_L g233 ( 
.A(n_198),
.Y(n_233)
);

BUFx3_ASAP7_75t_L g279 ( 
.A(n_233),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_191),
.B(n_140),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g283 ( 
.A(n_234),
.B(n_237),
.Y(n_283)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_196),
.Y(n_236)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_236),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_191),
.B(n_154),
.Y(n_237)
);

NAND2xp33_ASAP7_75t_SL g269 ( 
.A(n_238),
.B(n_241),
.Y(n_269)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_201),
.Y(n_239)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_239),
.Y(n_274)
);

A2O1A1Ixp33_ASAP7_75t_L g240 ( 
.A1(n_219),
.A2(n_168),
.B(n_149),
.C(n_147),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_185),
.A2(n_164),
.B1(n_165),
.B2(n_182),
.Y(n_243)
);

MAJx2_ASAP7_75t_L g244 ( 
.A(n_183),
.B(n_155),
.C(n_169),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_244),
.B(n_192),
.Y(n_272)
);

INVxp67_ASAP7_75t_L g246 ( 
.A(n_199),
.Y(n_246)
);

INVx13_ASAP7_75t_L g268 ( 
.A(n_246),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_197),
.B(n_137),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g288 ( 
.A(n_247),
.B(n_248),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_197),
.B(n_202),
.Y(n_248)
);

INVxp67_ASAP7_75t_L g249 ( 
.A(n_199),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_249),
.B(n_258),
.Y(n_267)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_201),
.Y(n_250)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_250),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_195),
.A2(n_175),
.B1(n_172),
.B2(n_181),
.Y(n_251)
);

INVx5_ASAP7_75t_L g252 ( 
.A(n_198),
.Y(n_252)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_252),
.Y(n_277)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_217),
.Y(n_253)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_253),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_190),
.A2(n_138),
.B1(n_11),
.B2(n_12),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_254),
.A2(n_187),
.B1(n_189),
.B2(n_188),
.Y(n_282)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_217),
.Y(n_255)
);

CKINVDCx16_ASAP7_75t_R g261 ( 
.A(n_255),
.Y(n_261)
);

BUFx3_ASAP7_75t_L g256 ( 
.A(n_198),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_256),
.Y(n_263)
);

OAI22x1_ASAP7_75t_L g257 ( 
.A1(n_216),
.A2(n_10),
.B1(n_13),
.B2(n_207),
.Y(n_257)
);

OAI22xp33_ASAP7_75t_L g280 ( 
.A1(n_257),
.A2(n_207),
.B1(n_209),
.B2(n_212),
.Y(n_280)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_193),
.Y(n_258)
);

OR2x2_ASAP7_75t_L g260 ( 
.A(n_257),
.B(n_216),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_260),
.B(n_264),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g306 ( 
.A(n_262),
.B(n_272),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_224),
.B(n_205),
.Y(n_264)
);

BUFx24_ASAP7_75t_SL g266 ( 
.A(n_246),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_266),
.B(n_290),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_SL g270 ( 
.A(n_249),
.B(n_222),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_SL g292 ( 
.A(n_270),
.B(n_273),
.Y(n_292)
);

OAI32xp33_ASAP7_75t_L g271 ( 
.A1(n_224),
.A2(n_212),
.A3(n_214),
.B1(n_222),
.B2(n_192),
.Y(n_271)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_271),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_SL g273 ( 
.A(n_232),
.B(n_205),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_229),
.B(n_223),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_278),
.B(n_284),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_280),
.A2(n_206),
.B1(n_218),
.B2(n_204),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_281),
.B(n_245),
.C(n_238),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_L g305 ( 
.A1(n_282),
.A2(n_235),
.B1(n_242),
.B2(n_190),
.Y(n_305)
);

OR2x2_ASAP7_75t_L g284 ( 
.A(n_243),
.B(n_223),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_251),
.B(n_184),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_SL g313 ( 
.A(n_286),
.B(n_186),
.Y(n_313)
);

AND2x6_ASAP7_75t_L g290 ( 
.A(n_244),
.B(n_221),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_291),
.B(n_297),
.C(n_299),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_283),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g339 ( 
.A(n_296),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_281),
.B(n_240),
.C(n_241),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_SL g298 ( 
.A1(n_260),
.A2(n_226),
.B(n_227),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_298),
.B(n_303),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_273),
.B(n_272),
.C(n_262),
.Y(n_299)
);

XOR2xp5_ASAP7_75t_L g301 ( 
.A(n_264),
.B(n_225),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_301),
.B(n_309),
.C(n_315),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_288),
.B(n_236),
.Y(n_302)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_302),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_279),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_265),
.Y(n_304)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_304),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_SL g324 ( 
.A1(n_305),
.A2(n_285),
.B1(n_276),
.B2(n_282),
.Y(n_324)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_279),
.Y(n_307)
);

INVx2_ASAP7_75t_L g320 ( 
.A(n_307),
.Y(n_320)
);

OAI21xp5_ASAP7_75t_SL g308 ( 
.A1(n_260),
.A2(n_227),
.B(n_221),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_308),
.B(n_313),
.Y(n_330)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_287),
.B(n_235),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_265),
.Y(n_310)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_310),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_267),
.B(n_239),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_311),
.B(n_314),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_SL g331 ( 
.A1(n_312),
.A2(n_274),
.B1(n_275),
.B2(n_259),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_270),
.B(n_258),
.Y(n_314)
);

XOR2xp5_ASAP7_75t_L g315 ( 
.A(n_287),
.B(n_193),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_268),
.B(n_213),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_316),
.B(n_213),
.Y(n_337)
);

AO22x1_ASAP7_75t_L g317 ( 
.A1(n_298),
.A2(n_271),
.B1(n_269),
.B2(n_284),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_317),
.Y(n_357)
);

AND2x6_ASAP7_75t_L g319 ( 
.A(n_300),
.B(n_268),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_319),
.B(n_327),
.Y(n_355)
);

OAI22xp5_ASAP7_75t_SL g344 ( 
.A1(n_324),
.A2(n_312),
.B1(n_295),
.B2(n_305),
.Y(n_344)
);

A2O1A1Ixp33_ASAP7_75t_SL g325 ( 
.A1(n_308),
.A2(n_269),
.B(n_284),
.C(n_290),
.Y(n_325)
);

AOI21xp5_ASAP7_75t_L g341 ( 
.A1(n_325),
.A2(n_309),
.B(n_294),
.Y(n_341)
);

OA21x2_ASAP7_75t_L g327 ( 
.A1(n_293),
.A2(n_278),
.B(n_268),
.Y(n_327)
);

OA21x2_ASAP7_75t_L g329 ( 
.A1(n_293),
.A2(n_277),
.B(n_276),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_329),
.B(n_303),
.Y(n_356)
);

AOI22xp5_ASAP7_75t_L g350 ( 
.A1(n_331),
.A2(n_333),
.B1(n_334),
.B2(n_310),
.Y(n_350)
);

OAI22xp5_ASAP7_75t_SL g333 ( 
.A1(n_295),
.A2(n_274),
.B1(n_275),
.B2(n_259),
.Y(n_333)
);

AOI211xp5_ASAP7_75t_L g334 ( 
.A1(n_294),
.A2(n_263),
.B(n_277),
.C(n_261),
.Y(n_334)
);

XOR2xp5_ASAP7_75t_L g335 ( 
.A(n_291),
.B(n_289),
.Y(n_335)
);

XOR2xp5_ASAP7_75t_L g342 ( 
.A(n_335),
.B(n_315),
.Y(n_342)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_299),
.B(n_261),
.C(n_289),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g351 ( 
.A(n_336),
.B(n_306),
.C(n_311),
.Y(n_351)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_337),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_292),
.B(n_188),
.Y(n_338)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_338),
.Y(n_348)
);

XNOR2xp5_ASAP7_75t_SL g369 ( 
.A(n_341),
.B(n_350),
.Y(n_369)
);

XOR2xp5_ASAP7_75t_L g371 ( 
.A(n_342),
.B(n_322),
.Y(n_371)
);

OAI21x1_ASAP7_75t_L g343 ( 
.A1(n_330),
.A2(n_292),
.B(n_314),
.Y(n_343)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_343),
.Y(n_361)
);

AOI22xp5_ASAP7_75t_L g370 ( 
.A1(n_344),
.A2(n_334),
.B1(n_326),
.B2(n_329),
.Y(n_370)
);

INVx3_ASAP7_75t_L g345 ( 
.A(n_339),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_345),
.B(n_346),
.Y(n_359)
);

BUFx5_ASAP7_75t_L g346 ( 
.A(n_320),
.Y(n_346)
);

AOI21xp5_ASAP7_75t_L g347 ( 
.A1(n_318),
.A2(n_297),
.B(n_301),
.Y(n_347)
);

OAI21xp5_ASAP7_75t_SL g363 ( 
.A1(n_347),
.A2(n_332),
.B(n_317),
.Y(n_363)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_333),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_349),
.B(n_350),
.Y(n_362)
);

MAJIxp5_ASAP7_75t_L g366 ( 
.A(n_351),
.B(n_352),
.C(n_353),
.Y(n_366)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_335),
.B(n_306),
.C(n_302),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g353 ( 
.A(n_328),
.B(n_304),
.C(n_296),
.Y(n_353)
);

XNOR2xp5_ASAP7_75t_L g354 ( 
.A(n_332),
.B(n_263),
.Y(n_354)
);

XNOR2xp5_ASAP7_75t_L g364 ( 
.A(n_354),
.B(n_342),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_356),
.B(n_322),
.Y(n_365)
);

MAJIxp5_ASAP7_75t_L g358 ( 
.A(n_328),
.B(n_256),
.C(n_233),
.Y(n_358)
);

MAJIxp5_ASAP7_75t_L g368 ( 
.A(n_358),
.B(n_331),
.C(n_324),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_SL g360 ( 
.A(n_340),
.B(n_336),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_SL g377 ( 
.A(n_360),
.B(n_367),
.Y(n_377)
);

AOI21xp5_ASAP7_75t_L g378 ( 
.A1(n_363),
.A2(n_341),
.B(n_347),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_L g383 ( 
.A(n_364),
.B(n_369),
.Y(n_383)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_365),
.Y(n_380)
);

XNOR2xp5_ASAP7_75t_L g367 ( 
.A(n_354),
.B(n_317),
.Y(n_367)
);

MAJIxp5_ASAP7_75t_L g376 ( 
.A(n_368),
.B(n_371),
.C(n_372),
.Y(n_376)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_370),
.Y(n_382)
);

MAJIxp5_ASAP7_75t_L g372 ( 
.A(n_358),
.B(n_326),
.C(n_319),
.Y(n_372)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_353),
.B(n_325),
.C(n_323),
.Y(n_373)
);

MAJIxp5_ASAP7_75t_L g379 ( 
.A(n_373),
.B(n_352),
.C(n_351),
.Y(n_379)
);

AOI21xp5_ASAP7_75t_L g374 ( 
.A1(n_361),
.A2(n_355),
.B(n_356),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_SL g391 ( 
.A(n_374),
.B(n_381),
.Y(n_391)
);

OR2x2_ASAP7_75t_L g375 ( 
.A(n_362),
.B(n_348),
.Y(n_375)
);

OAI22xp5_ASAP7_75t_SL g394 ( 
.A1(n_375),
.A2(n_384),
.B1(n_368),
.B2(n_325),
.Y(n_394)
);

XOR2xp5_ASAP7_75t_L g392 ( 
.A(n_378),
.B(n_373),
.Y(n_392)
);

XNOR2xp5_ASAP7_75t_L g386 ( 
.A(n_379),
.B(n_366),
.Y(n_386)
);

MAJIxp5_ASAP7_75t_L g381 ( 
.A(n_366),
.B(n_355),
.C(n_344),
.Y(n_381)
);

AOI22xp5_ASAP7_75t_L g384 ( 
.A1(n_369),
.A2(n_357),
.B1(n_329),
.B2(n_345),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_359),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_385),
.B(n_346),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_386),
.B(n_387),
.Y(n_401)
);

AOI22xp5_ASAP7_75t_L g387 ( 
.A1(n_382),
.A2(n_321),
.B1(n_371),
.B2(n_357),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_388),
.B(n_389),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_L g389 ( 
.A(n_375),
.B(n_381),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_380),
.B(n_372),
.Y(n_390)
);

XNOR2xp5_ASAP7_75t_L g396 ( 
.A(n_390),
.B(n_393),
.Y(n_396)
);

OR2x2_ASAP7_75t_L g397 ( 
.A(n_392),
.B(n_395),
.Y(n_397)
);

XNOR2xp5_ASAP7_75t_L g393 ( 
.A(n_379),
.B(n_364),
.Y(n_393)
);

XOR2xp5_ASAP7_75t_L g399 ( 
.A(n_394),
.B(n_395),
.Y(n_399)
);

XNOR2xp5_ASAP7_75t_L g395 ( 
.A(n_376),
.B(n_327),
.Y(n_395)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_397),
.Y(n_405)
);

AOI322xp5_ASAP7_75t_L g398 ( 
.A1(n_391),
.A2(n_374),
.A3(n_384),
.B1(n_383),
.B2(n_377),
.C1(n_325),
.C2(n_327),
.Y(n_398)
);

OAI21xp5_ASAP7_75t_SL g403 ( 
.A1(n_398),
.A2(n_400),
.B(n_189),
.Y(n_403)
);

AOI322xp5_ASAP7_75t_L g400 ( 
.A1(n_392),
.A2(n_376),
.A3(n_320),
.B1(n_307),
.B2(n_252),
.C1(n_220),
.C2(n_203),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_403),
.B(n_406),
.Y(n_408)
);

AOI21xp5_ASAP7_75t_L g404 ( 
.A1(n_402),
.A2(n_396),
.B(n_386),
.Y(n_404)
);

AOI21xp5_ASAP7_75t_SL g409 ( 
.A1(n_404),
.A2(n_400),
.B(n_398),
.Y(n_409)
);

OAI22xp5_ASAP7_75t_SL g406 ( 
.A1(n_401),
.A2(n_189),
.B1(n_203),
.B2(n_220),
.Y(n_406)
);

XOR2xp5_ASAP7_75t_L g407 ( 
.A(n_399),
.B(n_189),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_407),
.B(n_10),
.Y(n_410)
);

OAI21xp33_ASAP7_75t_SL g412 ( 
.A1(n_409),
.A2(n_410),
.B(n_406),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_SL g411 ( 
.A(n_408),
.B(n_405),
.Y(n_411)
);

MAJIxp5_ASAP7_75t_L g413 ( 
.A(n_411),
.B(n_412),
.C(n_407),
.Y(n_413)
);

AOI21xp5_ASAP7_75t_L g414 ( 
.A1(n_413),
.A2(n_13),
.B(n_389),
.Y(n_414)
);

XNOR2xp5_ASAP7_75t_L g415 ( 
.A(n_414),
.B(n_13),
.Y(n_415)
);


endmodule