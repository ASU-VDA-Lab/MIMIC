module fake_jpeg_14768_n_347 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_347);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_347;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx3_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_11),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

INVx11_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_1),
.Y(n_21)
);

INVx1_ASAP7_75t_SL g22 ( 
.A(n_9),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

BUFx16f_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_10),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

BUFx16f_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

INVx5_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_3),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_1),
.Y(n_36)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_24),
.Y(n_37)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_37),
.Y(n_59)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_25),
.Y(n_38)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_38),
.Y(n_62)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_39),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_36),
.Y(n_40)
);

CKINVDCx6p67_ASAP7_75t_R g74 ( 
.A(n_40),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_24),
.Y(n_41)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_41),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_36),
.Y(n_42)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

BUFx24_ASAP7_75t_L g43 ( 
.A(n_25),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g70 ( 
.A(n_43),
.Y(n_70)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_24),
.Y(n_44)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_44),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_45),
.Y(n_72)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_29),
.Y(n_46)
);

BUFx5_ASAP7_75t_L g58 ( 
.A(n_46),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_47),
.Y(n_52)
);

BUFx24_ASAP7_75t_L g48 ( 
.A(n_25),
.Y(n_48)
);

INVx11_ASAP7_75t_L g68 ( 
.A(n_48),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_29),
.Y(n_49)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_49),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_29),
.Y(n_50)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_50),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g51 ( 
.A(n_43),
.B(n_25),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_51),
.A2(n_21),
.B1(n_31),
.B2(n_17),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_37),
.A2(n_33),
.B1(n_44),
.B2(n_22),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_53),
.A2(n_64),
.B1(n_35),
.B2(n_21),
.Y(n_97)
);

AND2x2_ASAP7_75t_SL g55 ( 
.A(n_43),
.B(n_32),
.Y(n_55)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_55),
.B(n_48),
.C(n_22),
.Y(n_88)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_49),
.Y(n_56)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_56),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_38),
.A2(n_22),
.B1(n_33),
.B2(n_20),
.Y(n_61)
);

AOI21xp5_ASAP7_75t_L g95 ( 
.A1(n_61),
.A2(n_32),
.B(n_1),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_41),
.B(n_18),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_63),
.B(n_65),
.Y(n_81)
);

OA22x2_ASAP7_75t_L g64 ( 
.A1(n_50),
.A2(n_33),
.B1(n_32),
.B2(n_20),
.Y(n_64)
);

INVx2_ASAP7_75t_R g65 ( 
.A(n_48),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_40),
.B(n_18),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_69),
.B(n_30),
.Y(n_85)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_46),
.Y(n_73)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_73),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_55),
.B(n_19),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_76),
.B(n_80),
.Y(n_114)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_57),
.Y(n_78)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_78),
.Y(n_110)
);

INVx11_ASAP7_75t_L g79 ( 
.A(n_74),
.Y(n_79)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_79),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_55),
.B(n_19),
.Y(n_80)
);

INVxp67_ASAP7_75t_L g82 ( 
.A(n_65),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_82),
.B(n_85),
.Y(n_121)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_70),
.Y(n_83)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_83),
.Y(n_139)
);

BUFx4f_ASAP7_75t_SL g84 ( 
.A(n_70),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_84),
.Y(n_126)
);

BUFx2_ASAP7_75t_L g86 ( 
.A(n_56),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_86),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_59),
.B(n_30),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_87),
.B(n_91),
.Y(n_137)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_88),
.B(n_101),
.Y(n_116)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_73),
.Y(n_89)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_89),
.Y(n_133)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_67),
.Y(n_90)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_90),
.Y(n_138)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_57),
.Y(n_91)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_67),
.Y(n_92)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_92),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_51),
.B(n_46),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_93),
.B(n_99),
.Y(n_122)
);

OAI22xp33_ASAP7_75t_L g94 ( 
.A1(n_60),
.A2(n_20),
.B1(n_45),
.B2(n_42),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_94),
.A2(n_98),
.B1(n_74),
.B2(n_1),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_SL g131 ( 
.A1(n_95),
.A2(n_26),
.B(n_23),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_65),
.B(n_47),
.C(n_32),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_96),
.B(n_106),
.C(n_27),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_97),
.A2(n_100),
.B1(n_68),
.B2(n_26),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_60),
.A2(n_66),
.B1(n_54),
.B2(n_72),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_59),
.B(n_35),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_54),
.A2(n_31),
.B1(n_29),
.B2(n_34),
.Y(n_100)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_72),
.Y(n_102)
);

CKINVDCx16_ASAP7_75t_R g112 ( 
.A(n_102),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_L g103 ( 
.A1(n_66),
.A2(n_31),
.B1(n_34),
.B2(n_28),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_103),
.A2(n_52),
.B1(n_71),
.B2(n_64),
.Y(n_113)
);

INVx2_ASAP7_75t_SL g104 ( 
.A(n_70),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_104),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_51),
.B(n_28),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_105),
.B(n_68),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_70),
.B(n_27),
.C(n_17),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_71),
.Y(n_107)
);

OR2x2_ASAP7_75t_L g111 ( 
.A(n_107),
.B(n_108),
.Y(n_111)
);

O2A1O1Ixp33_ASAP7_75t_L g108 ( 
.A1(n_64),
.A2(n_28),
.B(n_17),
.C(n_31),
.Y(n_108)
);

BUFx3_ASAP7_75t_L g109 ( 
.A(n_52),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_109),
.Y(n_132)
);

OAI22xp33_ASAP7_75t_SL g158 ( 
.A1(n_113),
.A2(n_86),
.B1(n_109),
.B2(n_75),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_117),
.B(n_96),
.Y(n_146)
);

O2A1O1Ixp33_ASAP7_75t_L g118 ( 
.A1(n_95),
.A2(n_64),
.B(n_74),
.C(n_62),
.Y(n_118)
);

CKINVDCx16_ASAP7_75t_R g149 ( 
.A(n_118),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_88),
.B(n_58),
.C(n_27),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_119),
.B(n_106),
.C(n_58),
.Y(n_162)
);

O2A1O1Ixp33_ASAP7_75t_SL g123 ( 
.A1(n_76),
.A2(n_74),
.B(n_62),
.C(n_34),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_SL g165 ( 
.A1(n_123),
.A2(n_86),
.B(n_26),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_124),
.A2(n_136),
.B1(n_100),
.B2(n_87),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_101),
.A2(n_108),
.B1(n_97),
.B2(n_93),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_125),
.A2(n_84),
.B1(n_13),
.B2(n_12),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_127),
.A2(n_98),
.B1(n_102),
.B2(n_91),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_128),
.B(n_107),
.Y(n_148)
);

BUFx5_ASAP7_75t_L g129 ( 
.A(n_84),
.Y(n_129)
);

INVx4_ASAP7_75t_L g143 ( 
.A(n_129),
.Y(n_143)
);

AOI21xp5_ASAP7_75t_L g150 ( 
.A1(n_131),
.A2(n_78),
.B(n_2),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_80),
.B(n_0),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_135),
.B(n_99),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_105),
.A2(n_11),
.B1(n_16),
.B2(n_15),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_140),
.A2(n_155),
.B1(n_158),
.B2(n_168),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_SL g185 ( 
.A(n_141),
.B(n_151),
.Y(n_185)
);

NOR2x1_ASAP7_75t_L g142 ( 
.A(n_111),
.B(n_81),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_L g175 ( 
.A1(n_142),
.A2(n_150),
.B(n_157),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_111),
.B(n_81),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_144),
.B(n_148),
.Y(n_174)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_134),
.Y(n_145)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_145),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_146),
.B(n_162),
.C(n_170),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_147),
.A2(n_166),
.B1(n_127),
.B2(n_122),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_137),
.B(n_90),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_110),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_152),
.B(n_163),
.Y(n_184)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_134),
.Y(n_153)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_153),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_111),
.B(n_92),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_154),
.B(n_160),
.Y(n_190)
);

AOI22xp33_ASAP7_75t_SL g155 ( 
.A1(n_126),
.A2(n_79),
.B1(n_104),
.B2(n_89),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_134),
.Y(n_156)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_156),
.Y(n_180)
);

AOI21xp5_ASAP7_75t_L g157 ( 
.A1(n_131),
.A2(n_77),
.B(n_75),
.Y(n_157)
);

INVx8_ASAP7_75t_L g159 ( 
.A(n_129),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_159),
.B(n_129),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_114),
.B(n_85),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_137),
.B(n_77),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_SL g191 ( 
.A(n_161),
.B(n_121),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_110),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_138),
.Y(n_164)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_164),
.Y(n_182)
);

AOI21xp5_ASAP7_75t_L g186 ( 
.A1(n_165),
.A2(n_171),
.B(n_116),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_124),
.A2(n_104),
.B1(n_23),
.B2(n_84),
.Y(n_166)
);

A2O1A1Ixp33_ASAP7_75t_L g167 ( 
.A1(n_114),
.A2(n_23),
.B(n_11),
.C(n_16),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_167),
.B(n_136),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_116),
.A2(n_8),
.B1(n_15),
.B2(n_14),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g188 ( 
.A(n_169),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_117),
.B(n_119),
.C(n_128),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_SL g171 ( 
.A1(n_116),
.A2(n_83),
.B(n_2),
.Y(n_171)
);

CKINVDCx14_ASAP7_75t_R g218 ( 
.A(n_173),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_161),
.B(n_126),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_SL g229 ( 
.A(n_177),
.B(n_179),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_143),
.B(n_139),
.Y(n_179)
);

CKINVDCx16_ASAP7_75t_R g181 ( 
.A(n_145),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_181),
.B(n_189),
.Y(n_213)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_153),
.Y(n_183)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_183),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_SL g230 ( 
.A1(n_186),
.A2(n_193),
.B(n_198),
.Y(n_230)
);

BUFx6f_ASAP7_75t_L g187 ( 
.A(n_159),
.Y(n_187)
);

INVx4_ASAP7_75t_L g227 ( 
.A(n_187),
.Y(n_227)
);

INVxp67_ASAP7_75t_L g189 ( 
.A(n_169),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_191),
.B(n_192),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_141),
.B(n_121),
.Y(n_192)
);

INVxp33_ASAP7_75t_SL g194 ( 
.A(n_142),
.Y(n_194)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_194),
.Y(n_216)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_156),
.Y(n_195)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_195),
.Y(n_217)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_151),
.Y(n_196)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_196),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_148),
.B(n_116),
.Y(n_197)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_197),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_149),
.A2(n_125),
.B1(n_118),
.B2(n_113),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_199),
.A2(n_204),
.B1(n_157),
.B2(n_150),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_140),
.A2(n_118),
.B1(n_122),
.B2(n_123),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_200),
.A2(n_206),
.B1(n_189),
.B2(n_188),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_170),
.B(n_135),
.C(n_120),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_202),
.B(n_171),
.C(n_160),
.Y(n_225)
);

INVx3_ASAP7_75t_SL g203 ( 
.A(n_164),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_203),
.B(n_120),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_149),
.A2(n_123),
.B1(n_130),
.B2(n_112),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_154),
.Y(n_205)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_205),
.Y(n_228)
);

AND2x2_ASAP7_75t_L g206 ( 
.A(n_142),
.B(n_130),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_SL g232 ( 
.A1(n_206),
.A2(n_191),
.B(n_197),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_185),
.B(n_144),
.Y(n_207)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_207),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_L g248 ( 
.A1(n_208),
.A2(n_215),
.B1(n_223),
.B2(n_199),
.Y(n_248)
);

CKINVDCx14_ASAP7_75t_R g247 ( 
.A(n_210),
.Y(n_247)
);

INVxp67_ASAP7_75t_L g211 ( 
.A(n_184),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_211),
.B(n_222),
.Y(n_242)
);

HB1xp67_ASAP7_75t_L g212 ( 
.A(n_176),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_212),
.B(n_195),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_188),
.A2(n_147),
.B1(n_166),
.B2(n_165),
.Y(n_215)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_220),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_185),
.B(n_152),
.Y(n_221)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_221),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_182),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_206),
.A2(n_162),
.B1(n_146),
.B2(n_163),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_225),
.B(n_226),
.C(n_202),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_201),
.B(n_186),
.Y(n_226)
);

AOI21xp5_ASAP7_75t_L g231 ( 
.A1(n_175),
.A2(n_205),
.B(n_196),
.Y(n_231)
);

AOI21xp5_ASAP7_75t_L g258 ( 
.A1(n_231),
.A2(n_232),
.B(n_235),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_187),
.B(n_143),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_233),
.B(n_211),
.Y(n_239)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_182),
.Y(n_234)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_234),
.Y(n_255)
);

OAI21xp5_ASAP7_75t_L g235 ( 
.A1(n_175),
.A2(n_167),
.B(n_168),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_208),
.A2(n_198),
.B1(n_174),
.B2(n_190),
.Y(n_236)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_236),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_221),
.B(n_190),
.Y(n_237)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_237),
.Y(n_270)
);

INVxp67_ASAP7_75t_L g238 ( 
.A(n_213),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_238),
.B(n_241),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_239),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_207),
.B(n_174),
.Y(n_241)
);

NAND2xp67_ASAP7_75t_SL g243 ( 
.A(n_232),
.B(n_193),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_243),
.B(n_246),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_226),
.B(n_201),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_244),
.B(n_210),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_245),
.B(n_249),
.C(n_257),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_219),
.B(n_203),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_248),
.A2(n_260),
.B1(n_216),
.B2(n_224),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_223),
.B(n_204),
.C(n_176),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_219),
.B(n_203),
.Y(n_250)
);

HB1xp67_ASAP7_75t_L g264 ( 
.A(n_250),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_231),
.B(n_172),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_251),
.B(n_252),
.C(n_215),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_230),
.B(n_159),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_256),
.B(n_214),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_225),
.B(n_183),
.C(n_180),
.Y(n_257)
);

AND2x6_ASAP7_75t_L g259 ( 
.A(n_230),
.B(n_180),
.Y(n_259)
);

OAI21xp5_ASAP7_75t_SL g273 ( 
.A1(n_259),
.A2(n_216),
.B(n_228),
.Y(n_273)
);

INVx1_ASAP7_75t_SL g260 ( 
.A(n_222),
.Y(n_260)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_261),
.Y(n_284)
);

XOR2xp5_ASAP7_75t_L g292 ( 
.A(n_265),
.B(n_268),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_244),
.B(n_245),
.C(n_257),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_266),
.B(n_272),
.C(n_274),
.Y(n_283)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_249),
.B(n_235),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_SL g298 ( 
.A(n_269),
.B(n_241),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_271),
.B(n_238),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_252),
.B(n_218),
.Y(n_272)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_273),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_251),
.B(n_228),
.C(n_224),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_247),
.A2(n_217),
.B1(n_209),
.B2(n_234),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_277),
.A2(n_255),
.B1(n_240),
.B2(n_237),
.Y(n_297)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_258),
.B(n_229),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_278),
.B(n_279),
.C(n_280),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_236),
.B(n_217),
.C(n_209),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_258),
.B(n_178),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_246),
.B(n_178),
.C(n_139),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_281),
.B(n_260),
.C(n_242),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_267),
.A2(n_243),
.B1(n_259),
.B2(n_254),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_282),
.A2(n_255),
.B1(n_268),
.B2(n_263),
.Y(n_299)
);

AND2x2_ASAP7_75t_L g286 ( 
.A(n_278),
.B(n_250),
.Y(n_286)
);

AOI21xp5_ASAP7_75t_L g300 ( 
.A1(n_286),
.A2(n_288),
.B(n_265),
.Y(n_300)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_281),
.Y(n_287)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_287),
.Y(n_302)
);

AND2x2_ASAP7_75t_L g288 ( 
.A(n_275),
.B(n_274),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_SL g310 ( 
.A(n_289),
.B(n_293),
.Y(n_310)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_262),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_290),
.B(n_291),
.Y(n_305)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_270),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_276),
.B(n_253),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_295),
.B(n_133),
.C(n_115),
.Y(n_312)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_279),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_296),
.B(n_288),
.Y(n_307)
);

INVxp67_ASAP7_75t_L g301 ( 
.A(n_297),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g311 ( 
.A(n_298),
.B(n_132),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_L g316 ( 
.A1(n_299),
.A2(n_294),
.B1(n_283),
.B2(n_292),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_SL g323 ( 
.A(n_300),
.B(n_307),
.C(n_13),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_286),
.A2(n_227),
.B1(n_264),
.B2(n_263),
.Y(n_303)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_303),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_SL g304 ( 
.A(n_282),
.B(n_266),
.Y(n_304)
);

XOR2xp5_ASAP7_75t_L g317 ( 
.A(n_304),
.B(n_308),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_295),
.B(n_227),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_306),
.B(n_309),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_SL g308 ( 
.A(n_298),
.B(n_112),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_285),
.B(n_138),
.Y(n_309)
);

XOR2xp5_ASAP7_75t_L g321 ( 
.A(n_311),
.B(n_133),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_312),
.B(n_292),
.Y(n_320)
);

BUFx2_ASAP7_75t_L g313 ( 
.A(n_284),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_313),
.B(n_294),
.Y(n_314)
);

XOR2xp5_ASAP7_75t_L g333 ( 
.A(n_314),
.B(n_320),
.Y(n_333)
);

AOI322xp5_ASAP7_75t_L g327 ( 
.A1(n_316),
.A2(n_324),
.A3(n_325),
.B1(n_304),
.B2(n_312),
.C1(n_9),
.C2(n_8),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_313),
.B(n_283),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_SL g326 ( 
.A(n_318),
.B(n_322),
.Y(n_326)
);

XOR2xp5_ASAP7_75t_L g328 ( 
.A(n_321),
.B(n_323),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_310),
.B(n_13),
.Y(n_322)
);

OAI211xp5_ASAP7_75t_L g324 ( 
.A1(n_305),
.A2(n_301),
.B(n_302),
.C(n_308),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_301),
.B(n_12),
.Y(n_325)
);

OR2x2_ASAP7_75t_L g340 ( 
.A(n_327),
.B(n_329),
.Y(n_340)
);

AOI322xp5_ASAP7_75t_L g329 ( 
.A1(n_319),
.A2(n_8),
.A3(n_2),
.B1(n_3),
.B2(n_4),
.C1(n_0),
.C2(n_6),
.Y(n_329)
);

OR2x2_ASAP7_75t_L g330 ( 
.A(n_323),
.B(n_0),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_330),
.B(n_332),
.Y(n_335)
);

NOR2x1_ASAP7_75t_SL g331 ( 
.A(n_321),
.B(n_2),
.Y(n_331)
);

NOR3xp33_ASAP7_75t_L g336 ( 
.A(n_331),
.B(n_5),
.C(n_6),
.Y(n_336)
);

OAI21xp5_ASAP7_75t_L g332 ( 
.A1(n_315),
.A2(n_4),
.B(n_5),
.Y(n_332)
);

XOR2xp5_ASAP7_75t_L g334 ( 
.A(n_317),
.B(n_4),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_334),
.B(n_317),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_336),
.B(n_337),
.Y(n_341)
);

OAI21xp5_ASAP7_75t_SL g338 ( 
.A1(n_326),
.A2(n_5),
.B(n_6),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_338),
.B(n_333),
.C(n_7),
.Y(n_343)
);

AOI22xp33_ASAP7_75t_SL g339 ( 
.A1(n_328),
.A2(n_7),
.B1(n_330),
.B2(n_334),
.Y(n_339)
);

AND2x2_ASAP7_75t_L g342 ( 
.A(n_339),
.B(n_328),
.Y(n_342)
);

AOI21xp5_ASAP7_75t_L g344 ( 
.A1(n_342),
.A2(n_343),
.B(n_335),
.Y(n_344)
);

XOR2xp5_ASAP7_75t_L g345 ( 
.A(n_344),
.B(n_341),
.Y(n_345)
);

AOI21xp5_ASAP7_75t_L g346 ( 
.A1(n_345),
.A2(n_340),
.B(n_7),
.Y(n_346)
);

XNOR2xp5_ASAP7_75t_L g347 ( 
.A(n_346),
.B(n_7),
.Y(n_347)
);


endmodule