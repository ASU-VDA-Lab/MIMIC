module fake_netlist_5_151_n_2092 (n_137, n_294, n_318, n_82, n_194, n_316, n_248, n_124, n_86, n_136, n_146, n_315, n_268, n_61, n_127, n_75, n_235, n_226, n_74, n_57, n_111, n_155, n_43, n_116, n_22, n_284, n_46, n_245, n_21, n_139, n_38, n_105, n_280, n_4, n_17, n_254, n_33, n_23, n_302, n_265, n_293, n_244, n_47, n_173, n_198, n_247, n_314, n_8, n_321, n_292, n_100, n_212, n_119, n_275, n_252, n_26, n_295, n_133, n_330, n_2, n_6, n_39, n_147, n_67, n_307, n_87, n_150, n_106, n_209, n_259, n_301, n_68, n_93, n_186, n_134, n_191, n_51, n_63, n_171, n_153, n_204, n_250, n_260, n_298, n_320, n_286, n_122, n_282, n_331, n_10, n_24, n_325, n_132, n_90, n_101, n_281, n_240, n_189, n_220, n_291, n_231, n_257, n_31, n_13, n_152, n_317, n_9, n_323, n_195, n_42, n_227, n_45, n_271, n_94, n_123, n_167, n_234, n_308, n_267, n_297, n_156, n_5, n_225, n_219, n_157, n_131, n_192, n_223, n_158, n_138, n_264, n_109, n_163, n_276, n_95, n_183, n_185, n_243, n_169, n_59, n_255, n_215, n_196, n_211, n_218, n_181, n_3, n_290, n_221, n_178, n_287, n_72, n_104, n_41, n_56, n_141, n_15, n_145, n_48, n_50, n_313, n_88, n_216, n_168, n_164, n_311, n_208, n_142, n_214, n_328, n_140, n_299, n_303, n_296, n_241, n_184, n_65, n_78, n_144, n_114, n_96, n_165, n_213, n_129, n_98, n_197, n_107, n_69, n_236, n_1, n_249, n_304, n_329, n_203, n_274, n_80, n_35, n_73, n_277, n_92, n_19, n_149, n_333, n_309, n_30, n_14, n_84, n_130, n_322, n_258, n_29, n_79, n_151, n_25, n_306, n_288, n_188, n_190, n_201, n_263, n_44, n_224, n_40, n_34, n_228, n_283, n_112, n_85, n_239, n_55, n_49, n_310, n_54, n_12, n_76, n_170, n_332, n_27, n_77, n_102, n_161, n_273, n_270, n_230, n_81, n_118, n_279, n_70, n_253, n_261, n_174, n_289, n_172, n_206, n_217, n_312, n_210, n_91, n_176, n_182, n_143, n_83, n_237, n_180, n_207, n_37, n_229, n_108, n_66, n_177, n_60, n_16, n_0, n_58, n_18, n_117, n_326, n_233, n_205, n_113, n_246, n_179, n_125, n_269, n_128, n_285, n_120, n_232, n_327, n_135, n_126, n_202, n_266, n_272, n_193, n_251, n_53, n_160, n_154, n_62, n_148, n_71, n_300, n_159, n_334, n_175, n_262, n_238, n_99, n_319, n_20, n_121, n_242, n_36, n_200, n_162, n_64, n_222, n_28, n_89, n_115, n_324, n_199, n_187, n_32, n_103, n_97, n_166, n_11, n_7, n_256, n_305, n_52, n_278, n_110, n_2092);

input n_137;
input n_294;
input n_318;
input n_82;
input n_194;
input n_316;
input n_248;
input n_124;
input n_86;
input n_136;
input n_146;
input n_315;
input n_268;
input n_61;
input n_127;
input n_75;
input n_235;
input n_226;
input n_74;
input n_57;
input n_111;
input n_155;
input n_43;
input n_116;
input n_22;
input n_284;
input n_46;
input n_245;
input n_21;
input n_139;
input n_38;
input n_105;
input n_280;
input n_4;
input n_17;
input n_254;
input n_33;
input n_23;
input n_302;
input n_265;
input n_293;
input n_244;
input n_47;
input n_173;
input n_198;
input n_247;
input n_314;
input n_8;
input n_321;
input n_292;
input n_100;
input n_212;
input n_119;
input n_275;
input n_252;
input n_26;
input n_295;
input n_133;
input n_330;
input n_2;
input n_6;
input n_39;
input n_147;
input n_67;
input n_307;
input n_87;
input n_150;
input n_106;
input n_209;
input n_259;
input n_301;
input n_68;
input n_93;
input n_186;
input n_134;
input n_191;
input n_51;
input n_63;
input n_171;
input n_153;
input n_204;
input n_250;
input n_260;
input n_298;
input n_320;
input n_286;
input n_122;
input n_282;
input n_331;
input n_10;
input n_24;
input n_325;
input n_132;
input n_90;
input n_101;
input n_281;
input n_240;
input n_189;
input n_220;
input n_291;
input n_231;
input n_257;
input n_31;
input n_13;
input n_152;
input n_317;
input n_9;
input n_323;
input n_195;
input n_42;
input n_227;
input n_45;
input n_271;
input n_94;
input n_123;
input n_167;
input n_234;
input n_308;
input n_267;
input n_297;
input n_156;
input n_5;
input n_225;
input n_219;
input n_157;
input n_131;
input n_192;
input n_223;
input n_158;
input n_138;
input n_264;
input n_109;
input n_163;
input n_276;
input n_95;
input n_183;
input n_185;
input n_243;
input n_169;
input n_59;
input n_255;
input n_215;
input n_196;
input n_211;
input n_218;
input n_181;
input n_3;
input n_290;
input n_221;
input n_178;
input n_287;
input n_72;
input n_104;
input n_41;
input n_56;
input n_141;
input n_15;
input n_145;
input n_48;
input n_50;
input n_313;
input n_88;
input n_216;
input n_168;
input n_164;
input n_311;
input n_208;
input n_142;
input n_214;
input n_328;
input n_140;
input n_299;
input n_303;
input n_296;
input n_241;
input n_184;
input n_65;
input n_78;
input n_144;
input n_114;
input n_96;
input n_165;
input n_213;
input n_129;
input n_98;
input n_197;
input n_107;
input n_69;
input n_236;
input n_1;
input n_249;
input n_304;
input n_329;
input n_203;
input n_274;
input n_80;
input n_35;
input n_73;
input n_277;
input n_92;
input n_19;
input n_149;
input n_333;
input n_309;
input n_30;
input n_14;
input n_84;
input n_130;
input n_322;
input n_258;
input n_29;
input n_79;
input n_151;
input n_25;
input n_306;
input n_288;
input n_188;
input n_190;
input n_201;
input n_263;
input n_44;
input n_224;
input n_40;
input n_34;
input n_228;
input n_283;
input n_112;
input n_85;
input n_239;
input n_55;
input n_49;
input n_310;
input n_54;
input n_12;
input n_76;
input n_170;
input n_332;
input n_27;
input n_77;
input n_102;
input n_161;
input n_273;
input n_270;
input n_230;
input n_81;
input n_118;
input n_279;
input n_70;
input n_253;
input n_261;
input n_174;
input n_289;
input n_172;
input n_206;
input n_217;
input n_312;
input n_210;
input n_91;
input n_176;
input n_182;
input n_143;
input n_83;
input n_237;
input n_180;
input n_207;
input n_37;
input n_229;
input n_108;
input n_66;
input n_177;
input n_60;
input n_16;
input n_0;
input n_58;
input n_18;
input n_117;
input n_326;
input n_233;
input n_205;
input n_113;
input n_246;
input n_179;
input n_125;
input n_269;
input n_128;
input n_285;
input n_120;
input n_232;
input n_327;
input n_135;
input n_126;
input n_202;
input n_266;
input n_272;
input n_193;
input n_251;
input n_53;
input n_160;
input n_154;
input n_62;
input n_148;
input n_71;
input n_300;
input n_159;
input n_334;
input n_175;
input n_262;
input n_238;
input n_99;
input n_319;
input n_20;
input n_121;
input n_242;
input n_36;
input n_200;
input n_162;
input n_64;
input n_222;
input n_28;
input n_89;
input n_115;
input n_324;
input n_199;
input n_187;
input n_32;
input n_103;
input n_97;
input n_166;
input n_11;
input n_7;
input n_256;
input n_305;
input n_52;
input n_278;
input n_110;

output n_2092;

wire n_924;
wire n_1263;
wire n_1378;
wire n_977;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1729;
wire n_1166;
wire n_1751;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1859;
wire n_1677;
wire n_1150;
wire n_1780;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1360;
wire n_1198;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1738;
wire n_2021;
wire n_1021;
wire n_1960;
wire n_551;
wire n_2059;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1695;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_1789;
wire n_1666;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_1545;
wire n_864;
wire n_859;
wire n_951;
wire n_1947;
wire n_1264;
wire n_447;
wire n_2001;
wire n_1494;
wire n_625;
wire n_854;
wire n_1462;
wire n_1799;
wire n_2069;
wire n_1580;
wire n_674;
wire n_417;
wire n_1939;
wire n_1806;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_1869;
wire n_1607;
wire n_1563;
wire n_606;
wire n_2011;
wire n_877;
wire n_2024;
wire n_1696;
wire n_755;
wire n_1118;
wire n_1686;
wire n_947;
wire n_1285;
wire n_373;
wire n_1860;
wire n_1359;
wire n_530;
wire n_1107;
wire n_1728;
wire n_556;
wire n_2031;
wire n_2076;
wire n_1230;
wire n_668;
wire n_375;
wire n_1896;
wire n_929;
wire n_1124;
wire n_1818;
wire n_902;
wire n_1576;
wire n_1104;
wire n_1294;
wire n_1705;
wire n_659;
wire n_1257;
wire n_1182;
wire n_579;
wire n_1698;
wire n_1261;
wire n_938;
wire n_1098;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_406;
wire n_519;
wire n_1016;
wire n_1243;
wire n_546;
wire n_2047;
wire n_1280;
wire n_1845;
wire n_2052;
wire n_2058;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_1236;
wire n_1633;
wire n_569;
wire n_1778;
wire n_920;
wire n_1289;
wire n_1517;
wire n_2091;
wire n_335;
wire n_2085;
wire n_1669;
wire n_370;
wire n_976;
wire n_1949;
wire n_343;
wire n_1449;
wire n_1946;
wire n_1566;
wire n_2032;
wire n_1078;
wire n_1670;
wire n_775;
wire n_600;
wire n_1484;
wire n_2071;
wire n_1374;
wire n_1328;
wire n_1948;
wire n_1984;
wire n_1877;
wire n_1831;
wire n_1598;
wire n_1723;
wire n_955;
wire n_1850;
wire n_339;
wire n_1146;
wire n_882;
wire n_1036;
wire n_1097;
wire n_1749;
wire n_347;
wire n_696;
wire n_550;
wire n_897;
wire n_350;
wire n_798;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_580;
wire n_1040;
wire n_1872;
wire n_1852;
wire n_578;
wire n_926;
wire n_344;
wire n_1218;
wire n_1931;
wire n_422;
wire n_1070;
wire n_1547;
wire n_777;
wire n_475;
wire n_2089;
wire n_1030;
wire n_1755;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1801;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_663;
wire n_845;
wire n_1862;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_1796;
wire n_680;
wire n_1473;
wire n_1587;
wire n_395;
wire n_901;
wire n_553;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_1748;
wire n_1672;
wire n_675;
wire n_888;
wire n_1880;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1384;
wire n_1556;
wire n_446;
wire n_1863;
wire n_1064;
wire n_858;
wire n_2079;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_1706;
wire n_468;
wire n_342;
wire n_464;
wire n_363;
wire n_1582;
wire n_1069;
wire n_1784;
wire n_1075;
wire n_1836;
wire n_1450;
wire n_1322;
wire n_1471;
wire n_1986;
wire n_2072;
wire n_1750;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_1700;
wire n_477;
wire n_1585;
wire n_571;
wire n_461;
wire n_1971;
wire n_1599;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_1950;
wire n_907;
wire n_1447;
wire n_1377;
wire n_989;
wire n_1039;
wire n_2055;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_2062;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_1667;
wire n_838;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1926;
wire n_1248;
wire n_1331;
wire n_953;
wire n_1014;
wire n_1241;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_1819;
wire n_476;
wire n_1527;
wire n_2042;
wire n_534;
wire n_1882;
wire n_884;
wire n_345;
wire n_944;
wire n_1754;
wire n_1623;
wire n_1854;
wire n_1565;
wire n_1809;
wire n_1856;
wire n_647;
wire n_407;
wire n_1072;
wire n_832;
wire n_857;
wire n_1319;
wire n_561;
wire n_1825;
wire n_1951;
wire n_1883;
wire n_1906;
wire n_1712;
wire n_1387;
wire n_1532;
wire n_1027;
wire n_971;
wire n_1156;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1775;
wire n_2028;
wire n_1368;
wire n_558;
wire n_1276;
wire n_702;
wire n_822;
wire n_1412;
wire n_1709;
wire n_728;
wire n_1162;
wire n_1538;
wire n_1838;
wire n_1199;
wire n_1847;
wire n_1779;
wire n_352;
wire n_1884;
wire n_1038;
wire n_1369;
wire n_520;
wire n_409;
wire n_1841;
wire n_1660;
wire n_887;
wire n_1905;
wire n_809;
wire n_870;
wire n_931;
wire n_599;
wire n_1711;
wire n_1662;
wire n_1891;
wire n_1481;
wire n_1942;
wire n_434;
wire n_1978;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1629;
wire n_1293;
wire n_965;
wire n_1876;
wire n_1743;
wire n_935;
wire n_817;
wire n_1175;
wire n_360;
wire n_1479;
wire n_1810;
wire n_1888;
wire n_2009;
wire n_759;
wire n_1892;
wire n_806;
wire n_1997;
wire n_1766;
wire n_1477;
wire n_1635;
wire n_1963;
wire n_1571;
wire n_1189;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_2064;
wire n_784;
wire n_1733;
wire n_1244;
wire n_431;
wire n_1925;
wire n_1194;
wire n_1815;
wire n_851;
wire n_615;
wire n_1759;
wire n_843;
wire n_1788;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_1679;
wire n_776;
wire n_1798;
wire n_2022;
wire n_1790;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1746;
wire n_1647;
wire n_1829;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_1674;
wire n_1833;
wire n_1830;
wire n_2073;
wire n_1710;
wire n_1128;
wire n_1734;
wire n_744;
wire n_590;
wire n_629;
wire n_1308;
wire n_1767;
wire n_1680;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_2005;
wire n_526;
wire n_1916;
wire n_372;
wire n_677;
wire n_1333;
wire n_1121;
wire n_433;
wire n_604;
wire n_368;
wire n_2007;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_2054;
wire n_498;
wire n_1468;
wire n_1559;
wire n_1765;
wire n_1866;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_624;
wire n_1380;
wire n_1744;
wire n_1617;
wire n_1010;
wire n_1994;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_1837;
wire n_1839;
wire n_610;
wire n_1760;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_1832;
wire n_448;
wire n_1851;
wire n_999;
wire n_758;
wire n_2046;
wire n_1933;
wire n_1656;
wire n_1158;
wire n_2045;
wire n_1509;
wire n_1874;
wire n_2040;
wire n_563;
wire n_2060;
wire n_1987;
wire n_1145;
wire n_878;
wire n_524;
wire n_394;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_1871;
wire n_1964;
wire n_906;
wire n_1163;
wire n_2039;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_1781;
wire n_2084;
wire n_2035;
wire n_658;
wire n_2061;
wire n_1740;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_1923;
wire n_1773;
wire n_592;
wire n_1169;
wire n_1596;
wire n_1692;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_1095;
wire n_1828;
wire n_1614;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_2038;
wire n_603;
wire n_1431;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_2087;
wire n_1640;
wire n_1732;
wire n_1009;
wire n_1148;
wire n_2051;
wire n_742;
wire n_750;
wire n_2029;
wire n_995;
wire n_454;
wire n_1609;
wire n_374;
wire n_1989;
wire n_396;
wire n_1887;
wire n_1383;
wire n_1073;
wire n_662;
wire n_459;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1920;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1721;
wire n_1959;
wire n_1758;
wire n_1574;
wire n_473;
wire n_2048;
wire n_1921;
wire n_1309;
wire n_1878;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_1800;
wire n_1548;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_743;
wire n_2081;
wire n_613;
wire n_1119;
wire n_1240;
wire n_1820;
wire n_829;
wire n_1612;
wire n_1416;
wire n_2077;
wire n_1724;
wire n_361;
wire n_700;
wire n_1237;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1785;
wire n_1568;
wire n_1006;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_2017;
wire n_2090;
wire n_1870;
wire n_512;
wire n_1591;
wire n_2033;
wire n_1682;
wire n_1980;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1927;
wire n_1349;
wire n_1093;
wire n_1031;
wire n_609;
wire n_1041;
wire n_1265;
wire n_1909;
wire n_1562;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_1965;
wire n_630;
wire n_1902;
wire n_1941;
wire n_1913;
wire n_504;
wire n_1823;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_2015;
wire n_1875;
wire n_1982;
wire n_1304;
wire n_1324;
wire n_987;
wire n_1846;
wire n_2066;
wire n_1885;
wire n_1455;
wire n_767;
wire n_993;
wire n_1903;
wire n_1407;
wire n_1551;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_1805;
wire n_1816;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_1849;
wire n_729;
wire n_1131;
wire n_1084;
wire n_1961;
wire n_970;
wire n_1935;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1534;
wire n_560;
wire n_1354;
wire n_340;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_2088;
wire n_405;
wire n_824;
wire n_359;
wire n_1645;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_1684;
wire n_1717;
wire n_572;
wire n_366;
wire n_815;
wire n_1795;
wire n_1821;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_1708;
wire n_426;
wire n_1438;
wire n_1082;
wire n_1840;
wire n_589;
wire n_1630;
wire n_716;
wire n_562;
wire n_1436;
wire n_1691;
wire n_952;
wire n_1229;
wire n_391;
wire n_1437;
wire n_701;
wire n_1023;
wire n_2075;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_1776;
wire n_531;
wire n_1757;
wire n_890;
wire n_1897;
wire n_764;
wire n_1919;
wire n_1056;
wire n_1424;
wire n_960;
wire n_1893;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_2053;
wire n_634;
wire n_1958;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_1519;
wire n_950;
wire n_1553;
wire n_1811;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1808;
wire n_1060;
wire n_1141;
wire n_389;
wire n_418;
wire n_912;
wire n_968;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_1699;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_1050;
wire n_841;
wire n_802;
wire n_1954;
wire n_1608;
wire n_983;
wire n_1844;
wire n_1305;
wire n_873;
wire n_1826;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_1644;
wire n_690;
wire n_1974;
wire n_583;
wire n_2086;
wire n_1343;
wire n_1203;
wire n_1631;
wire n_821;
wire n_1763;
wire n_1966;
wire n_1768;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1719;
wire n_1288;
wire n_385;
wire n_507;
wire n_1560;
wire n_1605;
wire n_1228;
wire n_972;
wire n_692;
wire n_2037;
wire n_1953;
wire n_1938;
wire n_820;
wire n_1200;
wire n_1911;
wire n_1363;
wire n_1301;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_1967;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_1688;
wire n_945;
wire n_492;
wire n_1504;
wire n_943;
wire n_341;
wire n_992;
wire n_1932;
wire n_543;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_2082;
wire n_1992;
wire n_1643;
wire n_883;
wire n_1983;
wire n_470;
wire n_449;
wire n_1594;
wire n_1400;
wire n_1342;
wire n_1214;
wire n_900;
wire n_856;
wire n_1793;
wire n_1976;
wire n_918;
wire n_942;
wire n_1804;
wire n_1147;
wire n_1557;
wire n_1977;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_356;
wire n_894;
wire n_1636;
wire n_2056;
wire n_1730;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1865;
wire n_1470;
wire n_1096;
wire n_1575;
wire n_1697;
wire n_1735;
wire n_833;
wire n_2020;
wire n_1646;
wire n_1307;
wire n_1881;
wire n_988;
wire n_2043;
wire n_1940;
wire n_814;
wire n_1549;
wire n_1934;
wire n_1201;
wire n_1114;
wire n_655;
wire n_2025;
wire n_1616;
wire n_1446;
wire n_1458;
wire n_472;
wire n_669;
wire n_1176;
wire n_1472;
wire n_1807;
wire n_387;
wire n_1149;
wire n_398;
wire n_1671;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_1824;
wire n_1917;
wire n_1219;
wire n_1204;
wire n_1814;
wire n_1035;
wire n_783;
wire n_555;
wire n_1848;
wire n_1928;
wire n_1188;
wire n_1722;
wire n_661;
wire n_1802;
wire n_849;
wire n_336;
wire n_584;
wire n_681;
wire n_1638;
wire n_1786;
wire n_430;
wire n_2002;
wire n_510;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_2080;
wire n_2068;
wire n_875;
wire n_357;
wire n_1110;
wire n_1655;
wire n_445;
wire n_749;
wire n_1895;
wire n_1134;
wire n_1358;
wire n_717;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_1401;
wire n_969;
wire n_1019;
wire n_1105;
wire n_1998;
wire n_1338;
wire n_577;
wire n_2016;
wire n_1522;
wire n_1687;
wire n_1637;
wire n_2034;
wire n_1419;
wire n_338;
wire n_1653;
wire n_693;
wire n_1506;
wire n_990;
wire n_836;
wire n_1886;
wire n_1389;
wire n_1894;
wire n_975;
wire n_1908;
wire n_1256;
wire n_1702;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_1843;
wire n_1499;
wire n_711;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1929;
wire n_1164;
wire n_1659;
wire n_1834;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_2063;
wire n_1572;
wire n_1968;
wire n_1516;
wire n_876;
wire n_1190;
wire n_1736;
wire n_1685;
wire n_601;
wire n_917;
wire n_1714;
wire n_966;
wire n_1116;
wire n_2000;
wire n_1661;
wire n_1212;
wire n_2074;
wire n_1541;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_1731;
wire n_818;
wire n_1970;
wire n_861;
wire n_1713;
wire n_1183;
wire n_1658;
wire n_899;
wire n_1253;
wire n_1737;
wire n_1904;
wire n_1993;
wire n_774;
wire n_1628;
wire n_1335;
wire n_1514;
wire n_1777;
wire n_1957;
wire n_1059;
wire n_1345;
wire n_1133;
wire n_1771;
wire n_1912;
wire n_1899;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_2067;
wire n_527;
wire n_1168;
wire n_707;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_1584;
wire n_665;
wire n_1726;
wire n_1835;
wire n_1440;
wire n_421;
wire n_1988;
wire n_1853;
wire n_1356;
wire n_1787;
wire n_910;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1774;
wire n_1725;
wire n_1313;
wire n_1136;
wire n_1491;
wire n_754;
wire n_1496;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_1812;
wire n_735;
wire n_1915;
wire n_1109;
wire n_895;
wire n_1310;
wire n_1803;
wire n_427;
wire n_1399;
wire n_1543;
wire n_1991;
wire n_1979;
wire n_791;
wire n_732;
wire n_1533;
wire n_808;
wire n_797;
wire n_1025;
wire n_1930;
wire n_1955;
wire n_500;
wire n_1067;
wire n_1720;
wire n_435;
wire n_2003;
wire n_1457;
wire n_766;
wire n_541;
wire n_538;
wire n_2008;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1742;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_2012;
wire n_594;
wire n_1291;
wire n_1297;
wire n_1753;
wire n_1782;
wire n_1155;
wire n_1418;
wire n_1972;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_985;
wire n_1855;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1703;
wire n_1352;
wire n_626;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_2023;
wire n_676;
wire n_653;
wire n_642;
wire n_1602;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_664;
wire n_1999;
wire n_503;
wire n_2065;
wire n_1372;
wire n_605;
wire n_1273;
wire n_1822;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_980;
wire n_703;
wire n_698;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_1783;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_1907;
wire n_501;
wire n_823;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_1985;
wire n_1898;
wire n_581;
wire n_382;
wire n_554;
wire n_1625;
wire n_898;
wire n_1762;
wire n_1013;
wire n_1452;
wire n_718;
wire n_1120;
wire n_719;
wire n_443;
wire n_1791;
wire n_1890;
wire n_1747;
wire n_714;
wire n_1683;
wire n_1817;
wire n_909;
wire n_1944;
wire n_1497;
wire n_1530;
wire n_997;
wire n_932;
wire n_612;
wire n_2078;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_1981;
wire n_508;
wire n_506;
wire n_1320;
wire n_1663;
wire n_737;
wire n_1718;
wire n_986;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1715;
wire n_1281;
wire n_1952;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_1889;
wire n_1792;
wire n_1564;
wire n_1868;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1922;
wire n_1376;
wire n_941;
wire n_981;
wire n_1569;
wire n_867;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_518;
wire n_505;
wire n_2057;
wire n_1772;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1861;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1901;
wire n_1900;
wire n_1620;
wire n_381;
wire n_390;
wire n_1330;
wire n_1867;
wire n_1945;
wire n_481;
wire n_1675;
wire n_1924;
wire n_1727;
wire n_1554;
wire n_1745;
wire n_769;
wire n_2006;
wire n_1995;
wire n_1046;
wire n_934;
wire n_1618;
wire n_826;
wire n_1813;
wire n_886;
wire n_2014;
wire n_1221;
wire n_654;
wire n_1172;
wire n_379;
wire n_428;
wire n_1341;
wire n_570;
wire n_1641;
wire n_1361;
wire n_1707;
wire n_853;
wire n_377;
wire n_751;
wire n_1973;
wire n_1083;
wire n_786;
wire n_1142;
wire n_1129;
wire n_392;
wire n_704;
wire n_787;
wire n_1770;
wire n_961;
wire n_1756;
wire n_771;
wire n_1716;
wire n_1225;
wire n_1520;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_1873;
wire n_1411;
wire n_622;
wire n_1962;
wire n_1577;
wire n_1087;
wire n_994;
wire n_386;
wire n_1701;
wire n_848;
wire n_1550;
wire n_1498;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1857;
wire n_1344;
wire n_2041;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_1797;
wire n_432;
wire n_1769;
wire n_839;
wire n_1210;
wire n_1364;
wire n_1250;
wire n_369;
wire n_1842;
wire n_871;
wire n_598;
wire n_685;
wire n_608;
wire n_928;
wire n_1367;
wire n_1943;
wire n_1460;
wire n_772;
wire n_2018;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_413;
wire n_402;
wire n_1086;
wire n_796;
wire n_1858;
wire n_1619;
wire n_1502;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_2030;
wire n_903;
wire n_1525;
wire n_1752;
wire n_740;
wire n_384;
wire n_1404;
wire n_1794;
wire n_1315;
wire n_1061;
wire n_1910;
wire n_1298;
wire n_1652;
wire n_462;
wire n_2050;
wire n_1193;
wire n_1676;
wire n_1255;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_844;
wire n_471;
wire n_852;
wire n_1487;
wire n_1864;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_1673;
wire n_465;
wire n_362;
wire n_1321;
wire n_1975;
wire n_2070;
wire n_1937;
wire n_585;
wire n_1739;
wire n_616;
wire n_1914;
wire n_745;
wire n_1654;
wire n_1103;
wire n_648;
wire n_1379;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_1761;
wire n_641;
wire n_730;
wire n_2036;
wire n_1325;
wire n_1595;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_2083;
wire n_695;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_1956;
wire n_1936;
wire n_437;
wire n_1642;
wire n_2027;
wire n_403;
wire n_453;
wire n_1130;
wire n_720;
wire n_1918;
wire n_1526;
wire n_863;
wire n_805;
wire n_1604;
wire n_1275;
wire n_1764;
wire n_712;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_2049;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1741;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_2004;
wire n_1621;
wire n_566;
wire n_565;
wire n_1448;
wire n_1507;
wire n_1398;
wire n_1879;
wire n_597;
wire n_1996;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_2019;
wire n_651;
wire n_1340;
wire n_811;
wire n_1558;
wire n_807;
wire n_835;
wire n_666;
wire n_1433;
wire n_1704;
wire n_1254;
wire n_1026;
wire n_2026;
wire n_1969;
wire n_1234;
wire n_2044;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_2013;
wire n_1990;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_1681;
wire n_2010;
wire n_1018;
wire n_1693;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_1180;
wire n_1827;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_52),
.Y(n_335)
);

BUFx6f_ASAP7_75t_L g336 ( 
.A(n_177),
.Y(n_336)
);

BUFx5_ASAP7_75t_L g337 ( 
.A(n_16),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_245),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_29),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_198),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_154),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_146),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_39),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_312),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_140),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_226),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_317),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_16),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_327),
.Y(n_349)
);

CKINVDCx20_ASAP7_75t_R g350 ( 
.A(n_98),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_315),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_264),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_117),
.Y(n_353)
);

BUFx10_ASAP7_75t_L g354 ( 
.A(n_149),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_67),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_290),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_199),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_34),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_318),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_188),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_330),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_197),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_11),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_273),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_120),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_241),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_52),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_180),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_174),
.Y(n_369)
);

CKINVDCx20_ASAP7_75t_R g370 ( 
.A(n_194),
.Y(n_370)
);

BUFx10_ASAP7_75t_L g371 ( 
.A(n_271),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_148),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_114),
.Y(n_373)
);

INVx2_ASAP7_75t_L g374 ( 
.A(n_239),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_14),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_214),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_235),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_281),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_257),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_323),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_269),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_300),
.Y(n_382)
);

INVx2_ASAP7_75t_L g383 ( 
.A(n_294),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_95),
.Y(n_384)
);

BUFx3_ASAP7_75t_L g385 ( 
.A(n_131),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_238),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_321),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_298),
.Y(n_388)
);

BUFx3_ASAP7_75t_L g389 ( 
.A(n_77),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_320),
.Y(n_390)
);

BUFx6f_ASAP7_75t_L g391 ( 
.A(n_292),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_218),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_297),
.Y(n_393)
);

CKINVDCx14_ASAP7_75t_R g394 ( 
.A(n_149),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_32),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_200),
.Y(n_396)
);

INVx2_ASAP7_75t_L g397 ( 
.A(n_233),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_41),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_19),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_170),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_222),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_68),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_316),
.Y(n_403)
);

CKINVDCx20_ASAP7_75t_R g404 ( 
.A(n_86),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_65),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_119),
.Y(n_406)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_28),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_210),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_63),
.Y(n_409)
);

CKINVDCx20_ASAP7_75t_R g410 ( 
.A(n_250),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_175),
.Y(n_411)
);

BUFx3_ASAP7_75t_L g412 ( 
.A(n_329),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_104),
.Y(n_413)
);

BUFx6f_ASAP7_75t_L g414 ( 
.A(n_304),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_212),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_246),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_128),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_39),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_232),
.Y(n_419)
);

CKINVDCx20_ASAP7_75t_R g420 ( 
.A(n_93),
.Y(n_420)
);

BUFx3_ASAP7_75t_L g421 ( 
.A(n_14),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_221),
.Y(n_422)
);

CKINVDCx14_ASAP7_75t_R g423 ( 
.A(n_128),
.Y(n_423)
);

BUFx2_ASAP7_75t_L g424 ( 
.A(n_256),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_301),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_172),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_331),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_38),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_24),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_27),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_18),
.Y(n_431)
);

INVx1_ASAP7_75t_SL g432 ( 
.A(n_293),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_283),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_91),
.Y(n_434)
);

CKINVDCx20_ASAP7_75t_R g435 ( 
.A(n_117),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_254),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_277),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_247),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_201),
.Y(n_439)
);

CKINVDCx20_ASAP7_75t_R g440 ( 
.A(n_267),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_280),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_203),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_190),
.Y(n_443)
);

INVx2_ASAP7_75t_L g444 ( 
.A(n_70),
.Y(n_444)
);

INVx1_ASAP7_75t_SL g445 ( 
.A(n_325),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_291),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_230),
.Y(n_447)
);

BUFx3_ASAP7_75t_L g448 ( 
.A(n_55),
.Y(n_448)
);

CKINVDCx20_ASAP7_75t_R g449 ( 
.A(n_161),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_207),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_1),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_286),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_74),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_193),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_287),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_146),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_252),
.Y(n_457)
);

BUFx6f_ASAP7_75t_L g458 ( 
.A(n_160),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_248),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_8),
.Y(n_460)
);

BUFx2_ASAP7_75t_L g461 ( 
.A(n_202),
.Y(n_461)
);

CKINVDCx5p33_ASAP7_75t_R g462 ( 
.A(n_249),
.Y(n_462)
);

INVx1_ASAP7_75t_SL g463 ( 
.A(n_79),
.Y(n_463)
);

INVx2_ASAP7_75t_SL g464 ( 
.A(n_124),
.Y(n_464)
);

CKINVDCx20_ASAP7_75t_R g465 ( 
.A(n_272),
.Y(n_465)
);

INVx1_ASAP7_75t_SL g466 ( 
.A(n_84),
.Y(n_466)
);

CKINVDCx5p33_ASAP7_75t_R g467 ( 
.A(n_33),
.Y(n_467)
);

CKINVDCx5p33_ASAP7_75t_R g468 ( 
.A(n_255),
.Y(n_468)
);

CKINVDCx5p33_ASAP7_75t_R g469 ( 
.A(n_289),
.Y(n_469)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_314),
.Y(n_470)
);

BUFx10_ASAP7_75t_L g471 ( 
.A(n_260),
.Y(n_471)
);

INVx2_ASAP7_75t_L g472 ( 
.A(n_206),
.Y(n_472)
);

CKINVDCx5p33_ASAP7_75t_R g473 ( 
.A(n_10),
.Y(n_473)
);

INVx2_ASAP7_75t_SL g474 ( 
.A(n_322),
.Y(n_474)
);

CKINVDCx5p33_ASAP7_75t_R g475 ( 
.A(n_187),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_262),
.Y(n_476)
);

CKINVDCx20_ASAP7_75t_R g477 ( 
.A(n_285),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_296),
.Y(n_478)
);

CKINVDCx16_ASAP7_75t_R g479 ( 
.A(n_47),
.Y(n_479)
);

CKINVDCx5p33_ASAP7_75t_R g480 ( 
.A(n_44),
.Y(n_480)
);

BUFx2_ASAP7_75t_SL g481 ( 
.A(n_179),
.Y(n_481)
);

INVx2_ASAP7_75t_SL g482 ( 
.A(n_110),
.Y(n_482)
);

CKINVDCx5p33_ASAP7_75t_R g483 ( 
.A(n_97),
.Y(n_483)
);

INVx2_ASAP7_75t_L g484 ( 
.A(n_50),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_105),
.Y(n_485)
);

HB1xp67_ASAP7_75t_L g486 ( 
.A(n_85),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_334),
.Y(n_487)
);

CKINVDCx5p33_ASAP7_75t_R g488 ( 
.A(n_9),
.Y(n_488)
);

CKINVDCx16_ASAP7_75t_R g489 ( 
.A(n_196),
.Y(n_489)
);

BUFx6f_ASAP7_75t_L g490 ( 
.A(n_64),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_44),
.Y(n_491)
);

BUFx5_ASAP7_75t_L g492 ( 
.A(n_303),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_54),
.Y(n_493)
);

CKINVDCx5p33_ASAP7_75t_R g494 ( 
.A(n_36),
.Y(n_494)
);

CKINVDCx14_ASAP7_75t_R g495 ( 
.A(n_237),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_328),
.Y(n_496)
);

CKINVDCx20_ASAP7_75t_R g497 ( 
.A(n_282),
.Y(n_497)
);

INVxp67_ASAP7_75t_L g498 ( 
.A(n_49),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_261),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_220),
.Y(n_500)
);

CKINVDCx14_ASAP7_75t_R g501 ( 
.A(n_223),
.Y(n_501)
);

CKINVDCx5p33_ASAP7_75t_R g502 ( 
.A(n_73),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_82),
.Y(n_503)
);

CKINVDCx5p33_ASAP7_75t_R g504 ( 
.A(n_123),
.Y(n_504)
);

CKINVDCx5p33_ASAP7_75t_R g505 ( 
.A(n_69),
.Y(n_505)
);

CKINVDCx5p33_ASAP7_75t_R g506 ( 
.A(n_152),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_26),
.Y(n_507)
);

CKINVDCx5p33_ASAP7_75t_R g508 ( 
.A(n_59),
.Y(n_508)
);

CKINVDCx5p33_ASAP7_75t_R g509 ( 
.A(n_111),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_142),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_219),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_158),
.Y(n_512)
);

CKINVDCx5p33_ASAP7_75t_R g513 ( 
.A(n_15),
.Y(n_513)
);

CKINVDCx5p33_ASAP7_75t_R g514 ( 
.A(n_114),
.Y(n_514)
);

CKINVDCx20_ASAP7_75t_R g515 ( 
.A(n_228),
.Y(n_515)
);

CKINVDCx5p33_ASAP7_75t_R g516 ( 
.A(n_216),
.Y(n_516)
);

INVx2_ASAP7_75t_L g517 ( 
.A(n_104),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_310),
.Y(n_518)
);

CKINVDCx5p33_ASAP7_75t_R g519 ( 
.A(n_263),
.Y(n_519)
);

CKINVDCx5p33_ASAP7_75t_R g520 ( 
.A(n_302),
.Y(n_520)
);

CKINVDCx20_ASAP7_75t_R g521 ( 
.A(n_46),
.Y(n_521)
);

CKINVDCx5p33_ASAP7_75t_R g522 ( 
.A(n_151),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_103),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_109),
.Y(n_524)
);

INVx2_ASAP7_75t_L g525 ( 
.A(n_324),
.Y(n_525)
);

CKINVDCx5p33_ASAP7_75t_R g526 ( 
.A(n_148),
.Y(n_526)
);

CKINVDCx5p33_ASAP7_75t_R g527 ( 
.A(n_22),
.Y(n_527)
);

CKINVDCx5p33_ASAP7_75t_R g528 ( 
.A(n_40),
.Y(n_528)
);

CKINVDCx20_ASAP7_75t_R g529 ( 
.A(n_243),
.Y(n_529)
);

CKINVDCx20_ASAP7_75t_R g530 ( 
.A(n_122),
.Y(n_530)
);

INVx2_ASAP7_75t_L g531 ( 
.A(n_251),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_173),
.Y(n_532)
);

CKINVDCx5p33_ASAP7_75t_R g533 ( 
.A(n_268),
.Y(n_533)
);

CKINVDCx5p33_ASAP7_75t_R g534 ( 
.A(n_213),
.Y(n_534)
);

CKINVDCx20_ASAP7_75t_R g535 ( 
.A(n_234),
.Y(n_535)
);

BUFx10_ASAP7_75t_L g536 ( 
.A(n_99),
.Y(n_536)
);

CKINVDCx5p33_ASAP7_75t_R g537 ( 
.A(n_26),
.Y(n_537)
);

CKINVDCx5p33_ASAP7_75t_R g538 ( 
.A(n_84),
.Y(n_538)
);

CKINVDCx5p33_ASAP7_75t_R g539 ( 
.A(n_37),
.Y(n_539)
);

CKINVDCx5p33_ASAP7_75t_R g540 ( 
.A(n_154),
.Y(n_540)
);

CKINVDCx5p33_ASAP7_75t_R g541 ( 
.A(n_77),
.Y(n_541)
);

BUFx3_ASAP7_75t_L g542 ( 
.A(n_189),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_275),
.Y(n_543)
);

CKINVDCx5p33_ASAP7_75t_R g544 ( 
.A(n_126),
.Y(n_544)
);

INVx2_ASAP7_75t_L g545 ( 
.A(n_313),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_309),
.Y(n_546)
);

BUFx2_ASAP7_75t_L g547 ( 
.A(n_47),
.Y(n_547)
);

CKINVDCx5p33_ASAP7_75t_R g548 ( 
.A(n_122),
.Y(n_548)
);

CKINVDCx5p33_ASAP7_75t_R g549 ( 
.A(n_82),
.Y(n_549)
);

CKINVDCx5p33_ASAP7_75t_R g550 ( 
.A(n_34),
.Y(n_550)
);

CKINVDCx5p33_ASAP7_75t_R g551 ( 
.A(n_100),
.Y(n_551)
);

CKINVDCx5p33_ASAP7_75t_R g552 ( 
.A(n_109),
.Y(n_552)
);

CKINVDCx20_ASAP7_75t_R g553 ( 
.A(n_217),
.Y(n_553)
);

BUFx10_ASAP7_75t_L g554 ( 
.A(n_76),
.Y(n_554)
);

CKINVDCx5p33_ASAP7_75t_R g555 ( 
.A(n_105),
.Y(n_555)
);

CKINVDCx5p33_ASAP7_75t_R g556 ( 
.A(n_191),
.Y(n_556)
);

BUFx2_ASAP7_75t_SL g557 ( 
.A(n_135),
.Y(n_557)
);

CKINVDCx5p33_ASAP7_75t_R g558 ( 
.A(n_42),
.Y(n_558)
);

CKINVDCx5p33_ASAP7_75t_R g559 ( 
.A(n_139),
.Y(n_559)
);

INVxp67_ASAP7_75t_L g560 ( 
.A(n_139),
.Y(n_560)
);

CKINVDCx5p33_ASAP7_75t_R g561 ( 
.A(n_64),
.Y(n_561)
);

CKINVDCx5p33_ASAP7_75t_R g562 ( 
.A(n_71),
.Y(n_562)
);

CKINVDCx5p33_ASAP7_75t_R g563 ( 
.A(n_205),
.Y(n_563)
);

CKINVDCx5p33_ASAP7_75t_R g564 ( 
.A(n_46),
.Y(n_564)
);

CKINVDCx5p33_ASAP7_75t_R g565 ( 
.A(n_66),
.Y(n_565)
);

CKINVDCx20_ASAP7_75t_R g566 ( 
.A(n_83),
.Y(n_566)
);

CKINVDCx5p33_ASAP7_75t_R g567 ( 
.A(n_136),
.Y(n_567)
);

INVx1_ASAP7_75t_SL g568 ( 
.A(n_137),
.Y(n_568)
);

CKINVDCx20_ASAP7_75t_R g569 ( 
.A(n_253),
.Y(n_569)
);

CKINVDCx5p33_ASAP7_75t_R g570 ( 
.A(n_81),
.Y(n_570)
);

CKINVDCx5p33_ASAP7_75t_R g571 ( 
.A(n_288),
.Y(n_571)
);

CKINVDCx20_ASAP7_75t_R g572 ( 
.A(n_306),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_6),
.Y(n_573)
);

CKINVDCx5p33_ASAP7_75t_R g574 ( 
.A(n_94),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_168),
.Y(n_575)
);

CKINVDCx5p33_ASAP7_75t_R g576 ( 
.A(n_178),
.Y(n_576)
);

INVx2_ASAP7_75t_SL g577 ( 
.A(n_259),
.Y(n_577)
);

CKINVDCx5p33_ASAP7_75t_R g578 ( 
.A(n_278),
.Y(n_578)
);

CKINVDCx5p33_ASAP7_75t_R g579 ( 
.A(n_15),
.Y(n_579)
);

CKINVDCx5p33_ASAP7_75t_R g580 ( 
.A(n_2),
.Y(n_580)
);

CKINVDCx16_ASAP7_75t_R g581 ( 
.A(n_231),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_9),
.Y(n_582)
);

CKINVDCx5p33_ASAP7_75t_R g583 ( 
.A(n_17),
.Y(n_583)
);

HB1xp67_ASAP7_75t_L g584 ( 
.A(n_284),
.Y(n_584)
);

CKINVDCx5p33_ASAP7_75t_R g585 ( 
.A(n_295),
.Y(n_585)
);

BUFx2_ASAP7_75t_L g586 ( 
.A(n_332),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_215),
.Y(n_587)
);

CKINVDCx5p33_ASAP7_75t_R g588 ( 
.A(n_92),
.Y(n_588)
);

CKINVDCx5p33_ASAP7_75t_R g589 ( 
.A(n_86),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_76),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_58),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_185),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_96),
.Y(n_593)
);

INVx1_ASAP7_75t_SL g594 ( 
.A(n_102),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_22),
.Y(n_595)
);

CKINVDCx5p33_ASAP7_75t_R g596 ( 
.A(n_120),
.Y(n_596)
);

INVx1_ASAP7_75t_SL g597 ( 
.A(n_244),
.Y(n_597)
);

INVxp67_ASAP7_75t_L g598 ( 
.A(n_87),
.Y(n_598)
);

CKINVDCx16_ASAP7_75t_R g599 ( 
.A(n_85),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_192),
.Y(n_600)
);

CKINVDCx16_ASAP7_75t_R g601 ( 
.A(n_5),
.Y(n_601)
);

CKINVDCx5p33_ASAP7_75t_R g602 ( 
.A(n_305),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_266),
.Y(n_603)
);

CKINVDCx5p33_ASAP7_75t_R g604 ( 
.A(n_3),
.Y(n_604)
);

CKINVDCx5p33_ASAP7_75t_R g605 ( 
.A(n_48),
.Y(n_605)
);

CKINVDCx5p33_ASAP7_75t_R g606 ( 
.A(n_60),
.Y(n_606)
);

CKINVDCx5p33_ASAP7_75t_R g607 ( 
.A(n_151),
.Y(n_607)
);

HB1xp67_ASAP7_75t_L g608 ( 
.A(n_153),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_308),
.Y(n_609)
);

BUFx6f_ASAP7_75t_L g610 ( 
.A(n_227),
.Y(n_610)
);

CKINVDCx5p33_ASAP7_75t_R g611 ( 
.A(n_106),
.Y(n_611)
);

CKINVDCx5p33_ASAP7_75t_R g612 ( 
.A(n_141),
.Y(n_612)
);

CKINVDCx5p33_ASAP7_75t_R g613 ( 
.A(n_72),
.Y(n_613)
);

CKINVDCx20_ASAP7_75t_R g614 ( 
.A(n_258),
.Y(n_614)
);

CKINVDCx5p33_ASAP7_75t_R g615 ( 
.A(n_72),
.Y(n_615)
);

CKINVDCx5p33_ASAP7_75t_R g616 ( 
.A(n_12),
.Y(n_616)
);

CKINVDCx5p33_ASAP7_75t_R g617 ( 
.A(n_155),
.Y(n_617)
);

CKINVDCx5p33_ASAP7_75t_R g618 ( 
.A(n_145),
.Y(n_618)
);

CKINVDCx5p33_ASAP7_75t_R g619 ( 
.A(n_108),
.Y(n_619)
);

BUFx3_ASAP7_75t_L g620 ( 
.A(n_204),
.Y(n_620)
);

INVx2_ASAP7_75t_SL g621 ( 
.A(n_224),
.Y(n_621)
);

INVx1_ASAP7_75t_SL g622 ( 
.A(n_98),
.Y(n_622)
);

CKINVDCx5p33_ASAP7_75t_R g623 ( 
.A(n_31),
.Y(n_623)
);

INVx2_ASAP7_75t_L g624 ( 
.A(n_35),
.Y(n_624)
);

CKINVDCx5p33_ASAP7_75t_R g625 ( 
.A(n_20),
.Y(n_625)
);

CKINVDCx5p33_ASAP7_75t_R g626 ( 
.A(n_30),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_145),
.Y(n_627)
);

CKINVDCx16_ASAP7_75t_R g628 ( 
.A(n_3),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_126),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_61),
.Y(n_630)
);

CKINVDCx5p33_ASAP7_75t_R g631 ( 
.A(n_211),
.Y(n_631)
);

CKINVDCx5p33_ASAP7_75t_R g632 ( 
.A(n_225),
.Y(n_632)
);

CKINVDCx5p33_ASAP7_75t_R g633 ( 
.A(n_1),
.Y(n_633)
);

CKINVDCx5p33_ASAP7_75t_R g634 ( 
.A(n_0),
.Y(n_634)
);

CKINVDCx5p33_ASAP7_75t_R g635 ( 
.A(n_279),
.Y(n_635)
);

CKINVDCx5p33_ASAP7_75t_R g636 ( 
.A(n_12),
.Y(n_636)
);

BUFx2_ASAP7_75t_R g637 ( 
.A(n_229),
.Y(n_637)
);

CKINVDCx5p33_ASAP7_75t_R g638 ( 
.A(n_394),
.Y(n_638)
);

BUFx6f_ASAP7_75t_L g639 ( 
.A(n_336),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_337),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_337),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_337),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_337),
.Y(n_643)
);

INVx1_ASAP7_75t_SL g644 ( 
.A(n_547),
.Y(n_644)
);

INVx2_ASAP7_75t_L g645 ( 
.A(n_337),
.Y(n_645)
);

INVxp67_ASAP7_75t_L g646 ( 
.A(n_486),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_337),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_337),
.Y(n_648)
);

INVxp67_ASAP7_75t_SL g649 ( 
.A(n_584),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_337),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_385),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_385),
.Y(n_652)
);

CKINVDCx20_ASAP7_75t_R g653 ( 
.A(n_350),
.Y(n_653)
);

BUFx2_ASAP7_75t_L g654 ( 
.A(n_423),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_389),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_389),
.Y(n_656)
);

INVxp67_ASAP7_75t_SL g657 ( 
.A(n_424),
.Y(n_657)
);

BUFx3_ASAP7_75t_L g658 ( 
.A(n_412),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_421),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_448),
.Y(n_660)
);

CKINVDCx14_ASAP7_75t_R g661 ( 
.A(n_495),
.Y(n_661)
);

INVxp67_ASAP7_75t_SL g662 ( 
.A(n_461),
.Y(n_662)
);

CKINVDCx14_ASAP7_75t_R g663 ( 
.A(n_501),
.Y(n_663)
);

INVx2_ASAP7_75t_L g664 ( 
.A(n_490),
.Y(n_664)
);

INVx3_ASAP7_75t_L g665 ( 
.A(n_490),
.Y(n_665)
);

CKINVDCx5p33_ASAP7_75t_R g666 ( 
.A(n_388),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_L g667 ( 
.A(n_474),
.B(n_577),
.Y(n_667)
);

INVxp33_ASAP7_75t_SL g668 ( 
.A(n_608),
.Y(n_668)
);

INVxp67_ASAP7_75t_SL g669 ( 
.A(n_586),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_341),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_343),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_365),
.Y(n_672)
);

CKINVDCx20_ASAP7_75t_R g673 ( 
.A(n_404),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_399),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_413),
.Y(n_675)
);

BUFx3_ASAP7_75t_L g676 ( 
.A(n_412),
.Y(n_676)
);

INVxp33_ASAP7_75t_SL g677 ( 
.A(n_335),
.Y(n_677)
);

BUFx2_ASAP7_75t_L g678 ( 
.A(n_335),
.Y(n_678)
);

CKINVDCx5p33_ASAP7_75t_R g679 ( 
.A(n_479),
.Y(n_679)
);

INVxp67_ASAP7_75t_L g680 ( 
.A(n_354),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_485),
.Y(n_681)
);

INVxp33_ASAP7_75t_L g682 ( 
.A(n_407),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_491),
.Y(n_683)
);

CKINVDCx16_ASAP7_75t_R g684 ( 
.A(n_599),
.Y(n_684)
);

CKINVDCx16_ASAP7_75t_R g685 ( 
.A(n_601),
.Y(n_685)
);

INVxp67_ASAP7_75t_L g686 ( 
.A(n_354),
.Y(n_686)
);

INVx2_ASAP7_75t_L g687 ( 
.A(n_492),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_493),
.Y(n_688)
);

INVx3_ASAP7_75t_L g689 ( 
.A(n_407),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_503),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_507),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_510),
.Y(n_692)
);

INVxp67_ASAP7_75t_SL g693 ( 
.A(n_542),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_512),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_523),
.Y(n_695)
);

CKINVDCx20_ASAP7_75t_R g696 ( 
.A(n_420),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_524),
.Y(n_697)
);

INVxp33_ASAP7_75t_L g698 ( 
.A(n_444),
.Y(n_698)
);

CKINVDCx5p33_ASAP7_75t_R g699 ( 
.A(n_393),
.Y(n_699)
);

CKINVDCx5p33_ASAP7_75t_R g700 ( 
.A(n_628),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_573),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_582),
.Y(n_702)
);

INVx1_ASAP7_75t_SL g703 ( 
.A(n_435),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_590),
.Y(n_704)
);

CKINVDCx5p33_ASAP7_75t_R g705 ( 
.A(n_400),
.Y(n_705)
);

CKINVDCx5p33_ASAP7_75t_R g706 ( 
.A(n_395),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_591),
.Y(n_707)
);

CKINVDCx20_ASAP7_75t_R g708 ( 
.A(n_521),
.Y(n_708)
);

CKINVDCx14_ASAP7_75t_R g709 ( 
.A(n_371),
.Y(n_709)
);

INVxp67_ASAP7_75t_SL g710 ( 
.A(n_542),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_593),
.Y(n_711)
);

INVxp67_ASAP7_75t_L g712 ( 
.A(n_354),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_627),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_629),
.Y(n_714)
);

BUFx6f_ASAP7_75t_L g715 ( 
.A(n_336),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_630),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_620),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_620),
.Y(n_718)
);

CKINVDCx5p33_ASAP7_75t_R g719 ( 
.A(n_398),
.Y(n_719)
);

CKINVDCx16_ASAP7_75t_R g720 ( 
.A(n_489),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_346),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_347),
.Y(n_722)
);

INVx4_ASAP7_75t_R g723 ( 
.A(n_474),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_356),
.Y(n_724)
);

CKINVDCx16_ASAP7_75t_R g725 ( 
.A(n_581),
.Y(n_725)
);

BUFx3_ASAP7_75t_L g726 ( 
.A(n_371),
.Y(n_726)
);

CKINVDCx16_ASAP7_75t_R g727 ( 
.A(n_536),
.Y(n_727)
);

CKINVDCx5p33_ASAP7_75t_R g728 ( 
.A(n_402),
.Y(n_728)
);

INVx1_ASAP7_75t_SL g729 ( 
.A(n_530),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_361),
.Y(n_730)
);

INVx2_ASAP7_75t_L g731 ( 
.A(n_492),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_362),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_378),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_379),
.Y(n_734)
);

CKINVDCx20_ASAP7_75t_R g735 ( 
.A(n_566),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_381),
.Y(n_736)
);

INVxp67_ASAP7_75t_SL g737 ( 
.A(n_390),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_392),
.Y(n_738)
);

INVxp33_ASAP7_75t_SL g739 ( 
.A(n_339),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_396),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_401),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_415),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_427),
.Y(n_743)
);

INVxp67_ASAP7_75t_L g744 ( 
.A(n_536),
.Y(n_744)
);

INVxp67_ASAP7_75t_SL g745 ( 
.A(n_437),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_439),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_442),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_446),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_450),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_454),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_457),
.Y(n_751)
);

HB1xp67_ASAP7_75t_L g752 ( 
.A(n_339),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_459),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_476),
.Y(n_754)
);

INVxp67_ASAP7_75t_SL g755 ( 
.A(n_478),
.Y(n_755)
);

INVxp67_ASAP7_75t_SL g756 ( 
.A(n_487),
.Y(n_756)
);

INVxp67_ASAP7_75t_SL g757 ( 
.A(n_496),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_499),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_500),
.Y(n_759)
);

CKINVDCx5p33_ASAP7_75t_R g760 ( 
.A(n_403),
.Y(n_760)
);

CKINVDCx5p33_ASAP7_75t_R g761 ( 
.A(n_405),
.Y(n_761)
);

CKINVDCx5p33_ASAP7_75t_R g762 ( 
.A(n_408),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_511),
.Y(n_763)
);

INVxp67_ASAP7_75t_SL g764 ( 
.A(n_518),
.Y(n_764)
);

CKINVDCx20_ASAP7_75t_R g765 ( 
.A(n_342),
.Y(n_765)
);

INVx2_ASAP7_75t_L g766 ( 
.A(n_492),
.Y(n_766)
);

INVxp33_ASAP7_75t_L g767 ( 
.A(n_444),
.Y(n_767)
);

BUFx6f_ASAP7_75t_L g768 ( 
.A(n_336),
.Y(n_768)
);

INVxp67_ASAP7_75t_SL g769 ( 
.A(n_532),
.Y(n_769)
);

INVxp33_ASAP7_75t_SL g770 ( 
.A(n_342),
.Y(n_770)
);

BUFx3_ASAP7_75t_L g771 ( 
.A(n_371),
.Y(n_771)
);

INVx2_ASAP7_75t_L g772 ( 
.A(n_492),
.Y(n_772)
);

CKINVDCx5p33_ASAP7_75t_R g773 ( 
.A(n_411),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_543),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_546),
.Y(n_775)
);

INVxp33_ASAP7_75t_SL g776 ( 
.A(n_345),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_575),
.Y(n_777)
);

BUFx3_ASAP7_75t_L g778 ( 
.A(n_471),
.Y(n_778)
);

CKINVDCx5p33_ASAP7_75t_R g779 ( 
.A(n_416),
.Y(n_779)
);

BUFx6f_ASAP7_75t_L g780 ( 
.A(n_336),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_587),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_592),
.Y(n_782)
);

CKINVDCx5p33_ASAP7_75t_R g783 ( 
.A(n_419),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_600),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_603),
.Y(n_785)
);

INVxp67_ASAP7_75t_SL g786 ( 
.A(n_609),
.Y(n_786)
);

CKINVDCx20_ASAP7_75t_R g787 ( 
.A(n_345),
.Y(n_787)
);

BUFx3_ASAP7_75t_L g788 ( 
.A(n_471),
.Y(n_788)
);

INVxp67_ASAP7_75t_L g789 ( 
.A(n_536),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_374),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_374),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_383),
.Y(n_792)
);

CKINVDCx20_ASAP7_75t_R g793 ( 
.A(n_348),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_383),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_397),
.Y(n_795)
);

INVxp33_ASAP7_75t_SL g796 ( 
.A(n_348),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_397),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_470),
.Y(n_798)
);

INVxp67_ASAP7_75t_SL g799 ( 
.A(n_470),
.Y(n_799)
);

INVxp67_ASAP7_75t_SL g800 ( 
.A(n_472),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_472),
.Y(n_801)
);

INVxp67_ASAP7_75t_SL g802 ( 
.A(n_525),
.Y(n_802)
);

INVxp67_ASAP7_75t_SL g803 ( 
.A(n_525),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_531),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_545),
.Y(n_805)
);

INVxp67_ASAP7_75t_SL g806 ( 
.A(n_545),
.Y(n_806)
);

CKINVDCx16_ASAP7_75t_R g807 ( 
.A(n_554),
.Y(n_807)
);

INVx2_ASAP7_75t_L g808 ( 
.A(n_492),
.Y(n_808)
);

INVxp33_ASAP7_75t_L g809 ( 
.A(n_484),
.Y(n_809)
);

INVxp67_ASAP7_75t_SL g810 ( 
.A(n_498),
.Y(n_810)
);

CKINVDCx14_ASAP7_75t_R g811 ( 
.A(n_471),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_484),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_517),
.Y(n_813)
);

HB1xp67_ASAP7_75t_L g814 ( 
.A(n_353),
.Y(n_814)
);

INVxp33_ASAP7_75t_SL g815 ( 
.A(n_353),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_595),
.Y(n_816)
);

CKINVDCx20_ASAP7_75t_R g817 ( 
.A(n_355),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_595),
.Y(n_818)
);

CKINVDCx16_ASAP7_75t_R g819 ( 
.A(n_554),
.Y(n_819)
);

CKINVDCx5p33_ASAP7_75t_R g820 ( 
.A(n_422),
.Y(n_820)
);

CKINVDCx16_ASAP7_75t_R g821 ( 
.A(n_554),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_624),
.Y(n_822)
);

INVxp33_ASAP7_75t_SL g823 ( 
.A(n_355),
.Y(n_823)
);

INVxp67_ASAP7_75t_SL g824 ( 
.A(n_560),
.Y(n_824)
);

INVxp33_ASAP7_75t_L g825 ( 
.A(n_336),
.Y(n_825)
);

CKINVDCx20_ASAP7_75t_R g826 ( 
.A(n_358),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_577),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_621),
.Y(n_828)
);

CKINVDCx5p33_ASAP7_75t_R g829 ( 
.A(n_406),
.Y(n_829)
);

CKINVDCx5p33_ASAP7_75t_R g830 ( 
.A(n_409),
.Y(n_830)
);

BUFx2_ASAP7_75t_L g831 ( 
.A(n_358),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_621),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_557),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_464),
.Y(n_834)
);

BUFx3_ASAP7_75t_L g835 ( 
.A(n_338),
.Y(n_835)
);

INVxp33_ASAP7_75t_L g836 ( 
.A(n_391),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_464),
.Y(n_837)
);

INVxp33_ASAP7_75t_L g838 ( 
.A(n_391),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_482),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_482),
.Y(n_840)
);

INVxp33_ASAP7_75t_SL g841 ( 
.A(n_363),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_417),
.Y(n_842)
);

BUFx6f_ASAP7_75t_L g843 ( 
.A(n_391),
.Y(n_843)
);

INVxp67_ASAP7_75t_SL g844 ( 
.A(n_598),
.Y(n_844)
);

INVxp67_ASAP7_75t_L g845 ( 
.A(n_363),
.Y(n_845)
);

INVxp33_ASAP7_75t_SL g846 ( 
.A(n_367),
.Y(n_846)
);

INVx2_ASAP7_75t_L g847 ( 
.A(n_492),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_418),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_428),
.Y(n_849)
);

CKINVDCx5p33_ASAP7_75t_R g850 ( 
.A(n_429),
.Y(n_850)
);

INVxp33_ASAP7_75t_SL g851 ( 
.A(n_367),
.Y(n_851)
);

INVxp67_ASAP7_75t_SL g852 ( 
.A(n_391),
.Y(n_852)
);

INVxp33_ASAP7_75t_L g853 ( 
.A(n_391),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_430),
.Y(n_854)
);

INVxp67_ASAP7_75t_SL g855 ( 
.A(n_414),
.Y(n_855)
);

BUFx5_ASAP7_75t_L g856 ( 
.A(n_492),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_431),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_434),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_451),
.Y(n_859)
);

CKINVDCx14_ASAP7_75t_R g860 ( 
.A(n_338),
.Y(n_860)
);

INVxp33_ASAP7_75t_L g861 ( 
.A(n_414),
.Y(n_861)
);

INVxp67_ASAP7_75t_L g862 ( 
.A(n_372),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_453),
.Y(n_863)
);

CKINVDCx5p33_ASAP7_75t_R g864 ( 
.A(n_456),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_460),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_467),
.Y(n_866)
);

CKINVDCx20_ASAP7_75t_R g867 ( 
.A(n_372),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_473),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_480),
.Y(n_869)
);

BUFx3_ASAP7_75t_L g870 ( 
.A(n_340),
.Y(n_870)
);

INVxp33_ASAP7_75t_SL g871 ( 
.A(n_373),
.Y(n_871)
);

CKINVDCx16_ASAP7_75t_R g872 ( 
.A(n_370),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_483),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_488),
.Y(n_874)
);

INVx1_ASAP7_75t_SL g875 ( 
.A(n_463),
.Y(n_875)
);

CKINVDCx14_ASAP7_75t_R g876 ( 
.A(n_340),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_494),
.Y(n_877)
);

INVx2_ASAP7_75t_L g878 ( 
.A(n_414),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_502),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_504),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_505),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_506),
.Y(n_882)
);

BUFx3_ASAP7_75t_L g883 ( 
.A(n_658),
.Y(n_883)
);

AND2x4_ASAP7_75t_L g884 ( 
.A(n_835),
.B(n_870),
.Y(n_884)
);

BUFx8_ASAP7_75t_L g885 ( 
.A(n_654),
.Y(n_885)
);

INVx2_ASAP7_75t_L g886 ( 
.A(n_664),
.Y(n_886)
);

BUFx6f_ASAP7_75t_L g887 ( 
.A(n_639),
.Y(n_887)
);

BUFx3_ASAP7_75t_L g888 ( 
.A(n_658),
.Y(n_888)
);

INVx4_ASAP7_75t_L g889 ( 
.A(n_666),
.Y(n_889)
);

HB1xp67_ASAP7_75t_L g890 ( 
.A(n_875),
.Y(n_890)
);

AND2x2_ASAP7_75t_L g891 ( 
.A(n_661),
.B(n_432),
.Y(n_891)
);

INVx2_ASAP7_75t_L g892 ( 
.A(n_664),
.Y(n_892)
);

CKINVDCx5p33_ASAP7_75t_R g893 ( 
.A(n_872),
.Y(n_893)
);

BUFx6f_ASAP7_75t_L g894 ( 
.A(n_715),
.Y(n_894)
);

BUFx8_ASAP7_75t_SL g895 ( 
.A(n_653),
.Y(n_895)
);

INVxp67_ASAP7_75t_L g896 ( 
.A(n_752),
.Y(n_896)
);

BUFx2_ASAP7_75t_L g897 ( 
.A(n_679),
.Y(n_897)
);

AND2x2_ASAP7_75t_L g898 ( 
.A(n_661),
.B(n_663),
.Y(n_898)
);

BUFx8_ASAP7_75t_SL g899 ( 
.A(n_653),
.Y(n_899)
);

AND2x4_ASAP7_75t_L g900 ( 
.A(n_835),
.B(n_445),
.Y(n_900)
);

INVxp67_ASAP7_75t_L g901 ( 
.A(n_814),
.Y(n_901)
);

INVx2_ASAP7_75t_L g902 ( 
.A(n_878),
.Y(n_902)
);

OA21x2_ASAP7_75t_L g903 ( 
.A1(n_878),
.A2(n_509),
.B(n_508),
.Y(n_903)
);

AND2x4_ASAP7_75t_L g904 ( 
.A(n_870),
.B(n_597),
.Y(n_904)
);

BUFx6f_ASAP7_75t_L g905 ( 
.A(n_715),
.Y(n_905)
);

AND2x4_ASAP7_75t_L g906 ( 
.A(n_726),
.B(n_344),
.Y(n_906)
);

CKINVDCx5p33_ASAP7_75t_R g907 ( 
.A(n_699),
.Y(n_907)
);

AOI22xp5_ASAP7_75t_L g908 ( 
.A1(n_668),
.A2(n_440),
.B1(n_449),
.B2(n_410),
.Y(n_908)
);

AND2x4_ASAP7_75t_L g909 ( 
.A(n_726),
.B(n_344),
.Y(n_909)
);

INVx2_ASAP7_75t_L g910 ( 
.A(n_665),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_721),
.Y(n_911)
);

HB1xp67_ASAP7_75t_L g912 ( 
.A(n_644),
.Y(n_912)
);

INVx2_ASAP7_75t_L g913 ( 
.A(n_768),
.Y(n_913)
);

BUFx6f_ASAP7_75t_L g914 ( 
.A(n_768),
.Y(n_914)
);

INVx2_ASAP7_75t_L g915 ( 
.A(n_768),
.Y(n_915)
);

INVxp33_ASAP7_75t_SL g916 ( 
.A(n_638),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_L g917 ( 
.A(n_705),
.B(n_425),
.Y(n_917)
);

BUFx12f_ASAP7_75t_L g918 ( 
.A(n_638),
.Y(n_918)
);

NOR2xp33_ASAP7_75t_L g919 ( 
.A(n_667),
.B(n_349),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_L g920 ( 
.A(n_760),
.B(n_426),
.Y(n_920)
);

INVx2_ASAP7_75t_SL g921 ( 
.A(n_706),
.Y(n_921)
);

BUFx6f_ASAP7_75t_L g922 ( 
.A(n_768),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_722),
.Y(n_923)
);

BUFx12f_ASAP7_75t_L g924 ( 
.A(n_679),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_724),
.Y(n_925)
);

BUFx12f_ASAP7_75t_L g926 ( 
.A(n_700),
.Y(n_926)
);

OR2x2_ASAP7_75t_L g927 ( 
.A(n_678),
.B(n_466),
.Y(n_927)
);

OAI21x1_ASAP7_75t_L g928 ( 
.A1(n_645),
.A2(n_641),
.B(n_640),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_730),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_732),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_L g931 ( 
.A(n_762),
.B(n_433),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_733),
.Y(n_932)
);

INVx2_ASAP7_75t_L g933 ( 
.A(n_780),
.Y(n_933)
);

BUFx6f_ASAP7_75t_L g934 ( 
.A(n_843),
.Y(n_934)
);

BUFx2_ASAP7_75t_L g935 ( 
.A(n_700),
.Y(n_935)
);

BUFx8_ASAP7_75t_SL g936 ( 
.A(n_673),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_L g937 ( 
.A(n_773),
.B(n_779),
.Y(n_937)
);

BUFx6f_ASAP7_75t_L g938 ( 
.A(n_843),
.Y(n_938)
);

BUFx8_ASAP7_75t_SL g939 ( 
.A(n_673),
.Y(n_939)
);

CKINVDCx5p33_ASAP7_75t_R g940 ( 
.A(n_783),
.Y(n_940)
);

BUFx6f_ASAP7_75t_L g941 ( 
.A(n_843),
.Y(n_941)
);

AND2x2_ASAP7_75t_L g942 ( 
.A(n_709),
.B(n_351),
.Y(n_942)
);

AOI22xp5_ASAP7_75t_L g943 ( 
.A1(n_668),
.A2(n_477),
.B1(n_497),
.B2(n_465),
.Y(n_943)
);

BUFx6f_ASAP7_75t_L g944 ( 
.A(n_645),
.Y(n_944)
);

BUFx6f_ASAP7_75t_L g945 ( 
.A(n_642),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_L g946 ( 
.A(n_820),
.B(n_436),
.Y(n_946)
);

AOI22x1_ASAP7_75t_SL g947 ( 
.A1(n_696),
.A2(n_375),
.B1(n_384),
.B2(n_373),
.Y(n_947)
);

INVx1_ASAP7_75t_L g948 ( 
.A(n_734),
.Y(n_948)
);

INVx2_ASAP7_75t_L g949 ( 
.A(n_643),
.Y(n_949)
);

INVx2_ASAP7_75t_L g950 ( 
.A(n_647),
.Y(n_950)
);

INVx2_ASAP7_75t_L g951 ( 
.A(n_648),
.Y(n_951)
);

BUFx6f_ASAP7_75t_L g952 ( 
.A(n_650),
.Y(n_952)
);

INVx1_ASAP7_75t_L g953 ( 
.A(n_736),
.Y(n_953)
);

NOR2xp33_ASAP7_75t_L g954 ( 
.A(n_799),
.B(n_351),
.Y(n_954)
);

AND2x4_ASAP7_75t_L g955 ( 
.A(n_771),
.B(n_352),
.Y(n_955)
);

BUFx6f_ASAP7_75t_L g956 ( 
.A(n_812),
.Y(n_956)
);

BUFx6f_ASAP7_75t_L g957 ( 
.A(n_813),
.Y(n_957)
);

INVx6_ASAP7_75t_L g958 ( 
.A(n_676),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_738),
.Y(n_959)
);

BUFx12f_ASAP7_75t_L g960 ( 
.A(n_706),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_740),
.Y(n_961)
);

AND2x2_ASAP7_75t_L g962 ( 
.A(n_709),
.B(n_352),
.Y(n_962)
);

OAI21x1_ASAP7_75t_L g963 ( 
.A1(n_687),
.A2(n_481),
.B(n_441),
.Y(n_963)
);

BUFx6f_ASAP7_75t_L g964 ( 
.A(n_816),
.Y(n_964)
);

BUFx12f_ASAP7_75t_L g965 ( 
.A(n_719),
.Y(n_965)
);

NOR2xp67_ASAP7_75t_L g966 ( 
.A(n_845),
.B(n_357),
.Y(n_966)
);

OAI21x1_ASAP7_75t_L g967 ( 
.A1(n_687),
.A2(n_443),
.B(n_438),
.Y(n_967)
);

HB1xp67_ASAP7_75t_L g968 ( 
.A(n_831),
.Y(n_968)
);

BUFx8_ASAP7_75t_L g969 ( 
.A(n_771),
.Y(n_969)
);

BUFx12f_ASAP7_75t_L g970 ( 
.A(n_719),
.Y(n_970)
);

BUFx6f_ASAP7_75t_L g971 ( 
.A(n_818),
.Y(n_971)
);

INVx2_ASAP7_75t_L g972 ( 
.A(n_790),
.Y(n_972)
);

CKINVDCx20_ASAP7_75t_R g973 ( 
.A(n_696),
.Y(n_973)
);

AND2x4_ASAP7_75t_L g974 ( 
.A(n_778),
.B(n_788),
.Y(n_974)
);

BUFx8_ASAP7_75t_L g975 ( 
.A(n_778),
.Y(n_975)
);

INVx3_ASAP7_75t_L g976 ( 
.A(n_689),
.Y(n_976)
);

BUFx12f_ASAP7_75t_L g977 ( 
.A(n_728),
.Y(n_977)
);

AND2x4_ASAP7_75t_L g978 ( 
.A(n_788),
.B(n_357),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_741),
.Y(n_979)
);

INVx1_ASAP7_75t_L g980 ( 
.A(n_742),
.Y(n_980)
);

HB1xp67_ASAP7_75t_L g981 ( 
.A(n_862),
.Y(n_981)
);

BUFx6f_ASAP7_75t_L g982 ( 
.A(n_822),
.Y(n_982)
);

INVx5_ASAP7_75t_L g983 ( 
.A(n_731),
.Y(n_983)
);

HB1xp67_ASAP7_75t_L g984 ( 
.A(n_676),
.Y(n_984)
);

INVx3_ASAP7_75t_L g985 ( 
.A(n_670),
.Y(n_985)
);

INVx1_ASAP7_75t_L g986 ( 
.A(n_743),
.Y(n_986)
);

INVx1_ASAP7_75t_L g987 ( 
.A(n_746),
.Y(n_987)
);

BUFx6f_ASAP7_75t_L g988 ( 
.A(n_671),
.Y(n_988)
);

OA21x2_ASAP7_75t_L g989 ( 
.A1(n_791),
.A2(n_514),
.B(n_513),
.Y(n_989)
);

INVx2_ASAP7_75t_L g990 ( 
.A(n_792),
.Y(n_990)
);

BUFx3_ASAP7_75t_L g991 ( 
.A(n_717),
.Y(n_991)
);

INVx1_ASAP7_75t_L g992 ( 
.A(n_747),
.Y(n_992)
);

INVx2_ASAP7_75t_L g993 ( 
.A(n_794),
.Y(n_993)
);

AND2x2_ASAP7_75t_L g994 ( 
.A(n_811),
.B(n_359),
.Y(n_994)
);

OAI22x1_ASAP7_75t_L g995 ( 
.A1(n_680),
.A2(n_384),
.B1(n_567),
.B2(n_375),
.Y(n_995)
);

BUFx3_ASAP7_75t_L g996 ( 
.A(n_718),
.Y(n_996)
);

BUFx3_ASAP7_75t_L g997 ( 
.A(n_651),
.Y(n_997)
);

BUFx3_ASAP7_75t_L g998 ( 
.A(n_652),
.Y(n_998)
);

INVx1_ASAP7_75t_L g999 ( 
.A(n_748),
.Y(n_999)
);

BUFx12f_ASAP7_75t_L g1000 ( 
.A(n_728),
.Y(n_1000)
);

INVx1_ASAP7_75t_L g1001 ( 
.A(n_749),
.Y(n_1001)
);

INVx1_ASAP7_75t_L g1002 ( 
.A(n_750),
.Y(n_1002)
);

BUFx8_ASAP7_75t_SL g1003 ( 
.A(n_708),
.Y(n_1003)
);

BUFx8_ASAP7_75t_SL g1004 ( 
.A(n_708),
.Y(n_1004)
);

BUFx8_ASAP7_75t_SL g1005 ( 
.A(n_735),
.Y(n_1005)
);

BUFx6f_ASAP7_75t_L g1006 ( 
.A(n_672),
.Y(n_1006)
);

OAI22xp33_ASAP7_75t_L g1007 ( 
.A1(n_646),
.A2(n_568),
.B1(n_622),
.B2(n_594),
.Y(n_1007)
);

BUFx6f_ASAP7_75t_L g1008 ( 
.A(n_674),
.Y(n_1008)
);

INVx2_ASAP7_75t_L g1009 ( 
.A(n_795),
.Y(n_1009)
);

CKINVDCx5p33_ASAP7_75t_R g1010 ( 
.A(n_720),
.Y(n_1010)
);

HB1xp67_ASAP7_75t_L g1011 ( 
.A(n_761),
.Y(n_1011)
);

BUFx12f_ASAP7_75t_L g1012 ( 
.A(n_761),
.Y(n_1012)
);

INVx2_ASAP7_75t_L g1013 ( 
.A(n_797),
.Y(n_1013)
);

INVx2_ASAP7_75t_L g1014 ( 
.A(n_798),
.Y(n_1014)
);

OAI22x1_ASAP7_75t_SL g1015 ( 
.A1(n_735),
.A2(n_787),
.B1(n_793),
.B2(n_765),
.Y(n_1015)
);

BUFx6f_ASAP7_75t_L g1016 ( 
.A(n_675),
.Y(n_1016)
);

INVx2_ASAP7_75t_L g1017 ( 
.A(n_801),
.Y(n_1017)
);

AND2x2_ASAP7_75t_L g1018 ( 
.A(n_811),
.B(n_359),
.Y(n_1018)
);

BUFx3_ASAP7_75t_L g1019 ( 
.A(n_655),
.Y(n_1019)
);

AND2x4_ASAP7_75t_L g1020 ( 
.A(n_693),
.B(n_360),
.Y(n_1020)
);

AND2x6_ASAP7_75t_L g1021 ( 
.A(n_766),
.B(n_458),
.Y(n_1021)
);

BUFx2_ASAP7_75t_L g1022 ( 
.A(n_765),
.Y(n_1022)
);

BUFx3_ASAP7_75t_L g1023 ( 
.A(n_656),
.Y(n_1023)
);

INVxp67_ASAP7_75t_L g1024 ( 
.A(n_842),
.Y(n_1024)
);

OAI22xp5_ASAP7_75t_L g1025 ( 
.A1(n_657),
.A2(n_570),
.B1(n_574),
.B2(n_567),
.Y(n_1025)
);

OA21x2_ASAP7_75t_L g1026 ( 
.A1(n_804),
.A2(n_526),
.B(n_522),
.Y(n_1026)
);

AND2x4_ASAP7_75t_L g1027 ( 
.A(n_710),
.B(n_360),
.Y(n_1027)
);

INVx1_ASAP7_75t_L g1028 ( 
.A(n_751),
.Y(n_1028)
);

BUFx8_ASAP7_75t_SL g1029 ( 
.A(n_787),
.Y(n_1029)
);

AND2x4_ASAP7_75t_L g1030 ( 
.A(n_848),
.B(n_364),
.Y(n_1030)
);

CKINVDCx20_ASAP7_75t_R g1031 ( 
.A(n_684),
.Y(n_1031)
);

OAI21x1_ASAP7_75t_L g1032 ( 
.A1(n_772),
.A2(n_452),
.B(n_447),
.Y(n_1032)
);

OA21x2_ASAP7_75t_L g1033 ( 
.A1(n_805),
.A2(n_528),
.B(n_527),
.Y(n_1033)
);

INVx1_ASAP7_75t_L g1034 ( 
.A(n_753),
.Y(n_1034)
);

CKINVDCx8_ASAP7_75t_R g1035 ( 
.A(n_685),
.Y(n_1035)
);

AOI22xp5_ASAP7_75t_L g1036 ( 
.A1(n_900),
.A2(n_662),
.B1(n_669),
.B2(n_649),
.Y(n_1036)
);

AND2x4_ASAP7_75t_L g1037 ( 
.A(n_883),
.B(n_827),
.Y(n_1037)
);

INVx2_ASAP7_75t_L g1038 ( 
.A(n_886),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_911),
.Y(n_1039)
);

INVxp67_ASAP7_75t_L g1040 ( 
.A(n_890),
.Y(n_1040)
);

INVx3_ASAP7_75t_L g1041 ( 
.A(n_944),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_923),
.Y(n_1042)
);

INVx3_ASAP7_75t_L g1043 ( 
.A(n_944),
.Y(n_1043)
);

AND2x2_ASAP7_75t_L g1044 ( 
.A(n_890),
.B(n_882),
.Y(n_1044)
);

AND2x4_ASAP7_75t_L g1045 ( 
.A(n_883),
.B(n_828),
.Y(n_1045)
);

INVx2_ASAP7_75t_L g1046 ( 
.A(n_892),
.Y(n_1046)
);

BUFx6f_ASAP7_75t_L g1047 ( 
.A(n_887),
.Y(n_1047)
);

INVx1_ASAP7_75t_L g1048 ( 
.A(n_925),
.Y(n_1048)
);

INVx1_ASAP7_75t_L g1049 ( 
.A(n_929),
.Y(n_1049)
);

HB1xp67_ASAP7_75t_L g1050 ( 
.A(n_912),
.Y(n_1050)
);

INVx1_ASAP7_75t_L g1051 ( 
.A(n_930),
.Y(n_1051)
);

INVx1_ASAP7_75t_L g1052 ( 
.A(n_932),
.Y(n_1052)
);

INVx3_ASAP7_75t_L g1053 ( 
.A(n_944),
.Y(n_1053)
);

AND2x4_ASAP7_75t_L g1054 ( 
.A(n_888),
.B(n_991),
.Y(n_1054)
);

INVx4_ASAP7_75t_L g1055 ( 
.A(n_983),
.Y(n_1055)
);

AND2x4_ASAP7_75t_L g1056 ( 
.A(n_888),
.B(n_832),
.Y(n_1056)
);

INVx1_ASAP7_75t_L g1057 ( 
.A(n_948),
.Y(n_1057)
);

INVxp67_ASAP7_75t_L g1058 ( 
.A(n_912),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_953),
.Y(n_1059)
);

INVx1_ASAP7_75t_L g1060 ( 
.A(n_959),
.Y(n_1060)
);

INVx1_ASAP7_75t_L g1061 ( 
.A(n_961),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_L g1062 ( 
.A(n_919),
.B(n_852),
.Y(n_1062)
);

BUFx3_ASAP7_75t_L g1063 ( 
.A(n_958),
.Y(n_1063)
);

INVx3_ASAP7_75t_L g1064 ( 
.A(n_887),
.Y(n_1064)
);

INVx1_ASAP7_75t_L g1065 ( 
.A(n_979),
.Y(n_1065)
);

NAND2xp5_ASAP7_75t_L g1066 ( 
.A(n_919),
.B(n_1024),
.Y(n_1066)
);

INVxp67_ASAP7_75t_L g1067 ( 
.A(n_984),
.Y(n_1067)
);

INVx1_ASAP7_75t_L g1068 ( 
.A(n_980),
.Y(n_1068)
);

AND2x2_ASAP7_75t_L g1069 ( 
.A(n_991),
.B(n_881),
.Y(n_1069)
);

INVx1_ASAP7_75t_L g1070 ( 
.A(n_986),
.Y(n_1070)
);

AND2x2_ASAP7_75t_L g1071 ( 
.A(n_984),
.B(n_860),
.Y(n_1071)
);

BUFx6f_ASAP7_75t_L g1072 ( 
.A(n_894),
.Y(n_1072)
);

BUFx2_ASAP7_75t_L g1073 ( 
.A(n_1031),
.Y(n_1073)
);

INVx1_ASAP7_75t_L g1074 ( 
.A(n_987),
.Y(n_1074)
);

BUFx3_ASAP7_75t_L g1075 ( 
.A(n_958),
.Y(n_1075)
);

INVx2_ASAP7_75t_L g1076 ( 
.A(n_902),
.Y(n_1076)
);

OAI22xp5_ASAP7_75t_SL g1077 ( 
.A1(n_908),
.A2(n_817),
.B1(n_826),
.B2(n_793),
.Y(n_1077)
);

OA21x2_ASAP7_75t_L g1078 ( 
.A1(n_928),
.A2(n_855),
.B(n_802),
.Y(n_1078)
);

INVx1_ASAP7_75t_L g1079 ( 
.A(n_992),
.Y(n_1079)
);

BUFx3_ASAP7_75t_L g1080 ( 
.A(n_958),
.Y(n_1080)
);

OAI21x1_ASAP7_75t_L g1081 ( 
.A1(n_963),
.A2(n_808),
.B(n_772),
.Y(n_1081)
);

AND2x2_ASAP7_75t_L g1082 ( 
.A(n_996),
.B(n_849),
.Y(n_1082)
);

INVx2_ASAP7_75t_L g1083 ( 
.A(n_902),
.Y(n_1083)
);

INVx2_ASAP7_75t_L g1084 ( 
.A(n_949),
.Y(n_1084)
);

AND2x2_ASAP7_75t_SL g1085 ( 
.A(n_989),
.B(n_458),
.Y(n_1085)
);

AND2x4_ASAP7_75t_L g1086 ( 
.A(n_996),
.B(n_681),
.Y(n_1086)
);

INVxp33_ASAP7_75t_SL g1087 ( 
.A(n_943),
.Y(n_1087)
);

AND2x4_ASAP7_75t_L g1088 ( 
.A(n_884),
.B(n_997),
.Y(n_1088)
);

INVx1_ASAP7_75t_L g1089 ( 
.A(n_999),
.Y(n_1089)
);

INVx2_ASAP7_75t_L g1090 ( 
.A(n_949),
.Y(n_1090)
);

INVx3_ASAP7_75t_L g1091 ( 
.A(n_894),
.Y(n_1091)
);

AND2x2_ASAP7_75t_L g1092 ( 
.A(n_972),
.B(n_854),
.Y(n_1092)
);

AND2x4_ASAP7_75t_L g1093 ( 
.A(n_884),
.B(n_683),
.Y(n_1093)
);

NAND2xp5_ASAP7_75t_L g1094 ( 
.A(n_1024),
.B(n_860),
.Y(n_1094)
);

INVx2_ASAP7_75t_L g1095 ( 
.A(n_950),
.Y(n_1095)
);

AND2x4_ASAP7_75t_L g1096 ( 
.A(n_997),
.B(n_688),
.Y(n_1096)
);

INVx1_ASAP7_75t_L g1097 ( 
.A(n_1001),
.Y(n_1097)
);

INVx1_ASAP7_75t_L g1098 ( 
.A(n_1002),
.Y(n_1098)
);

AND2x6_ASAP7_75t_L g1099 ( 
.A(n_898),
.B(n_458),
.Y(n_1099)
);

INVx2_ASAP7_75t_L g1100 ( 
.A(n_951),
.Y(n_1100)
);

INVx1_ASAP7_75t_L g1101 ( 
.A(n_1028),
.Y(n_1101)
);

NAND2xp5_ASAP7_75t_L g1102 ( 
.A(n_954),
.B(n_876),
.Y(n_1102)
);

INVx1_ASAP7_75t_L g1103 ( 
.A(n_1034),
.Y(n_1103)
);

INVx1_ASAP7_75t_L g1104 ( 
.A(n_951),
.Y(n_1104)
);

NAND2xp5_ASAP7_75t_L g1105 ( 
.A(n_954),
.B(n_876),
.Y(n_1105)
);

OAI21x1_ASAP7_75t_L g1106 ( 
.A1(n_967),
.A2(n_847),
.B(n_808),
.Y(n_1106)
);

INVx1_ASAP7_75t_L g1107 ( 
.A(n_945),
.Y(n_1107)
);

INVx1_ASAP7_75t_L g1108 ( 
.A(n_945),
.Y(n_1108)
);

NAND2xp5_ASAP7_75t_L g1109 ( 
.A(n_1020),
.B(n_737),
.Y(n_1109)
);

AND2x4_ASAP7_75t_L g1110 ( 
.A(n_998),
.B(n_690),
.Y(n_1110)
);

INVx2_ASAP7_75t_L g1111 ( 
.A(n_910),
.Y(n_1111)
);

OAI22xp5_ASAP7_75t_SL g1112 ( 
.A1(n_1031),
.A2(n_826),
.B1(n_867),
.B2(n_817),
.Y(n_1112)
);

INVx1_ASAP7_75t_L g1113 ( 
.A(n_952),
.Y(n_1113)
);

INVx3_ASAP7_75t_L g1114 ( 
.A(n_905),
.Y(n_1114)
);

AND2x2_ASAP7_75t_L g1115 ( 
.A(n_972),
.B(n_880),
.Y(n_1115)
);

INVx2_ASAP7_75t_L g1116 ( 
.A(n_910),
.Y(n_1116)
);

INVx6_ASAP7_75t_L g1117 ( 
.A(n_974),
.Y(n_1117)
);

NAND2xp5_ASAP7_75t_L g1118 ( 
.A(n_1020),
.B(n_1027),
.Y(n_1118)
);

INVx2_ASAP7_75t_L g1119 ( 
.A(n_913),
.Y(n_1119)
);

INVx1_ASAP7_75t_L g1120 ( 
.A(n_998),
.Y(n_1120)
);

NAND2xp5_ASAP7_75t_L g1121 ( 
.A(n_1027),
.B(n_745),
.Y(n_1121)
);

NOR2xp33_ASAP7_75t_L g1122 ( 
.A(n_981),
.B(n_677),
.Y(n_1122)
);

INVx1_ASAP7_75t_L g1123 ( 
.A(n_1019),
.Y(n_1123)
);

BUFx6f_ASAP7_75t_L g1124 ( 
.A(n_905),
.Y(n_1124)
);

INVx1_ASAP7_75t_L g1125 ( 
.A(n_1019),
.Y(n_1125)
);

INVx1_ASAP7_75t_L g1126 ( 
.A(n_1023),
.Y(n_1126)
);

AND2x2_ASAP7_75t_L g1127 ( 
.A(n_990),
.B(n_879),
.Y(n_1127)
);

INVx1_ASAP7_75t_L g1128 ( 
.A(n_1023),
.Y(n_1128)
);

INVx2_ASAP7_75t_L g1129 ( 
.A(n_915),
.Y(n_1129)
);

AND2x4_ASAP7_75t_L g1130 ( 
.A(n_985),
.B(n_691),
.Y(n_1130)
);

INVx1_ASAP7_75t_L g1131 ( 
.A(n_988),
.Y(n_1131)
);

INVx1_ASAP7_75t_L g1132 ( 
.A(n_988),
.Y(n_1132)
);

INVxp67_ASAP7_75t_L g1133 ( 
.A(n_927),
.Y(n_1133)
);

HB1xp67_ASAP7_75t_L g1134 ( 
.A(n_968),
.Y(n_1134)
);

INVx3_ASAP7_75t_L g1135 ( 
.A(n_905),
.Y(n_1135)
);

OA21x2_ASAP7_75t_L g1136 ( 
.A1(n_1032),
.A2(n_803),
.B(n_800),
.Y(n_1136)
);

INVx3_ASAP7_75t_L g1137 ( 
.A(n_905),
.Y(n_1137)
);

INVx1_ASAP7_75t_L g1138 ( 
.A(n_1006),
.Y(n_1138)
);

INVx2_ASAP7_75t_L g1139 ( 
.A(n_933),
.Y(n_1139)
);

NAND2xp5_ASAP7_75t_L g1140 ( 
.A(n_917),
.B(n_920),
.Y(n_1140)
);

INVx2_ASAP7_75t_L g1141 ( 
.A(n_933),
.Y(n_1141)
);

XNOR2xp5_ASAP7_75t_L g1142 ( 
.A(n_973),
.B(n_703),
.Y(n_1142)
);

INVx3_ASAP7_75t_L g1143 ( 
.A(n_914),
.Y(n_1143)
);

AND2x4_ASAP7_75t_L g1144 ( 
.A(n_985),
.B(n_692),
.Y(n_1144)
);

INVx1_ASAP7_75t_L g1145 ( 
.A(n_1008),
.Y(n_1145)
);

BUFx2_ASAP7_75t_L g1146 ( 
.A(n_893),
.Y(n_1146)
);

INVx1_ASAP7_75t_L g1147 ( 
.A(n_1008),
.Y(n_1147)
);

NAND2xp5_ASAP7_75t_L g1148 ( 
.A(n_931),
.B(n_755),
.Y(n_1148)
);

INVx1_ASAP7_75t_L g1149 ( 
.A(n_1008),
.Y(n_1149)
);

BUFx6f_ASAP7_75t_L g1150 ( 
.A(n_914),
.Y(n_1150)
);

AND2x2_ASAP7_75t_L g1151 ( 
.A(n_993),
.B(n_857),
.Y(n_1151)
);

AND2x2_ASAP7_75t_L g1152 ( 
.A(n_981),
.B(n_725),
.Y(n_1152)
);

INVx1_ASAP7_75t_L g1153 ( 
.A(n_1016),
.Y(n_1153)
);

AND2x2_ASAP7_75t_L g1154 ( 
.A(n_891),
.B(n_829),
.Y(n_1154)
);

INVx3_ASAP7_75t_L g1155 ( 
.A(n_922),
.Y(n_1155)
);

BUFx6f_ASAP7_75t_L g1156 ( 
.A(n_922),
.Y(n_1156)
);

INVx3_ASAP7_75t_L g1157 ( 
.A(n_922),
.Y(n_1157)
);

AND2x2_ASAP7_75t_L g1158 ( 
.A(n_1050),
.B(n_974),
.Y(n_1158)
);

INVx2_ASAP7_75t_SL g1159 ( 
.A(n_1050),
.Y(n_1159)
);

NOR2xp33_ASAP7_75t_L g1160 ( 
.A(n_1066),
.B(n_937),
.Y(n_1160)
);

AOI22xp33_ASAP7_75t_L g1161 ( 
.A1(n_1085),
.A2(n_1026),
.B1(n_1033),
.B2(n_989),
.Y(n_1161)
);

BUFx10_ASAP7_75t_L g1162 ( 
.A(n_1122),
.Y(n_1162)
);

INVx4_ASAP7_75t_L g1163 ( 
.A(n_1117),
.Y(n_1163)
);

OR2x6_ASAP7_75t_L g1164 ( 
.A(n_1146),
.B(n_924),
.Y(n_1164)
);

NAND2xp5_ASAP7_75t_L g1165 ( 
.A(n_1062),
.B(n_900),
.Y(n_1165)
);

NAND2xp5_ASAP7_75t_L g1166 ( 
.A(n_1140),
.B(n_1148),
.Y(n_1166)
);

INVx2_ASAP7_75t_L g1167 ( 
.A(n_1038),
.Y(n_1167)
);

NAND2xp5_ASAP7_75t_SL g1168 ( 
.A(n_1085),
.B(n_904),
.Y(n_1168)
);

BUFx6f_ASAP7_75t_L g1169 ( 
.A(n_1063),
.Y(n_1169)
);

INVx1_ASAP7_75t_L g1170 ( 
.A(n_1039),
.Y(n_1170)
);

BUFx10_ASAP7_75t_L g1171 ( 
.A(n_1122),
.Y(n_1171)
);

NAND2xp5_ASAP7_75t_L g1172 ( 
.A(n_1109),
.B(n_904),
.Y(n_1172)
);

NOR2xp33_ASAP7_75t_L g1173 ( 
.A(n_1067),
.B(n_889),
.Y(n_1173)
);

INVx1_ASAP7_75t_L g1174 ( 
.A(n_1042),
.Y(n_1174)
);

INVx2_ASAP7_75t_L g1175 ( 
.A(n_1046),
.Y(n_1175)
);

NAND2xp5_ASAP7_75t_SL g1176 ( 
.A(n_1118),
.B(n_921),
.Y(n_1176)
);

NAND2xp5_ASAP7_75t_SL g1177 ( 
.A(n_1121),
.B(n_940),
.Y(n_1177)
);

OAI22xp33_ASAP7_75t_SL g1178 ( 
.A1(n_1087),
.A2(n_739),
.B1(n_770),
.B2(n_677),
.Y(n_1178)
);

OR2x2_ASAP7_75t_L g1179 ( 
.A(n_1133),
.B(n_729),
.Y(n_1179)
);

NOR2xp33_ASAP7_75t_L g1180 ( 
.A(n_1102),
.B(n_889),
.Y(n_1180)
);

INVx6_ASAP7_75t_L g1181 ( 
.A(n_1117),
.Y(n_1181)
);

BUFx2_ASAP7_75t_L g1182 ( 
.A(n_1058),
.Y(n_1182)
);

NAND2xp5_ASAP7_75t_SL g1183 ( 
.A(n_1105),
.B(n_940),
.Y(n_1183)
);

INVx2_ASAP7_75t_SL g1184 ( 
.A(n_1093),
.Y(n_1184)
);

NAND2xp5_ASAP7_75t_L g1185 ( 
.A(n_1048),
.B(n_946),
.Y(n_1185)
);

AOI22xp33_ASAP7_75t_L g1186 ( 
.A1(n_1078),
.A2(n_1026),
.B1(n_1033),
.B2(n_989),
.Y(n_1186)
);

INVxp67_ASAP7_75t_L g1187 ( 
.A(n_1044),
.Y(n_1187)
);

BUFx3_ASAP7_75t_L g1188 ( 
.A(n_1075),
.Y(n_1188)
);

NAND2xp5_ASAP7_75t_L g1189 ( 
.A(n_1049),
.B(n_1051),
.Y(n_1189)
);

NAND2xp5_ASAP7_75t_L g1190 ( 
.A(n_1052),
.B(n_903),
.Y(n_1190)
);

NOR3xp33_ASAP7_75t_L g1191 ( 
.A(n_1094),
.B(n_1007),
.C(n_901),
.Y(n_1191)
);

INVx1_ASAP7_75t_L g1192 ( 
.A(n_1057),
.Y(n_1192)
);

BUFx2_ASAP7_75t_L g1193 ( 
.A(n_1040),
.Y(n_1193)
);

INVx3_ASAP7_75t_L g1194 ( 
.A(n_1119),
.Y(n_1194)
);

CKINVDCx6p67_ASAP7_75t_R g1195 ( 
.A(n_1073),
.Y(n_1195)
);

BUFx3_ASAP7_75t_L g1196 ( 
.A(n_1075),
.Y(n_1196)
);

AND3x2_ASAP7_75t_L g1197 ( 
.A(n_1134),
.B(n_1011),
.C(n_935),
.Y(n_1197)
);

INVx1_ASAP7_75t_L g1198 ( 
.A(n_1059),
.Y(n_1198)
);

INVx1_ASAP7_75t_L g1199 ( 
.A(n_1060),
.Y(n_1199)
);

BUFx6f_ASAP7_75t_SL g1200 ( 
.A(n_1093),
.Y(n_1200)
);

AOI22xp33_ASAP7_75t_L g1201 ( 
.A1(n_1078),
.A2(n_1033),
.B1(n_1026),
.B2(n_903),
.Y(n_1201)
);

AND2x2_ASAP7_75t_L g1202 ( 
.A(n_1044),
.B(n_942),
.Y(n_1202)
);

CKINVDCx5p33_ASAP7_75t_R g1203 ( 
.A(n_1142),
.Y(n_1203)
);

INVx1_ASAP7_75t_L g1204 ( 
.A(n_1061),
.Y(n_1204)
);

NAND2x1p5_ASAP7_75t_L g1205 ( 
.A(n_1088),
.B(n_903),
.Y(n_1205)
);

AND2x2_ASAP7_75t_L g1206 ( 
.A(n_1154),
.B(n_962),
.Y(n_1206)
);

NAND2xp5_ASAP7_75t_SL g1207 ( 
.A(n_1088),
.B(n_907),
.Y(n_1207)
);

INVx1_ASAP7_75t_L g1208 ( 
.A(n_1065),
.Y(n_1208)
);

CKINVDCx20_ASAP7_75t_R g1209 ( 
.A(n_1112),
.Y(n_1209)
);

BUFx2_ASAP7_75t_L g1210 ( 
.A(n_1134),
.Y(n_1210)
);

NAND3xp33_ASAP7_75t_SL g1211 ( 
.A(n_1036),
.B(n_867),
.C(n_830),
.Y(n_1211)
);

INVx1_ASAP7_75t_L g1212 ( 
.A(n_1068),
.Y(n_1212)
);

NAND2xp5_ASAP7_75t_SL g1213 ( 
.A(n_1088),
.B(n_966),
.Y(n_1213)
);

INVx2_ASAP7_75t_L g1214 ( 
.A(n_1076),
.Y(n_1214)
);

NOR2xp33_ASAP7_75t_L g1215 ( 
.A(n_1070),
.B(n_896),
.Y(n_1215)
);

OAI22xp33_ASAP7_75t_L g1216 ( 
.A1(n_1087),
.A2(n_698),
.B1(n_767),
.B2(n_682),
.Y(n_1216)
);

NOR2xp33_ASAP7_75t_L g1217 ( 
.A(n_1074),
.B(n_896),
.Y(n_1217)
);

INVx1_ASAP7_75t_L g1218 ( 
.A(n_1079),
.Y(n_1218)
);

NAND2xp5_ASAP7_75t_L g1219 ( 
.A(n_1089),
.B(n_994),
.Y(n_1219)
);

AO22x2_ASAP7_75t_L g1220 ( 
.A1(n_1152),
.A2(n_947),
.B1(n_1025),
.B2(n_901),
.Y(n_1220)
);

INVx2_ASAP7_75t_L g1221 ( 
.A(n_1083),
.Y(n_1221)
);

INVx2_ASAP7_75t_L g1222 ( 
.A(n_1111),
.Y(n_1222)
);

NAND2xp33_ASAP7_75t_SL g1223 ( 
.A(n_1071),
.B(n_515),
.Y(n_1223)
);

INVx2_ASAP7_75t_L g1224 ( 
.A(n_1111),
.Y(n_1224)
);

BUFx4f_ASAP7_75t_L g1225 ( 
.A(n_1117),
.Y(n_1225)
);

INVx1_ASAP7_75t_L g1226 ( 
.A(n_1097),
.Y(n_1226)
);

INVx2_ASAP7_75t_L g1227 ( 
.A(n_1116),
.Y(n_1227)
);

NAND2xp5_ASAP7_75t_L g1228 ( 
.A(n_1098),
.B(n_1018),
.Y(n_1228)
);

NAND2xp5_ASAP7_75t_SL g1229 ( 
.A(n_1054),
.B(n_1011),
.Y(n_1229)
);

INVx1_ASAP7_75t_L g1230 ( 
.A(n_1101),
.Y(n_1230)
);

INVx2_ASAP7_75t_L g1231 ( 
.A(n_1116),
.Y(n_1231)
);

AND2x4_ASAP7_75t_L g1232 ( 
.A(n_1080),
.B(n_1054),
.Y(n_1232)
);

AOI22xp33_ASAP7_75t_L g1233 ( 
.A1(n_1078),
.A2(n_1007),
.B1(n_806),
.B2(n_682),
.Y(n_1233)
);

INVxp67_ASAP7_75t_SL g1234 ( 
.A(n_1092),
.Y(n_1234)
);

INVx2_ASAP7_75t_L g1235 ( 
.A(n_1084),
.Y(n_1235)
);

INVx2_ASAP7_75t_L g1236 ( 
.A(n_1090),
.Y(n_1236)
);

INVx2_ASAP7_75t_L g1237 ( 
.A(n_1090),
.Y(n_1237)
);

INVx2_ASAP7_75t_L g1238 ( 
.A(n_1095),
.Y(n_1238)
);

INVx4_ASAP7_75t_L g1239 ( 
.A(n_1080),
.Y(n_1239)
);

INVx1_ASAP7_75t_L g1240 ( 
.A(n_1103),
.Y(n_1240)
);

INVx5_ASAP7_75t_L g1241 ( 
.A(n_1055),
.Y(n_1241)
);

NOR2xp33_ASAP7_75t_L g1242 ( 
.A(n_1069),
.B(n_1030),
.Y(n_1242)
);

NOR2xp33_ASAP7_75t_L g1243 ( 
.A(n_1069),
.B(n_1030),
.Y(n_1243)
);

INVx2_ASAP7_75t_L g1244 ( 
.A(n_1095),
.Y(n_1244)
);

INVx4_ASAP7_75t_L g1245 ( 
.A(n_1054),
.Y(n_1245)
);

INVx2_ASAP7_75t_SL g1246 ( 
.A(n_1037),
.Y(n_1246)
);

NAND3xp33_ASAP7_75t_L g1247 ( 
.A(n_1082),
.B(n_830),
.C(n_829),
.Y(n_1247)
);

OAI22xp33_ASAP7_75t_SL g1248 ( 
.A1(n_1120),
.A2(n_739),
.B1(n_776),
.B2(n_770),
.Y(n_1248)
);

INVx2_ASAP7_75t_SL g1249 ( 
.A(n_1037),
.Y(n_1249)
);

OAI22xp5_ASAP7_75t_L g1250 ( 
.A1(n_1123),
.A2(n_535),
.B1(n_553),
.B2(n_529),
.Y(n_1250)
);

NOR2xp33_ASAP7_75t_R g1251 ( 
.A(n_1125),
.B(n_893),
.Y(n_1251)
);

INVx4_ASAP7_75t_L g1252 ( 
.A(n_1037),
.Y(n_1252)
);

INVx4_ASAP7_75t_L g1253 ( 
.A(n_1045),
.Y(n_1253)
);

OAI22xp33_ASAP7_75t_L g1254 ( 
.A1(n_1126),
.A2(n_767),
.B1(n_809),
.B2(n_698),
.Y(n_1254)
);

INVx6_ASAP7_75t_L g1255 ( 
.A(n_1045),
.Y(n_1255)
);

NAND2xp5_ASAP7_75t_L g1256 ( 
.A(n_1092),
.B(n_906),
.Y(n_1256)
);

CKINVDCx5p33_ASAP7_75t_R g1257 ( 
.A(n_1077),
.Y(n_1257)
);

NAND2xp5_ASAP7_75t_L g1258 ( 
.A(n_1115),
.B(n_906),
.Y(n_1258)
);

AO22x2_ASAP7_75t_L g1259 ( 
.A1(n_1082),
.A2(n_712),
.B1(n_744),
.B2(n_686),
.Y(n_1259)
);

AND3x2_ASAP7_75t_L g1260 ( 
.A(n_1045),
.B(n_897),
.C(n_968),
.Y(n_1260)
);

NAND2xp5_ASAP7_75t_L g1261 ( 
.A(n_1115),
.B(n_909),
.Y(n_1261)
);

NAND2xp5_ASAP7_75t_L g1262 ( 
.A(n_1127),
.B(n_909),
.Y(n_1262)
);

BUFx3_ASAP7_75t_L g1263 ( 
.A(n_1056),
.Y(n_1263)
);

INVx2_ASAP7_75t_L g1264 ( 
.A(n_1100),
.Y(n_1264)
);

INVx2_ASAP7_75t_L g1265 ( 
.A(n_1129),
.Y(n_1265)
);

NOR2xp33_ASAP7_75t_L g1266 ( 
.A(n_1128),
.B(n_776),
.Y(n_1266)
);

NOR2xp33_ASAP7_75t_L g1267 ( 
.A(n_1127),
.B(n_796),
.Y(n_1267)
);

INVx1_ASAP7_75t_L g1268 ( 
.A(n_1151),
.Y(n_1268)
);

INVx1_ASAP7_75t_L g1269 ( 
.A(n_1151),
.Y(n_1269)
);

NOR2xp33_ASAP7_75t_L g1270 ( 
.A(n_1086),
.B(n_796),
.Y(n_1270)
);

BUFx10_ASAP7_75t_L g1271 ( 
.A(n_1086),
.Y(n_1271)
);

INVx1_ASAP7_75t_L g1272 ( 
.A(n_1096),
.Y(n_1272)
);

INVx2_ASAP7_75t_L g1273 ( 
.A(n_1139),
.Y(n_1273)
);

INVx1_ASAP7_75t_L g1274 ( 
.A(n_1096),
.Y(n_1274)
);

INVx1_ASAP7_75t_L g1275 ( 
.A(n_1096),
.Y(n_1275)
);

AND2x4_ASAP7_75t_L g1276 ( 
.A(n_1110),
.B(n_955),
.Y(n_1276)
);

INVx1_ASAP7_75t_L g1277 ( 
.A(n_1110),
.Y(n_1277)
);

INVxp67_ASAP7_75t_SL g1278 ( 
.A(n_1047),
.Y(n_1278)
);

INVx1_ASAP7_75t_L g1279 ( 
.A(n_1110),
.Y(n_1279)
);

INVx1_ASAP7_75t_L g1280 ( 
.A(n_1130),
.Y(n_1280)
);

BUFx6f_ASAP7_75t_L g1281 ( 
.A(n_1047),
.Y(n_1281)
);

INVx1_ASAP7_75t_L g1282 ( 
.A(n_1130),
.Y(n_1282)
);

INVx1_ASAP7_75t_L g1283 ( 
.A(n_1130),
.Y(n_1283)
);

INVx1_ASAP7_75t_L g1284 ( 
.A(n_1144),
.Y(n_1284)
);

INVx1_ASAP7_75t_SL g1285 ( 
.A(n_1144),
.Y(n_1285)
);

AND2x2_ASAP7_75t_L g1286 ( 
.A(n_1187),
.B(n_955),
.Y(n_1286)
);

BUFx3_ASAP7_75t_L g1287 ( 
.A(n_1188),
.Y(n_1287)
);

NAND2xp5_ASAP7_75t_SL g1288 ( 
.A(n_1166),
.B(n_1145),
.Y(n_1288)
);

NAND2xp5_ASAP7_75t_SL g1289 ( 
.A(n_1160),
.B(n_1147),
.Y(n_1289)
);

NAND2xp5_ASAP7_75t_SL g1290 ( 
.A(n_1160),
.B(n_1149),
.Y(n_1290)
);

BUFx2_ASAP7_75t_L g1291 ( 
.A(n_1210),
.Y(n_1291)
);

AND2x4_ASAP7_75t_L g1292 ( 
.A(n_1188),
.B(n_1196),
.Y(n_1292)
);

INVx2_ASAP7_75t_L g1293 ( 
.A(n_1224),
.Y(n_1293)
);

CKINVDCx5p33_ASAP7_75t_R g1294 ( 
.A(n_1203),
.Y(n_1294)
);

INVx3_ASAP7_75t_L g1295 ( 
.A(n_1245),
.Y(n_1295)
);

BUFx2_ASAP7_75t_L g1296 ( 
.A(n_1159),
.Y(n_1296)
);

INVx1_ASAP7_75t_L g1297 ( 
.A(n_1235),
.Y(n_1297)
);

INVx1_ASAP7_75t_L g1298 ( 
.A(n_1236),
.Y(n_1298)
);

AND2x4_ASAP7_75t_L g1299 ( 
.A(n_1196),
.B(n_1144),
.Y(n_1299)
);

NOR2xp33_ASAP7_75t_L g1300 ( 
.A(n_1187),
.B(n_916),
.Y(n_1300)
);

BUFx6f_ASAP7_75t_L g1301 ( 
.A(n_1169),
.Y(n_1301)
);

INVx5_ASAP7_75t_L g1302 ( 
.A(n_1281),
.Y(n_1302)
);

INVx3_ASAP7_75t_L g1303 ( 
.A(n_1232),
.Y(n_1303)
);

BUFx6f_ASAP7_75t_L g1304 ( 
.A(n_1169),
.Y(n_1304)
);

AOI22xp33_ASAP7_75t_L g1305 ( 
.A1(n_1168),
.A2(n_824),
.B1(n_844),
.B2(n_810),
.Y(n_1305)
);

NOR2xp33_ASAP7_75t_L g1306 ( 
.A(n_1165),
.B(n_916),
.Y(n_1306)
);

HB1xp67_ASAP7_75t_L g1307 ( 
.A(n_1234),
.Y(n_1307)
);

INVx1_ASAP7_75t_L g1308 ( 
.A(n_1237),
.Y(n_1308)
);

NAND2x1p5_ASAP7_75t_L g1309 ( 
.A(n_1163),
.B(n_1225),
.Y(n_1309)
);

AND2x4_ASAP7_75t_SL g1310 ( 
.A(n_1271),
.B(n_973),
.Y(n_1310)
);

INVx2_ASAP7_75t_L g1311 ( 
.A(n_1224),
.Y(n_1311)
);

NAND2xp5_ASAP7_75t_L g1312 ( 
.A(n_1234),
.B(n_1104),
.Y(n_1312)
);

INVx2_ASAP7_75t_L g1313 ( 
.A(n_1227),
.Y(n_1313)
);

NAND2xp33_ASAP7_75t_L g1314 ( 
.A(n_1168),
.B(n_1099),
.Y(n_1314)
);

NOR2xp33_ASAP7_75t_SL g1315 ( 
.A(n_1225),
.B(n_637),
.Y(n_1315)
);

INVx8_ASAP7_75t_L g1316 ( 
.A(n_1200),
.Y(n_1316)
);

BUFx2_ASAP7_75t_L g1317 ( 
.A(n_1158),
.Y(n_1317)
);

INVx1_ASAP7_75t_L g1318 ( 
.A(n_1238),
.Y(n_1318)
);

INVx4_ASAP7_75t_L g1319 ( 
.A(n_1169),
.Y(n_1319)
);

AND2x4_ASAP7_75t_L g1320 ( 
.A(n_1232),
.B(n_978),
.Y(n_1320)
);

NOR2x1p5_ASAP7_75t_L g1321 ( 
.A(n_1195),
.B(n_918),
.Y(n_1321)
);

INVx1_ASAP7_75t_SL g1322 ( 
.A(n_1182),
.Y(n_1322)
);

INVx1_ASAP7_75t_L g1323 ( 
.A(n_1244),
.Y(n_1323)
);

INVx1_ASAP7_75t_L g1324 ( 
.A(n_1244),
.Y(n_1324)
);

INVx2_ASAP7_75t_L g1325 ( 
.A(n_1227),
.Y(n_1325)
);

AND2x4_ASAP7_75t_L g1326 ( 
.A(n_1263),
.B(n_978),
.Y(n_1326)
);

INVx2_ASAP7_75t_L g1327 ( 
.A(n_1231),
.Y(n_1327)
);

NAND2xp5_ASAP7_75t_L g1328 ( 
.A(n_1172),
.B(n_1041),
.Y(n_1328)
);

INVx2_ASAP7_75t_L g1329 ( 
.A(n_1231),
.Y(n_1329)
);

BUFx4f_ASAP7_75t_L g1330 ( 
.A(n_1164),
.Y(n_1330)
);

INVx3_ASAP7_75t_L g1331 ( 
.A(n_1252),
.Y(n_1331)
);

NOR2xp33_ASAP7_75t_L g1332 ( 
.A(n_1267),
.B(n_815),
.Y(n_1332)
);

AND2x4_ASAP7_75t_L g1333 ( 
.A(n_1263),
.B(n_1131),
.Y(n_1333)
);

INVx2_ASAP7_75t_L g1334 ( 
.A(n_1167),
.Y(n_1334)
);

OR2x6_ASAP7_75t_L g1335 ( 
.A(n_1164),
.B(n_1022),
.Y(n_1335)
);

XOR2xp5_ASAP7_75t_L g1336 ( 
.A(n_1247),
.B(n_1015),
.Y(n_1336)
);

AND2x4_ASAP7_75t_L g1337 ( 
.A(n_1184),
.B(n_1132),
.Y(n_1337)
);

BUFx3_ASAP7_75t_L g1338 ( 
.A(n_1193),
.Y(n_1338)
);

INVx2_ASAP7_75t_L g1339 ( 
.A(n_1175),
.Y(n_1339)
);

NOR2xp33_ASAP7_75t_L g1340 ( 
.A(n_1267),
.B(n_815),
.Y(n_1340)
);

AOI22x1_ASAP7_75t_L g1341 ( 
.A1(n_1205),
.A2(n_995),
.B1(n_1141),
.B2(n_1107),
.Y(n_1341)
);

INVx1_ASAP7_75t_SL g1342 ( 
.A(n_1179),
.Y(n_1342)
);

CKINVDCx8_ASAP7_75t_R g1343 ( 
.A(n_1164),
.Y(n_1343)
);

NAND2xp5_ASAP7_75t_L g1344 ( 
.A(n_1185),
.B(n_1043),
.Y(n_1344)
);

INVx3_ASAP7_75t_L g1345 ( 
.A(n_1253),
.Y(n_1345)
);

OR2x2_ASAP7_75t_L g1346 ( 
.A(n_1250),
.B(n_1010),
.Y(n_1346)
);

NAND2xp5_ASAP7_75t_SL g1347 ( 
.A(n_1256),
.B(n_1153),
.Y(n_1347)
);

BUFx6f_ASAP7_75t_L g1348 ( 
.A(n_1281),
.Y(n_1348)
);

NAND2xp5_ASAP7_75t_L g1349 ( 
.A(n_1268),
.B(n_1043),
.Y(n_1349)
);

NOR2xp33_ASAP7_75t_L g1350 ( 
.A(n_1177),
.B(n_1162),
.Y(n_1350)
);

INVxp67_ASAP7_75t_SL g1351 ( 
.A(n_1281),
.Y(n_1351)
);

NAND2xp5_ASAP7_75t_SL g1352 ( 
.A(n_1258),
.B(n_1138),
.Y(n_1352)
);

AND2x4_ASAP7_75t_L g1353 ( 
.A(n_1246),
.B(n_1249),
.Y(n_1353)
);

INVx4_ASAP7_75t_L g1354 ( 
.A(n_1181),
.Y(n_1354)
);

NAND2xp5_ASAP7_75t_L g1355 ( 
.A(n_1269),
.B(n_1043),
.Y(n_1355)
);

AND2x2_ASAP7_75t_L g1356 ( 
.A(n_1202),
.B(n_850),
.Y(n_1356)
);

BUFx6f_ASAP7_75t_L g1357 ( 
.A(n_1271),
.Y(n_1357)
);

INVx4_ASAP7_75t_L g1358 ( 
.A(n_1181),
.Y(n_1358)
);

NAND3xp33_ASAP7_75t_L g1359 ( 
.A(n_1191),
.B(n_864),
.C(n_850),
.Y(n_1359)
);

INVxp67_ASAP7_75t_L g1360 ( 
.A(n_1242),
.Y(n_1360)
);

AND2x2_ASAP7_75t_L g1361 ( 
.A(n_1206),
.B(n_864),
.Y(n_1361)
);

AND2x6_ASAP7_75t_L g1362 ( 
.A(n_1242),
.B(n_1141),
.Y(n_1362)
);

OAI22xp5_ASAP7_75t_L g1363 ( 
.A1(n_1233),
.A2(n_572),
.B1(n_614),
.B2(n_569),
.Y(n_1363)
);

BUFx3_ASAP7_75t_L g1364 ( 
.A(n_1181),
.Y(n_1364)
);

INVxp67_ASAP7_75t_SL g1365 ( 
.A(n_1278),
.Y(n_1365)
);

INVx3_ASAP7_75t_L g1366 ( 
.A(n_1253),
.Y(n_1366)
);

NOR2xp33_ASAP7_75t_L g1367 ( 
.A(n_1177),
.B(n_823),
.Y(n_1367)
);

AOI22xp33_ASAP7_75t_L g1368 ( 
.A1(n_1191),
.A2(n_756),
.B1(n_764),
.B2(n_757),
.Y(n_1368)
);

OR2x2_ASAP7_75t_SL g1369 ( 
.A(n_1211),
.B(n_727),
.Y(n_1369)
);

NAND2xp5_ASAP7_75t_L g1370 ( 
.A(n_1243),
.B(n_1053),
.Y(n_1370)
);

AND2x2_ASAP7_75t_L g1371 ( 
.A(n_1332),
.B(n_1215),
.Y(n_1371)
);

NOR2xp33_ASAP7_75t_L g1372 ( 
.A(n_1360),
.B(n_1162),
.Y(n_1372)
);

INVx1_ASAP7_75t_L g1373 ( 
.A(n_1297),
.Y(n_1373)
);

INVx2_ASAP7_75t_L g1374 ( 
.A(n_1293),
.Y(n_1374)
);

NAND2xp5_ASAP7_75t_L g1375 ( 
.A(n_1307),
.B(n_1360),
.Y(n_1375)
);

INVx2_ASAP7_75t_L g1376 ( 
.A(n_1311),
.Y(n_1376)
);

NAND2xp5_ASAP7_75t_L g1377 ( 
.A(n_1307),
.B(n_1180),
.Y(n_1377)
);

OAI22xp5_ASAP7_75t_L g1378 ( 
.A1(n_1365),
.A2(n_1243),
.B1(n_1262),
.B2(n_1261),
.Y(n_1378)
);

AOI22xp33_ASAP7_75t_L g1379 ( 
.A1(n_1332),
.A2(n_1233),
.B1(n_1190),
.B2(n_1220),
.Y(n_1379)
);

BUFx6f_ASAP7_75t_L g1380 ( 
.A(n_1348),
.Y(n_1380)
);

NOR2xp33_ASAP7_75t_L g1381 ( 
.A(n_1340),
.B(n_1171),
.Y(n_1381)
);

AND2x4_ASAP7_75t_SL g1382 ( 
.A(n_1357),
.B(n_1276),
.Y(n_1382)
);

NAND2xp5_ASAP7_75t_L g1383 ( 
.A(n_1365),
.B(n_1180),
.Y(n_1383)
);

NAND2xp5_ASAP7_75t_L g1384 ( 
.A(n_1306),
.B(n_1173),
.Y(n_1384)
);

AOI22xp5_ASAP7_75t_L g1385 ( 
.A1(n_1363),
.A2(n_1183),
.B1(n_1176),
.B2(n_1270),
.Y(n_1385)
);

NAND2xp5_ASAP7_75t_L g1386 ( 
.A(n_1306),
.B(n_1173),
.Y(n_1386)
);

NAND2xp5_ASAP7_75t_L g1387 ( 
.A(n_1340),
.B(n_1285),
.Y(n_1387)
);

NAND2xp5_ASAP7_75t_L g1388 ( 
.A(n_1363),
.B(n_1215),
.Y(n_1388)
);

NAND2xp5_ASAP7_75t_L g1389 ( 
.A(n_1312),
.B(n_1217),
.Y(n_1389)
);

NAND2xp5_ASAP7_75t_L g1390 ( 
.A(n_1312),
.B(n_1344),
.Y(n_1390)
);

NAND2xp5_ASAP7_75t_L g1391 ( 
.A(n_1344),
.B(n_1217),
.Y(n_1391)
);

AND2x2_ASAP7_75t_L g1392 ( 
.A(n_1356),
.B(n_1171),
.Y(n_1392)
);

NOR2xp33_ASAP7_75t_L g1393 ( 
.A(n_1342),
.B(n_1183),
.Y(n_1393)
);

CKINVDCx5p33_ASAP7_75t_R g1394 ( 
.A(n_1294),
.Y(n_1394)
);

AOI22xp33_ASAP7_75t_L g1395 ( 
.A1(n_1367),
.A2(n_1220),
.B1(n_1257),
.B2(n_1280),
.Y(n_1395)
);

INVx2_ASAP7_75t_L g1396 ( 
.A(n_1313),
.Y(n_1396)
);

AOI22xp33_ASAP7_75t_SL g1397 ( 
.A1(n_1315),
.A2(n_1367),
.B1(n_1350),
.B2(n_1178),
.Y(n_1397)
);

CKINVDCx20_ASAP7_75t_R g1398 ( 
.A(n_1294),
.Y(n_1398)
);

AOI22xp5_ASAP7_75t_L g1399 ( 
.A1(n_1350),
.A2(n_1176),
.B1(n_1270),
.B2(n_1223),
.Y(n_1399)
);

INVx8_ASAP7_75t_L g1400 ( 
.A(n_1316),
.Y(n_1400)
);

OAI22xp5_ASAP7_75t_SL g1401 ( 
.A1(n_1336),
.A2(n_1209),
.B1(n_819),
.B2(n_821),
.Y(n_1401)
);

AOI22xp5_ASAP7_75t_L g1402 ( 
.A1(n_1300),
.A2(n_1223),
.B1(n_1276),
.B2(n_1213),
.Y(n_1402)
);

INVx2_ASAP7_75t_SL g1403 ( 
.A(n_1338),
.Y(n_1403)
);

NAND2xp5_ASAP7_75t_L g1404 ( 
.A(n_1286),
.B(n_1328),
.Y(n_1404)
);

NAND2xp5_ASAP7_75t_L g1405 ( 
.A(n_1328),
.B(n_1216),
.Y(n_1405)
);

AOI22xp5_ASAP7_75t_L g1406 ( 
.A1(n_1300),
.A2(n_1213),
.B1(n_1229),
.B2(n_1207),
.Y(n_1406)
);

OAI22xp5_ASAP7_75t_L g1407 ( 
.A1(n_1370),
.A2(n_1255),
.B1(n_1205),
.B2(n_1228),
.Y(n_1407)
);

NAND2xp5_ASAP7_75t_L g1408 ( 
.A(n_1289),
.B(n_1216),
.Y(n_1408)
);

NAND2xp5_ASAP7_75t_SL g1409 ( 
.A(n_1302),
.B(n_1161),
.Y(n_1409)
);

NAND2xp5_ASAP7_75t_SL g1410 ( 
.A(n_1322),
.B(n_1219),
.Y(n_1410)
);

NAND2xp5_ASAP7_75t_SL g1411 ( 
.A(n_1322),
.B(n_1229),
.Y(n_1411)
);

NAND2xp5_ASAP7_75t_SL g1412 ( 
.A(n_1342),
.B(n_1207),
.Y(n_1412)
);

NAND2xp5_ASAP7_75t_SL g1413 ( 
.A(n_1299),
.B(n_1266),
.Y(n_1413)
);

INVx2_ASAP7_75t_L g1414 ( 
.A(n_1325),
.Y(n_1414)
);

NAND2xp5_ASAP7_75t_L g1415 ( 
.A(n_1289),
.B(n_1170),
.Y(n_1415)
);

INVx2_ASAP7_75t_L g1416 ( 
.A(n_1327),
.Y(n_1416)
);

NOR2xp33_ASAP7_75t_L g1417 ( 
.A(n_1317),
.B(n_1266),
.Y(n_1417)
);

CKINVDCx5p33_ASAP7_75t_R g1418 ( 
.A(n_1316),
.Y(n_1418)
);

NAND2xp5_ASAP7_75t_SL g1419 ( 
.A(n_1299),
.B(n_1254),
.Y(n_1419)
);

AOI22xp33_ASAP7_75t_L g1420 ( 
.A1(n_1362),
.A2(n_1220),
.B1(n_1283),
.B2(n_1282),
.Y(n_1420)
);

NAND2xp5_ASAP7_75t_L g1421 ( 
.A(n_1290),
.B(n_1174),
.Y(n_1421)
);

OAI22xp5_ASAP7_75t_SL g1422 ( 
.A1(n_1369),
.A2(n_807),
.B1(n_1010),
.B2(n_841),
.Y(n_1422)
);

INVx3_ASAP7_75t_L g1423 ( 
.A(n_1301),
.Y(n_1423)
);

AND2x2_ASAP7_75t_L g1424 ( 
.A(n_1361),
.B(n_1272),
.Y(n_1424)
);

NAND2xp5_ASAP7_75t_SL g1425 ( 
.A(n_1302),
.B(n_1161),
.Y(n_1425)
);

AOI22xp5_ASAP7_75t_L g1426 ( 
.A1(n_1359),
.A2(n_1275),
.B1(n_1277),
.B2(n_1274),
.Y(n_1426)
);

AND2x6_ASAP7_75t_SL g1427 ( 
.A(n_1335),
.B(n_895),
.Y(n_1427)
);

OAI21xp5_ASAP7_75t_L g1428 ( 
.A1(n_1290),
.A2(n_1201),
.B(n_1186),
.Y(n_1428)
);

INVx2_ASAP7_75t_L g1429 ( 
.A(n_1329),
.Y(n_1429)
);

AOI21xp5_ASAP7_75t_L g1430 ( 
.A1(n_1302),
.A2(n_1278),
.B(n_1241),
.Y(n_1430)
);

AND2x2_ASAP7_75t_L g1431 ( 
.A(n_1305),
.B(n_1279),
.Y(n_1431)
);

INVx2_ASAP7_75t_L g1432 ( 
.A(n_1334),
.Y(n_1432)
);

OAI22xp33_ASAP7_75t_L g1433 ( 
.A1(n_1315),
.A2(n_1284),
.B1(n_1189),
.B2(n_1198),
.Y(n_1433)
);

NAND2xp5_ASAP7_75t_SL g1434 ( 
.A(n_1302),
.B(n_1248),
.Y(n_1434)
);

INVx2_ASAP7_75t_SL g1435 ( 
.A(n_1291),
.Y(n_1435)
);

NAND2xp5_ASAP7_75t_L g1436 ( 
.A(n_1368),
.B(n_1192),
.Y(n_1436)
);

NAND2xp5_ASAP7_75t_L g1437 ( 
.A(n_1368),
.B(n_1199),
.Y(n_1437)
);

NAND2xp5_ASAP7_75t_L g1438 ( 
.A(n_1370),
.B(n_1288),
.Y(n_1438)
);

OAI21xp33_ASAP7_75t_L g1439 ( 
.A1(n_1305),
.A2(n_841),
.B(n_823),
.Y(n_1439)
);

AOI22xp33_ASAP7_75t_L g1440 ( 
.A1(n_1388),
.A2(n_1341),
.B1(n_1326),
.B2(n_1346),
.Y(n_1440)
);

INVx1_ASAP7_75t_L g1441 ( 
.A(n_1374),
.Y(n_1441)
);

NAND2xp5_ASAP7_75t_L g1442 ( 
.A(n_1371),
.B(n_1353),
.Y(n_1442)
);

OR2x6_ASAP7_75t_L g1443 ( 
.A(n_1404),
.B(n_1309),
.Y(n_1443)
);

INVx2_ASAP7_75t_L g1444 ( 
.A(n_1374),
.Y(n_1444)
);

AND2x4_ASAP7_75t_L g1445 ( 
.A(n_1382),
.B(n_1303),
.Y(n_1445)
);

BUFx12f_ASAP7_75t_L g1446 ( 
.A(n_1418),
.Y(n_1446)
);

O2A1O1Ixp5_ASAP7_75t_L g1447 ( 
.A1(n_1384),
.A2(n_1386),
.B(n_1381),
.C(n_1434),
.Y(n_1447)
);

INVx3_ASAP7_75t_L g1448 ( 
.A(n_1380),
.Y(n_1448)
);

NAND2xp5_ASAP7_75t_L g1449 ( 
.A(n_1389),
.B(n_1353),
.Y(n_1449)
);

AOI22xp5_ASAP7_75t_SL g1450 ( 
.A1(n_1381),
.A2(n_846),
.B1(n_871),
.B2(n_851),
.Y(n_1450)
);

AND2x2_ASAP7_75t_L g1451 ( 
.A(n_1391),
.B(n_1339),
.Y(n_1451)
);

INVx1_ASAP7_75t_L g1452 ( 
.A(n_1376),
.Y(n_1452)
);

INVx1_ASAP7_75t_L g1453 ( 
.A(n_1376),
.Y(n_1453)
);

HB1xp67_ASAP7_75t_L g1454 ( 
.A(n_1435),
.Y(n_1454)
);

AND2x4_ASAP7_75t_L g1455 ( 
.A(n_1382),
.B(n_1303),
.Y(n_1455)
);

INVx2_ASAP7_75t_L g1456 ( 
.A(n_1396),
.Y(n_1456)
);

INVx1_ASAP7_75t_L g1457 ( 
.A(n_1396),
.Y(n_1457)
);

INVx2_ASAP7_75t_L g1458 ( 
.A(n_1414),
.Y(n_1458)
);

AOI22xp33_ASAP7_75t_L g1459 ( 
.A1(n_1397),
.A2(n_1326),
.B1(n_1320),
.B2(n_1200),
.Y(n_1459)
);

INVxp67_ASAP7_75t_L g1460 ( 
.A(n_1393),
.Y(n_1460)
);

INVx1_ASAP7_75t_SL g1461 ( 
.A(n_1398),
.Y(n_1461)
);

INVx2_ASAP7_75t_SL g1462 ( 
.A(n_1403),
.Y(n_1462)
);

BUFx2_ASAP7_75t_L g1463 ( 
.A(n_1375),
.Y(n_1463)
);

BUFx2_ASAP7_75t_L g1464 ( 
.A(n_1380),
.Y(n_1464)
);

NAND2xp5_ASAP7_75t_L g1465 ( 
.A(n_1387),
.B(n_1383),
.Y(n_1465)
);

OAI21xp5_ASAP7_75t_L g1466 ( 
.A1(n_1405),
.A2(n_1288),
.B(n_1347),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_1416),
.Y(n_1467)
);

INVx2_ASAP7_75t_L g1468 ( 
.A(n_1416),
.Y(n_1468)
);

AOI22xp33_ASAP7_75t_L g1469 ( 
.A1(n_1379),
.A2(n_1320),
.B1(n_1333),
.B2(n_1337),
.Y(n_1469)
);

INVx5_ASAP7_75t_L g1470 ( 
.A(n_1380),
.Y(n_1470)
);

INVx2_ASAP7_75t_L g1471 ( 
.A(n_1429),
.Y(n_1471)
);

AOI22xp5_ASAP7_75t_L g1472 ( 
.A1(n_1385),
.A2(n_1259),
.B1(n_1208),
.B2(n_1212),
.Y(n_1472)
);

BUFx6f_ASAP7_75t_L g1473 ( 
.A(n_1400),
.Y(n_1473)
);

HB1xp67_ASAP7_75t_L g1474 ( 
.A(n_1424),
.Y(n_1474)
);

AOI22xp33_ASAP7_75t_L g1475 ( 
.A1(n_1379),
.A2(n_1439),
.B1(n_1419),
.B2(n_1393),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_1429),
.Y(n_1476)
);

INVx1_ASAP7_75t_SL g1477 ( 
.A(n_1392),
.Y(n_1477)
);

O2A1O1Ixp33_ASAP7_75t_L g1478 ( 
.A1(n_1433),
.A2(n_1218),
.B(n_1226),
.C(n_1204),
.Y(n_1478)
);

HB1xp67_ASAP7_75t_L g1479 ( 
.A(n_1423),
.Y(n_1479)
);

INVxp67_ASAP7_75t_L g1480 ( 
.A(n_1417),
.Y(n_1480)
);

INVx2_ASAP7_75t_L g1481 ( 
.A(n_1432),
.Y(n_1481)
);

NAND2xp5_ASAP7_75t_L g1482 ( 
.A(n_1377),
.B(n_1390),
.Y(n_1482)
);

INVxp67_ASAP7_75t_SL g1483 ( 
.A(n_1409),
.Y(n_1483)
);

NAND2xp5_ASAP7_75t_L g1484 ( 
.A(n_1408),
.B(n_1292),
.Y(n_1484)
);

BUFx2_ASAP7_75t_L g1485 ( 
.A(n_1423),
.Y(n_1485)
);

AOI21xp5_ASAP7_75t_L g1486 ( 
.A1(n_1482),
.A2(n_1425),
.B(n_1409),
.Y(n_1486)
);

INVx2_ASAP7_75t_L g1487 ( 
.A(n_1444),
.Y(n_1487)
);

INVx2_ASAP7_75t_L g1488 ( 
.A(n_1444),
.Y(n_1488)
);

NOR2xp33_ASAP7_75t_L g1489 ( 
.A(n_1480),
.B(n_1417),
.Y(n_1489)
);

O2A1O1Ixp33_ASAP7_75t_L g1490 ( 
.A1(n_1447),
.A2(n_1413),
.B(n_1434),
.C(n_1412),
.Y(n_1490)
);

AOI21xp5_ASAP7_75t_L g1491 ( 
.A1(n_1465),
.A2(n_1425),
.B(n_1428),
.Y(n_1491)
);

NOR2xp33_ASAP7_75t_L g1492 ( 
.A(n_1460),
.B(n_1399),
.Y(n_1492)
);

AOI22xp33_ASAP7_75t_L g1493 ( 
.A1(n_1475),
.A2(n_1395),
.B1(n_1259),
.B2(n_1431),
.Y(n_1493)
);

BUFx3_ASAP7_75t_L g1494 ( 
.A(n_1473),
.Y(n_1494)
);

BUFx6f_ASAP7_75t_L g1495 ( 
.A(n_1470),
.Y(n_1495)
);

AO21x1_ASAP7_75t_L g1496 ( 
.A1(n_1472),
.A2(n_1378),
.B(n_1407),
.Y(n_1496)
);

BUFx3_ASAP7_75t_L g1497 ( 
.A(n_1473),
.Y(n_1497)
);

NAND2xp5_ASAP7_75t_L g1498 ( 
.A(n_1449),
.B(n_1484),
.Y(n_1498)
);

AOI21xp5_ASAP7_75t_L g1499 ( 
.A1(n_1466),
.A2(n_1314),
.B(n_1438),
.Y(n_1499)
);

OAI22xp5_ASAP7_75t_L g1500 ( 
.A1(n_1477),
.A2(n_1395),
.B1(n_1406),
.B2(n_1420),
.Y(n_1500)
);

NAND2xp5_ASAP7_75t_L g1501 ( 
.A(n_1442),
.B(n_1372),
.Y(n_1501)
);

BUFx6f_ASAP7_75t_L g1502 ( 
.A(n_1470),
.Y(n_1502)
);

AND2x2_ASAP7_75t_L g1503 ( 
.A(n_1474),
.B(n_1292),
.Y(n_1503)
);

NOR2xp33_ASAP7_75t_L g1504 ( 
.A(n_1477),
.B(n_1372),
.Y(n_1504)
);

OAI22xp5_ASAP7_75t_L g1505 ( 
.A1(n_1450),
.A2(n_1420),
.B1(n_1402),
.B2(n_1436),
.Y(n_1505)
);

INVx2_ASAP7_75t_L g1506 ( 
.A(n_1444),
.Y(n_1506)
);

OAI22xp5_ASAP7_75t_L g1507 ( 
.A1(n_1450),
.A2(n_1437),
.B1(n_1410),
.B2(n_1330),
.Y(n_1507)
);

INVx2_ASAP7_75t_L g1508 ( 
.A(n_1456),
.Y(n_1508)
);

NAND2xp5_ASAP7_75t_L g1509 ( 
.A(n_1463),
.B(n_1254),
.Y(n_1509)
);

OR2x6_ASAP7_75t_L g1510 ( 
.A(n_1443),
.B(n_1400),
.Y(n_1510)
);

NAND2xp5_ASAP7_75t_L g1511 ( 
.A(n_1463),
.B(n_1394),
.Y(n_1511)
);

O2A1O1Ixp33_ASAP7_75t_L g1512 ( 
.A1(n_1478),
.A2(n_1411),
.B(n_833),
.C(n_859),
.Y(n_1512)
);

NAND2xp5_ASAP7_75t_L g1513 ( 
.A(n_1451),
.B(n_1415),
.Y(n_1513)
);

NOR3xp33_ASAP7_75t_SL g1514 ( 
.A(n_1483),
.B(n_1422),
.C(n_1401),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_1441),
.Y(n_1515)
);

AND2x2_ASAP7_75t_L g1516 ( 
.A(n_1451),
.B(n_1287),
.Y(n_1516)
);

NAND2xp5_ASAP7_75t_L g1517 ( 
.A(n_1472),
.B(n_1421),
.Y(n_1517)
);

INVx2_ASAP7_75t_SL g1518 ( 
.A(n_1462),
.Y(n_1518)
);

NAND2xp5_ASAP7_75t_L g1519 ( 
.A(n_1440),
.B(n_1296),
.Y(n_1519)
);

AOI22xp5_ASAP7_75t_SL g1520 ( 
.A1(n_1461),
.A2(n_574),
.B1(n_579),
.B2(n_570),
.Y(n_1520)
);

A2O1A1Ixp33_ASAP7_75t_L g1521 ( 
.A1(n_1469),
.A2(n_1314),
.B(n_1426),
.C(n_1230),
.Y(n_1521)
);

BUFx8_ASAP7_75t_L g1522 ( 
.A(n_1446),
.Y(n_1522)
);

INVx2_ASAP7_75t_L g1523 ( 
.A(n_1456),
.Y(n_1523)
);

OR2x2_ASAP7_75t_L g1524 ( 
.A(n_1454),
.B(n_1373),
.Y(n_1524)
);

AND2x4_ASAP7_75t_L g1525 ( 
.A(n_1473),
.B(n_1287),
.Y(n_1525)
);

AOI21xp5_ASAP7_75t_L g1526 ( 
.A1(n_1443),
.A2(n_1430),
.B(n_1351),
.Y(n_1526)
);

INVx2_ASAP7_75t_L g1527 ( 
.A(n_1456),
.Y(n_1527)
);

BUFx3_ASAP7_75t_L g1528 ( 
.A(n_1473),
.Y(n_1528)
);

BUFx6f_ASAP7_75t_L g1529 ( 
.A(n_1470),
.Y(n_1529)
);

BUFx6f_ASAP7_75t_L g1530 ( 
.A(n_1470),
.Y(n_1530)
);

NAND2xp5_ASAP7_75t_L g1531 ( 
.A(n_1459),
.B(n_1310),
.Y(n_1531)
);

INVx2_ASAP7_75t_L g1532 ( 
.A(n_1458),
.Y(n_1532)
);

O2A1O1Ixp33_ASAP7_75t_L g1533 ( 
.A1(n_1462),
.A2(n_858),
.B(n_865),
.C(n_863),
.Y(n_1533)
);

INVx1_ASAP7_75t_L g1534 ( 
.A(n_1441),
.Y(n_1534)
);

BUFx2_ASAP7_75t_L g1535 ( 
.A(n_1516),
.Y(n_1535)
);

INVx2_ASAP7_75t_L g1536 ( 
.A(n_1487),
.Y(n_1536)
);

AOI22xp5_ASAP7_75t_L g1537 ( 
.A1(n_1507),
.A2(n_965),
.B1(n_970),
.B2(n_960),
.Y(n_1537)
);

BUFx6f_ASAP7_75t_L g1538 ( 
.A(n_1495),
.Y(n_1538)
);

BUFx6f_ASAP7_75t_L g1539 ( 
.A(n_1495),
.Y(n_1539)
);

AOI22xp5_ASAP7_75t_L g1540 ( 
.A1(n_1492),
.A2(n_965),
.B1(n_970),
.B2(n_960),
.Y(n_1540)
);

NOR2xp33_ASAP7_75t_SL g1541 ( 
.A(n_1522),
.B(n_1446),
.Y(n_1541)
);

INVx3_ASAP7_75t_L g1542 ( 
.A(n_1494),
.Y(n_1542)
);

INVx2_ASAP7_75t_SL g1543 ( 
.A(n_1518),
.Y(n_1543)
);

AOI22xp33_ASAP7_75t_L g1544 ( 
.A1(n_1493),
.A2(n_1259),
.B1(n_580),
.B2(n_583),
.Y(n_1544)
);

AND2x2_ASAP7_75t_L g1545 ( 
.A(n_1503),
.B(n_1485),
.Y(n_1545)
);

INVx2_ASAP7_75t_SL g1546 ( 
.A(n_1524),
.Y(n_1546)
);

BUFx3_ASAP7_75t_L g1547 ( 
.A(n_1525),
.Y(n_1547)
);

INVx2_ASAP7_75t_SL g1548 ( 
.A(n_1522),
.Y(n_1548)
);

BUFx2_ASAP7_75t_L g1549 ( 
.A(n_1511),
.Y(n_1549)
);

AOI22xp33_ASAP7_75t_L g1550 ( 
.A1(n_1493),
.A2(n_1492),
.B1(n_1500),
.B2(n_1505),
.Y(n_1550)
);

BUFx4f_ASAP7_75t_L g1551 ( 
.A(n_1525),
.Y(n_1551)
);

INVx2_ASAP7_75t_L g1552 ( 
.A(n_1487),
.Y(n_1552)
);

NAND2x1p5_ASAP7_75t_L g1553 ( 
.A(n_1495),
.B(n_1470),
.Y(n_1553)
);

AND2x4_ASAP7_75t_L g1554 ( 
.A(n_1510),
.B(n_1473),
.Y(n_1554)
);

BUFx12f_ASAP7_75t_L g1555 ( 
.A(n_1495),
.Y(n_1555)
);

AND2x4_ASAP7_75t_L g1556 ( 
.A(n_1510),
.B(n_1473),
.Y(n_1556)
);

A2O1A1Ixp33_ASAP7_75t_L g1557 ( 
.A1(n_1490),
.A2(n_1330),
.B(n_1351),
.C(n_1445),
.Y(n_1557)
);

HB1xp67_ASAP7_75t_L g1558 ( 
.A(n_1515),
.Y(n_1558)
);

BUFx6f_ASAP7_75t_L g1559 ( 
.A(n_1502),
.Y(n_1559)
);

OAI22xp5_ASAP7_75t_L g1560 ( 
.A1(n_1504),
.A2(n_1343),
.B1(n_1335),
.B2(n_1443),
.Y(n_1560)
);

INVx2_ASAP7_75t_SL g1561 ( 
.A(n_1494),
.Y(n_1561)
);

INVx2_ASAP7_75t_L g1562 ( 
.A(n_1488),
.Y(n_1562)
);

NAND2xp5_ASAP7_75t_L g1563 ( 
.A(n_1498),
.B(n_1452),
.Y(n_1563)
);

HB1xp67_ASAP7_75t_L g1564 ( 
.A(n_1534),
.Y(n_1564)
);

INVx1_ASAP7_75t_L g1565 ( 
.A(n_1488),
.Y(n_1565)
);

AOI21xp5_ASAP7_75t_L g1566 ( 
.A1(n_1499),
.A2(n_1443),
.B(n_1345),
.Y(n_1566)
);

INVx1_ASAP7_75t_L g1567 ( 
.A(n_1506),
.Y(n_1567)
);

BUFx6f_ASAP7_75t_L g1568 ( 
.A(n_1502),
.Y(n_1568)
);

CKINVDCx20_ASAP7_75t_R g1569 ( 
.A(n_1514),
.Y(n_1569)
);

HB1xp67_ASAP7_75t_L g1570 ( 
.A(n_1510),
.Y(n_1570)
);

INVx2_ASAP7_75t_SL g1571 ( 
.A(n_1497),
.Y(n_1571)
);

BUFx2_ASAP7_75t_L g1572 ( 
.A(n_1497),
.Y(n_1572)
);

AOI221xp5_ASAP7_75t_L g1573 ( 
.A1(n_1512),
.A2(n_789),
.B1(n_851),
.B2(n_871),
.C(n_846),
.Y(n_1573)
);

INVx4_ASAP7_75t_L g1574 ( 
.A(n_1502),
.Y(n_1574)
);

INVx3_ASAP7_75t_L g1575 ( 
.A(n_1528),
.Y(n_1575)
);

CKINVDCx6p67_ASAP7_75t_R g1576 ( 
.A(n_1528),
.Y(n_1576)
);

CKINVDCx5p33_ASAP7_75t_R g1577 ( 
.A(n_1489),
.Y(n_1577)
);

INVx3_ASAP7_75t_L g1578 ( 
.A(n_1502),
.Y(n_1578)
);

INVx2_ASAP7_75t_L g1579 ( 
.A(n_1506),
.Y(n_1579)
);

BUFx6f_ASAP7_75t_L g1580 ( 
.A(n_1529),
.Y(n_1580)
);

NOR3xp33_ASAP7_75t_L g1581 ( 
.A(n_1531),
.B(n_868),
.C(n_866),
.Y(n_1581)
);

OR2x6_ASAP7_75t_L g1582 ( 
.A(n_1526),
.B(n_1443),
.Y(n_1582)
);

INVx1_ASAP7_75t_L g1583 ( 
.A(n_1508),
.Y(n_1583)
);

NAND2xp5_ASAP7_75t_L g1584 ( 
.A(n_1501),
.B(n_1452),
.Y(n_1584)
);

BUFx6f_ASAP7_75t_L g1585 ( 
.A(n_1529),
.Y(n_1585)
);

BUFx8_ASAP7_75t_SL g1586 ( 
.A(n_1529),
.Y(n_1586)
);

NAND3xp33_ASAP7_75t_L g1587 ( 
.A(n_1514),
.B(n_975),
.C(n_969),
.Y(n_1587)
);

AND2x4_ASAP7_75t_L g1588 ( 
.A(n_1508),
.B(n_1448),
.Y(n_1588)
);

AOI22xp33_ASAP7_75t_L g1589 ( 
.A1(n_1517),
.A2(n_580),
.B1(n_583),
.B2(n_579),
.Y(n_1589)
);

NAND2xp5_ASAP7_75t_L g1590 ( 
.A(n_1513),
.B(n_1453),
.Y(n_1590)
);

INVx1_ASAP7_75t_L g1591 ( 
.A(n_1527),
.Y(n_1591)
);

AND2x2_ASAP7_75t_L g1592 ( 
.A(n_1504),
.B(n_1485),
.Y(n_1592)
);

AND2x4_ASAP7_75t_L g1593 ( 
.A(n_1527),
.B(n_1448),
.Y(n_1593)
);

CKINVDCx5p33_ASAP7_75t_R g1594 ( 
.A(n_1520),
.Y(n_1594)
);

BUFx3_ASAP7_75t_L g1595 ( 
.A(n_1529),
.Y(n_1595)
);

CKINVDCx5p33_ASAP7_75t_R g1596 ( 
.A(n_1509),
.Y(n_1596)
);

INVx3_ASAP7_75t_L g1597 ( 
.A(n_1530),
.Y(n_1597)
);

BUFx3_ASAP7_75t_L g1598 ( 
.A(n_1530),
.Y(n_1598)
);

A2O1A1Ixp33_ASAP7_75t_L g1599 ( 
.A1(n_1537),
.A2(n_1521),
.B(n_1519),
.C(n_1491),
.Y(n_1599)
);

NAND2xp5_ASAP7_75t_L g1600 ( 
.A(n_1546),
.B(n_1486),
.Y(n_1600)
);

INVx1_ASAP7_75t_L g1601 ( 
.A(n_1558),
.Y(n_1601)
);

O2A1O1Ixp33_ASAP7_75t_SL g1602 ( 
.A1(n_1569),
.A2(n_1587),
.B(n_1540),
.C(n_1548),
.Y(n_1602)
);

A2O1A1Ixp33_ASAP7_75t_L g1603 ( 
.A1(n_1550),
.A2(n_1521),
.B(n_1533),
.C(n_1455),
.Y(n_1603)
);

NAND3xp33_ASAP7_75t_L g1604 ( 
.A(n_1589),
.B(n_975),
.C(n_969),
.Y(n_1604)
);

OAI21x1_ASAP7_75t_L g1605 ( 
.A1(n_1566),
.A2(n_1496),
.B(n_1523),
.Y(n_1605)
);

INVx1_ASAP7_75t_L g1606 ( 
.A(n_1558),
.Y(n_1606)
);

OAI21xp5_ASAP7_75t_L g1607 ( 
.A1(n_1581),
.A2(n_1352),
.B(n_1347),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_1564),
.Y(n_1608)
);

AOI221xp5_ASAP7_75t_SL g1609 ( 
.A1(n_1569),
.A2(n_610),
.B1(n_839),
.B2(n_837),
.C(n_834),
.Y(n_1609)
);

NAND2xp5_ASAP7_75t_L g1610 ( 
.A(n_1549),
.B(n_1532),
.Y(n_1610)
);

OAI21x1_ASAP7_75t_L g1611 ( 
.A1(n_1578),
.A2(n_1352),
.B(n_1106),
.Y(n_1611)
);

INVx2_ASAP7_75t_L g1612 ( 
.A(n_1536),
.Y(n_1612)
);

NOR2x1_ASAP7_75t_R g1613 ( 
.A(n_1594),
.B(n_977),
.Y(n_1613)
);

BUFx3_ASAP7_75t_L g1614 ( 
.A(n_1535),
.Y(n_1614)
);

OAI22xp33_ASAP7_75t_L g1615 ( 
.A1(n_1596),
.A2(n_1335),
.B1(n_1000),
.B2(n_1012),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_1564),
.Y(n_1616)
);

OAI22xp5_ASAP7_75t_L g1617 ( 
.A1(n_1550),
.A2(n_1455),
.B1(n_1445),
.B2(n_1446),
.Y(n_1617)
);

INVx4_ASAP7_75t_L g1618 ( 
.A(n_1542),
.Y(n_1618)
);

OAI222xp33_ASAP7_75t_L g1619 ( 
.A1(n_1544),
.A2(n_634),
.B1(n_589),
.B2(n_636),
.C1(n_633),
.C2(n_588),
.Y(n_1619)
);

A2O1A1Ixp33_ASAP7_75t_L g1620 ( 
.A1(n_1544),
.A2(n_1455),
.B(n_1445),
.C(n_589),
.Y(n_1620)
);

INVx4_ASAP7_75t_L g1621 ( 
.A(n_1542),
.Y(n_1621)
);

AOI21xp5_ASAP7_75t_L g1622 ( 
.A1(n_1557),
.A2(n_1530),
.B(n_1345),
.Y(n_1622)
);

OAI22xp5_ASAP7_75t_L g1623 ( 
.A1(n_1589),
.A2(n_1455),
.B1(n_1445),
.B2(n_1000),
.Y(n_1623)
);

AOI21xp5_ASAP7_75t_L g1624 ( 
.A1(n_1557),
.A2(n_1530),
.B(n_1366),
.Y(n_1624)
);

AO31x2_ASAP7_75t_L g1625 ( 
.A1(n_1536),
.A2(n_1471),
.A3(n_1481),
.B(n_1468),
.Y(n_1625)
);

AOI22xp33_ASAP7_75t_L g1626 ( 
.A1(n_1596),
.A2(n_1012),
.B1(n_977),
.B2(n_899),
.Y(n_1626)
);

NAND3xp33_ASAP7_75t_L g1627 ( 
.A(n_1573),
.B(n_1560),
.C(n_1577),
.Y(n_1627)
);

AOI22xp33_ASAP7_75t_L g1628 ( 
.A1(n_1570),
.A2(n_899),
.B1(n_936),
.B2(n_895),
.Y(n_1628)
);

OAI21xp5_ASAP7_75t_L g1629 ( 
.A1(n_1584),
.A2(n_873),
.B(n_869),
.Y(n_1629)
);

OAI22xp5_ASAP7_75t_L g1630 ( 
.A1(n_1543),
.A2(n_1035),
.B1(n_1309),
.B2(n_1321),
.Y(n_1630)
);

INVxp67_ASAP7_75t_SL g1631 ( 
.A(n_1552),
.Y(n_1631)
);

NAND2xp5_ASAP7_75t_SL g1632 ( 
.A(n_1551),
.B(n_1357),
.Y(n_1632)
);

AOI21xp5_ASAP7_75t_L g1633 ( 
.A1(n_1582),
.A2(n_1366),
.B(n_1331),
.Y(n_1633)
);

AOI21xp5_ASAP7_75t_L g1634 ( 
.A1(n_1582),
.A2(n_1331),
.B(n_1295),
.Y(n_1634)
);

AOI22xp33_ASAP7_75t_L g1635 ( 
.A1(n_1570),
.A2(n_939),
.B1(n_1003),
.B2(n_936),
.Y(n_1635)
);

AND2x2_ASAP7_75t_L g1636 ( 
.A(n_1592),
.B(n_1464),
.Y(n_1636)
);

AOI22xp33_ASAP7_75t_L g1637 ( 
.A1(n_1547),
.A2(n_1003),
.B1(n_1004),
.B2(n_939),
.Y(n_1637)
);

CKINVDCx5p33_ASAP7_75t_R g1638 ( 
.A(n_1586),
.Y(n_1638)
);

AO32x2_ASAP7_75t_L g1639 ( 
.A1(n_1561),
.A2(n_1571),
.A3(n_1574),
.B1(n_1582),
.B2(n_1579),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_1565),
.Y(n_1640)
);

NOR2xp33_ASAP7_75t_L g1641 ( 
.A(n_1545),
.B(n_1004),
.Y(n_1641)
);

AO21x2_ASAP7_75t_L g1642 ( 
.A1(n_1567),
.A2(n_1251),
.B(n_1453),
.Y(n_1642)
);

AOI21xp5_ASAP7_75t_L g1643 ( 
.A1(n_1551),
.A2(n_1295),
.B(n_1470),
.Y(n_1643)
);

AOI21xp5_ASAP7_75t_L g1644 ( 
.A1(n_1563),
.A2(n_1590),
.B(n_1553),
.Y(n_1644)
);

AND2x4_ASAP7_75t_L g1645 ( 
.A(n_1554),
.B(n_1464),
.Y(n_1645)
);

BUFx6f_ASAP7_75t_L g1646 ( 
.A(n_1538),
.Y(n_1646)
);

AOI221xp5_ASAP7_75t_SL g1647 ( 
.A1(n_1572),
.A2(n_610),
.B1(n_840),
.B2(n_877),
.C(n_874),
.Y(n_1647)
);

O2A1O1Ixp33_ASAP7_75t_L g1648 ( 
.A1(n_1541),
.A2(n_695),
.B(n_697),
.C(n_694),
.Y(n_1648)
);

AND2x4_ASAP7_75t_L g1649 ( 
.A(n_1554),
.B(n_1448),
.Y(n_1649)
);

OR2x6_ASAP7_75t_L g1650 ( 
.A(n_1554),
.B(n_1400),
.Y(n_1650)
);

BUFx6f_ASAP7_75t_L g1651 ( 
.A(n_1538),
.Y(n_1651)
);

NAND2xp5_ASAP7_75t_L g1652 ( 
.A(n_1583),
.B(n_1457),
.Y(n_1652)
);

NAND2xp5_ASAP7_75t_L g1653 ( 
.A(n_1591),
.B(n_1457),
.Y(n_1653)
);

INVx1_ASAP7_75t_L g1654 ( 
.A(n_1552),
.Y(n_1654)
);

OAI21x1_ASAP7_75t_L g1655 ( 
.A1(n_1597),
.A2(n_1081),
.B(n_1349),
.Y(n_1655)
);

BUFx12f_ASAP7_75t_L g1656 ( 
.A(n_1555),
.Y(n_1656)
);

O2A1O1Ixp33_ASAP7_75t_SL g1657 ( 
.A1(n_1575),
.A2(n_1479),
.B(n_1476),
.C(n_1467),
.Y(n_1657)
);

OAI21xp5_ASAP7_75t_L g1658 ( 
.A1(n_1556),
.A2(n_1240),
.B(n_1186),
.Y(n_1658)
);

AOI21xp5_ASAP7_75t_L g1659 ( 
.A1(n_1556),
.A2(n_1201),
.B(n_1319),
.Y(n_1659)
);

OAI21x1_ASAP7_75t_L g1660 ( 
.A1(n_1562),
.A2(n_1355),
.B(n_1349),
.Y(n_1660)
);

BUFx10_ASAP7_75t_L g1661 ( 
.A(n_1538),
.Y(n_1661)
);

INVx1_ASAP7_75t_L g1662 ( 
.A(n_1562),
.Y(n_1662)
);

CKINVDCx5p33_ASAP7_75t_R g1663 ( 
.A(n_1586),
.Y(n_1663)
);

INVxp67_ASAP7_75t_L g1664 ( 
.A(n_1547),
.Y(n_1664)
);

A2O1A1Ixp33_ASAP7_75t_L g1665 ( 
.A1(n_1598),
.A2(n_633),
.B(n_634),
.C(n_588),
.Y(n_1665)
);

AOI21xp5_ASAP7_75t_L g1666 ( 
.A1(n_1538),
.A2(n_1304),
.B(n_1301),
.Y(n_1666)
);

BUFx5_ASAP7_75t_L g1667 ( 
.A(n_1555),
.Y(n_1667)
);

BUFx2_ASAP7_75t_L g1668 ( 
.A(n_1576),
.Y(n_1668)
);

A2O1A1Ixp33_ASAP7_75t_L g1669 ( 
.A1(n_1595),
.A2(n_636),
.B(n_809),
.C(n_758),
.Y(n_1669)
);

BUFx12f_ASAP7_75t_L g1670 ( 
.A(n_1539),
.Y(n_1670)
);

AOI21xp5_ASAP7_75t_L g1671 ( 
.A1(n_1539),
.A2(n_1304),
.B(n_1301),
.Y(n_1671)
);

CKINVDCx16_ASAP7_75t_R g1672 ( 
.A(n_1598),
.Y(n_1672)
);

NAND2xp5_ASAP7_75t_L g1673 ( 
.A(n_1588),
.B(n_1467),
.Y(n_1673)
);

O2A1O1Ixp33_ASAP7_75t_L g1674 ( 
.A1(n_1588),
.A2(n_702),
.B(n_704),
.C(n_701),
.Y(n_1674)
);

AOI22xp33_ASAP7_75t_L g1675 ( 
.A1(n_1588),
.A2(n_1005),
.B1(n_926),
.B2(n_924),
.Y(n_1675)
);

AOI22xp33_ASAP7_75t_L g1676 ( 
.A1(n_1593),
.A2(n_1005),
.B1(n_926),
.B2(n_1029),
.Y(n_1676)
);

NAND3xp33_ASAP7_75t_L g1677 ( 
.A(n_1627),
.B(n_610),
.C(n_538),
.Y(n_1677)
);

BUFx3_ASAP7_75t_L g1678 ( 
.A(n_1614),
.Y(n_1678)
);

OR2x6_ASAP7_75t_L g1679 ( 
.A(n_1644),
.B(n_1579),
.Y(n_1679)
);

INVx1_ASAP7_75t_L g1680 ( 
.A(n_1601),
.Y(n_1680)
);

NAND2x1p5_ASAP7_75t_L g1681 ( 
.A(n_1618),
.B(n_1539),
.Y(n_1681)
);

OR2x2_ASAP7_75t_L g1682 ( 
.A(n_1606),
.B(n_1593),
.Y(n_1682)
);

OAI22xp5_ASAP7_75t_L g1683 ( 
.A1(n_1604),
.A2(n_1568),
.B1(n_1580),
.B2(n_1559),
.Y(n_1683)
);

INVx4_ASAP7_75t_L g1684 ( 
.A(n_1656),
.Y(n_1684)
);

INVx2_ASAP7_75t_L g1685 ( 
.A(n_1612),
.Y(n_1685)
);

AOI22xp5_ASAP7_75t_L g1686 ( 
.A1(n_1623),
.A2(n_1362),
.B1(n_539),
.B2(n_540),
.Y(n_1686)
);

INVx1_ASAP7_75t_L g1687 ( 
.A(n_1608),
.Y(n_1687)
);

INVx2_ASAP7_75t_L g1688 ( 
.A(n_1654),
.Y(n_1688)
);

AOI221xp5_ASAP7_75t_L g1689 ( 
.A1(n_1619),
.A2(n_544),
.B1(n_548),
.B2(n_541),
.C(n_537),
.Y(n_1689)
);

NOR2xp33_ASAP7_75t_L g1690 ( 
.A(n_1615),
.B(n_1427),
.Y(n_1690)
);

AOI22xp33_ASAP7_75t_L g1691 ( 
.A1(n_1617),
.A2(n_1029),
.B1(n_1362),
.B2(n_610),
.Y(n_1691)
);

OR2x6_ASAP7_75t_L g1692 ( 
.A(n_1650),
.B(n_1559),
.Y(n_1692)
);

NOR2x1_ASAP7_75t_SL g1693 ( 
.A(n_1642),
.B(n_1559),
.Y(n_1693)
);

INVx1_ASAP7_75t_L g1694 ( 
.A(n_1616),
.Y(n_1694)
);

HB1xp67_ASAP7_75t_L g1695 ( 
.A(n_1600),
.Y(n_1695)
);

AOI22xp5_ASAP7_75t_L g1696 ( 
.A1(n_1620),
.A2(n_1362),
.B1(n_550),
.B2(n_551),
.Y(n_1696)
);

OAI22xp5_ASAP7_75t_L g1697 ( 
.A1(n_1603),
.A2(n_1568),
.B1(n_1580),
.B2(n_1559),
.Y(n_1697)
);

CKINVDCx5p33_ASAP7_75t_R g1698 ( 
.A(n_1638),
.Y(n_1698)
);

INVx2_ASAP7_75t_L g1699 ( 
.A(n_1662),
.Y(n_1699)
);

INVx2_ASAP7_75t_L g1700 ( 
.A(n_1640),
.Y(n_1700)
);

NAND3xp33_ASAP7_75t_L g1701 ( 
.A(n_1599),
.B(n_552),
.C(n_549),
.Y(n_1701)
);

BUFx12f_ASAP7_75t_L g1702 ( 
.A(n_1663),
.Y(n_1702)
);

AND2x2_ASAP7_75t_L g1703 ( 
.A(n_1672),
.B(n_1593),
.Y(n_1703)
);

AOI22xp5_ASAP7_75t_L g1704 ( 
.A1(n_1602),
.A2(n_1609),
.B1(n_1607),
.B2(n_1630),
.Y(n_1704)
);

OR2x6_ASAP7_75t_L g1705 ( 
.A(n_1650),
.B(n_1668),
.Y(n_1705)
);

NAND2x1_ASAP7_75t_L g1706 ( 
.A(n_1621),
.B(n_1568),
.Y(n_1706)
);

INVx1_ASAP7_75t_L g1707 ( 
.A(n_1631),
.Y(n_1707)
);

CKINVDCx11_ASAP7_75t_R g1708 ( 
.A(n_1670),
.Y(n_1708)
);

NOR2xp33_ASAP7_75t_L g1709 ( 
.A(n_1641),
.B(n_918),
.Y(n_1709)
);

INVx1_ASAP7_75t_SL g1710 ( 
.A(n_1636),
.Y(n_1710)
);

INVx1_ASAP7_75t_L g1711 ( 
.A(n_1610),
.Y(n_1711)
);

AO21x2_ASAP7_75t_L g1712 ( 
.A1(n_1605),
.A2(n_1251),
.B(n_1476),
.Y(n_1712)
);

OAI22xp5_ASAP7_75t_L g1713 ( 
.A1(n_1626),
.A2(n_1580),
.B1(n_1585),
.B2(n_1568),
.Y(n_1713)
);

BUFx3_ASAP7_75t_L g1714 ( 
.A(n_1646),
.Y(n_1714)
);

AOI21xp5_ASAP7_75t_L g1715 ( 
.A1(n_1643),
.A2(n_1585),
.B(n_1580),
.Y(n_1715)
);

BUFx2_ASAP7_75t_L g1716 ( 
.A(n_1664),
.Y(n_1716)
);

AOI22xp33_ASAP7_75t_L g1717 ( 
.A1(n_1645),
.A2(n_1362),
.B1(n_711),
.B2(n_713),
.Y(n_1717)
);

INVx1_ASAP7_75t_L g1718 ( 
.A(n_1639),
.Y(n_1718)
);

INVx1_ASAP7_75t_L g1719 ( 
.A(n_1639),
.Y(n_1719)
);

AND2x4_ASAP7_75t_L g1720 ( 
.A(n_1645),
.B(n_1585),
.Y(n_1720)
);

CKINVDCx20_ASAP7_75t_R g1721 ( 
.A(n_1632),
.Y(n_1721)
);

OAI22xp5_ASAP7_75t_L g1722 ( 
.A1(n_1675),
.A2(n_1635),
.B1(n_1628),
.B2(n_1676),
.Y(n_1722)
);

INVx1_ASAP7_75t_L g1723 ( 
.A(n_1639),
.Y(n_1723)
);

INVx4_ASAP7_75t_L g1724 ( 
.A(n_1646),
.Y(n_1724)
);

AOI221xp5_ASAP7_75t_L g1725 ( 
.A1(n_1648),
.A2(n_559),
.B1(n_561),
.B2(n_558),
.C(n_555),
.Y(n_1725)
);

INVx1_ASAP7_75t_SL g1726 ( 
.A(n_1649),
.Y(n_1726)
);

AND2x4_ASAP7_75t_L g1727 ( 
.A(n_1649),
.B(n_1585),
.Y(n_1727)
);

AOI22xp33_ASAP7_75t_L g1728 ( 
.A1(n_1637),
.A2(n_714),
.B1(n_716),
.B2(n_707),
.Y(n_1728)
);

INVx4_ASAP7_75t_L g1729 ( 
.A(n_1646),
.Y(n_1729)
);

CKINVDCx8_ASAP7_75t_R g1730 ( 
.A(n_1651),
.Y(n_1730)
);

INVx1_ASAP7_75t_L g1731 ( 
.A(n_1652),
.Y(n_1731)
);

BUFx3_ASAP7_75t_L g1732 ( 
.A(n_1651),
.Y(n_1732)
);

INVx1_ASAP7_75t_L g1733 ( 
.A(n_1653),
.Y(n_1733)
);

OAI21xp5_ASAP7_75t_SL g1734 ( 
.A1(n_1669),
.A2(n_1197),
.B(n_1260),
.Y(n_1734)
);

OAI21x1_ASAP7_75t_L g1735 ( 
.A1(n_1718),
.A2(n_1634),
.B(n_1633),
.Y(n_1735)
);

INVx2_ASAP7_75t_L g1736 ( 
.A(n_1719),
.Y(n_1736)
);

BUFx12f_ASAP7_75t_L g1737 ( 
.A(n_1684),
.Y(n_1737)
);

OAI21x1_ASAP7_75t_L g1738 ( 
.A1(n_1723),
.A2(n_1624),
.B(n_1622),
.Y(n_1738)
);

OAI21x1_ASAP7_75t_L g1739 ( 
.A1(n_1715),
.A2(n_1660),
.B(n_1655),
.Y(n_1739)
);

INVx1_ASAP7_75t_L g1740 ( 
.A(n_1680),
.Y(n_1740)
);

HB1xp67_ASAP7_75t_L g1741 ( 
.A(n_1695),
.Y(n_1741)
);

AND2x4_ASAP7_75t_L g1742 ( 
.A(n_1679),
.B(n_1625),
.Y(n_1742)
);

AOI22xp33_ASAP7_75t_L g1743 ( 
.A1(n_1701),
.A2(n_1629),
.B1(n_564),
.B2(n_565),
.Y(n_1743)
);

INVx1_ASAP7_75t_L g1744 ( 
.A(n_1687),
.Y(n_1744)
);

INVx1_ASAP7_75t_L g1745 ( 
.A(n_1694),
.Y(n_1745)
);

AOI21xp5_ASAP7_75t_L g1746 ( 
.A1(n_1701),
.A2(n_1657),
.B(n_1659),
.Y(n_1746)
);

INVx2_ASAP7_75t_L g1747 ( 
.A(n_1688),
.Y(n_1747)
);

OR2x2_ASAP7_75t_L g1748 ( 
.A(n_1707),
.B(n_1673),
.Y(n_1748)
);

NAND2xp5_ASAP7_75t_L g1749 ( 
.A(n_1711),
.B(n_1625),
.Y(n_1749)
);

NAND2xp5_ASAP7_75t_L g1750 ( 
.A(n_1731),
.B(n_1625),
.Y(n_1750)
);

INVx1_ASAP7_75t_L g1751 ( 
.A(n_1700),
.Y(n_1751)
);

INVx2_ASAP7_75t_L g1752 ( 
.A(n_1699),
.Y(n_1752)
);

INVx1_ASAP7_75t_L g1753 ( 
.A(n_1685),
.Y(n_1753)
);

NAND2xp33_ASAP7_75t_L g1754 ( 
.A(n_1677),
.B(n_1667),
.Y(n_1754)
);

INVx2_ASAP7_75t_L g1755 ( 
.A(n_1679),
.Y(n_1755)
);

INVx3_ASAP7_75t_L g1756 ( 
.A(n_1679),
.Y(n_1756)
);

INVx2_ASAP7_75t_L g1757 ( 
.A(n_1733),
.Y(n_1757)
);

NAND2xp5_ASAP7_75t_L g1758 ( 
.A(n_1710),
.B(n_1647),
.Y(n_1758)
);

AND2x2_ASAP7_75t_L g1759 ( 
.A(n_1682),
.B(n_1726),
.Y(n_1759)
);

INVx2_ASAP7_75t_L g1760 ( 
.A(n_1712),
.Y(n_1760)
);

AND2x2_ASAP7_75t_L g1761 ( 
.A(n_1716),
.B(n_1661),
.Y(n_1761)
);

CKINVDCx20_ASAP7_75t_R g1762 ( 
.A(n_1708),
.Y(n_1762)
);

INVx2_ASAP7_75t_SL g1763 ( 
.A(n_1705),
.Y(n_1763)
);

INVx3_ASAP7_75t_L g1764 ( 
.A(n_1712),
.Y(n_1764)
);

INVx2_ASAP7_75t_L g1765 ( 
.A(n_1693),
.Y(n_1765)
);

INVx1_ASAP7_75t_L g1766 ( 
.A(n_1703),
.Y(n_1766)
);

INVx2_ASAP7_75t_L g1767 ( 
.A(n_1727),
.Y(n_1767)
);

INVx1_ASAP7_75t_L g1768 ( 
.A(n_1720),
.Y(n_1768)
);

OAI21x1_ASAP7_75t_L g1769 ( 
.A1(n_1697),
.A2(n_1706),
.B(n_1611),
.Y(n_1769)
);

AOI222xp33_ASAP7_75t_L g1770 ( 
.A1(n_1743),
.A2(n_1677),
.B1(n_1689),
.B2(n_1722),
.C1(n_1725),
.C2(n_1690),
.Y(n_1770)
);

AOI22xp33_ASAP7_75t_L g1771 ( 
.A1(n_1743),
.A2(n_1686),
.B1(n_1691),
.B2(n_1683),
.Y(n_1771)
);

AOI321xp33_ASAP7_75t_L g1772 ( 
.A1(n_1746),
.A2(n_1704),
.A3(n_1713),
.B1(n_1686),
.B2(n_1758),
.C(n_1696),
.Y(n_1772)
);

OAI22xp33_ASAP7_75t_L g1773 ( 
.A1(n_1746),
.A2(n_1704),
.B1(n_1705),
.B2(n_1692),
.Y(n_1773)
);

INVxp67_ASAP7_75t_L g1774 ( 
.A(n_1741),
.Y(n_1774)
);

NAND2xp5_ASAP7_75t_L g1775 ( 
.A(n_1741),
.B(n_1748),
.Y(n_1775)
);

OAI22xp5_ASAP7_75t_L g1776 ( 
.A1(n_1758),
.A2(n_1721),
.B1(n_1692),
.B2(n_1696),
.Y(n_1776)
);

AOI22xp33_ASAP7_75t_L g1777 ( 
.A1(n_1754),
.A2(n_1684),
.B1(n_1709),
.B2(n_1678),
.Y(n_1777)
);

AOI21xp5_ASAP7_75t_L g1778 ( 
.A1(n_1754),
.A2(n_1734),
.B(n_1658),
.Y(n_1778)
);

OAI22xp5_ASAP7_75t_L g1779 ( 
.A1(n_1763),
.A2(n_1730),
.B1(n_1727),
.B2(n_1720),
.Y(n_1779)
);

INVx1_ASAP7_75t_L g1780 ( 
.A(n_1740),
.Y(n_1780)
);

AOI22xp33_ASAP7_75t_SL g1781 ( 
.A1(n_1762),
.A2(n_885),
.B1(n_1667),
.B2(n_1702),
.Y(n_1781)
);

INVx2_ASAP7_75t_L g1782 ( 
.A(n_1747),
.Y(n_1782)
);

AOI22xp33_ASAP7_75t_L g1783 ( 
.A1(n_1763),
.A2(n_1717),
.B1(n_1728),
.B2(n_1714),
.Y(n_1783)
);

AND2x2_ASAP7_75t_L g1784 ( 
.A(n_1767),
.B(n_1763),
.Y(n_1784)
);

AO21x2_ASAP7_75t_L g1785 ( 
.A1(n_1760),
.A2(n_1671),
.B(n_1666),
.Y(n_1785)
);

INVx1_ASAP7_75t_L g1786 ( 
.A(n_1747),
.Y(n_1786)
);

AO22x1_ASAP7_75t_L g1787 ( 
.A1(n_1765),
.A2(n_1698),
.B1(n_1729),
.B2(n_1724),
.Y(n_1787)
);

AND2x4_ASAP7_75t_L g1788 ( 
.A(n_1756),
.B(n_1724),
.Y(n_1788)
);

AND2x4_ASAP7_75t_L g1789 ( 
.A(n_1756),
.B(n_1755),
.Y(n_1789)
);

AOI22xp33_ASAP7_75t_L g1790 ( 
.A1(n_1737),
.A2(n_1767),
.B1(n_1768),
.B2(n_1766),
.Y(n_1790)
);

INVx2_ASAP7_75t_L g1791 ( 
.A(n_1747),
.Y(n_1791)
);

AOI21xp33_ASAP7_75t_L g1792 ( 
.A1(n_1755),
.A2(n_1613),
.B(n_1674),
.Y(n_1792)
);

OAI22xp33_ASAP7_75t_L g1793 ( 
.A1(n_1767),
.A2(n_1681),
.B1(n_1729),
.B2(n_1732),
.Y(n_1793)
);

INVx2_ASAP7_75t_L g1794 ( 
.A(n_1747),
.Y(n_1794)
);

INVx1_ASAP7_75t_L g1795 ( 
.A(n_1780),
.Y(n_1795)
);

OR2x2_ASAP7_75t_L g1796 ( 
.A(n_1775),
.B(n_1774),
.Y(n_1796)
);

INVx1_ASAP7_75t_L g1797 ( 
.A(n_1786),
.Y(n_1797)
);

INVx1_ASAP7_75t_L g1798 ( 
.A(n_1786),
.Y(n_1798)
);

INVx1_ASAP7_75t_L g1799 ( 
.A(n_1782),
.Y(n_1799)
);

AOI221xp5_ASAP7_75t_L g1800 ( 
.A1(n_1773),
.A2(n_604),
.B1(n_605),
.B2(n_596),
.C(n_562),
.Y(n_1800)
);

AND2x2_ASAP7_75t_L g1801 ( 
.A(n_1784),
.B(n_1767),
.Y(n_1801)
);

AOI211xp5_ASAP7_75t_L g1802 ( 
.A1(n_1778),
.A2(n_1665),
.B(n_607),
.C(n_611),
.Y(n_1802)
);

AOI22xp33_ASAP7_75t_L g1803 ( 
.A1(n_1770),
.A2(n_1737),
.B1(n_1755),
.B2(n_1756),
.Y(n_1803)
);

INVx1_ASAP7_75t_L g1804 ( 
.A(n_1782),
.Y(n_1804)
);

INVx1_ASAP7_75t_L g1805 ( 
.A(n_1791),
.Y(n_1805)
);

INVx2_ASAP7_75t_L g1806 ( 
.A(n_1791),
.Y(n_1806)
);

AO31x2_ASAP7_75t_L g1807 ( 
.A1(n_1794),
.A2(n_1760),
.A3(n_1765),
.B(n_1736),
.Y(n_1807)
);

AND2x2_ASAP7_75t_L g1808 ( 
.A(n_1784),
.B(n_1736),
.Y(n_1808)
);

INVx1_ASAP7_75t_L g1809 ( 
.A(n_1789),
.Y(n_1809)
);

INVx2_ASAP7_75t_L g1810 ( 
.A(n_1789),
.Y(n_1810)
);

AND2x4_ASAP7_75t_L g1811 ( 
.A(n_1789),
.B(n_1756),
.Y(n_1811)
);

AND2x2_ASAP7_75t_L g1812 ( 
.A(n_1788),
.B(n_1736),
.Y(n_1812)
);

AND2x4_ASAP7_75t_SL g1813 ( 
.A(n_1788),
.B(n_1762),
.Y(n_1813)
);

HB1xp67_ASAP7_75t_L g1814 ( 
.A(n_1785),
.Y(n_1814)
);

AND2x2_ASAP7_75t_L g1815 ( 
.A(n_1788),
.B(n_1736),
.Y(n_1815)
);

HB1xp67_ASAP7_75t_L g1816 ( 
.A(n_1785),
.Y(n_1816)
);

INVx2_ASAP7_75t_L g1817 ( 
.A(n_1785),
.Y(n_1817)
);

NAND2xp5_ASAP7_75t_L g1818 ( 
.A(n_1790),
.B(n_1757),
.Y(n_1818)
);

INVx1_ASAP7_75t_L g1819 ( 
.A(n_1779),
.Y(n_1819)
);

NAND3xp33_ASAP7_75t_L g1820 ( 
.A(n_1772),
.B(n_1760),
.C(n_1764),
.Y(n_1820)
);

OR2x2_ASAP7_75t_L g1821 ( 
.A(n_1787),
.B(n_1748),
.Y(n_1821)
);

BUFx3_ASAP7_75t_L g1822 ( 
.A(n_1776),
.Y(n_1822)
);

OA21x2_ASAP7_75t_L g1823 ( 
.A1(n_1792),
.A2(n_1760),
.B(n_1735),
.Y(n_1823)
);

INVx1_ASAP7_75t_L g1824 ( 
.A(n_1793),
.Y(n_1824)
);

NAND2xp33_ASAP7_75t_L g1825 ( 
.A(n_1777),
.B(n_1765),
.Y(n_1825)
);

BUFx3_ASAP7_75t_L g1826 ( 
.A(n_1813),
.Y(n_1826)
);

INVx1_ASAP7_75t_L g1827 ( 
.A(n_1795),
.Y(n_1827)
);

NAND2xp5_ASAP7_75t_L g1828 ( 
.A(n_1803),
.B(n_1822),
.Y(n_1828)
);

INVx2_ASAP7_75t_L g1829 ( 
.A(n_1811),
.Y(n_1829)
);

AOI22xp33_ASAP7_75t_L g1830 ( 
.A1(n_1822),
.A2(n_1771),
.B1(n_1764),
.B2(n_1783),
.Y(n_1830)
);

OAI22xp33_ASAP7_75t_L g1831 ( 
.A1(n_1820),
.A2(n_1800),
.B1(n_1824),
.B2(n_1819),
.Y(n_1831)
);

OA211x2_ASAP7_75t_L g1832 ( 
.A1(n_1818),
.A2(n_1787),
.B(n_1781),
.C(n_1749),
.Y(n_1832)
);

OAI21xp33_ASAP7_75t_L g1833 ( 
.A1(n_1824),
.A2(n_1764),
.B(n_1756),
.Y(n_1833)
);

OAI33xp33_ASAP7_75t_L g1834 ( 
.A1(n_1796),
.A2(n_615),
.A3(n_612),
.B1(n_616),
.B2(n_613),
.B3(n_606),
.Y(n_1834)
);

OAI22xp5_ASAP7_75t_L g1835 ( 
.A1(n_1813),
.A2(n_1768),
.B1(n_1764),
.B2(n_1748),
.Y(n_1835)
);

AOI221xp5_ASAP7_75t_L g1836 ( 
.A1(n_1819),
.A2(n_619),
.B1(n_623),
.B2(n_618),
.C(n_617),
.Y(n_1836)
);

AOI22xp5_ASAP7_75t_L g1837 ( 
.A1(n_1825),
.A2(n_1737),
.B1(n_1764),
.B2(n_1761),
.Y(n_1837)
);

OAI22xp33_ASAP7_75t_L g1838 ( 
.A1(n_1821),
.A2(n_1766),
.B1(n_1757),
.B2(n_1749),
.Y(n_1838)
);

OAI31xp33_ASAP7_75t_L g1839 ( 
.A1(n_1821),
.A2(n_1761),
.A3(n_1742),
.B(n_1744),
.Y(n_1839)
);

AOI222xp33_ASAP7_75t_L g1840 ( 
.A1(n_1802),
.A2(n_625),
.B1(n_626),
.B2(n_1742),
.C1(n_763),
.C2(n_759),
.Y(n_1840)
);

OA222x2_ASAP7_75t_L g1841 ( 
.A1(n_1809),
.A2(n_1757),
.B1(n_1740),
.B2(n_1745),
.C1(n_1744),
.C2(n_1750),
.Y(n_1841)
);

INVx1_ASAP7_75t_L g1842 ( 
.A(n_1795),
.Y(n_1842)
);

INVx2_ASAP7_75t_L g1843 ( 
.A(n_1811),
.Y(n_1843)
);

INVx1_ASAP7_75t_SL g1844 ( 
.A(n_1796),
.Y(n_1844)
);

INVx2_ASAP7_75t_L g1845 ( 
.A(n_1811),
.Y(n_1845)
);

OAI21x1_ASAP7_75t_L g1846 ( 
.A1(n_1810),
.A2(n_1769),
.B(n_1735),
.Y(n_1846)
);

NAND3xp33_ASAP7_75t_L g1847 ( 
.A(n_1802),
.B(n_885),
.C(n_1742),
.Y(n_1847)
);

OR2x2_ASAP7_75t_L g1848 ( 
.A(n_1844),
.B(n_1809),
.Y(n_1848)
);

INVx1_ASAP7_75t_L g1849 ( 
.A(n_1827),
.Y(n_1849)
);

NAND2xp5_ASAP7_75t_L g1850 ( 
.A(n_1830),
.B(n_1810),
.Y(n_1850)
);

NAND2xp5_ASAP7_75t_L g1851 ( 
.A(n_1830),
.B(n_1801),
.Y(n_1851)
);

AND2x2_ASAP7_75t_L g1852 ( 
.A(n_1826),
.B(n_1812),
.Y(n_1852)
);

INVx1_ASAP7_75t_L g1853 ( 
.A(n_1842),
.Y(n_1853)
);

INVx2_ASAP7_75t_L g1854 ( 
.A(n_1829),
.Y(n_1854)
);

AND2x2_ASAP7_75t_L g1855 ( 
.A(n_1826),
.B(n_1812),
.Y(n_1855)
);

INVx2_ASAP7_75t_L g1856 ( 
.A(n_1843),
.Y(n_1856)
);

AND2x2_ASAP7_75t_L g1857 ( 
.A(n_1845),
.B(n_1815),
.Y(n_1857)
);

AND2x2_ASAP7_75t_L g1858 ( 
.A(n_1837),
.B(n_1815),
.Y(n_1858)
);

AND2x2_ASAP7_75t_L g1859 ( 
.A(n_1841),
.B(n_1811),
.Y(n_1859)
);

INVx2_ASAP7_75t_L g1860 ( 
.A(n_1846),
.Y(n_1860)
);

AND2x2_ASAP7_75t_L g1861 ( 
.A(n_1833),
.B(n_1801),
.Y(n_1861)
);

INVx1_ASAP7_75t_SL g1862 ( 
.A(n_1828),
.Y(n_1862)
);

INVx2_ASAP7_75t_L g1863 ( 
.A(n_1835),
.Y(n_1863)
);

AND2x2_ASAP7_75t_L g1864 ( 
.A(n_1839),
.B(n_1808),
.Y(n_1864)
);

INVx1_ASAP7_75t_L g1865 ( 
.A(n_1849),
.Y(n_1865)
);

AOI22xp5_ASAP7_75t_L g1866 ( 
.A1(n_1862),
.A2(n_1831),
.B1(n_1832),
.B2(n_1840),
.Y(n_1866)
);

INVx2_ASAP7_75t_L g1867 ( 
.A(n_1852),
.Y(n_1867)
);

INVx2_ASAP7_75t_SL g1868 ( 
.A(n_1852),
.Y(n_1868)
);

OAI211xp5_ASAP7_75t_L g1869 ( 
.A1(n_1851),
.A2(n_1847),
.B(n_1836),
.C(n_1831),
.Y(n_1869)
);

NAND2xp5_ASAP7_75t_L g1870 ( 
.A(n_1855),
.B(n_1838),
.Y(n_1870)
);

INVx1_ASAP7_75t_L g1871 ( 
.A(n_1853),
.Y(n_1871)
);

NAND2xp5_ASAP7_75t_L g1872 ( 
.A(n_1855),
.B(n_1838),
.Y(n_1872)
);

AOI221xp5_ASAP7_75t_L g1873 ( 
.A1(n_1850),
.A2(n_1834),
.B1(n_1816),
.B2(n_1814),
.C(n_1817),
.Y(n_1873)
);

AND2x4_ASAP7_75t_L g1874 ( 
.A(n_1868),
.B(n_1854),
.Y(n_1874)
);

AND2x2_ASAP7_75t_L g1875 ( 
.A(n_1867),
.B(n_1858),
.Y(n_1875)
);

INVx1_ASAP7_75t_L g1876 ( 
.A(n_1865),
.Y(n_1876)
);

NAND2xp5_ASAP7_75t_L g1877 ( 
.A(n_1866),
.B(n_1854),
.Y(n_1877)
);

AND2x2_ASAP7_75t_L g1878 ( 
.A(n_1870),
.B(n_1858),
.Y(n_1878)
);

INVx2_ASAP7_75t_L g1879 ( 
.A(n_1871),
.Y(n_1879)
);

INVx1_ASAP7_75t_L g1880 ( 
.A(n_1872),
.Y(n_1880)
);

NAND2xp5_ASAP7_75t_L g1881 ( 
.A(n_1874),
.B(n_1869),
.Y(n_1881)
);

NOR2xp33_ASAP7_75t_L g1882 ( 
.A(n_1877),
.B(n_1848),
.Y(n_1882)
);

NAND2xp5_ASAP7_75t_L g1883 ( 
.A(n_1874),
.B(n_1875),
.Y(n_1883)
);

AOI22xp5_ASAP7_75t_L g1884 ( 
.A1(n_1878),
.A2(n_1859),
.B1(n_1863),
.B2(n_1873),
.Y(n_1884)
);

AND2x2_ASAP7_75t_L g1885 ( 
.A(n_1875),
.B(n_1863),
.Y(n_1885)
);

INVx2_ASAP7_75t_SL g1886 ( 
.A(n_1883),
.Y(n_1886)
);

OR2x2_ASAP7_75t_L g1887 ( 
.A(n_1881),
.B(n_1880),
.Y(n_1887)
);

INVx1_ASAP7_75t_L g1888 ( 
.A(n_1885),
.Y(n_1888)
);

INVx1_ASAP7_75t_L g1889 ( 
.A(n_1888),
.Y(n_1889)
);

NAND2xp33_ASAP7_75t_SL g1890 ( 
.A(n_1886),
.B(n_1874),
.Y(n_1890)
);

OAI211xp5_ASAP7_75t_L g1891 ( 
.A1(n_1890),
.A2(n_1884),
.B(n_1882),
.C(n_1887),
.Y(n_1891)
);

INVx1_ASAP7_75t_L g1892 ( 
.A(n_1889),
.Y(n_1892)
);

INVx1_ASAP7_75t_L g1893 ( 
.A(n_1892),
.Y(n_1893)
);

NAND2xp5_ASAP7_75t_L g1894 ( 
.A(n_1891),
.B(n_1879),
.Y(n_1894)
);

AOI221xp5_ASAP7_75t_L g1895 ( 
.A1(n_1894),
.A2(n_1876),
.B1(n_1879),
.B2(n_1859),
.C(n_1856),
.Y(n_1895)
);

AOI211xp5_ASAP7_75t_L g1896 ( 
.A1(n_1893),
.A2(n_1856),
.B(n_1834),
.C(n_1864),
.Y(n_1896)
);

NAND2xp5_ASAP7_75t_L g1897 ( 
.A(n_1894),
.B(n_1857),
.Y(n_1897)
);

AO22x2_ASAP7_75t_L g1898 ( 
.A1(n_1897),
.A2(n_1860),
.B1(n_1857),
.B2(n_1864),
.Y(n_1898)
);

XOR2x2_ASAP7_75t_L g1899 ( 
.A(n_1895),
.B(n_1896),
.Y(n_1899)
);

INVx1_ASAP7_75t_L g1900 ( 
.A(n_1897),
.Y(n_1900)
);

OAI21xp33_ASAP7_75t_L g1901 ( 
.A1(n_1899),
.A2(n_1861),
.B(n_1804),
.Y(n_1901)
);

INVx1_ASAP7_75t_L g1902 ( 
.A(n_1898),
.Y(n_1902)
);

NOR2xp67_ASAP7_75t_L g1903 ( 
.A(n_1900),
.B(n_2),
.Y(n_1903)
);

INVx1_ASAP7_75t_L g1904 ( 
.A(n_1903),
.Y(n_1904)
);

AOI31xp33_ASAP7_75t_L g1905 ( 
.A1(n_1902),
.A2(n_1316),
.A3(n_659),
.B(n_660),
.Y(n_1905)
);

AOI22xp5_ASAP7_75t_L g1906 ( 
.A1(n_1901),
.A2(n_1823),
.B1(n_1806),
.B2(n_1805),
.Y(n_1906)
);

INVx2_ASAP7_75t_SL g1907 ( 
.A(n_1902),
.Y(n_1907)
);

AOI22xp5_ASAP7_75t_L g1908 ( 
.A1(n_1901),
.A2(n_1823),
.B1(n_1799),
.B2(n_1798),
.Y(n_1908)
);

AOI22xp5_ASAP7_75t_L g1909 ( 
.A1(n_1901),
.A2(n_1799),
.B1(n_1798),
.B2(n_1797),
.Y(n_1909)
);

NAND3x1_ASAP7_75t_SL g1910 ( 
.A(n_1905),
.B(n_723),
.C(n_0),
.Y(n_1910)
);

INVx1_ASAP7_75t_L g1911 ( 
.A(n_1908),
.Y(n_1911)
);

AND2x4_ASAP7_75t_L g1912 ( 
.A(n_1909),
.B(n_1807),
.Y(n_1912)
);

OAI21xp5_ASAP7_75t_L g1913 ( 
.A1(n_1906),
.A2(n_774),
.B(n_754),
.Y(n_1913)
);

NAND2xp33_ASAP7_75t_L g1914 ( 
.A(n_1904),
.B(n_1016),
.Y(n_1914)
);

NAND3xp33_ASAP7_75t_L g1915 ( 
.A(n_1907),
.B(n_777),
.C(n_775),
.Y(n_1915)
);

NAND3xp33_ASAP7_75t_L g1916 ( 
.A(n_1907),
.B(n_782),
.C(n_781),
.Y(n_1916)
);

NAND3xp33_ASAP7_75t_L g1917 ( 
.A(n_1907),
.B(n_785),
.C(n_784),
.Y(n_1917)
);

AND4x1_ASAP7_75t_L g1918 ( 
.A(n_1904),
.B(n_7),
.C(n_4),
.D(n_6),
.Y(n_1918)
);

NOR3xp33_ASAP7_75t_L g1919 ( 
.A(n_1907),
.B(n_976),
.C(n_769),
.Y(n_1919)
);

INVx2_ASAP7_75t_SL g1920 ( 
.A(n_1904),
.Y(n_1920)
);

NOR2x1_ASAP7_75t_L g1921 ( 
.A(n_1904),
.B(n_1239),
.Y(n_1921)
);

NAND2xp5_ASAP7_75t_L g1922 ( 
.A(n_1907),
.B(n_1807),
.Y(n_1922)
);

CKINVDCx5p33_ASAP7_75t_R g1923 ( 
.A(n_1904),
.Y(n_1923)
);

NOR3xp33_ASAP7_75t_L g1924 ( 
.A(n_1907),
.B(n_786),
.C(n_1009),
.Y(n_1924)
);

NOR3xp33_ASAP7_75t_L g1925 ( 
.A(n_1907),
.B(n_1013),
.C(n_1009),
.Y(n_1925)
);

NOR3xp33_ASAP7_75t_L g1926 ( 
.A(n_1907),
.B(n_1017),
.C(n_1014),
.Y(n_1926)
);

NOR2xp67_ASAP7_75t_L g1927 ( 
.A(n_1904),
.B(n_13),
.Y(n_1927)
);

OAI211xp5_ASAP7_75t_L g1928 ( 
.A1(n_1927),
.A2(n_368),
.B(n_369),
.C(n_366),
.Y(n_1928)
);

INVx1_ASAP7_75t_L g1929 ( 
.A(n_1918),
.Y(n_1929)
);

INVx1_ASAP7_75t_L g1930 ( 
.A(n_1910),
.Y(n_1930)
);

AO22x1_ASAP7_75t_L g1931 ( 
.A1(n_1921),
.A2(n_1364),
.B1(n_376),
.B2(n_377),
.Y(n_1931)
);

OAI21x1_ASAP7_75t_SL g1932 ( 
.A1(n_1913),
.A2(n_1358),
.B(n_1354),
.Y(n_1932)
);

XOR2xp5_ASAP7_75t_L g1933 ( 
.A(n_1915),
.B(n_21),
.Y(n_1933)
);

INVx1_ASAP7_75t_L g1934 ( 
.A(n_1916),
.Y(n_1934)
);

OAI221xp5_ASAP7_75t_SL g1935 ( 
.A1(n_1924),
.A2(n_27),
.B1(n_23),
.B2(n_25),
.C(n_28),
.Y(n_1935)
);

AOI221xp5_ASAP7_75t_L g1936 ( 
.A1(n_1919),
.A2(n_386),
.B1(n_387),
.B2(n_382),
.C(n_380),
.Y(n_1936)
);

AOI221xp5_ASAP7_75t_L g1937 ( 
.A1(n_1912),
.A2(n_578),
.B1(n_585),
.B2(n_576),
.C(n_571),
.Y(n_1937)
);

NAND2xp5_ASAP7_75t_L g1938 ( 
.A(n_1925),
.B(n_1926),
.Y(n_1938)
);

INVx1_ASAP7_75t_L g1939 ( 
.A(n_1917),
.Y(n_1939)
);

OR3x2_ASAP7_75t_L g1940 ( 
.A(n_1914),
.B(n_23),
.C(n_29),
.Y(n_1940)
);

OAI221xp5_ASAP7_75t_L g1941 ( 
.A1(n_1927),
.A2(n_635),
.B1(n_632),
.B2(n_631),
.C(n_1354),
.Y(n_1941)
);

OR2x2_ASAP7_75t_L g1942 ( 
.A(n_1920),
.B(n_41),
.Y(n_1942)
);

INVx1_ASAP7_75t_L g1943 ( 
.A(n_1927),
.Y(n_1943)
);

INVx1_ASAP7_75t_L g1944 ( 
.A(n_1927),
.Y(n_1944)
);

INVx1_ASAP7_75t_L g1945 ( 
.A(n_1927),
.Y(n_1945)
);

AND2x2_ASAP7_75t_L g1946 ( 
.A(n_1920),
.B(n_1759),
.Y(n_1946)
);

AND2x2_ASAP7_75t_L g1947 ( 
.A(n_1920),
.B(n_1759),
.Y(n_1947)
);

OAI211xp5_ASAP7_75t_SL g1948 ( 
.A1(n_1911),
.A2(n_45),
.B(n_42),
.C(n_43),
.Y(n_1948)
);

OAI22xp5_ASAP7_75t_L g1949 ( 
.A1(n_1923),
.A2(n_1753),
.B1(n_1751),
.B2(n_1752),
.Y(n_1949)
);

AND2x2_ASAP7_75t_L g1950 ( 
.A(n_1920),
.B(n_1752),
.Y(n_1950)
);

INVx1_ASAP7_75t_L g1951 ( 
.A(n_1927),
.Y(n_1951)
);

INVx1_ASAP7_75t_L g1952 ( 
.A(n_1927),
.Y(n_1952)
);

OAI211xp5_ASAP7_75t_L g1953 ( 
.A1(n_1927),
.A2(n_54),
.B(n_51),
.C(n_53),
.Y(n_1953)
);

INVx1_ASAP7_75t_L g1954 ( 
.A(n_1927),
.Y(n_1954)
);

NOR2xp67_ASAP7_75t_L g1955 ( 
.A(n_1927),
.B(n_56),
.Y(n_1955)
);

NOR2x1_ASAP7_75t_L g1956 ( 
.A(n_1927),
.B(n_57),
.Y(n_1956)
);

AOI211xp5_ASAP7_75t_L g1957 ( 
.A1(n_1927),
.A2(n_836),
.B(n_838),
.C(n_825),
.Y(n_1957)
);

O2A1O1Ixp5_ASAP7_75t_L g1958 ( 
.A1(n_1922),
.A2(n_838),
.B(n_853),
.C(n_825),
.Y(n_1958)
);

AOI211xp5_ASAP7_75t_L g1959 ( 
.A1(n_1927),
.A2(n_861),
.B(n_853),
.C(n_63),
.Y(n_1959)
);

NOR2xp67_ASAP7_75t_L g1960 ( 
.A(n_1927),
.B(n_62),
.Y(n_1960)
);

OAI221xp5_ASAP7_75t_L g1961 ( 
.A1(n_1927),
.A2(n_468),
.B1(n_469),
.B2(n_462),
.C(n_455),
.Y(n_1961)
);

NOR2xp67_ASAP7_75t_L g1962 ( 
.A(n_1927),
.B(n_66),
.Y(n_1962)
);

AND2x4_ASAP7_75t_L g1963 ( 
.A(n_1955),
.B(n_1960),
.Y(n_1963)
);

NAND2x1p5_ASAP7_75t_L g1964 ( 
.A(n_1956),
.B(n_1337),
.Y(n_1964)
);

NOR4xp25_ASAP7_75t_L g1965 ( 
.A(n_1928),
.B(n_1930),
.C(n_1929),
.D(n_1943),
.Y(n_1965)
);

HB1xp67_ASAP7_75t_L g1966 ( 
.A(n_1962),
.Y(n_1966)
);

NOR3xp33_ASAP7_75t_SL g1967 ( 
.A(n_1941),
.B(n_516),
.C(n_475),
.Y(n_1967)
);

INVx1_ASAP7_75t_SL g1968 ( 
.A(n_1942),
.Y(n_1968)
);

NAND3xp33_ASAP7_75t_SL g1969 ( 
.A(n_1959),
.B(n_520),
.C(n_519),
.Y(n_1969)
);

NAND2xp5_ASAP7_75t_L g1970 ( 
.A(n_1946),
.B(n_73),
.Y(n_1970)
);

NAND2xp5_ASAP7_75t_L g1971 ( 
.A(n_1947),
.B(n_75),
.Y(n_1971)
);

NAND4xp75_ASAP7_75t_L g1972 ( 
.A(n_1944),
.B(n_1951),
.C(n_1952),
.D(n_1945),
.Y(n_1972)
);

AOI211xp5_ASAP7_75t_L g1973 ( 
.A1(n_1948),
.A2(n_861),
.B(n_81),
.C(n_78),
.Y(n_1973)
);

AOI21x1_ASAP7_75t_L g1974 ( 
.A1(n_1931),
.A2(n_80),
.B(n_83),
.Y(n_1974)
);

NOR3xp33_ASAP7_75t_L g1975 ( 
.A(n_1954),
.B(n_534),
.C(n_533),
.Y(n_1975)
);

NOR3x1_ASAP7_75t_L g1976 ( 
.A(n_1953),
.B(n_88),
.C(n_89),
.Y(n_1976)
);

NOR3x1_ASAP7_75t_L g1977 ( 
.A(n_1961),
.B(n_90),
.C(n_92),
.Y(n_1977)
);

AOI211xp5_ASAP7_75t_L g1978 ( 
.A1(n_1935),
.A2(n_95),
.B(n_93),
.C(n_94),
.Y(n_1978)
);

OAI22xp5_ASAP7_75t_L g1979 ( 
.A1(n_1940),
.A2(n_563),
.B1(n_602),
.B2(n_556),
.Y(n_1979)
);

AND3x2_ASAP7_75t_L g1980 ( 
.A(n_1957),
.B(n_96),
.C(n_97),
.Y(n_1980)
);

OR2x2_ASAP7_75t_L g1981 ( 
.A(n_1950),
.B(n_101),
.Y(n_1981)
);

CKINVDCx20_ASAP7_75t_R g1982 ( 
.A(n_1933),
.Y(n_1982)
);

BUFx3_ASAP7_75t_L g1983 ( 
.A(n_1934),
.Y(n_1983)
);

INVxp33_ASAP7_75t_L g1984 ( 
.A(n_1938),
.Y(n_1984)
);

CKINVDCx5p33_ASAP7_75t_R g1985 ( 
.A(n_1939),
.Y(n_1985)
);

AOI222xp33_ASAP7_75t_L g1986 ( 
.A1(n_1937),
.A2(n_107),
.B1(n_110),
.B2(n_111),
.C1(n_112),
.C2(n_113),
.Y(n_1986)
);

NOR3xp33_ASAP7_75t_L g1987 ( 
.A(n_1936),
.B(n_115),
.C(n_116),
.Y(n_1987)
);

AOI222xp33_ASAP7_75t_L g1988 ( 
.A1(n_1932),
.A2(n_115),
.B1(n_116),
.B2(n_118),
.C1(n_119),
.C2(n_121),
.Y(n_1988)
);

INVx2_ASAP7_75t_L g1989 ( 
.A(n_1981),
.Y(n_1989)
);

NOR3xp33_ASAP7_75t_L g1990 ( 
.A(n_1972),
.B(n_1958),
.C(n_1949),
.Y(n_1990)
);

NAND3xp33_ASAP7_75t_L g1991 ( 
.A(n_1978),
.B(n_957),
.C(n_956),
.Y(n_1991)
);

NAND4xp25_ASAP7_75t_L g1992 ( 
.A(n_1976),
.B(n_129),
.C(n_125),
.D(n_127),
.Y(n_1992)
);

AND2x4_ASAP7_75t_L g1993 ( 
.A(n_1963),
.B(n_130),
.Y(n_1993)
);

AND4x1_ASAP7_75t_L g1994 ( 
.A(n_1965),
.B(n_134),
.C(n_132),
.D(n_133),
.Y(n_1994)
);

XNOR2xp5_ASAP7_75t_L g1995 ( 
.A(n_1982),
.B(n_135),
.Y(n_1995)
);

AND3x2_ASAP7_75t_L g1996 ( 
.A(n_1966),
.B(n_137),
.C(n_138),
.Y(n_1996)
);

INVxp33_ASAP7_75t_SL g1997 ( 
.A(n_1968),
.Y(n_1997)
);

INVx1_ASAP7_75t_L g1998 ( 
.A(n_1970),
.Y(n_1998)
);

NAND2xp5_ASAP7_75t_L g1999 ( 
.A(n_1980),
.B(n_143),
.Y(n_1999)
);

NAND4xp25_ASAP7_75t_L g2000 ( 
.A(n_1973),
.B(n_147),
.C(n_143),
.D(n_144),
.Y(n_2000)
);

BUFx2_ASAP7_75t_L g2001 ( 
.A(n_1964),
.Y(n_2001)
);

AND4x1_ASAP7_75t_L g2002 ( 
.A(n_1977),
.B(n_155),
.C(n_147),
.D(n_150),
.Y(n_2002)
);

NOR3xp33_ASAP7_75t_SL g2003 ( 
.A(n_1985),
.B(n_150),
.C(n_156),
.Y(n_2003)
);

XOR2xp5_ASAP7_75t_L g2004 ( 
.A(n_1984),
.B(n_1971),
.Y(n_2004)
);

NAND4xp25_ASAP7_75t_L g2005 ( 
.A(n_1988),
.B(n_159),
.C(n_157),
.D(n_158),
.Y(n_2005)
);

INVxp33_ASAP7_75t_L g2006 ( 
.A(n_1987),
.Y(n_2006)
);

AND3x2_ASAP7_75t_L g2007 ( 
.A(n_1975),
.B(n_157),
.C(n_159),
.Y(n_2007)
);

AOI22xp5_ASAP7_75t_L g2008 ( 
.A1(n_1983),
.A2(n_1667),
.B1(n_964),
.B2(n_971),
.Y(n_2008)
);

INVx3_ASAP7_75t_L g2009 ( 
.A(n_1974),
.Y(n_2009)
);

AND4x1_ASAP7_75t_L g2010 ( 
.A(n_1986),
.B(n_164),
.C(n_162),
.D(n_163),
.Y(n_2010)
);

XOR2xp5_ASAP7_75t_L g2011 ( 
.A(n_1969),
.B(n_1979),
.Y(n_2011)
);

XNOR2xp5_ASAP7_75t_L g2012 ( 
.A(n_1967),
.B(n_165),
.Y(n_2012)
);

NAND2xp5_ASAP7_75t_L g2013 ( 
.A(n_1996),
.B(n_1994),
.Y(n_2013)
);

AO22x2_ASAP7_75t_L g2014 ( 
.A1(n_2009),
.A2(n_169),
.B1(n_166),
.B2(n_167),
.Y(n_2014)
);

AND2x4_ASAP7_75t_L g2015 ( 
.A(n_1989),
.B(n_982),
.Y(n_2015)
);

NAND2xp5_ASAP7_75t_L g2016 ( 
.A(n_2002),
.B(n_171),
.Y(n_2016)
);

INVx2_ASAP7_75t_SL g2017 ( 
.A(n_1993),
.Y(n_2017)
);

INVx1_ASAP7_75t_L g2018 ( 
.A(n_1999),
.Y(n_2018)
);

NAND2xp5_ASAP7_75t_L g2019 ( 
.A(n_2007),
.B(n_176),
.Y(n_2019)
);

INVx1_ASAP7_75t_L g2020 ( 
.A(n_1995),
.Y(n_2020)
);

OA21x2_ASAP7_75t_L g2021 ( 
.A1(n_1998),
.A2(n_1264),
.B(n_1222),
.Y(n_2021)
);

AOI22xp5_ASAP7_75t_L g2022 ( 
.A1(n_2005),
.A2(n_1738),
.B1(n_1298),
.B2(n_1308),
.Y(n_2022)
);

INVx2_ASAP7_75t_L g2023 ( 
.A(n_2012),
.Y(n_2023)
);

OAI211xp5_ASAP7_75t_L g2024 ( 
.A1(n_2004),
.A2(n_2000),
.B(n_1990),
.C(n_2008),
.Y(n_2024)
);

NOR2x1_ASAP7_75t_L g2025 ( 
.A(n_1991),
.B(n_1264),
.Y(n_2025)
);

AOI21xp5_ASAP7_75t_L g2026 ( 
.A1(n_2006),
.A2(n_1136),
.B(n_1108),
.Y(n_2026)
);

OAI22xp5_ASAP7_75t_SL g2027 ( 
.A1(n_2001),
.A2(n_1136),
.B1(n_182),
.B2(n_183),
.Y(n_2027)
);

AOI22x1_ASAP7_75t_L g2028 ( 
.A1(n_2011),
.A2(n_181),
.B1(n_184),
.B2(n_186),
.Y(n_2028)
);

AOI22xp33_ASAP7_75t_SL g2029 ( 
.A1(n_1997),
.A2(n_1661),
.B1(n_856),
.B2(n_1738),
.Y(n_2029)
);

NAND2xp5_ASAP7_75t_L g2030 ( 
.A(n_1996),
.B(n_195),
.Y(n_2030)
);

AND2x2_ASAP7_75t_L g2031 ( 
.A(n_2003),
.B(n_1739),
.Y(n_2031)
);

OR2x2_ASAP7_75t_L g2032 ( 
.A(n_1992),
.B(n_208),
.Y(n_2032)
);

AOI211x1_ASAP7_75t_L g2033 ( 
.A1(n_2010),
.A2(n_1318),
.B(n_1323),
.C(n_1324),
.Y(n_2033)
);

NAND2xp5_ASAP7_75t_L g2034 ( 
.A(n_1996),
.B(n_209),
.Y(n_2034)
);

OAI221xp5_ASAP7_75t_L g2035 ( 
.A1(n_2030),
.A2(n_2034),
.B1(n_2019),
.B2(n_2017),
.C(n_2013),
.Y(n_2035)
);

INVx1_ASAP7_75t_L g2036 ( 
.A(n_2016),
.Y(n_2036)
);

NOR4xp25_ASAP7_75t_L g2037 ( 
.A(n_2024),
.B(n_236),
.C(n_240),
.D(n_242),
.Y(n_2037)
);

INVx1_ASAP7_75t_L g2038 ( 
.A(n_2032),
.Y(n_2038)
);

NAND2x1p5_ASAP7_75t_L g2039 ( 
.A(n_2020),
.B(n_1194),
.Y(n_2039)
);

AND2x4_ASAP7_75t_L g2040 ( 
.A(n_2018),
.B(n_265),
.Y(n_2040)
);

NAND2xp5_ASAP7_75t_L g2041 ( 
.A(n_2033),
.B(n_270),
.Y(n_2041)
);

NOR3xp33_ASAP7_75t_L g2042 ( 
.A(n_2023),
.B(n_1113),
.C(n_1221),
.Y(n_2042)
);

AND3x4_ASAP7_75t_L g2043 ( 
.A(n_2025),
.B(n_274),
.C(n_276),
.Y(n_2043)
);

INVx1_ASAP7_75t_L g2044 ( 
.A(n_2015),
.Y(n_2044)
);

INVx3_ASAP7_75t_L g2045 ( 
.A(n_2014),
.Y(n_2045)
);

AND2x4_ASAP7_75t_L g2046 ( 
.A(n_2031),
.B(n_299),
.Y(n_2046)
);

XNOR2xp5_ASAP7_75t_L g2047 ( 
.A(n_2028),
.B(n_307),
.Y(n_2047)
);

BUFx2_ASAP7_75t_SL g2048 ( 
.A(n_2045),
.Y(n_2048)
);

HB1xp67_ASAP7_75t_L g2049 ( 
.A(n_2043),
.Y(n_2049)
);

INVx3_ASAP7_75t_L g2050 ( 
.A(n_2046),
.Y(n_2050)
);

INVx2_ASAP7_75t_L g2051 ( 
.A(n_2040),
.Y(n_2051)
);

INVx1_ASAP7_75t_L g2052 ( 
.A(n_2041),
.Y(n_2052)
);

INVx1_ASAP7_75t_L g2053 ( 
.A(n_2047),
.Y(n_2053)
);

NAND2xp5_ASAP7_75t_L g2054 ( 
.A(n_2044),
.B(n_2021),
.Y(n_2054)
);

INVx1_ASAP7_75t_L g2055 ( 
.A(n_2039),
.Y(n_2055)
);

OR2x2_ASAP7_75t_L g2056 ( 
.A(n_2037),
.B(n_2021),
.Y(n_2056)
);

AND2x4_ASAP7_75t_L g2057 ( 
.A(n_2036),
.B(n_2022),
.Y(n_2057)
);

NOR2xp33_ASAP7_75t_R g2058 ( 
.A(n_2038),
.B(n_2014),
.Y(n_2058)
);

OAI22xp5_ASAP7_75t_L g2059 ( 
.A1(n_2035),
.A2(n_2026),
.B1(n_2027),
.B2(n_2029),
.Y(n_2059)
);

OR2x2_ASAP7_75t_SL g2060 ( 
.A(n_2056),
.B(n_2042),
.Y(n_2060)
);

NAND2xp5_ASAP7_75t_L g2061 ( 
.A(n_2048),
.B(n_311),
.Y(n_2061)
);

HB1xp67_ASAP7_75t_L g2062 ( 
.A(n_2058),
.Y(n_2062)
);

XNOR2xp5_ASAP7_75t_L g2063 ( 
.A(n_2049),
.B(n_319),
.Y(n_2063)
);

NAND3x1_ASAP7_75t_L g2064 ( 
.A(n_2050),
.B(n_326),
.C(n_333),
.Y(n_2064)
);

AOI22xp5_ASAP7_75t_L g2065 ( 
.A1(n_2052),
.A2(n_2051),
.B1(n_2053),
.B2(n_2057),
.Y(n_2065)
);

OAI22xp5_ASAP7_75t_SL g2066 ( 
.A1(n_2061),
.A2(n_2055),
.B1(n_2054),
.B2(n_2059),
.Y(n_2066)
);

CKINVDCx20_ASAP7_75t_R g2067 ( 
.A(n_2065),
.Y(n_2067)
);

INVx1_ASAP7_75t_SL g2068 ( 
.A(n_2062),
.Y(n_2068)
);

INVx2_ASAP7_75t_L g2069 ( 
.A(n_2064),
.Y(n_2069)
);

BUFx2_ASAP7_75t_L g2070 ( 
.A(n_2060),
.Y(n_2070)
);

NOR2xp67_ASAP7_75t_L g2071 ( 
.A(n_2069),
.B(n_2063),
.Y(n_2071)
);

INVxp67_ASAP7_75t_L g2072 ( 
.A(n_2070),
.Y(n_2072)
);

INVx1_ASAP7_75t_L g2073 ( 
.A(n_2067),
.Y(n_2073)
);

HB1xp67_ASAP7_75t_L g2074 ( 
.A(n_2068),
.Y(n_2074)
);

OAI22x1_ASAP7_75t_L g2075 ( 
.A1(n_2066),
.A2(n_1214),
.B1(n_1091),
.B2(n_1135),
.Y(n_2075)
);

AO21x2_ASAP7_75t_L g2076 ( 
.A1(n_2071),
.A2(n_1273),
.B(n_1265),
.Y(n_2076)
);

OAI22xp33_ASAP7_75t_L g2077 ( 
.A1(n_2072),
.A2(n_941),
.B1(n_938),
.B2(n_934),
.Y(n_2077)
);

INVx1_ASAP7_75t_L g2078 ( 
.A(n_2074),
.Y(n_2078)
);

AOI22xp5_ASAP7_75t_L g2079 ( 
.A1(n_2073),
.A2(n_1021),
.B1(n_938),
.B2(n_934),
.Y(n_2079)
);

HB1xp67_ASAP7_75t_L g2080 ( 
.A(n_2078),
.Y(n_2080)
);

INVx1_ASAP7_75t_L g2081 ( 
.A(n_2076),
.Y(n_2081)
);

HB1xp67_ASAP7_75t_L g2082 ( 
.A(n_2077),
.Y(n_2082)
);

AOI22xp33_ASAP7_75t_L g2083 ( 
.A1(n_2080),
.A2(n_2075),
.B1(n_2079),
.B2(n_934),
.Y(n_2083)
);

AOI22xp5_ASAP7_75t_L g2084 ( 
.A1(n_2081),
.A2(n_1137),
.B1(n_1157),
.B2(n_1155),
.Y(n_2084)
);

INVx1_ASAP7_75t_L g2085 ( 
.A(n_2082),
.Y(n_2085)
);

OAI31xp33_ASAP7_75t_L g2086 ( 
.A1(n_2085),
.A2(n_1137),
.A3(n_1157),
.B(n_1155),
.Y(n_2086)
);

OR2x6_ASAP7_75t_L g2087 ( 
.A(n_2083),
.B(n_1124),
.Y(n_2087)
);

XOR2xp5_ASAP7_75t_L g2088 ( 
.A(n_2084),
.B(n_1124),
.Y(n_2088)
);

OR2x2_ASAP7_75t_L g2089 ( 
.A(n_2087),
.B(n_1143),
.Y(n_2089)
);

AOI221xp5_ASAP7_75t_L g2090 ( 
.A1(n_2088),
.A2(n_1114),
.B1(n_1091),
.B2(n_1064),
.C(n_1072),
.Y(n_2090)
);

AOI21xp5_ASAP7_75t_L g2091 ( 
.A1(n_2089),
.A2(n_2090),
.B(n_2086),
.Y(n_2091)
);

AOI211xp5_ASAP7_75t_L g2092 ( 
.A1(n_2091),
.A2(n_1124),
.B(n_1156),
.C(n_1150),
.Y(n_2092)
);


endmodule