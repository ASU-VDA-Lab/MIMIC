module fake_jpeg_3061_n_555 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_555);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_555;

wire n_529;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx4_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_13),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_15),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

INVx11_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_6),
.Y(n_36)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_7),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_7),
.Y(n_38)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_14),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_3),
.Y(n_41)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_11),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_7),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_1),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_9),
.Y(n_45)
);

INVx1_ASAP7_75t_SL g46 ( 
.A(n_17),
.Y(n_46)
);

INVx1_ASAP7_75t_SL g47 ( 
.A(n_3),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_9),
.Y(n_48)
);

BUFx5_ASAP7_75t_L g49 ( 
.A(n_4),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_14),
.Y(n_50)
);

BUFx5_ASAP7_75t_L g51 ( 
.A(n_4),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_28),
.B(n_18),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_52),
.B(n_57),
.Y(n_113)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_28),
.Y(n_53)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_53),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_32),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_54),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_32),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_55),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_32),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_56),
.B(n_59),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_23),
.B(n_17),
.Y(n_57)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_58),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_23),
.B(n_18),
.Y(n_59)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_30),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_60),
.Y(n_148)
);

INVx4_ASAP7_75t_SL g61 ( 
.A(n_24),
.Y(n_61)
);

INVx5_ASAP7_75t_SL g125 ( 
.A(n_61),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_25),
.B(n_14),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_62),
.B(n_75),
.Y(n_136)
);

BUFx5_ASAP7_75t_L g63 ( 
.A(n_49),
.Y(n_63)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_63),
.Y(n_109)
);

BUFx12_ASAP7_75t_L g64 ( 
.A(n_24),
.Y(n_64)
);

BUFx12f_ASAP7_75t_L g142 ( 
.A(n_64),
.Y(n_142)
);

BUFx2_ASAP7_75t_L g65 ( 
.A(n_34),
.Y(n_65)
);

BUFx2_ASAP7_75t_L g146 ( 
.A(n_65),
.Y(n_146)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_34),
.Y(n_66)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_66),
.Y(n_124)
);

BUFx12f_ASAP7_75t_L g67 ( 
.A(n_34),
.Y(n_67)
);

INVx5_ASAP7_75t_L g110 ( 
.A(n_67),
.Y(n_110)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_37),
.Y(n_68)
);

INVx3_ASAP7_75t_L g167 ( 
.A(n_68),
.Y(n_167)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_24),
.Y(n_69)
);

INVx5_ASAP7_75t_L g160 ( 
.A(n_69),
.Y(n_160)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_37),
.Y(n_70)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_70),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_25),
.B(n_16),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_71),
.B(n_46),
.Y(n_144)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_19),
.Y(n_72)
);

INVx4_ASAP7_75t_L g123 ( 
.A(n_72),
.Y(n_123)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_22),
.Y(n_73)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_73),
.Y(n_115)
);

BUFx2_ASAP7_75t_L g74 ( 
.A(n_19),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g106 ( 
.A(n_74),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_32),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_30),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_76),
.Y(n_152)
);

INVx11_ASAP7_75t_L g77 ( 
.A(n_24),
.Y(n_77)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_77),
.Y(n_127)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_30),
.Y(n_78)
);

BUFx3_ASAP7_75t_L g150 ( 
.A(n_78),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_50),
.B(n_16),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_79),
.B(n_84),
.Y(n_151)
);

INVx8_ASAP7_75t_L g80 ( 
.A(n_24),
.Y(n_80)
);

INVx3_ASAP7_75t_SL g155 ( 
.A(n_80),
.Y(n_155)
);

BUFx5_ASAP7_75t_L g81 ( 
.A(n_49),
.Y(n_81)
);

INVx4_ASAP7_75t_L g147 ( 
.A(n_81),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_30),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_82),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_20),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_83),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_21),
.Y(n_84)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_51),
.Y(n_85)
);

INVx4_ASAP7_75t_L g140 ( 
.A(n_85),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_20),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_86),
.Y(n_161)
);

BUFx3_ASAP7_75t_L g87 ( 
.A(n_20),
.Y(n_87)
);

INVx4_ASAP7_75t_L g154 ( 
.A(n_87),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_44),
.Y(n_88)
);

INVx6_ASAP7_75t_L g114 ( 
.A(n_88),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_44),
.Y(n_89)
);

INVx6_ASAP7_75t_L g139 ( 
.A(n_89),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_44),
.Y(n_90)
);

INVx8_ASAP7_75t_L g119 ( 
.A(n_90),
.Y(n_119)
);

BUFx5_ASAP7_75t_L g91 ( 
.A(n_49),
.Y(n_91)
);

BUFx5_ASAP7_75t_L g116 ( 
.A(n_91),
.Y(n_116)
);

BUFx12f_ASAP7_75t_L g92 ( 
.A(n_39),
.Y(n_92)
);

INVx8_ASAP7_75t_L g130 ( 
.A(n_92),
.Y(n_130)
);

HB1xp67_ASAP7_75t_L g93 ( 
.A(n_19),
.Y(n_93)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_93),
.Y(n_129)
);

BUFx12f_ASAP7_75t_L g94 ( 
.A(n_39),
.Y(n_94)
);

INVx8_ASAP7_75t_L g138 ( 
.A(n_94),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_21),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_95),
.B(n_96),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_21),
.Y(n_96)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_39),
.Y(n_97)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_97),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_33),
.Y(n_98)
);

BUFx12f_ASAP7_75t_L g166 ( 
.A(n_98),
.Y(n_166)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_42),
.Y(n_99)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_99),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_33),
.Y(n_100)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_100),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_33),
.Y(n_101)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_101),
.Y(n_165)
);

INVx13_ASAP7_75t_L g102 ( 
.A(n_47),
.Y(n_102)
);

INVx6_ASAP7_75t_SL g105 ( 
.A(n_102),
.Y(n_105)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_42),
.Y(n_103)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_103),
.Y(n_120)
);

BUFx12f_ASAP7_75t_L g104 ( 
.A(n_42),
.Y(n_104)
);

BUFx12_ASAP7_75t_L g141 ( 
.A(n_104),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_61),
.A2(n_47),
.B1(n_46),
.B2(n_27),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g185 ( 
.A1(n_108),
.A2(n_134),
.B1(n_162),
.B2(n_77),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_65),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g203 ( 
.A(n_112),
.B(n_122),
.Y(n_203)
);

A2O1A1Ixp33_ASAP7_75t_L g117 ( 
.A1(n_102),
.A2(n_50),
.B(n_40),
.C(n_22),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_117),
.B(n_48),
.Y(n_186)
);

INVx6_ASAP7_75t_SL g121 ( 
.A(n_64),
.Y(n_121)
);

INVx13_ASAP7_75t_L g192 ( 
.A(n_121),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_74),
.Y(n_122)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_72),
.Y(n_131)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_131),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_85),
.A2(n_47),
.B1(n_46),
.B2(n_27),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_68),
.B(n_35),
.C(n_40),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_135),
.B(n_29),
.C(n_45),
.Y(n_168)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_58),
.Y(n_137)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_137),
.Y(n_175)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_60),
.Y(n_143)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_143),
.Y(n_204)
);

NAND3xp33_ASAP7_75t_L g217 ( 
.A(n_144),
.B(n_38),
.C(n_48),
.Y(n_217)
);

INVx6_ASAP7_75t_SL g145 ( 
.A(n_64),
.Y(n_145)
);

INVx13_ASAP7_75t_L g211 ( 
.A(n_145),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_98),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_156),
.B(n_163),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_SL g162 ( 
.A1(n_67),
.A2(n_27),
.B1(n_26),
.B2(n_35),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_100),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_92),
.B(n_26),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_164),
.B(n_26),
.Y(n_179)
);

AND2x2_ASAP7_75t_L g232 ( 
.A(n_168),
.B(n_224),
.Y(n_232)
);

BUFx5_ASAP7_75t_L g169 ( 
.A(n_105),
.Y(n_169)
);

INVx4_ASAP7_75t_L g243 ( 
.A(n_169),
.Y(n_243)
);

AOI21xp5_ASAP7_75t_L g170 ( 
.A1(n_108),
.A2(n_91),
.B(n_29),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_L g245 ( 
.A1(n_170),
.A2(n_199),
.B(n_209),
.Y(n_245)
);

CKINVDCx16_ASAP7_75t_R g172 ( 
.A(n_125),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_172),
.B(n_195),
.Y(n_264)
);

INVx4_ASAP7_75t_L g173 ( 
.A(n_160),
.Y(n_173)
);

INVx3_ASAP7_75t_L g262 ( 
.A(n_173),
.Y(n_262)
);

INVx4_ASAP7_75t_L g176 ( 
.A(n_154),
.Y(n_176)
);

INVx1_ASAP7_75t_SL g247 ( 
.A(n_176),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_115),
.B(n_104),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_SL g231 ( 
.A(n_177),
.B(n_190),
.Y(n_231)
);

BUFx3_ASAP7_75t_L g178 ( 
.A(n_110),
.Y(n_178)
);

BUFx3_ASAP7_75t_L g229 ( 
.A(n_178),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_179),
.B(n_191),
.Y(n_251)
);

INVx6_ASAP7_75t_L g180 ( 
.A(n_159),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g244 ( 
.A(n_180),
.Y(n_244)
);

INVx4_ASAP7_75t_L g181 ( 
.A(n_154),
.Y(n_181)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_181),
.Y(n_235)
);

INVx5_ASAP7_75t_L g182 ( 
.A(n_130),
.Y(n_182)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_182),
.Y(n_261)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_129),
.Y(n_183)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_183),
.Y(n_273)
);

INVx6_ASAP7_75t_L g184 ( 
.A(n_159),
.Y(n_184)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_184),
.Y(n_274)
);

INVxp67_ASAP7_75t_L g238 ( 
.A(n_185),
.Y(n_238)
);

CKINVDCx14_ASAP7_75t_R g260 ( 
.A(n_186),
.Y(n_260)
);

AND2x2_ASAP7_75t_L g187 ( 
.A(n_113),
.B(n_67),
.Y(n_187)
);

CKINVDCx16_ASAP7_75t_R g271 ( 
.A(n_187),
.Y(n_271)
);

AOI22xp33_ASAP7_75t_SL g188 ( 
.A1(n_109),
.A2(n_104),
.B1(n_94),
.B2(n_92),
.Y(n_188)
);

AOI22xp33_ASAP7_75t_SL g266 ( 
.A1(n_188),
.A2(n_127),
.B1(n_138),
.B2(n_166),
.Y(n_266)
);

BUFx12f_ASAP7_75t_L g189 ( 
.A(n_141),
.Y(n_189)
);

INVx13_ASAP7_75t_L g275 ( 
.A(n_189),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_126),
.B(n_94),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_136),
.B(n_151),
.Y(n_191)
);

INVx11_ASAP7_75t_L g193 ( 
.A(n_166),
.Y(n_193)
);

INVxp67_ASAP7_75t_L g277 ( 
.A(n_193),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_157),
.B(n_80),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_194),
.B(n_197),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_107),
.B(n_31),
.Y(n_195)
);

BUFx12f_ASAP7_75t_L g196 ( 
.A(n_141),
.Y(n_196)
);

INVx6_ASAP7_75t_L g254 ( 
.A(n_196),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_120),
.B(n_69),
.Y(n_197)
);

OR2x2_ASAP7_75t_L g198 ( 
.A(n_125),
.B(n_45),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g268 ( 
.A(n_198),
.B(n_219),
.Y(n_268)
);

AOI21xp5_ASAP7_75t_L g199 ( 
.A1(n_134),
.A2(n_31),
.B(n_51),
.Y(n_199)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_133),
.Y(n_200)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_200),
.Y(n_239)
);

AND2x2_ASAP7_75t_L g201 ( 
.A(n_128),
.B(n_78),
.Y(n_201)
);

CKINVDCx16_ASAP7_75t_R g279 ( 
.A(n_201),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_149),
.B(n_140),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_202),
.B(n_217),
.Y(n_278)
);

INVx2_ASAP7_75t_SL g205 ( 
.A(n_146),
.Y(n_205)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_205),
.Y(n_236)
);

INVx4_ASAP7_75t_L g206 ( 
.A(n_130),
.Y(n_206)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_206),
.Y(n_241)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_124),
.Y(n_207)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_207),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_158),
.A2(n_54),
.B1(n_55),
.B2(n_89),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g252 ( 
.A1(n_208),
.A2(n_114),
.B1(n_139),
.B2(n_153),
.Y(n_252)
);

AOI21xp5_ASAP7_75t_L g209 ( 
.A1(n_162),
.A2(n_51),
.B(n_36),
.Y(n_209)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_167),
.Y(n_210)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_210),
.Y(n_248)
);

CKINVDCx16_ASAP7_75t_R g212 ( 
.A(n_146),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g281 ( 
.A(n_212),
.B(n_222),
.Y(n_281)
);

INVx3_ASAP7_75t_L g213 ( 
.A(n_106),
.Y(n_213)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_213),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_118),
.B(n_87),
.C(n_101),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_214),
.B(n_215),
.C(n_147),
.Y(n_259)
);

AND2x2_ASAP7_75t_SL g215 ( 
.A(n_140),
.B(n_82),
.Y(n_215)
);

INVx13_ASAP7_75t_L g216 ( 
.A(n_142),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_216),
.Y(n_249)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_165),
.Y(n_218)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_218),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_123),
.B(n_36),
.Y(n_219)
);

INVx3_ASAP7_75t_L g220 ( 
.A(n_106),
.Y(n_220)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_220),
.Y(n_267)
);

INVx6_ASAP7_75t_L g221 ( 
.A(n_161),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_221),
.Y(n_263)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_155),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_155),
.B(n_43),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_223),
.B(n_227),
.Y(n_237)
);

INVx5_ASAP7_75t_L g224 ( 
.A(n_138),
.Y(n_224)
);

CKINVDCx12_ASAP7_75t_R g225 ( 
.A(n_142),
.Y(n_225)
);

AND2x2_ASAP7_75t_L g242 ( 
.A(n_225),
.B(n_226),
.Y(n_242)
);

INVx2_ASAP7_75t_SL g226 ( 
.A(n_150),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_111),
.B(n_43),
.Y(n_227)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_114),
.Y(n_228)
);

AND2x2_ASAP7_75t_L g280 ( 
.A(n_228),
.B(n_0),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_185),
.A2(n_86),
.B1(n_83),
.B2(n_88),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g319 ( 
.A1(n_230),
.A2(n_270),
.B1(n_276),
.B2(n_0),
.Y(n_319)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_209),
.A2(n_148),
.B1(n_90),
.B2(n_161),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_L g316 ( 
.A1(n_233),
.A2(n_234),
.B1(n_250),
.B2(n_196),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_199),
.A2(n_148),
.B1(n_76),
.B2(n_152),
.Y(n_234)
);

A2O1A1Ixp33_ASAP7_75t_L g240 ( 
.A1(n_187),
.A2(n_41),
.B(n_38),
.C(n_116),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_L g283 ( 
.A1(n_240),
.A2(n_203),
.B(n_192),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_170),
.A2(n_153),
.B1(n_152),
.B2(n_111),
.Y(n_250)
);

AOI22xp33_ASAP7_75t_L g330 ( 
.A1(n_252),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_330)
);

AND2x2_ASAP7_75t_SL g253 ( 
.A(n_168),
.B(n_142),
.Y(n_253)
);

INVx1_ASAP7_75t_SL g315 ( 
.A(n_253),
.Y(n_315)
);

AOI22xp33_ASAP7_75t_L g255 ( 
.A1(n_171),
.A2(n_41),
.B1(n_132),
.B2(n_150),
.Y(n_255)
);

OAI22xp33_ASAP7_75t_SL g321 ( 
.A1(n_255),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_321)
);

AND2x2_ASAP7_75t_L g289 ( 
.A(n_259),
.B(n_265),
.Y(n_289)
);

AO22x2_ASAP7_75t_L g265 ( 
.A1(n_215),
.A2(n_127),
.B1(n_119),
.B2(n_166),
.Y(n_265)
);

INVxp67_ASAP7_75t_L g310 ( 
.A(n_266),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_215),
.B(n_139),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_269),
.B(n_173),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_L g270 ( 
.A1(n_208),
.A2(n_119),
.B1(n_132),
.B2(n_16),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_SL g272 ( 
.A(n_214),
.B(n_12),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_272),
.B(n_196),
.C(n_1),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_L g276 ( 
.A1(n_198),
.A2(n_12),
.B1(n_11),
.B2(n_10),
.Y(n_276)
);

AND2x2_ASAP7_75t_L g300 ( 
.A(n_280),
.B(n_206),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_238),
.A2(n_228),
.B1(n_201),
.B2(n_188),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_282),
.B(n_291),
.Y(n_331)
);

INVxp33_ASAP7_75t_SL g340 ( 
.A(n_283),
.Y(n_340)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_242),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g355 ( 
.A(n_284),
.B(n_285),
.Y(n_355)
);

AND2x6_ASAP7_75t_L g285 ( 
.A(n_253),
.B(n_192),
.Y(n_285)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_274),
.Y(n_286)
);

INVx2_ASAP7_75t_L g333 ( 
.A(n_286),
.Y(n_333)
);

CKINVDCx12_ASAP7_75t_R g287 ( 
.A(n_242),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_SL g342 ( 
.A(n_287),
.B(n_297),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_SL g288 ( 
.A(n_268),
.B(n_174),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_SL g339 ( 
.A(n_288),
.B(n_290),
.Y(n_339)
);

CKINVDCx16_ASAP7_75t_R g290 ( 
.A(n_242),
.Y(n_290)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_274),
.Y(n_292)
);

INVx2_ASAP7_75t_L g369 ( 
.A(n_292),
.Y(n_369)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_236),
.Y(n_293)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_293),
.Y(n_351)
);

AND2x2_ASAP7_75t_SL g294 ( 
.A(n_232),
.B(n_204),
.Y(n_294)
);

INVx1_ASAP7_75t_SL g361 ( 
.A(n_294),
.Y(n_361)
);

OAI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_238),
.A2(n_180),
.B1(n_221),
.B2(n_184),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_295),
.B(n_302),
.Y(n_338)
);

OAI21xp5_ASAP7_75t_L g296 ( 
.A1(n_245),
.A2(n_175),
.B(n_226),
.Y(n_296)
);

OAI21xp5_ASAP7_75t_SL g336 ( 
.A1(n_296),
.A2(n_234),
.B(n_250),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_231),
.B(n_205),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_SL g298 ( 
.A(n_251),
.B(n_176),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g356 ( 
.A(n_298),
.B(n_301),
.Y(n_356)
);

CKINVDCx10_ASAP7_75t_R g299 ( 
.A(n_275),
.Y(n_299)
);

INVx1_ASAP7_75t_SL g365 ( 
.A(n_299),
.Y(n_365)
);

INVx1_ASAP7_75t_SL g370 ( 
.A(n_300),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_256),
.B(n_264),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_272),
.B(n_181),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_278),
.B(n_220),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_SL g371 ( 
.A(n_303),
.B(n_313),
.Y(n_371)
);

XNOR2xp5_ASAP7_75t_L g304 ( 
.A(n_253),
.B(n_232),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_304),
.B(n_329),
.C(n_267),
.Y(n_347)
);

AND2x6_ASAP7_75t_L g305 ( 
.A(n_260),
.B(n_211),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_305),
.B(n_307),
.Y(n_345)
);

OR2x2_ASAP7_75t_L g306 ( 
.A(n_245),
.B(n_211),
.Y(n_306)
);

OAI21xp5_ASAP7_75t_L g353 ( 
.A1(n_306),
.A2(n_277),
.B(n_247),
.Y(n_353)
);

OAI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_233),
.A2(n_213),
.B1(n_224),
.B2(n_182),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_236),
.Y(n_308)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_308),
.Y(n_358)
);

AOI21xp5_ASAP7_75t_L g309 ( 
.A1(n_240),
.A2(n_169),
.B(n_216),
.Y(n_309)
);

AOI21xp5_ASAP7_75t_L g344 ( 
.A1(n_309),
.A2(n_322),
.B(n_280),
.Y(n_344)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_246),
.Y(n_311)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_311),
.Y(n_360)
);

AOI22xp33_ASAP7_75t_SL g312 ( 
.A1(n_230),
.A2(n_193),
.B1(n_178),
.B2(n_189),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_L g332 ( 
.A1(n_312),
.A2(n_319),
.B1(n_328),
.B2(n_330),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_237),
.B(n_189),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_232),
.B(n_0),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_314),
.B(n_317),
.Y(n_346)
);

AOI22xp33_ASAP7_75t_L g335 ( 
.A1(n_316),
.A2(n_321),
.B1(n_269),
.B2(n_279),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_281),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_SL g318 ( 
.A(n_237),
.B(n_12),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_318),
.B(n_327),
.Y(n_348)
);

XNOR2xp5_ASAP7_75t_SL g373 ( 
.A(n_320),
.B(n_235),
.Y(n_373)
);

AOI21xp5_ASAP7_75t_L g322 ( 
.A1(n_259),
.A2(n_1),
.B(n_3),
.Y(n_322)
);

CKINVDCx12_ASAP7_75t_R g323 ( 
.A(n_275),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_323),
.Y(n_334)
);

INVx4_ASAP7_75t_L g324 ( 
.A(n_262),
.Y(n_324)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_324),
.Y(n_359)
);

INVx5_ASAP7_75t_L g325 ( 
.A(n_244),
.Y(n_325)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_325),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_249),
.B(n_3),
.Y(n_326)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_326),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_243),
.B(n_4),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_243),
.B(n_4),
.Y(n_328)
);

XNOR2xp5_ASAP7_75t_L g329 ( 
.A(n_271),
.B(n_5),
.Y(n_329)
);

INVxp33_ASAP7_75t_L g401 ( 
.A(n_335),
.Y(n_401)
);

OAI21xp5_ASAP7_75t_SL g385 ( 
.A1(n_336),
.A2(n_354),
.B(n_362),
.Y(n_385)
);

OAI22xp5_ASAP7_75t_L g337 ( 
.A1(n_316),
.A2(n_317),
.B1(n_283),
.B2(n_319),
.Y(n_337)
);

AOI22xp5_ASAP7_75t_SL g382 ( 
.A1(n_337),
.A2(n_298),
.B1(n_282),
.B2(n_295),
.Y(n_382)
);

XNOR2xp5_ASAP7_75t_L g341 ( 
.A(n_304),
.B(n_239),
.Y(n_341)
);

MAJIxp5_ASAP7_75t_L g380 ( 
.A(n_341),
.B(n_349),
.C(n_352),
.Y(n_380)
);

OAI22xp5_ASAP7_75t_SL g343 ( 
.A1(n_289),
.A2(n_265),
.B1(n_263),
.B2(n_280),
.Y(n_343)
);

AOI22xp5_ASAP7_75t_L g404 ( 
.A1(n_343),
.A2(n_350),
.B1(n_372),
.B2(n_292),
.Y(n_404)
);

INVx1_ASAP7_75t_SL g383 ( 
.A(n_344),
.Y(n_383)
);

XNOR2xp5_ASAP7_75t_L g375 ( 
.A(n_347),
.B(n_294),
.Y(n_375)
);

XNOR2xp5_ASAP7_75t_L g349 ( 
.A(n_315),
.B(n_246),
.Y(n_349)
);

OAI22xp5_ASAP7_75t_SL g350 ( 
.A1(n_289),
.A2(n_265),
.B1(n_244),
.B2(n_241),
.Y(n_350)
);

XOR2xp5_ASAP7_75t_L g352 ( 
.A(n_315),
.B(n_265),
.Y(n_352)
);

AOI21xp5_ASAP7_75t_SL g393 ( 
.A1(n_353),
.A2(n_364),
.B(n_367),
.Y(n_393)
);

OAI21xp5_ASAP7_75t_L g354 ( 
.A1(n_306),
.A2(n_296),
.B(n_309),
.Y(n_354)
);

MAJIxp5_ASAP7_75t_L g357 ( 
.A(n_289),
.B(n_248),
.C(n_258),
.Y(n_357)
);

MAJIxp5_ASAP7_75t_L g384 ( 
.A(n_357),
.B(n_293),
.C(n_308),
.Y(n_384)
);

OAI21xp5_ASAP7_75t_SL g362 ( 
.A1(n_306),
.A2(n_257),
.B(n_267),
.Y(n_362)
);

OA22x2_ASAP7_75t_L g363 ( 
.A1(n_285),
.A2(n_261),
.B1(n_262),
.B2(n_257),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_363),
.B(n_307),
.Y(n_379)
);

OAI21xp5_ASAP7_75t_SL g364 ( 
.A1(n_302),
.A2(n_261),
.B(n_247),
.Y(n_364)
);

OAI21xp5_ASAP7_75t_L g367 ( 
.A1(n_284),
.A2(n_248),
.B(n_277),
.Y(n_367)
);

OAI22xp5_ASAP7_75t_SL g372 ( 
.A1(n_294),
.A2(n_258),
.B1(n_273),
.B2(n_235),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_SL g394 ( 
.A(n_373),
.B(n_329),
.Y(n_394)
);

CKINVDCx20_ASAP7_75t_R g374 ( 
.A(n_334),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_374),
.Y(n_410)
);

XOR2xp5_ASAP7_75t_L g431 ( 
.A(n_375),
.B(n_394),
.Y(n_431)
);

OAI22xp5_ASAP7_75t_SL g376 ( 
.A1(n_331),
.A2(n_291),
.B1(n_310),
.B2(n_314),
.Y(n_376)
);

AOI22xp5_ASAP7_75t_L g418 ( 
.A1(n_376),
.A2(n_381),
.B1(n_361),
.B2(n_343),
.Y(n_418)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_351),
.Y(n_377)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_377),
.Y(n_413)
);

CKINVDCx20_ASAP7_75t_R g378 ( 
.A(n_367),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_378),
.Y(n_412)
);

AOI22xp33_ASAP7_75t_L g421 ( 
.A1(n_379),
.A2(n_407),
.B1(n_408),
.B2(n_338),
.Y(n_421)
);

OAI22xp5_ASAP7_75t_SL g381 ( 
.A1(n_331),
.A2(n_310),
.B1(n_322),
.B2(n_290),
.Y(n_381)
);

OAI22xp5_ASAP7_75t_L g414 ( 
.A1(n_382),
.A2(n_404),
.B1(n_379),
.B2(n_338),
.Y(n_414)
);

MAJIxp5_ASAP7_75t_L g416 ( 
.A(n_384),
.B(n_395),
.C(n_397),
.Y(n_416)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_358),
.Y(n_386)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_386),
.Y(n_422)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_360),
.Y(n_387)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_387),
.Y(n_425)
);

AND2x6_ASAP7_75t_L g388 ( 
.A(n_355),
.B(n_305),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_388),
.B(n_391),
.Y(n_426)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_333),
.Y(n_389)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_389),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_346),
.B(n_300),
.Y(n_390)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_390),
.Y(n_411)
);

INVxp67_ASAP7_75t_L g391 ( 
.A(n_353),
.Y(n_391)
);

NOR2xp33_ASAP7_75t_L g392 ( 
.A(n_342),
.B(n_288),
.Y(n_392)
);

NOR2xp33_ASAP7_75t_SL g434 ( 
.A(n_392),
.B(n_403),
.Y(n_434)
);

XNOR2xp5_ASAP7_75t_L g395 ( 
.A(n_341),
.B(n_320),
.Y(n_395)
);

CKINVDCx16_ASAP7_75t_R g396 ( 
.A(n_371),
.Y(n_396)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_396),
.Y(n_437)
);

XNOR2xp5_ASAP7_75t_L g397 ( 
.A(n_347),
.B(n_300),
.Y(n_397)
);

CKINVDCx20_ASAP7_75t_R g398 ( 
.A(n_356),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_L g423 ( 
.A(n_398),
.B(n_400),
.Y(n_423)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_333),
.Y(n_399)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_399),
.Y(n_427)
);

MAJIxp5_ASAP7_75t_L g400 ( 
.A(n_357),
.B(n_311),
.C(n_273),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_346),
.B(n_318),
.Y(n_402)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_402),
.Y(n_432)
);

CKINVDCx20_ASAP7_75t_R g403 ( 
.A(n_372),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_SL g405 ( 
.A(n_339),
.B(n_299),
.Y(n_405)
);

OR2x2_ASAP7_75t_L g419 ( 
.A(n_405),
.B(n_406),
.Y(n_419)
);

NOR2xp33_ASAP7_75t_L g406 ( 
.A(n_368),
.B(n_229),
.Y(n_406)
);

CKINVDCx20_ASAP7_75t_R g407 ( 
.A(n_363),
.Y(n_407)
);

CKINVDCx20_ASAP7_75t_R g408 ( 
.A(n_363),
.Y(n_408)
);

AOI22xp5_ASAP7_75t_SL g409 ( 
.A1(n_350),
.A2(n_324),
.B1(n_325),
.B2(n_286),
.Y(n_409)
);

AND2x2_ASAP7_75t_L g420 ( 
.A(n_409),
.B(n_332),
.Y(n_420)
);

OAI22xp5_ASAP7_75t_L g442 ( 
.A1(n_414),
.A2(n_418),
.B1(n_430),
.B2(n_438),
.Y(n_442)
);

INVx1_ASAP7_75t_SL g415 ( 
.A(n_389),
.Y(n_415)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_415),
.Y(n_456)
);

INVxp67_ASAP7_75t_L g417 ( 
.A(n_385),
.Y(n_417)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_417),
.Y(n_448)
);

HB1xp67_ASAP7_75t_L g458 ( 
.A(n_420),
.Y(n_458)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_421),
.Y(n_444)
);

BUFx2_ASAP7_75t_L g424 ( 
.A(n_409),
.Y(n_424)
);

CKINVDCx14_ASAP7_75t_R g443 ( 
.A(n_424),
.Y(n_443)
);

OAI22xp5_ASAP7_75t_SL g428 ( 
.A1(n_382),
.A2(n_345),
.B1(n_354),
.B2(n_340),
.Y(n_428)
);

AOI22xp5_ASAP7_75t_L g464 ( 
.A1(n_428),
.A2(n_366),
.B1(n_365),
.B2(n_369),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_390),
.B(n_345),
.Y(n_429)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_429),
.Y(n_453)
);

AOI22xp5_ASAP7_75t_SL g430 ( 
.A1(n_383),
.A2(n_361),
.B1(n_370),
.B2(n_363),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_402),
.B(n_404),
.Y(n_435)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_435),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_384),
.B(n_362),
.Y(n_436)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_436),
.Y(n_466)
);

AOI22xp5_ASAP7_75t_L g438 ( 
.A1(n_401),
.A2(n_352),
.B1(n_344),
.B2(n_336),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_400),
.B(n_364),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_439),
.B(n_440),
.Y(n_445)
);

INVx2_ASAP7_75t_SL g440 ( 
.A(n_399),
.Y(n_440)
);

AOI22xp33_ASAP7_75t_L g441 ( 
.A1(n_401),
.A2(n_370),
.B1(n_348),
.B2(n_359),
.Y(n_441)
);

OAI22xp5_ASAP7_75t_L g450 ( 
.A1(n_441),
.A2(n_393),
.B1(n_391),
.B2(n_383),
.Y(n_450)
);

OA21x2_ASAP7_75t_L g446 ( 
.A1(n_428),
.A2(n_393),
.B(n_385),
.Y(n_446)
);

OAI21xp5_ASAP7_75t_SL g482 ( 
.A1(n_446),
.A2(n_454),
.B(n_412),
.Y(n_482)
);

XNOR2xp5_ASAP7_75t_L g447 ( 
.A(n_416),
.B(n_397),
.Y(n_447)
);

XNOR2xp5_ASAP7_75t_L g486 ( 
.A(n_447),
.B(n_455),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_432),
.B(n_376),
.Y(n_449)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_449),
.Y(n_477)
);

OAI22xp5_ASAP7_75t_L g478 ( 
.A1(n_450),
.A2(n_464),
.B1(n_465),
.B2(n_424),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_432),
.B(n_387),
.Y(n_451)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_451),
.Y(n_484)
);

MAJIxp5_ASAP7_75t_L g452 ( 
.A(n_416),
.B(n_431),
.C(n_436),
.Y(n_452)
);

MAJIxp5_ASAP7_75t_L g472 ( 
.A(n_452),
.B(n_455),
.C(n_457),
.Y(n_472)
);

AOI21xp5_ASAP7_75t_L g454 ( 
.A1(n_417),
.A2(n_381),
.B(n_388),
.Y(n_454)
);

MAJIxp5_ASAP7_75t_L g455 ( 
.A(n_431),
.B(n_380),
.C(n_375),
.Y(n_455)
);

MAJIxp5_ASAP7_75t_L g457 ( 
.A(n_423),
.B(n_380),
.C(n_395),
.Y(n_457)
);

MAJIxp5_ASAP7_75t_L g459 ( 
.A(n_439),
.B(n_373),
.C(n_349),
.Y(n_459)
);

MAJIxp5_ASAP7_75t_L g476 ( 
.A(n_459),
.B(n_460),
.C(n_462),
.Y(n_476)
);

MAJIxp5_ASAP7_75t_L g460 ( 
.A(n_411),
.B(n_386),
.C(n_377),
.Y(n_460)
);

MAJIxp5_ASAP7_75t_L g462 ( 
.A(n_411),
.B(n_359),
.C(n_366),
.Y(n_462)
);

NOR2xp33_ASAP7_75t_L g463 ( 
.A(n_410),
.B(n_348),
.Y(n_463)
);

NOR2xp33_ASAP7_75t_SL g485 ( 
.A(n_463),
.B(n_467),
.Y(n_485)
);

OAI22xp5_ASAP7_75t_L g465 ( 
.A1(n_434),
.A2(n_365),
.B1(n_369),
.B2(n_254),
.Y(n_465)
);

CKINVDCx20_ASAP7_75t_R g467 ( 
.A(n_410),
.Y(n_467)
);

CKINVDCx16_ASAP7_75t_R g468 ( 
.A(n_419),
.Y(n_468)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_468),
.Y(n_487)
);

OAI22xp5_ASAP7_75t_L g469 ( 
.A1(n_444),
.A2(n_435),
.B1(n_426),
.B2(n_418),
.Y(n_469)
);

OAI22xp5_ASAP7_75t_L g494 ( 
.A1(n_469),
.A2(n_475),
.B1(n_483),
.B2(n_464),
.Y(n_494)
);

AOI21xp5_ASAP7_75t_L g470 ( 
.A1(n_454),
.A2(n_426),
.B(n_444),
.Y(n_470)
);

AOI21xp5_ASAP7_75t_L g497 ( 
.A1(n_470),
.A2(n_482),
.B(n_442),
.Y(n_497)
);

OAI22xp5_ASAP7_75t_SL g471 ( 
.A1(n_461),
.A2(n_438),
.B1(n_429),
.B2(n_420),
.Y(n_471)
);

AOI22xp5_ASAP7_75t_L g503 ( 
.A1(n_471),
.A2(n_458),
.B1(n_449),
.B2(n_453),
.Y(n_503)
);

INVx11_ASAP7_75t_L g473 ( 
.A(n_443),
.Y(n_473)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_473),
.Y(n_507)
);

OAI21xp5_ASAP7_75t_L g474 ( 
.A1(n_446),
.A2(n_430),
.B(n_412),
.Y(n_474)
);

OAI21xp5_ASAP7_75t_L g504 ( 
.A1(n_474),
.A2(n_448),
.B(n_453),
.Y(n_504)
);

CKINVDCx14_ASAP7_75t_R g475 ( 
.A(n_451),
.Y(n_475)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_478),
.Y(n_493)
);

MAJIxp5_ASAP7_75t_L g479 ( 
.A(n_447),
.B(n_420),
.C(n_415),
.Y(n_479)
);

MAJIxp5_ASAP7_75t_L g492 ( 
.A(n_479),
.B(n_481),
.C(n_488),
.Y(n_492)
);

INVx2_ASAP7_75t_L g480 ( 
.A(n_456),
.Y(n_480)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_480),
.Y(n_498)
);

MAJIxp5_ASAP7_75t_L g481 ( 
.A(n_452),
.B(n_440),
.C(n_427),
.Y(n_481)
);

CKINVDCx20_ASAP7_75t_R g483 ( 
.A(n_445),
.Y(n_483)
);

HB1xp67_ASAP7_75t_L g509 ( 
.A(n_486),
.Y(n_509)
);

MAJIxp5_ASAP7_75t_L g488 ( 
.A(n_457),
.B(n_440),
.C(n_427),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_460),
.Y(n_489)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_489),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_445),
.B(n_419),
.Y(n_490)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_490),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_461),
.B(n_433),
.Y(n_491)
);

CKINVDCx16_ASAP7_75t_R g505 ( 
.A(n_491),
.Y(n_505)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_494),
.Y(n_514)
);

NOR2xp33_ASAP7_75t_L g495 ( 
.A(n_485),
.B(n_437),
.Y(n_495)
);

AOI22xp5_ASAP7_75t_L g512 ( 
.A1(n_495),
.A2(n_487),
.B1(n_489),
.B2(n_485),
.Y(n_512)
);

MAJIxp5_ASAP7_75t_L g496 ( 
.A(n_476),
.B(n_466),
.C(n_462),
.Y(n_496)
);

MAJIxp5_ASAP7_75t_L g513 ( 
.A(n_496),
.B(n_508),
.C(n_472),
.Y(n_513)
);

OAI21xp5_ASAP7_75t_L g510 ( 
.A1(n_497),
.A2(n_504),
.B(n_506),
.Y(n_510)
);

NOR2xp33_ASAP7_75t_SL g499 ( 
.A(n_487),
.B(n_466),
.Y(n_499)
);

NOR2xp33_ASAP7_75t_L g519 ( 
.A(n_499),
.B(n_413),
.Y(n_519)
);

XOR2xp5_ASAP7_75t_L g500 ( 
.A(n_479),
.B(n_446),
.Y(n_500)
);

XNOR2xp5_ASAP7_75t_L g515 ( 
.A(n_500),
.B(n_474),
.Y(n_515)
);

OAI22xp5_ASAP7_75t_SL g520 ( 
.A1(n_503),
.A2(n_483),
.B1(n_484),
.B2(n_477),
.Y(n_520)
);

OAI21xp5_ASAP7_75t_L g506 ( 
.A1(n_482),
.A2(n_448),
.B(n_459),
.Y(n_506)
);

MAJIxp5_ASAP7_75t_L g508 ( 
.A(n_476),
.B(n_425),
.C(n_422),
.Y(n_508)
);

MAJIxp5_ASAP7_75t_SL g511 ( 
.A(n_501),
.B(n_472),
.C(n_486),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_511),
.B(n_517),
.Y(n_530)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_512),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_SL g531 ( 
.A(n_513),
.B(n_518),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_515),
.B(n_516),
.Y(n_525)
);

XOR2xp5_ASAP7_75t_L g516 ( 
.A(n_500),
.B(n_481),
.Y(n_516)
);

AOI22xp5_ASAP7_75t_L g517 ( 
.A1(n_493),
.A2(n_490),
.B1(n_469),
.B2(n_484),
.Y(n_517)
);

MAJIxp5_ASAP7_75t_L g518 ( 
.A(n_492),
.B(n_488),
.C(n_470),
.Y(n_518)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_519),
.Y(n_534)
);

AOI22xp5_ASAP7_75t_L g526 ( 
.A1(n_520),
.A2(n_523),
.B1(n_504),
.B2(n_505),
.Y(n_526)
);

BUFx24_ASAP7_75t_SL g521 ( 
.A(n_501),
.Y(n_521)
);

NOR2xp33_ASAP7_75t_L g528 ( 
.A(n_521),
.B(n_522),
.Y(n_528)
);

AOI22xp5_ASAP7_75t_L g522 ( 
.A1(n_493),
.A2(n_477),
.B1(n_471),
.B2(n_480),
.Y(n_522)
);

OAI22xp5_ASAP7_75t_L g523 ( 
.A1(n_502),
.A2(n_473),
.B1(n_491),
.B2(n_254),
.Y(n_523)
);

MAJIxp5_ASAP7_75t_L g524 ( 
.A(n_492),
.B(n_229),
.C(n_6),
.Y(n_524)
);

MAJIxp5_ASAP7_75t_L g532 ( 
.A(n_524),
.B(n_506),
.C(n_508),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_L g538 ( 
.A(n_526),
.B(n_527),
.Y(n_538)
);

CKINVDCx20_ASAP7_75t_R g527 ( 
.A(n_510),
.Y(n_527)
);

NOR2xp33_ASAP7_75t_L g541 ( 
.A(n_532),
.B(n_524),
.Y(n_541)
);

AOI22xp5_ASAP7_75t_L g533 ( 
.A1(n_514),
.A2(n_502),
.B1(n_497),
.B2(n_503),
.Y(n_533)
);

AND2x2_ASAP7_75t_L g536 ( 
.A(n_533),
.B(n_535),
.Y(n_536)
);

AOI22xp5_ASAP7_75t_L g535 ( 
.A1(n_510),
.A2(n_498),
.B1(n_507),
.B2(n_496),
.Y(n_535)
);

NOR2xp33_ASAP7_75t_L g537 ( 
.A(n_534),
.B(n_498),
.Y(n_537)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_537),
.Y(n_543)
);

AOI21xp5_ASAP7_75t_L g539 ( 
.A1(n_530),
.A2(n_513),
.B(n_518),
.Y(n_539)
);

OAI21xp5_ASAP7_75t_L g545 ( 
.A1(n_539),
.A2(n_540),
.B(n_525),
.Y(n_545)
);

AOI21xp5_ASAP7_75t_SL g540 ( 
.A1(n_531),
.A2(n_509),
.B(n_516),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_L g546 ( 
.A(n_541),
.B(n_542),
.Y(n_546)
);

MAJIxp5_ASAP7_75t_L g542 ( 
.A(n_525),
.B(n_515),
.C(n_8),
.Y(n_542)
);

NOR2xp33_ASAP7_75t_L g544 ( 
.A(n_537),
.B(n_535),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_L g548 ( 
.A(n_544),
.B(n_528),
.Y(n_548)
);

AOI21xp5_ASAP7_75t_L g547 ( 
.A1(n_545),
.A2(n_538),
.B(n_536),
.Y(n_547)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_547),
.Y(n_550)
);

NOR2xp33_ASAP7_75t_L g549 ( 
.A(n_548),
.B(n_543),
.Y(n_549)
);

MAJIxp5_ASAP7_75t_L g551 ( 
.A(n_549),
.B(n_546),
.C(n_529),
.Y(n_551)
);

MAJIxp5_ASAP7_75t_L g552 ( 
.A(n_551),
.B(n_550),
.C(n_533),
.Y(n_552)
);

NOR3xp33_ASAP7_75t_L g553 ( 
.A(n_552),
.B(n_532),
.C(n_526),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_553),
.B(n_9),
.Y(n_554)
);

OAI22xp5_ASAP7_75t_L g555 ( 
.A1(n_554),
.A2(n_5),
.B1(n_8),
.B2(n_9),
.Y(n_555)
);


endmodule