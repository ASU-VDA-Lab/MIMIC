module fake_jpeg_1338_n_181 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_181);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_181;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_93;
wire n_54;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g45 ( 
.A(n_11),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_32),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_43),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_16),
.Y(n_49)
);

INVx8_ASAP7_75t_SL g50 ( 
.A(n_19),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_25),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_9),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_26),
.Y(n_53)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_34),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_15),
.Y(n_55)
);

INVx13_ASAP7_75t_L g56 ( 
.A(n_29),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_13),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_15),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_7),
.Y(n_59)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_11),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_18),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_9),
.Y(n_62)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_41),
.Y(n_63)
);

INVx11_ASAP7_75t_L g64 ( 
.A(n_50),
.Y(n_64)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_64),
.Y(n_73)
);

INVx11_ASAP7_75t_L g65 ( 
.A(n_56),
.Y(n_65)
);

BUFx8_ASAP7_75t_L g83 ( 
.A(n_65),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_53),
.Y(n_66)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_66),
.Y(n_79)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_60),
.Y(n_67)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_67),
.Y(n_81)
);

BUFx12f_ASAP7_75t_L g68 ( 
.A(n_56),
.Y(n_68)
);

INVx5_ASAP7_75t_L g75 ( 
.A(n_68),
.Y(n_75)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_63),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_69),
.B(n_71),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_53),
.Y(n_70)
);

INVx5_ASAP7_75t_L g80 ( 
.A(n_70),
.Y(n_80)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_60),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_67),
.A2(n_52),
.B1(n_57),
.B2(n_45),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_72),
.A2(n_74),
.B1(n_68),
.B2(n_64),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_71),
.A2(n_52),
.B1(n_57),
.B2(n_45),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_69),
.A2(n_66),
.B1(n_70),
.B2(n_63),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_77),
.A2(n_79),
.B1(n_76),
.B2(n_80),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_71),
.B(n_58),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_78),
.B(n_51),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_70),
.B(n_46),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_82),
.B(n_61),
.Y(n_86)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_81),
.Y(n_84)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_84),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_82),
.B(n_46),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_85),
.B(n_86),
.Y(n_102)
);

OAI22xp33_ASAP7_75t_L g87 ( 
.A1(n_81),
.A2(n_66),
.B1(n_65),
.B2(n_59),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_87),
.A2(n_89),
.B1(n_92),
.B2(n_94),
.Y(n_103)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_79),
.Y(n_88)
);

INVx4_ASAP7_75t_L g115 ( 
.A(n_88),
.Y(n_115)
);

OAI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_76),
.A2(n_66),
.B1(n_65),
.B2(n_64),
.Y(n_89)
);

OA22x2_ASAP7_75t_L g109 ( 
.A1(n_90),
.A2(n_95),
.B1(n_96),
.B2(n_68),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_91),
.B(n_0),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_78),
.B(n_47),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_93),
.B(n_98),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_77),
.A2(n_59),
.B1(n_48),
.B2(n_47),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_L g95 ( 
.A1(n_80),
.A2(n_55),
.B1(n_49),
.B2(n_62),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_75),
.A2(n_55),
.B1(n_49),
.B2(n_48),
.Y(n_96)
);

A2O1A1Ixp33_ASAP7_75t_L g97 ( 
.A1(n_83),
.A2(n_68),
.B(n_1),
.C(n_2),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_97),
.B(n_99),
.Y(n_107)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_73),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_83),
.Y(n_99)
);

BUFx2_ASAP7_75t_L g100 ( 
.A(n_75),
.Y(n_100)
);

CKINVDCx16_ASAP7_75t_R g114 ( 
.A(n_100),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_100),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_101),
.B(n_110),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_92),
.A2(n_61),
.B1(n_73),
.B2(n_83),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_105),
.A2(n_120),
.B1(n_33),
.B2(n_42),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_85),
.B(n_73),
.C(n_83),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_106),
.B(n_111),
.C(n_28),
.Y(n_123)
);

NOR2x1_ASAP7_75t_L g108 ( 
.A(n_96),
.B(n_68),
.Y(n_108)
);

CKINVDCx16_ASAP7_75t_R g131 ( 
.A(n_108),
.Y(n_131)
);

CKINVDCx16_ASAP7_75t_R g134 ( 
.A(n_109),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_L g111 ( 
.A(n_94),
.B(n_54),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_88),
.B(n_0),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_112),
.B(n_116),
.Y(n_126)
);

OAI32xp33_ASAP7_75t_L g113 ( 
.A1(n_97),
.A2(n_54),
.A3(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_113),
.B(n_8),
.Y(n_124)
);

CKINVDCx16_ASAP7_75t_R g116 ( 
.A(n_98),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_87),
.B(n_1),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_117),
.B(n_119),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_85),
.B(n_3),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_92),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_104),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_121),
.B(n_124),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_103),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_122),
.A2(n_129),
.B1(n_136),
.B2(n_22),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_123),
.B(n_132),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_115),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_128),
.B(n_135),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_103),
.A2(n_8),
.B1(n_10),
.B2(n_12),
.Y(n_129)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_118),
.Y(n_130)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_130),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g132 ( 
.A(n_102),
.B(n_30),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_115),
.Y(n_133)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_133),
.Y(n_154)
);

CKINVDCx16_ASAP7_75t_R g135 ( 
.A(n_108),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_107),
.A2(n_10),
.B1(n_12),
.B2(n_13),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_137),
.A2(n_17),
.B1(n_20),
.B2(n_21),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_106),
.B(n_31),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_138),
.B(n_24),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_109),
.A2(n_14),
.B1(n_16),
.B2(n_17),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_139),
.Y(n_151)
);

AOI322xp5_ASAP7_75t_L g140 ( 
.A1(n_124),
.A2(n_120),
.A3(n_111),
.B1(n_109),
.B2(n_105),
.C1(n_114),
.C2(n_23),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_140),
.B(n_141),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g141 ( 
.A(n_125),
.B(n_14),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_143),
.A2(n_145),
.B1(n_147),
.B2(n_37),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_126),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_146),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_134),
.A2(n_131),
.B1(n_127),
.B2(n_122),
.Y(n_147)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_148),
.Y(n_155)
);

AOI21xp5_ASAP7_75t_L g149 ( 
.A1(n_138),
.A2(n_44),
.B(n_36),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_L g161 ( 
.A1(n_149),
.A2(n_38),
.B(n_39),
.Y(n_161)
);

HB1xp67_ASAP7_75t_L g152 ( 
.A(n_133),
.Y(n_152)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_152),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_153),
.B(n_123),
.C(n_132),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_156),
.B(n_157),
.C(n_161),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_153),
.B(n_136),
.C(n_129),
.Y(n_157)
);

XOR2xp5_ASAP7_75t_L g158 ( 
.A(n_150),
.B(n_27),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_SL g165 ( 
.A(n_158),
.B(n_149),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_159),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_156),
.B(n_148),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_164),
.B(n_165),
.C(n_168),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_155),
.B(n_144),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_162),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_169),
.B(n_163),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_170),
.B(n_172),
.Y(n_173)
);

NOR3xp33_ASAP7_75t_L g172 ( 
.A(n_166),
.B(n_142),
.C(n_151),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_171),
.B(n_167),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_SL g175 ( 
.A(n_174),
.B(n_157),
.Y(n_175)
);

AOI21xp5_ASAP7_75t_L g176 ( 
.A1(n_175),
.A2(n_174),
.B(n_173),
.Y(n_176)
);

AOI21xp5_ASAP7_75t_L g177 ( 
.A1(n_176),
.A2(n_158),
.B(n_160),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_177),
.B(n_165),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_178),
.B(n_151),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_179),
.B(n_145),
.C(n_154),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_180),
.B(n_40),
.Y(n_181)
);


endmodule