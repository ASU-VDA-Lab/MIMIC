module fake_jpeg_13362_n_132 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_132);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_132;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

INVx2_ASAP7_75t_L g14 ( 
.A(n_4),
.Y(n_14)
);

BUFx2_ASAP7_75t_L g15 ( 
.A(n_9),
.Y(n_15)
);

BUFx12_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_2),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

INVx5_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_11),
.B(n_3),
.Y(n_20)
);

BUFx16f_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_11),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_8),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_10),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_28),
.Y(n_29)
);

HB1xp67_ASAP7_75t_L g55 ( 
.A(n_29),
.Y(n_55)
);

INVx2_ASAP7_75t_SL g30 ( 
.A(n_19),
.Y(n_30)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_30),
.Y(n_46)
);

BUFx10_ASAP7_75t_L g31 ( 
.A(n_21),
.Y(n_31)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_31),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_20),
.B(n_1),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_SL g43 ( 
.A(n_32),
.B(n_17),
.Y(n_43)
);

INVx5_ASAP7_75t_L g33 ( 
.A(n_28),
.Y(n_33)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_33),
.Y(n_48)
);

A2O1A1Ixp33_ASAP7_75t_L g34 ( 
.A1(n_20),
.A2(n_1),
.B(n_2),
.C(n_3),
.Y(n_34)
);

NOR2x1_ASAP7_75t_L g60 ( 
.A(n_34),
.B(n_18),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g35 ( 
.A1(n_14),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_35),
.A2(n_36),
.B1(n_17),
.B2(n_19),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_L g36 ( 
.A1(n_15),
.A2(n_13),
.B1(n_6),
.B2(n_7),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_16),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_37),
.B(n_21),
.Y(n_47)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_15),
.Y(n_38)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_23),
.B(n_25),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_39),
.B(n_41),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_22),
.Y(n_40)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_23),
.B(n_5),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_15),
.Y(n_42)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_43),
.B(n_47),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_32),
.B(n_14),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_44),
.B(n_61),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_37),
.B(n_25),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_49),
.B(n_53),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_50),
.A2(n_26),
.B1(n_30),
.B2(n_27),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g52 ( 
.A(n_29),
.B(n_18),
.Y(n_52)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_52),
.B(n_62),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g53 ( 
.A(n_34),
.B(n_24),
.Y(n_53)
);

MAJIxp5_ASAP7_75t_L g56 ( 
.A(n_38),
.B(n_26),
.C(n_22),
.Y(n_56)
);

FAx1_ASAP7_75t_SL g67 ( 
.A(n_56),
.B(n_31),
.CI(n_62),
.CON(n_67),
.SN(n_67)
);

NOR2xp33_ASAP7_75t_SL g59 ( 
.A(n_31),
.B(n_24),
.Y(n_59)
);

OR2x2_ASAP7_75t_L g79 ( 
.A(n_59),
.B(n_60),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_35),
.B(n_18),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_42),
.B(n_18),
.Y(n_62)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_51),
.Y(n_64)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_64),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_61),
.A2(n_53),
.B1(n_44),
.B2(n_60),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_65),
.A2(n_70),
.B1(n_72),
.B2(n_75),
.Y(n_89)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_51),
.Y(n_66)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_66),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_67),
.B(n_77),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_55),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_68),
.B(n_54),
.Y(n_90)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_58),
.Y(n_69)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_69),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_56),
.A2(n_33),
.B1(n_30),
.B2(n_40),
.Y(n_72)
);

OAI21xp5_ASAP7_75t_SL g73 ( 
.A1(n_52),
.A2(n_31),
.B(n_27),
.Y(n_73)
);

AOI21xp5_ASAP7_75t_L g93 ( 
.A1(n_73),
.A2(n_76),
.B(n_57),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_52),
.A2(n_40),
.B1(n_21),
.B2(n_16),
.Y(n_75)
);

OAI21xp5_ASAP7_75t_SL g76 ( 
.A1(n_58),
.A2(n_16),
.B(n_40),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_46),
.A2(n_16),
.B1(n_7),
.B2(n_12),
.Y(n_77)
);

INVxp67_ASAP7_75t_L g80 ( 
.A(n_76),
.Y(n_80)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_80),
.Y(n_95)
);

XOR2xp5_ASAP7_75t_L g83 ( 
.A(n_63),
.B(n_74),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_83),
.B(n_87),
.C(n_69),
.Y(n_101)
);

CKINVDCx14_ASAP7_75t_R g85 ( 
.A(n_71),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_SL g100 ( 
.A1(n_85),
.A2(n_88),
.B(n_70),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_63),
.B(n_46),
.C(n_54),
.Y(n_87)
);

OR2x2_ASAP7_75t_L g88 ( 
.A(n_73),
.B(n_43),
.Y(n_88)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_90),
.Y(n_102)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_64),
.Y(n_91)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_91),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_67),
.B(n_45),
.Y(n_92)
);

XNOR2xp5_ASAP7_75t_SL g94 ( 
.A(n_92),
.B(n_78),
.Y(n_94)
);

A2O1A1Ixp33_ASAP7_75t_SL g97 ( 
.A1(n_93),
.A2(n_67),
.B(n_72),
.C(n_79),
.Y(n_97)
);

XNOR2xp5_ASAP7_75t_SL g107 ( 
.A(n_94),
.B(n_101),
.Y(n_107)
);

AOI21xp5_ASAP7_75t_L g96 ( 
.A1(n_80),
.A2(n_79),
.B(n_74),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_96),
.B(n_86),
.C(n_88),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_97),
.A2(n_86),
.B1(n_87),
.B2(n_89),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_82),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_98),
.B(n_100),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_L g99 ( 
.A1(n_92),
.A2(n_74),
.B(n_66),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_99),
.B(n_104),
.C(n_93),
.Y(n_106)
);

XNOR2xp5_ASAP7_75t_SL g104 ( 
.A(n_83),
.B(n_77),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_103),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_105),
.B(n_111),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_106),
.B(n_109),
.C(n_110),
.Y(n_117)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_102),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_101),
.B(n_91),
.C(n_82),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_112),
.B(n_97),
.C(n_99),
.Y(n_119)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_95),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_113),
.B(n_84),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_114),
.B(n_118),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g115 ( 
.A(n_108),
.B(n_94),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_115),
.B(n_116),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_107),
.B(n_104),
.Y(n_116)
);

BUFx24_ASAP7_75t_SL g118 ( 
.A(n_107),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_119),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_L g123 ( 
.A1(n_117),
.A2(n_106),
.B(n_97),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_123),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_120),
.A2(n_97),
.B1(n_84),
.B2(n_81),
.Y(n_124)
);

OR2x2_ASAP7_75t_L g128 ( 
.A(n_124),
.B(n_75),
.Y(n_128)
);

AOI31xp67_ASAP7_75t_L g126 ( 
.A1(n_125),
.A2(n_122),
.A3(n_121),
.B(n_81),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_126),
.B(n_122),
.C(n_57),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_128),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_130),
.A2(n_127),
.B1(n_48),
.B2(n_13),
.Y(n_131)
);

A2O1A1O1Ixp25_ASAP7_75t_L g132 ( 
.A1(n_131),
.A2(n_129),
.B(n_12),
.C(n_6),
.D(n_48),
.Y(n_132)
);


endmodule