module fake_jpeg_5538_n_342 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_342);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_342;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g16 ( 
.A(n_15),
.Y(n_16)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_9),
.Y(n_18)
);

INVxp67_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_6),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_13),
.Y(n_25)
);

INVx13_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

INVxp67_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_13),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_15),
.Y(n_34)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_22),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_35),
.B(n_36),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_25),
.Y(n_36)
);

INVx11_ASAP7_75t_L g37 ( 
.A(n_20),
.Y(n_37)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_37),
.Y(n_60)
);

INVx3_ASAP7_75t_SL g38 ( 
.A(n_30),
.Y(n_38)
);

HB1xp67_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_22),
.Y(n_39)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_22),
.Y(n_41)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_30),
.Y(n_42)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

INVx11_ASAP7_75t_L g43 ( 
.A(n_20),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_43),
.A2(n_44),
.B1(n_46),
.B2(n_47),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_25),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_17),
.Y(n_45)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_45),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g46 ( 
.A(n_18),
.B(n_0),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_23),
.B(n_0),
.Y(n_47)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_38),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_48),
.B(n_50),
.Y(n_73)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_51),
.B(n_53),
.Y(n_80)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_54),
.B(n_55),
.Y(n_82)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_42),
.A2(n_17),
.B1(n_31),
.B2(n_32),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_59),
.A2(n_64),
.B1(n_69),
.B2(n_70),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_42),
.A2(n_17),
.B1(n_31),
.B2(n_32),
.Y(n_64)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_39),
.Y(n_65)
);

INVx6_ASAP7_75t_L g96 ( 
.A(n_65),
.Y(n_96)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_35),
.Y(n_66)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_66),
.Y(n_78)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_45),
.Y(n_67)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_67),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_L g68 ( 
.A1(n_36),
.A2(n_31),
.B1(n_33),
.B2(n_34),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_68),
.A2(n_34),
.B1(n_33),
.B2(n_36),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_42),
.A2(n_31),
.B1(n_32),
.B2(n_16),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_42),
.A2(n_16),
.B1(n_18),
.B2(n_21),
.Y(n_70)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_45),
.Y(n_71)
);

INVx1_ASAP7_75t_SL g90 ( 
.A(n_71),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_61),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_72),
.B(n_83),
.Y(n_110)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_63),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_74),
.B(n_77),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_49),
.B(n_46),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_75),
.B(n_76),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_61),
.B(n_46),
.Y(n_76)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_63),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_58),
.B(n_41),
.C(n_45),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_79),
.B(n_104),
.C(n_53),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_58),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_84),
.A2(n_23),
.B1(n_27),
.B2(n_47),
.Y(n_107)
);

A2O1A1Ixp33_ASAP7_75t_L g86 ( 
.A1(n_71),
.A2(n_44),
.B(n_46),
.C(n_28),
.Y(n_86)
);

AOI21xp5_ASAP7_75t_L g119 ( 
.A1(n_86),
.A2(n_97),
.B(n_19),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_60),
.Y(n_87)
);

BUFx3_ASAP7_75t_L g116 ( 
.A(n_87),
.Y(n_116)
);

CKINVDCx16_ASAP7_75t_R g88 ( 
.A(n_57),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_88),
.B(n_91),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_52),
.B(n_46),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_89),
.B(n_92),
.Y(n_113)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_55),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_52),
.B(n_46),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_L g93 ( 
.A1(n_60),
.A2(n_43),
.B1(n_37),
.B2(n_44),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_93),
.A2(n_98),
.B1(n_43),
.B2(n_62),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_67),
.B(n_47),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_94),
.B(n_27),
.Y(n_124)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_54),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_95),
.B(n_99),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_48),
.A2(n_35),
.B1(n_16),
.B2(n_37),
.Y(n_97)
);

OAI22xp33_ASAP7_75t_L g98 ( 
.A1(n_60),
.A2(n_37),
.B1(n_43),
.B2(n_35),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_50),
.B(n_21),
.Y(n_99)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_65),
.Y(n_100)
);

INVx5_ASAP7_75t_SL g129 ( 
.A(n_100),
.Y(n_129)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_55),
.Y(n_101)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_101),
.Y(n_128)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_62),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_102),
.Y(n_112)
);

INVx1_ASAP7_75t_SL g103 ( 
.A(n_57),
.Y(n_103)
);

CKINVDCx14_ASAP7_75t_R g126 ( 
.A(n_103),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_51),
.B(n_41),
.C(n_35),
.Y(n_104)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_105),
.B(n_109),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_107),
.A2(n_29),
.B1(n_24),
.B2(n_87),
.Y(n_159)
);

CKINVDCx16_ASAP7_75t_R g108 ( 
.A(n_82),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_108),
.B(n_111),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g109 ( 
.A(n_75),
.B(n_92),
.Y(n_109)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_84),
.Y(n_111)
);

OAI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_114),
.A2(n_74),
.B1(n_77),
.B2(n_88),
.Y(n_136)
);

INVx13_ASAP7_75t_L g115 ( 
.A(n_78),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_115),
.B(n_118),
.Y(n_156)
);

OAI32xp33_ASAP7_75t_L g117 ( 
.A1(n_89),
.A2(n_27),
.A3(n_23),
.B1(n_62),
.B2(n_40),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_117),
.B(n_124),
.Y(n_157)
);

OA21x2_ASAP7_75t_L g118 ( 
.A1(n_73),
.A2(n_40),
.B(n_66),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_L g138 ( 
.A1(n_119),
.A2(n_102),
.B1(n_96),
.B2(n_100),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_85),
.A2(n_72),
.B1(n_86),
.B2(n_76),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_121),
.A2(n_132),
.B1(n_95),
.B2(n_90),
.Y(n_146)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_94),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_122),
.B(n_123),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_83),
.Y(n_123)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_99),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_125),
.B(n_110),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_80),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_130),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_104),
.A2(n_24),
.B1(n_20),
.B2(n_40),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_L g133 ( 
.A1(n_79),
.A2(n_40),
.B(n_26),
.Y(n_133)
);

AOI21xp5_ASAP7_75t_L g139 ( 
.A1(n_133),
.A2(n_110),
.B(n_106),
.Y(n_139)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_124),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_134),
.B(n_135),
.Y(n_196)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_127),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_136),
.A2(n_142),
.B1(n_143),
.B2(n_155),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_138),
.A2(n_146),
.B1(n_150),
.B2(n_152),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_L g168 ( 
.A1(n_139),
.A2(n_144),
.B(n_131),
.Y(n_168)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_127),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_140),
.B(n_145),
.Y(n_171)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_129),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_141),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_111),
.A2(n_98),
.B1(n_81),
.B2(n_96),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_122),
.A2(n_81),
.B1(n_78),
.B2(n_91),
.Y(n_143)
);

NAND2xp33_ASAP7_75t_SL g144 ( 
.A(n_133),
.B(n_103),
.Y(n_144)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_120),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_148),
.B(n_158),
.Y(n_172)
);

INVx8_ASAP7_75t_L g149 ( 
.A(n_116),
.Y(n_149)
);

CKINVDCx14_ASAP7_75t_R g192 ( 
.A(n_149),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_121),
.A2(n_90),
.B1(n_101),
.B2(n_56),
.Y(n_150)
);

INVx4_ASAP7_75t_L g151 ( 
.A(n_116),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_151),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_105),
.A2(n_56),
.B1(n_87),
.B2(n_24),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_125),
.B(n_26),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_153),
.B(n_129),
.Y(n_182)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_129),
.Y(n_154)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_154),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_106),
.A2(n_56),
.B1(n_24),
.B2(n_20),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_120),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_159),
.A2(n_164),
.B1(n_126),
.B2(n_128),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_109),
.B(n_113),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_160),
.B(n_139),
.C(n_165),
.Y(n_178)
);

CKINVDCx14_ASAP7_75t_R g162 ( 
.A(n_131),
.Y(n_162)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_162),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_119),
.A2(n_29),
.B1(n_26),
.B2(n_3),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_105),
.A2(n_114),
.B1(n_113),
.B2(n_132),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_165),
.A2(n_146),
.B1(n_134),
.B2(n_164),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_168),
.B(n_177),
.Y(n_206)
);

AOI21xp5_ASAP7_75t_L g169 ( 
.A1(n_144),
.A2(n_117),
.B(n_108),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g218 ( 
.A1(n_169),
.A2(n_179),
.B1(n_1),
.B2(n_2),
.Y(n_218)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_161),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_173),
.B(n_174),
.Y(n_211)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_143),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_163),
.B(n_107),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_175),
.B(n_178),
.C(n_137),
.Y(n_204)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_147),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_176),
.B(n_181),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_163),
.B(n_130),
.Y(n_177)
);

AOI21xp5_ASAP7_75t_L g179 ( 
.A1(n_157),
.A2(n_118),
.B(n_123),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_L g180 ( 
.A1(n_157),
.A2(n_126),
.B(n_118),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_180),
.B(n_29),
.Y(n_212)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_142),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_182),
.B(n_186),
.Y(n_208)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_152),
.Y(n_183)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_183),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_160),
.B(n_118),
.Y(n_185)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_185),
.Y(n_209)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_155),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_156),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_187),
.B(n_188),
.Y(n_215)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_147),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_145),
.Y(n_189)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_189),
.Y(n_217)
);

INVxp67_ASAP7_75t_L g191 ( 
.A(n_150),
.Y(n_191)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_191),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_193),
.B(n_1),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_195),
.A2(n_112),
.B1(n_128),
.B2(n_149),
.Y(n_210)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_153),
.Y(n_197)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_197),
.Y(n_229)
);

OR2x2_ASAP7_75t_SL g198 ( 
.A(n_137),
.B(n_11),
.Y(n_198)
);

OAI21xp33_ASAP7_75t_L g228 ( 
.A1(n_198),
.A2(n_14),
.B(n_12),
.Y(n_228)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_159),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_199),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_158),
.A2(n_112),
.B1(n_128),
.B2(n_29),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_200),
.A2(n_154),
.B1(n_141),
.B2(n_148),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_201),
.A2(n_213),
.B1(n_226),
.B2(n_195),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_204),
.B(n_216),
.C(n_224),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_181),
.A2(n_140),
.B1(n_135),
.B2(n_149),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_207),
.B(n_219),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_210),
.A2(n_218),
.B1(n_167),
.B2(n_196),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_212),
.B(n_223),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_193),
.A2(n_116),
.B1(n_151),
.B2(n_115),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_191),
.A2(n_183),
.B1(n_174),
.B2(n_185),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_214),
.A2(n_205),
.B1(n_203),
.B2(n_208),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_178),
.B(n_115),
.C(n_26),
.Y(n_216)
);

INVxp67_ASAP7_75t_L g221 ( 
.A(n_200),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_221),
.B(n_222),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_166),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_177),
.B(n_175),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_168),
.B(n_15),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_179),
.B(n_14),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_225),
.B(n_198),
.Y(n_250)
);

OA21x2_ASAP7_75t_L g226 ( 
.A1(n_182),
.A2(n_2),
.B(n_3),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_169),
.B(n_14),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_227),
.B(n_171),
.C(n_188),
.Y(n_232)
);

CKINVDCx16_ASAP7_75t_R g246 ( 
.A(n_228),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_232),
.B(n_236),
.C(n_239),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_211),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_233),
.B(n_234),
.Y(n_276)
);

CKINVDCx14_ASAP7_75t_R g234 ( 
.A(n_201),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_217),
.B(n_172),
.Y(n_235)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_235),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_204),
.B(n_180),
.C(n_184),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_237),
.A2(n_253),
.B1(n_220),
.B2(n_226),
.Y(n_262)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_213),
.Y(n_238)
);

INVx11_ASAP7_75t_L g271 ( 
.A(n_238),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_209),
.B(n_184),
.C(n_186),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_SL g240 ( 
.A(n_206),
.B(n_190),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_240),
.B(n_252),
.Y(n_269)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_241),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_214),
.A2(n_199),
.B1(n_187),
.B2(n_190),
.Y(n_242)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_242),
.Y(n_263)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_215),
.Y(n_243)
);

AOI21xp5_ASAP7_75t_L g272 ( 
.A1(n_243),
.A2(n_248),
.B(n_251),
.Y(n_272)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_244),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_216),
.B(n_192),
.C(n_170),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_247),
.B(n_224),
.C(n_227),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_229),
.B(n_194),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_250),
.B(n_255),
.Y(n_261)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_202),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_223),
.B(n_194),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_207),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_221),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_254)
);

INVxp67_ASAP7_75t_L g259 ( 
.A(n_254),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_206),
.B(n_12),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_260),
.B(n_264),
.C(n_266),
.Y(n_279)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_262),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_230),
.B(n_219),
.C(n_212),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_230),
.B(n_225),
.C(n_226),
.Y(n_266)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_231),
.Y(n_267)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_267),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_240),
.B(n_228),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_268),
.B(n_255),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_236),
.B(n_2),
.C(n_4),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_270),
.B(n_275),
.C(n_232),
.Y(n_280)
);

FAx1_ASAP7_75t_SL g273 ( 
.A(n_245),
.B(n_5),
.CI(n_6),
.CON(n_273),
.SN(n_273)
);

NAND2xp5_ASAP7_75t_SL g283 ( 
.A(n_273),
.B(n_274),
.Y(n_283)
);

AOI211xp5_ASAP7_75t_L g274 ( 
.A1(n_245),
.A2(n_11),
.B(n_6),
.C(n_7),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_252),
.B(n_5),
.C(n_7),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_SL g296 ( 
.A(n_277),
.B(n_287),
.Y(n_296)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_280),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_257),
.B(n_247),
.C(n_239),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_281),
.B(n_285),
.C(n_289),
.Y(n_295)
);

CKINVDCx16_ASAP7_75t_R g282 ( 
.A(n_276),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_282),
.B(n_286),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_269),
.B(n_249),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_SL g286 ( 
.A(n_259),
.B(n_242),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_272),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_275),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_SL g305 ( 
.A(n_288),
.B(n_292),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_257),
.B(n_249),
.C(n_241),
.Y(n_289)
);

INVx13_ASAP7_75t_L g290 ( 
.A(n_258),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_290),
.B(n_271),
.Y(n_297)
);

AOI21xp5_ASAP7_75t_SL g291 ( 
.A1(n_263),
.A2(n_246),
.B(n_250),
.Y(n_291)
);

AOI22xp33_ASAP7_75t_SL g299 ( 
.A1(n_291),
.A2(n_273),
.B1(n_271),
.B2(n_268),
.Y(n_299)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_270),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_265),
.A2(n_5),
.B1(n_7),
.B2(n_8),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_293),
.A2(n_259),
.B1(n_266),
.B2(n_273),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_278),
.B(n_256),
.Y(n_294)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_294),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_297),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_299),
.A2(n_280),
.B1(n_284),
.B2(n_291),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_300),
.B(n_302),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_290),
.B(n_261),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_289),
.B(n_269),
.C(n_264),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_303),
.B(n_307),
.C(n_295),
.Y(n_314)
);

OAI221xp5_ASAP7_75t_L g304 ( 
.A1(n_283),
.A2(n_261),
.B1(n_260),
.B2(n_9),
.C(n_10),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g308 ( 
.A(n_304),
.B(n_293),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_284),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_306),
.A2(n_8),
.B1(n_10),
.B2(n_277),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_281),
.B(n_8),
.C(n_9),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_308),
.B(n_300),
.Y(n_320)
);

XOR2xp5_ASAP7_75t_L g309 ( 
.A(n_295),
.B(n_285),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_309),
.B(n_314),
.C(n_306),
.Y(n_322)
);

XNOR2xp5_ASAP7_75t_L g328 ( 
.A(n_311),
.B(n_319),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_301),
.B(n_294),
.Y(n_312)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_312),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_313),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_305),
.B(n_279),
.Y(n_315)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_315),
.Y(n_327)
);

AND2x2_ASAP7_75t_L g316 ( 
.A(n_307),
.B(n_279),
.Y(n_316)
);

OAI21xp5_ASAP7_75t_SL g321 ( 
.A1(n_316),
.A2(n_298),
.B(n_296),
.Y(n_321)
);

XNOR2xp5_ASAP7_75t_L g319 ( 
.A(n_303),
.B(n_10),
.Y(n_319)
);

OAI21xp5_ASAP7_75t_L g329 ( 
.A1(n_320),
.A2(n_321),
.B(n_322),
.Y(n_329)
);

OAI21xp5_ASAP7_75t_SL g325 ( 
.A1(n_314),
.A2(n_310),
.B(n_316),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_325),
.B(n_326),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_318),
.B(n_317),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_328),
.B(n_308),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_331),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_328),
.B(n_319),
.Y(n_332)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_332),
.Y(n_336)
);

OR2x2_ASAP7_75t_L g333 ( 
.A(n_324),
.B(n_309),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_333),
.B(n_334),
.Y(n_337)
);

INVxp67_ASAP7_75t_L g334 ( 
.A(n_321),
.Y(n_334)
);

OAI21xp5_ASAP7_75t_SL g338 ( 
.A1(n_336),
.A2(n_322),
.B(n_330),
.Y(n_338)
);

OAI22xp5_ASAP7_75t_L g339 ( 
.A1(n_338),
.A2(n_335),
.B1(n_333),
.B2(n_337),
.Y(n_339)
);

AOI21xp5_ASAP7_75t_L g340 ( 
.A1(n_339),
.A2(n_329),
.B(n_327),
.Y(n_340)
);

BUFx24_ASAP7_75t_SL g341 ( 
.A(n_340),
.Y(n_341)
);

XOR2xp5_ASAP7_75t_L g342 ( 
.A(n_341),
.B(n_323),
.Y(n_342)
);


endmodule