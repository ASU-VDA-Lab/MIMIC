module fake_jpeg_13304_n_85 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_26, n_9, n_5, n_11, n_17, n_25, n_2, n_12, n_8, n_15, n_7, n_85);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_85;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_44;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_35;
wire n_48;
wire n_46;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_3),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_15),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_22),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_3),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_20),
.B(n_27),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_8),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_6),
.Y(n_36)
);

INVx11_ASAP7_75t_SL g37 ( 
.A(n_12),
.Y(n_37)
);

BUFx16f_ASAP7_75t_L g38 ( 
.A(n_9),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_24),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_28),
.B(n_0),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_40),
.B(n_42),
.Y(n_49)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_30),
.Y(n_41)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_33),
.B(n_0),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_43),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g44 ( 
.A(n_36),
.B(n_1),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_44),
.B(n_45),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_35),
.B(n_2),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_29),
.B(n_2),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g47 ( 
.A(n_46),
.B(n_4),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_47),
.B(n_52),
.Y(n_64)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_43),
.Y(n_51)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_51),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_41),
.B(n_29),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_41),
.A2(n_30),
.B1(n_37),
.B2(n_38),
.Y(n_53)
);

OAI21xp5_ASAP7_75t_L g61 ( 
.A1(n_53),
.A2(n_38),
.B(n_32),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_54),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_55),
.B(n_56),
.Y(n_67)
);

BUFx8_ASAP7_75t_L g56 ( 
.A(n_48),
.Y(n_56)
);

XNOR2xp5_ASAP7_75t_L g57 ( 
.A(n_49),
.B(n_34),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_57),
.B(n_62),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_49),
.B(n_31),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_58),
.B(n_4),
.Y(n_70)
);

A2O1A1Ixp33_ASAP7_75t_L g60 ( 
.A1(n_50),
.A2(n_38),
.B(n_37),
.C(n_30),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_60),
.B(n_51),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_61),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_73)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_54),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_53),
.A2(n_39),
.B1(n_5),
.B2(n_6),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_63),
.A2(n_65),
.B1(n_47),
.B2(n_48),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_50),
.A2(n_14),
.B1(n_25),
.B2(n_23),
.Y(n_65)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_68),
.Y(n_77)
);

XOR2xp5_ASAP7_75t_L g75 ( 
.A(n_69),
.B(n_71),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_70),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_64),
.B(n_7),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_SL g72 ( 
.A(n_57),
.B(n_7),
.C(n_8),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_60),
.B(n_59),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_75),
.B(n_74),
.Y(n_78)
);

AOI21xp5_ASAP7_75t_L g80 ( 
.A1(n_78),
.A2(n_79),
.B(n_72),
.Y(n_80)
);

OAI21x1_ASAP7_75t_L g79 ( 
.A1(n_75),
.A2(n_66),
.B(n_67),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_80),
.A2(n_76),
.B1(n_77),
.B2(n_68),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_81),
.B(n_56),
.Y(n_82)
);

AOI21xp5_ASAP7_75t_L g83 ( 
.A1(n_82),
.A2(n_73),
.B(n_56),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_83),
.B(n_73),
.C(n_13),
.Y(n_84)
);

AOI322xp5_ASAP7_75t_L g85 ( 
.A1(n_84),
.A2(n_26),
.A3(n_16),
.B1(n_17),
.B2(n_18),
.C1(n_19),
.C2(n_21),
.Y(n_85)
);


endmodule