module fake_jpeg_24533_n_335 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_335);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_335;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_145;
wire n_18;
wire n_20;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx5_ASAP7_75t_L g15 ( 
.A(n_4),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_12),
.Y(n_16)
);

BUFx3_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

BUFx8_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

INVx2_ASAP7_75t_SL g22 ( 
.A(n_9),
.Y(n_22)
);

OR2x2_ASAP7_75t_L g23 ( 
.A(n_9),
.B(n_11),
.Y(n_23)
);

BUFx12_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_14),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_23),
.B(n_0),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_32),
.B(n_23),
.Y(n_45)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_26),
.Y(n_33)
);

INVx11_ASAP7_75t_L g48 ( 
.A(n_33),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_34),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_30),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_35),
.B(n_36),
.Y(n_43)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_37),
.B(n_38),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_30),
.Y(n_38)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_16),
.Y(n_39)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_39),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_23),
.B(n_0),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_40),
.B(n_41),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_30),
.Y(n_41)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_17),
.Y(n_42)
);

INVx13_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_45),
.B(n_52),
.Y(n_91)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_42),
.Y(n_47)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_47),
.Y(n_76)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_40),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_50),
.B(n_55),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_32),
.B(n_23),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_51),
.B(n_53),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_32),
.B(n_31),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_40),
.B(n_41),
.Y(n_53)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_42),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_56),
.B(n_57),
.Y(n_75)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_42),
.Y(n_57)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_34),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_59),
.B(n_61),
.Y(n_87)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_34),
.Y(n_60)
);

CKINVDCx14_ASAP7_75t_R g70 ( 
.A(n_60),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_35),
.B(n_38),
.Y(n_61)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_34),
.Y(n_62)
);

HB1xp67_ASAP7_75t_L g90 ( 
.A(n_62),
.Y(n_90)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_39),
.Y(n_63)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_63),
.Y(n_66)
);

AOI21xp5_ASAP7_75t_L g64 ( 
.A1(n_34),
.A2(n_28),
.B(n_25),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_64),
.A2(n_65),
.B1(n_22),
.B2(n_28),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_39),
.A2(n_26),
.B1(n_22),
.B2(n_28),
.Y(n_65)
);

OAI22xp33_ASAP7_75t_L g67 ( 
.A1(n_48),
.A2(n_39),
.B1(n_26),
.B2(n_25),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_67),
.A2(n_80),
.B1(n_37),
.B2(n_33),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_60),
.Y(n_68)
);

INVx6_ASAP7_75t_L g105 ( 
.A(n_68),
.Y(n_105)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_60),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_69),
.B(n_72),
.Y(n_96)
);

CKINVDCx9p33_ASAP7_75t_R g71 ( 
.A(n_48),
.Y(n_71)
);

HB1xp67_ASAP7_75t_L g110 ( 
.A(n_71),
.Y(n_110)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_48),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_61),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_74),
.B(n_81),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_45),
.A2(n_37),
.B1(n_33),
.B2(n_36),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_77),
.A2(n_78),
.B1(n_79),
.B2(n_82),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_50),
.A2(n_51),
.B1(n_52),
.B2(n_25),
.Y(n_78)
);

A2O1A1Ixp33_ASAP7_75t_SL g80 ( 
.A1(n_64),
.A2(n_17),
.B(n_15),
.C(n_27),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_46),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_L g82 ( 
.A1(n_49),
.A2(n_27),
.B1(n_17),
.B2(n_15),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_46),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_83),
.Y(n_97)
);

BUFx12f_ASAP7_75t_L g84 ( 
.A(n_57),
.Y(n_84)
);

INVx8_ASAP7_75t_L g94 ( 
.A(n_84),
.Y(n_94)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_54),
.Y(n_85)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_85),
.Y(n_95)
);

BUFx3_ASAP7_75t_L g86 ( 
.A(n_62),
.Y(n_86)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_86),
.Y(n_92)
);

INVx13_ASAP7_75t_L g88 ( 
.A(n_58),
.Y(n_88)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_88),
.Y(n_103)
);

INVx2_ASAP7_75t_SL g93 ( 
.A(n_90),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_93),
.B(n_101),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_74),
.B(n_49),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_99),
.B(n_115),
.Y(n_133)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_86),
.Y(n_100)
);

INVx6_ASAP7_75t_L g124 ( 
.A(n_100),
.Y(n_124)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_84),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_L g134 ( 
.A1(n_102),
.A2(n_107),
.B1(n_85),
.B2(n_54),
.Y(n_134)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_75),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_104),
.B(n_112),
.Y(n_139)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_84),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_106),
.B(n_111),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_81),
.A2(n_37),
.B1(n_33),
.B2(n_36),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_91),
.B(n_53),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_108),
.B(n_117),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_87),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_73),
.Y(n_112)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_77),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_113),
.B(n_114),
.Y(n_138)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_89),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g115 ( 
.A(n_89),
.B(n_43),
.Y(n_115)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_84),
.Y(n_116)
);

HB1xp67_ASAP7_75t_L g141 ( 
.A(n_116),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_91),
.B(n_43),
.Y(n_117)
);

INVx4_ASAP7_75t_L g118 ( 
.A(n_110),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_118),
.B(n_120),
.Y(n_152)
);

AND2x6_ASAP7_75t_L g119 ( 
.A(n_97),
.B(n_80),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_119),
.B(n_135),
.Y(n_151)
);

BUFx5_ASAP7_75t_L g120 ( 
.A(n_101),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_SL g122 ( 
.A1(n_117),
.A2(n_83),
.B(n_80),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_SL g165 ( 
.A1(n_122),
.A2(n_129),
.B(n_56),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_114),
.B(n_91),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_123),
.B(n_127),
.Y(n_145)
);

XOR2xp5_ASAP7_75t_L g125 ( 
.A(n_108),
.B(n_78),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_125),
.B(n_59),
.C(n_95),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_97),
.B(n_76),
.Y(n_127)
);

OR2x6_ASAP7_75t_L g129 ( 
.A(n_109),
.B(n_80),
.Y(n_129)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_96),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_130),
.B(n_132),
.Y(n_169)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_94),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_131),
.Y(n_156)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_107),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_134),
.A2(n_71),
.B1(n_95),
.B2(n_44),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g135 ( 
.A(n_98),
.B(n_80),
.Y(n_135)
);

INVx13_ASAP7_75t_L g136 ( 
.A(n_106),
.Y(n_136)
);

CKINVDCx14_ASAP7_75t_R g150 ( 
.A(n_136),
.Y(n_150)
);

INVx13_ASAP7_75t_L g137 ( 
.A(n_116),
.Y(n_137)
);

INVxp67_ASAP7_75t_L g158 ( 
.A(n_137),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_111),
.B(n_76),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_140),
.B(n_142),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_112),
.B(n_88),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_102),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_143),
.B(n_144),
.Y(n_168)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_93),
.Y(n_144)
);

XOR2xp5_ASAP7_75t_L g146 ( 
.A(n_125),
.B(n_113),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_146),
.B(n_153),
.C(n_160),
.Y(n_172)
);

INVx5_ASAP7_75t_L g147 ( 
.A(n_124),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_147),
.B(n_148),
.Y(n_195)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_126),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_143),
.A2(n_104),
.B1(n_27),
.B2(n_103),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_149),
.A2(n_155),
.B1(n_171),
.B2(n_118),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_122),
.B(n_121),
.Y(n_153)
);

AOI21xp5_ASAP7_75t_SL g154 ( 
.A1(n_129),
.A2(n_103),
.B(n_19),
.Y(n_154)
);

HAxp5_ASAP7_75t_SL g193 ( 
.A(n_154),
.B(n_165),
.CON(n_193),
.SN(n_193)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_129),
.A2(n_36),
.B1(n_63),
.B2(n_44),
.Y(n_155)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_127),
.Y(n_157)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_157),
.Y(n_173)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_120),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_159),
.B(n_161),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g161 ( 
.A(n_141),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_128),
.Y(n_162)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_162),
.Y(n_183)
);

MAJx2_ASAP7_75t_L g164 ( 
.A(n_129),
.B(n_17),
.C(n_88),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_164),
.B(n_123),
.C(n_140),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_129),
.A2(n_119),
.B1(n_132),
.B2(n_135),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_166),
.A2(n_170),
.B1(n_58),
.B2(n_144),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_139),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_167),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_138),
.A2(n_72),
.B1(n_93),
.B2(n_66),
.Y(n_171)
);

AND2x6_ASAP7_75t_L g175 ( 
.A(n_151),
.B(n_121),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_L g216 ( 
.A1(n_175),
.A2(n_181),
.B(n_184),
.Y(n_216)
);

CKINVDCx14_ASAP7_75t_R g220 ( 
.A(n_176),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_156),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_178),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_179),
.B(n_153),
.Y(n_200)
);

INVx13_ASAP7_75t_L g180 ( 
.A(n_158),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_180),
.B(n_186),
.Y(n_219)
);

OR2x4_ASAP7_75t_L g181 ( 
.A(n_164),
.B(n_154),
.Y(n_181)
);

HB1xp67_ASAP7_75t_L g182 ( 
.A(n_147),
.Y(n_182)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_182),
.Y(n_199)
);

AND2x6_ASAP7_75t_L g184 ( 
.A(n_151),
.B(n_133),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_185),
.A2(n_187),
.B1(n_196),
.B2(n_197),
.Y(n_209)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_168),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_168),
.A2(n_142),
.B1(n_130),
.B2(n_133),
.Y(n_187)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_158),
.Y(n_188)
);

INVx6_ASAP7_75t_L g207 ( 
.A(n_188),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_146),
.B(n_70),
.C(n_131),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_189),
.B(n_190),
.C(n_163),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_160),
.B(n_145),
.C(n_166),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_152),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_191),
.B(n_192),
.Y(n_204)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_163),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_149),
.A2(n_105),
.B1(n_124),
.B2(n_66),
.Y(n_194)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_194),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_165),
.A2(n_105),
.B1(n_55),
.B2(n_47),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_155),
.A2(n_55),
.B1(n_47),
.B2(n_58),
.Y(n_197)
);

INVx6_ASAP7_75t_L g198 ( 
.A(n_159),
.Y(n_198)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_198),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_200),
.B(n_94),
.Y(n_241)
);

INVxp67_ASAP7_75t_L g201 ( 
.A(n_177),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_201),
.B(n_205),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_203),
.B(n_190),
.C(n_189),
.Y(n_225)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_195),
.Y(n_205)
);

INVxp67_ASAP7_75t_L g206 ( 
.A(n_177),
.Y(n_206)
);

AOI21xp5_ASAP7_75t_L g234 ( 
.A1(n_206),
.A2(n_213),
.B(n_214),
.Y(n_234)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_187),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_208),
.B(n_211),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_172),
.B(n_145),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_210),
.B(n_174),
.Y(n_230)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_196),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_185),
.A2(n_169),
.B1(n_171),
.B2(n_161),
.Y(n_212)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_212),
.Y(n_229)
);

AOI21xp5_ASAP7_75t_L g213 ( 
.A1(n_181),
.A2(n_150),
.B(n_69),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_188),
.Y(n_214)
);

AO22x1_ASAP7_75t_L g215 ( 
.A1(n_193),
.A2(n_67),
.B1(n_16),
.B2(n_29),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_L g242 ( 
.A1(n_215),
.A2(n_100),
.B1(n_92),
.B2(n_136),
.Y(n_242)
);

CKINVDCx16_ASAP7_75t_R g217 ( 
.A(n_197),
.Y(n_217)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_217),
.Y(n_231)
);

AO21x1_ASAP7_75t_L g218 ( 
.A1(n_193),
.A2(n_18),
.B(n_19),
.Y(n_218)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_218),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_173),
.B(n_137),
.Y(n_222)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_222),
.Y(n_243)
);

INVx1_ASAP7_75t_SL g223 ( 
.A(n_180),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_L g233 ( 
.A1(n_223),
.A2(n_183),
.B(n_19),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_225),
.B(n_226),
.C(n_228),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_203),
.B(n_172),
.C(n_179),
.Y(n_226)
);

CKINVDCx14_ASAP7_75t_R g227 ( 
.A(n_219),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_227),
.B(n_244),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_216),
.B(n_175),
.C(n_184),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_230),
.B(n_237),
.Y(n_247)
);

CKINVDCx14_ASAP7_75t_R g260 ( 
.A(n_233),
.Y(n_260)
);

BUFx6f_ASAP7_75t_L g235 ( 
.A(n_223),
.Y(n_235)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_235),
.Y(n_254)
);

HB1xp67_ASAP7_75t_L g236 ( 
.A(n_215),
.Y(n_236)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_236),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_200),
.B(n_198),
.Y(n_237)
);

INVxp67_ASAP7_75t_L g238 ( 
.A(n_222),
.Y(n_238)
);

OAI21xp5_ASAP7_75t_SL g265 ( 
.A1(n_238),
.A2(n_18),
.B(n_21),
.Y(n_265)
);

BUFx24_ASAP7_75t_SL g240 ( 
.A(n_210),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_240),
.B(n_221),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_241),
.B(n_68),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_242),
.A2(n_212),
.B1(n_215),
.B2(n_207),
.Y(n_256)
);

NOR3xp33_ASAP7_75t_SL g244 ( 
.A(n_216),
.B(n_41),
.C(n_38),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_213),
.B(n_68),
.C(n_92),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_246),
.B(n_237),
.C(n_243),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_250),
.B(n_253),
.C(n_266),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_241),
.B(n_209),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_251),
.B(n_264),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_L g252 ( 
.A1(n_231),
.A2(n_220),
.B1(n_202),
.B2(n_201),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_252),
.A2(n_262),
.B1(n_22),
.B2(n_16),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_238),
.B(n_206),
.Y(n_255)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_255),
.Y(n_269)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_256),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_229),
.A2(n_209),
.B1(n_224),
.B2(n_204),
.Y(n_258)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_258),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_239),
.Y(n_259)
);

OAI21xp5_ASAP7_75t_SL g278 ( 
.A1(n_259),
.A2(n_18),
.B(n_31),
.Y(n_278)
);

BUFx3_ASAP7_75t_L g261 ( 
.A(n_235),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_261),
.B(n_0),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_245),
.A2(n_204),
.B1(n_207),
.B2(n_199),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_244),
.B(n_218),
.Y(n_263)
);

AOI21xp5_ASAP7_75t_L g281 ( 
.A1(n_263),
.A2(n_265),
.B(n_21),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_225),
.B(n_16),
.Y(n_266)
);

HAxp5_ASAP7_75t_SL g267 ( 
.A(n_257),
.B(n_234),
.CON(n_267),
.SN(n_267)
);

OAI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_267),
.A2(n_281),
.B1(n_8),
.B2(n_13),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_253),
.B(n_230),
.C(n_226),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_268),
.B(n_270),
.C(n_271),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_249),
.B(n_228),
.C(n_246),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_249),
.B(n_232),
.C(n_31),
.Y(n_271)
);

AND2x2_ASAP7_75t_L g272 ( 
.A(n_251),
.B(n_12),
.Y(n_272)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_272),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_SL g273 ( 
.A(n_247),
.B(n_11),
.C(n_14),
.Y(n_273)
);

OAI21xp5_ASAP7_75t_SL g293 ( 
.A1(n_273),
.A2(n_9),
.B(n_14),
.Y(n_293)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_278),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_247),
.B(n_21),
.C(n_1),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_279),
.B(n_270),
.C(n_271),
.Y(n_295)
);

BUFx12_ASAP7_75t_L g280 ( 
.A(n_261),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_280),
.B(n_282),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_SL g291 ( 
.A(n_283),
.B(n_1),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_274),
.B(n_264),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_284),
.B(n_287),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_276),
.A2(n_260),
.B1(n_254),
.B2(n_256),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_285),
.A2(n_289),
.B1(n_294),
.B2(n_29),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_274),
.B(n_258),
.Y(n_287)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_268),
.B(n_266),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_288),
.B(n_296),
.C(n_7),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_277),
.A2(n_248),
.B1(n_262),
.B2(n_265),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_291),
.B(n_293),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_269),
.A2(n_22),
.B1(n_35),
.B2(n_29),
.Y(n_294)
);

OAI21xp5_ASAP7_75t_SL g300 ( 
.A1(n_295),
.A2(n_279),
.B(n_272),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_275),
.B(n_1),
.C(n_2),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_298),
.A2(n_267),
.B1(n_22),
.B2(n_280),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_300),
.B(n_303),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_290),
.B(n_280),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_SL g313 ( 
.A(n_302),
.B(n_304),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_297),
.B(n_29),
.Y(n_304)
);

OAI21xp5_ASAP7_75t_L g305 ( 
.A1(n_286),
.A2(n_292),
.B(n_295),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_SL g314 ( 
.A(n_305),
.B(n_306),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_307),
.A2(n_284),
.B1(n_288),
.B2(n_20),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_296),
.B(n_24),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_308),
.B(n_24),
.Y(n_312)
);

A2O1A1Ixp33_ASAP7_75t_L g309 ( 
.A1(n_287),
.A2(n_6),
.B(n_10),
.C(n_8),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_L g319 ( 
.A1(n_309),
.A2(n_310),
.B1(n_2),
.B2(n_3),
.Y(n_319)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_292),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_311),
.B(n_306),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_312),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_301),
.B(n_8),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_SL g323 ( 
.A(n_315),
.B(n_316),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_310),
.B(n_10),
.Y(n_316)
);

AND2x2_ASAP7_75t_SL g318 ( 
.A(n_305),
.B(n_10),
.Y(n_318)
);

OAI21xp5_ASAP7_75t_L g326 ( 
.A1(n_318),
.A2(n_5),
.B(n_20),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_SL g325 ( 
.A(n_319),
.B(n_5),
.Y(n_325)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_320),
.Y(n_328)
);

AOI322xp5_ASAP7_75t_L g321 ( 
.A1(n_314),
.A2(n_299),
.A3(n_309),
.B1(n_5),
.B2(n_3),
.C1(n_4),
.C2(n_24),
.Y(n_321)
);

OR2x2_ASAP7_75t_L g327 ( 
.A(n_321),
.B(n_322),
.Y(n_327)
);

OAI21xp33_ASAP7_75t_L g322 ( 
.A1(n_317),
.A2(n_4),
.B(n_5),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_325),
.B(n_326),
.C(n_323),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_SL g330 ( 
.A(n_329),
.B(n_313),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_330),
.B(n_328),
.Y(n_331)
);

AOI322xp5_ASAP7_75t_L g332 ( 
.A1(n_331),
.A2(n_20),
.A3(n_24),
.B1(n_318),
.B2(n_324),
.C1(n_327),
.C2(n_328),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_332),
.B(n_20),
.Y(n_333)
);

AOI21xp5_ASAP7_75t_SL g334 ( 
.A1(n_333),
.A2(n_20),
.B(n_24),
.Y(n_334)
);

XOR2xp5_ASAP7_75t_L g335 ( 
.A(n_334),
.B(n_20),
.Y(n_335)
);


endmodule