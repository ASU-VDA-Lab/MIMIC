module fake_netlist_1_7943_n_692 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_6, n_4, n_40, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_692);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_6;
input n_4;
input n_40;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_692;
wire n_117;
wire n_663;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_85;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_490;
wire n_247;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_446;
wire n_423;
wire n_342;
wire n_420;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_357;
wire n_90;
wire n_653;
wire n_260;
wire n_78;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_684;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_84;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g78 ( .A(n_37), .Y(n_78) );
BUFx3_ASAP7_75t_L g79 ( .A(n_39), .Y(n_79) );
INVx1_ASAP7_75t_L g80 ( .A(n_55), .Y(n_80) );
INVx1_ASAP7_75t_L g81 ( .A(n_64), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_25), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_1), .Y(n_83) );
CKINVDCx14_ASAP7_75t_R g84 ( .A(n_52), .Y(n_84) );
INVx2_ASAP7_75t_L g85 ( .A(n_32), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_15), .Y(n_86) );
CKINVDCx5p33_ASAP7_75t_R g87 ( .A(n_56), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_3), .Y(n_88) );
INVxp67_ASAP7_75t_L g89 ( .A(n_17), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_34), .Y(n_90) );
INVx2_ASAP7_75t_SL g91 ( .A(n_44), .Y(n_91) );
INVx2_ASAP7_75t_L g92 ( .A(n_1), .Y(n_92) );
INVx2_ASAP7_75t_L g93 ( .A(n_20), .Y(n_93) );
INVxp67_ASAP7_75t_L g94 ( .A(n_46), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_75), .Y(n_95) );
INVx2_ASAP7_75t_L g96 ( .A(n_77), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_62), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_24), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_66), .Y(n_99) );
INVxp33_ASAP7_75t_SL g100 ( .A(n_19), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_28), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_16), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_67), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_22), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_12), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_53), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_72), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_59), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_16), .Y(n_109) );
INVx4_ASAP7_75t_R g110 ( .A(n_12), .Y(n_110) );
CKINVDCx20_ASAP7_75t_R g111 ( .A(n_10), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_48), .Y(n_112) );
INVxp67_ASAP7_75t_SL g113 ( .A(n_4), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_73), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_15), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_65), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_35), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_29), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_31), .Y(n_119) );
INVx2_ASAP7_75t_L g120 ( .A(n_63), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_69), .Y(n_121) );
CKINVDCx14_ASAP7_75t_R g122 ( .A(n_17), .Y(n_122) );
INVxp33_ASAP7_75t_L g123 ( .A(n_68), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_60), .Y(n_124) );
CKINVDCx5p33_ASAP7_75t_R g125 ( .A(n_0), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_8), .Y(n_126) );
INVx2_ASAP7_75t_L g127 ( .A(n_85), .Y(n_127) );
INVx2_ASAP7_75t_L g128 ( .A(n_85), .Y(n_128) );
AND2x2_ASAP7_75t_L g129 ( .A(n_122), .B(n_0), .Y(n_129) );
BUFx8_ASAP7_75t_L g130 ( .A(n_91), .Y(n_130) );
INVx1_ASAP7_75t_L g131 ( .A(n_78), .Y(n_131) );
AND2x6_ASAP7_75t_L g132 ( .A(n_79), .B(n_38), .Y(n_132) );
NAND2xp5_ASAP7_75t_L g133 ( .A(n_91), .B(n_2), .Y(n_133) );
BUFx6f_ASAP7_75t_L g134 ( .A(n_79), .Y(n_134) );
AND2x2_ASAP7_75t_L g135 ( .A(n_123), .B(n_2), .Y(n_135) );
AND2x2_ASAP7_75t_L g136 ( .A(n_84), .B(n_3), .Y(n_136) );
CKINVDCx5p33_ASAP7_75t_R g137 ( .A(n_87), .Y(n_137) );
INVxp67_ASAP7_75t_L g138 ( .A(n_102), .Y(n_138) );
INVx3_ASAP7_75t_L g139 ( .A(n_92), .Y(n_139) );
NAND2xp5_ASAP7_75t_L g140 ( .A(n_89), .B(n_4), .Y(n_140) );
CKINVDCx5p33_ASAP7_75t_R g141 ( .A(n_87), .Y(n_141) );
AND2x6_ASAP7_75t_L g142 ( .A(n_80), .B(n_41), .Y(n_142) );
INVx2_ASAP7_75t_L g143 ( .A(n_93), .Y(n_143) );
BUFx2_ASAP7_75t_L g144 ( .A(n_125), .Y(n_144) );
CKINVDCx5p33_ASAP7_75t_R g145 ( .A(n_100), .Y(n_145) );
OR2x2_ASAP7_75t_SL g146 ( .A(n_92), .B(n_5), .Y(n_146) );
NOR2xp33_ASAP7_75t_L g147 ( .A(n_97), .B(n_5), .Y(n_147) );
CKINVDCx5p33_ASAP7_75t_R g148 ( .A(n_100), .Y(n_148) );
INVx3_ASAP7_75t_L g149 ( .A(n_80), .Y(n_149) );
INVx1_ASAP7_75t_L g150 ( .A(n_81), .Y(n_150) );
INVx1_ASAP7_75t_L g151 ( .A(n_81), .Y(n_151) );
INVx1_ASAP7_75t_L g152 ( .A(n_82), .Y(n_152) );
INVx2_ASAP7_75t_L g153 ( .A(n_93), .Y(n_153) );
BUFx2_ASAP7_75t_L g154 ( .A(n_125), .Y(n_154) );
INVx1_ASAP7_75t_L g155 ( .A(n_82), .Y(n_155) );
AND2x4_ASAP7_75t_L g156 ( .A(n_83), .B(n_6), .Y(n_156) );
INVx2_ASAP7_75t_L g157 ( .A(n_96), .Y(n_157) );
BUFx6f_ASAP7_75t_L g158 ( .A(n_96), .Y(n_158) );
INVx1_ASAP7_75t_L g159 ( .A(n_90), .Y(n_159) );
INVx2_ASAP7_75t_L g160 ( .A(n_120), .Y(n_160) );
HB1xp67_ASAP7_75t_L g161 ( .A(n_83), .Y(n_161) );
NAND2xp5_ASAP7_75t_L g162 ( .A(n_105), .B(n_6), .Y(n_162) );
INVx1_ASAP7_75t_L g163 ( .A(n_90), .Y(n_163) );
XOR2xp5_ASAP7_75t_L g164 ( .A(n_111), .B(n_7), .Y(n_164) );
INVx1_ASAP7_75t_L g165 ( .A(n_95), .Y(n_165) );
NOR2xp33_ASAP7_75t_R g166 ( .A(n_98), .B(n_43), .Y(n_166) );
NOR2xp33_ASAP7_75t_L g167 ( .A(n_99), .B(n_7), .Y(n_167) );
CKINVDCx5p33_ASAP7_75t_R g168 ( .A(n_94), .Y(n_168) );
CKINVDCx5p33_ASAP7_75t_R g169 ( .A(n_101), .Y(n_169) );
INVx2_ASAP7_75t_L g170 ( .A(n_120), .Y(n_170) );
CKINVDCx5p33_ASAP7_75t_R g171 ( .A(n_103), .Y(n_171) );
NAND2xp5_ASAP7_75t_L g172 ( .A(n_109), .B(n_8), .Y(n_172) );
INVx1_ASAP7_75t_L g173 ( .A(n_158), .Y(n_173) );
INVx3_ASAP7_75t_L g174 ( .A(n_156), .Y(n_174) );
INVx3_ASAP7_75t_L g175 ( .A(n_156), .Y(n_175) );
NAND2xp5_ASAP7_75t_SL g176 ( .A(n_168), .B(n_108), .Y(n_176) );
AND2x4_ASAP7_75t_L g177 ( .A(n_156), .B(n_126), .Y(n_177) );
INVx5_ASAP7_75t_L g178 ( .A(n_132), .Y(n_178) );
INVx8_ASAP7_75t_L g179 ( .A(n_132), .Y(n_179) );
INVx1_ASAP7_75t_L g180 ( .A(n_158), .Y(n_180) );
NOR2xp33_ASAP7_75t_L g181 ( .A(n_145), .B(n_114), .Y(n_181) );
AND2x4_ASAP7_75t_L g182 ( .A(n_156), .B(n_126), .Y(n_182) );
INVx1_ASAP7_75t_L g183 ( .A(n_158), .Y(n_183) );
INVx1_ASAP7_75t_L g184 ( .A(n_158), .Y(n_184) );
INVx4_ASAP7_75t_L g185 ( .A(n_132), .Y(n_185) );
NAND2xp5_ASAP7_75t_SL g186 ( .A(n_137), .B(n_112), .Y(n_186) );
INVx2_ASAP7_75t_L g187 ( .A(n_158), .Y(n_187) );
NAND2xp5_ASAP7_75t_L g188 ( .A(n_144), .B(n_104), .Y(n_188) );
INVx2_ASAP7_75t_L g189 ( .A(n_134), .Y(n_189) );
INVx3_ASAP7_75t_L g190 ( .A(n_149), .Y(n_190) );
NAND2xp33_ASAP7_75t_L g191 ( .A(n_132), .B(n_124), .Y(n_191) );
INVx1_ASAP7_75t_L g192 ( .A(n_149), .Y(n_192) );
INVx1_ASAP7_75t_L g193 ( .A(n_149), .Y(n_193) );
INVx3_ASAP7_75t_L g194 ( .A(n_149), .Y(n_194) );
INVx2_ASAP7_75t_L g195 ( .A(n_134), .Y(n_195) );
NAND2xp5_ASAP7_75t_L g196 ( .A(n_144), .B(n_107), .Y(n_196) );
INVx1_ASAP7_75t_SL g197 ( .A(n_154), .Y(n_197) );
BUFx6f_ASAP7_75t_L g198 ( .A(n_132), .Y(n_198) );
BUFx2_ASAP7_75t_L g199 ( .A(n_154), .Y(n_199) );
OR2x6_ASAP7_75t_L g200 ( .A(n_129), .B(n_86), .Y(n_200) );
AOI22xp5_ASAP7_75t_L g201 ( .A1(n_148), .A2(n_115), .B1(n_86), .B2(n_88), .Y(n_201) );
INVx2_ASAP7_75t_L g202 ( .A(n_134), .Y(n_202) );
INVx2_ASAP7_75t_L g203 ( .A(n_134), .Y(n_203) );
INVx1_ASAP7_75t_L g204 ( .A(n_131), .Y(n_204) );
AO22x1_ASAP7_75t_L g205 ( .A1(n_142), .A2(n_124), .B1(n_121), .B2(n_119), .Y(n_205) );
INVx1_ASAP7_75t_L g206 ( .A(n_131), .Y(n_206) );
INVx1_ASAP7_75t_L g207 ( .A(n_143), .Y(n_207) );
NOR2x1p5_ASAP7_75t_L g208 ( .A(n_141), .B(n_113), .Y(n_208) );
INVx1_ASAP7_75t_L g209 ( .A(n_143), .Y(n_209) );
INVx2_ASAP7_75t_SL g210 ( .A(n_130), .Y(n_210) );
HB1xp67_ASAP7_75t_SL g211 ( .A(n_164), .Y(n_211) );
BUFx3_ASAP7_75t_L g212 ( .A(n_130), .Y(n_212) );
INVx2_ASAP7_75t_L g213 ( .A(n_134), .Y(n_213) );
INVxp67_ASAP7_75t_SL g214 ( .A(n_136), .Y(n_214) );
INVx1_ASAP7_75t_L g215 ( .A(n_143), .Y(n_215) );
INVx1_ASAP7_75t_L g216 ( .A(n_157), .Y(n_216) );
INVx5_ASAP7_75t_L g217 ( .A(n_132), .Y(n_217) );
AO22x2_ASAP7_75t_L g218 ( .A1(n_164), .A2(n_121), .B1(n_119), .B2(n_118), .Y(n_218) );
BUFx2_ASAP7_75t_L g219 ( .A(n_136), .Y(n_219) );
INVx1_ASAP7_75t_L g220 ( .A(n_157), .Y(n_220) );
NOR2xp33_ASAP7_75t_L g221 ( .A(n_169), .B(n_106), .Y(n_221) );
AND2x4_ASAP7_75t_L g222 ( .A(n_161), .B(n_88), .Y(n_222) );
HB1xp67_ASAP7_75t_L g223 ( .A(n_129), .Y(n_223) );
AND2x4_ASAP7_75t_SL g224 ( .A(n_135), .B(n_118), .Y(n_224) );
INVx1_ASAP7_75t_L g225 ( .A(n_157), .Y(n_225) );
INVx8_ASAP7_75t_L g226 ( .A(n_132), .Y(n_226) );
AOI22xp5_ASAP7_75t_L g227 ( .A1(n_135), .A2(n_117), .B1(n_116), .B2(n_95), .Y(n_227) );
INVx2_ASAP7_75t_L g228 ( .A(n_170), .Y(n_228) );
INVx2_ASAP7_75t_L g229 ( .A(n_170), .Y(n_229) );
INVx2_ASAP7_75t_L g230 ( .A(n_170), .Y(n_230) );
INVx2_ASAP7_75t_L g231 ( .A(n_127), .Y(n_231) );
INVx2_ASAP7_75t_L g232 ( .A(n_127), .Y(n_232) );
INVx1_ASAP7_75t_L g233 ( .A(n_150), .Y(n_233) );
HB1xp67_ASAP7_75t_L g234 ( .A(n_197), .Y(n_234) );
AOI22xp5_ASAP7_75t_L g235 ( .A1(n_222), .A2(n_171), .B1(n_138), .B2(n_140), .Y(n_235) );
INVx1_ASAP7_75t_L g236 ( .A(n_190), .Y(n_236) );
INVx2_ASAP7_75t_SL g237 ( .A(n_212), .Y(n_237) );
INVx1_ASAP7_75t_L g238 ( .A(n_194), .Y(n_238) );
INVx2_ASAP7_75t_L g239 ( .A(n_194), .Y(n_239) );
NOR2xp33_ASAP7_75t_R g240 ( .A(n_179), .B(n_142), .Y(n_240) );
NAND2xp5_ASAP7_75t_L g241 ( .A(n_214), .B(n_130), .Y(n_241) );
BUFx6f_ASAP7_75t_L g242 ( .A(n_212), .Y(n_242) );
INVx1_ASAP7_75t_L g243 ( .A(n_194), .Y(n_243) );
NAND2xp5_ASAP7_75t_L g244 ( .A(n_222), .B(n_130), .Y(n_244) );
INVx5_ASAP7_75t_L g245 ( .A(n_179), .Y(n_245) );
INVx2_ASAP7_75t_L g246 ( .A(n_192), .Y(n_246) );
NOR3xp33_ASAP7_75t_SL g247 ( .A(n_186), .B(n_172), .C(n_162), .Y(n_247) );
NOR3xp33_ASAP7_75t_SL g248 ( .A(n_176), .B(n_167), .C(n_147), .Y(n_248) );
INVx1_ASAP7_75t_L g249 ( .A(n_207), .Y(n_249) );
OAI22xp5_ASAP7_75t_L g250 ( .A1(n_200), .A2(n_146), .B1(n_165), .B2(n_163), .Y(n_250) );
INVx6_ASAP7_75t_L g251 ( .A(n_177), .Y(n_251) );
INVx1_ASAP7_75t_L g252 ( .A(n_207), .Y(n_252) );
AND2x2_ASAP7_75t_L g253 ( .A(n_219), .B(n_151), .Y(n_253) );
INVx2_ASAP7_75t_L g254 ( .A(n_193), .Y(n_254) );
INVx2_ASAP7_75t_SL g255 ( .A(n_179), .Y(n_255) );
NAND2xp5_ASAP7_75t_L g256 ( .A(n_222), .B(n_151), .Y(n_256) );
NOR2xp33_ASAP7_75t_R g257 ( .A(n_179), .B(n_142), .Y(n_257) );
INVx4_ASAP7_75t_L g258 ( .A(n_210), .Y(n_258) );
NOR2xp33_ASAP7_75t_R g259 ( .A(n_226), .B(n_142), .Y(n_259) );
INVx1_ASAP7_75t_L g260 ( .A(n_209), .Y(n_260) );
AOI22x1_ASAP7_75t_L g261 ( .A1(n_185), .A2(n_150), .B1(n_165), .B2(n_163), .Y(n_261) );
NOR3xp33_ASAP7_75t_SL g262 ( .A(n_181), .B(n_133), .C(n_159), .Y(n_262) );
NOR2xp33_ASAP7_75t_L g263 ( .A(n_188), .B(n_152), .Y(n_263) );
BUFx2_ASAP7_75t_L g264 ( .A(n_199), .Y(n_264) );
INVx2_ASAP7_75t_L g265 ( .A(n_228), .Y(n_265) );
BUFx3_ASAP7_75t_L g266 ( .A(n_210), .Y(n_266) );
INVxp67_ASAP7_75t_L g267 ( .A(n_199), .Y(n_267) );
INVx1_ASAP7_75t_L g268 ( .A(n_209), .Y(n_268) );
NOR3xp33_ASAP7_75t_SL g269 ( .A(n_221), .B(n_196), .C(n_152), .Y(n_269) );
AOI211xp5_ASAP7_75t_L g270 ( .A1(n_223), .A2(n_159), .B(n_155), .C(n_117), .Y(n_270) );
AND2x2_ASAP7_75t_L g271 ( .A(n_219), .B(n_155), .Y(n_271) );
INVx4_ASAP7_75t_L g272 ( .A(n_226), .Y(n_272) );
INVx1_ASAP7_75t_L g273 ( .A(n_215), .Y(n_273) );
NOR2xp33_ASAP7_75t_L g274 ( .A(n_227), .B(n_139), .Y(n_274) );
INVx1_ASAP7_75t_L g275 ( .A(n_215), .Y(n_275) );
NAND2xp5_ASAP7_75t_L g276 ( .A(n_204), .B(n_206), .Y(n_276) );
INVx2_ASAP7_75t_L g277 ( .A(n_228), .Y(n_277) );
AND2x2_ASAP7_75t_L g278 ( .A(n_200), .B(n_139), .Y(n_278) );
INVx1_ASAP7_75t_SL g279 ( .A(n_224), .Y(n_279) );
AND2x2_ASAP7_75t_L g280 ( .A(n_200), .B(n_139), .Y(n_280) );
NOR2xp33_ASAP7_75t_R g281 ( .A(n_226), .B(n_142), .Y(n_281) );
NAND3xp33_ASAP7_75t_SL g282 ( .A(n_201), .B(n_166), .C(n_116), .Y(n_282) );
HB1xp67_ASAP7_75t_L g283 ( .A(n_200), .Y(n_283) );
OAI22xp5_ASAP7_75t_SL g284 ( .A1(n_211), .A2(n_146), .B1(n_139), .B2(n_110), .Y(n_284) );
HB1xp67_ASAP7_75t_L g285 ( .A(n_224), .Y(n_285) );
INVx1_ASAP7_75t_L g286 ( .A(n_216), .Y(n_286) );
INVx2_ASAP7_75t_L g287 ( .A(n_229), .Y(n_287) );
NOR2xp33_ASAP7_75t_L g288 ( .A(n_177), .B(n_160), .Y(n_288) );
CKINVDCx5p33_ASAP7_75t_R g289 ( .A(n_208), .Y(n_289) );
BUFx6f_ASAP7_75t_L g290 ( .A(n_198), .Y(n_290) );
INVx1_ASAP7_75t_SL g291 ( .A(n_216), .Y(n_291) );
NAND2xp5_ASAP7_75t_L g292 ( .A(n_233), .B(n_160), .Y(n_292) );
BUFx2_ASAP7_75t_L g293 ( .A(n_218), .Y(n_293) );
NAND2xp5_ASAP7_75t_L g294 ( .A(n_177), .B(n_153), .Y(n_294) );
INVx1_ASAP7_75t_L g295 ( .A(n_220), .Y(n_295) );
NAND2xp5_ASAP7_75t_SL g296 ( .A(n_185), .B(n_153), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g297 ( .A(n_182), .B(n_128), .Y(n_297) );
INVx1_ASAP7_75t_L g298 ( .A(n_220), .Y(n_298) );
INVx2_ASAP7_75t_L g299 ( .A(n_229), .Y(n_299) );
INVx1_ASAP7_75t_L g300 ( .A(n_249), .Y(n_300) );
BUFx3_ASAP7_75t_L g301 ( .A(n_242), .Y(n_301) );
AND2x2_ASAP7_75t_L g302 ( .A(n_234), .B(n_218), .Y(n_302) );
AOI21xp33_ASAP7_75t_L g303 ( .A1(n_244), .A2(n_191), .B(n_226), .Y(n_303) );
AND2x4_ASAP7_75t_L g304 ( .A(n_280), .B(n_278), .Y(n_304) );
INVx1_ASAP7_75t_L g305 ( .A(n_252), .Y(n_305) );
INVx2_ASAP7_75t_L g306 ( .A(n_265), .Y(n_306) );
NAND2xp5_ASAP7_75t_SL g307 ( .A(n_237), .B(n_185), .Y(n_307) );
BUFx12f_ASAP7_75t_L g308 ( .A(n_264), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g309 ( .A(n_263), .B(n_182), .Y(n_309) );
BUFx12f_ASAP7_75t_L g310 ( .A(n_289), .Y(n_310) );
AOI22xp33_ASAP7_75t_L g311 ( .A1(n_280), .A2(n_175), .B1(n_174), .B2(n_218), .Y(n_311) );
CKINVDCx6p67_ASAP7_75t_R g312 ( .A(n_279), .Y(n_312) );
NAND2x1_ASAP7_75t_L g313 ( .A(n_251), .B(n_175), .Y(n_313) );
BUFx2_ASAP7_75t_L g314 ( .A(n_283), .Y(n_314) );
AND2x2_ASAP7_75t_L g315 ( .A(n_253), .B(n_218), .Y(n_315) );
BUFx12f_ASAP7_75t_L g316 ( .A(n_289), .Y(n_316) );
INVx3_ASAP7_75t_SL g317 ( .A(n_245), .Y(n_317) );
BUFx3_ASAP7_75t_L g318 ( .A(n_242), .Y(n_318) );
INVx2_ASAP7_75t_L g319 ( .A(n_265), .Y(n_319) );
INVx2_ASAP7_75t_L g320 ( .A(n_277), .Y(n_320) );
INVx2_ASAP7_75t_L g321 ( .A(n_277), .Y(n_321) );
INVx1_ASAP7_75t_L g322 ( .A(n_260), .Y(n_322) );
AND2x2_ASAP7_75t_L g323 ( .A(n_253), .B(n_174), .Y(n_323) );
INVx1_ASAP7_75t_L g324 ( .A(n_268), .Y(n_324) );
INVx4_ASAP7_75t_SL g325 ( .A(n_251), .Y(n_325) );
AND2x4_ASAP7_75t_L g326 ( .A(n_245), .B(n_174), .Y(n_326) );
INVx2_ASAP7_75t_L g327 ( .A(n_287), .Y(n_327) );
BUFx3_ASAP7_75t_L g328 ( .A(n_242), .Y(n_328) );
AND2x6_ASAP7_75t_L g329 ( .A(n_266), .B(n_198), .Y(n_329) );
INVx1_ASAP7_75t_L g330 ( .A(n_273), .Y(n_330) );
BUFx2_ASAP7_75t_SL g331 ( .A(n_245), .Y(n_331) );
INVx6_ASAP7_75t_L g332 ( .A(n_251), .Y(n_332) );
HB1xp67_ASAP7_75t_L g333 ( .A(n_267), .Y(n_333) );
INVx2_ASAP7_75t_L g334 ( .A(n_287), .Y(n_334) );
NAND2xp5_ASAP7_75t_L g335 ( .A(n_256), .B(n_175), .Y(n_335) );
BUFx6f_ASAP7_75t_L g336 ( .A(n_290), .Y(n_336) );
NOR2xp33_ASAP7_75t_L g337 ( .A(n_235), .B(n_198), .Y(n_337) );
AND3x1_ASAP7_75t_SL g338 ( .A(n_284), .B(n_293), .C(n_247), .Y(n_338) );
AND2x4_ASAP7_75t_L g339 ( .A(n_245), .B(n_217), .Y(n_339) );
CKINVDCx14_ASAP7_75t_R g340 ( .A(n_285), .Y(n_340) );
AOI22xp5_ASAP7_75t_L g341 ( .A1(n_250), .A2(n_191), .B1(n_205), .B2(n_225), .Y(n_341) );
INVx2_ASAP7_75t_L g342 ( .A(n_299), .Y(n_342) );
INVx1_ASAP7_75t_SL g343 ( .A(n_271), .Y(n_343) );
BUFx2_ASAP7_75t_L g344 ( .A(n_291), .Y(n_344) );
INVx4_ASAP7_75t_L g345 ( .A(n_245), .Y(n_345) );
AND2x4_ASAP7_75t_L g346 ( .A(n_272), .B(n_217), .Y(n_346) );
AOI22xp33_ASAP7_75t_L g347 ( .A1(n_274), .A2(n_198), .B1(n_225), .B2(n_232), .Y(n_347) );
O2A1O1Ixp33_ASAP7_75t_L g348 ( .A1(n_274), .A2(n_230), .B(n_232), .C(n_231), .Y(n_348) );
NOR2xp33_ASAP7_75t_R g349 ( .A(n_282), .B(n_198), .Y(n_349) );
INVx1_ASAP7_75t_L g350 ( .A(n_275), .Y(n_350) );
BUFx3_ASAP7_75t_L g351 ( .A(n_242), .Y(n_351) );
AND2x2_ASAP7_75t_L g352 ( .A(n_269), .B(n_230), .Y(n_352) );
NAND2xp5_ASAP7_75t_L g353 ( .A(n_270), .B(n_205), .Y(n_353) );
INVx2_ASAP7_75t_SL g354 ( .A(n_237), .Y(n_354) );
CKINVDCx5p33_ASAP7_75t_R g355 ( .A(n_262), .Y(n_355) );
OAI22xp33_ASAP7_75t_L g356 ( .A1(n_344), .A2(n_241), .B1(n_276), .B2(n_297), .Y(n_356) );
BUFx6f_ASAP7_75t_L g357 ( .A(n_336), .Y(n_357) );
NAND3xp33_ASAP7_75t_SL g358 ( .A(n_355), .B(n_248), .C(n_294), .Y(n_358) );
NAND2xp5_ASAP7_75t_L g359 ( .A(n_344), .B(n_288), .Y(n_359) );
OAI221xp5_ASAP7_75t_L g360 ( .A1(n_311), .A2(n_288), .B1(n_261), .B2(n_238), .C(n_236), .Y(n_360) );
OR2x2_ASAP7_75t_L g361 ( .A(n_343), .B(n_286), .Y(n_361) );
NAND2xp5_ASAP7_75t_L g362 ( .A(n_323), .B(n_295), .Y(n_362) );
INVx5_ASAP7_75t_L g363 ( .A(n_329), .Y(n_363) );
AND2x6_ASAP7_75t_SL g364 ( .A(n_302), .B(n_315), .Y(n_364) );
OAI21x1_ASAP7_75t_L g365 ( .A1(n_348), .A2(n_296), .B(n_292), .Y(n_365) );
OAI22xp5_ASAP7_75t_L g366 ( .A1(n_309), .A2(n_298), .B1(n_258), .B2(n_299), .Y(n_366) );
INVx1_ASAP7_75t_SL g367 ( .A(n_308), .Y(n_367) );
A2O1A1Ixp33_ASAP7_75t_L g368 ( .A1(n_300), .A2(n_246), .B(n_254), .C(n_231), .Y(n_368) );
AND2x2_ASAP7_75t_L g369 ( .A(n_315), .B(n_239), .Y(n_369) );
AND2x2_ASAP7_75t_L g370 ( .A(n_323), .B(n_246), .Y(n_370) );
INVx1_ASAP7_75t_L g371 ( .A(n_300), .Y(n_371) );
AOI21xp5_ASAP7_75t_L g372 ( .A1(n_303), .A2(n_296), .B(n_178), .Y(n_372) );
OAI22xp5_ASAP7_75t_L g373 ( .A1(n_341), .A2(n_258), .B1(n_254), .B2(n_272), .Y(n_373) );
AND2x2_ASAP7_75t_L g374 ( .A(n_305), .B(n_243), .Y(n_374) );
OAI22xp5_ASAP7_75t_L g375 ( .A1(n_341), .A2(n_258), .B1(n_272), .B2(n_255), .Y(n_375) );
OAI211xp5_ASAP7_75t_SL g376 ( .A1(n_333), .A2(n_128), .B(n_173), .C(n_180), .Y(n_376) );
AND2x2_ASAP7_75t_L g377 ( .A(n_305), .B(n_281), .Y(n_377) );
CKINVDCx6p67_ASAP7_75t_R g378 ( .A(n_308), .Y(n_378) );
OAI21x1_ASAP7_75t_L g379 ( .A1(n_322), .A2(n_202), .B(n_189), .Y(n_379) );
INVx6_ASAP7_75t_L g380 ( .A(n_325), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_322), .Y(n_381) );
INVx2_ASAP7_75t_L g382 ( .A(n_306), .Y(n_382) );
INVx2_ASAP7_75t_L g383 ( .A(n_306), .Y(n_383) );
AOI22xp5_ASAP7_75t_L g384 ( .A1(n_355), .A2(n_255), .B1(n_178), .B2(n_217), .Y(n_384) );
NAND2xp5_ASAP7_75t_L g385 ( .A(n_314), .B(n_281), .Y(n_385) );
AND2x2_ASAP7_75t_L g386 ( .A(n_324), .B(n_259), .Y(n_386) );
OAI221xp5_ASAP7_75t_L g387 ( .A1(n_353), .A2(n_178), .B1(n_217), .B2(n_189), .C(n_202), .Y(n_387) );
OAI221xp5_ASAP7_75t_L g388 ( .A1(n_314), .A2(n_178), .B1(n_217), .B2(n_203), .C(n_213), .Y(n_388) );
CKINVDCx11_ASAP7_75t_R g389 ( .A(n_312), .Y(n_389) );
AOI22xp33_ASAP7_75t_L g390 ( .A1(n_358), .A2(n_352), .B1(n_304), .B2(n_337), .Y(n_390) );
AND2x4_ASAP7_75t_L g391 ( .A(n_371), .B(n_304), .Y(n_391) );
OAI221xp5_ASAP7_75t_L g392 ( .A1(n_359), .A2(n_352), .B1(n_335), .B2(n_347), .C(n_313), .Y(n_392) );
INVxp67_ASAP7_75t_L g393 ( .A(n_361), .Y(n_393) );
NAND2xp5_ASAP7_75t_L g394 ( .A(n_361), .B(n_304), .Y(n_394) );
INVx1_ASAP7_75t_L g395 ( .A(n_381), .Y(n_395) );
AOI22xp33_ASAP7_75t_SL g396 ( .A1(n_377), .A2(n_340), .B1(n_331), .B2(n_304), .Y(n_396) );
BUFx3_ASAP7_75t_L g397 ( .A(n_380), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_374), .Y(n_398) );
O2A1O1Ixp33_ASAP7_75t_SL g399 ( .A1(n_356), .A2(n_350), .B(n_324), .C(n_330), .Y(n_399) );
NOR2xp33_ASAP7_75t_L g400 ( .A(n_367), .B(n_312), .Y(n_400) );
OR2x2_ASAP7_75t_L g401 ( .A(n_369), .B(n_330), .Y(n_401) );
AND2x2_ASAP7_75t_SL g402 ( .A(n_377), .B(n_345), .Y(n_402) );
AND2x2_ASAP7_75t_L g403 ( .A(n_370), .B(n_350), .Y(n_403) );
NOR2xp33_ASAP7_75t_L g404 ( .A(n_364), .B(n_310), .Y(n_404) );
INVx2_ASAP7_75t_L g405 ( .A(n_382), .Y(n_405) );
OR2x2_ASAP7_75t_L g406 ( .A(n_369), .B(n_319), .Y(n_406) );
HB1xp67_ASAP7_75t_L g407 ( .A(n_378), .Y(n_407) );
AOI22xp33_ASAP7_75t_L g408 ( .A1(n_370), .A2(n_313), .B1(n_332), .B2(n_326), .Y(n_408) );
AO21x2_ASAP7_75t_L g409 ( .A1(n_368), .A2(n_349), .B(n_240), .Y(n_409) );
AOI222xp33_ASAP7_75t_L g410 ( .A1(n_389), .A2(n_310), .B1(n_316), .B2(n_325), .C1(n_338), .C2(n_332), .Y(n_410) );
INVx3_ASAP7_75t_L g411 ( .A(n_363), .Y(n_411) );
OAI22xp5_ASAP7_75t_L g412 ( .A1(n_362), .A2(n_354), .B1(n_321), .B2(n_320), .Y(n_412) );
INVx1_ASAP7_75t_L g413 ( .A(n_374), .Y(n_413) );
OAI22xp5_ASAP7_75t_L g414 ( .A1(n_386), .A2(n_354), .B1(n_321), .B2(n_320), .Y(n_414) );
INVx1_ASAP7_75t_L g415 ( .A(n_382), .Y(n_415) );
BUFx6f_ASAP7_75t_L g416 ( .A(n_357), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_383), .Y(n_417) );
INVx3_ASAP7_75t_L g418 ( .A(n_411), .Y(n_418) );
OR2x2_ASAP7_75t_L g419 ( .A(n_393), .B(n_383), .Y(n_419) );
AOI221xp5_ASAP7_75t_L g420 ( .A1(n_398), .A2(n_360), .B1(n_376), .B2(n_368), .C(n_385), .Y(n_420) );
NOR3xp33_ASAP7_75t_L g421 ( .A(n_392), .B(n_389), .C(n_388), .Y(n_421) );
AND2x4_ASAP7_75t_L g422 ( .A(n_398), .B(n_363), .Y(n_422) );
AOI22xp33_ASAP7_75t_L g423 ( .A1(n_390), .A2(n_386), .B1(n_378), .B2(n_366), .Y(n_423) );
AOI33xp33_ASAP7_75t_L g424 ( .A1(n_395), .A2(n_184), .A3(n_180), .B1(n_183), .B2(n_173), .B3(n_195), .Y(n_424) );
AND2x2_ASAP7_75t_L g425 ( .A(n_403), .B(n_319), .Y(n_425) );
INVx2_ASAP7_75t_L g426 ( .A(n_405), .Y(n_426) );
AOI221xp5_ASAP7_75t_L g427 ( .A1(n_413), .A2(n_373), .B1(n_334), .B2(n_342), .C(n_327), .Y(n_427) );
BUFx3_ASAP7_75t_L g428 ( .A(n_397), .Y(n_428) );
BUFx3_ASAP7_75t_L g429 ( .A(n_397), .Y(n_429) );
AND2x2_ASAP7_75t_L g430 ( .A(n_403), .B(n_327), .Y(n_430) );
AND2x4_ASAP7_75t_L g431 ( .A(n_413), .B(n_363), .Y(n_431) );
OAI31xp33_ASAP7_75t_L g432 ( .A1(n_399), .A2(n_375), .A3(n_326), .B(n_342), .Y(n_432) );
NOR2xp33_ASAP7_75t_L g433 ( .A(n_407), .B(n_316), .Y(n_433) );
INVx2_ASAP7_75t_L g434 ( .A(n_405), .Y(n_434) );
INVx1_ASAP7_75t_L g435 ( .A(n_415), .Y(n_435) );
AND2x2_ASAP7_75t_L g436 ( .A(n_415), .B(n_365), .Y(n_436) );
NOR2xp33_ASAP7_75t_L g437 ( .A(n_404), .B(n_332), .Y(n_437) );
AND2x2_ASAP7_75t_L g438 ( .A(n_417), .B(n_365), .Y(n_438) );
AO21x2_ASAP7_75t_L g439 ( .A1(n_409), .A2(n_379), .B(n_372), .Y(n_439) );
BUFx3_ASAP7_75t_L g440 ( .A(n_402), .Y(n_440) );
INVx2_ASAP7_75t_L g441 ( .A(n_417), .Y(n_441) );
CKINVDCx5p33_ASAP7_75t_R g442 ( .A(n_400), .Y(n_442) );
OAI211xp5_ASAP7_75t_L g443 ( .A1(n_410), .A2(n_363), .B(n_345), .C(n_257), .Y(n_443) );
NAND4xp25_ASAP7_75t_L g444 ( .A(n_396), .B(n_183), .C(n_184), .D(n_195), .Y(n_444) );
INVx1_ASAP7_75t_L g445 ( .A(n_395), .Y(n_445) );
OAI21xp5_ASAP7_75t_L g446 ( .A1(n_412), .A2(n_387), .B(n_379), .Y(n_446) );
OAI211xp5_ASAP7_75t_L g447 ( .A1(n_408), .A2(n_363), .B(n_345), .C(n_240), .Y(n_447) );
BUFx3_ASAP7_75t_L g448 ( .A(n_402), .Y(n_448) );
OAI21xp33_ASAP7_75t_L g449 ( .A1(n_394), .A2(n_203), .B(n_213), .Y(n_449) );
AO21x1_ASAP7_75t_L g450 ( .A1(n_414), .A2(n_307), .B(n_187), .Y(n_450) );
AND2x4_ASAP7_75t_L g451 ( .A(n_411), .B(n_357), .Y(n_451) );
OR2x6_ASAP7_75t_L g452 ( .A(n_411), .B(n_380), .Y(n_452) );
AND2x2_ASAP7_75t_L g453 ( .A(n_441), .B(n_406), .Y(n_453) );
AND2x2_ASAP7_75t_L g454 ( .A(n_441), .B(n_406), .Y(n_454) );
INVx3_ASAP7_75t_L g455 ( .A(n_451), .Y(n_455) );
AND2x4_ASAP7_75t_L g456 ( .A(n_436), .B(n_416), .Y(n_456) );
HB1xp67_ASAP7_75t_L g457 ( .A(n_441), .Y(n_457) );
INVx2_ASAP7_75t_L g458 ( .A(n_426), .Y(n_458) );
INVx1_ASAP7_75t_L g459 ( .A(n_445), .Y(n_459) );
AND2x2_ASAP7_75t_L g460 ( .A(n_445), .B(n_435), .Y(n_460) );
NAND2xp5_ASAP7_75t_L g461 ( .A(n_425), .B(n_401), .Y(n_461) );
BUFx6f_ASAP7_75t_L g462 ( .A(n_451), .Y(n_462) );
OR2x2_ASAP7_75t_L g463 ( .A(n_435), .B(n_401), .Y(n_463) );
INVx2_ASAP7_75t_L g464 ( .A(n_426), .Y(n_464) );
INVx1_ASAP7_75t_L g465 ( .A(n_436), .Y(n_465) );
OA211x2_ASAP7_75t_L g466 ( .A1(n_432), .A2(n_409), .B(n_380), .C(n_11), .Y(n_466) );
INVx2_ASAP7_75t_L g467 ( .A(n_426), .Y(n_467) );
INVx1_ASAP7_75t_L g468 ( .A(n_438), .Y(n_468) );
INVx2_ASAP7_75t_L g469 ( .A(n_434), .Y(n_469) );
NAND2xp5_ASAP7_75t_SL g470 ( .A(n_440), .B(n_416), .Y(n_470) );
AOI21xp5_ASAP7_75t_L g471 ( .A1(n_446), .A2(n_357), .B(n_416), .Y(n_471) );
NOR3xp33_ASAP7_75t_L g472 ( .A(n_421), .B(n_391), .C(n_187), .Y(n_472) );
INVx1_ASAP7_75t_L g473 ( .A(n_438), .Y(n_473) );
OAI31xp33_ASAP7_75t_SL g474 ( .A1(n_443), .A2(n_391), .A3(n_10), .B(n_11), .Y(n_474) );
AOI221xp5_ASAP7_75t_L g475 ( .A1(n_437), .A2(n_328), .B1(n_301), .B2(n_351), .C(n_318), .Y(n_475) );
OAI21x1_ASAP7_75t_L g476 ( .A1(n_450), .A2(n_416), .B(n_384), .Y(n_476) );
OAI22xp5_ASAP7_75t_L g477 ( .A1(n_440), .A2(n_416), .B1(n_328), .B2(n_351), .Y(n_477) );
CKINVDCx5p33_ASAP7_75t_R g478 ( .A(n_442), .Y(n_478) );
INVx2_ASAP7_75t_L g479 ( .A(n_434), .Y(n_479) );
AOI22xp33_ASAP7_75t_L g480 ( .A1(n_440), .A2(n_318), .B1(n_301), .B2(n_329), .Y(n_480) );
HB1xp67_ASAP7_75t_L g481 ( .A(n_419), .Y(n_481) );
AND2x2_ASAP7_75t_L g482 ( .A(n_425), .B(n_9), .Y(n_482) );
INVx1_ASAP7_75t_SL g483 ( .A(n_419), .Y(n_483) );
INVx2_ASAP7_75t_L g484 ( .A(n_434), .Y(n_484) );
OR2x2_ASAP7_75t_L g485 ( .A(n_448), .B(n_9), .Y(n_485) );
INVx1_ASAP7_75t_L g486 ( .A(n_418), .Y(n_486) );
INVx2_ASAP7_75t_L g487 ( .A(n_439), .Y(n_487) );
INVxp67_ASAP7_75t_SL g488 ( .A(n_448), .Y(n_488) );
AND2x2_ASAP7_75t_L g489 ( .A(n_430), .B(n_13), .Y(n_489) );
AOI31xp33_ASAP7_75t_L g490 ( .A1(n_433), .A2(n_13), .A3(n_14), .B(n_18), .Y(n_490) );
NOR2x1_ASAP7_75t_L g491 ( .A(n_418), .B(n_357), .Y(n_491) );
OR2x2_ASAP7_75t_L g492 ( .A(n_430), .B(n_14), .Y(n_492) );
INVx1_ASAP7_75t_L g493 ( .A(n_418), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_423), .B(n_18), .Y(n_494) );
OAI31xp33_ASAP7_75t_L g495 ( .A1(n_443), .A2(n_339), .A3(n_346), .B(n_325), .Y(n_495) );
INVx2_ASAP7_75t_L g496 ( .A(n_439), .Y(n_496) );
BUFx2_ASAP7_75t_L g497 ( .A(n_451), .Y(n_497) );
OR2x2_ASAP7_75t_L g498 ( .A(n_418), .B(n_317), .Y(n_498) );
AND2x2_ASAP7_75t_L g499 ( .A(n_422), .B(n_21), .Y(n_499) );
OR2x2_ASAP7_75t_L g500 ( .A(n_483), .B(n_439), .Y(n_500) );
OR2x4_ASAP7_75t_L g501 ( .A(n_490), .B(n_432), .Y(n_501) );
INVx1_ASAP7_75t_L g502 ( .A(n_460), .Y(n_502) );
INVx1_ASAP7_75t_L g503 ( .A(n_459), .Y(n_503) );
INVx1_ASAP7_75t_L g504 ( .A(n_459), .Y(n_504) );
AO21x2_ASAP7_75t_L g505 ( .A1(n_476), .A2(n_450), .B(n_439), .Y(n_505) );
INVx1_ASAP7_75t_L g506 ( .A(n_481), .Y(n_506) );
INVx2_ASAP7_75t_SL g507 ( .A(n_457), .Y(n_507) );
INVx2_ASAP7_75t_SL g508 ( .A(n_462), .Y(n_508) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_483), .B(n_422), .Y(n_509) );
AND2x2_ASAP7_75t_L g510 ( .A(n_465), .B(n_422), .Y(n_510) );
AND2x2_ASAP7_75t_L g511 ( .A(n_465), .B(n_431), .Y(n_511) );
NAND3x1_ASAP7_75t_SL g512 ( .A(n_495), .B(n_427), .C(n_420), .Y(n_512) );
AND5x1_ASAP7_75t_L g513 ( .A(n_474), .B(n_420), .C(n_427), .D(n_444), .E(n_452), .Y(n_513) );
INVx1_ASAP7_75t_L g514 ( .A(n_463), .Y(n_514) );
INVx2_ASAP7_75t_L g515 ( .A(n_458), .Y(n_515) );
INVx1_ASAP7_75t_L g516 ( .A(n_463), .Y(n_516) );
AND2x2_ASAP7_75t_L g517 ( .A(n_468), .B(n_431), .Y(n_517) );
INVx2_ASAP7_75t_L g518 ( .A(n_458), .Y(n_518) );
NOR2xp33_ASAP7_75t_R g519 ( .A(n_478), .B(n_429), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_453), .B(n_431), .Y(n_520) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_453), .B(n_429), .Y(n_521) );
INVx1_ASAP7_75t_L g522 ( .A(n_454), .Y(n_522) );
BUFx2_ASAP7_75t_L g523 ( .A(n_488), .Y(n_523) );
NAND2xp5_ASAP7_75t_SL g524 ( .A(n_495), .B(n_451), .Y(n_524) );
AND2x2_ASAP7_75t_L g525 ( .A(n_468), .B(n_429), .Y(n_525) );
INVx2_ASAP7_75t_L g526 ( .A(n_458), .Y(n_526) );
OR2x2_ASAP7_75t_L g527 ( .A(n_473), .B(n_428), .Y(n_527) );
AND2x2_ASAP7_75t_SL g528 ( .A(n_485), .B(n_424), .Y(n_528) );
AND2x2_ASAP7_75t_L g529 ( .A(n_473), .B(n_428), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_454), .B(n_428), .Y(n_530) );
INVx1_ASAP7_75t_L g531 ( .A(n_485), .Y(n_531) );
INVx1_ASAP7_75t_L g532 ( .A(n_492), .Y(n_532) );
AND2x2_ASAP7_75t_L g533 ( .A(n_456), .B(n_452), .Y(n_533) );
INVx1_ASAP7_75t_L g534 ( .A(n_492), .Y(n_534) );
INVx1_ASAP7_75t_SL g535 ( .A(n_482), .Y(n_535) );
INVx1_ASAP7_75t_L g536 ( .A(n_464), .Y(n_536) );
INVx1_ASAP7_75t_L g537 ( .A(n_464), .Y(n_537) );
INVx1_ASAP7_75t_L g538 ( .A(n_464), .Y(n_538) );
AND2x2_ASAP7_75t_L g539 ( .A(n_456), .B(n_467), .Y(n_539) );
AND2x2_ASAP7_75t_L g540 ( .A(n_456), .B(n_452), .Y(n_540) );
AOI22xp33_ASAP7_75t_L g541 ( .A1(n_472), .A2(n_452), .B1(n_449), .B2(n_329), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_482), .B(n_452), .Y(n_542) );
NAND2xp33_ASAP7_75t_R g543 ( .A(n_499), .B(n_259), .Y(n_543) );
INVx2_ASAP7_75t_L g544 ( .A(n_467), .Y(n_544) );
INVx2_ASAP7_75t_L g545 ( .A(n_467), .Y(n_545) );
INVx2_ASAP7_75t_SL g546 ( .A(n_462), .Y(n_546) );
AND2x4_ASAP7_75t_L g547 ( .A(n_455), .B(n_23), .Y(n_547) );
OR2x2_ASAP7_75t_L g548 ( .A(n_461), .B(n_449), .Y(n_548) );
INVx2_ASAP7_75t_SL g549 ( .A(n_462), .Y(n_549) );
AND2x2_ASAP7_75t_L g550 ( .A(n_456), .B(n_26), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g551 ( .A(n_489), .B(n_447), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g552 ( .A(n_489), .B(n_447), .Y(n_552) );
INVx3_ASAP7_75t_L g553 ( .A(n_462), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g554 ( .A(n_469), .B(n_325), .Y(n_554) );
OR2x2_ASAP7_75t_L g555 ( .A(n_469), .B(n_27), .Y(n_555) );
AOI22xp5_ASAP7_75t_L g556 ( .A1(n_501), .A2(n_494), .B1(n_466), .B2(n_497), .Y(n_556) );
NAND3xp33_ASAP7_75t_SL g557 ( .A(n_519), .B(n_499), .C(n_498), .Y(n_557) );
AOI21xp33_ASAP7_75t_SL g558 ( .A1(n_524), .A2(n_470), .B(n_498), .Y(n_558) );
INVx1_ASAP7_75t_L g559 ( .A(n_503), .Y(n_559) );
INVx1_ASAP7_75t_SL g560 ( .A(n_519), .Y(n_560) );
INVx1_ASAP7_75t_L g561 ( .A(n_504), .Y(n_561) );
INVx2_ASAP7_75t_L g562 ( .A(n_507), .Y(n_562) );
OAI22xp33_ASAP7_75t_SL g563 ( .A1(n_535), .A2(n_497), .B1(n_493), .B2(n_486), .Y(n_563) );
INVx1_ASAP7_75t_L g564 ( .A(n_506), .Y(n_564) );
INVx1_ASAP7_75t_L g565 ( .A(n_502), .Y(n_565) );
AND2x2_ASAP7_75t_L g566 ( .A(n_510), .B(n_455), .Y(n_566) );
OR2x2_ASAP7_75t_L g567 ( .A(n_507), .B(n_479), .Y(n_567) );
O2A1O1Ixp33_ASAP7_75t_L g568 ( .A1(n_532), .A2(n_534), .B(n_524), .C(n_551), .Y(n_568) );
OAI21xp5_ASAP7_75t_L g569 ( .A1(n_528), .A2(n_493), .B(n_486), .Y(n_569) );
INVx1_ASAP7_75t_L g570 ( .A(n_514), .Y(n_570) );
INVx1_ASAP7_75t_L g571 ( .A(n_516), .Y(n_571) );
AOI21xp5_ASAP7_75t_L g572 ( .A1(n_501), .A2(n_471), .B(n_477), .Y(n_572) );
INVx1_ASAP7_75t_SL g573 ( .A(n_523), .Y(n_573) );
OR2x2_ASAP7_75t_L g574 ( .A(n_522), .B(n_479), .Y(n_574) );
OR2x2_ASAP7_75t_L g575 ( .A(n_521), .B(n_479), .Y(n_575) );
INVx1_ASAP7_75t_L g576 ( .A(n_527), .Y(n_576) );
INVx1_ASAP7_75t_L g577 ( .A(n_527), .Y(n_577) );
O2A1O1Ixp33_ASAP7_75t_L g578 ( .A1(n_552), .A2(n_496), .B(n_487), .C(n_455), .Y(n_578) );
OR2x6_ASAP7_75t_L g579 ( .A(n_547), .B(n_455), .Y(n_579) );
INVx1_ASAP7_75t_SL g580 ( .A(n_553), .Y(n_580) );
AOI22xp33_ASAP7_75t_SL g581 ( .A1(n_528), .A2(n_462), .B1(n_487), .B2(n_496), .Y(n_581) );
AOI22xp5_ASAP7_75t_L g582 ( .A1(n_543), .A2(n_466), .B1(n_462), .B2(n_484), .Y(n_582) );
INVx1_ASAP7_75t_L g583 ( .A(n_525), .Y(n_583) );
OAI21xp5_ASAP7_75t_L g584 ( .A1(n_541), .A2(n_491), .B(n_480), .Y(n_584) );
O2A1O1Ixp33_ASAP7_75t_SL g585 ( .A1(n_542), .A2(n_484), .B(n_469), .C(n_475), .Y(n_585) );
AND2x2_ASAP7_75t_L g586 ( .A(n_510), .B(n_484), .Y(n_586) );
OAI22xp5_ASAP7_75t_L g587 ( .A1(n_530), .A2(n_548), .B1(n_520), .B2(n_509), .Y(n_587) );
HB1xp67_ASAP7_75t_L g588 ( .A(n_529), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g589 ( .A(n_531), .B(n_491), .Y(n_589) );
INVx2_ASAP7_75t_L g590 ( .A(n_515), .Y(n_590) );
AOI32xp33_ASAP7_75t_L g591 ( .A1(n_529), .A2(n_339), .A3(n_346), .B1(n_36), .B2(n_40), .Y(n_591) );
INVx2_ASAP7_75t_SL g592 ( .A(n_511), .Y(n_592) );
AOI22xp5_ASAP7_75t_L g593 ( .A1(n_543), .A2(n_329), .B1(n_336), .B2(n_178), .Y(n_593) );
AOI221xp5_ASAP7_75t_L g594 ( .A1(n_517), .A2(n_257), .B1(n_336), .B2(n_42), .C(n_45), .Y(n_594) );
AND2x4_ASAP7_75t_SL g595 ( .A(n_517), .B(n_336), .Y(n_595) );
INVx2_ASAP7_75t_L g596 ( .A(n_515), .Y(n_596) );
INVxp67_ASAP7_75t_L g597 ( .A(n_550), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g598 ( .A(n_539), .B(n_30), .Y(n_598) );
OAI22xp33_ASAP7_75t_L g599 ( .A1(n_555), .A2(n_33), .B1(n_47), .B2(n_49), .Y(n_599) );
NOR2xp33_ASAP7_75t_L g600 ( .A(n_533), .B(n_50), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g601 ( .A(n_536), .B(n_51), .Y(n_601) );
INVx1_ASAP7_75t_L g602 ( .A(n_537), .Y(n_602) );
OAI222xp33_ASAP7_75t_L g603 ( .A1(n_560), .A2(n_540), .B1(n_533), .B2(n_500), .C1(n_550), .C2(n_549), .Y(n_603) );
XNOR2xp5_ASAP7_75t_L g604 ( .A(n_560), .B(n_512), .Y(n_604) );
INVx2_ASAP7_75t_L g605 ( .A(n_567), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g606 ( .A(n_587), .B(n_538), .Y(n_606) );
NAND2xp5_ASAP7_75t_SL g607 ( .A(n_563), .B(n_547), .Y(n_607) );
NOR2xp33_ASAP7_75t_L g608 ( .A(n_573), .B(n_553), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g609 ( .A(n_576), .B(n_545), .Y(n_609) );
NOR2xp33_ASAP7_75t_L g610 ( .A(n_573), .B(n_553), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g611 ( .A(n_577), .B(n_544), .Y(n_611) );
NOR3xp33_ASAP7_75t_SL g612 ( .A(n_557), .B(n_513), .C(n_554), .Y(n_612) );
INVx1_ASAP7_75t_L g613 ( .A(n_559), .Y(n_613) );
INVx2_ASAP7_75t_L g614 ( .A(n_562), .Y(n_614) );
OA21x2_ASAP7_75t_L g615 ( .A1(n_569), .A2(n_526), .B(n_545), .Y(n_615) );
NAND2xp5_ASAP7_75t_L g616 ( .A(n_565), .B(n_526), .Y(n_616) );
INVx1_ASAP7_75t_L g617 ( .A(n_561), .Y(n_617) );
OAI21xp33_ASAP7_75t_L g618 ( .A1(n_581), .A2(n_549), .B(n_546), .Y(n_618) );
INVx1_ASAP7_75t_L g619 ( .A(n_564), .Y(n_619) );
INVx2_ASAP7_75t_SL g620 ( .A(n_588), .Y(n_620) );
INVx3_ASAP7_75t_L g621 ( .A(n_579), .Y(n_621) );
OAI21xp5_ASAP7_75t_L g622 ( .A1(n_568), .A2(n_555), .B(n_546), .Y(n_622) );
OAI21xp33_ASAP7_75t_L g623 ( .A1(n_563), .A2(n_508), .B(n_540), .Y(n_623) );
OAI22xp5_ASAP7_75t_L g624 ( .A1(n_579), .A2(n_518), .B1(n_512), .B2(n_505), .Y(n_624) );
NAND2xp5_ASAP7_75t_SL g625 ( .A(n_558), .B(n_505), .Y(n_625) );
NAND2xp33_ASAP7_75t_L g626 ( .A(n_591), .B(n_329), .Y(n_626) );
NAND2xp33_ASAP7_75t_R g627 ( .A(n_579), .B(n_54), .Y(n_627) );
NAND4xp75_ASAP7_75t_L g628 ( .A(n_572), .B(n_57), .C(n_58), .D(n_61), .Y(n_628) );
INVx2_ASAP7_75t_L g629 ( .A(n_590), .Y(n_629) );
INVx2_ASAP7_75t_L g630 ( .A(n_596), .Y(n_630) );
INVx1_ASAP7_75t_L g631 ( .A(n_570), .Y(n_631) );
AOI21xp33_ASAP7_75t_L g632 ( .A1(n_578), .A2(n_70), .B(n_71), .Y(n_632) );
INVx2_ASAP7_75t_L g633 ( .A(n_575), .Y(n_633) );
A2O1A1Ixp33_ASAP7_75t_L g634 ( .A1(n_556), .A2(n_74), .B(n_76), .C(n_329), .Y(n_634) );
INVxp33_ASAP7_75t_L g635 ( .A(n_600), .Y(n_635) );
INVxp67_ASAP7_75t_L g636 ( .A(n_571), .Y(n_636) );
INVx2_ASAP7_75t_L g637 ( .A(n_602), .Y(n_637) );
INVx1_ASAP7_75t_SL g638 ( .A(n_620), .Y(n_638) );
XNOR2xp5_ASAP7_75t_L g639 ( .A(n_604), .B(n_583), .Y(n_639) );
CKINVDCx5p33_ASAP7_75t_R g640 ( .A(n_627), .Y(n_640) );
XNOR2x1_ASAP7_75t_L g641 ( .A(n_624), .B(n_566), .Y(n_641) );
NOR2xp33_ASAP7_75t_L g642 ( .A(n_635), .B(n_592), .Y(n_642) );
NAND2xp5_ASAP7_75t_L g643 ( .A(n_637), .B(n_574), .Y(n_643) );
XOR2x2_ASAP7_75t_SL g644 ( .A(n_627), .B(n_582), .Y(n_644) );
INVx1_ASAP7_75t_L g645 ( .A(n_613), .Y(n_645) );
INVx1_ASAP7_75t_L g646 ( .A(n_617), .Y(n_646) );
CKINVDCx20_ASAP7_75t_R g647 ( .A(n_633), .Y(n_647) );
INVx1_ASAP7_75t_L g648 ( .A(n_619), .Y(n_648) );
INVx1_ASAP7_75t_L g649 ( .A(n_631), .Y(n_649) );
XNOR2x1_ASAP7_75t_L g650 ( .A(n_621), .B(n_586), .Y(n_650) );
INVx1_ASAP7_75t_L g651 ( .A(n_606), .Y(n_651) );
AND2x2_ASAP7_75t_L g652 ( .A(n_605), .B(n_597), .Y(n_652) );
NAND2xp5_ASAP7_75t_L g653 ( .A(n_636), .B(n_589), .Y(n_653) );
INVxp67_ASAP7_75t_L g654 ( .A(n_608), .Y(n_654) );
NAND4xp75_ASAP7_75t_L g655 ( .A(n_607), .B(n_584), .C(n_594), .D(n_598), .Y(n_655) );
BUFx2_ASAP7_75t_L g656 ( .A(n_614), .Y(n_656) );
AND3x4_ASAP7_75t_L g657 ( .A(n_612), .B(n_585), .C(n_599), .Y(n_657) );
INVx1_ASAP7_75t_L g658 ( .A(n_616), .Y(n_658) );
AOI21xp33_ASAP7_75t_L g659 ( .A1(n_635), .A2(n_601), .B(n_580), .Y(n_659) );
INVx2_ASAP7_75t_SL g660 ( .A(n_608), .Y(n_660) );
AO22x2_ASAP7_75t_L g661 ( .A1(n_638), .A2(n_607), .B1(n_621), .B2(n_625), .Y(n_661) );
AOI22xp5_ASAP7_75t_L g662 ( .A1(n_640), .A2(n_626), .B1(n_623), .B2(n_610), .Y(n_662) );
AOI22xp5_ASAP7_75t_L g663 ( .A1(n_655), .A2(n_622), .B1(n_612), .B2(n_610), .Y(n_663) );
INVx2_ASAP7_75t_SL g664 ( .A(n_647), .Y(n_664) );
OAI211xp5_ASAP7_75t_SL g665 ( .A1(n_651), .A2(n_634), .B(n_618), .C(n_632), .Y(n_665) );
XNOR2xp5_ASAP7_75t_L g666 ( .A(n_639), .B(n_628), .Y(n_666) );
NOR2xp33_ASAP7_75t_L g667 ( .A(n_653), .B(n_603), .Y(n_667) );
INVx1_ASAP7_75t_SL g668 ( .A(n_656), .Y(n_668) );
BUFx2_ASAP7_75t_L g669 ( .A(n_644), .Y(n_669) );
INVx1_ASAP7_75t_L g670 ( .A(n_658), .Y(n_670) );
CKINVDCx5p33_ASAP7_75t_R g671 ( .A(n_642), .Y(n_671) );
AOI22xp5_ASAP7_75t_L g672 ( .A1(n_657), .A2(n_609), .B1(n_611), .B2(n_615), .Y(n_672) );
AOI211xp5_ASAP7_75t_L g673 ( .A1(n_659), .A2(n_580), .B(n_630), .C(n_629), .Y(n_673) );
OAI22xp5_ASAP7_75t_L g674 ( .A1(n_641), .A2(n_595), .B1(n_615), .B2(n_593), .Y(n_674) );
OAI22xp5_ASAP7_75t_L g675 ( .A1(n_650), .A2(n_290), .B1(n_329), .B2(n_654), .Y(n_675) );
OAI321xp33_ASAP7_75t_L g676 ( .A1(n_660), .A2(n_645), .A3(n_646), .B1(n_648), .B2(n_649), .C(n_643), .Y(n_676) );
AOI221xp5_ASAP7_75t_SL g677 ( .A1(n_652), .A2(n_654), .B1(n_639), .B2(n_607), .C(n_638), .Y(n_677) );
OAI22xp5_ASAP7_75t_L g678 ( .A1(n_659), .A2(n_640), .B1(n_560), .B2(n_647), .Y(n_678) );
INVx1_ASAP7_75t_L g679 ( .A(n_670), .Y(n_679) );
BUFx4f_ASAP7_75t_SL g680 ( .A(n_664), .Y(n_680) );
BUFx2_ASAP7_75t_L g681 ( .A(n_669), .Y(n_681) );
AOI22xp5_ASAP7_75t_L g682 ( .A1(n_677), .A2(n_674), .B1(n_663), .B2(n_678), .Y(n_682) );
HB1xp67_ASAP7_75t_L g683 ( .A(n_668), .Y(n_683) );
NAND5xp2_ASAP7_75t_L g684 ( .A(n_682), .B(n_663), .C(n_662), .D(n_676), .E(n_667), .Y(n_684) );
INVx1_ASAP7_75t_L g685 ( .A(n_683), .Y(n_685) );
AND3x1_ASAP7_75t_L g686 ( .A(n_681), .B(n_672), .C(n_673), .Y(n_686) );
BUFx2_ASAP7_75t_L g687 ( .A(n_685), .Y(n_687) );
OR3x1_ASAP7_75t_L g688 ( .A(n_684), .B(n_681), .C(n_665), .Y(n_688) );
HB1xp67_ASAP7_75t_L g689 ( .A(n_687), .Y(n_689) );
HB1xp67_ASAP7_75t_L g690 ( .A(n_688), .Y(n_690) );
AOI322xp5_ASAP7_75t_L g691 ( .A1(n_690), .A2(n_685), .A3(n_688), .B1(n_686), .B2(n_679), .C1(n_671), .C2(n_680), .Y(n_691) );
AOI221xp5_ASAP7_75t_L g692 ( .A1(n_691), .A2(n_689), .B1(n_661), .B2(n_666), .C(n_675), .Y(n_692) );
endmodule