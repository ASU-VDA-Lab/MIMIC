module fake_jpeg_17752_n_45 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_45);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_45;

wire n_21;
wire n_33;
wire n_23;
wire n_27;
wire n_22;
wire n_40;
wire n_19;
wire n_20;
wire n_35;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_31;
wire n_25;
wire n_29;
wire n_37;
wire n_43;
wire n_32;

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_16),
.B(n_5),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_2),
.B(n_11),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_17),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_1),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_2),
.B(n_10),
.Y(n_25)
);

AOI22xp33_ASAP7_75t_L g26 ( 
.A1(n_23),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_26)
);

XOR2xp5_ASAP7_75t_L g34 ( 
.A(n_26),
.B(n_28),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_19),
.B(n_0),
.Y(n_27)
);

OAI21xp5_ASAP7_75t_L g33 ( 
.A1(n_27),
.A2(n_31),
.B(n_20),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_L g28 ( 
.A1(n_19),
.A2(n_8),
.B1(n_15),
.B2(n_13),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_24),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_29),
.B(n_30),
.Y(n_32)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_22),
.Y(n_30)
);

CKINVDCx14_ASAP7_75t_R g31 ( 
.A(n_25),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_SL g39 ( 
.A(n_33),
.B(n_3),
.Y(n_39)
);

MAJIxp5_ASAP7_75t_L g35 ( 
.A(n_29),
.B(n_24),
.C(n_21),
.Y(n_35)
);

XOR2xp5_ASAP7_75t_L g37 ( 
.A(n_35),
.B(n_36),
.Y(n_37)
);

XNOR2xp5_ASAP7_75t_L g36 ( 
.A(n_27),
.B(n_28),
.Y(n_36)
);

BUFx24_ASAP7_75t_SL g38 ( 
.A(n_34),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_SL g41 ( 
.A(n_38),
.B(n_39),
.Y(n_41)
);

XNOR2xp5_ASAP7_75t_L g40 ( 
.A(n_37),
.B(n_34),
.Y(n_40)
);

OAI21xp5_ASAP7_75t_SL g42 ( 
.A1(n_40),
.A2(n_32),
.B(n_22),
.Y(n_42)
);

O2A1O1Ixp33_ASAP7_75t_SL g43 ( 
.A1(n_42),
.A2(n_41),
.B(n_30),
.C(n_6),
.Y(n_43)
);

OAI21x1_ASAP7_75t_L g44 ( 
.A1(n_43),
.A2(n_4),
.B(n_5),
.Y(n_44)
);

OAI321xp33_ASAP7_75t_L g45 ( 
.A1(n_44),
.A2(n_4),
.A3(n_6),
.B1(n_7),
.B2(n_12),
.C(n_18),
.Y(n_45)
);


endmodule