module fake_jpeg_12077_n_561 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_561);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_561;

wire n_529;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_349;
wire n_21;
wire n_288;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_7),
.Y(n_19)
);

INVx4_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_8),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

BUFx24_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

INVx5_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_7),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_11),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_9),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_6),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_15),
.Y(n_35)
);

INVxp67_ASAP7_75t_L g36 ( 
.A(n_2),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_14),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_0),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_12),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_6),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_10),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_18),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_1),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_10),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_9),
.Y(n_45)
);

INVx11_ASAP7_75t_L g46 ( 
.A(n_7),
.Y(n_46)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_15),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_16),
.Y(n_48)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_1),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_10),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_13),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_0),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_11),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_11),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_2),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_3),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_1),
.Y(n_57)
);

INVx11_ASAP7_75t_SL g58 ( 
.A(n_6),
.Y(n_58)
);

INVx1_ASAP7_75t_SL g59 ( 
.A(n_24),
.Y(n_59)
);

INVx13_ASAP7_75t_L g144 ( 
.A(n_59),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_46),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_60),
.B(n_61),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_46),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_22),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_62),
.Y(n_129)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_24),
.Y(n_63)
);

INVx5_ASAP7_75t_L g138 ( 
.A(n_63),
.Y(n_138)
);

BUFx2_ASAP7_75t_L g64 ( 
.A(n_24),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g140 ( 
.A(n_64),
.Y(n_140)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_27),
.Y(n_65)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_65),
.Y(n_139)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_26),
.Y(n_66)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_66),
.Y(n_130)
);

INVx2_ASAP7_75t_SL g67 ( 
.A(n_24),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g204 ( 
.A(n_67),
.Y(n_204)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_22),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_68),
.Y(n_131)
);

BUFx16f_ASAP7_75t_L g69 ( 
.A(n_28),
.Y(n_69)
);

CKINVDCx16_ASAP7_75t_R g142 ( 
.A(n_69),
.Y(n_142)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_28),
.Y(n_70)
);

INVx4_ASAP7_75t_L g143 ( 
.A(n_70),
.Y(n_143)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_27),
.Y(n_71)
);

INVx3_ASAP7_75t_L g152 ( 
.A(n_71),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_37),
.B(n_18),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_72),
.B(n_77),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_37),
.B(n_18),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_73),
.B(n_84),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_46),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_74),
.B(n_83),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_22),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_75),
.Y(n_156)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_26),
.Y(n_76)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_76),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_35),
.B(n_17),
.Y(n_77)
);

INVx8_ASAP7_75t_L g78 ( 
.A(n_23),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g170 ( 
.A(n_78),
.Y(n_170)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_47),
.Y(n_79)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_79),
.Y(n_160)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_28),
.Y(n_80)
);

INVx4_ASAP7_75t_L g147 ( 
.A(n_80),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_35),
.B(n_17),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g199 ( 
.A(n_81),
.B(n_97),
.Y(n_199)
);

INVx8_ASAP7_75t_L g82 ( 
.A(n_23),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g180 ( 
.A(n_82),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_48),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_19),
.B(n_17),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_23),
.Y(n_85)
);

INVx6_ASAP7_75t_L g145 ( 
.A(n_85),
.Y(n_145)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_48),
.Y(n_86)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_86),
.Y(n_132)
);

BUFx12_ASAP7_75t_L g87 ( 
.A(n_58),
.Y(n_87)
);

INVx2_ASAP7_75t_SL g197 ( 
.A(n_87),
.Y(n_197)
);

BUFx16f_ASAP7_75t_L g88 ( 
.A(n_28),
.Y(n_88)
);

INVx3_ASAP7_75t_L g207 ( 
.A(n_88),
.Y(n_207)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_32),
.Y(n_89)
);

INVx6_ASAP7_75t_L g188 ( 
.A(n_89),
.Y(n_188)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_47),
.Y(n_90)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_90),
.Y(n_137)
);

INVx1_ASAP7_75t_SL g91 ( 
.A(n_52),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_91),
.B(n_92),
.Y(n_149)
);

NAND2xp33_ASAP7_75t_SL g92 ( 
.A(n_36),
.B(n_0),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_19),
.B(n_16),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_93),
.B(n_99),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_32),
.Y(n_94)
);

INVx8_ASAP7_75t_L g163 ( 
.A(n_94),
.Y(n_163)
);

INVx8_ASAP7_75t_L g95 ( 
.A(n_32),
.Y(n_95)
);

INVx3_ASAP7_75t_SL g134 ( 
.A(n_95),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_21),
.B(n_16),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_96),
.B(n_102),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_21),
.B(n_14),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_38),
.Y(n_98)
);

INVx3_ASAP7_75t_SL g208 ( 
.A(n_98),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_20),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_38),
.Y(n_100)
);

INVx4_ASAP7_75t_L g155 ( 
.A(n_100),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_38),
.Y(n_101)
);

INVx4_ASAP7_75t_L g174 ( 
.A(n_101),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_30),
.B(n_14),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_20),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_103),
.B(n_108),
.Y(n_159)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_20),
.Y(n_104)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_104),
.Y(n_172)
);

INVx5_ASAP7_75t_L g105 ( 
.A(n_25),
.Y(n_105)
);

INVx4_ASAP7_75t_L g183 ( 
.A(n_105),
.Y(n_183)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_41),
.Y(n_106)
);

INVx4_ASAP7_75t_L g184 ( 
.A(n_106),
.Y(n_184)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_39),
.Y(n_107)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_107),
.Y(n_175)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_39),
.Y(n_108)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_43),
.Y(n_109)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_109),
.Y(n_176)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_27),
.Y(n_110)
);

INVx4_ASAP7_75t_L g186 ( 
.A(n_110),
.Y(n_186)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_43),
.Y(n_111)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_111),
.Y(n_141)
);

BUFx12f_ASAP7_75t_L g112 ( 
.A(n_41),
.Y(n_112)
);

INVx4_ASAP7_75t_L g189 ( 
.A(n_112),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_41),
.Y(n_113)
);

INVx4_ASAP7_75t_L g200 ( 
.A(n_113),
.Y(n_200)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_56),
.Y(n_114)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_114),
.Y(n_182)
);

INVx2_ASAP7_75t_R g115 ( 
.A(n_30),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_115),
.B(n_124),
.Y(n_167)
);

INVx8_ASAP7_75t_L g116 ( 
.A(n_44),
.Y(n_116)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_116),
.Y(n_185)
);

INVx4_ASAP7_75t_L g117 ( 
.A(n_52),
.Y(n_117)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_117),
.Y(n_187)
);

INVx6_ASAP7_75t_L g118 ( 
.A(n_44),
.Y(n_118)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_118),
.Y(n_191)
);

INVx8_ASAP7_75t_L g119 ( 
.A(n_44),
.Y(n_119)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_119),
.Y(n_194)
);

INVx6_ASAP7_75t_L g120 ( 
.A(n_51),
.Y(n_120)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_120),
.Y(n_195)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_51),
.Y(n_121)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_121),
.Y(n_196)
);

INVx8_ASAP7_75t_L g122 ( 
.A(n_51),
.Y(n_122)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_122),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_31),
.B(n_0),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_123),
.B(n_1),
.Y(n_166)
);

BUFx3_ASAP7_75t_L g124 ( 
.A(n_52),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_56),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_125),
.B(n_45),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_118),
.A2(n_42),
.B1(n_29),
.B2(n_49),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g264 ( 
.A1(n_126),
.A2(n_133),
.B1(n_135),
.B2(n_153),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_120),
.A2(n_42),
.B1(n_29),
.B2(n_49),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_62),
.A2(n_42),
.B1(n_29),
.B2(n_49),
.Y(n_135)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_108),
.Y(n_150)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_150),
.Y(n_211)
);

AOI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_59),
.A2(n_25),
.B1(n_53),
.B2(n_52),
.Y(n_153)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_104),
.Y(n_158)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_158),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_75),
.A2(n_53),
.B1(n_57),
.B2(n_33),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_161),
.A2(n_164),
.B1(n_190),
.B2(n_193),
.Y(n_253)
);

AOI22xp33_ASAP7_75t_SL g162 ( 
.A1(n_63),
.A2(n_53),
.B1(n_57),
.B2(n_33),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_SL g209 ( 
.A1(n_162),
.A2(n_179),
.B1(n_67),
.B2(n_124),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_85),
.A2(n_55),
.B1(n_54),
.B2(n_50),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_L g165 ( 
.A1(n_89),
.A2(n_55),
.B1(n_54),
.B2(n_50),
.Y(n_165)
);

OA22x2_ASAP7_75t_L g230 ( 
.A1(n_165),
.A2(n_173),
.B1(n_177),
.B2(n_201),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_166),
.B(n_192),
.Y(n_274)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_115),
.Y(n_168)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_168),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_169),
.B(n_199),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_69),
.B(n_45),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_SL g212 ( 
.A(n_171),
.B(n_178),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_94),
.A2(n_40),
.B1(n_34),
.B2(n_31),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_L g177 ( 
.A1(n_98),
.A2(n_40),
.B1(n_34),
.B2(n_4),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_69),
.B(n_2),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_SL g179 ( 
.A1(n_64),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_88),
.B(n_92),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_SL g252 ( 
.A(n_181),
.B(n_198),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_100),
.A2(n_13),
.B1(n_4),
.B2(n_5),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_91),
.B(n_3),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_101),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_87),
.Y(n_198)
);

OAI22xp33_ASAP7_75t_SL g201 ( 
.A1(n_106),
.A2(n_5),
.B1(n_9),
.B2(n_12),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_88),
.B(n_5),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_202),
.B(n_205),
.Y(n_213)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_65),
.Y(n_203)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_203),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_70),
.B(n_9),
.Y(n_205)
);

OAI22xp33_ASAP7_75t_SL g206 ( 
.A1(n_113),
.A2(n_12),
.B1(n_13),
.B2(n_121),
.Y(n_206)
);

AO22x1_ASAP7_75t_L g261 ( 
.A1(n_206),
.A2(n_201),
.B1(n_177),
.B2(n_165),
.Y(n_261)
);

INVxp67_ASAP7_75t_L g301 ( 
.A(n_209),
.Y(n_301)
);

INVx6_ASAP7_75t_L g210 ( 
.A(n_129),
.Y(n_210)
);

BUFx6f_ASAP7_75t_L g305 ( 
.A(n_210),
.Y(n_305)
);

AND2x2_ASAP7_75t_L g214 ( 
.A(n_149),
.B(n_117),
.Y(n_214)
);

OAI21xp33_ASAP7_75t_L g314 ( 
.A1(n_214),
.A2(n_217),
.B(n_233),
.Y(n_314)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_191),
.Y(n_216)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_216),
.Y(n_280)
);

AND2x2_ASAP7_75t_L g217 ( 
.A(n_160),
.B(n_71),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_218),
.B(n_224),
.Y(n_303)
);

INVx8_ASAP7_75t_L g220 ( 
.A(n_131),
.Y(n_220)
);

BUFx2_ASAP7_75t_L g292 ( 
.A(n_220),
.Y(n_292)
);

INVx5_ASAP7_75t_L g221 ( 
.A(n_207),
.Y(n_221)
);

BUFx2_ASAP7_75t_L g296 ( 
.A(n_221),
.Y(n_296)
);

INVx6_ASAP7_75t_L g222 ( 
.A(n_129),
.Y(n_222)
);

INVx3_ASAP7_75t_L g307 ( 
.A(n_222),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_136),
.B(n_110),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_223),
.B(n_258),
.Y(n_286)
);

CKINVDCx14_ASAP7_75t_R g224 ( 
.A(n_144),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_148),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_225),
.B(n_237),
.Y(n_310)
);

INVx8_ASAP7_75t_L g227 ( 
.A(n_131),
.Y(n_227)
);

INVx3_ASAP7_75t_L g312 ( 
.A(n_227),
.Y(n_312)
);

INVx4_ASAP7_75t_L g228 ( 
.A(n_189),
.Y(n_228)
);

INVx3_ASAP7_75t_L g313 ( 
.A(n_228),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_157),
.B(n_105),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g331 ( 
.A(n_229),
.B(n_231),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_151),
.B(n_80),
.Y(n_231)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_195),
.Y(n_232)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_232),
.Y(n_284)
);

AND2x2_ASAP7_75t_L g233 ( 
.A(n_130),
.B(n_112),
.Y(n_233)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_196),
.Y(n_234)
);

INVx2_ASAP7_75t_L g306 ( 
.A(n_234),
.Y(n_306)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_132),
.Y(n_235)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_235),
.Y(n_281)
);

INVx4_ASAP7_75t_L g236 ( 
.A(n_189),
.Y(n_236)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_236),
.Y(n_315)
);

INVxp67_ASAP7_75t_L g237 ( 
.A(n_167),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_128),
.B(n_112),
.Y(n_238)
);

INVxp67_ASAP7_75t_L g316 ( 
.A(n_238),
.Y(n_316)
);

INVx3_ASAP7_75t_L g239 ( 
.A(n_140),
.Y(n_239)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_239),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_127),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_240),
.B(n_243),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_159),
.B(n_68),
.Y(n_241)
);

INVxp67_ASAP7_75t_L g320 ( 
.A(n_241),
.Y(n_320)
);

INVx4_ASAP7_75t_L g242 ( 
.A(n_140),
.Y(n_242)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_242),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_141),
.Y(n_243)
);

A2O1A1Ixp33_ASAP7_75t_L g244 ( 
.A1(n_137),
.A2(n_87),
.B(n_122),
.C(n_78),
.Y(n_244)
);

NOR2x1_ASAP7_75t_L g294 ( 
.A(n_244),
.B(n_277),
.Y(n_294)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_139),
.Y(n_245)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_245),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_142),
.B(n_82),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_246),
.B(n_249),
.Y(n_327)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_175),
.Y(n_247)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_247),
.Y(n_332)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_176),
.Y(n_248)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_248),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_154),
.B(n_95),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_204),
.B(n_116),
.Y(n_250)
);

CKINVDCx16_ASAP7_75t_R g288 ( 
.A(n_250),
.Y(n_288)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_182),
.Y(n_251)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_251),
.Y(n_289)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_139),
.Y(n_254)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_254),
.Y(n_290)
);

INVx3_ASAP7_75t_L g255 ( 
.A(n_185),
.Y(n_255)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_255),
.Y(n_295)
);

BUFx2_ASAP7_75t_L g256 ( 
.A(n_138),
.Y(n_256)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_256),
.Y(n_298)
);

INVxp67_ASAP7_75t_L g257 ( 
.A(n_144),
.Y(n_257)
);

CKINVDCx16_ASAP7_75t_R g319 ( 
.A(n_257),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_172),
.B(n_119),
.Y(n_258)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_152),
.Y(n_259)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_259),
.Y(n_318)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_146),
.Y(n_260)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_260),
.Y(n_322)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_261),
.A2(n_208),
.B1(n_145),
.B2(n_188),
.Y(n_282)
);

AOI22xp33_ASAP7_75t_L g262 ( 
.A1(n_206),
.A2(n_174),
.B1(n_200),
.B2(n_184),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_L g304 ( 
.A1(n_262),
.A2(n_156),
.B1(n_273),
.B2(n_253),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_186),
.B(n_187),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_263),
.B(n_265),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_186),
.B(n_152),
.Y(n_265)
);

INVx3_ASAP7_75t_L g266 ( 
.A(n_194),
.Y(n_266)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_266),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_163),
.B(n_174),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_267),
.B(n_269),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_204),
.B(n_207),
.Y(n_268)
);

AND2x2_ASAP7_75t_L g328 ( 
.A(n_268),
.B(n_270),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_163),
.B(n_200),
.Y(n_269)
);

BUFx3_ASAP7_75t_L g270 ( 
.A(n_197),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_197),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_271),
.Y(n_291)
);

AND2x2_ASAP7_75t_SL g272 ( 
.A(n_143),
.B(n_147),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g330 ( 
.A(n_272),
.B(n_273),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_153),
.B(n_133),
.C(n_134),
.Y(n_273)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_155),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_275),
.Y(n_302)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_155),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_276),
.Y(n_333)
);

AOI21xp33_ASAP7_75t_SL g277 ( 
.A1(n_143),
.A2(n_147),
.B(n_138),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_179),
.B(n_162),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_278),
.B(n_279),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_208),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_L g337 ( 
.A1(n_282),
.A2(n_308),
.B1(n_210),
.B2(n_222),
.Y(n_337)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_253),
.A2(n_188),
.B1(n_145),
.B2(n_184),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g340 ( 
.A1(n_287),
.A2(n_304),
.B1(n_317),
.B2(n_272),
.Y(n_340)
);

AOI21xp5_ASAP7_75t_L g293 ( 
.A1(n_278),
.A2(n_183),
.B(n_134),
.Y(n_293)
);

AOI21xp5_ASAP7_75t_L g361 ( 
.A1(n_293),
.A2(n_242),
.B(n_228),
.Y(n_361)
);

OAI21xp5_ASAP7_75t_L g297 ( 
.A1(n_252),
.A2(n_170),
.B(n_180),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_L g342 ( 
.A1(n_297),
.A2(n_309),
.B(n_233),
.Y(n_342)
);

AOI22xp33_ASAP7_75t_SL g299 ( 
.A1(n_237),
.A2(n_183),
.B1(n_170),
.B2(n_180),
.Y(n_299)
);

CKINVDCx14_ASAP7_75t_R g356 ( 
.A(n_299),
.Y(n_356)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_264),
.A2(n_156),
.B1(n_261),
.B2(n_230),
.Y(n_308)
);

O2A1O1Ixp33_ASAP7_75t_L g309 ( 
.A1(n_244),
.A2(n_214),
.B(n_272),
.C(n_257),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_223),
.A2(n_230),
.B1(n_213),
.B2(n_274),
.Y(n_317)
);

FAx1_ASAP7_75t_SL g329 ( 
.A(n_214),
.B(n_263),
.CI(n_265),
.CON(n_329),
.SN(n_329)
);

NOR2xp33_ASAP7_75t_SL g364 ( 
.A(n_329),
.B(n_236),
.Y(n_364)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_321),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_334),
.B(n_345),
.Y(n_376)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_285),
.Y(n_335)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_335),
.Y(n_380)
);

OAI22xp5_ASAP7_75t_SL g336 ( 
.A1(n_308),
.A2(n_230),
.B1(n_269),
.B2(n_267),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_L g393 ( 
.A1(n_336),
.A2(n_337),
.B1(n_339),
.B2(n_341),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_SL g338 ( 
.A(n_310),
.B(n_219),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_SL g395 ( 
.A(n_338),
.B(n_346),
.Y(n_395)
);

OAI22xp5_ASAP7_75t_L g339 ( 
.A1(n_293),
.A2(n_230),
.B1(n_212),
.B2(n_220),
.Y(n_339)
);

OAI22xp5_ASAP7_75t_L g391 ( 
.A1(n_340),
.A2(n_348),
.B1(n_374),
.B2(n_366),
.Y(n_391)
);

OAI22xp5_ASAP7_75t_L g341 ( 
.A1(n_323),
.A2(n_227),
.B1(n_232),
.B2(n_216),
.Y(n_341)
);

OAI21xp5_ASAP7_75t_SL g382 ( 
.A1(n_342),
.A2(n_344),
.B(n_361),
.Y(n_382)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_285),
.Y(n_343)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_343),
.Y(n_396)
);

A2O1A1O1Ixp25_ASAP7_75t_L g344 ( 
.A1(n_325),
.A2(n_215),
.B(n_211),
.C(n_226),
.D(n_217),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_317),
.B(n_217),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_331),
.B(n_270),
.Y(n_346)
);

OAI22xp5_ASAP7_75t_SL g347 ( 
.A1(n_325),
.A2(n_234),
.B1(n_266),
.B2(n_255),
.Y(n_347)
);

AOI22xp5_ASAP7_75t_SL g389 ( 
.A1(n_347),
.A2(n_351),
.B1(n_375),
.B2(n_324),
.Y(n_389)
);

AOI22xp5_ASAP7_75t_L g348 ( 
.A1(n_287),
.A2(n_233),
.B1(n_259),
.B2(n_245),
.Y(n_348)
);

BUFx24_ASAP7_75t_SL g349 ( 
.A(n_303),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_SL g403 ( 
.A(n_349),
.B(n_363),
.Y(n_403)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_289),
.Y(n_350)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_350),
.Y(n_405)
);

OAI22xp5_ASAP7_75t_SL g351 ( 
.A1(n_323),
.A2(n_254),
.B1(n_275),
.B2(n_276),
.Y(n_351)
);

INVx2_ASAP7_75t_L g352 ( 
.A(n_280),
.Y(n_352)
);

HB1xp67_ASAP7_75t_L g409 ( 
.A(n_352),
.Y(n_409)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_289),
.Y(n_353)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_353),
.Y(n_394)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_290),
.Y(n_354)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_354),
.Y(n_404)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_290),
.Y(n_355)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_355),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_286),
.B(n_256),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_357),
.B(n_359),
.Y(n_377)
);

XNOR2xp5_ASAP7_75t_SL g358 ( 
.A(n_330),
.B(n_221),
.Y(n_358)
);

XNOR2xp5_ASAP7_75t_SL g385 ( 
.A(n_358),
.B(n_372),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_286),
.B(n_239),
.Y(n_359)
);

INVx2_ASAP7_75t_L g360 ( 
.A(n_280),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_360),
.B(n_362),
.Y(n_388)
);

CKINVDCx20_ASAP7_75t_R g362 ( 
.A(n_291),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_318),
.Y(n_363)
);

XOR2x2_ASAP7_75t_SL g397 ( 
.A(n_364),
.B(n_365),
.Y(n_397)
);

AND2x2_ASAP7_75t_L g365 ( 
.A(n_309),
.B(n_314),
.Y(n_365)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_328),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_366),
.B(n_367),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_SL g367 ( 
.A(n_300),
.B(n_320),
.Y(n_367)
);

CKINVDCx20_ASAP7_75t_R g368 ( 
.A(n_328),
.Y(n_368)
);

CKINVDCx20_ASAP7_75t_R g378 ( 
.A(n_368),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_300),
.B(n_329),
.Y(n_369)
);

XNOR2xp5_ASAP7_75t_L g379 ( 
.A(n_369),
.B(n_297),
.Y(n_379)
);

MAJx2_ASAP7_75t_L g370 ( 
.A(n_330),
.B(n_327),
.C(n_316),
.Y(n_370)
);

MAJIxp5_ASAP7_75t_L g384 ( 
.A(n_370),
.B(n_322),
.C(n_332),
.Y(n_384)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_318),
.Y(n_371)
);

AOI22xp33_ASAP7_75t_SL g381 ( 
.A1(n_371),
.A2(n_292),
.B1(n_296),
.B2(n_301),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_SL g372 ( 
.A(n_288),
.B(n_320),
.Y(n_372)
);

INVx1_ASAP7_75t_SL g373 ( 
.A(n_328),
.Y(n_373)
);

BUFx24_ASAP7_75t_L g401 ( 
.A(n_373),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_L g374 ( 
.A(n_281),
.B(n_316),
.Y(n_374)
);

OAI22xp5_ASAP7_75t_SL g375 ( 
.A1(n_301),
.A2(n_282),
.B1(n_294),
.B2(n_329),
.Y(n_375)
);

XNOR2xp5_ASAP7_75t_L g413 ( 
.A(n_379),
.B(n_384),
.Y(n_413)
);

INVxp67_ASAP7_75t_L g419 ( 
.A(n_381),
.Y(n_419)
);

OAI22xp5_ASAP7_75t_SL g383 ( 
.A1(n_340),
.A2(n_294),
.B1(n_307),
.B2(n_322),
.Y(n_383)
);

AOI22xp5_ASAP7_75t_L g414 ( 
.A1(n_383),
.A2(n_386),
.B1(n_391),
.B2(n_400),
.Y(n_414)
);

OAI22xp33_ASAP7_75t_SL g386 ( 
.A1(n_373),
.A2(n_312),
.B1(n_292),
.B2(n_307),
.Y(n_386)
);

MAJIxp5_ASAP7_75t_L g387 ( 
.A(n_358),
.B(n_283),
.C(n_324),
.Y(n_387)
);

MAJIxp5_ASAP7_75t_L g428 ( 
.A(n_387),
.B(n_390),
.C(n_392),
.Y(n_428)
);

OAI22xp33_ASAP7_75t_SL g411 ( 
.A1(n_389),
.A2(n_348),
.B1(n_336),
.B2(n_337),
.Y(n_411)
);

MAJIxp5_ASAP7_75t_L g390 ( 
.A(n_370),
.B(n_283),
.C(n_295),
.Y(n_390)
);

XNOR2xp5_ASAP7_75t_L g392 ( 
.A(n_369),
.B(n_295),
.Y(n_392)
);

XNOR2xp5_ASAP7_75t_L g398 ( 
.A(n_367),
.B(n_311),
.Y(n_398)
);

XNOR2xp5_ASAP7_75t_L g417 ( 
.A(n_398),
.B(n_399),
.Y(n_417)
);

MAJIxp5_ASAP7_75t_L g399 ( 
.A(n_365),
.B(n_326),
.C(n_319),
.Y(n_399)
);

OAI22xp5_ASAP7_75t_SL g400 ( 
.A1(n_345),
.A2(n_312),
.B1(n_305),
.B2(n_298),
.Y(n_400)
);

MAJIxp5_ASAP7_75t_L g406 ( 
.A(n_365),
.B(n_368),
.C(n_361),
.Y(n_406)
);

INVxp67_ASAP7_75t_L g422 ( 
.A(n_406),
.Y(n_422)
);

OAI22xp5_ASAP7_75t_L g408 ( 
.A1(n_357),
.A2(n_305),
.B1(n_302),
.B2(n_333),
.Y(n_408)
);

AOI22xp5_ASAP7_75t_L g421 ( 
.A1(n_408),
.A2(n_341),
.B1(n_351),
.B2(n_347),
.Y(n_421)
);

OAI21xp5_ASAP7_75t_SL g410 ( 
.A1(n_406),
.A2(n_356),
.B(n_342),
.Y(n_410)
);

OAI21xp5_ASAP7_75t_L g442 ( 
.A1(n_410),
.A2(n_416),
.B(n_436),
.Y(n_442)
);

AOI22xp5_ASAP7_75t_L g456 ( 
.A1(n_411),
.A2(n_425),
.B1(n_426),
.B2(n_400),
.Y(n_456)
);

CKINVDCx20_ASAP7_75t_R g412 ( 
.A(n_388),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_412),
.B(n_415),
.Y(n_447)
);

OA21x2_ASAP7_75t_L g415 ( 
.A1(n_383),
.A2(n_375),
.B(n_359),
.Y(n_415)
);

OAI21xp5_ASAP7_75t_SL g416 ( 
.A1(n_382),
.A2(n_362),
.B(n_344),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_L g418 ( 
.A(n_378),
.B(n_334),
.Y(n_418)
);

CKINVDCx14_ASAP7_75t_R g441 ( 
.A(n_418),
.Y(n_441)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_394),
.Y(n_420)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_420),
.Y(n_452)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_421),
.Y(n_459)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_394),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_SL g461 ( 
.A(n_423),
.B(n_424),
.Y(n_461)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_404),
.Y(n_424)
);

OA21x2_ASAP7_75t_L g425 ( 
.A1(n_393),
.A2(n_339),
.B(n_364),
.Y(n_425)
);

OAI22xp5_ASAP7_75t_SL g426 ( 
.A1(n_393),
.A2(n_389),
.B1(n_376),
.B2(n_377),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_404),
.Y(n_427)
);

CKINVDCx20_ASAP7_75t_R g445 ( 
.A(n_427),
.Y(n_445)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_407),
.Y(n_429)
);

CKINVDCx20_ASAP7_75t_R g462 ( 
.A(n_429),
.Y(n_462)
);

NOR2xp33_ASAP7_75t_L g430 ( 
.A(n_403),
.B(n_296),
.Y(n_430)
);

NOR2xp33_ASAP7_75t_SL g449 ( 
.A(n_430),
.B(n_395),
.Y(n_449)
);

OR2x2_ASAP7_75t_L g431 ( 
.A(n_397),
.B(n_350),
.Y(n_431)
);

CKINVDCx20_ASAP7_75t_R g463 ( 
.A(n_431),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_377),
.B(n_353),
.Y(n_432)
);

AO21x1_ASAP7_75t_L g443 ( 
.A1(n_432),
.A2(n_434),
.B(n_435),
.Y(n_443)
);

INVx2_ASAP7_75t_L g433 ( 
.A(n_407),
.Y(n_433)
);

CKINVDCx16_ASAP7_75t_R g450 ( 
.A(n_433),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_376),
.B(n_343),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_402),
.B(n_388),
.Y(n_435)
);

AOI22xp33_ASAP7_75t_SL g436 ( 
.A1(n_401),
.A2(n_371),
.B1(n_363),
.B2(n_355),
.Y(n_436)
);

AND2x2_ASAP7_75t_L g437 ( 
.A(n_401),
.B(n_354),
.Y(n_437)
);

CKINVDCx20_ASAP7_75t_R g453 ( 
.A(n_437),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_402),
.B(n_335),
.Y(n_438)
);

CKINVDCx20_ASAP7_75t_R g457 ( 
.A(n_438),
.Y(n_457)
);

CKINVDCx20_ASAP7_75t_R g439 ( 
.A(n_409),
.Y(n_439)
);

CKINVDCx16_ASAP7_75t_R g455 ( 
.A(n_439),
.Y(n_455)
);

XOR2xp5_ASAP7_75t_L g440 ( 
.A(n_413),
.B(n_385),
.Y(n_440)
);

XOR2xp5_ASAP7_75t_L g477 ( 
.A(n_440),
.B(n_451),
.Y(n_477)
);

XNOR2xp5_ASAP7_75t_SL g444 ( 
.A(n_413),
.B(n_385),
.Y(n_444)
);

XNOR2xp5_ASAP7_75t_SL g470 ( 
.A(n_444),
.B(n_446),
.Y(n_470)
);

XNOR2xp5_ASAP7_75t_SL g446 ( 
.A(n_417),
.B(n_398),
.Y(n_446)
);

XOR2x2_ASAP7_75t_L g448 ( 
.A(n_422),
.B(n_379),
.Y(n_448)
);

NOR2xp33_ASAP7_75t_L g476 ( 
.A(n_448),
.B(n_415),
.Y(n_476)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_449),
.Y(n_468)
);

XNOR2xp5_ASAP7_75t_SL g451 ( 
.A(n_417),
.B(n_392),
.Y(n_451)
);

XOR2xp5_ASAP7_75t_L g454 ( 
.A(n_428),
.B(n_387),
.Y(n_454)
);

XOR2xp5_ASAP7_75t_L g483 ( 
.A(n_454),
.B(n_458),
.Y(n_483)
);

OAI22xp5_ASAP7_75t_L g482 ( 
.A1(n_456),
.A2(n_432),
.B1(n_421),
.B2(n_439),
.Y(n_482)
);

XNOR2xp5_ASAP7_75t_L g458 ( 
.A(n_428),
.B(n_397),
.Y(n_458)
);

OAI21xp5_ASAP7_75t_L g460 ( 
.A1(n_431),
.A2(n_382),
.B(n_401),
.Y(n_460)
);

AOI21xp5_ASAP7_75t_L g481 ( 
.A1(n_460),
.A2(n_435),
.B(n_437),
.Y(n_481)
);

OAI22xp5_ASAP7_75t_SL g464 ( 
.A1(n_414),
.A2(n_390),
.B1(n_399),
.B2(n_384),
.Y(n_464)
);

AOI22xp5_ASAP7_75t_L g467 ( 
.A1(n_464),
.A2(n_415),
.B1(n_426),
.B2(n_425),
.Y(n_467)
);

MAJIxp5_ASAP7_75t_L g465 ( 
.A(n_410),
.B(n_405),
.C(n_396),
.Y(n_465)
);

MAJIxp5_ASAP7_75t_L g480 ( 
.A(n_465),
.B(n_437),
.C(n_420),
.Y(n_480)
);

XOR2xp5_ASAP7_75t_L g466 ( 
.A(n_431),
.B(n_380),
.Y(n_466)
);

XOR2xp5_ASAP7_75t_L g484 ( 
.A(n_466),
.B(n_429),
.Y(n_484)
);

MAJIxp5_ASAP7_75t_L g496 ( 
.A(n_467),
.B(n_480),
.C(n_486),
.Y(n_496)
);

NOR2xp33_ASAP7_75t_SL g469 ( 
.A(n_458),
.B(n_418),
.Y(n_469)
);

NOR2xp33_ASAP7_75t_L g500 ( 
.A(n_469),
.B(n_472),
.Y(n_500)
);

AOI22xp5_ASAP7_75t_L g471 ( 
.A1(n_459),
.A2(n_425),
.B1(n_415),
.B2(n_412),
.Y(n_471)
);

OAI22xp5_ASAP7_75t_SL g494 ( 
.A1(n_471),
.A2(n_473),
.B1(n_478),
.B2(n_456),
.Y(n_494)
);

CKINVDCx16_ASAP7_75t_R g472 ( 
.A(n_447),
.Y(n_472)
);

AOI22xp33_ASAP7_75t_SL g473 ( 
.A1(n_459),
.A2(n_419),
.B1(n_427),
.B2(n_424),
.Y(n_473)
);

OR2x2_ASAP7_75t_L g474 ( 
.A(n_441),
.B(n_416),
.Y(n_474)
);

AOI21xp5_ASAP7_75t_L g495 ( 
.A1(n_474),
.A2(n_442),
.B(n_443),
.Y(n_495)
);

AND2x2_ASAP7_75t_L g475 ( 
.A(n_453),
.B(n_414),
.Y(n_475)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_475),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_SL g503 ( 
.A(n_476),
.B(n_455),
.Y(n_503)
);

AOI22xp5_ASAP7_75t_SL g478 ( 
.A1(n_465),
.A2(n_425),
.B1(n_434),
.B2(n_438),
.Y(n_478)
);

INVx2_ASAP7_75t_L g479 ( 
.A(n_452),
.Y(n_479)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_479),
.Y(n_502)
);

NAND4xp25_ASAP7_75t_L g507 ( 
.A(n_481),
.B(n_487),
.C(n_471),
.D(n_467),
.Y(n_507)
);

AOI22xp5_ASAP7_75t_L g491 ( 
.A1(n_482),
.A2(n_466),
.B1(n_447),
.B2(n_463),
.Y(n_491)
);

XOR2xp5_ASAP7_75t_L g492 ( 
.A(n_484),
.B(n_446),
.Y(n_492)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_461),
.Y(n_485)
);

NOR2xp33_ASAP7_75t_L g504 ( 
.A(n_485),
.B(n_445),
.Y(n_504)
);

MAJIxp5_ASAP7_75t_L g486 ( 
.A(n_454),
.B(n_448),
.C(n_440),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_457),
.B(n_433),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_487),
.B(n_462),
.Y(n_498)
);

MAJIxp5_ASAP7_75t_L g488 ( 
.A(n_464),
.B(n_423),
.C(n_315),
.Y(n_488)
);

MAJIxp5_ASAP7_75t_L g497 ( 
.A(n_488),
.B(n_489),
.C(n_450),
.Y(n_497)
);

MAJIxp5_ASAP7_75t_L g489 ( 
.A(n_451),
.B(n_315),
.C(n_313),
.Y(n_489)
);

FAx1_ASAP7_75t_SL g490 ( 
.A(n_474),
.B(n_463),
.CI(n_460),
.CON(n_490),
.SN(n_490)
);

NOR2xp33_ASAP7_75t_L g509 ( 
.A(n_490),
.B(n_481),
.Y(n_509)
);

OAI22xp5_ASAP7_75t_SL g511 ( 
.A1(n_491),
.A2(n_484),
.B1(n_489),
.B2(n_475),
.Y(n_511)
);

XOR2xp5_ASAP7_75t_L g520 ( 
.A(n_492),
.B(n_493),
.Y(n_520)
);

XOR2xp5_ASAP7_75t_L g493 ( 
.A(n_477),
.B(n_442),
.Y(n_493)
);

NOR2xp67_ASAP7_75t_SL g516 ( 
.A(n_494),
.B(n_507),
.Y(n_516)
);

OAI21xp5_ASAP7_75t_SL g512 ( 
.A1(n_495),
.A2(n_475),
.B(n_479),
.Y(n_512)
);

MAJIxp5_ASAP7_75t_L g508 ( 
.A(n_497),
.B(n_505),
.C(n_483),
.Y(n_508)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_498),
.Y(n_517)
);

OAI22xp5_ASAP7_75t_SL g499 ( 
.A1(n_478),
.A2(n_443),
.B1(n_462),
.B2(n_445),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_499),
.B(n_504),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_SL g518 ( 
.A(n_503),
.B(n_506),
.Y(n_518)
);

MAJIxp5_ASAP7_75t_L g505 ( 
.A(n_483),
.B(n_444),
.C(n_452),
.Y(n_505)
);

NOR2xp33_ASAP7_75t_L g506 ( 
.A(n_468),
.B(n_352),
.Y(n_506)
);

XNOR2xp5_ASAP7_75t_L g530 ( 
.A(n_508),
.B(n_492),
.Y(n_530)
);

OAI21xp5_ASAP7_75t_L g526 ( 
.A1(n_509),
.A2(n_512),
.B(n_514),
.Y(n_526)
);

MAJIxp5_ASAP7_75t_L g510 ( 
.A(n_496),
.B(n_488),
.C(n_480),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_SL g533 ( 
.A(n_510),
.B(n_513),
.Y(n_533)
);

AOI22xp5_ASAP7_75t_L g522 ( 
.A1(n_511),
.A2(n_494),
.B1(n_499),
.B2(n_501),
.Y(n_522)
);

MAJIxp5_ASAP7_75t_L g513 ( 
.A(n_496),
.B(n_486),
.C(n_477),
.Y(n_513)
);

AOI21xp5_ASAP7_75t_L g514 ( 
.A1(n_495),
.A2(n_470),
.B(n_298),
.Y(n_514)
);

NOR2xp33_ASAP7_75t_L g515 ( 
.A(n_500),
.B(n_360),
.Y(n_515)
);

CKINVDCx16_ASAP7_75t_R g525 ( 
.A(n_515),
.Y(n_525)
);

INVx11_ASAP7_75t_L g519 ( 
.A(n_507),
.Y(n_519)
);

AOI22xp5_ASAP7_75t_L g527 ( 
.A1(n_519),
.A2(n_501),
.B1(n_498),
.B2(n_502),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g534 ( 
.A(n_522),
.B(n_523),
.Y(n_534)
);

NOR2xp33_ASAP7_75t_L g523 ( 
.A(n_521),
.B(n_503),
.Y(n_523)
);

NOR2xp33_ASAP7_75t_L g524 ( 
.A(n_521),
.B(n_506),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g538 ( 
.A(n_524),
.B(n_527),
.Y(n_538)
);

OAI22xp5_ASAP7_75t_L g528 ( 
.A1(n_519),
.A2(n_491),
.B1(n_502),
.B2(n_490),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_528),
.B(n_530),
.Y(n_540)
);

XOR2xp5_ASAP7_75t_L g529 ( 
.A(n_520),
.B(n_505),
.Y(n_529)
);

MAJIxp5_ASAP7_75t_L g542 ( 
.A(n_529),
.B(n_514),
.C(n_518),
.Y(n_542)
);

NOR2xp33_ASAP7_75t_L g531 ( 
.A(n_510),
.B(n_497),
.Y(n_531)
);

NOR2xp33_ASAP7_75t_L g535 ( 
.A(n_531),
.B(n_508),
.Y(n_535)
);

XOR2xp5_ASAP7_75t_L g532 ( 
.A(n_520),
.B(n_493),
.Y(n_532)
);

MAJIxp5_ASAP7_75t_L g537 ( 
.A(n_532),
.B(n_513),
.C(n_470),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_535),
.B(n_537),
.Y(n_543)
);

NOR3xp33_ASAP7_75t_L g536 ( 
.A(n_526),
.B(n_516),
.C(n_518),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g544 ( 
.A(n_536),
.B(n_526),
.Y(n_544)
);

MAJIxp5_ASAP7_75t_L g539 ( 
.A(n_533),
.B(n_511),
.C(n_512),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_L g546 ( 
.A(n_539),
.B(n_541),
.Y(n_546)
);

AOI22xp5_ASAP7_75t_SL g541 ( 
.A1(n_525),
.A2(n_517),
.B1(n_516),
.B2(n_490),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_L g547 ( 
.A(n_542),
.B(n_530),
.Y(n_547)
);

INVxp33_ASAP7_75t_L g553 ( 
.A(n_544),
.Y(n_553)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_538),
.Y(n_545)
);

NOR2xp33_ASAP7_75t_L g551 ( 
.A(n_545),
.B(n_548),
.Y(n_551)
);

MAJIxp5_ASAP7_75t_L g550 ( 
.A(n_547),
.B(n_540),
.C(n_529),
.Y(n_550)
);

NOR2x1_ASAP7_75t_L g548 ( 
.A(n_534),
.B(n_517),
.Y(n_548)
);

NOR2xp33_ASAP7_75t_L g549 ( 
.A(n_535),
.B(n_522),
.Y(n_549)
);

NOR2xp33_ASAP7_75t_L g552 ( 
.A(n_549),
.B(n_532),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_SL g554 ( 
.A(n_550),
.B(n_552),
.Y(n_554)
);

NOR3xp33_ASAP7_75t_L g555 ( 
.A(n_551),
.B(n_544),
.C(n_546),
.Y(n_555)
);

NAND3xp33_ASAP7_75t_L g557 ( 
.A(n_555),
.B(n_556),
.C(n_313),
.Y(n_557)
);

OAI21xp5_ASAP7_75t_SL g556 ( 
.A1(n_553),
.A2(n_543),
.B(n_548),
.Y(n_556)
);

BUFx24_ASAP7_75t_SL g559 ( 
.A(n_557),
.Y(n_559)
);

OAI22xp5_ASAP7_75t_L g558 ( 
.A1(n_554),
.A2(n_284),
.B1(n_306),
.B2(n_544),
.Y(n_558)
);

OAI21xp5_ASAP7_75t_SL g560 ( 
.A1(n_559),
.A2(n_558),
.B(n_284),
.Y(n_560)
);

INVxp67_ASAP7_75t_L g561 ( 
.A(n_560),
.Y(n_561)
);


endmodule