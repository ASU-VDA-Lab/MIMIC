module fake_jpeg_496_n_77 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_77);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_77;

wire n_10;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_40;
wire n_71;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_61;
wire n_45;
wire n_20;
wire n_18;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_11;
wire n_56;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_22;
wire n_35;
wire n_48;
wire n_46;
wire n_36;
wire n_62;
wire n_43;
wire n_32;

BUFx4f_ASAP7_75t_SL g10 ( 
.A(n_5),
.Y(n_10)
);

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_3),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_8),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_5),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_0),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_4),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_4),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_6),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

AND2x2_ASAP7_75t_L g33 ( 
.A(n_20),
.B(n_21),
.Y(n_33)
);

INVx5_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_SL g22 ( 
.A(n_13),
.B(n_0),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_SL g40 ( 
.A(n_22),
.B(n_27),
.Y(n_40)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_23),
.Y(n_31)
);

INVx8_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

INVxp67_ASAP7_75t_L g34 ( 
.A(n_24),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_19),
.B(n_9),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_25),
.B(n_26),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_19),
.B(n_12),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_11),
.B(n_18),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_11),
.B(n_9),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_28),
.B(n_29),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

MAJIxp5_ASAP7_75t_L g30 ( 
.A(n_23),
.B(n_17),
.C(n_15),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_30),
.B(n_36),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g32 ( 
.A1(n_22),
.A2(n_18),
.B1(n_17),
.B2(n_15),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_32),
.A2(n_39),
.B1(n_38),
.B2(n_35),
.Y(n_49)
);

INVxp67_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

MAJIxp5_ASAP7_75t_L g38 ( 
.A(n_29),
.B(n_14),
.C(n_13),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_SL g43 ( 
.A(n_38),
.B(n_21),
.Y(n_43)
);

OAI22xp33_ASAP7_75t_SL g39 ( 
.A1(n_28),
.A2(n_14),
.B1(n_16),
.B2(n_12),
.Y(n_39)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_31),
.Y(n_41)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_41),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_36),
.B(n_25),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_42),
.B(n_43),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g44 ( 
.A(n_40),
.B(n_16),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_44),
.B(n_46),
.Y(n_54)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_37),
.B(n_7),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_47),
.B(n_49),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_30),
.B(n_20),
.Y(n_48)
);

XNOR2xp5_ASAP7_75t_SL g56 ( 
.A(n_48),
.B(n_20),
.Y(n_56)
);

A2O1A1Ixp33_ASAP7_75t_L g50 ( 
.A1(n_33),
.A2(n_20),
.B(n_24),
.C(n_7),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_50),
.B(n_33),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_41),
.Y(n_52)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_52),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_55),
.A2(n_45),
.B1(n_49),
.B2(n_43),
.Y(n_61)
);

XNOR2xp5_ASAP7_75t_L g60 ( 
.A(n_56),
.B(n_48),
.Y(n_60)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_53),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_58),
.B(n_54),
.Y(n_64)
);

BUFx2_ASAP7_75t_L g59 ( 
.A(n_53),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_59),
.Y(n_63)
);

MAJIxp5_ASAP7_75t_L g66 ( 
.A(n_60),
.B(n_61),
.C(n_45),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_64),
.B(n_66),
.Y(n_68)
);

OAI21xp5_ASAP7_75t_L g65 ( 
.A1(n_60),
.A2(n_51),
.B(n_55),
.Y(n_65)
);

AOI21xp5_ASAP7_75t_L g67 ( 
.A1(n_65),
.A2(n_57),
.B(n_44),
.Y(n_67)
);

INVxp67_ASAP7_75t_L g71 ( 
.A(n_67),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_63),
.A2(n_62),
.B1(n_59),
.B2(n_56),
.Y(n_69)
);

AOI321xp33_ASAP7_75t_L g70 ( 
.A1(n_69),
.A2(n_50),
.A3(n_46),
.B1(n_34),
.B2(n_24),
.C(n_4),
.Y(n_70)
);

AOI21xp5_ASAP7_75t_SL g72 ( 
.A1(n_70),
.A2(n_68),
.B(n_6),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_72),
.B(n_73),
.C(n_1),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_71),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_74),
.A2(n_2),
.B1(n_3),
.B2(n_5),
.Y(n_75)
);

AOI21xp5_ASAP7_75t_L g76 ( 
.A1(n_75),
.A2(n_2),
.B(n_3),
.Y(n_76)
);

XOR2xp5_ASAP7_75t_L g77 ( 
.A(n_76),
.B(n_46),
.Y(n_77)
);


endmodule