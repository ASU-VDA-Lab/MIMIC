module fake_jpeg_13657_n_540 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_540);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_540;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_419;
wire n_378;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_260;
wire n_199;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_6),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

BUFx4f_ASAP7_75t_SL g22 ( 
.A(n_8),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_17),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_17),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

INVx11_ASAP7_75t_SL g26 ( 
.A(n_2),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_17),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_15),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_4),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_18),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_1),
.Y(n_33)
);

BUFx10_ASAP7_75t_L g34 ( 
.A(n_17),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_3),
.B(n_18),
.Y(n_36)
);

INVx11_ASAP7_75t_L g37 ( 
.A(n_11),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_1),
.Y(n_38)
);

BUFx10_ASAP7_75t_L g39 ( 
.A(n_10),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_2),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_6),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_9),
.Y(n_42)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_3),
.Y(n_43)
);

INVx11_ASAP7_75t_SL g44 ( 
.A(n_4),
.Y(n_44)
);

BUFx5_ASAP7_75t_L g45 ( 
.A(n_16),
.Y(n_45)
);

BUFx10_ASAP7_75t_L g46 ( 
.A(n_12),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_3),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_14),
.Y(n_48)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_10),
.Y(n_49)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_4),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_7),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_12),
.Y(n_52)
);

AOI21xp33_ASAP7_75t_L g53 ( 
.A1(n_36),
.A2(n_18),
.B(n_1),
.Y(n_53)
);

AOI21xp33_ASAP7_75t_L g107 ( 
.A1(n_53),
.A2(n_52),
.B(n_20),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_36),
.B(n_0),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_54),
.B(n_60),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_22),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_55),
.Y(n_133)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_21),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g108 ( 
.A(n_56),
.Y(n_108)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_50),
.Y(n_57)
);

INVx5_ASAP7_75t_L g118 ( 
.A(n_57),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_22),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_58),
.Y(n_140)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_50),
.Y(n_59)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_59),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_30),
.B(n_0),
.Y(n_60)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_21),
.Y(n_61)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_61),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_22),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_62),
.Y(n_143)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_50),
.Y(n_63)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_63),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_22),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_64),
.Y(n_148)
);

INVx3_ASAP7_75t_SL g65 ( 
.A(n_34),
.Y(n_65)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_65),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_22),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_66),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_30),
.B(n_0),
.Y(n_67)
);

AND2x2_ASAP7_75t_L g131 ( 
.A(n_67),
.B(n_91),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_19),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_68),
.Y(n_153)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_25),
.Y(n_69)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_69),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_19),
.Y(n_70)
);

INVx6_ASAP7_75t_L g112 ( 
.A(n_70),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_19),
.Y(n_71)
);

INVx6_ASAP7_75t_L g114 ( 
.A(n_71),
.Y(n_114)
);

BUFx12f_ASAP7_75t_L g72 ( 
.A(n_21),
.Y(n_72)
);

INVx5_ASAP7_75t_L g163 ( 
.A(n_72),
.Y(n_163)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_25),
.Y(n_73)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_73),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_19),
.Y(n_74)
);

INVx6_ASAP7_75t_L g135 ( 
.A(n_74),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_32),
.Y(n_75)
);

INVx6_ASAP7_75t_L g136 ( 
.A(n_75),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_32),
.Y(n_76)
);

INVx6_ASAP7_75t_L g151 ( 
.A(n_76),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_32),
.Y(n_77)
);

INVx6_ASAP7_75t_L g155 ( 
.A(n_77),
.Y(n_155)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_25),
.Y(n_78)
);

INVx3_ASAP7_75t_L g144 ( 
.A(n_78),
.Y(n_144)
);

INVx3_ASAP7_75t_SL g79 ( 
.A(n_34),
.Y(n_79)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_79),
.Y(n_122)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_45),
.Y(n_80)
);

INVx4_ASAP7_75t_L g116 ( 
.A(n_80),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_32),
.Y(n_81)
);

INVx4_ASAP7_75t_L g120 ( 
.A(n_81),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_35),
.Y(n_82)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_82),
.Y(n_127)
);

BUFx5_ASAP7_75t_L g83 ( 
.A(n_45),
.Y(n_83)
);

INVx4_ASAP7_75t_L g157 ( 
.A(n_83),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_35),
.Y(n_84)
);

INVx3_ASAP7_75t_L g156 ( 
.A(n_84),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_35),
.Y(n_85)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_85),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_35),
.Y(n_86)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_86),
.Y(n_129)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_41),
.Y(n_87)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_87),
.Y(n_134)
);

INVx11_ASAP7_75t_L g88 ( 
.A(n_34),
.Y(n_88)
);

HB1xp67_ASAP7_75t_L g109 ( 
.A(n_88),
.Y(n_109)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_23),
.Y(n_89)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_89),
.Y(n_110)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_41),
.Y(n_90)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_90),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_52),
.B(n_0),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_40),
.Y(n_92)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_92),
.Y(n_146)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_41),
.Y(n_93)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_93),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_40),
.Y(n_94)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_94),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_40),
.Y(n_95)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_95),
.Y(n_121)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_23),
.Y(n_96)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_96),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_40),
.Y(n_97)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_97),
.Y(n_141)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_31),
.Y(n_98)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_98),
.Y(n_142)
);

INVx6_ASAP7_75t_L g99 ( 
.A(n_47),
.Y(n_99)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_99),
.Y(n_152)
);

BUFx12f_ASAP7_75t_L g100 ( 
.A(n_45),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_100),
.B(n_102),
.Y(n_119)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_49),
.Y(n_101)
);

NAND2xp33_ASAP7_75t_SL g125 ( 
.A(n_101),
.B(n_104),
.Y(n_125)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_31),
.Y(n_102)
);

INVx5_ASAP7_75t_L g103 ( 
.A(n_49),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_103),
.B(n_56),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_47),
.Y(n_104)
);

AND2x2_ASAP7_75t_L g171 ( 
.A(n_107),
.B(n_147),
.Y(n_171)
);

CKINVDCx14_ASAP7_75t_R g199 ( 
.A(n_124),
.Y(n_199)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_65),
.A2(n_49),
.B1(n_46),
.B2(n_39),
.Y(n_126)
);

OAI22x1_ASAP7_75t_L g205 ( 
.A1(n_126),
.A2(n_160),
.B1(n_46),
.B2(n_39),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_60),
.B(n_24),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_128),
.B(n_130),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_67),
.B(n_91),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_79),
.B(n_48),
.C(n_38),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_145),
.B(n_46),
.C(n_39),
.Y(n_213)
);

AND2x2_ASAP7_75t_SL g147 ( 
.A(n_55),
.B(n_34),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_58),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_149),
.B(n_64),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_72),
.B(n_24),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_154),
.B(n_162),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_68),
.A2(n_43),
.B1(n_51),
.B2(n_47),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_158),
.A2(n_161),
.B1(n_51),
.B2(n_97),
.Y(n_204)
);

AOI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_62),
.A2(n_34),
.B1(n_46),
.B2(n_39),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_L g161 ( 
.A1(n_70),
.A2(n_43),
.B1(n_47),
.B2(n_51),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_100),
.B(n_20),
.Y(n_162)
);

INVx11_ASAP7_75t_L g164 ( 
.A(n_157),
.Y(n_164)
);

BUFx2_ASAP7_75t_L g264 ( 
.A(n_164),
.Y(n_264)
);

INVx3_ASAP7_75t_L g165 ( 
.A(n_133),
.Y(n_165)
);

INVx1_ASAP7_75t_SL g225 ( 
.A(n_165),
.Y(n_225)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_110),
.Y(n_166)
);

INVx1_ASAP7_75t_SL g252 ( 
.A(n_166),
.Y(n_252)
);

INVx3_ASAP7_75t_L g167 ( 
.A(n_133),
.Y(n_167)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_167),
.Y(n_234)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_152),
.Y(n_168)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_168),
.Y(n_236)
);

INVx4_ASAP7_75t_L g169 ( 
.A(n_140),
.Y(n_169)
);

INVx5_ASAP7_75t_L g250 ( 
.A(n_169),
.Y(n_250)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_123),
.Y(n_172)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_172),
.Y(n_239)
);

CKINVDCx16_ASAP7_75t_R g173 ( 
.A(n_119),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_173),
.B(n_179),
.Y(n_223)
);

INVx4_ASAP7_75t_L g174 ( 
.A(n_140),
.Y(n_174)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_174),
.Y(n_241)
);

INVx3_ASAP7_75t_L g175 ( 
.A(n_143),
.Y(n_175)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_175),
.Y(n_248)
);

INVx3_ASAP7_75t_L g176 ( 
.A(n_143),
.Y(n_176)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_176),
.Y(n_253)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_129),
.Y(n_177)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_177),
.Y(n_224)
);

BUFx3_ASAP7_75t_L g178 ( 
.A(n_108),
.Y(n_178)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_178),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_109),
.Y(n_179)
);

INVx6_ASAP7_75t_L g180 ( 
.A(n_153),
.Y(n_180)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_180),
.Y(n_231)
);

INVx8_ASAP7_75t_L g181 ( 
.A(n_148),
.Y(n_181)
);

INVxp67_ASAP7_75t_L g260 ( 
.A(n_181),
.Y(n_260)
);

AOI22xp33_ASAP7_75t_SL g182 ( 
.A1(n_157),
.A2(n_37),
.B1(n_38),
.B2(n_48),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_SL g244 ( 
.A1(n_182),
.A2(n_205),
.B1(n_221),
.B2(n_135),
.Y(n_244)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_146),
.Y(n_183)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_183),
.Y(n_232)
);

CKINVDCx16_ASAP7_75t_R g240 ( 
.A(n_184),
.Y(n_240)
);

INVx5_ASAP7_75t_L g185 ( 
.A(n_148),
.Y(n_185)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_185),
.Y(n_233)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_137),
.Y(n_186)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_186),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_106),
.B(n_42),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_187),
.B(n_192),
.Y(n_242)
);

BUFx2_ASAP7_75t_L g188 ( 
.A(n_150),
.Y(n_188)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_188),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_131),
.B(n_142),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_189),
.B(n_190),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_131),
.B(n_42),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_115),
.Y(n_191)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_191),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_109),
.Y(n_192)
);

HB1xp67_ASAP7_75t_L g193 ( 
.A(n_122),
.Y(n_193)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_193),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_134),
.B(n_33),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_194),
.B(n_195),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_138),
.B(n_159),
.Y(n_195)
);

INVx6_ASAP7_75t_SL g196 ( 
.A(n_118),
.Y(n_196)
);

CKINVDCx14_ASAP7_75t_R g238 ( 
.A(n_196),
.Y(n_238)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_111),
.Y(n_197)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_197),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_147),
.A2(n_43),
.B1(n_39),
.B2(n_34),
.Y(n_198)
);

AOI21xp5_ASAP7_75t_L g254 ( 
.A1(n_198),
.A2(n_215),
.B(n_222),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_161),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_200),
.B(n_203),
.Y(n_255)
);

INVx3_ASAP7_75t_L g201 ( 
.A(n_150),
.Y(n_201)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_201),
.Y(n_268)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_121),
.Y(n_202)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_202),
.Y(n_269)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_141),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_204),
.A2(n_155),
.B1(n_151),
.B2(n_136),
.Y(n_230)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_132),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_206),
.B(n_207),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_120),
.Y(n_207)
);

NAND2x1_ASAP7_75t_SL g208 ( 
.A(n_113),
.B(n_66),
.Y(n_208)
);

OR2x6_ASAP7_75t_L g235 ( 
.A(n_208),
.B(n_37),
.Y(n_235)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_156),
.Y(n_209)
);

AND2x2_ASAP7_75t_L g245 ( 
.A(n_209),
.B(n_210),
.Y(n_245)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_139),
.Y(n_210)
);

CKINVDCx14_ASAP7_75t_R g211 ( 
.A(n_163),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_211),
.B(n_214),
.Y(n_261)
);

AND2x2_ASAP7_75t_L g265 ( 
.A(n_213),
.B(n_219),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_144),
.B(n_33),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_116),
.A2(n_46),
.B1(n_39),
.B2(n_44),
.Y(n_215)
);

BUFx3_ASAP7_75t_L g216 ( 
.A(n_108),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_216),
.B(n_218),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_125),
.B(n_29),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_217),
.B(n_28),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_120),
.Y(n_218)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_127),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_105),
.Y(n_220)
);

INVxp33_ASAP7_75t_L g256 ( 
.A(n_220),
.Y(n_256)
);

BUFx6f_ASAP7_75t_L g221 ( 
.A(n_153),
.Y(n_221)
);

AOI21xp5_ASAP7_75t_L g222 ( 
.A1(n_126),
.A2(n_46),
.B(n_37),
.Y(n_222)
);

OAI22xp33_ASAP7_75t_SL g228 ( 
.A1(n_215),
.A2(n_160),
.B1(n_127),
.B2(n_117),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_SL g319 ( 
.A1(n_228),
.A2(n_229),
.B1(n_235),
.B2(n_260),
.Y(n_319)
);

OAI22xp33_ASAP7_75t_SL g229 ( 
.A1(n_217),
.A2(n_116),
.B1(n_81),
.B2(n_104),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_L g308 ( 
.A1(n_230),
.A2(n_237),
.B1(n_270),
.B2(n_272),
.Y(n_308)
);

CKINVDCx14_ASAP7_75t_R g302 ( 
.A(n_235),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_204),
.A2(n_155),
.B1(n_151),
.B2(n_136),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_171),
.B(n_135),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_243),
.B(n_208),
.C(n_209),
.Y(n_277)
);

INVxp67_ASAP7_75t_L g301 ( 
.A(n_244),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_SL g310 ( 
.A(n_246),
.B(n_27),
.Y(n_310)
);

AOI22xp33_ASAP7_75t_SL g249 ( 
.A1(n_205),
.A2(n_114),
.B1(n_112),
.B2(n_28),
.Y(n_249)
);

INVxp67_ASAP7_75t_L g313 ( 
.A(n_249),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_189),
.B(n_213),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_267),
.B(n_273),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_171),
.A2(n_114),
.B1(n_112),
.B2(n_95),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_171),
.A2(n_26),
.B1(n_44),
.B2(n_51),
.Y(n_271)
);

OAI21xp5_ASAP7_75t_L g288 ( 
.A1(n_271),
.A2(n_27),
.B(n_178),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_190),
.A2(n_94),
.B1(n_92),
.B2(n_86),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_212),
.B(n_29),
.Y(n_273)
);

AND2x2_ASAP7_75t_L g274 ( 
.A(n_265),
.B(n_255),
.Y(n_274)
);

INVxp67_ASAP7_75t_L g361 ( 
.A(n_274),
.Y(n_361)
);

OAI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_254),
.A2(n_222),
.B1(n_198),
.B2(n_170),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_275),
.A2(n_287),
.B1(n_288),
.B2(n_311),
.Y(n_321)
);

AOI22xp33_ASAP7_75t_SL g276 ( 
.A1(n_225),
.A2(n_196),
.B1(n_164),
.B2(n_188),
.Y(n_276)
);

OAI21xp5_ASAP7_75t_L g324 ( 
.A1(n_276),
.A2(n_291),
.B(n_316),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_277),
.B(n_293),
.C(n_297),
.Y(n_345)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_243),
.A2(n_199),
.B1(n_210),
.B2(n_177),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_SL g323 ( 
.A1(n_279),
.A2(n_285),
.B1(n_289),
.B2(n_305),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_265),
.B(n_202),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_280),
.B(n_290),
.Y(n_328)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_269),
.Y(n_281)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_281),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_247),
.B(n_168),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_SL g347 ( 
.A(n_282),
.B(n_310),
.Y(n_347)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_245),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_283),
.B(n_286),
.Y(n_322)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_269),
.Y(n_284)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_284),
.Y(n_335)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_265),
.A2(n_172),
.B1(n_183),
.B2(n_180),
.Y(n_285)
);

CKINVDCx16_ASAP7_75t_R g286 ( 
.A(n_245),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_254),
.A2(n_75),
.B1(n_85),
.B2(n_84),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_267),
.A2(n_246),
.B1(n_240),
.B2(n_230),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_226),
.B(n_219),
.Y(n_290)
);

AOI22xp33_ASAP7_75t_SL g291 ( 
.A1(n_225),
.A2(n_216),
.B1(n_181),
.B2(n_201),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_259),
.Y(n_292)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_292),
.Y(n_338)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_226),
.B(n_242),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_223),
.B(n_174),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_294),
.B(n_298),
.Y(n_329)
);

BUFx3_ASAP7_75t_L g295 ( 
.A(n_227),
.Y(n_295)
);

INVx5_ASAP7_75t_L g337 ( 
.A(n_295),
.Y(n_337)
);

AND2x2_ASAP7_75t_L g296 ( 
.A(n_270),
.B(n_165),
.Y(n_296)
);

OAI21xp5_ASAP7_75t_SL g350 ( 
.A1(n_296),
.A2(n_319),
.B(n_241),
.Y(n_350)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_251),
.B(n_167),
.C(n_176),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_262),
.B(n_169),
.Y(n_298)
);

INVxp67_ASAP7_75t_SL g299 ( 
.A(n_227),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_299),
.B(n_303),
.Y(n_325)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_259),
.Y(n_300)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_300),
.Y(n_342)
);

NAND3xp33_ASAP7_75t_L g303 ( 
.A(n_261),
.B(n_2),
.C(n_3),
.Y(n_303)
);

BUFx8_ASAP7_75t_L g304 ( 
.A(n_238),
.Y(n_304)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_304),
.Y(n_343)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_237),
.A2(n_175),
.B1(n_71),
.B2(n_76),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_273),
.B(n_185),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_306),
.B(n_260),
.Y(n_331)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_268),
.Y(n_307)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_307),
.Y(n_353)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_224),
.Y(n_309)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_309),
.Y(n_357)
);

OAI22xp33_ASAP7_75t_SL g311 ( 
.A1(n_235),
.A2(n_221),
.B1(n_82),
.B2(n_77),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_L g312 ( 
.A1(n_235),
.A2(n_74),
.B1(n_26),
.B2(n_5),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g334 ( 
.A1(n_312),
.A2(n_231),
.B1(n_233),
.B2(n_250),
.Y(n_334)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_271),
.B(n_258),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g348 ( 
.A(n_314),
.B(n_232),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_SL g315 ( 
.A(n_252),
.B(n_251),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_SL g362 ( 
.A(n_315),
.B(n_239),
.Y(n_362)
);

AOI22xp33_ASAP7_75t_SL g316 ( 
.A1(n_268),
.A2(n_233),
.B1(n_235),
.B2(n_248),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_252),
.B(n_2),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_317),
.B(n_318),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_256),
.B(n_266),
.Y(n_318)
);

AOI22xp33_ASAP7_75t_L g320 ( 
.A1(n_235),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_320),
.Y(n_326)
);

OAI21xp5_ASAP7_75t_L g327 ( 
.A1(n_302),
.A2(n_266),
.B(n_245),
.Y(n_327)
);

OAI21xp5_ASAP7_75t_L g374 ( 
.A1(n_327),
.A2(n_332),
.B(n_284),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_331),
.B(n_336),
.Y(n_363)
);

OAI21xp5_ASAP7_75t_L g332 ( 
.A1(n_274),
.A2(n_263),
.B(n_236),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_L g373 ( 
.A1(n_334),
.A2(n_349),
.B1(n_305),
.B2(n_296),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_SL g336 ( 
.A(n_293),
.B(n_263),
.Y(n_336)
);

AOI21xp5_ASAP7_75t_L g339 ( 
.A1(n_313),
.A2(n_264),
.B(n_257),
.Y(n_339)
);

AOI21xp5_ASAP7_75t_L g394 ( 
.A1(n_339),
.A2(n_354),
.B(n_356),
.Y(n_394)
);

OAI22xp5_ASAP7_75t_SL g340 ( 
.A1(n_319),
.A2(n_272),
.B1(n_231),
.B2(n_257),
.Y(n_340)
);

AOI22xp5_ASAP7_75t_L g379 ( 
.A1(n_340),
.A2(n_323),
.B1(n_326),
.B2(n_359),
.Y(n_379)
);

CKINVDCx20_ASAP7_75t_R g341 ( 
.A(n_298),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g386 ( 
.A(n_341),
.B(n_344),
.Y(n_386)
);

CKINVDCx20_ASAP7_75t_R g344 ( 
.A(n_294),
.Y(n_344)
);

OAI32xp33_ASAP7_75t_L g346 ( 
.A1(n_278),
.A2(n_224),
.A3(n_232),
.B1(n_253),
.B2(n_248),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_346),
.B(n_355),
.Y(n_375)
);

XNOR2xp5_ASAP7_75t_SL g398 ( 
.A(n_348),
.B(n_13),
.Y(n_398)
);

AOI22xp5_ASAP7_75t_L g349 ( 
.A1(n_275),
.A2(n_308),
.B1(n_313),
.B2(n_287),
.Y(n_349)
);

OR2x2_ASAP7_75t_L g381 ( 
.A(n_350),
.B(n_234),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_289),
.B(n_306),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_SL g378 ( 
.A(n_351),
.B(n_352),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_L g352 ( 
.A(n_310),
.B(n_236),
.Y(n_352)
);

AOI21xp5_ASAP7_75t_L g354 ( 
.A1(n_301),
.A2(n_264),
.B(n_250),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_L g355 ( 
.A(n_278),
.B(n_239),
.Y(n_355)
);

AOI21xp5_ASAP7_75t_L g356 ( 
.A1(n_301),
.A2(n_264),
.B(n_253),
.Y(n_356)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_292),
.Y(n_358)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_358),
.Y(n_369)
);

AO22x1_ASAP7_75t_SL g359 ( 
.A1(n_308),
.A2(n_296),
.B1(n_312),
.B2(n_279),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_359),
.B(n_350),
.Y(n_389)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_300),
.Y(n_360)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_360),
.Y(n_382)
);

NOR2xp33_ASAP7_75t_L g391 ( 
.A(n_362),
.B(n_12),
.Y(n_391)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_345),
.B(n_280),
.C(n_274),
.Y(n_364)
);

MAJIxp5_ASAP7_75t_L g413 ( 
.A(n_364),
.B(n_370),
.C(n_371),
.Y(n_413)
);

AOI22xp5_ASAP7_75t_SL g365 ( 
.A1(n_361),
.A2(n_344),
.B1(n_341),
.B2(n_340),
.Y(n_365)
);

OAI21xp5_ASAP7_75t_SL g415 ( 
.A1(n_365),
.A2(n_381),
.B(n_390),
.Y(n_415)
);

OAI22xp5_ASAP7_75t_SL g366 ( 
.A1(n_349),
.A2(n_290),
.B1(n_277),
.B2(n_283),
.Y(n_366)
);

AOI22xp5_ASAP7_75t_L g427 ( 
.A1(n_366),
.A2(n_373),
.B1(n_380),
.B2(n_383),
.Y(n_427)
);

INVx3_ASAP7_75t_L g367 ( 
.A(n_337),
.Y(n_367)
);

BUFx2_ASAP7_75t_L g420 ( 
.A(n_367),
.Y(n_420)
);

INVx2_ASAP7_75t_L g368 ( 
.A(n_330),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_368),
.B(n_376),
.Y(n_417)
);

MAJIxp5_ASAP7_75t_L g370 ( 
.A(n_345),
.B(n_285),
.C(n_314),
.Y(n_370)
);

MAJIxp5_ASAP7_75t_L g371 ( 
.A(n_336),
.B(n_297),
.C(n_309),
.Y(n_371)
);

XNOR2xp5_ASAP7_75t_L g372 ( 
.A(n_348),
.B(n_288),
.Y(n_372)
);

MAJIxp5_ASAP7_75t_L g419 ( 
.A(n_372),
.B(n_384),
.C(n_398),
.Y(n_419)
);

AO21x1_ASAP7_75t_L g410 ( 
.A1(n_374),
.A2(n_377),
.B(n_388),
.Y(n_410)
);

CKINVDCx20_ASAP7_75t_R g376 ( 
.A(n_331),
.Y(n_376)
);

OAI21xp5_ASAP7_75t_L g377 ( 
.A1(n_322),
.A2(n_281),
.B(n_307),
.Y(n_377)
);

OAI22xp5_ASAP7_75t_L g423 ( 
.A1(n_379),
.A2(n_387),
.B1(n_389),
.B2(n_397),
.Y(n_423)
);

OAI22xp5_ASAP7_75t_L g380 ( 
.A1(n_321),
.A2(n_295),
.B1(n_234),
.B2(n_304),
.Y(n_380)
);

OAI22xp5_ASAP7_75t_SL g383 ( 
.A1(n_321),
.A2(n_241),
.B1(n_304),
.B2(n_8),
.Y(n_383)
);

MAJIxp5_ASAP7_75t_L g384 ( 
.A(n_322),
.B(n_304),
.C(n_7),
.Y(n_384)
);

OAI22xp5_ASAP7_75t_SL g385 ( 
.A1(n_351),
.A2(n_5),
.B1(n_7),
.B2(n_8),
.Y(n_385)
);

AOI22xp5_ASAP7_75t_L g428 ( 
.A1(n_385),
.A2(n_392),
.B1(n_342),
.B2(n_357),
.Y(n_428)
);

AOI22xp5_ASAP7_75t_L g387 ( 
.A1(n_323),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_387)
);

OAI21xp5_ASAP7_75t_L g388 ( 
.A1(n_327),
.A2(n_9),
.B(n_10),
.Y(n_388)
);

A2O1A1O1Ixp25_ASAP7_75t_L g390 ( 
.A1(n_328),
.A2(n_9),
.B(n_10),
.C(n_11),
.D(n_12),
.Y(n_390)
);

CKINVDCx14_ASAP7_75t_R g409 ( 
.A(n_391),
.Y(n_409)
);

OAI22xp5_ASAP7_75t_SL g392 ( 
.A1(n_359),
.A2(n_328),
.B1(n_355),
.B2(n_326),
.Y(n_392)
);

CKINVDCx20_ASAP7_75t_R g393 ( 
.A(n_329),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_393),
.B(n_395),
.Y(n_411)
);

CKINVDCx20_ASAP7_75t_R g395 ( 
.A(n_329),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_338),
.Y(n_396)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_396),
.Y(n_406)
);

AOI22xp5_ASAP7_75t_SL g397 ( 
.A1(n_359),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_397)
);

XNOR2xp5_ASAP7_75t_L g401 ( 
.A(n_398),
.B(n_333),
.Y(n_401)
);

OAI22xp5_ASAP7_75t_SL g399 ( 
.A1(n_379),
.A2(n_339),
.B1(n_356),
.B2(n_354),
.Y(n_399)
);

AOI22xp5_ASAP7_75t_SL g431 ( 
.A1(n_399),
.A2(n_402),
.B1(n_405),
.B2(n_422),
.Y(n_431)
);

AOI21xp5_ASAP7_75t_L g400 ( 
.A1(n_394),
.A2(n_324),
.B(n_332),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_400),
.B(n_416),
.Y(n_432)
);

XNOR2xp5_ASAP7_75t_L g443 ( 
.A(n_401),
.B(n_419),
.Y(n_443)
);

OAI22xp5_ASAP7_75t_SL g402 ( 
.A1(n_365),
.A2(n_389),
.B1(n_375),
.B2(n_397),
.Y(n_402)
);

XOR2xp5_ASAP7_75t_L g403 ( 
.A(n_364),
.B(n_346),
.Y(n_403)
);

XOR2xp5_ASAP7_75t_L g437 ( 
.A(n_403),
.B(n_404),
.Y(n_437)
);

XNOR2xp5_ASAP7_75t_L g404 ( 
.A(n_372),
.B(n_362),
.Y(n_404)
);

OAI22xp5_ASAP7_75t_SL g405 ( 
.A1(n_375),
.A2(n_334),
.B1(n_324),
.B2(n_347),
.Y(n_405)
);

CKINVDCx16_ASAP7_75t_R g407 ( 
.A(n_377),
.Y(n_407)
);

CKINVDCx14_ASAP7_75t_R g441 ( 
.A(n_407),
.Y(n_441)
);

BUFx3_ASAP7_75t_L g408 ( 
.A(n_367),
.Y(n_408)
);

BUFx6f_ASAP7_75t_L g454 ( 
.A(n_408),
.Y(n_454)
);

XNOR2xp5_ASAP7_75t_L g412 ( 
.A(n_370),
.B(n_352),
.Y(n_412)
);

MAJIxp5_ASAP7_75t_L g433 ( 
.A(n_412),
.B(n_418),
.C(n_426),
.Y(n_433)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_368),
.Y(n_414)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_414),
.Y(n_430)
);

CKINVDCx14_ASAP7_75t_R g416 ( 
.A(n_378),
.Y(n_416)
);

XNOR2xp5_ASAP7_75t_L g418 ( 
.A(n_371),
.B(n_333),
.Y(n_418)
);

FAx1_ASAP7_75t_SL g421 ( 
.A(n_363),
.B(n_347),
.CI(n_325),
.CON(n_421),
.SN(n_421)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_421),
.B(n_385),
.Y(n_445)
);

OAI22xp5_ASAP7_75t_SL g422 ( 
.A1(n_393),
.A2(n_360),
.B1(n_358),
.B2(n_338),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_SL g424 ( 
.A(n_386),
.B(n_325),
.Y(n_424)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_424),
.Y(n_434)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_369),
.Y(n_425)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_425),
.Y(n_438)
);

MAJIxp5_ASAP7_75t_L g426 ( 
.A(n_366),
.B(n_353),
.C(n_342),
.Y(n_426)
);

OAI22xp5_ASAP7_75t_SL g435 ( 
.A1(n_428),
.A2(n_381),
.B1(n_376),
.B2(n_387),
.Y(n_435)
);

NOR2xp33_ASAP7_75t_SL g429 ( 
.A(n_395),
.B(n_363),
.Y(n_429)
);

CKINVDCx20_ASAP7_75t_R g436 ( 
.A(n_429),
.Y(n_436)
);

AOI22xp5_ASAP7_75t_L g477 ( 
.A1(n_435),
.A2(n_442),
.B1(n_453),
.B2(n_15),
.Y(n_477)
);

AOI22xp5_ASAP7_75t_SL g439 ( 
.A1(n_405),
.A2(n_392),
.B1(n_380),
.B2(n_383),
.Y(n_439)
);

OAI22xp5_ASAP7_75t_SL g459 ( 
.A1(n_439),
.A2(n_410),
.B1(n_400),
.B2(n_423),
.Y(n_459)
);

MAJIxp5_ASAP7_75t_L g440 ( 
.A(n_413),
.B(n_374),
.C(n_394),
.Y(n_440)
);

MAJIxp5_ASAP7_75t_L g462 ( 
.A(n_440),
.B(n_450),
.C(n_455),
.Y(n_462)
);

OAI22xp5_ASAP7_75t_SL g442 ( 
.A1(n_427),
.A2(n_396),
.B1(n_382),
.B2(n_369),
.Y(n_442)
);

CKINVDCx20_ASAP7_75t_R g444 ( 
.A(n_411),
.Y(n_444)
);

CKINVDCx20_ASAP7_75t_R g473 ( 
.A(n_444),
.Y(n_473)
);

OAI22xp5_ASAP7_75t_L g457 ( 
.A1(n_445),
.A2(n_451),
.B1(n_410),
.B2(n_426),
.Y(n_457)
);

XNOR2xp5_ASAP7_75t_L g446 ( 
.A(n_412),
.B(n_384),
.Y(n_446)
);

XNOR2xp5_ASAP7_75t_L g458 ( 
.A(n_446),
.B(n_452),
.Y(n_458)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_422),
.Y(n_447)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_447),
.Y(n_456)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_411),
.Y(n_448)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_448),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_417),
.B(n_382),
.Y(n_449)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_449),
.Y(n_463)
);

MAJIxp5_ASAP7_75t_L g450 ( 
.A(n_413),
.B(n_353),
.C(n_357),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_406),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_428),
.B(n_335),
.Y(n_452)
);

OAI22xp5_ASAP7_75t_SL g453 ( 
.A1(n_427),
.A2(n_388),
.B1(n_335),
.B2(n_330),
.Y(n_453)
);

MAJIxp5_ASAP7_75t_L g455 ( 
.A(n_403),
.B(n_343),
.C(n_337),
.Y(n_455)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_457),
.Y(n_491)
);

HB1xp67_ASAP7_75t_L g488 ( 
.A(n_459),
.Y(n_488)
);

XOR2xp5_ASAP7_75t_L g461 ( 
.A(n_440),
.B(n_418),
.Y(n_461)
);

XOR2xp5_ASAP7_75t_L g485 ( 
.A(n_461),
.B(n_467),
.Y(n_485)
);

INVx11_ASAP7_75t_L g464 ( 
.A(n_441),
.Y(n_464)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_464),
.Y(n_493)
);

MAJIxp5_ASAP7_75t_L g465 ( 
.A(n_450),
.B(n_404),
.C(n_419),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_SL g492 ( 
.A(n_465),
.B(n_468),
.Y(n_492)
);

OAI22xp5_ASAP7_75t_L g466 ( 
.A1(n_436),
.A2(n_409),
.B1(n_421),
.B2(n_415),
.Y(n_466)
);

HB1xp67_ASAP7_75t_L g490 ( 
.A(n_466),
.Y(n_490)
);

FAx1_ASAP7_75t_L g467 ( 
.A(n_431),
.B(n_402),
.CI(n_399),
.CON(n_467),
.SN(n_467)
);

MAJIxp5_ASAP7_75t_L g468 ( 
.A(n_433),
.B(n_401),
.C(n_415),
.Y(n_468)
);

XNOR2xp5_ASAP7_75t_L g469 ( 
.A(n_433),
.B(n_343),
.Y(n_469)
);

XNOR2xp5_ASAP7_75t_L g483 ( 
.A(n_469),
.B(n_471),
.Y(n_483)
);

MAJIxp5_ASAP7_75t_L g470 ( 
.A(n_437),
.B(n_420),
.C(n_421),
.Y(n_470)
);

MAJIxp5_ASAP7_75t_L g478 ( 
.A(n_470),
.B(n_443),
.C(n_446),
.Y(n_478)
);

XNOR2xp5_ASAP7_75t_L g471 ( 
.A(n_443),
.B(n_390),
.Y(n_471)
);

OAI21xp5_ASAP7_75t_SL g472 ( 
.A1(n_432),
.A2(n_420),
.B(n_408),
.Y(n_472)
);

AOI21xp5_ASAP7_75t_L g482 ( 
.A1(n_472),
.A2(n_430),
.B(n_451),
.Y(n_482)
);

XOR2xp5_ASAP7_75t_L g474 ( 
.A(n_455),
.B(n_13),
.Y(n_474)
);

XNOR2xp5_ASAP7_75t_L g484 ( 
.A(n_474),
.B(n_476),
.Y(n_484)
);

FAx1_ASAP7_75t_SL g475 ( 
.A(n_445),
.B(n_13),
.CI(n_14),
.CON(n_475),
.SN(n_475)
);

OAI22xp5_ASAP7_75t_SL g479 ( 
.A1(n_475),
.A2(n_477),
.B1(n_439),
.B2(n_431),
.Y(n_479)
);

XOR2xp5_ASAP7_75t_L g476 ( 
.A(n_437),
.B(n_14),
.Y(n_476)
);

NOR2xp67_ASAP7_75t_SL g506 ( 
.A(n_478),
.B(n_465),
.Y(n_506)
);

AOI22xp5_ASAP7_75t_L g504 ( 
.A1(n_479),
.A2(n_481),
.B1(n_494),
.B2(n_459),
.Y(n_504)
);

MAJIxp5_ASAP7_75t_L g480 ( 
.A(n_462),
.B(n_447),
.C(n_432),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_SL g501 ( 
.A(n_480),
.B(n_486),
.Y(n_501)
);

OAI22xp5_ASAP7_75t_SL g481 ( 
.A1(n_477),
.A2(n_448),
.B1(n_452),
.B2(n_449),
.Y(n_481)
);

AOI21xp5_ASAP7_75t_L g495 ( 
.A1(n_482),
.A2(n_487),
.B(n_489),
.Y(n_495)
);

MAJIxp5_ASAP7_75t_L g486 ( 
.A(n_462),
.B(n_442),
.C(n_453),
.Y(n_486)
);

AOI21xp5_ASAP7_75t_L g487 ( 
.A1(n_470),
.A2(n_472),
.B(n_469),
.Y(n_487)
);

AOI21xp5_ASAP7_75t_L g489 ( 
.A1(n_464),
.A2(n_434),
.B(n_438),
.Y(n_489)
);

OAI22xp5_ASAP7_75t_SL g494 ( 
.A1(n_473),
.A2(n_435),
.B1(n_454),
.B2(n_15),
.Y(n_494)
);

NOR2xp33_ASAP7_75t_L g496 ( 
.A(n_480),
.B(n_454),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_496),
.B(n_499),
.Y(n_510)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_494),
.Y(n_497)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_497),
.Y(n_517)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_493),
.Y(n_498)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_498),
.Y(n_519)
);

XNOR2xp5_ASAP7_75t_L g499 ( 
.A(n_478),
.B(n_458),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_481),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_500),
.B(n_502),
.Y(n_512)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_491),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_490),
.Y(n_503)
);

NOR2xp33_ASAP7_75t_L g511 ( 
.A(n_503),
.B(n_475),
.Y(n_511)
);

OAI22xp5_ASAP7_75t_SL g515 ( 
.A1(n_504),
.A2(n_467),
.B1(n_485),
.B2(n_471),
.Y(n_515)
);

OAI21xp5_ASAP7_75t_SL g505 ( 
.A1(n_488),
.A2(n_456),
.B(n_460),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_SL g516 ( 
.A(n_505),
.B(n_506),
.Y(n_516)
);

NOR2xp33_ASAP7_75t_L g507 ( 
.A(n_486),
.B(n_458),
.Y(n_507)
);

NOR2xp33_ASAP7_75t_SL g518 ( 
.A(n_507),
.B(n_509),
.Y(n_518)
);

OAI22xp5_ASAP7_75t_SL g508 ( 
.A1(n_479),
.A2(n_463),
.B1(n_467),
.B2(n_468),
.Y(n_508)
);

XNOR2xp5_ASAP7_75t_L g514 ( 
.A(n_508),
.B(n_485),
.Y(n_514)
);

NOR2xp33_ASAP7_75t_L g509 ( 
.A(n_492),
.B(n_475),
.Y(n_509)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_511),
.Y(n_527)
);

OAI21xp5_ASAP7_75t_SL g513 ( 
.A1(n_495),
.A2(n_504),
.B(n_500),
.Y(n_513)
);

AND2x2_ASAP7_75t_SL g523 ( 
.A(n_513),
.B(n_514),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_SL g521 ( 
.A(n_515),
.B(n_508),
.Y(n_521)
);

NOR2xp33_ASAP7_75t_L g520 ( 
.A(n_501),
.B(n_461),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_520),
.B(n_512),
.Y(n_526)
);

NOR3xp33_ASAP7_75t_L g528 ( 
.A(n_521),
.B(n_526),
.C(n_512),
.Y(n_528)
);

OAI21xp5_ASAP7_75t_SL g522 ( 
.A1(n_516),
.A2(n_495),
.B(n_499),
.Y(n_522)
);

XNOR2xp5_ASAP7_75t_L g529 ( 
.A(n_522),
.B(n_524),
.Y(n_529)
);

XOR2xp5_ASAP7_75t_L g524 ( 
.A(n_510),
.B(n_483),
.Y(n_524)
);

AOI21xp5_ASAP7_75t_L g525 ( 
.A1(n_518),
.A2(n_505),
.B(n_483),
.Y(n_525)
);

OAI21xp5_ASAP7_75t_SL g531 ( 
.A1(n_525),
.A2(n_517),
.B(n_519),
.Y(n_531)
);

AOI21x1_ASAP7_75t_SL g534 ( 
.A1(n_528),
.A2(n_531),
.B(n_497),
.Y(n_534)
);

INVxp67_ASAP7_75t_L g530 ( 
.A(n_521),
.Y(n_530)
);

MAJIxp5_ASAP7_75t_L g532 ( 
.A(n_530),
.B(n_523),
.C(n_527),
.Y(n_532)
);

MAJx2_ASAP7_75t_L g535 ( 
.A(n_532),
.B(n_533),
.C(n_514),
.Y(n_535)
);

MAJIxp5_ASAP7_75t_L g533 ( 
.A(n_529),
.B(n_523),
.C(n_513),
.Y(n_533)
);

MAJIxp5_ASAP7_75t_L g536 ( 
.A(n_534),
.B(n_515),
.C(n_474),
.Y(n_536)
);

OAI21xp5_ASAP7_75t_L g537 ( 
.A1(n_535),
.A2(n_536),
.B(n_476),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g538 ( 
.A(n_537),
.B(n_484),
.Y(n_538)
);

MAJIxp5_ASAP7_75t_L g539 ( 
.A(n_538),
.B(n_484),
.C(n_16),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_SL g540 ( 
.A(n_539),
.B(n_16),
.Y(n_540)
);


endmodule