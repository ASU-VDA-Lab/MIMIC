module fake_netlist_1_3130_n_520 (n_53, n_67, n_45, n_20, n_2, n_38, n_44, n_64, n_54, n_62, n_36, n_47, n_37, n_69, n_34, n_5, n_23, n_8, n_28, n_31, n_22, n_46, n_48, n_58, n_57, n_11, n_25, n_16, n_26, n_13, n_30, n_33, n_50, n_52, n_49, n_59, n_73, n_3, n_18, n_60, n_66, n_32, n_0, n_41, n_1, n_35, n_55, n_65, n_12, n_9, n_70, n_17, n_63, n_14, n_10, n_15, n_56, n_71, n_42, n_24, n_19, n_61, n_21, n_6, n_4, n_74, n_72, n_51, n_29, n_43, n_7, n_68, n_40, n_27, n_39, n_520);
input n_53;
input n_67;
input n_45;
input n_20;
input n_2;
input n_38;
input n_44;
input n_64;
input n_54;
input n_62;
input n_36;
input n_47;
input n_37;
input n_69;
input n_34;
input n_5;
input n_23;
input n_8;
input n_28;
input n_31;
input n_22;
input n_46;
input n_48;
input n_58;
input n_57;
input n_11;
input n_25;
input n_16;
input n_26;
input n_13;
input n_30;
input n_33;
input n_50;
input n_52;
input n_49;
input n_59;
input n_73;
input n_3;
input n_18;
input n_60;
input n_66;
input n_32;
input n_0;
input n_41;
input n_1;
input n_35;
input n_55;
input n_65;
input n_12;
input n_9;
input n_70;
input n_17;
input n_63;
input n_14;
input n_10;
input n_15;
input n_56;
input n_71;
input n_42;
input n_24;
input n_19;
input n_61;
input n_21;
input n_6;
input n_4;
input n_74;
input n_72;
input n_51;
input n_29;
input n_43;
input n_7;
input n_68;
input n_40;
input n_27;
input n_39;
output n_520;
wire n_117;
wire n_361;
wire n_513;
wire n_185;
wire n_407;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_154;
wire n_328;
wire n_468;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_353;
wire n_206;
wire n_288;
wire n_383;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_211;
wire n_334;
wire n_389;
wire n_436;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_231;
wire n_452;
wire n_518;
wire n_298;
wire n_411;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_228;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_366;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_244;
wire n_119;
wire n_141;
wire n_517;
wire n_479;
wire n_97;
wire n_167;
wire n_447;
wire n_171;
wire n_196;
wire n_192;
wire n_502;
wire n_312;
wire n_455;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_367;
wire n_250;
wire n_85;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_293;
wire n_506;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_381;
wire n_304;
wire n_399;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_77;
wire n_404;
wire n_369;
wire n_509;
wire n_172;
wire n_329;
wire n_251;
wire n_218;
wire n_507;
wire n_271;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_133;
wire n_149;
wire n_81;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_107;
wire n_403;
wire n_516;
wire n_254;
wire n_262;
wire n_239;
wire n_439;
wire n_87;
wire n_379;
wire n_98;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_370;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_245;
wire n_90;
wire n_357;
wire n_260;
wire n_78;
wire n_197;
wire n_201;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_265;
wire n_264;
wire n_200;
wire n_208;
wire n_126;
wire n_178;
wire n_118;
wire n_365;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_75;
wire n_376;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_76;
wire n_435;
wire n_216;
wire n_147;
wire n_148;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_225;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_121;
wire n_497;
wire n_339;
wire n_240;
wire n_378;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_335;
wire n_272;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_198;
wire n_169;
wire n_424;
wire n_156;
wire n_124;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_418;
wire n_493;
wire n_380;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_487;
wire n_451;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_258;
wire n_253;
wire n_515;
wire n_84;
wire n_266;
wire n_213;
wire n_182;
wire n_492;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_469;
wire n_123;
wire n_457;
wire n_223;
wire n_494;
wire n_480;
wire n_372;
wire n_453;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_425;
wire n_332;
wire n_414;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_406;
wire n_395;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
HB1xp67_ASAP7_75t_L g75 ( .A(n_31), .Y(n_75) );
CKINVDCx20_ASAP7_75t_R g76 ( .A(n_56), .Y(n_76) );
INVx1_ASAP7_75t_L g77 ( .A(n_24), .Y(n_77) );
INVxp33_ASAP7_75t_SL g78 ( .A(n_30), .Y(n_78) );
INVxp33_ASAP7_75t_L g79 ( .A(n_60), .Y(n_79) );
CKINVDCx5p33_ASAP7_75t_R g80 ( .A(n_0), .Y(n_80) );
CKINVDCx5p33_ASAP7_75t_R g81 ( .A(n_28), .Y(n_81) );
CKINVDCx5p33_ASAP7_75t_R g82 ( .A(n_8), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_72), .Y(n_83) );
CKINVDCx14_ASAP7_75t_R g84 ( .A(n_51), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_74), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_69), .Y(n_86) );
INVx2_ASAP7_75t_L g87 ( .A(n_16), .Y(n_87) );
INVx2_ASAP7_75t_L g88 ( .A(n_11), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_27), .Y(n_89) );
INVx2_ASAP7_75t_L g90 ( .A(n_36), .Y(n_90) );
INVx2_ASAP7_75t_L g91 ( .A(n_26), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_1), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_21), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_61), .Y(n_94) );
INVxp33_ASAP7_75t_SL g95 ( .A(n_39), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_0), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_70), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_49), .Y(n_98) );
CKINVDCx16_ASAP7_75t_R g99 ( .A(n_6), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_1), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_7), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_41), .Y(n_102) );
INVxp67_ASAP7_75t_SL g103 ( .A(n_5), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_11), .Y(n_104) );
CKINVDCx16_ASAP7_75t_R g105 ( .A(n_9), .Y(n_105) );
INVx2_ASAP7_75t_L g106 ( .A(n_2), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_5), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_6), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_88), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_88), .Y(n_110) );
AND2x4_ASAP7_75t_L g111 ( .A(n_88), .B(n_2), .Y(n_111) );
INVx2_ASAP7_75t_L g112 ( .A(n_90), .Y(n_112) );
AND2x2_ASAP7_75t_L g113 ( .A(n_99), .B(n_3), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_106), .Y(n_114) );
AND2x2_ASAP7_75t_L g115 ( .A(n_99), .B(n_3), .Y(n_115) );
AND2x2_ASAP7_75t_L g116 ( .A(n_105), .B(n_4), .Y(n_116) );
INVx2_ASAP7_75t_L g117 ( .A(n_90), .Y(n_117) );
NAND2xp5_ASAP7_75t_SL g118 ( .A(n_79), .B(n_4), .Y(n_118) );
CKINVDCx5p33_ASAP7_75t_R g119 ( .A(n_76), .Y(n_119) );
INVx2_ASAP7_75t_L g120 ( .A(n_90), .Y(n_120) );
INVx2_ASAP7_75t_L g121 ( .A(n_91), .Y(n_121) );
BUFx6f_ASAP7_75t_L g122 ( .A(n_91), .Y(n_122) );
NAND2xp5_ASAP7_75t_L g123 ( .A(n_75), .B(n_7), .Y(n_123) );
BUFx2_ASAP7_75t_L g124 ( .A(n_84), .Y(n_124) );
BUFx3_ASAP7_75t_L g125 ( .A(n_91), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_106), .Y(n_126) );
INVx1_ASAP7_75t_L g127 ( .A(n_106), .Y(n_127) );
NAND2xp5_ASAP7_75t_SL g128 ( .A(n_77), .B(n_8), .Y(n_128) );
BUFx3_ASAP7_75t_L g129 ( .A(n_77), .Y(n_129) );
INVx2_ASAP7_75t_L g130 ( .A(n_83), .Y(n_130) );
OA21x2_ASAP7_75t_L g131 ( .A1(n_83), .A2(n_9), .B(n_10), .Y(n_131) );
AND2x4_ASAP7_75t_L g132 ( .A(n_111), .B(n_87), .Y(n_132) );
OR2x6_ASAP7_75t_L g133 ( .A(n_113), .B(n_92), .Y(n_133) );
INVx1_ASAP7_75t_L g134 ( .A(n_120), .Y(n_134) );
BUFx3_ASAP7_75t_L g135 ( .A(n_111), .Y(n_135) );
AND2x4_ASAP7_75t_L g136 ( .A(n_111), .B(n_87), .Y(n_136) );
INVx2_ASAP7_75t_L g137 ( .A(n_122), .Y(n_137) );
BUFx2_ASAP7_75t_L g138 ( .A(n_124), .Y(n_138) );
CKINVDCx5p33_ASAP7_75t_R g139 ( .A(n_119), .Y(n_139) );
CKINVDCx20_ASAP7_75t_R g140 ( .A(n_124), .Y(n_140) );
INVx2_ASAP7_75t_L g141 ( .A(n_122), .Y(n_141) );
NAND2x1p5_ASAP7_75t_L g142 ( .A(n_131), .B(n_85), .Y(n_142) );
INVx1_ASAP7_75t_SL g143 ( .A(n_113), .Y(n_143) );
NAND2xp5_ASAP7_75t_L g144 ( .A(n_129), .B(n_85), .Y(n_144) );
INVx1_ASAP7_75t_L g145 ( .A(n_120), .Y(n_145) );
OAI22xp5_ASAP7_75t_L g146 ( .A1(n_113), .A2(n_105), .B1(n_107), .B2(n_108), .Y(n_146) );
INVx1_ASAP7_75t_L g147 ( .A(n_120), .Y(n_147) );
INVx1_ASAP7_75t_L g148 ( .A(n_120), .Y(n_148) );
BUFx3_ASAP7_75t_L g149 ( .A(n_111), .Y(n_149) );
INVx1_ASAP7_75t_L g150 ( .A(n_112), .Y(n_150) );
INVx4_ASAP7_75t_L g151 ( .A(n_111), .Y(n_151) );
HB1xp67_ASAP7_75t_L g152 ( .A(n_124), .Y(n_152) );
NAND2xp5_ASAP7_75t_SL g153 ( .A(n_129), .B(n_81), .Y(n_153) );
INVx2_ASAP7_75t_L g154 ( .A(n_122), .Y(n_154) );
AND2x4_ASAP7_75t_L g155 ( .A(n_129), .B(n_92), .Y(n_155) );
NAND2xp5_ASAP7_75t_L g156 ( .A(n_129), .B(n_102), .Y(n_156) );
INVx1_ASAP7_75t_L g157 ( .A(n_112), .Y(n_157) );
AND2x4_ASAP7_75t_L g158 ( .A(n_133), .B(n_115), .Y(n_158) );
INVx1_ASAP7_75t_L g159 ( .A(n_134), .Y(n_159) );
BUFx3_ASAP7_75t_L g160 ( .A(n_135), .Y(n_160) );
CKINVDCx5p33_ASAP7_75t_R g161 ( .A(n_139), .Y(n_161) );
NAND2xp5_ASAP7_75t_SL g162 ( .A(n_138), .B(n_123), .Y(n_162) );
NAND2xp5_ASAP7_75t_L g163 ( .A(n_143), .B(n_123), .Y(n_163) );
INVx1_ASAP7_75t_L g164 ( .A(n_134), .Y(n_164) );
AND2x6_ASAP7_75t_L g165 ( .A(n_135), .B(n_115), .Y(n_165) );
INVx1_ASAP7_75t_L g166 ( .A(n_145), .Y(n_166) );
A2O1A1Ixp33_ASAP7_75t_L g167 ( .A1(n_135), .A2(n_125), .B(n_130), .C(n_117), .Y(n_167) );
INVx1_ASAP7_75t_L g168 ( .A(n_145), .Y(n_168) );
NAND2xp5_ASAP7_75t_L g169 ( .A(n_143), .B(n_115), .Y(n_169) );
INVx1_ASAP7_75t_L g170 ( .A(n_147), .Y(n_170) );
INVxp67_ASAP7_75t_SL g171 ( .A(n_152), .Y(n_171) );
NAND2xp5_ASAP7_75t_L g172 ( .A(n_151), .B(n_116), .Y(n_172) );
NAND2xp5_ASAP7_75t_L g173 ( .A(n_151), .B(n_116), .Y(n_173) );
AND2x4_ASAP7_75t_L g174 ( .A(n_133), .B(n_116), .Y(n_174) );
HB1xp67_ASAP7_75t_L g175 ( .A(n_152), .Y(n_175) );
HB1xp67_ASAP7_75t_L g176 ( .A(n_138), .Y(n_176) );
INVx2_ASAP7_75t_L g177 ( .A(n_147), .Y(n_177) );
INVx1_ASAP7_75t_L g178 ( .A(n_148), .Y(n_178) );
INVx2_ASAP7_75t_L g179 ( .A(n_148), .Y(n_179) );
BUFx6f_ASAP7_75t_L g180 ( .A(n_149), .Y(n_180) );
AND2x4_ASAP7_75t_L g181 ( .A(n_133), .B(n_128), .Y(n_181) );
BUFx6f_ASAP7_75t_L g182 ( .A(n_149), .Y(n_182) );
AOI22x1_ASAP7_75t_SL g183 ( .A1(n_140), .A2(n_80), .B1(n_82), .B2(n_103), .Y(n_183) );
AOI22xp5_ASAP7_75t_L g184 ( .A1(n_133), .A2(n_118), .B1(n_128), .B2(n_95), .Y(n_184) );
INVx1_ASAP7_75t_L g185 ( .A(n_151), .Y(n_185) );
BUFx6f_ASAP7_75t_L g186 ( .A(n_149), .Y(n_186) );
OR2x4_ASAP7_75t_L g187 ( .A(n_146), .B(n_96), .Y(n_187) );
INVx1_ASAP7_75t_L g188 ( .A(n_151), .Y(n_188) );
INVx1_ASAP7_75t_L g189 ( .A(n_150), .Y(n_189) );
AND2x4_ASAP7_75t_L g190 ( .A(n_133), .B(n_118), .Y(n_190) );
INVx2_ASAP7_75t_L g191 ( .A(n_142), .Y(n_191) );
INVx2_ASAP7_75t_L g192 ( .A(n_177), .Y(n_192) );
BUFx3_ASAP7_75t_L g193 ( .A(n_180), .Y(n_193) );
INVx2_ASAP7_75t_L g194 ( .A(n_177), .Y(n_194) );
NAND2xp5_ASAP7_75t_L g195 ( .A(n_163), .B(n_133), .Y(n_195) );
INVx2_ASAP7_75t_SL g196 ( .A(n_158), .Y(n_196) );
OR2x6_ASAP7_75t_L g197 ( .A(n_158), .B(n_132), .Y(n_197) );
BUFx2_ASAP7_75t_SL g198 ( .A(n_158), .Y(n_198) );
BUFx3_ASAP7_75t_L g199 ( .A(n_180), .Y(n_199) );
AOI22xp33_ASAP7_75t_L g200 ( .A1(n_174), .A2(n_146), .B1(n_132), .B2(n_136), .Y(n_200) );
BUFx3_ASAP7_75t_L g201 ( .A(n_165), .Y(n_201) );
INVx1_ASAP7_75t_L g202 ( .A(n_159), .Y(n_202) );
INVx3_ASAP7_75t_L g203 ( .A(n_180), .Y(n_203) );
NAND2x1_ASAP7_75t_L g204 ( .A(n_179), .B(n_132), .Y(n_204) );
BUFx6f_ASAP7_75t_L g205 ( .A(n_180), .Y(n_205) );
INVx1_ASAP7_75t_L g206 ( .A(n_159), .Y(n_206) );
NAND2xp5_ASAP7_75t_L g207 ( .A(n_172), .B(n_155), .Y(n_207) );
INVx1_ASAP7_75t_L g208 ( .A(n_164), .Y(n_208) );
INVx2_ASAP7_75t_SL g209 ( .A(n_174), .Y(n_209) );
AOI22xp5_ASAP7_75t_L g210 ( .A1(n_174), .A2(n_155), .B1(n_132), .B2(n_136), .Y(n_210) );
NAND2xp5_ASAP7_75t_L g211 ( .A(n_173), .B(n_155), .Y(n_211) );
INVx1_ASAP7_75t_L g212 ( .A(n_164), .Y(n_212) );
INVx1_ASAP7_75t_L g213 ( .A(n_166), .Y(n_213) );
INVx4_ASAP7_75t_L g214 ( .A(n_165), .Y(n_214) );
BUFx6f_ASAP7_75t_L g215 ( .A(n_180), .Y(n_215) );
BUFx2_ASAP7_75t_L g216 ( .A(n_165), .Y(n_216) );
NAND2xp5_ASAP7_75t_L g217 ( .A(n_169), .B(n_155), .Y(n_217) );
INVx1_ASAP7_75t_L g218 ( .A(n_166), .Y(n_218) );
INVx1_ASAP7_75t_L g219 ( .A(n_168), .Y(n_219) );
NAND2xp5_ASAP7_75t_L g220 ( .A(n_165), .B(n_136), .Y(n_220) );
INVx1_ASAP7_75t_SL g221 ( .A(n_176), .Y(n_221) );
CKINVDCx5p33_ASAP7_75t_R g222 ( .A(n_161), .Y(n_222) );
A2O1A1Ixp33_ASAP7_75t_L g223 ( .A1(n_168), .A2(n_144), .B(n_156), .C(n_136), .Y(n_223) );
AOI21xp5_ASAP7_75t_L g224 ( .A1(n_191), .A2(n_153), .B(n_142), .Y(n_224) );
NAND2xp5_ASAP7_75t_L g225 ( .A(n_202), .B(n_165), .Y(n_225) );
CKINVDCx20_ASAP7_75t_R g226 ( .A(n_222), .Y(n_226) );
AOI22xp33_ASAP7_75t_L g227 ( .A1(n_197), .A2(n_165), .B1(n_190), .B2(n_181), .Y(n_227) );
O2A1O1Ixp33_ASAP7_75t_SL g228 ( .A1(n_223), .A2(n_167), .B(n_189), .C(n_170), .Y(n_228) );
AND2x2_ASAP7_75t_L g229 ( .A(n_198), .B(n_179), .Y(n_229) );
OR2x6_ASAP7_75t_L g230 ( .A(n_198), .B(n_181), .Y(n_230) );
AOI22xp33_ASAP7_75t_L g231 ( .A1(n_197), .A2(n_165), .B1(n_190), .B2(n_181), .Y(n_231) );
INVx3_ASAP7_75t_L g232 ( .A(n_214), .Y(n_232) );
BUFx3_ASAP7_75t_L g233 ( .A(n_201), .Y(n_233) );
CKINVDCx6p67_ASAP7_75t_R g234 ( .A(n_201), .Y(n_234) );
AOI22xp33_ASAP7_75t_L g235 ( .A1(n_197), .A2(n_190), .B1(n_181), .B2(n_175), .Y(n_235) );
AOI221xp5_ASAP7_75t_L g236 ( .A1(n_200), .A2(n_171), .B1(n_162), .B2(n_161), .C(n_187), .Y(n_236) );
AOI21xp5_ASAP7_75t_L g237 ( .A1(n_224), .A2(n_191), .B(n_189), .Y(n_237) );
NAND2xp5_ASAP7_75t_L g238 ( .A(n_202), .B(n_170), .Y(n_238) );
AOI22xp33_ASAP7_75t_L g239 ( .A1(n_197), .A2(n_160), .B1(n_188), .B2(n_185), .Y(n_239) );
AOI22xp33_ASAP7_75t_L g240 ( .A1(n_197), .A2(n_160), .B1(n_188), .B2(n_185), .Y(n_240) );
AOI21xp5_ASAP7_75t_L g241 ( .A1(n_206), .A2(n_178), .B(n_142), .Y(n_241) );
O2A1O1Ixp33_ASAP7_75t_L g242 ( .A1(n_195), .A2(n_144), .B(n_156), .C(n_130), .Y(n_242) );
OR2x2_ASAP7_75t_L g243 ( .A(n_221), .B(n_178), .Y(n_243) );
OAI211xp5_ASAP7_75t_L g244 ( .A1(n_210), .A2(n_184), .B(n_204), .C(n_217), .Y(n_244) );
AOI22xp33_ASAP7_75t_L g245 ( .A1(n_214), .A2(n_186), .B1(n_182), .B2(n_142), .Y(n_245) );
INVx2_ASAP7_75t_L g246 ( .A(n_192), .Y(n_246) );
AO31x2_ASAP7_75t_L g247 ( .A1(n_206), .A2(n_130), .A3(n_121), .B(n_117), .Y(n_247) );
AOI22xp33_ASAP7_75t_L g248 ( .A1(n_214), .A2(n_186), .B1(n_182), .B2(n_78), .Y(n_248) );
INVx1_ASAP7_75t_L g249 ( .A(n_208), .Y(n_249) );
AOI221xp5_ASAP7_75t_L g250 ( .A1(n_236), .A2(n_244), .B1(n_228), .B2(n_235), .C(n_249), .Y(n_250) );
AOI332xp33_ASAP7_75t_L g251 ( .A1(n_249), .A2(n_96), .A3(n_100), .B1(n_101), .B2(n_104), .B3(n_107), .C1(n_108), .C2(n_114), .Y(n_251) );
BUFx2_ASAP7_75t_L g252 ( .A(n_230), .Y(n_252) );
AOI22xp33_ASAP7_75t_L g253 ( .A1(n_227), .A2(n_214), .B1(n_216), .B2(n_209), .Y(n_253) );
OAI221xp5_ASAP7_75t_L g254 ( .A1(n_231), .A2(n_210), .B1(n_220), .B2(n_209), .C(n_196), .Y(n_254) );
AOI22xp33_ASAP7_75t_L g255 ( .A1(n_230), .A2(n_216), .B1(n_196), .B2(n_218), .Y(n_255) );
AOI221xp5_ASAP7_75t_L g256 ( .A1(n_243), .A2(n_211), .B1(n_207), .B2(n_213), .C(n_212), .Y(n_256) );
OAI22xp5_ASAP7_75t_L g257 ( .A1(n_238), .A2(n_219), .B1(n_218), .B2(n_208), .Y(n_257) );
OAI21xp5_ASAP7_75t_L g258 ( .A1(n_241), .A2(n_219), .B(n_212), .Y(n_258) );
AND2x4_ASAP7_75t_L g259 ( .A(n_230), .B(n_213), .Y(n_259) );
OR2x2_ASAP7_75t_L g260 ( .A(n_243), .B(n_192), .Y(n_260) );
HB1xp67_ASAP7_75t_L g261 ( .A(n_229), .Y(n_261) );
INVx2_ASAP7_75t_L g262 ( .A(n_246), .Y(n_262) );
AOI21xp5_ASAP7_75t_L g263 ( .A1(n_238), .A2(n_194), .B(n_204), .Y(n_263) );
OAI211xp5_ASAP7_75t_SL g264 ( .A1(n_239), .A2(n_104), .B(n_100), .C(n_101), .Y(n_264) );
OAI22xp5_ASAP7_75t_L g265 ( .A1(n_230), .A2(n_187), .B1(n_194), .B2(n_193), .Y(n_265) );
OAI22xp5_ASAP7_75t_L g266 ( .A1(n_230), .A2(n_187), .B1(n_199), .B2(n_193), .Y(n_266) );
AOI22xp33_ASAP7_75t_L g267 ( .A1(n_229), .A2(n_186), .B1(n_182), .B2(n_199), .Y(n_267) );
NAND2xp5_ASAP7_75t_L g268 ( .A(n_246), .B(n_203), .Y(n_268) );
AOI22xp33_ASAP7_75t_L g269 ( .A1(n_225), .A2(n_186), .B1(n_182), .B2(n_199), .Y(n_269) );
OAI22xp5_ASAP7_75t_L g270 ( .A1(n_225), .A2(n_193), .B1(n_215), .B2(n_205), .Y(n_270) );
NAND2xp5_ASAP7_75t_L g271 ( .A(n_260), .B(n_246), .Y(n_271) );
AOI21xp5_ASAP7_75t_SL g272 ( .A1(n_257), .A2(n_233), .B(n_242), .Y(n_272) );
OAI22xp5_ASAP7_75t_L g273 ( .A1(n_256), .A2(n_234), .B1(n_240), .B2(n_245), .Y(n_273) );
OAI211xp5_ASAP7_75t_L g274 ( .A1(n_251), .A2(n_109), .B(n_110), .C(n_114), .Y(n_274) );
INVx2_ASAP7_75t_L g275 ( .A(n_262), .Y(n_275) );
AOI21xp5_ASAP7_75t_L g276 ( .A1(n_263), .A2(n_237), .B(n_205), .Y(n_276) );
AOI221xp5_ASAP7_75t_SL g277 ( .A1(n_250), .A2(n_248), .B1(n_109), .B2(n_110), .C(n_127), .Y(n_277) );
NAND2xp5_ASAP7_75t_L g278 ( .A(n_260), .B(n_247), .Y(n_278) );
INVx2_ASAP7_75t_L g279 ( .A(n_262), .Y(n_279) );
NOR2xp33_ASAP7_75t_L g280 ( .A(n_254), .B(n_183), .Y(n_280) );
AOI221xp5_ASAP7_75t_L g281 ( .A1(n_264), .A2(n_127), .B1(n_126), .B2(n_125), .C(n_112), .Y(n_281) );
AND2x2_ASAP7_75t_L g282 ( .A(n_261), .B(n_247), .Y(n_282) );
OAI33xp33_ASAP7_75t_L g283 ( .A1(n_265), .A2(n_126), .A3(n_89), .B1(n_93), .B2(n_94), .B3(n_97), .Y(n_283) );
INVx2_ASAP7_75t_L g284 ( .A(n_259), .Y(n_284) );
OAI221xp5_ASAP7_75t_L g285 ( .A1(n_255), .A2(n_117), .B1(n_121), .B2(n_183), .C(n_125), .Y(n_285) );
BUFx2_ASAP7_75t_L g286 ( .A(n_252), .Y(n_286) );
OAI211xp5_ASAP7_75t_L g287 ( .A1(n_251), .A2(n_131), .B(n_89), .C(n_98), .Y(n_287) );
NAND2xp5_ASAP7_75t_SL g288 ( .A(n_259), .B(n_226), .Y(n_288) );
INVx3_ASAP7_75t_SL g289 ( .A(n_259), .Y(n_289) );
INVx1_ASAP7_75t_L g290 ( .A(n_258), .Y(n_290) );
INVx1_ASAP7_75t_L g291 ( .A(n_258), .Y(n_291) );
AOI31xp33_ASAP7_75t_L g292 ( .A1(n_266), .A2(n_86), .A3(n_93), .B(n_94), .Y(n_292) );
AND2x2_ASAP7_75t_L g293 ( .A(n_275), .B(n_247), .Y(n_293) );
INVx1_ASAP7_75t_SL g294 ( .A(n_289), .Y(n_294) );
AOI22xp33_ASAP7_75t_L g295 ( .A1(n_280), .A2(n_252), .B1(n_253), .B2(n_233), .Y(n_295) );
AND2x2_ASAP7_75t_SL g296 ( .A(n_286), .B(n_267), .Y(n_296) );
BUFx2_ASAP7_75t_L g297 ( .A(n_286), .Y(n_297) );
INVx3_ASAP7_75t_L g298 ( .A(n_275), .Y(n_298) );
INVx5_ASAP7_75t_L g299 ( .A(n_275), .Y(n_299) );
AND2x2_ASAP7_75t_L g300 ( .A(n_279), .B(n_247), .Y(n_300) );
AND2x2_ASAP7_75t_L g301 ( .A(n_279), .B(n_247), .Y(n_301) );
INVx1_ASAP7_75t_SL g302 ( .A(n_289), .Y(n_302) );
AND2x2_ASAP7_75t_L g303 ( .A(n_279), .B(n_131), .Y(n_303) );
INVx1_ASAP7_75t_L g304 ( .A(n_290), .Y(n_304) );
AOI211xp5_ASAP7_75t_L g305 ( .A1(n_287), .A2(n_86), .B(n_97), .C(n_98), .Y(n_305) );
AOI22xp33_ASAP7_75t_L g306 ( .A1(n_283), .A2(n_125), .B1(n_102), .B2(n_269), .Y(n_306) );
AOI22xp33_ASAP7_75t_L g307 ( .A1(n_273), .A2(n_233), .B1(n_121), .B2(n_270), .Y(n_307) );
OAI22xp33_ASAP7_75t_L g308 ( .A1(n_292), .A2(n_234), .B1(n_268), .B2(n_232), .Y(n_308) );
INVxp67_ASAP7_75t_L g309 ( .A(n_278), .Y(n_309) );
INVx2_ASAP7_75t_L g310 ( .A(n_290), .Y(n_310) );
AND2x2_ASAP7_75t_L g311 ( .A(n_291), .B(n_131), .Y(n_311) );
INVx1_ASAP7_75t_SL g312 ( .A(n_289), .Y(n_312) );
AOI22xp5_ASAP7_75t_L g313 ( .A1(n_277), .A2(n_131), .B1(n_232), .B2(n_157), .Y(n_313) );
AND2x2_ASAP7_75t_SL g314 ( .A(n_282), .B(n_232), .Y(n_314) );
INVx1_ASAP7_75t_L g315 ( .A(n_291), .Y(n_315) );
INVx1_ASAP7_75t_L g316 ( .A(n_282), .Y(n_316) );
AOI33xp33_ASAP7_75t_L g317 ( .A1(n_284), .A2(n_150), .A3(n_157), .B1(n_137), .B2(n_154), .B3(n_141), .Y(n_317) );
INVx1_ASAP7_75t_L g318 ( .A(n_284), .Y(n_318) );
AND2x2_ASAP7_75t_L g319 ( .A(n_284), .B(n_131), .Y(n_319) );
NAND2xp5_ASAP7_75t_SL g320 ( .A(n_292), .B(n_122), .Y(n_320) );
AND2x2_ASAP7_75t_L g321 ( .A(n_271), .B(n_122), .Y(n_321) );
AOI221xp5_ASAP7_75t_L g322 ( .A1(n_285), .A2(n_122), .B1(n_182), .B2(n_186), .C(n_203), .Y(n_322) );
AOI22xp33_ASAP7_75t_L g323 ( .A1(n_273), .A2(n_203), .B1(n_205), .B2(n_215), .Y(n_323) );
NOR3xp33_ASAP7_75t_SL g324 ( .A(n_308), .B(n_288), .C(n_274), .Y(n_324) );
INVx2_ASAP7_75t_L g325 ( .A(n_298), .Y(n_325) );
NAND4xp25_ASAP7_75t_SL g326 ( .A(n_294), .B(n_272), .C(n_277), .D(n_281), .Y(n_326) );
INVx1_ASAP7_75t_L g327 ( .A(n_316), .Y(n_327) );
OR2x2_ASAP7_75t_L g328 ( .A(n_309), .B(n_272), .Y(n_328) );
NOR2x1_ASAP7_75t_L g329 ( .A(n_308), .B(n_122), .Y(n_329) );
INVx1_ASAP7_75t_L g330 ( .A(n_318), .Y(n_330) );
INVx2_ASAP7_75t_L g331 ( .A(n_298), .Y(n_331) );
INVx1_ASAP7_75t_SL g332 ( .A(n_294), .Y(n_332) );
INVx1_ASAP7_75t_L g333 ( .A(n_318), .Y(n_333) );
OAI322xp33_ASAP7_75t_L g334 ( .A1(n_309), .A2(n_122), .A3(n_12), .B1(n_13), .B2(n_14), .C1(n_15), .C2(n_10), .Y(n_334) );
OR2x2_ASAP7_75t_L g335 ( .A(n_316), .B(n_12), .Y(n_335) );
OR2x2_ASAP7_75t_L g336 ( .A(n_297), .B(n_13), .Y(n_336) );
OAI21xp33_ASAP7_75t_L g337 ( .A1(n_323), .A2(n_154), .B(n_141), .Y(n_337) );
NAND2xp5_ASAP7_75t_SL g338 ( .A(n_302), .B(n_276), .Y(n_338) );
NAND2xp5_ASAP7_75t_L g339 ( .A(n_293), .B(n_14), .Y(n_339) );
AND2x2_ASAP7_75t_L g340 ( .A(n_293), .B(n_15), .Y(n_340) );
AND2x4_ASAP7_75t_SL g341 ( .A(n_293), .B(n_215), .Y(n_341) );
AND2x2_ASAP7_75t_SL g342 ( .A(n_314), .B(n_215), .Y(n_342) );
AND2x2_ASAP7_75t_L g343 ( .A(n_300), .B(n_16), .Y(n_343) );
HB1xp67_ASAP7_75t_L g344 ( .A(n_297), .Y(n_344) );
INVx1_ASAP7_75t_L g345 ( .A(n_321), .Y(n_345) );
NOR3xp33_ASAP7_75t_L g346 ( .A(n_320), .B(n_137), .C(n_141), .Y(n_346) );
NAND2xp5_ASAP7_75t_L g347 ( .A(n_300), .B(n_301), .Y(n_347) );
NAND4xp25_ASAP7_75t_L g348 ( .A(n_307), .B(n_154), .C(n_137), .D(n_19), .Y(n_348) );
INVx2_ASAP7_75t_L g349 ( .A(n_298), .Y(n_349) );
NAND2xp5_ASAP7_75t_L g350 ( .A(n_300), .B(n_17), .Y(n_350) );
INVx1_ASAP7_75t_L g351 ( .A(n_304), .Y(n_351) );
INVx2_ASAP7_75t_L g352 ( .A(n_298), .Y(n_352) );
NAND2xp5_ASAP7_75t_L g353 ( .A(n_301), .B(n_17), .Y(n_353) );
NOR2xp33_ASAP7_75t_L g354 ( .A(n_302), .B(n_18), .Y(n_354) );
AND2x2_ASAP7_75t_L g355 ( .A(n_301), .B(n_18), .Y(n_355) );
INVx1_ASAP7_75t_L g356 ( .A(n_304), .Y(n_356) );
HB1xp67_ASAP7_75t_L g357 ( .A(n_299), .Y(n_357) );
INVx1_ASAP7_75t_L g358 ( .A(n_321), .Y(n_358) );
OR2x2_ASAP7_75t_L g359 ( .A(n_315), .B(n_19), .Y(n_359) );
INVx1_ASAP7_75t_SL g360 ( .A(n_312), .Y(n_360) );
NAND2xp5_ASAP7_75t_L g361 ( .A(n_321), .B(n_20), .Y(n_361) );
BUFx2_ASAP7_75t_L g362 ( .A(n_299), .Y(n_362) );
AND2x2_ASAP7_75t_L g363 ( .A(n_310), .B(n_20), .Y(n_363) );
INVx1_ASAP7_75t_L g364 ( .A(n_315), .Y(n_364) );
AND2x2_ASAP7_75t_L g365 ( .A(n_310), .B(n_22), .Y(n_365) );
INVx3_ASAP7_75t_L g366 ( .A(n_299), .Y(n_366) );
INVx2_ASAP7_75t_L g367 ( .A(n_299), .Y(n_367) );
OR2x2_ASAP7_75t_L g368 ( .A(n_310), .B(n_203), .Y(n_368) );
AOI22xp5_ASAP7_75t_L g369 ( .A1(n_295), .A2(n_215), .B1(n_205), .B2(n_29), .Y(n_369) );
AND2x2_ASAP7_75t_L g370 ( .A(n_347), .B(n_314), .Y(n_370) );
OR2x2_ASAP7_75t_L g371 ( .A(n_344), .B(n_312), .Y(n_371) );
NOR2xp33_ASAP7_75t_L g372 ( .A(n_332), .B(n_314), .Y(n_372) );
INVx3_ASAP7_75t_L g373 ( .A(n_366), .Y(n_373) );
NOR2xp33_ASAP7_75t_L g374 ( .A(n_360), .B(n_296), .Y(n_374) );
OR2x2_ASAP7_75t_L g375 ( .A(n_327), .B(n_328), .Y(n_375) );
INVx1_ASAP7_75t_L g376 ( .A(n_351), .Y(n_376) );
NOR2xp33_ASAP7_75t_L g377 ( .A(n_354), .B(n_296), .Y(n_377) );
NAND2xp5_ASAP7_75t_L g378 ( .A(n_340), .B(n_299), .Y(n_378) );
NAND2xp5_ASAP7_75t_L g379 ( .A(n_340), .B(n_299), .Y(n_379) );
AND2x2_ASAP7_75t_L g380 ( .A(n_351), .B(n_356), .Y(n_380) );
OR2x2_ASAP7_75t_L g381 ( .A(n_328), .B(n_299), .Y(n_381) );
AND2x2_ASAP7_75t_L g382 ( .A(n_356), .B(n_311), .Y(n_382) );
NAND2xp5_ASAP7_75t_L g383 ( .A(n_343), .B(n_296), .Y(n_383) );
NAND2xp5_ASAP7_75t_L g384 ( .A(n_343), .B(n_307), .Y(n_384) );
INVxp67_ASAP7_75t_L g385 ( .A(n_357), .Y(n_385) );
AND2x2_ASAP7_75t_L g386 ( .A(n_364), .B(n_311), .Y(n_386) );
NOR2xp33_ASAP7_75t_L g387 ( .A(n_361), .B(n_23), .Y(n_387) );
NAND2xp5_ASAP7_75t_L g388 ( .A(n_355), .B(n_311), .Y(n_388) );
OR2x2_ASAP7_75t_L g389 ( .A(n_345), .B(n_313), .Y(n_389) );
AOI221xp5_ASAP7_75t_L g390 ( .A1(n_334), .A2(n_339), .B1(n_353), .B2(n_350), .C(n_355), .Y(n_390) );
INVx1_ASAP7_75t_SL g391 ( .A(n_362), .Y(n_391) );
OA21x2_ASAP7_75t_L g392 ( .A1(n_338), .A2(n_303), .B(n_313), .Y(n_392) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_358), .B(n_305), .Y(n_393) );
O2A1O1Ixp33_ASAP7_75t_L g394 ( .A1(n_336), .A2(n_305), .B(n_306), .C(n_322), .Y(n_394) );
INVx1_ASAP7_75t_L g395 ( .A(n_364), .Y(n_395) );
NAND2x1p5_ASAP7_75t_L g396 ( .A(n_329), .B(n_303), .Y(n_396) );
INVx1_ASAP7_75t_SL g397 ( .A(n_362), .Y(n_397) );
AND2x2_ASAP7_75t_L g398 ( .A(n_330), .B(n_303), .Y(n_398) );
CKINVDCx5p33_ASAP7_75t_R g399 ( .A(n_324), .Y(n_399) );
AOI22xp33_ASAP7_75t_L g400 ( .A1(n_326), .A2(n_306), .B1(n_322), .B2(n_319), .Y(n_400) );
NAND2x1p5_ASAP7_75t_L g401 ( .A(n_342), .B(n_319), .Y(n_401) );
AND2x2_ASAP7_75t_L g402 ( .A(n_333), .B(n_319), .Y(n_402) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_363), .B(n_317), .Y(n_403) );
NAND2xp5_ASAP7_75t_L g404 ( .A(n_363), .B(n_25), .Y(n_404) );
INVx2_ASAP7_75t_L g405 ( .A(n_333), .Y(n_405) );
INVxp67_ASAP7_75t_L g406 ( .A(n_336), .Y(n_406) );
INVx1_ASAP7_75t_L g407 ( .A(n_368), .Y(n_407) );
OAI31xp33_ASAP7_75t_L g408 ( .A1(n_348), .A2(n_32), .A3(n_33), .B(n_34), .Y(n_408) );
INVx1_ASAP7_75t_L g409 ( .A(n_368), .Y(n_409) );
AND2x2_ASAP7_75t_L g410 ( .A(n_325), .B(n_35), .Y(n_410) );
AND2x2_ASAP7_75t_L g411 ( .A(n_325), .B(n_37), .Y(n_411) );
AOI22xp33_ASAP7_75t_L g412 ( .A1(n_342), .A2(n_215), .B1(n_205), .B2(n_42), .Y(n_412) );
AND2x2_ASAP7_75t_L g413 ( .A(n_331), .B(n_38), .Y(n_413) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_335), .B(n_40), .Y(n_414) );
AND2x2_ASAP7_75t_L g415 ( .A(n_349), .B(n_43), .Y(n_415) );
AND2x2_ASAP7_75t_L g416 ( .A(n_349), .B(n_44), .Y(n_416) );
NAND2xp5_ASAP7_75t_L g417 ( .A(n_335), .B(n_45), .Y(n_417) );
NAND2xp5_ASAP7_75t_L g418 ( .A(n_359), .B(n_46), .Y(n_418) );
NAND2xp5_ASAP7_75t_L g419 ( .A(n_375), .B(n_359), .Y(n_419) );
INVx1_ASAP7_75t_L g420 ( .A(n_380), .Y(n_420) );
NAND2xp5_ASAP7_75t_L g421 ( .A(n_375), .B(n_366), .Y(n_421) );
NOR2xp33_ASAP7_75t_L g422 ( .A(n_399), .B(n_367), .Y(n_422) );
NAND2xp5_ASAP7_75t_SL g423 ( .A(n_373), .B(n_366), .Y(n_423) );
NAND2xp5_ASAP7_75t_L g424 ( .A(n_406), .B(n_352), .Y(n_424) );
NOR2xp33_ASAP7_75t_L g425 ( .A(n_399), .B(n_367), .Y(n_425) );
INVx1_ASAP7_75t_L g426 ( .A(n_380), .Y(n_426) );
INVx1_ASAP7_75t_L g427 ( .A(n_376), .Y(n_427) );
INVx1_ASAP7_75t_L g428 ( .A(n_376), .Y(n_428) );
NOR2xp67_ASAP7_75t_L g429 ( .A(n_373), .B(n_352), .Y(n_429) );
OAI21xp5_ASAP7_75t_L g430 ( .A1(n_408), .A2(n_346), .B(n_369), .Y(n_430) );
AND2x2_ASAP7_75t_L g431 ( .A(n_370), .B(n_341), .Y(n_431) );
INVx1_ASAP7_75t_L g432 ( .A(n_395), .Y(n_432) );
INVx2_ASAP7_75t_SL g433 ( .A(n_391), .Y(n_433) );
AOI22xp5_ASAP7_75t_L g434 ( .A1(n_377), .A2(n_390), .B1(n_374), .B2(n_383), .Y(n_434) );
INVx1_ASAP7_75t_L g435 ( .A(n_395), .Y(n_435) );
NAND3xp33_ASAP7_75t_L g436 ( .A(n_385), .B(n_365), .C(n_337), .Y(n_436) );
AND2x2_ASAP7_75t_L g437 ( .A(n_402), .B(n_341), .Y(n_437) );
AND2x2_ASAP7_75t_L g438 ( .A(n_370), .B(n_365), .Y(n_438) );
AO211x2_ASAP7_75t_L g439 ( .A1(n_403), .A2(n_47), .B(n_48), .C(n_50), .Y(n_439) );
NOR2xp33_ASAP7_75t_SL g440 ( .A(n_408), .B(n_205), .Y(n_440) );
NAND2xp5_ASAP7_75t_L g441 ( .A(n_382), .B(n_52), .Y(n_441) );
INVx1_ASAP7_75t_L g442 ( .A(n_405), .Y(n_442) );
AND2x2_ASAP7_75t_L g443 ( .A(n_371), .B(n_53), .Y(n_443) );
INVx1_ASAP7_75t_L g444 ( .A(n_405), .Y(n_444) );
INVx1_ASAP7_75t_L g445 ( .A(n_407), .Y(n_445) );
NAND2xp5_ASAP7_75t_L g446 ( .A(n_382), .B(n_54), .Y(n_446) );
INVx1_ASAP7_75t_L g447 ( .A(n_407), .Y(n_447) );
INVx1_ASAP7_75t_L g448 ( .A(n_409), .Y(n_448) );
INVxp67_ASAP7_75t_L g449 ( .A(n_371), .Y(n_449) );
NAND2x1p5_ASAP7_75t_L g450 ( .A(n_391), .B(n_55), .Y(n_450) );
OR2x2_ASAP7_75t_L g451 ( .A(n_388), .B(n_57), .Y(n_451) );
INVx1_ASAP7_75t_L g452 ( .A(n_409), .Y(n_452) );
INVx2_ASAP7_75t_L g453 ( .A(n_373), .Y(n_453) );
OAI22xp5_ASAP7_75t_L g454 ( .A1(n_396), .A2(n_58), .B1(n_59), .B2(n_62), .Y(n_454) );
XOR2x2_ASAP7_75t_L g455 ( .A(n_396), .B(n_63), .Y(n_455) );
NAND2xp5_ASAP7_75t_L g456 ( .A(n_386), .B(n_64), .Y(n_456) );
NAND2xp5_ASAP7_75t_L g457 ( .A(n_386), .B(n_65), .Y(n_457) );
INVx1_ASAP7_75t_L g458 ( .A(n_398), .Y(n_458) );
BUFx6f_ASAP7_75t_L g459 ( .A(n_410), .Y(n_459) );
AOI22xp5_ASAP7_75t_L g460 ( .A1(n_372), .A2(n_66), .B1(n_67), .B2(n_68), .Y(n_460) );
A2O1A1Ixp33_ASAP7_75t_SL g461 ( .A1(n_387), .A2(n_71), .B(n_73), .C(n_417), .Y(n_461) );
INVx1_ASAP7_75t_SL g462 ( .A(n_397), .Y(n_462) );
XNOR2xp5_ASAP7_75t_L g463 ( .A(n_378), .B(n_379), .Y(n_463) );
NAND3xp33_ASAP7_75t_L g464 ( .A(n_381), .B(n_400), .C(n_389), .Y(n_464) );
CKINVDCx11_ASAP7_75t_R g465 ( .A(n_396), .Y(n_465) );
OAI21xp5_ASAP7_75t_SL g466 ( .A1(n_401), .A2(n_394), .B(n_384), .Y(n_466) );
NAND2xp5_ASAP7_75t_SL g467 ( .A(n_401), .B(n_381), .Y(n_467) );
XNOR2xp5_ASAP7_75t_L g468 ( .A(n_401), .B(n_402), .Y(n_468) );
NAND4xp25_ASAP7_75t_SL g469 ( .A(n_412), .B(n_393), .C(n_414), .D(n_418), .Y(n_469) );
AOI22xp5_ASAP7_75t_L g470 ( .A1(n_398), .A2(n_389), .B1(n_404), .B2(n_392), .Y(n_470) );
INVx2_ASAP7_75t_L g471 ( .A(n_392), .Y(n_471) );
INVx1_ASAP7_75t_SL g472 ( .A(n_416), .Y(n_472) );
AOI22xp33_ASAP7_75t_L g473 ( .A1(n_392), .A2(n_411), .B1(n_413), .B2(n_415), .Y(n_473) );
NOR3x1_ASAP7_75t_L g474 ( .A(n_392), .B(n_415), .C(n_416), .Y(n_474) );
INVx1_ASAP7_75t_SL g475 ( .A(n_371), .Y(n_475) );
INVx1_ASAP7_75t_L g476 ( .A(n_380), .Y(n_476) );
NAND2xp5_ASAP7_75t_L g477 ( .A(n_375), .B(n_406), .Y(n_477) );
NOR2xp33_ASAP7_75t_L g478 ( .A(n_399), .B(n_406), .Y(n_478) );
INVx1_ASAP7_75t_SL g479 ( .A(n_371), .Y(n_479) );
NAND2xp5_ASAP7_75t_L g480 ( .A(n_380), .B(n_382), .Y(n_480) );
XNOR2xp5_ASAP7_75t_L g481 ( .A(n_399), .B(n_226), .Y(n_481) );
AOI22xp33_ASAP7_75t_L g482 ( .A1(n_464), .A2(n_469), .B1(n_455), .B2(n_478), .Y(n_482) );
AND2x2_ASAP7_75t_L g483 ( .A(n_479), .B(n_475), .Y(n_483) );
O2A1O1Ixp33_ASAP7_75t_L g484 ( .A1(n_466), .A2(n_440), .B(n_461), .C(n_430), .Y(n_484) );
XOR2xp5_ASAP7_75t_L g485 ( .A(n_481), .B(n_455), .Y(n_485) );
OAI21xp33_ASAP7_75t_L g486 ( .A1(n_434), .A2(n_470), .B(n_477), .Y(n_486) );
AND2x2_ASAP7_75t_L g487 ( .A(n_462), .B(n_449), .Y(n_487) );
INVx1_ASAP7_75t_L g488 ( .A(n_480), .Y(n_488) );
AOI211xp5_ASAP7_75t_SL g489 ( .A1(n_422), .A2(n_425), .B(n_454), .C(n_457), .Y(n_489) );
AOI21xp5_ASAP7_75t_L g490 ( .A1(n_423), .A2(n_467), .B(n_425), .Y(n_490) );
OAI22xp5_ASAP7_75t_L g491 ( .A1(n_468), .A2(n_422), .B1(n_463), .B2(n_449), .Y(n_491) );
OAI321xp33_ASAP7_75t_L g492 ( .A1(n_450), .A2(n_423), .A3(n_436), .B1(n_419), .B2(n_473), .C(n_471), .Y(n_492) );
AOI22xp5_ASAP7_75t_L g493 ( .A1(n_465), .A2(n_421), .B1(n_437), .B2(n_458), .Y(n_493) );
INVx1_ASAP7_75t_L g494 ( .A(n_480), .Y(n_494) );
AOI22xp5_ASAP7_75t_L g495 ( .A1(n_437), .A2(n_431), .B1(n_448), .B2(n_452), .Y(n_495) );
AOI22xp5_ASAP7_75t_L g496 ( .A1(n_445), .A2(n_447), .B1(n_476), .B2(n_426), .Y(n_496) );
AOI221xp5_ASAP7_75t_L g497 ( .A1(n_420), .A2(n_424), .B1(n_428), .B2(n_427), .C(n_435), .Y(n_497) );
CKINVDCx16_ASAP7_75t_R g498 ( .A(n_485), .Y(n_498) );
NOR2xp33_ASAP7_75t_SL g499 ( .A(n_484), .B(n_450), .Y(n_499) );
OAI22xp33_ASAP7_75t_SL g500 ( .A1(n_491), .A2(n_433), .B1(n_453), .B2(n_457), .Y(n_500) );
INVx1_ASAP7_75t_L g501 ( .A(n_488), .Y(n_501) );
NOR2x1p5_ASAP7_75t_L g502 ( .A(n_487), .B(n_453), .Y(n_502) );
INVx1_ASAP7_75t_L g503 ( .A(n_494), .Y(n_503) );
AOI221xp5_ASAP7_75t_L g504 ( .A1(n_486), .A2(n_433), .B1(n_432), .B2(n_472), .C(n_444), .Y(n_504) );
AOI211x1_ASAP7_75t_SL g505 ( .A1(n_490), .A2(n_429), .B(n_456), .C(n_446), .Y(n_505) );
OAI22xp5_ASAP7_75t_L g506 ( .A1(n_482), .A2(n_459), .B1(n_438), .B2(n_451), .Y(n_506) );
INVx1_ASAP7_75t_L g507 ( .A(n_501), .Y(n_507) );
AO22x1_ASAP7_75t_L g508 ( .A1(n_506), .A2(n_474), .B1(n_489), .B2(n_483), .Y(n_508) );
NOR3xp33_ASAP7_75t_L g509 ( .A(n_498), .B(n_492), .C(n_497), .Y(n_509) );
OAI21xp33_ASAP7_75t_L g510 ( .A1(n_499), .A2(n_493), .B(n_495), .Y(n_510) );
XOR2xp5_ASAP7_75t_L g511 ( .A(n_505), .B(n_496), .Y(n_511) );
OAI211xp5_ASAP7_75t_SL g512 ( .A1(n_509), .A2(n_504), .B(n_503), .C(n_500), .Y(n_512) );
OAI22xp5_ASAP7_75t_L g513 ( .A1(n_511), .A2(n_502), .B1(n_492), .B2(n_460), .Y(n_513) );
NOR3xp33_ASAP7_75t_L g514 ( .A(n_508), .B(n_441), .C(n_443), .Y(n_514) );
XNOR2xp5_ASAP7_75t_L g515 ( .A(n_513), .B(n_507), .Y(n_515) );
NAND3xp33_ASAP7_75t_L g516 ( .A(n_514), .B(n_510), .C(n_442), .Y(n_516) );
AND2x2_ASAP7_75t_L g517 ( .A(n_515), .B(n_512), .Y(n_517) );
INVx2_ASAP7_75t_SL g518 ( .A(n_517), .Y(n_518) );
INVx1_ASAP7_75t_L g519 ( .A(n_518), .Y(n_519) );
AOI21xp5_ASAP7_75t_L g520 ( .A1(n_519), .A2(n_516), .B(n_439), .Y(n_520) );
endmodule