module fake_jpeg_24059_n_63 (n_13, n_21, n_1, n_10, n_23, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_9, n_5, n_11, n_17, n_25, n_2, n_12, n_8, n_15, n_7, n_63);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_63;

wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_27;
wire n_55;
wire n_47;
wire n_51;
wire n_40;
wire n_59;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_44;
wire n_28;
wire n_38;
wire n_26;
wire n_36;
wire n_62;
wire n_31;
wire n_56;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_32;

INVx1_ASAP7_75t_L g26 ( 
.A(n_25),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_7),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_21),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_17),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_18),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_22),
.Y(n_32)
);

INVx11_ASAP7_75t_L g33 ( 
.A(n_23),
.Y(n_33)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_33),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_34),
.B(n_32),
.Y(n_43)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_29),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_35),
.B(n_36),
.Y(n_41)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_SL g37 ( 
.A1(n_35),
.A2(n_33),
.B1(n_29),
.B2(n_0),
.Y(n_37)
);

AOI21xp5_ASAP7_75t_L g46 ( 
.A1(n_37),
.A2(n_40),
.B(n_43),
.Y(n_46)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_34),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_38),
.B(n_39),
.Y(n_48)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_34),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_34),
.B(n_0),
.Y(n_40)
);

BUFx2_ASAP7_75t_L g42 ( 
.A(n_34),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_42),
.B(n_1),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g44 ( 
.A1(n_41),
.A2(n_30),
.B1(n_31),
.B2(n_28),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g51 ( 
.A1(n_44),
.A2(n_47),
.B1(n_4),
.B2(n_5),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_45),
.B(n_46),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g47 ( 
.A1(n_40),
.A2(n_27),
.B1(n_2),
.B2(n_3),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_48),
.B(n_1),
.Y(n_49)
);

MAJIxp5_ASAP7_75t_L g54 ( 
.A(n_49),
.B(n_52),
.C(n_53),
.Y(n_54)
);

CKINVDCx14_ASAP7_75t_R g56 ( 
.A(n_50),
.Y(n_56)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_51),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_47),
.A2(n_6),
.B1(n_8),
.B2(n_9),
.Y(n_52)
);

XNOR2xp5_ASAP7_75t_L g53 ( 
.A(n_44),
.B(n_10),
.Y(n_53)
);

XNOR2xp5_ASAP7_75t_L g57 ( 
.A(n_54),
.B(n_24),
.Y(n_57)
);

AOI21xp5_ASAP7_75t_L g58 ( 
.A1(n_57),
.A2(n_55),
.B(n_56),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_58),
.B(n_11),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_59),
.B(n_12),
.Y(n_60)
);

AO21x1_ASAP7_75t_L g61 ( 
.A1(n_60),
.A2(n_13),
.B(n_14),
.Y(n_61)
);

OAI21xp5_ASAP7_75t_SL g62 ( 
.A1(n_61),
.A2(n_16),
.B(n_19),
.Y(n_62)
);

XNOR2xp5_ASAP7_75t_L g63 ( 
.A(n_62),
.B(n_20),
.Y(n_63)
);


endmodule