module fake_netlist_6_1442_n_72 (n_7, n_6, n_12, n_4, n_2, n_15, n_16, n_3, n_5, n_1, n_14, n_13, n_0, n_9, n_11, n_8, n_17, n_10, n_72);

input n_7;
input n_6;
input n_12;
input n_4;
input n_2;
input n_15;
input n_16;
input n_3;
input n_5;
input n_1;
input n_14;
input n_13;
input n_0;
input n_9;
input n_11;
input n_8;
input n_17;
input n_10;

output n_72;

wire n_41;
wire n_52;
wire n_45;
wire n_46;
wire n_34;
wire n_42;
wire n_70;
wire n_21;
wire n_18;
wire n_24;
wire n_71;
wire n_37;
wire n_54;
wire n_33;
wire n_67;
wire n_27;
wire n_38;
wire n_61;
wire n_39;
wire n_63;
wire n_60;
wire n_59;
wire n_32;
wire n_66;
wire n_36;
wire n_22;
wire n_26;
wire n_68;
wire n_55;
wire n_35;
wire n_28;
wire n_23;
wire n_58;
wire n_69;
wire n_20;
wire n_50;
wire n_49;
wire n_30;
wire n_64;
wire n_43;
wire n_48;
wire n_19;
wire n_62;
wire n_29;
wire n_47;
wire n_31;
wire n_65;
wire n_40;
wire n_25;
wire n_57;
wire n_53;
wire n_51;
wire n_44;
wire n_56;

OA21x2_ASAP7_75t_L g18 ( 
.A1(n_3),
.A2(n_12),
.B(n_16),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

BUFx8_ASAP7_75t_SL g20 ( 
.A(n_7),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_17),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_8),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_2),
.B(n_13),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_22),
.B(n_27),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_22),
.B(n_1),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_27),
.B(n_2),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_21),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_21),
.Y(n_36)
);

AOI21xp5_ASAP7_75t_L g37 ( 
.A1(n_32),
.A2(n_29),
.B(n_28),
.Y(n_37)
);

INVx2_ASAP7_75t_SL g38 ( 
.A(n_36),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g39 ( 
.A(n_33),
.B(n_21),
.Y(n_39)
);

INVxp67_ASAP7_75t_L g40 ( 
.A(n_35),
.Y(n_40)
);

NAND2xp33_ASAP7_75t_R g41 ( 
.A(n_34),
.B(n_18),
.Y(n_41)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_35),
.Y(n_42)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_39),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g44 ( 
.A1(n_37),
.A2(n_26),
.B1(n_24),
.B2(n_30),
.Y(n_44)
);

AND2x2_ASAP7_75t_L g45 ( 
.A(n_40),
.B(n_24),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_42),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_38),
.Y(n_47)
);

AND2x4_ASAP7_75t_L g48 ( 
.A(n_42),
.B(n_23),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_41),
.Y(n_49)
);

AND2x4_ASAP7_75t_SL g50 ( 
.A(n_45),
.B(n_25),
.Y(n_50)
);

AND2x2_ASAP7_75t_L g51 ( 
.A(n_48),
.B(n_19),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_L g52 ( 
.A1(n_49),
.A2(n_18),
.B1(n_30),
.B2(n_19),
.Y(n_52)
);

AND2x2_ASAP7_75t_L g53 ( 
.A(n_48),
.B(n_23),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_L g54 ( 
.A1(n_44),
.A2(n_18),
.B1(n_31),
.B2(n_21),
.Y(n_54)
);

INVxp67_ASAP7_75t_L g55 ( 
.A(n_53),
.Y(n_55)
);

BUFx2_ASAP7_75t_L g56 ( 
.A(n_51),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_52),
.B(n_54),
.Y(n_57)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_50),
.Y(n_58)
);

INVxp67_ASAP7_75t_L g59 ( 
.A(n_56),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_L g60 ( 
.A1(n_57),
.A2(n_52),
.B1(n_46),
.B2(n_43),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_55),
.B(n_43),
.Y(n_61)
);

NOR2x1_ASAP7_75t_SL g62 ( 
.A(n_60),
.B(n_58),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_59),
.B(n_55),
.Y(n_63)
);

AOI21xp5_ASAP7_75t_L g64 ( 
.A1(n_62),
.A2(n_61),
.B(n_58),
.Y(n_64)
);

OAI32xp33_ASAP7_75t_L g65 ( 
.A1(n_63),
.A2(n_47),
.A3(n_46),
.B1(n_20),
.B2(n_5),
.Y(n_65)
);

OR2x2_ASAP7_75t_L g66 ( 
.A(n_64),
.B(n_31),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_65),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_66),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_67),
.A2(n_31),
.B1(n_20),
.B2(n_5),
.Y(n_69)
);

AO22x2_ASAP7_75t_L g70 ( 
.A1(n_68),
.A2(n_69),
.B1(n_4),
.B2(n_3),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_70),
.B(n_31),
.Y(n_71)
);

OR2x6_ASAP7_75t_L g72 ( 
.A(n_71),
.B(n_15),
.Y(n_72)
);


endmodule