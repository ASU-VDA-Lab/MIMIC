module fake_jpeg_12518_n_467 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_467);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_467;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx4_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

BUFx16f_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_10),
.Y(n_22)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

BUFx16f_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_SL g26 ( 
.A(n_2),
.B(n_4),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_SL g27 ( 
.A(n_4),
.B(n_12),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_6),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_5),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_17),
.Y(n_33)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_2),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_15),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_13),
.Y(n_37)
);

INVx11_ASAP7_75t_SL g38 ( 
.A(n_1),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_14),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_0),
.Y(n_40)
);

INVx6_ASAP7_75t_SL g41 ( 
.A(n_5),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_3),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_6),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_13),
.B(n_0),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_1),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_6),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_10),
.Y(n_47)
);

INVx11_ASAP7_75t_L g48 ( 
.A(n_3),
.Y(n_48)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_9),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_0),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_8),
.Y(n_51)
);

BUFx8_ASAP7_75t_L g52 ( 
.A(n_16),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_16),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_11),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_19),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g160 ( 
.A(n_55),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_27),
.B(n_17),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_56),
.B(n_57),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g57 ( 
.A(n_27),
.B(n_17),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_58),
.B(n_59),
.Y(n_120)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_37),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_47),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_60),
.B(n_61),
.Y(n_121)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_47),
.Y(n_61)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_52),
.Y(n_62)
);

INVx3_ASAP7_75t_L g163 ( 
.A(n_62),
.Y(n_163)
);

BUFx5_ASAP7_75t_L g63 ( 
.A(n_41),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g129 ( 
.A(n_63),
.Y(n_129)
);

INVx1_ASAP7_75t_SL g64 ( 
.A(n_28),
.Y(n_64)
);

AND2x2_ASAP7_75t_L g149 ( 
.A(n_64),
.B(n_71),
.Y(n_149)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_28),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g184 ( 
.A(n_65),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_26),
.B(n_16),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_66),
.B(n_70),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_19),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g180 ( 
.A(n_67),
.Y(n_180)
);

INVx5_ASAP7_75t_SL g68 ( 
.A(n_41),
.Y(n_68)
);

CKINVDCx16_ASAP7_75t_R g140 ( 
.A(n_68),
.Y(n_140)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_19),
.Y(n_69)
);

INVx3_ASAP7_75t_SL g173 ( 
.A(n_69),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_44),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_44),
.B(n_15),
.Y(n_71)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_24),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g169 ( 
.A(n_72),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_24),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g196 ( 
.A(n_73),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_24),
.Y(n_74)
);

INVx6_ASAP7_75t_L g185 ( 
.A(n_74),
.Y(n_185)
);

BUFx12f_ASAP7_75t_L g75 ( 
.A(n_52),
.Y(n_75)
);

INVx4_ASAP7_75t_L g138 ( 
.A(n_75),
.Y(n_138)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_36),
.Y(n_76)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_76),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_48),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_77),
.B(n_83),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_22),
.B(n_53),
.Y(n_78)
);

AND2x2_ASAP7_75t_L g161 ( 
.A(n_78),
.B(n_79),
.Y(n_161)
);

INVx4_ASAP7_75t_SL g79 ( 
.A(n_48),
.Y(n_79)
);

BUFx12_ASAP7_75t_L g80 ( 
.A(n_48),
.Y(n_80)
);

BUFx4f_ASAP7_75t_SL g166 ( 
.A(n_80),
.Y(n_166)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_28),
.Y(n_81)
);

INVx4_ASAP7_75t_L g178 ( 
.A(n_81),
.Y(n_178)
);

BUFx2_ASAP7_75t_L g82 ( 
.A(n_18),
.Y(n_82)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_82),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_26),
.B(n_15),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_40),
.Y(n_84)
);

INVx8_ASAP7_75t_L g137 ( 
.A(n_84),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_22),
.B(n_53),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_85),
.B(n_86),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_39),
.B(n_14),
.Y(n_86)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_18),
.Y(n_87)
);

HB1xp67_ASAP7_75t_L g148 ( 
.A(n_87),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_40),
.Y(n_88)
);

INVx4_ASAP7_75t_L g187 ( 
.A(n_88),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_40),
.Y(n_89)
);

INVx4_ASAP7_75t_L g197 ( 
.A(n_89),
.Y(n_197)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_36),
.Y(n_90)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_90),
.Y(n_134)
);

INVx2_ASAP7_75t_SL g91 ( 
.A(n_28),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g194 ( 
.A(n_91),
.B(n_106),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_46),
.Y(n_92)
);

INVx3_ASAP7_75t_L g195 ( 
.A(n_92),
.Y(n_195)
);

INVx8_ASAP7_75t_L g93 ( 
.A(n_46),
.Y(n_93)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_93),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_39),
.B(n_12),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_94),
.B(n_95),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_39),
.B(n_12),
.Y(n_95)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_18),
.Y(n_96)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_96),
.Y(n_145)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_34),
.Y(n_97)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_97),
.Y(n_147)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_21),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_98),
.B(n_104),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_46),
.Y(n_99)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_99),
.Y(n_170)
);

BUFx12f_ASAP7_75t_L g100 ( 
.A(n_52),
.Y(n_100)
);

BUFx2_ASAP7_75t_SL g159 ( 
.A(n_100),
.Y(n_159)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_34),
.Y(n_101)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_101),
.Y(n_177)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_34),
.Y(n_102)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_102),
.Y(n_181)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_21),
.Y(n_103)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_103),
.Y(n_193)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_29),
.Y(n_104)
);

INVx11_ASAP7_75t_L g105 ( 
.A(n_38),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_105),
.Y(n_167)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_52),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_39),
.B(n_11),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_107),
.B(n_108),
.Y(n_157)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_20),
.Y(n_108)
);

INVx4_ASAP7_75t_SL g109 ( 
.A(n_32),
.Y(n_109)
);

OR2x2_ASAP7_75t_L g192 ( 
.A(n_109),
.B(n_110),
.Y(n_192)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_29),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_49),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_111),
.B(n_112),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_54),
.B(n_11),
.Y(n_112)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_45),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_113),
.B(n_115),
.Y(n_183)
);

BUFx5_ASAP7_75t_L g114 ( 
.A(n_49),
.Y(n_114)
);

NOR2x1_ASAP7_75t_L g133 ( 
.A(n_114),
.B(n_25),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_30),
.B(n_31),
.Y(n_115)
);

INVx8_ASAP7_75t_L g116 ( 
.A(n_49),
.Y(n_116)
);

AND2x4_ASAP7_75t_SL g182 ( 
.A(n_116),
.B(n_117),
.Y(n_182)
);

INVx6_ASAP7_75t_L g117 ( 
.A(n_32),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_30),
.B(n_9),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_118),
.B(n_0),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_64),
.B(n_32),
.C(n_33),
.Y(n_122)
);

AOI21xp5_ASAP7_75t_L g205 ( 
.A1(n_122),
.A2(n_146),
.B(n_151),
.Y(n_205)
);

AOI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_62),
.A2(n_23),
.B1(n_54),
.B2(n_33),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g211 ( 
.A1(n_124),
.A2(n_130),
.B1(n_131),
.B2(n_136),
.Y(n_211)
);

OAI22xp33_ASAP7_75t_L g126 ( 
.A1(n_117),
.A2(n_33),
.B1(n_54),
.B2(n_45),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_126),
.A2(n_141),
.B1(n_154),
.B2(n_179),
.Y(n_236)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_75),
.A2(n_23),
.B1(n_51),
.B2(n_50),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_75),
.A2(n_23),
.B1(n_51),
.B2(n_50),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_L g132 ( 
.A1(n_55),
.A2(n_43),
.B1(n_42),
.B2(n_35),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_132),
.A2(n_135),
.B1(n_155),
.B2(n_175),
.Y(n_230)
);

INVxp67_ASAP7_75t_L g258 ( 
.A(n_133),
.Y(n_258)
);

AOI22xp33_ASAP7_75t_L g135 ( 
.A1(n_67),
.A2(n_43),
.B1(n_42),
.B2(n_35),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_100),
.A2(n_31),
.B1(n_25),
.B2(n_20),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_73),
.A2(n_89),
.B1(n_88),
.B2(n_84),
.Y(n_141)
);

AND2x2_ASAP7_75t_SL g142 ( 
.A(n_87),
.B(n_0),
.Y(n_142)
);

AND2x2_ASAP7_75t_L g223 ( 
.A(n_142),
.B(n_162),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_91),
.B(n_25),
.C(n_20),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_100),
.A2(n_25),
.B1(n_20),
.B2(n_5),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_SL g234 ( 
.A1(n_150),
.A2(n_152),
.B1(n_156),
.B2(n_164),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_82),
.B(n_1),
.C(n_2),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_69),
.A2(n_2),
.B1(n_5),
.B2(n_7),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_111),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_L g155 ( 
.A1(n_74),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_SL g156 ( 
.A1(n_72),
.A2(n_93),
.B1(n_116),
.B2(n_65),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_92),
.B(n_99),
.C(n_68),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_SL g164 ( 
.A1(n_81),
.A2(n_105),
.B1(n_109),
.B2(n_79),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_80),
.B(n_76),
.C(n_90),
.Y(n_165)
);

AND2x2_ASAP7_75t_L g249 ( 
.A(n_165),
.B(n_168),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_80),
.B(n_76),
.C(n_90),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_SL g171 ( 
.A1(n_62),
.A2(n_18),
.B1(n_23),
.B2(n_34),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_SL g239 ( 
.A1(n_171),
.A2(n_172),
.B1(n_174),
.B2(n_176),
.Y(n_239)
);

AOI22xp33_ASAP7_75t_SL g172 ( 
.A1(n_62),
.A2(n_18),
.B1(n_23),
.B2(n_34),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_SL g174 ( 
.A1(n_62),
.A2(n_18),
.B1(n_23),
.B2(n_34),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_70),
.A2(n_117),
.B1(n_76),
.B2(n_90),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_SL g176 ( 
.A1(n_62),
.A2(n_18),
.B1(n_23),
.B2(n_34),
.Y(n_176)
);

OAI22xp33_ASAP7_75t_SL g179 ( 
.A1(n_76),
.A2(n_90),
.B1(n_36),
.B2(n_111),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_SL g186 ( 
.A1(n_62),
.A2(n_18),
.B1(n_23),
.B2(n_34),
.Y(n_186)
);

AOI22xp33_ASAP7_75t_SL g245 ( 
.A1(n_186),
.A2(n_191),
.B1(n_173),
.B2(n_163),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_188),
.B(n_184),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_70),
.A2(n_90),
.B1(n_76),
.B2(n_117),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_189),
.A2(n_190),
.B1(n_154),
.B2(n_173),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_70),
.A2(n_117),
.B1(n_76),
.B2(n_90),
.Y(n_190)
);

AOI22xp33_ASAP7_75t_SL g191 ( 
.A1(n_62),
.A2(n_18),
.B1(n_23),
.B2(n_34),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_139),
.B(n_128),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_SL g279 ( 
.A(n_198),
.B(n_213),
.Y(n_279)
);

INVx3_ASAP7_75t_L g199 ( 
.A(n_144),
.Y(n_199)
);

CKINVDCx14_ASAP7_75t_R g200 ( 
.A(n_194),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_200),
.B(n_201),
.Y(n_267)
);

CKINVDCx16_ASAP7_75t_R g201 ( 
.A(n_194),
.Y(n_201)
);

INVx1_ASAP7_75t_SL g202 ( 
.A(n_194),
.Y(n_202)
);

AND2x2_ASAP7_75t_L g282 ( 
.A(n_202),
.B(n_233),
.Y(n_282)
);

A2O1A1Ixp33_ASAP7_75t_SL g203 ( 
.A1(n_182),
.A2(n_142),
.B(n_133),
.C(n_141),
.Y(n_203)
);

OA21x2_ASAP7_75t_L g274 ( 
.A1(n_203),
.A2(n_204),
.B(n_220),
.Y(n_274)
);

OA22x2_ASAP7_75t_L g204 ( 
.A1(n_182),
.A2(n_175),
.B1(n_142),
.B2(n_193),
.Y(n_204)
);

INVx13_ASAP7_75t_L g206 ( 
.A(n_140),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_183),
.B(n_188),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_207),
.B(n_225),
.Y(n_284)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_170),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_SL g209 ( 
.A(n_119),
.B(n_127),
.Y(n_209)
);

OR2x2_ASAP7_75t_L g277 ( 
.A(n_209),
.B(n_229),
.Y(n_277)
);

INVx11_ASAP7_75t_L g210 ( 
.A(n_166),
.Y(n_210)
);

BUFx10_ASAP7_75t_L g269 ( 
.A(n_210),
.Y(n_269)
);

BUFx12_ASAP7_75t_L g212 ( 
.A(n_159),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_143),
.B(n_153),
.Y(n_213)
);

CKINVDCx11_ASAP7_75t_R g214 ( 
.A(n_140),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_214),
.B(n_215),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_120),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_121),
.B(n_157),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_SL g280 ( 
.A(n_216),
.B(n_217),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_161),
.B(n_183),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_193),
.Y(n_218)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_218),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_161),
.B(n_149),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_SL g293 ( 
.A(n_219),
.B(n_222),
.Y(n_293)
);

AO21x2_ASAP7_75t_SL g220 ( 
.A1(n_182),
.A2(n_126),
.B(n_192),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_125),
.Y(n_221)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_221),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_161),
.B(n_149),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_149),
.B(n_158),
.Y(n_224)
);

INVxp67_ASAP7_75t_L g291 ( 
.A(n_224),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_151),
.B(n_189),
.Y(n_225)
);

BUFx6f_ASAP7_75t_L g226 ( 
.A(n_160),
.Y(n_226)
);

BUFx6f_ASAP7_75t_L g278 ( 
.A(n_226),
.Y(n_278)
);

CKINVDCx16_ASAP7_75t_R g227 ( 
.A(n_148),
.Y(n_227)
);

INVxp33_ASAP7_75t_L g264 ( 
.A(n_227),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_165),
.B(n_168),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_228),
.B(n_248),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_SL g229 ( 
.A(n_129),
.B(n_167),
.Y(n_229)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_170),
.Y(n_231)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_231),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_192),
.B(n_167),
.Y(n_232)
);

INVxp67_ASAP7_75t_L g297 ( 
.A(n_232),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_123),
.B(n_134),
.Y(n_233)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_123),
.Y(n_235)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_235),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_SL g237 ( 
.A(n_190),
.B(n_138),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_237),
.A2(n_245),
.B1(n_202),
.B2(n_239),
.Y(n_283)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_145),
.Y(n_238)
);

AND2x2_ASAP7_75t_L g287 ( 
.A(n_238),
.B(n_242),
.Y(n_287)
);

INVx4_ASAP7_75t_L g240 ( 
.A(n_138),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_L g299 ( 
.A1(n_241),
.A2(n_251),
.B1(n_236),
.B2(n_220),
.Y(n_299)
);

OA22x2_ASAP7_75t_L g242 ( 
.A1(n_162),
.A2(n_134),
.B1(n_195),
.B2(n_177),
.Y(n_242)
);

NAND2x1p5_ASAP7_75t_L g243 ( 
.A(n_146),
.B(n_122),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_L g265 ( 
.A1(n_243),
.A2(n_205),
.B(n_228),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_SL g244 ( 
.A(n_129),
.B(n_166),
.Y(n_244)
);

NOR3xp33_ASAP7_75t_SL g300 ( 
.A(n_244),
.B(n_262),
.C(n_263),
.Y(n_300)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_195),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_163),
.B(n_177),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_247),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_147),
.B(n_181),
.Y(n_248)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_145),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_250),
.B(n_252),
.Y(n_292)
);

AOI22xp33_ASAP7_75t_L g251 ( 
.A1(n_187),
.A2(n_197),
.B1(n_137),
.B2(n_185),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_147),
.B(n_181),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_144),
.B(n_137),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_253),
.B(n_256),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_185),
.A2(n_197),
.B1(n_187),
.B2(n_196),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_254),
.A2(n_259),
.B1(n_256),
.B2(n_220),
.Y(n_275)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_178),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_173),
.Y(n_256)
);

OA22x2_ASAP7_75t_L g257 ( 
.A1(n_169),
.A2(n_196),
.B1(n_180),
.B2(n_160),
.Y(n_257)
);

AND2x2_ASAP7_75t_SL g268 ( 
.A(n_257),
.B(n_259),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_196),
.A2(n_180),
.B1(n_169),
.B2(n_178),
.Y(n_259)
);

BUFx5_ASAP7_75t_L g260 ( 
.A(n_169),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_184),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_261),
.B(n_262),
.Y(n_295)
);

BUFx24_ASAP7_75t_L g262 ( 
.A(n_166),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_265),
.B(n_281),
.C(n_266),
.Y(n_330)
);

AOI21xp5_ASAP7_75t_L g266 ( 
.A1(n_243),
.A2(n_223),
.B(n_258),
.Y(n_266)
);

AOI21xp5_ASAP7_75t_L g312 ( 
.A1(n_266),
.A2(n_270),
.B(n_290),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_268),
.A2(n_299),
.B1(n_257),
.B2(n_246),
.Y(n_317)
);

OAI21xp5_ASAP7_75t_SL g270 ( 
.A1(n_223),
.A2(n_225),
.B(n_205),
.Y(n_270)
);

AND2x6_ASAP7_75t_L g272 ( 
.A(n_243),
.B(n_258),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_SL g309 ( 
.A(n_272),
.B(n_296),
.Y(n_309)
);

AOI22xp33_ASAP7_75t_L g321 ( 
.A1(n_275),
.A2(n_231),
.B1(n_226),
.B2(n_255),
.Y(n_321)
);

AND2x2_ASAP7_75t_SL g281 ( 
.A(n_204),
.B(n_223),
.Y(n_281)
);

OAI21xp5_ASAP7_75t_SL g336 ( 
.A1(n_283),
.A2(n_267),
.B(n_274),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_230),
.A2(n_237),
.B1(n_220),
.B2(n_203),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_L g318 ( 
.A1(n_289),
.A2(n_235),
.B1(n_199),
.B2(n_208),
.Y(n_318)
);

OAI21xp5_ASAP7_75t_SL g290 ( 
.A1(n_249),
.A2(n_241),
.B(n_204),
.Y(n_290)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_295),
.Y(n_310)
);

AND2x6_ASAP7_75t_L g296 ( 
.A(n_249),
.B(n_203),
.Y(n_296)
);

OAI21xp5_ASAP7_75t_SL g301 ( 
.A1(n_249),
.A2(n_204),
.B(n_203),
.Y(n_301)
);

OR2x2_ASAP7_75t_L g313 ( 
.A(n_301),
.B(n_218),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_207),
.B(n_242),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_302),
.B(n_303),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_242),
.B(n_253),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_280),
.B(n_215),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_SL g355 ( 
.A(n_304),
.B(n_315),
.Y(n_355)
);

XOR2xp5_ASAP7_75t_L g305 ( 
.A(n_265),
.B(n_242),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g363 ( 
.A(n_305),
.B(n_298),
.C(n_288),
.Y(n_363)
);

OAI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_289),
.A2(n_303),
.B1(n_284),
.B2(n_302),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_306),
.B(n_308),
.Y(n_341)
);

AOI22xp33_ASAP7_75t_SL g307 ( 
.A1(n_275),
.A2(n_211),
.B1(n_234),
.B2(n_262),
.Y(n_307)
);

INVxp67_ASAP7_75t_L g349 ( 
.A(n_307),
.Y(n_349)
);

OAI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_284),
.A2(n_236),
.B1(n_254),
.B2(n_257),
.Y(n_308)
);

AOI22xp33_ASAP7_75t_SL g311 ( 
.A1(n_283),
.A2(n_210),
.B1(n_261),
.B2(n_257),
.Y(n_311)
);

INVxp67_ASAP7_75t_L g351 ( 
.A(n_311),
.Y(n_351)
);

OAI21xp5_ASAP7_75t_SL g361 ( 
.A1(n_313),
.A2(n_336),
.B(n_339),
.Y(n_361)
);

OAI21xp5_ASAP7_75t_L g314 ( 
.A1(n_281),
.A2(n_301),
.B(n_290),
.Y(n_314)
);

INVxp67_ASAP7_75t_L g353 ( 
.A(n_314),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_280),
.B(n_250),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_279),
.B(n_238),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_SL g356 ( 
.A(n_316),
.B(n_324),
.Y(n_356)
);

OAI22xp5_ASAP7_75t_L g360 ( 
.A1(n_317),
.A2(n_321),
.B1(n_325),
.B2(n_334),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_318),
.B(n_326),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_SL g320 ( 
.A(n_286),
.B(n_221),
.Y(n_320)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_273),
.Y(n_322)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_322),
.Y(n_340)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_273),
.Y(n_323)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_323),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_SL g324 ( 
.A(n_297),
.B(n_206),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_L g325 ( 
.A1(n_287),
.A2(n_240),
.B1(n_260),
.B2(n_212),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_276),
.B(n_277),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_276),
.B(n_277),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_327),
.B(n_328),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_286),
.B(n_294),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_271),
.B(n_297),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_329),
.B(n_331),
.Y(n_345)
);

XNOR2xp5_ASAP7_75t_L g343 ( 
.A(n_330),
.B(n_282),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_295),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_294),
.B(n_270),
.Y(n_332)
);

A2O1A1O1Ixp25_ASAP7_75t_L g348 ( 
.A1(n_332),
.A2(n_335),
.B(n_272),
.C(n_296),
.D(n_282),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_264),
.B(n_292),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g350 ( 
.A(n_333),
.B(n_338),
.Y(n_350)
);

AOI22xp5_ASAP7_75t_L g334 ( 
.A1(n_287),
.A2(n_268),
.B1(n_274),
.B2(n_281),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_292),
.B(n_287),
.Y(n_335)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_285),
.Y(n_337)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_337),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_SL g338 ( 
.A(n_291),
.B(n_293),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_293),
.B(n_291),
.Y(n_339)
);

XOR2xp5_ASAP7_75t_L g342 ( 
.A(n_330),
.B(n_274),
.Y(n_342)
);

XNOR2xp5_ASAP7_75t_L g378 ( 
.A(n_342),
.B(n_343),
.Y(n_378)
);

CKINVDCx16_ASAP7_75t_R g346 ( 
.A(n_329),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_SL g372 ( 
.A(n_346),
.B(n_347),
.Y(n_372)
);

XNOR2xp5_ASAP7_75t_L g347 ( 
.A(n_330),
.B(n_282),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_SL g389 ( 
.A(n_348),
.B(n_362),
.Y(n_389)
);

CKINVDCx20_ASAP7_75t_R g357 ( 
.A(n_326),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_L g373 ( 
.A(n_357),
.B(n_364),
.Y(n_373)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_322),
.Y(n_359)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_359),
.Y(n_370)
);

NOR3xp33_ASAP7_75t_SL g362 ( 
.A(n_332),
.B(n_300),
.C(n_269),
.Y(n_362)
);

OAI21xp5_ASAP7_75t_SL g381 ( 
.A1(n_363),
.A2(n_312),
.B(n_313),
.Y(n_381)
);

CKINVDCx20_ASAP7_75t_R g364 ( 
.A(n_327),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_323),
.Y(n_365)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_365),
.Y(n_375)
);

BUFx10_ASAP7_75t_L g366 ( 
.A(n_311),
.Y(n_366)
);

HB1xp67_ASAP7_75t_L g382 ( 
.A(n_366),
.Y(n_382)
);

OAI22xp5_ASAP7_75t_L g367 ( 
.A1(n_317),
.A2(n_268),
.B1(n_300),
.B2(n_278),
.Y(n_367)
);

AOI22xp5_ASAP7_75t_L g377 ( 
.A1(n_367),
.A2(n_351),
.B1(n_360),
.B2(n_305),
.Y(n_377)
);

OAI22xp5_ASAP7_75t_SL g368 ( 
.A1(n_341),
.A2(n_334),
.B1(n_319),
.B2(n_307),
.Y(n_368)
);

AOI22xp5_ASAP7_75t_L g396 ( 
.A1(n_368),
.A2(n_383),
.B1(n_306),
.B2(n_305),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_SL g369 ( 
.A(n_357),
.B(n_331),
.Y(n_369)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_369),
.Y(n_397)
);

NOR2xp33_ASAP7_75t_SL g371 ( 
.A(n_364),
.B(n_339),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_SL g408 ( 
.A(n_371),
.B(n_304),
.Y(n_408)
);

CKINVDCx20_ASAP7_75t_R g374 ( 
.A(n_345),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_374),
.B(n_386),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_352),
.B(n_310),
.Y(n_376)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_376),
.Y(n_395)
);

OAI22xp5_ASAP7_75t_L g410 ( 
.A1(n_377),
.A2(n_380),
.B1(n_390),
.B2(n_313),
.Y(n_410)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_340),
.Y(n_379)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_379),
.Y(n_404)
);

CKINVDCx14_ASAP7_75t_R g380 ( 
.A(n_356),
.Y(n_380)
);

XOR2xp5_ASAP7_75t_L g392 ( 
.A(n_381),
.B(n_342),
.Y(n_392)
);

OAI22xp5_ASAP7_75t_SL g383 ( 
.A1(n_341),
.A2(n_334),
.B1(n_319),
.B2(n_317),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_340),
.Y(n_384)
);

INVx1_ASAP7_75t_SL g401 ( 
.A(n_384),
.Y(n_401)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_354),
.Y(n_385)
);

INVxp67_ASAP7_75t_L g393 ( 
.A(n_385),
.Y(n_393)
);

CKINVDCx20_ASAP7_75t_R g386 ( 
.A(n_350),
.Y(n_386)
);

AOI21xp5_ASAP7_75t_L g387 ( 
.A1(n_353),
.A2(n_336),
.B(n_314),
.Y(n_387)
);

INVxp67_ASAP7_75t_L g402 ( 
.A(n_387),
.Y(n_402)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_354),
.Y(n_388)
);

INVxp67_ASAP7_75t_L g406 ( 
.A(n_388),
.Y(n_406)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_358),
.Y(n_390)
);

HB1xp67_ASAP7_75t_L g391 ( 
.A(n_344),
.Y(n_391)
);

INVxp33_ASAP7_75t_L g409 ( 
.A(n_391),
.Y(n_409)
);

XOR2xp5_ASAP7_75t_L g425 ( 
.A(n_392),
.B(n_403),
.Y(n_425)
);

OAI22xp5_ASAP7_75t_SL g416 ( 
.A1(n_396),
.A2(n_400),
.B1(n_407),
.B2(n_411),
.Y(n_416)
);

MAJIxp5_ASAP7_75t_L g398 ( 
.A(n_378),
.B(n_363),
.C(n_343),
.Y(n_398)
);

MAJIxp5_ASAP7_75t_L g412 ( 
.A(n_398),
.B(n_405),
.C(n_361),
.Y(n_412)
);

OAI22xp5_ASAP7_75t_SL g399 ( 
.A1(n_377),
.A2(n_351),
.B1(n_366),
.B2(n_349),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_399),
.B(n_410),
.Y(n_423)
);

AOI22xp5_ASAP7_75t_L g400 ( 
.A1(n_368),
.A2(n_366),
.B1(n_349),
.B2(n_344),
.Y(n_400)
);

XNOR2xp5_ASAP7_75t_L g403 ( 
.A(n_378),
.B(n_372),
.Y(n_403)
);

MAJIxp5_ASAP7_75t_L g405 ( 
.A(n_381),
.B(n_347),
.C(n_312),
.Y(n_405)
);

AOI22xp5_ASAP7_75t_L g407 ( 
.A1(n_383),
.A2(n_366),
.B1(n_308),
.B2(n_353),
.Y(n_407)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_408),
.Y(n_424)
);

OAI22xp5_ASAP7_75t_SL g411 ( 
.A1(n_387),
.A2(n_314),
.B1(n_352),
.B2(n_309),
.Y(n_411)
);

XNOR2xp5_ASAP7_75t_L g430 ( 
.A(n_412),
.B(n_417),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_SL g413 ( 
.A(n_394),
.B(n_374),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_413),
.B(n_414),
.Y(n_432)
);

NOR2xp33_ASAP7_75t_L g414 ( 
.A(n_394),
.B(n_355),
.Y(n_414)
);

CKINVDCx20_ASAP7_75t_R g415 ( 
.A(n_401),
.Y(n_415)
);

AOI22xp5_ASAP7_75t_L g427 ( 
.A1(n_415),
.A2(n_421),
.B1(n_409),
.B2(n_395),
.Y(n_427)
);

NOR2xp33_ASAP7_75t_L g417 ( 
.A(n_397),
.B(n_355),
.Y(n_417)
);

AND2x2_ASAP7_75t_L g418 ( 
.A(n_399),
.B(n_382),
.Y(n_418)
);

NOR2xp67_ASAP7_75t_SL g436 ( 
.A(n_418),
.B(n_356),
.Y(n_436)
);

MAJIxp5_ASAP7_75t_L g419 ( 
.A(n_398),
.B(n_328),
.C(n_361),
.Y(n_419)
);

MAJIxp5_ASAP7_75t_L g434 ( 
.A(n_419),
.B(n_420),
.C(n_426),
.Y(n_434)
);

MAJIxp5_ASAP7_75t_L g420 ( 
.A(n_392),
.B(n_389),
.C(n_320),
.Y(n_420)
);

OAI22xp5_ASAP7_75t_SL g421 ( 
.A1(n_407),
.A2(n_400),
.B1(n_396),
.B2(n_395),
.Y(n_421)
);

XNOR2xp5_ASAP7_75t_L g422 ( 
.A(n_403),
.B(n_411),
.Y(n_422)
);

XOR2xp5_ASAP7_75t_L g428 ( 
.A(n_422),
.B(n_373),
.Y(n_428)
);

MAJIxp5_ASAP7_75t_L g426 ( 
.A(n_405),
.B(n_369),
.C(n_376),
.Y(n_426)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_427),
.Y(n_443)
);

XNOR2xp5_ASAP7_75t_L g439 ( 
.A(n_428),
.B(n_429),
.Y(n_439)
);

XOR2xp5_ASAP7_75t_L g429 ( 
.A(n_425),
.B(n_402),
.Y(n_429)
);

OAI21xp5_ASAP7_75t_L g431 ( 
.A1(n_426),
.A2(n_348),
.B(n_402),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_431),
.B(n_435),
.Y(n_445)
);

XOR2xp5_ASAP7_75t_L g433 ( 
.A(n_425),
.B(n_309),
.Y(n_433)
);

AND2x2_ASAP7_75t_L g446 ( 
.A(n_433),
.B(n_420),
.Y(n_446)
);

OR2x2_ASAP7_75t_L g435 ( 
.A(n_424),
.B(n_371),
.Y(n_435)
);

INVxp67_ASAP7_75t_L g441 ( 
.A(n_436),
.Y(n_441)
);

AOI22xp5_ASAP7_75t_L g437 ( 
.A1(n_421),
.A2(n_386),
.B1(n_401),
.B2(n_318),
.Y(n_437)
);

NOR2xp33_ASAP7_75t_L g444 ( 
.A(n_437),
.B(n_416),
.Y(n_444)
);

MAJIxp5_ASAP7_75t_L g438 ( 
.A(n_412),
.B(n_406),
.C(n_393),
.Y(n_438)
);

MAJIxp5_ASAP7_75t_L g440 ( 
.A(n_438),
.B(n_429),
.C(n_434),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_L g450 ( 
.A(n_440),
.B(n_447),
.Y(n_450)
);

A2O1A1Ixp33_ASAP7_75t_SL g442 ( 
.A1(n_433),
.A2(n_416),
.B(n_418),
.C(n_423),
.Y(n_442)
);

OAI21xp5_ASAP7_75t_SL g448 ( 
.A1(n_442),
.A2(n_418),
.B(n_438),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_444),
.Y(n_449)
);

XNOR2xp5_ASAP7_75t_L g454 ( 
.A(n_446),
.B(n_434),
.Y(n_454)
);

NOR2xp33_ASAP7_75t_SL g447 ( 
.A(n_432),
.B(n_316),
.Y(n_447)
);

AOI21xp5_ASAP7_75t_L g457 ( 
.A1(n_448),
.A2(n_444),
.B(n_422),
.Y(n_457)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_443),
.Y(n_451)
);

NOR2xp33_ASAP7_75t_L g459 ( 
.A(n_451),
.B(n_452),
.Y(n_459)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_441),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_445),
.Y(n_453)
);

OR2x2_ASAP7_75t_L g456 ( 
.A(n_453),
.B(n_454),
.Y(n_456)
);

MAJIxp5_ASAP7_75t_L g455 ( 
.A(n_454),
.B(n_430),
.C(n_442),
.Y(n_455)
);

AOI21xp5_ASAP7_75t_L g461 ( 
.A1(n_455),
.A2(n_457),
.B(n_458),
.Y(n_461)
);

AOI21xp5_ASAP7_75t_SL g458 ( 
.A1(n_450),
.A2(n_435),
.B(n_419),
.Y(n_458)
);

AOI322xp5_ASAP7_75t_L g460 ( 
.A1(n_459),
.A2(n_449),
.A3(n_448),
.B1(n_393),
.B2(n_406),
.C1(n_442),
.C2(n_404),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_460),
.B(n_462),
.Y(n_464)
);

AOI322xp5_ASAP7_75t_L g462 ( 
.A1(n_456),
.A2(n_384),
.A3(n_370),
.B1(n_390),
.B2(n_388),
.C1(n_385),
.C2(n_375),
.Y(n_462)
);

INVxp67_ASAP7_75t_L g463 ( 
.A(n_461),
.Y(n_463)
);

MAJIxp5_ASAP7_75t_L g465 ( 
.A(n_463),
.B(n_464),
.C(n_428),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_465),
.Y(n_466)
);

XOR2xp5_ASAP7_75t_L g467 ( 
.A(n_466),
.B(n_439),
.Y(n_467)
);


endmodule