module fake_netlist_5_180_n_541 (n_91, n_82, n_10, n_24, n_86, n_83, n_61, n_90, n_75, n_65, n_78, n_74, n_57, n_96, n_37, n_31, n_13, n_66, n_60, n_16, n_43, n_0, n_58, n_9, n_69, n_18, n_42, n_22, n_1, n_45, n_46, n_21, n_94, n_38, n_80, n_4, n_35, n_73, n_17, n_92, n_19, n_30, n_5, n_33, n_14, n_84, n_23, n_29, n_79, n_47, n_25, n_53, n_8, n_44, n_40, n_34, n_62, n_71, n_85, n_95, n_59, n_26, n_55, n_2, n_3, n_49, n_20, n_6, n_39, n_54, n_12, n_67, n_36, n_76, n_87, n_27, n_64, n_77, n_81, n_28, n_89, n_70, n_68, n_93, n_72, n_32, n_41, n_56, n_51, n_63, n_11, n_7, n_15, n_48, n_50, n_52, n_88, n_541);

input n_91;
input n_82;
input n_10;
input n_24;
input n_86;
input n_83;
input n_61;
input n_90;
input n_75;
input n_65;
input n_78;
input n_74;
input n_57;
input n_96;
input n_37;
input n_31;
input n_13;
input n_66;
input n_60;
input n_16;
input n_43;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_42;
input n_22;
input n_1;
input n_45;
input n_46;
input n_21;
input n_94;
input n_38;
input n_80;
input n_4;
input n_35;
input n_73;
input n_17;
input n_92;
input n_19;
input n_30;
input n_5;
input n_33;
input n_14;
input n_84;
input n_23;
input n_29;
input n_79;
input n_47;
input n_25;
input n_53;
input n_8;
input n_44;
input n_40;
input n_34;
input n_62;
input n_71;
input n_85;
input n_95;
input n_59;
input n_26;
input n_55;
input n_2;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_12;
input n_67;
input n_36;
input n_76;
input n_87;
input n_27;
input n_64;
input n_77;
input n_81;
input n_28;
input n_89;
input n_70;
input n_68;
input n_93;
input n_72;
input n_32;
input n_41;
input n_56;
input n_51;
input n_63;
input n_11;
input n_7;
input n_15;
input n_48;
input n_50;
input n_52;
input n_88;

output n_541;

wire n_137;
wire n_294;
wire n_431;
wire n_318;
wire n_380;
wire n_419;
wire n_444;
wire n_469;
wire n_194;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_136;
wire n_146;
wire n_124;
wire n_315;
wire n_268;
wire n_523;
wire n_451;
wire n_532;
wire n_408;
wire n_376;
wire n_503;
wire n_127;
wire n_235;
wire n_226;
wire n_515;
wire n_353;
wire n_351;
wire n_367;
wire n_452;
wire n_397;
wire n_493;
wire n_111;
wire n_525;
wire n_483;
wire n_155;
wire n_116;
wire n_467;
wire n_423;
wire n_284;
wire n_245;
wire n_501;
wire n_139;
wire n_105;
wire n_280;
wire n_378;
wire n_382;
wire n_254;
wire n_302;
wire n_265;
wire n_526;
wire n_293;
wire n_372;
wire n_443;
wire n_244;
wire n_173;
wire n_198;
wire n_447;
wire n_247;
wire n_314;
wire n_368;
wire n_433;
wire n_321;
wire n_292;
wire n_100;
wire n_455;
wire n_417;
wire n_212;
wire n_385;
wire n_498;
wire n_516;
wire n_507;
wire n_119;
wire n_497;
wire n_275;
wire n_252;
wire n_295;
wire n_133;
wire n_330;
wire n_508;
wire n_506;
wire n_509;
wire n_147;
wire n_373;
wire n_307;
wire n_439;
wire n_150;
wire n_530;
wire n_106;
wire n_209;
wire n_259;
wire n_448;
wire n_375;
wire n_301;
wire n_186;
wire n_537;
wire n_134;
wire n_191;
wire n_492;
wire n_171;
wire n_153;
wire n_524;
wire n_399;
wire n_341;
wire n_204;
wire n_394;
wire n_250;
wire n_260;
wire n_298;
wire n_320;
wire n_518;
wire n_505;
wire n_286;
wire n_122;
wire n_282;
wire n_331;
wire n_406;
wire n_519;
wire n_470;
wire n_325;
wire n_449;
wire n_132;
wire n_101;
wire n_281;
wire n_240;
wire n_381;
wire n_189;
wire n_220;
wire n_291;
wire n_231;
wire n_257;
wire n_390;
wire n_456;
wire n_371;
wire n_481;
wire n_535;
wire n_152;
wire n_540;
wire n_317;
wire n_323;
wire n_195;
wire n_356;
wire n_227;
wire n_271;
wire n_335;
wire n_123;
wire n_370;
wire n_167;
wire n_234;
wire n_343;
wire n_308;
wire n_379;
wire n_428;
wire n_267;
wire n_514;
wire n_457;
wire n_297;
wire n_156;
wire n_225;
wire n_377;
wire n_484;
wire n_219;
wire n_442;
wire n_157;
wire n_131;
wire n_192;
wire n_223;
wire n_392;
wire n_158;
wire n_138;
wire n_264;
wire n_109;
wire n_472;
wire n_454;
wire n_387;
wire n_374;
wire n_163;
wire n_276;
wire n_339;
wire n_183;
wire n_185;
wire n_243;
wire n_398;
wire n_396;
wire n_347;
wire n_169;
wire n_522;
wire n_255;
wire n_215;
wire n_350;
wire n_196;
wire n_459;
wire n_211;
wire n_218;
wire n_400;
wire n_181;
wire n_436;
wire n_290;
wire n_221;
wire n_178;
wire n_386;
wire n_287;
wire n_344;
wire n_473;
wire n_422;
wire n_475;
wire n_104;
wire n_415;
wire n_141;
wire n_485;
wire n_496;
wire n_355;
wire n_486;
wire n_336;
wire n_145;
wire n_521;
wire n_337;
wire n_430;
wire n_313;
wire n_528;
wire n_479;
wire n_510;
wire n_216;
wire n_168;
wire n_395;
wire n_164;
wire n_432;
wire n_311;
wire n_208;
wire n_142;
wire n_214;
wire n_328;
wire n_140;
wire n_299;
wire n_303;
wire n_369;
wire n_296;
wire n_241;
wire n_357;
wire n_184;
wire n_446;
wire n_445;
wire n_144;
wire n_114;
wire n_165;
wire n_468;
wire n_499;
wire n_213;
wire n_129;
wire n_342;
wire n_482;
wire n_517;
wire n_98;
wire n_361;
wire n_464;
wire n_363;
wire n_413;
wire n_402;
wire n_197;
wire n_107;
wire n_236;
wire n_388;
wire n_249;
wire n_304;
wire n_329;
wire n_203;
wire n_274;
wire n_384;
wire n_460;
wire n_277;
wire n_338;
wire n_149;
wire n_477;
wire n_461;
wire n_333;
wire n_309;
wire n_512;
wire n_462;
wire n_130;
wire n_322;
wire n_258;
wire n_151;
wire n_306;
wire n_458;
wire n_288;
wire n_188;
wire n_190;
wire n_201;
wire n_263;
wire n_471;
wire n_224;
wire n_228;
wire n_283;
wire n_383;
wire n_474;
wire n_112;
wire n_488;
wire n_463;
wire n_502;
wire n_239;
wire n_466;
wire n_420;
wire n_489;
wire n_310;
wire n_504;
wire n_511;
wire n_465;
wire n_358;
wire n_362;
wire n_170;
wire n_332;
wire n_102;
wire n_161;
wire n_273;
wire n_349;
wire n_270;
wire n_230;
wire n_118;
wire n_279;
wire n_253;
wire n_261;
wire n_174;
wire n_289;
wire n_206;
wire n_172;
wire n_217;
wire n_440;
wire n_478;
wire n_441;
wire n_450;
wire n_312;
wire n_476;
wire n_429;
wire n_534;
wire n_345;
wire n_210;
wire n_494;
wire n_365;
wire n_176;
wire n_182;
wire n_143;
wire n_354;
wire n_480;
wire n_237;
wire n_425;
wire n_513;
wire n_407;
wire n_527;
wire n_180;
wire n_340;
wire n_207;
wire n_346;
wire n_393;
wire n_229;
wire n_108;
wire n_495;
wire n_487;
wire n_437;
wire n_177;
wire n_403;
wire n_453;
wire n_421;
wire n_405;
wire n_359;
wire n_490;
wire n_117;
wire n_326;
wire n_233;
wire n_404;
wire n_205;
wire n_366;
wire n_113;
wire n_246;
wire n_179;
wire n_125;
wire n_410;
wire n_269;
wire n_529;
wire n_128;
wire n_285;
wire n_412;
wire n_120;
wire n_232;
wire n_327;
wire n_135;
wire n_126;
wire n_202;
wire n_266;
wire n_272;
wire n_491;
wire n_427;
wire n_193;
wire n_251;
wire n_352;
wire n_160;
wire n_426;
wire n_520;
wire n_409;
wire n_500;
wire n_154;
wire n_148;
wire n_300;
wire n_435;
wire n_159;
wire n_334;
wire n_391;
wire n_434;
wire n_539;
wire n_175;
wire n_538;
wire n_262;
wire n_238;
wire n_99;
wire n_411;
wire n_414;
wire n_319;
wire n_364;
wire n_536;
wire n_531;
wire n_121;
wire n_242;
wire n_360;
wire n_200;
wire n_162;
wire n_222;
wire n_438;
wire n_115;
wire n_324;
wire n_416;
wire n_199;
wire n_187;
wire n_401;
wire n_103;
wire n_348;
wire n_97;
wire n_166;
wire n_424;
wire n_256;
wire n_305;
wire n_533;
wire n_278;
wire n_110;

CKINVDCx14_ASAP7_75t_R g97 ( 
.A(n_89),
.Y(n_97)
);

CKINVDCx5p33_ASAP7_75t_R g98 ( 
.A(n_18),
.Y(n_98)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_31),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_49),
.Y(n_100)
);

CKINVDCx5p33_ASAP7_75t_R g101 ( 
.A(n_76),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_36),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_88),
.Y(n_103)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_67),
.Y(n_104)
);

CKINVDCx5p33_ASAP7_75t_R g105 ( 
.A(n_21),
.Y(n_105)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_71),
.Y(n_106)
);

CKINVDCx5p33_ASAP7_75t_R g107 ( 
.A(n_43),
.Y(n_107)
);

CKINVDCx5p33_ASAP7_75t_R g108 ( 
.A(n_87),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_20),
.Y(n_109)
);

INVx1_ASAP7_75t_SL g110 ( 
.A(n_34),
.Y(n_110)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_14),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_51),
.Y(n_112)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_46),
.Y(n_113)
);

BUFx10_ASAP7_75t_L g114 ( 
.A(n_26),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_95),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_1),
.Y(n_116)
);

INVx1_ASAP7_75t_SL g117 ( 
.A(n_13),
.Y(n_117)
);

BUFx3_ASAP7_75t_L g118 ( 
.A(n_60),
.Y(n_118)
);

CKINVDCx5p33_ASAP7_75t_R g119 ( 
.A(n_81),
.Y(n_119)
);

CKINVDCx5p33_ASAP7_75t_R g120 ( 
.A(n_29),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_55),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_64),
.Y(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_8),
.Y(n_123)
);

CKINVDCx5p33_ASAP7_75t_R g124 ( 
.A(n_73),
.Y(n_124)
);

CKINVDCx5p33_ASAP7_75t_R g125 ( 
.A(n_75),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_23),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_91),
.Y(n_127)
);

CKINVDCx5p33_ASAP7_75t_R g128 ( 
.A(n_2),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_53),
.Y(n_129)
);

CKINVDCx5p33_ASAP7_75t_R g130 ( 
.A(n_32),
.Y(n_130)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_40),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_72),
.Y(n_132)
);

CKINVDCx5p33_ASAP7_75t_R g133 ( 
.A(n_1),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_86),
.Y(n_134)
);

NOR2xp67_ASAP7_75t_L g135 ( 
.A(n_47),
.B(n_54),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_62),
.Y(n_136)
);

INVxp67_ASAP7_75t_SL g137 ( 
.A(n_11),
.Y(n_137)
);

CKINVDCx5p33_ASAP7_75t_R g138 ( 
.A(n_24),
.Y(n_138)
);

CKINVDCx5p33_ASAP7_75t_R g139 ( 
.A(n_37),
.Y(n_139)
);

CKINVDCx5p33_ASAP7_75t_R g140 ( 
.A(n_58),
.Y(n_140)
);

CKINVDCx5p33_ASAP7_75t_R g141 ( 
.A(n_84),
.Y(n_141)
);

CKINVDCx5p33_ASAP7_75t_R g142 ( 
.A(n_83),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_50),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_90),
.Y(n_144)
);

CKINVDCx5p33_ASAP7_75t_R g145 ( 
.A(n_44),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_69),
.Y(n_146)
);

CKINVDCx5p33_ASAP7_75t_R g147 ( 
.A(n_27),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_48),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_9),
.Y(n_149)
);

CKINVDCx16_ASAP7_75t_R g150 ( 
.A(n_3),
.Y(n_150)
);

CKINVDCx5p33_ASAP7_75t_R g151 ( 
.A(n_79),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_2),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_8),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_61),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_19),
.Y(n_155)
);

BUFx3_ASAP7_75t_L g156 ( 
.A(n_15),
.Y(n_156)
);

NOR2xp67_ASAP7_75t_L g157 ( 
.A(n_25),
.B(n_59),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_15),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_35),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_10),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_80),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_92),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_22),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_33),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_78),
.Y(n_165)
);

CKINVDCx16_ASAP7_75t_R g166 ( 
.A(n_10),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_16),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_38),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_5),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_7),
.Y(n_170)
);

HB1xp67_ASAP7_75t_L g171 ( 
.A(n_41),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_82),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_12),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_45),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_16),
.Y(n_175)
);

BUFx10_ASAP7_75t_L g176 ( 
.A(n_57),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_74),
.Y(n_177)
);

BUFx2_ASAP7_75t_L g178 ( 
.A(n_14),
.Y(n_178)
);

INVxp67_ASAP7_75t_SL g179 ( 
.A(n_96),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_63),
.Y(n_180)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_30),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_6),
.Y(n_182)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_6),
.Y(n_183)
);

BUFx5_ASAP7_75t_L g184 ( 
.A(n_5),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g185 ( 
.A(n_70),
.Y(n_185)
);

HB1xp67_ASAP7_75t_L g186 ( 
.A(n_93),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_94),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_3),
.Y(n_188)
);

INVx1_ASAP7_75t_SL g189 ( 
.A(n_12),
.Y(n_189)
);

BUFx2_ASAP7_75t_L g190 ( 
.A(n_13),
.Y(n_190)
);

BUFx6f_ASAP7_75t_L g191 ( 
.A(n_144),
.Y(n_191)
);

BUFx6f_ASAP7_75t_L g192 ( 
.A(n_144),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_171),
.B(n_0),
.Y(n_193)
);

OA21x2_ASAP7_75t_L g194 ( 
.A1(n_111),
.A2(n_0),
.B(n_4),
.Y(n_194)
);

INVx3_ASAP7_75t_L g195 ( 
.A(n_118),
.Y(n_195)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_184),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_150),
.B(n_4),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_171),
.B(n_7),
.Y(n_198)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_111),
.Y(n_199)
);

BUFx12f_ASAP7_75t_L g200 ( 
.A(n_114),
.Y(n_200)
);

BUFx3_ASAP7_75t_L g201 ( 
.A(n_118),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_183),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_183),
.Y(n_203)
);

INVx3_ASAP7_75t_L g204 ( 
.A(n_99),
.Y(n_204)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_116),
.Y(n_205)
);

INVx6_ASAP7_75t_L g206 ( 
.A(n_114),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_182),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_156),
.Y(n_208)
);

BUFx6f_ASAP7_75t_L g209 ( 
.A(n_144),
.Y(n_209)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_123),
.Y(n_210)
);

AND2x2_ASAP7_75t_SL g211 ( 
.A(n_166),
.B(n_9),
.Y(n_211)
);

OA21x2_ASAP7_75t_L g212 ( 
.A1(n_149),
.A2(n_11),
.B(n_17),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_186),
.B(n_28),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_122),
.B(n_39),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_97),
.A2(n_42),
.B1(n_52),
.B2(n_56),
.Y(n_215)
);

BUFx6f_ASAP7_75t_L g216 ( 
.A(n_144),
.Y(n_216)
);

BUFx3_ASAP7_75t_L g217 ( 
.A(n_176),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_156),
.Y(n_218)
);

BUFx2_ASAP7_75t_L g219 ( 
.A(n_178),
.Y(n_219)
);

BUFx8_ASAP7_75t_SL g220 ( 
.A(n_182),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_97),
.A2(n_65),
.B1(n_66),
.B2(n_68),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_190),
.A2(n_77),
.B1(n_85),
.B2(n_128),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_152),
.Y(n_223)
);

AND2x2_ASAP7_75t_L g224 ( 
.A(n_153),
.B(n_170),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_117),
.A2(n_189),
.B1(n_137),
.B2(n_167),
.Y(n_225)
);

HB1xp67_ASAP7_75t_L g226 ( 
.A(n_133),
.Y(n_226)
);

AND2x4_ASAP7_75t_L g227 ( 
.A(n_99),
.B(n_131),
.Y(n_227)
);

AND2x4_ASAP7_75t_L g228 ( 
.A(n_131),
.B(n_181),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_173),
.Y(n_229)
);

AND2x2_ASAP7_75t_L g230 ( 
.A(n_175),
.B(n_176),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_181),
.B(n_102),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_103),
.B(n_104),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_110),
.B(n_106),
.Y(n_233)
);

INVx3_ASAP7_75t_L g234 ( 
.A(n_185),
.Y(n_234)
);

BUFx2_ASAP7_75t_L g235 ( 
.A(n_158),
.Y(n_235)
);

AND2x4_ASAP7_75t_L g236 ( 
.A(n_109),
.B(n_187),
.Y(n_236)
);

BUFx6f_ASAP7_75t_L g237 ( 
.A(n_185),
.Y(n_237)
);

HB1xp67_ASAP7_75t_L g238 ( 
.A(n_160),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_112),
.B(n_148),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_113),
.Y(n_240)
);

BUFx3_ASAP7_75t_L g241 ( 
.A(n_115),
.Y(n_241)
);

AND2x4_ASAP7_75t_L g242 ( 
.A(n_121),
.B(n_146),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_126),
.Y(n_243)
);

BUFx6f_ASAP7_75t_L g244 ( 
.A(n_127),
.Y(n_244)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_129),
.Y(n_245)
);

OA21x2_ASAP7_75t_L g246 ( 
.A1(n_132),
.A2(n_143),
.B(n_134),
.Y(n_246)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_136),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_154),
.B(n_174),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_155),
.B(n_168),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_162),
.Y(n_250)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_163),
.Y(n_251)
);

HB1xp67_ASAP7_75t_L g252 ( 
.A(n_169),
.Y(n_252)
);

INVxp67_ASAP7_75t_L g253 ( 
.A(n_188),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_98),
.Y(n_254)
);

BUFx6f_ASAP7_75t_L g255 ( 
.A(n_101),
.Y(n_255)
);

OA21x2_ASAP7_75t_L g256 ( 
.A1(n_179),
.A2(n_157),
.B(n_135),
.Y(n_256)
);

INVxp67_ASAP7_75t_SL g257 ( 
.A(n_195),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_245),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_254),
.B(n_140),
.Y(n_259)
);

XOR2x2_ASAP7_75t_L g260 ( 
.A(n_211),
.B(n_100),
.Y(n_260)
);

INVx4_ASAP7_75t_L g261 ( 
.A(n_255),
.Y(n_261)
);

AOI22xp33_ASAP7_75t_L g262 ( 
.A1(n_227),
.A2(n_100),
.B1(n_159),
.B2(n_107),
.Y(n_262)
);

INVx1_ASAP7_75t_SL g263 ( 
.A(n_220),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_255),
.B(n_233),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_247),
.Y(n_265)
);

AND2x6_ASAP7_75t_L g266 ( 
.A(n_191),
.B(n_159),
.Y(n_266)
);

AND3x2_ASAP7_75t_L g267 ( 
.A(n_193),
.B(n_105),
.C(n_108),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_247),
.Y(n_268)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_234),
.Y(n_269)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_234),
.Y(n_270)
);

INVx2_ASAP7_75t_SL g271 ( 
.A(n_206),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_211),
.B(n_119),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_255),
.B(n_180),
.Y(n_273)
);

INVx4_ASAP7_75t_L g274 ( 
.A(n_256),
.Y(n_274)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_234),
.Y(n_275)
);

OR2x6_ASAP7_75t_L g276 ( 
.A(n_197),
.B(n_120),
.Y(n_276)
);

NOR2x1p5_ASAP7_75t_L g277 ( 
.A(n_200),
.B(n_124),
.Y(n_277)
);

BUFx6f_ASAP7_75t_L g278 ( 
.A(n_191),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_253),
.B(n_125),
.Y(n_279)
);

INVx3_ASAP7_75t_L g280 ( 
.A(n_191),
.Y(n_280)
);

INVx2_ASAP7_75t_SL g281 ( 
.A(n_206),
.Y(n_281)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_196),
.Y(n_282)
);

INVx2_ASAP7_75t_SL g283 ( 
.A(n_206),
.Y(n_283)
);

BUFx3_ASAP7_75t_L g284 ( 
.A(n_201),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_198),
.B(n_130),
.Y(n_285)
);

OR2x2_ASAP7_75t_L g286 ( 
.A(n_235),
.B(n_138),
.Y(n_286)
);

BUFx8_ASAP7_75t_SL g287 ( 
.A(n_220),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_251),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_251),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_195),
.B(n_177),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_195),
.B(n_139),
.Y(n_291)
);

INVx3_ASAP7_75t_L g292 ( 
.A(n_191),
.Y(n_292)
);

AOI21x1_ASAP7_75t_L g293 ( 
.A1(n_231),
.A2(n_172),
.B(n_142),
.Y(n_293)
);

INVx2_ASAP7_75t_SL g294 ( 
.A(n_206),
.Y(n_294)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_196),
.Y(n_295)
);

NAND3xp33_ASAP7_75t_L g296 ( 
.A(n_232),
.B(n_141),
.C(n_145),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_SL g297 ( 
.A(n_213),
.B(n_147),
.Y(n_297)
);

NAND2xp33_ASAP7_75t_SL g298 ( 
.A(n_230),
.B(n_151),
.Y(n_298)
);

OR2x6_ASAP7_75t_L g299 ( 
.A(n_215),
.B(n_161),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_SL g300 ( 
.A(n_222),
.B(n_164),
.Y(n_300)
);

BUFx3_ASAP7_75t_L g301 ( 
.A(n_201),
.Y(n_301)
);

NAND3xp33_ASAP7_75t_L g302 ( 
.A(n_239),
.B(n_165),
.C(n_248),
.Y(n_302)
);

INVx3_ASAP7_75t_L g303 ( 
.A(n_191),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_257),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_269),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_264),
.B(n_226),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_259),
.B(n_238),
.Y(n_307)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_280),
.Y(n_308)
);

BUFx8_ASAP7_75t_L g309 ( 
.A(n_266),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_270),
.Y(n_310)
);

INVxp67_ASAP7_75t_L g311 ( 
.A(n_286),
.Y(n_311)
);

INVxp33_ASAP7_75t_L g312 ( 
.A(n_287),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_270),
.Y(n_313)
);

OAI221xp5_ASAP7_75t_L g314 ( 
.A1(n_262),
.A2(n_249),
.B1(n_250),
.B2(n_240),
.C(n_243),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_290),
.B(n_256),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_291),
.B(n_242),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_273),
.B(n_242),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_261),
.B(n_236),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_L g319 ( 
.A1(n_272),
.A2(n_252),
.B1(n_235),
.B2(n_219),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_SL g320 ( 
.A(n_298),
.B(n_217),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_275),
.Y(n_321)
);

BUFx8_ASAP7_75t_L g322 ( 
.A(n_266),
.Y(n_322)
);

AND2x2_ASAP7_75t_L g323 ( 
.A(n_284),
.B(n_217),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_302),
.B(n_241),
.Y(n_324)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_292),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_SL g326 ( 
.A(n_274),
.B(n_214),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_SL g327 ( 
.A(n_298),
.B(n_200),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_279),
.B(n_241),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_SL g329 ( 
.A(n_284),
.B(n_225),
.Y(n_329)
);

INVxp67_ASAP7_75t_L g330 ( 
.A(n_301),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_297),
.B(n_246),
.Y(n_331)
);

CKINVDCx8_ASAP7_75t_R g332 ( 
.A(n_266),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_285),
.B(n_246),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_296),
.B(n_208),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_SL g335 ( 
.A(n_301),
.B(n_221),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_271),
.B(n_227),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_SL g337 ( 
.A(n_271),
.B(n_228),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_275),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_287),
.Y(n_339)
);

OAI22xp5_ASAP7_75t_L g340 ( 
.A1(n_276),
.A2(n_228),
.B1(n_227),
.B2(n_218),
.Y(n_340)
);

INVx2_ASAP7_75t_L g341 ( 
.A(n_292),
.Y(n_341)
);

BUFx3_ASAP7_75t_L g342 ( 
.A(n_294),
.Y(n_342)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_303),
.Y(n_343)
);

INVx3_ASAP7_75t_L g344 ( 
.A(n_278),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_L g345 ( 
.A1(n_276),
.A2(n_208),
.B1(n_218),
.B2(n_229),
.Y(n_345)
);

INVx8_ASAP7_75t_L g346 ( 
.A(n_266),
.Y(n_346)
);

BUFx6f_ASAP7_75t_L g347 ( 
.A(n_278),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g348 ( 
.A(n_300),
.B(n_250),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_328),
.B(n_266),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_SL g350 ( 
.A(n_307),
.B(n_306),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_328),
.B(n_266),
.Y(n_351)
);

NOR3xp33_ASAP7_75t_L g352 ( 
.A(n_314),
.B(n_329),
.C(n_311),
.Y(n_352)
);

OAI21xp5_ASAP7_75t_L g353 ( 
.A1(n_315),
.A2(n_293),
.B(n_295),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_317),
.B(n_316),
.Y(n_354)
);

AND2x2_ASAP7_75t_L g355 ( 
.A(n_306),
.B(n_283),
.Y(n_355)
);

INVx2_ASAP7_75t_L g356 ( 
.A(n_305),
.Y(n_356)
);

AND2x4_ASAP7_75t_L g357 ( 
.A(n_330),
.B(n_283),
.Y(n_357)
);

AOI22xp33_ASAP7_75t_SL g358 ( 
.A1(n_348),
.A2(n_276),
.B1(n_207),
.B2(n_260),
.Y(n_358)
);

AND2x2_ASAP7_75t_L g359 ( 
.A(n_311),
.B(n_281),
.Y(n_359)
);

O2A1O1Ixp33_ASAP7_75t_L g360 ( 
.A1(n_326),
.A2(n_243),
.B(n_240),
.C(n_300),
.Y(n_360)
);

INVxp67_ASAP7_75t_L g361 ( 
.A(n_307),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_SL g362 ( 
.A(n_332),
.B(n_299),
.Y(n_362)
);

INVx2_ASAP7_75t_L g363 ( 
.A(n_310),
.Y(n_363)
);

AOI22xp5_ASAP7_75t_L g364 ( 
.A1(n_324),
.A2(n_299),
.B1(n_260),
.B2(n_267),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_334),
.B(n_282),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_336),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_334),
.B(n_282),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_SL g368 ( 
.A(n_345),
.B(n_258),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_SL g369 ( 
.A(n_319),
.B(n_288),
.Y(n_369)
);

OAI22xp5_ASAP7_75t_L g370 ( 
.A1(n_335),
.A2(n_299),
.B1(n_194),
.B2(n_223),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_L g371 ( 
.A(n_330),
.B(n_299),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_313),
.Y(n_372)
);

HB1xp67_ASAP7_75t_L g373 ( 
.A(n_337),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_321),
.B(n_338),
.Y(n_374)
);

INVxp67_ASAP7_75t_L g375 ( 
.A(n_320),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_308),
.Y(n_376)
);

OR2x6_ASAP7_75t_SL g377 ( 
.A(n_339),
.B(n_207),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_344),
.B(n_289),
.Y(n_378)
);

AOI22xp5_ASAP7_75t_L g379 ( 
.A1(n_327),
.A2(n_277),
.B1(n_265),
.B2(n_268),
.Y(n_379)
);

OR2x2_ASAP7_75t_L g380 ( 
.A(n_342),
.B(n_263),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_325),
.B(n_244),
.Y(n_381)
);

AND2x2_ASAP7_75t_L g382 ( 
.A(n_341),
.B(n_224),
.Y(n_382)
);

OAI22xp5_ASAP7_75t_L g383 ( 
.A1(n_343),
.A2(n_194),
.B1(n_223),
.B2(n_205),
.Y(n_383)
);

OAI22xp5_ASAP7_75t_L g384 ( 
.A1(n_312),
.A2(n_205),
.B1(n_210),
.B2(n_199),
.Y(n_384)
);

INVx1_ASAP7_75t_SL g385 ( 
.A(n_347),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_R g386 ( 
.A(n_309),
.B(n_204),
.Y(n_386)
);

HB1xp67_ASAP7_75t_L g387 ( 
.A(n_322),
.Y(n_387)
);

OR2x6_ASAP7_75t_L g388 ( 
.A(n_322),
.B(n_199),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_L g389 ( 
.A(n_307),
.B(n_244),
.Y(n_389)
);

AOI21xp5_ASAP7_75t_L g390 ( 
.A1(n_318),
.A2(n_192),
.B(n_237),
.Y(n_390)
);

AOI21xp5_ASAP7_75t_L g391 ( 
.A1(n_318),
.A2(n_192),
.B(n_237),
.Y(n_391)
);

BUFx6f_ASAP7_75t_L g392 ( 
.A(n_342),
.Y(n_392)
);

BUFx2_ASAP7_75t_SL g393 ( 
.A(n_323),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_328),
.B(n_244),
.Y(n_394)
);

AOI22xp5_ASAP7_75t_L g395 ( 
.A1(n_348),
.A2(n_212),
.B1(n_204),
.B2(n_203),
.Y(n_395)
);

AOI21xp5_ASAP7_75t_L g396 ( 
.A1(n_318),
.A2(n_192),
.B(n_209),
.Y(n_396)
);

NOR2xp67_ASAP7_75t_L g397 ( 
.A(n_311),
.B(n_204),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_304),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_328),
.B(n_192),
.Y(n_399)
);

INVx3_ASAP7_75t_L g400 ( 
.A(n_344),
.Y(n_400)
);

AOI21xp5_ASAP7_75t_L g401 ( 
.A1(n_354),
.A2(n_209),
.B(n_216),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_SL g402 ( 
.A(n_361),
.B(n_202),
.Y(n_402)
);

INVx2_ASAP7_75t_SL g403 ( 
.A(n_359),
.Y(n_403)
);

AO21x2_ASAP7_75t_L g404 ( 
.A1(n_349),
.A2(n_351),
.B(n_395),
.Y(n_404)
);

INVx5_ASAP7_75t_L g405 ( 
.A(n_388),
.Y(n_405)
);

INVx2_ASAP7_75t_L g406 ( 
.A(n_356),
.Y(n_406)
);

AO32x2_ASAP7_75t_L g407 ( 
.A1(n_383),
.A2(n_370),
.A3(n_384),
.B1(n_360),
.B2(n_362),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_389),
.B(n_366),
.Y(n_408)
);

AOI21x1_ASAP7_75t_L g409 ( 
.A1(n_365),
.A2(n_367),
.B(n_399),
.Y(n_409)
);

BUFx6f_ASAP7_75t_L g410 ( 
.A(n_392),
.Y(n_410)
);

A2O1A1Ixp33_ASAP7_75t_L g411 ( 
.A1(n_352),
.A2(n_371),
.B(n_375),
.C(n_398),
.Y(n_411)
);

BUFx6f_ASAP7_75t_L g412 ( 
.A(n_392),
.Y(n_412)
);

BUFx3_ASAP7_75t_L g413 ( 
.A(n_392),
.Y(n_413)
);

OAI22x1_ASAP7_75t_L g414 ( 
.A1(n_364),
.A2(n_358),
.B1(n_355),
.B2(n_379),
.Y(n_414)
);

NOR2xp33_ASAP7_75t_L g415 ( 
.A(n_393),
.B(n_362),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_394),
.B(n_397),
.Y(n_416)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_363),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_372),
.B(n_382),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_SL g419 ( 
.A(n_357),
.B(n_373),
.Y(n_419)
);

BUFx6f_ASAP7_75t_L g420 ( 
.A(n_388),
.Y(n_420)
);

AOI22xp5_ASAP7_75t_L g421 ( 
.A1(n_357),
.A2(n_369),
.B1(n_368),
.B2(n_376),
.Y(n_421)
);

AOI21xp5_ASAP7_75t_L g422 ( 
.A1(n_385),
.A2(n_378),
.B(n_381),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_385),
.B(n_400),
.Y(n_423)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_384),
.Y(n_424)
);

AND2x2_ASAP7_75t_L g425 ( 
.A(n_380),
.B(n_387),
.Y(n_425)
);

INVx3_ASAP7_75t_SL g426 ( 
.A(n_377),
.Y(n_426)
);

AOI21xp5_ASAP7_75t_L g427 ( 
.A1(n_390),
.A2(n_391),
.B(n_396),
.Y(n_427)
);

AOI21xp5_ASAP7_75t_L g428 ( 
.A1(n_386),
.A2(n_346),
.B(n_354),
.Y(n_428)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_356),
.Y(n_429)
);

INVx2_ASAP7_75t_L g430 ( 
.A(n_356),
.Y(n_430)
);

BUFx3_ASAP7_75t_L g431 ( 
.A(n_392),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_374),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_354),
.B(n_361),
.Y(n_433)
);

BUFx6f_ASAP7_75t_L g434 ( 
.A(n_392),
.Y(n_434)
);

BUFx2_ASAP7_75t_L g435 ( 
.A(n_359),
.Y(n_435)
);

AO22x2_ASAP7_75t_L g436 ( 
.A1(n_350),
.A2(n_361),
.B1(n_370),
.B2(n_340),
.Y(n_436)
);

BUFx6f_ASAP7_75t_L g437 ( 
.A(n_392),
.Y(n_437)
);

OAI21xp5_ASAP7_75t_L g438 ( 
.A1(n_353),
.A2(n_331),
.B(n_333),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_354),
.B(n_361),
.Y(n_439)
);

OR2x6_ASAP7_75t_L g440 ( 
.A(n_388),
.B(n_393),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_L g441 ( 
.A(n_361),
.B(n_350),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_354),
.B(n_361),
.Y(n_442)
);

NAND3xp33_ASAP7_75t_SL g443 ( 
.A(n_350),
.B(n_358),
.C(n_361),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_374),
.Y(n_444)
);

CKINVDCx14_ASAP7_75t_R g445 ( 
.A(n_377),
.Y(n_445)
);

OAI21xp5_ASAP7_75t_L g446 ( 
.A1(n_353),
.A2(n_331),
.B(n_333),
.Y(n_446)
);

NAND3xp33_ASAP7_75t_L g447 ( 
.A(n_350),
.B(n_361),
.C(n_262),
.Y(n_447)
);

NAND3xp33_ASAP7_75t_L g448 ( 
.A(n_447),
.B(n_411),
.C(n_439),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_406),
.Y(n_449)
);

OR2x2_ASAP7_75t_L g450 ( 
.A(n_433),
.B(n_442),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_417),
.Y(n_451)
);

NOR2xp67_ASAP7_75t_L g452 ( 
.A(n_443),
.B(n_403),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_432),
.B(n_444),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_441),
.B(n_408),
.Y(n_454)
);

AOI21x1_ASAP7_75t_L g455 ( 
.A1(n_409),
.A2(n_416),
.B(n_422),
.Y(n_455)
);

BUFx6f_ASAP7_75t_L g456 ( 
.A(n_410),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_429),
.Y(n_457)
);

AND2x4_ASAP7_75t_L g458 ( 
.A(n_413),
.B(n_431),
.Y(n_458)
);

AOI21x1_ASAP7_75t_L g459 ( 
.A1(n_438),
.A2(n_446),
.B(n_427),
.Y(n_459)
);

O2A1O1Ixp33_ASAP7_75t_L g460 ( 
.A1(n_424),
.A2(n_402),
.B(n_415),
.C(n_418),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_436),
.B(n_421),
.Y(n_461)
);

AND2x2_ASAP7_75t_L g462 ( 
.A(n_435),
.B(n_425),
.Y(n_462)
);

OAI21xp5_ASAP7_75t_L g463 ( 
.A1(n_401),
.A2(n_423),
.B(n_428),
.Y(n_463)
);

AND2x2_ASAP7_75t_L g464 ( 
.A(n_419),
.B(n_414),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_436),
.B(n_430),
.Y(n_465)
);

HB1xp67_ASAP7_75t_L g466 ( 
.A(n_410),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_412),
.B(n_434),
.Y(n_467)
);

AO21x1_ASAP7_75t_L g468 ( 
.A1(n_407),
.A2(n_404),
.B(n_440),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_412),
.Y(n_469)
);

OAI21x1_ASAP7_75t_L g470 ( 
.A1(n_407),
.A2(n_405),
.B(n_440),
.Y(n_470)
);

INVx6_ASAP7_75t_L g471 ( 
.A(n_412),
.Y(n_471)
);

INVx2_ASAP7_75t_L g472 ( 
.A(n_434),
.Y(n_472)
);

OAI21x1_ASAP7_75t_L g473 ( 
.A1(n_405),
.A2(n_420),
.B(n_437),
.Y(n_473)
);

INVx2_ASAP7_75t_L g474 ( 
.A(n_437),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_437),
.Y(n_475)
);

NOR2xp33_ASAP7_75t_R g476 ( 
.A(n_450),
.B(n_445),
.Y(n_476)
);

OAI21x1_ASAP7_75t_SL g477 ( 
.A1(n_468),
.A2(n_405),
.B(n_420),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_453),
.Y(n_478)
);

AOI21x1_ASAP7_75t_L g479 ( 
.A1(n_455),
.A2(n_420),
.B(n_426),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_465),
.Y(n_480)
);

INVx1_ASAP7_75t_SL g481 ( 
.A(n_462),
.Y(n_481)
);

INVx2_ASAP7_75t_L g482 ( 
.A(n_459),
.Y(n_482)
);

BUFx10_ASAP7_75t_L g483 ( 
.A(n_458),
.Y(n_483)
);

HB1xp67_ASAP7_75t_L g484 ( 
.A(n_466),
.Y(n_484)
);

OR2x2_ASAP7_75t_L g485 ( 
.A(n_454),
.B(n_448),
.Y(n_485)
);

OR2x2_ASAP7_75t_L g486 ( 
.A(n_461),
.B(n_464),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_449),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g488 ( 
.A(n_460),
.B(n_452),
.Y(n_488)
);

HB1xp67_ASAP7_75t_L g489 ( 
.A(n_466),
.Y(n_489)
);

INVx3_ASAP7_75t_L g490 ( 
.A(n_473),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_451),
.Y(n_491)
);

AND2x2_ASAP7_75t_L g492 ( 
.A(n_457),
.B(n_470),
.Y(n_492)
);

HB1xp67_ASAP7_75t_L g493 ( 
.A(n_492),
.Y(n_493)
);

INVx1_ASAP7_75t_SL g494 ( 
.A(n_481),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_492),
.Y(n_495)
);

AND2x2_ASAP7_75t_L g496 ( 
.A(n_480),
.B(n_486),
.Y(n_496)
);

AND2x2_ASAP7_75t_L g497 ( 
.A(n_478),
.B(n_485),
.Y(n_497)
);

AND2x2_ASAP7_75t_L g498 ( 
.A(n_485),
.B(n_474),
.Y(n_498)
);

OR2x2_ASAP7_75t_L g499 ( 
.A(n_486),
.B(n_467),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_488),
.B(n_472),
.Y(n_500)
);

INVxp67_ASAP7_75t_L g501 ( 
.A(n_484),
.Y(n_501)
);

BUFx2_ASAP7_75t_L g502 ( 
.A(n_493),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_495),
.Y(n_503)
);

AND2x4_ASAP7_75t_L g504 ( 
.A(n_498),
.B(n_490),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_497),
.B(n_489),
.Y(n_505)
);

NOR2xp33_ASAP7_75t_L g506 ( 
.A(n_494),
.B(n_458),
.Y(n_506)
);

AND2x2_ASAP7_75t_L g507 ( 
.A(n_496),
.B(n_482),
.Y(n_507)
);

OR2x2_ASAP7_75t_L g508 ( 
.A(n_502),
.B(n_499),
.Y(n_508)
);

INVxp67_ASAP7_75t_L g509 ( 
.A(n_506),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_505),
.B(n_497),
.Y(n_510)
);

OR2x2_ASAP7_75t_L g511 ( 
.A(n_502),
.B(n_499),
.Y(n_511)
);

AND2x4_ASAP7_75t_L g512 ( 
.A(n_504),
.B(n_503),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_503),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_513),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_508),
.Y(n_515)
);

OAI22xp5_ASAP7_75t_L g516 ( 
.A1(n_509),
.A2(n_494),
.B1(n_501),
.B2(n_500),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_511),
.Y(n_517)
);

AOI21xp33_ASAP7_75t_L g518 ( 
.A1(n_510),
.A2(n_477),
.B(n_500),
.Y(n_518)
);

INVxp67_ASAP7_75t_L g519 ( 
.A(n_512),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_512),
.B(n_507),
.Y(n_520)
);

INVx2_ASAP7_75t_L g521 ( 
.A(n_512),
.Y(n_521)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_521),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_514),
.Y(n_523)
);

INVx2_ASAP7_75t_L g524 ( 
.A(n_515),
.Y(n_524)
);

INVx1_ASAP7_75t_SL g525 ( 
.A(n_517),
.Y(n_525)
);

HB1xp67_ASAP7_75t_L g526 ( 
.A(n_525),
.Y(n_526)
);

AOI211x1_ASAP7_75t_SL g527 ( 
.A1(n_526),
.A2(n_516),
.B(n_518),
.C(n_524),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_527),
.B(n_525),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_528),
.B(n_523),
.Y(n_529)
);

AOI221xp5_ASAP7_75t_L g530 ( 
.A1(n_529),
.A2(n_516),
.B1(n_522),
.B2(n_519),
.C(n_501),
.Y(n_530)
);

NAND3x1_ASAP7_75t_L g531 ( 
.A(n_529),
.B(n_476),
.C(n_479),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_530),
.B(n_520),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_531),
.Y(n_533)
);

AOI22x1_ASAP7_75t_L g534 ( 
.A1(n_533),
.A2(n_477),
.B1(n_458),
.B2(n_456),
.Y(n_534)
);

CKINVDCx16_ASAP7_75t_R g535 ( 
.A(n_534),
.Y(n_535)
);

AOI21xp5_ASAP7_75t_L g536 ( 
.A1(n_534),
.A2(n_532),
.B(n_487),
.Y(n_536)
);

OA21x2_ASAP7_75t_L g537 ( 
.A1(n_536),
.A2(n_463),
.B(n_491),
.Y(n_537)
);

AND2x2_ASAP7_75t_L g538 ( 
.A(n_537),
.B(n_535),
.Y(n_538)
);

AOI22xp33_ASAP7_75t_SL g539 ( 
.A1(n_538),
.A2(n_471),
.B1(n_456),
.B2(n_483),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_539),
.B(n_475),
.Y(n_540)
);

AOI22xp5_ASAP7_75t_L g541 ( 
.A1(n_540),
.A2(n_471),
.B1(n_456),
.B2(n_469),
.Y(n_541)
);


endmodule