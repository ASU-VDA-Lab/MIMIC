module fake_jpeg_9573_n_172 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_172);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_172;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_57;
wire n_21;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g14 ( 
.A(n_13),
.Y(n_14)
);

INVx6_ASAP7_75t_L g15 ( 
.A(n_2),
.Y(n_15)
);

BUFx12_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

BUFx10_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_8),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_27),
.Y(n_30)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_30),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_22),
.B(n_0),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_31),
.B(n_35),
.Y(n_49)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_27),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_32),
.B(n_34),
.Y(n_53)
);

INVx5_ASAP7_75t_L g33 ( 
.A(n_18),
.Y(n_33)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_16),
.B(n_0),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_22),
.B(n_1),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_24),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_23),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_37),
.B(n_20),
.Y(n_47)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_24),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_38),
.B(n_17),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

AOI21xp33_ASAP7_75t_L g40 ( 
.A1(n_31),
.A2(n_15),
.B(n_20),
.Y(n_40)
);

AND2x2_ASAP7_75t_L g60 ( 
.A(n_40),
.B(n_45),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g41 ( 
.A1(n_38),
.A2(n_29),
.B1(n_15),
.B2(n_26),
.Y(n_41)
);

INVxp67_ASAP7_75t_L g65 ( 
.A(n_41),
.Y(n_65)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_42),
.B(n_50),
.Y(n_58)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_45),
.B(n_47),
.Y(n_63)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_46),
.Y(n_62)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_34),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_48),
.B(n_54),
.Y(n_72)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

BUFx2_ASAP7_75t_L g51 ( 
.A(n_30),
.Y(n_51)
);

CKINVDCx16_ASAP7_75t_R g59 ( 
.A(n_51),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_32),
.A2(n_29),
.B1(n_15),
.B2(n_26),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_52),
.A2(n_19),
.B1(n_28),
.B2(n_25),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_37),
.B(n_17),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_49),
.B(n_14),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_57),
.B(n_16),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_60),
.B(n_64),
.Y(n_79)
);

HB1xp67_ASAP7_75t_L g61 ( 
.A(n_51),
.Y(n_61)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_61),
.Y(n_76)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_54),
.Y(n_64)
);

INVx1_ASAP7_75t_SL g66 ( 
.A(n_42),
.Y(n_66)
);

CKINVDCx16_ASAP7_75t_R g89 ( 
.A(n_66),
.Y(n_89)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_47),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_67),
.B(n_1),
.Y(n_90)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_51),
.Y(n_68)
);

INVxp67_ASAP7_75t_L g78 ( 
.A(n_68),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_L g69 ( 
.A1(n_49),
.A2(n_19),
.B1(n_26),
.B2(n_28),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_69),
.A2(n_19),
.B1(n_56),
.B2(n_44),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_L g82 ( 
.A1(n_70),
.A2(n_56),
.B1(n_44),
.B2(n_50),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_48),
.B(n_23),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_71),
.B(n_73),
.C(n_53),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_53),
.B(n_14),
.C(n_25),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_74),
.A2(n_77),
.B1(n_88),
.B2(n_59),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_75),
.B(n_86),
.Y(n_101)
);

O2A1O1Ixp33_ASAP7_75t_L g77 ( 
.A1(n_70),
.A2(n_43),
.B(n_39),
.C(n_36),
.Y(n_77)
);

XNOR2xp5_ASAP7_75t_L g80 ( 
.A(n_72),
.B(n_43),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_80),
.B(n_81),
.C(n_73),
.Y(n_94)
);

XOR2xp5_ASAP7_75t_L g81 ( 
.A(n_72),
.B(n_18),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_82),
.A2(n_66),
.B1(n_62),
.B2(n_55),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_L g83 ( 
.A1(n_64),
.A2(n_21),
.B(n_18),
.Y(n_83)
);

OAI21xp5_ASAP7_75t_L g93 ( 
.A1(n_83),
.A2(n_65),
.B(n_59),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_60),
.B(n_39),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_84),
.B(n_85),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_60),
.B(n_63),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_58),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_87),
.B(n_90),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_65),
.A2(n_44),
.B1(n_55),
.B2(n_21),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_63),
.B(n_55),
.Y(n_91)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_91),
.Y(n_103)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_71),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_92),
.B(n_16),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_SL g124 ( 
.A(n_93),
.B(n_87),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_L g118 ( 
.A(n_94),
.B(n_85),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_88),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_95),
.Y(n_115)
);

NOR3xp33_ASAP7_75t_SL g96 ( 
.A(n_79),
.B(n_71),
.C(n_67),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_96),
.B(n_106),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_97),
.A2(n_98),
.B1(n_89),
.B2(n_76),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_81),
.B(n_62),
.C(n_68),
.Y(n_99)
);

XOR2xp5_ASAP7_75t_L g119 ( 
.A(n_99),
.B(n_105),
.Y(n_119)
);

AND2x2_ASAP7_75t_SL g102 ( 
.A(n_84),
.B(n_21),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_102),
.B(n_108),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_86),
.B(n_16),
.Y(n_104)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_104),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_80),
.B(n_30),
.C(n_21),
.Y(n_105)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_91),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_90),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_109),
.B(n_92),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_110),
.A2(n_122),
.B1(n_123),
.B2(n_96),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_112),
.B(n_121),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_103),
.B(n_79),
.Y(n_114)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_114),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_103),
.B(n_106),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_116),
.B(n_100),
.Y(n_131)
);

BUFx5_ASAP7_75t_L g117 ( 
.A(n_101),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_117),
.B(n_99),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_118),
.B(n_124),
.C(n_94),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_98),
.Y(n_121)
);

AOI21xp5_ASAP7_75t_L g122 ( 
.A1(n_93),
.A2(n_83),
.B(n_89),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_95),
.A2(n_77),
.B1(n_74),
.B2(n_75),
.Y(n_123)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_126),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_128),
.B(n_129),
.C(n_119),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_119),
.B(n_100),
.C(n_105),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_115),
.A2(n_97),
.B1(n_108),
.B2(n_102),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_130),
.A2(n_135),
.B1(n_113),
.B2(n_114),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_131),
.B(n_132),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_111),
.B(n_107),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_113),
.B(n_76),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_SL g146 ( 
.A1(n_133),
.A2(n_136),
.B(n_1),
.Y(n_146)
);

AOI21xp5_ASAP7_75t_L g141 ( 
.A1(n_134),
.A2(n_120),
.B(n_117),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_115),
.A2(n_102),
.B1(n_78),
.B2(n_21),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_116),
.Y(n_136)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_138),
.Y(n_147)
);

XOR2x1_ASAP7_75t_SL g139 ( 
.A(n_130),
.B(n_122),
.Y(n_139)
);

AOI31xp67_ASAP7_75t_L g151 ( 
.A1(n_139),
.A2(n_135),
.A3(n_125),
.B(n_4),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_140),
.B(n_142),
.C(n_11),
.Y(n_152)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_141),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_128),
.B(n_118),
.C(n_124),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_SL g143 ( 
.A(n_131),
.B(n_121),
.Y(n_143)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_143),
.B(n_145),
.Y(n_153)
);

XOR2xp5_ASAP7_75t_L g145 ( 
.A(n_129),
.B(n_12),
.Y(n_145)
);

AOI21xp5_ASAP7_75t_SL g150 ( 
.A1(n_146),
.A2(n_125),
.B(n_12),
.Y(n_150)
);

HB1xp67_ASAP7_75t_L g148 ( 
.A(n_139),
.Y(n_148)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_148),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g149 ( 
.A(n_140),
.B(n_127),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_149),
.B(n_137),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_150),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_151),
.A2(n_154),
.B1(n_147),
.B2(n_4),
.Y(n_157)
);

AOI21xp5_ASAP7_75t_L g158 ( 
.A1(n_152),
.A2(n_144),
.B(n_142),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_SL g165 ( 
.A(n_155),
.B(n_158),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_157),
.B(n_5),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_148),
.A2(n_143),
.B1(n_138),
.B2(n_145),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_159),
.B(n_2),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_SL g161 ( 
.A1(n_160),
.A2(n_153),
.B(n_3),
.Y(n_161)
);

AOI21xp5_ASAP7_75t_L g167 ( 
.A1(n_161),
.A2(n_162),
.B(n_6),
.Y(n_167)
);

AOI21xp5_ASAP7_75t_L g163 ( 
.A1(n_156),
.A2(n_2),
.B(n_3),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_L g166 ( 
.A1(n_163),
.A2(n_6),
.B(n_7),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_164),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_166),
.B(n_167),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_L g170 ( 
.A1(n_168),
.A2(n_165),
.B(n_162),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_170),
.B(n_9),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_171),
.B(n_169),
.Y(n_172)
);


endmodule