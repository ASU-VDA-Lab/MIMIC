module fake_netlist_6_651_n_2098 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_193, n_147, n_154, n_191, n_88, n_3, n_209, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_199, n_138, n_22, n_161, n_208, n_68, n_166, n_28, n_184, n_50, n_158, n_49, n_7, n_210, n_83, n_206, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_188, n_102, n_186, n_204, n_0, n_87, n_195, n_189, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_197, n_11, n_137, n_17, n_23, n_203, n_142, n_20, n_143, n_207, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_205, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_202, n_94, n_97, n_108, n_58, n_116, n_211, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_196, n_200, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_198, n_104, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_190, n_14, n_123, n_136, n_72, n_187, n_89, n_173, n_201, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_194, n_171, n_31, n_192, n_57, n_169, n_53, n_51, n_44, n_56, n_2098);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_193;
input n_147;
input n_154;
input n_191;
input n_88;
input n_3;
input n_209;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_199;
input n_138;
input n_22;
input n_161;
input n_208;
input n_68;
input n_166;
input n_28;
input n_184;
input n_50;
input n_158;
input n_49;
input n_7;
input n_210;
input n_83;
input n_206;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_188;
input n_102;
input n_186;
input n_204;
input n_0;
input n_87;
input n_195;
input n_189;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_197;
input n_11;
input n_137;
input n_17;
input n_23;
input n_203;
input n_142;
input n_20;
input n_143;
input n_207;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_205;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_202;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_211;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_196;
input n_200;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_190;
input n_14;
input n_123;
input n_136;
input n_72;
input n_187;
input n_89;
input n_173;
input n_201;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_194;
input n_171;
input n_31;
input n_192;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_2098;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_2003;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_1853;
wire n_783;
wire n_1738;
wire n_798;
wire n_1575;
wire n_1854;
wire n_1923;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_2051;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1688;
wire n_1691;
wire n_1975;
wire n_1009;
wire n_1743;
wire n_1930;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1991;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_1844;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_1985;
wire n_447;
wire n_1803;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1867;
wire n_1704;
wire n_1078;
wire n_250;
wire n_544;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_2019;
wire n_836;
wire n_375;
wire n_2074;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_2018;
wire n_2094;
wire n_1903;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_616;
wire n_658;
wire n_1874;
wire n_1119;
wire n_2013;
wire n_428;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_2044;
wire n_1954;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_1971;
wire n_2058;
wire n_2090;
wire n_405;
wire n_213;
wire n_538;
wire n_2004;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_1936;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1961;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_1894;
wire n_1231;
wire n_1978;
wire n_2085;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_1815;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1967;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1911;
wire n_1956;
wire n_1644;
wire n_2011;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_1986;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_1918;
wire n_577;
wire n_1843;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1909;
wire n_2080;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_2093;
wire n_483;
wire n_1970;
wire n_608;
wire n_261;
wire n_630;
wire n_2059;
wire n_541;
wire n_512;
wire n_2073;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_1957;
wire n_219;
wire n_1907;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1876;
wire n_1895;
wire n_1697;
wire n_243;
wire n_979;
wire n_1873;
wire n_905;
wire n_1866;
wire n_1680;
wire n_322;
wire n_993;
wire n_689;
wire n_2031;
wire n_354;
wire n_1413;
wire n_1330;
wire n_1605;
wire n_1988;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_2009;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_2068;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_2072;
wire n_1354;
wire n_586;
wire n_423;
wire n_1875;
wire n_1865;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_1950;
wire n_530;
wire n_1563;
wire n_1912;
wire n_277;
wire n_1982;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_1927;
wire n_2028;
wire n_1069;
wire n_1722;
wire n_1664;
wire n_612;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_2008;
wire n_1926;
wire n_1175;
wire n_328;
wire n_1386;
wire n_1896;
wire n_429;
wire n_1747;
wire n_1012;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1977;
wire n_1802;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_928;
wire n_835;
wire n_1214;
wire n_690;
wire n_850;
wire n_1801;
wire n_1886;
wire n_2092;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_2096;
wire n_1965;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_697;
wire n_687;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_484;
wire n_2036;
wire n_1709;
wire n_1825;
wire n_1757;
wire n_1796;
wire n_1792;
wire n_891;
wire n_2067;
wire n_2082;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_2075;
wire n_1987;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_462;
wire n_1052;
wire n_1033;
wire n_1296;
wire n_1990;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_2078;
wire n_595;
wire n_297;
wire n_627;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1858;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_382;
wire n_673;
wire n_1969;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_1968;
wire n_898;
wire n_255;
wire n_284;
wire n_1952;
wire n_865;
wire n_925;
wire n_1932;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_1839;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_1863;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_1308;
wire n_2089;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_1913;
wire n_510;
wire n_837;
wire n_2097;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_1947;
wire n_536;
wire n_1788;
wire n_1999;
wire n_622;
wire n_1469;
wire n_2060;
wire n_1838;
wire n_1835;
wire n_1766;
wire n_1776;
wire n_1959;
wire n_2002;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_1878;
wire n_899;
wire n_738;
wire n_2012;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_2069;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_1181;
wire n_1822;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_1992;
wire n_648;
wire n_657;
wire n_1049;
wire n_2057;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_1817;
wire n_927;
wire n_1849;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_552;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_216;
wire n_912;
wire n_1857;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_1955;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_683;
wire n_527;
wire n_811;
wire n_1207;
wire n_312;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_1897;
wire n_2064;
wire n_880;
wire n_2053;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_1942;
wire n_1966;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_1837;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_2063;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_1483;
wire n_1834;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1993;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1919;
wire n_1080;
wire n_723;
wire n_1877;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1939;
wire n_2030;
wire n_1769;
wire n_1220;
wire n_1893;
wire n_556;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_2025;
wire n_1125;
wire n_970;
wire n_1980;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_1951;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_1286;
wire n_1773;
wire n_1775;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_1745;
wire n_914;
wire n_759;
wire n_1831;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_1901;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1892;
wire n_1933;
wire n_1135;
wire n_1179;
wire n_1169;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1917;
wire n_2000;
wire n_1580;
wire n_1425;
wire n_1881;
wire n_1281;
wire n_1267;
wire n_1806;
wire n_983;
wire n_2023;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_2087;
wire n_1855;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_1832;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_2049;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1995;
wire n_1594;
wire n_664;
wire n_1869;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_1889;
wire n_435;
wire n_1905;
wire n_2016;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_1937;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_575;
wire n_368;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1934;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_1871;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_1859;
wire n_238;
wire n_1095;
wire n_2024;
wire n_1595;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_1916;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_1847;
wire n_2052;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1841;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_1997;
wire n_340;
wire n_710;
wire n_1108;
wire n_1818;
wire n_1182;
wire n_1298;
wire n_2088;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1960;
wire n_2061;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1943;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1983;
wire n_1938;
wire n_1262;
wire n_218;
wire n_1891;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_239;
wire n_2037;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_1472;
wire n_2050;
wire n_1081;
wire n_402;
wire n_1870;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_2006;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_2017;
wire n_370;
wire n_1695;
wire n_1828;
wire n_2046;
wire n_650;
wire n_1046;
wire n_1940;
wire n_1979;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_1963;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1883;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_2084;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_1823;
wire n_227;
wire n_1974;
wire n_1720;
wire n_934;
wire n_482;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_1964;
wire n_1920;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_2007;
wire n_2039;
wire n_1946;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_1846;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_1676;
wire n_833;
wire n_1830;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_1900;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_2021;
wire n_1086;
wire n_1066;
wire n_1948;
wire n_2026;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1906;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_1758;
wire n_1925;
wire n_737;
wire n_1318;
wire n_1914;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_2056;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1984;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_1931;
wire n_2083;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_1941;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1962;
wire n_1559;
wire n_1725;
wire n_1928;
wire n_1872;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1746;
wire n_1325;
wire n_1002;
wire n_1741;
wire n_1949;
wire n_545;
wire n_489;
wire n_1804;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_2054;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_2062;
wire n_2041;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1860;
wire n_1904;
wire n_1200;
wire n_2070;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1908;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_2045;
wire n_817;
wire n_262;
wire n_897;
wire n_846;
wire n_2066;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1800;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1882;
wire n_1076;
wire n_1118;
wire n_1007;
wire n_1807;
wire n_1929;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_1879;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_680;
wire n_367;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_1953;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1976;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_2029;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_1810;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_2020;
wire n_1729;
wire n_669;
wire n_2048;
wire n_300;
wire n_222;
wire n_2005;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_2076;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1785;
wire n_763;
wire n_1147;
wire n_1848;
wire n_360;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_1994;
wire n_895;
wire n_866;
wire n_1227;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_1924;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_1174;
wire n_1944;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_2081;
wire n_234;
wire n_2022;
wire n_1945;
wire n_910;
wire n_1721;
wire n_1656;
wire n_1460;
wire n_911;
wire n_1464;
wire n_653;
wire n_236;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_2034;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_1922;
wire n_563;
wire n_2032;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_1973;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_2015;
wire n_390;
wire n_1148;
wire n_334;
wire n_1989;
wire n_1161;
wire n_1085;
wire n_232;
wire n_2014;
wire n_2042;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1972;
wire n_1525;
wire n_455;
wire n_1585;
wire n_1851;
wire n_363;
wire n_1799;
wire n_1090;
wire n_592;
wire n_1816;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_1829;
wire n_503;
wire n_2035;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_2033;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_2071;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_2010;
wire n_1651;
wire n_1198;
wire n_2047;
wire n_2095;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1998;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1981;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_1996;
wire n_249;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_2043;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1921;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_2065;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_271;
wire n_404;
wire n_2001;
wire n_1884;
wire n_2040;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1819;
wire n_2055;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_2038;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_373;
wire n_1632;
wire n_1890;
wire n_1805;
wire n_257;
wire n_1557;
wire n_1888;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_1850;
wire n_1898;
wire n_1868;
wire n_2079;
wire n_1089;
wire n_1887;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_1242;
wire n_2086;
wire n_1836;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1899;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1862;
wire n_1856;
wire n_1958;
wire n_2077;
wire n_339;
wire n_784;
wire n_434;
wire n_315;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_1423;
wire n_1935;
wire n_2027;
wire n_457;
wire n_2091;
wire n_364;
wire n_1915;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1885;
wire n_1013;
wire n_1259;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

INVx1_ASAP7_75t_L g212 ( 
.A(n_76),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_44),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_96),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_170),
.Y(n_215)
);

BUFx8_ASAP7_75t_SL g216 ( 
.A(n_194),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_12),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_95),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_176),
.Y(n_219)
);

INVxp67_ASAP7_75t_L g220 ( 
.A(n_23),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_46),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_193),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_168),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_164),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_100),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_104),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_33),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_149),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_137),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_129),
.Y(n_230)
);

BUFx10_ASAP7_75t_L g231 ( 
.A(n_157),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_87),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_10),
.Y(n_233)
);

BUFx6f_ASAP7_75t_L g234 ( 
.A(n_8),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_90),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_97),
.Y(n_236)
);

BUFx6f_ASAP7_75t_L g237 ( 
.A(n_22),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_159),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_21),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_143),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_116),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_22),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_0),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_88),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_108),
.Y(n_245)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_62),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_83),
.Y(n_247)
);

BUFx5_ASAP7_75t_L g248 ( 
.A(n_78),
.Y(n_248)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_40),
.Y(n_249)
);

BUFx10_ASAP7_75t_L g250 ( 
.A(n_148),
.Y(n_250)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_133),
.Y(n_251)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_39),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_37),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_101),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_66),
.Y(n_255)
);

INVxp67_ASAP7_75t_L g256 ( 
.A(n_167),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_171),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_177),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_131),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_158),
.Y(n_260)
);

BUFx10_ASAP7_75t_L g261 ( 
.A(n_32),
.Y(n_261)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_112),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_65),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_173),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_115),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_169),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_89),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_106),
.Y(n_268)
);

INVx1_ASAP7_75t_SL g269 ( 
.A(n_47),
.Y(n_269)
);

BUFx3_ASAP7_75t_L g270 ( 
.A(n_0),
.Y(n_270)
);

BUFx3_ASAP7_75t_L g271 ( 
.A(n_207),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_132),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_203),
.Y(n_273)
);

CKINVDCx16_ASAP7_75t_R g274 ( 
.A(n_183),
.Y(n_274)
);

BUFx3_ASAP7_75t_L g275 ( 
.A(n_27),
.Y(n_275)
);

BUFx2_ASAP7_75t_L g276 ( 
.A(n_206),
.Y(n_276)
);

INVx1_ASAP7_75t_SL g277 ( 
.A(n_210),
.Y(n_277)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_86),
.Y(n_278)
);

BUFx6f_ASAP7_75t_L g279 ( 
.A(n_40),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_59),
.Y(n_280)
);

INVxp67_ASAP7_75t_L g281 ( 
.A(n_47),
.Y(n_281)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_105),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_188),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_46),
.Y(n_284)
);

INVxp67_ASAP7_75t_L g285 ( 
.A(n_127),
.Y(n_285)
);

BUFx10_ASAP7_75t_L g286 ( 
.A(n_14),
.Y(n_286)
);

INVx1_ASAP7_75t_SL g287 ( 
.A(n_191),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_1),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_20),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_8),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_134),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_190),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_7),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_202),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_24),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_99),
.Y(n_296)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_64),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_181),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_165),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_80),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_120),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_156),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_43),
.Y(n_303)
);

CKINVDCx16_ASAP7_75t_R g304 ( 
.A(n_33),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_51),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_142),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_144),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_102),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_56),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_130),
.Y(n_310)
);

BUFx3_ASAP7_75t_L g311 ( 
.A(n_24),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_82),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_20),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_13),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_52),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_198),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_65),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_18),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_32),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_14),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_98),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_84),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_1),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_74),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_57),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_93),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_135),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_110),
.Y(n_328)
);

CKINVDCx16_ASAP7_75t_R g329 ( 
.A(n_53),
.Y(n_329)
);

CKINVDCx16_ASAP7_75t_R g330 ( 
.A(n_175),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_155),
.Y(n_331)
);

BUFx6f_ASAP7_75t_L g332 ( 
.A(n_51),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_182),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_211),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_28),
.Y(n_335)
);

BUFx3_ASAP7_75t_L g336 ( 
.A(n_54),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_39),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_66),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_25),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_208),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_146),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_5),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_117),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_166),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_62),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_45),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g347 ( 
.A(n_189),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_54),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_49),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_114),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_7),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_29),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_9),
.Y(n_353)
);

BUFx3_ASAP7_75t_L g354 ( 
.A(n_180),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_195),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_124),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_201),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_27),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_187),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g360 ( 
.A(n_125),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_2),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_186),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_209),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g364 ( 
.A(n_161),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_13),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_52),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_150),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_123),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_60),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_196),
.Y(n_370)
);

CKINVDCx16_ASAP7_75t_R g371 ( 
.A(n_11),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_126),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_147),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_73),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_151),
.Y(n_375)
);

CKINVDCx20_ASAP7_75t_R g376 ( 
.A(n_28),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_63),
.Y(n_377)
);

BUFx5_ASAP7_75t_L g378 ( 
.A(n_174),
.Y(n_378)
);

INVx1_ASAP7_75t_SL g379 ( 
.A(n_119),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_122),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_53),
.Y(n_381)
);

INVx2_ASAP7_75t_SL g382 ( 
.A(n_61),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_9),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_92),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_26),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_18),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_200),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_154),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_58),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_107),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_163),
.Y(n_391)
);

CKINVDCx20_ASAP7_75t_R g392 ( 
.A(n_36),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_60),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_178),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_59),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_3),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_121),
.Y(n_397)
);

INVx2_ASAP7_75t_L g398 ( 
.A(n_68),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_38),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_34),
.Y(n_400)
);

HB1xp67_ASAP7_75t_L g401 ( 
.A(n_153),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_75),
.Y(n_402)
);

INVx1_ASAP7_75t_SL g403 ( 
.A(n_192),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_71),
.Y(n_404)
);

INVx2_ASAP7_75t_L g405 ( 
.A(n_58),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_10),
.Y(n_406)
);

BUFx2_ASAP7_75t_SL g407 ( 
.A(n_30),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_55),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_138),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_140),
.Y(n_410)
);

CKINVDCx16_ASAP7_75t_R g411 ( 
.A(n_128),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_77),
.Y(n_412)
);

BUFx2_ASAP7_75t_L g413 ( 
.A(n_37),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_42),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_139),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_34),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_35),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_35),
.Y(n_418)
);

BUFx2_ASAP7_75t_L g419 ( 
.A(n_91),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_234),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_L g421 ( 
.A(n_276),
.B(n_419),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_234),
.Y(n_422)
);

NOR2xp33_ASAP7_75t_L g423 ( 
.A(n_401),
.B(n_2),
.Y(n_423)
);

CKINVDCx20_ASAP7_75t_R g424 ( 
.A(n_218),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_304),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_329),
.Y(n_426)
);

NOR2xp33_ASAP7_75t_L g427 ( 
.A(n_256),
.B(n_3),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_371),
.Y(n_428)
);

CKINVDCx20_ASAP7_75t_R g429 ( 
.A(n_347),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_263),
.Y(n_430)
);

CKINVDCx20_ASAP7_75t_R g431 ( 
.A(n_360),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_280),
.Y(n_432)
);

CKINVDCx20_ASAP7_75t_R g433 ( 
.A(n_364),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_270),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_270),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_293),
.Y(n_436)
);

BUFx2_ASAP7_75t_L g437 ( 
.A(n_413),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_275),
.Y(n_438)
);

CKINVDCx16_ASAP7_75t_R g439 ( 
.A(n_274),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_295),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_275),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_303),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_305),
.Y(n_443)
);

HB1xp67_ASAP7_75t_L g444 ( 
.A(n_217),
.Y(n_444)
);

AND2x2_ASAP7_75t_L g445 ( 
.A(n_311),
.B(n_4),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_234),
.Y(n_446)
);

INVx2_ASAP7_75t_L g447 ( 
.A(n_234),
.Y(n_447)
);

BUFx2_ASAP7_75t_SL g448 ( 
.A(n_382),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_234),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_319),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_320),
.Y(n_451)
);

CKINVDCx20_ASAP7_75t_R g452 ( 
.A(n_216),
.Y(n_452)
);

CKINVDCx20_ASAP7_75t_R g453 ( 
.A(n_330),
.Y(n_453)
);

CKINVDCx20_ASAP7_75t_R g454 ( 
.A(n_411),
.Y(n_454)
);

BUFx3_ASAP7_75t_L g455 ( 
.A(n_271),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_251),
.B(n_4),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_311),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_336),
.Y(n_458)
);

NOR2xp33_ASAP7_75t_R g459 ( 
.A(n_260),
.B(n_205),
.Y(n_459)
);

NOR2xp67_ASAP7_75t_L g460 ( 
.A(n_220),
.B(n_5),
.Y(n_460)
);

CKINVDCx20_ASAP7_75t_R g461 ( 
.A(n_264),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_336),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_237),
.Y(n_463)
);

CKINVDCx5p33_ASAP7_75t_R g464 ( 
.A(n_323),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_237),
.Y(n_465)
);

CKINVDCx20_ASAP7_75t_R g466 ( 
.A(n_266),
.Y(n_466)
);

CKINVDCx5p33_ASAP7_75t_R g467 ( 
.A(n_335),
.Y(n_467)
);

CKINVDCx20_ASAP7_75t_R g468 ( 
.A(n_268),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_237),
.Y(n_469)
);

INVxp33_ASAP7_75t_SL g470 ( 
.A(n_217),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_251),
.B(n_6),
.Y(n_471)
);

INVxp67_ASAP7_75t_SL g472 ( 
.A(n_271),
.Y(n_472)
);

HB1xp67_ASAP7_75t_L g473 ( 
.A(n_221),
.Y(n_473)
);

CKINVDCx20_ASAP7_75t_R g474 ( 
.A(n_283),
.Y(n_474)
);

CKINVDCx5p33_ASAP7_75t_R g475 ( 
.A(n_338),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_237),
.Y(n_476)
);

NOR2xp33_ASAP7_75t_L g477 ( 
.A(n_285),
.B(n_6),
.Y(n_477)
);

INVx2_ASAP7_75t_L g478 ( 
.A(n_237),
.Y(n_478)
);

CKINVDCx20_ASAP7_75t_R g479 ( 
.A(n_292),
.Y(n_479)
);

CKINVDCx20_ASAP7_75t_R g480 ( 
.A(n_298),
.Y(n_480)
);

INVx2_ASAP7_75t_L g481 ( 
.A(n_279),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_279),
.Y(n_482)
);

NOR2xp67_ASAP7_75t_L g483 ( 
.A(n_281),
.B(n_11),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_262),
.B(n_12),
.Y(n_484)
);

CKINVDCx20_ASAP7_75t_R g485 ( 
.A(n_299),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_279),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_279),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_279),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_332),
.Y(n_489)
);

INVxp67_ASAP7_75t_SL g490 ( 
.A(n_354),
.Y(n_490)
);

CKINVDCx5p33_ASAP7_75t_R g491 ( 
.A(n_342),
.Y(n_491)
);

CKINVDCx5p33_ASAP7_75t_R g492 ( 
.A(n_345),
.Y(n_492)
);

INVx2_ASAP7_75t_L g493 ( 
.A(n_332),
.Y(n_493)
);

INVxp67_ASAP7_75t_L g494 ( 
.A(n_261),
.Y(n_494)
);

CKINVDCx20_ASAP7_75t_R g495 ( 
.A(n_300),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_332),
.Y(n_496)
);

CKINVDCx5p33_ASAP7_75t_R g497 ( 
.A(n_346),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_332),
.Y(n_498)
);

CKINVDCx16_ASAP7_75t_R g499 ( 
.A(n_261),
.Y(n_499)
);

BUFx6f_ASAP7_75t_SL g500 ( 
.A(n_231),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_332),
.Y(n_501)
);

INVxp67_ASAP7_75t_L g502 ( 
.A(n_261),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_213),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_284),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_288),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_289),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_290),
.Y(n_507)
);

CKINVDCx20_ASAP7_75t_R g508 ( 
.A(n_301),
.Y(n_508)
);

CKINVDCx20_ASAP7_75t_R g509 ( 
.A(n_308),
.Y(n_509)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_248),
.Y(n_510)
);

CKINVDCx5p33_ASAP7_75t_R g511 ( 
.A(n_348),
.Y(n_511)
);

CKINVDCx5p33_ASAP7_75t_R g512 ( 
.A(n_349),
.Y(n_512)
);

CKINVDCx5p33_ASAP7_75t_R g513 ( 
.A(n_351),
.Y(n_513)
);

BUFx2_ASAP7_75t_L g514 ( 
.A(n_221),
.Y(n_514)
);

BUFx2_ASAP7_75t_L g515 ( 
.A(n_227),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_313),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_246),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_246),
.Y(n_518)
);

CKINVDCx5p33_ASAP7_75t_R g519 ( 
.A(n_352),
.Y(n_519)
);

NOR2xp67_ASAP7_75t_L g520 ( 
.A(n_382),
.B(n_15),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_249),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_249),
.Y(n_522)
);

CKINVDCx20_ASAP7_75t_R g523 ( 
.A(n_322),
.Y(n_523)
);

NOR2xp33_ASAP7_75t_L g524 ( 
.A(n_262),
.B(n_15),
.Y(n_524)
);

CKINVDCx16_ASAP7_75t_R g525 ( 
.A(n_286),
.Y(n_525)
);

CKINVDCx5p33_ASAP7_75t_R g526 ( 
.A(n_353),
.Y(n_526)
);

CKINVDCx5p33_ASAP7_75t_R g527 ( 
.A(n_361),
.Y(n_527)
);

CKINVDCx20_ASAP7_75t_R g528 ( 
.A(n_424),
.Y(n_528)
);

CKINVDCx5p33_ASAP7_75t_R g529 ( 
.A(n_452),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_420),
.Y(n_530)
);

INVx3_ASAP7_75t_L g531 ( 
.A(n_447),
.Y(n_531)
);

INVx3_ASAP7_75t_L g532 ( 
.A(n_447),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_420),
.Y(n_533)
);

OA21x2_ASAP7_75t_L g534 ( 
.A1(n_456),
.A2(n_282),
.B(n_278),
.Y(n_534)
);

NOR2xp33_ASAP7_75t_L g535 ( 
.A(n_421),
.B(n_277),
.Y(n_535)
);

CKINVDCx5p33_ASAP7_75t_R g536 ( 
.A(n_461),
.Y(n_536)
);

NAND2x1_ASAP7_75t_L g537 ( 
.A(n_422),
.B(n_278),
.Y(n_537)
);

CKINVDCx20_ASAP7_75t_R g538 ( 
.A(n_429),
.Y(n_538)
);

AND2x2_ASAP7_75t_L g539 ( 
.A(n_472),
.B(n_252),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_422),
.Y(n_540)
);

CKINVDCx5p33_ASAP7_75t_R g541 ( 
.A(n_466),
.Y(n_541)
);

BUFx6f_ASAP7_75t_L g542 ( 
.A(n_478),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_446),
.Y(n_543)
);

BUFx6f_ASAP7_75t_L g544 ( 
.A(n_478),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_446),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_449),
.Y(n_546)
);

AND2x4_ASAP7_75t_L g547 ( 
.A(n_445),
.B(n_354),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_SL g548 ( 
.A(n_439),
.B(n_231),
.Y(n_548)
);

INVx2_ASAP7_75t_L g549 ( 
.A(n_481),
.Y(n_549)
);

CKINVDCx20_ASAP7_75t_R g550 ( 
.A(n_431),
.Y(n_550)
);

BUFx10_ASAP7_75t_L g551 ( 
.A(n_500),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_449),
.Y(n_552)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_481),
.Y(n_553)
);

BUFx2_ASAP7_75t_L g554 ( 
.A(n_425),
.Y(n_554)
);

OA21x2_ASAP7_75t_L g555 ( 
.A1(n_471),
.A2(n_282),
.B(n_224),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_L g556 ( 
.A(n_490),
.B(n_212),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_493),
.Y(n_557)
);

INVx4_ASAP7_75t_L g558 ( 
.A(n_510),
.Y(n_558)
);

INVx2_ASAP7_75t_L g559 ( 
.A(n_493),
.Y(n_559)
);

CKINVDCx5p33_ASAP7_75t_R g560 ( 
.A(n_468),
.Y(n_560)
);

CKINVDCx20_ASAP7_75t_R g561 ( 
.A(n_433),
.Y(n_561)
);

CKINVDCx5p33_ASAP7_75t_R g562 ( 
.A(n_474),
.Y(n_562)
);

BUFx8_ASAP7_75t_L g563 ( 
.A(n_500),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_L g564 ( 
.A(n_455),
.B(n_240),
.Y(n_564)
);

HB1xp67_ASAP7_75t_L g565 ( 
.A(n_425),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_463),
.Y(n_566)
);

INVx3_ASAP7_75t_L g567 ( 
.A(n_510),
.Y(n_567)
);

CKINVDCx20_ASAP7_75t_R g568 ( 
.A(n_479),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_SL g569 ( 
.A(n_499),
.B(n_231),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_465),
.Y(n_570)
);

CKINVDCx5p33_ASAP7_75t_R g571 ( 
.A(n_480),
.Y(n_571)
);

CKINVDCx20_ASAP7_75t_R g572 ( 
.A(n_485),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_469),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_476),
.Y(n_574)
);

INVx3_ASAP7_75t_L g575 ( 
.A(n_482),
.Y(n_575)
);

AND2x4_ASAP7_75t_L g576 ( 
.A(n_445),
.B(n_247),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_486),
.Y(n_577)
);

AND2x4_ASAP7_75t_L g578 ( 
.A(n_487),
.B(n_488),
.Y(n_578)
);

INVx3_ASAP7_75t_L g579 ( 
.A(n_489),
.Y(n_579)
);

INVx2_ASAP7_75t_L g580 ( 
.A(n_496),
.Y(n_580)
);

INVx2_ASAP7_75t_L g581 ( 
.A(n_498),
.Y(n_581)
);

CKINVDCx5p33_ASAP7_75t_R g582 ( 
.A(n_495),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_501),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_517),
.Y(n_584)
);

NOR2xp33_ASAP7_75t_R g585 ( 
.A(n_508),
.B(n_327),
.Y(n_585)
);

CKINVDCx5p33_ASAP7_75t_R g586 ( 
.A(n_509),
.Y(n_586)
);

CKINVDCx20_ASAP7_75t_R g587 ( 
.A(n_523),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_517),
.Y(n_588)
);

CKINVDCx5p33_ASAP7_75t_R g589 ( 
.A(n_430),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_518),
.Y(n_590)
);

CKINVDCx5p33_ASAP7_75t_R g591 ( 
.A(n_430),
.Y(n_591)
);

CKINVDCx5p33_ASAP7_75t_R g592 ( 
.A(n_432),
.Y(n_592)
);

CKINVDCx5p33_ASAP7_75t_R g593 ( 
.A(n_432),
.Y(n_593)
);

HB1xp67_ASAP7_75t_L g594 ( 
.A(n_426),
.Y(n_594)
);

CKINVDCx5p33_ASAP7_75t_R g595 ( 
.A(n_436),
.Y(n_595)
);

INVx2_ASAP7_75t_L g596 ( 
.A(n_518),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_521),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_521),
.Y(n_598)
);

CKINVDCx5p33_ASAP7_75t_R g599 ( 
.A(n_436),
.Y(n_599)
);

CKINVDCx5p33_ASAP7_75t_R g600 ( 
.A(n_440),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_522),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_522),
.Y(n_602)
);

BUFx6f_ASAP7_75t_L g603 ( 
.A(n_484),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_503),
.Y(n_604)
);

CKINVDCx5p33_ASAP7_75t_R g605 ( 
.A(n_440),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g606 ( 
.A(n_455),
.B(n_265),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_L g607 ( 
.A(n_434),
.B(n_267),
.Y(n_607)
);

AND2x4_ASAP7_75t_L g608 ( 
.A(n_435),
.B(n_272),
.Y(n_608)
);

BUFx6f_ASAP7_75t_L g609 ( 
.A(n_504),
.Y(n_609)
);

CKINVDCx5p33_ASAP7_75t_R g610 ( 
.A(n_442),
.Y(n_610)
);

INVx3_ASAP7_75t_L g611 ( 
.A(n_505),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_506),
.Y(n_612)
);

INVx2_ASAP7_75t_L g613 ( 
.A(n_507),
.Y(n_613)
);

NAND3xp33_ASAP7_75t_L g614 ( 
.A(n_535),
.B(n_423),
.C(n_442),
.Y(n_614)
);

AND2x4_ASAP7_75t_L g615 ( 
.A(n_547),
.B(n_516),
.Y(n_615)
);

INVx3_ASAP7_75t_L g616 ( 
.A(n_558),
.Y(n_616)
);

AND2x4_ASAP7_75t_L g617 ( 
.A(n_547),
.B(n_438),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_603),
.B(n_443),
.Y(n_618)
);

NOR2xp33_ASAP7_75t_L g619 ( 
.A(n_556),
.B(n_470),
.Y(n_619)
);

BUFx3_ASAP7_75t_L g620 ( 
.A(n_603),
.Y(n_620)
);

BUFx3_ASAP7_75t_L g621 ( 
.A(n_603),
.Y(n_621)
);

INVx2_ASAP7_75t_L g622 ( 
.A(n_549),
.Y(n_622)
);

NOR2xp33_ASAP7_75t_L g623 ( 
.A(n_548),
.B(n_443),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_SL g624 ( 
.A(n_551),
.B(n_525),
.Y(n_624)
);

INVx3_ASAP7_75t_L g625 ( 
.A(n_558),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_L g626 ( 
.A(n_603),
.B(n_450),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_604),
.Y(n_627)
);

INVx3_ASAP7_75t_L g628 ( 
.A(n_558),
.Y(n_628)
);

INVx4_ASAP7_75t_L g629 ( 
.A(n_558),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_L g630 ( 
.A(n_603),
.B(n_450),
.Y(n_630)
);

INVx2_ASAP7_75t_L g631 ( 
.A(n_549),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_578),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_SL g633 ( 
.A(n_551),
.B(n_451),
.Y(n_633)
);

INVx4_ASAP7_75t_L g634 ( 
.A(n_603),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_L g635 ( 
.A(n_547),
.B(n_451),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_L g636 ( 
.A(n_547),
.B(n_464),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_SL g637 ( 
.A(n_551),
.B(n_464),
.Y(n_637)
);

AND2x2_ASAP7_75t_L g638 ( 
.A(n_539),
.B(n_448),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_L g639 ( 
.A(n_576),
.B(n_467),
.Y(n_639)
);

BUFx10_ASAP7_75t_L g640 ( 
.A(n_589),
.Y(n_640)
);

INVx2_ASAP7_75t_L g641 ( 
.A(n_553),
.Y(n_641)
);

AOI22xp33_ASAP7_75t_L g642 ( 
.A1(n_576),
.A2(n_524),
.B1(n_437),
.B2(n_477),
.Y(n_642)
);

AND2x6_ASAP7_75t_L g643 ( 
.A(n_576),
.B(n_273),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_L g644 ( 
.A(n_576),
.B(n_467),
.Y(n_644)
);

NOR2xp33_ASAP7_75t_L g645 ( 
.A(n_591),
.B(n_475),
.Y(n_645)
);

INVx3_ASAP7_75t_L g646 ( 
.A(n_567),
.Y(n_646)
);

OR2x2_ASAP7_75t_L g647 ( 
.A(n_564),
.B(n_514),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_578),
.Y(n_648)
);

BUFx10_ASAP7_75t_L g649 ( 
.A(n_592),
.Y(n_649)
);

INVx2_ASAP7_75t_L g650 ( 
.A(n_553),
.Y(n_650)
);

NOR2xp33_ASAP7_75t_L g651 ( 
.A(n_593),
.B(n_475),
.Y(n_651)
);

AND2x4_ASAP7_75t_L g652 ( 
.A(n_608),
.B(n_539),
.Y(n_652)
);

INVx2_ASAP7_75t_SL g653 ( 
.A(n_608),
.Y(n_653)
);

NOR2xp33_ASAP7_75t_L g654 ( 
.A(n_595),
.B(n_491),
.Y(n_654)
);

OR2x2_ASAP7_75t_L g655 ( 
.A(n_606),
.B(n_514),
.Y(n_655)
);

AND2x4_ASAP7_75t_L g656 ( 
.A(n_608),
.B(n_441),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_604),
.Y(n_657)
);

NOR2x1p5_ASAP7_75t_L g658 ( 
.A(n_599),
.B(n_426),
.Y(n_658)
);

BUFx6f_ASAP7_75t_L g659 ( 
.A(n_609),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_SL g660 ( 
.A(n_551),
.B(n_491),
.Y(n_660)
);

CKINVDCx5p33_ASAP7_75t_R g661 ( 
.A(n_585),
.Y(n_661)
);

AND2x2_ASAP7_75t_SL g662 ( 
.A(n_555),
.B(n_427),
.Y(n_662)
);

INVx5_ASAP7_75t_L g663 ( 
.A(n_567),
.Y(n_663)
);

INVx2_ASAP7_75t_L g664 ( 
.A(n_559),
.Y(n_664)
);

OR2x2_ASAP7_75t_L g665 ( 
.A(n_554),
.B(n_515),
.Y(n_665)
);

INVx4_ASAP7_75t_L g666 ( 
.A(n_542),
.Y(n_666)
);

AND2x2_ASAP7_75t_L g667 ( 
.A(n_608),
.B(n_448),
.Y(n_667)
);

INVxp67_ASAP7_75t_SL g668 ( 
.A(n_567),
.Y(n_668)
);

AND2x4_ASAP7_75t_L g669 ( 
.A(n_612),
.B(n_457),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_578),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_578),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_SL g672 ( 
.A(n_563),
.B(n_492),
.Y(n_672)
);

NAND2xp33_ASAP7_75t_R g673 ( 
.A(n_600),
.B(n_428),
.Y(n_673)
);

OAI22xp33_ASAP7_75t_L g674 ( 
.A1(n_569),
.A2(n_269),
.B1(n_520),
.B2(n_437),
.Y(n_674)
);

NOR2x1p5_ASAP7_75t_L g675 ( 
.A(n_605),
.B(n_428),
.Y(n_675)
);

BUFx3_ASAP7_75t_L g676 ( 
.A(n_537),
.Y(n_676)
);

INVx2_ASAP7_75t_SL g677 ( 
.A(n_555),
.Y(n_677)
);

BUFx3_ASAP7_75t_L g678 ( 
.A(n_537),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_L g679 ( 
.A(n_530),
.B(n_533),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_612),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_L g681 ( 
.A(n_530),
.B(n_492),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_611),
.Y(n_682)
);

INVx5_ASAP7_75t_L g683 ( 
.A(n_567),
.Y(n_683)
);

INVx4_ASAP7_75t_L g684 ( 
.A(n_542),
.Y(n_684)
);

CKINVDCx5p33_ASAP7_75t_R g685 ( 
.A(n_536),
.Y(n_685)
);

BUFx2_ASAP7_75t_L g686 ( 
.A(n_554),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_SL g687 ( 
.A(n_563),
.B(n_497),
.Y(n_687)
);

OAI22xp33_ASAP7_75t_L g688 ( 
.A1(n_607),
.A2(n_460),
.B1(n_483),
.B2(n_369),
.Y(n_688)
);

OAI22xp5_ASAP7_75t_L g689 ( 
.A1(n_610),
.A2(n_453),
.B1(n_454),
.B2(n_519),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_533),
.B(n_497),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_L g691 ( 
.A(n_540),
.B(n_511),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_L g692 ( 
.A(n_540),
.B(n_543),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_L g693 ( 
.A(n_543),
.B(n_511),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_611),
.Y(n_694)
);

INVx2_ASAP7_75t_SL g695 ( 
.A(n_555),
.Y(n_695)
);

AND3x2_ASAP7_75t_L g696 ( 
.A(n_565),
.B(n_297),
.C(n_252),
.Y(n_696)
);

INVx3_ASAP7_75t_L g697 ( 
.A(n_542),
.Y(n_697)
);

XOR2xp5_ASAP7_75t_L g698 ( 
.A(n_528),
.B(n_538),
.Y(n_698)
);

AOI22xp33_ASAP7_75t_L g699 ( 
.A1(n_555),
.A2(n_297),
.B1(n_398),
.B2(n_405),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_611),
.Y(n_700)
);

INVx3_ASAP7_75t_L g701 ( 
.A(n_542),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_L g702 ( 
.A(n_545),
.B(n_512),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_L g703 ( 
.A(n_545),
.B(n_512),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_L g704 ( 
.A(n_546),
.B(n_513),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_611),
.Y(n_705)
);

INVx3_ASAP7_75t_L g706 ( 
.A(n_542),
.Y(n_706)
);

HB1xp67_ASAP7_75t_L g707 ( 
.A(n_594),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_546),
.Y(n_708)
);

INVx2_ASAP7_75t_L g709 ( 
.A(n_559),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_L g710 ( 
.A(n_552),
.B(n_513),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_552),
.Y(n_711)
);

NOR2x1p5_ASAP7_75t_L g712 ( 
.A(n_563),
.B(n_519),
.Y(n_712)
);

INVxp33_ASAP7_75t_SL g713 ( 
.A(n_541),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_566),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_566),
.Y(n_715)
);

AND2x2_ASAP7_75t_L g716 ( 
.A(n_584),
.B(n_458),
.Y(n_716)
);

BUFx3_ASAP7_75t_L g717 ( 
.A(n_609),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_570),
.Y(n_718)
);

BUFx3_ASAP7_75t_L g719 ( 
.A(n_609),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_570),
.B(n_526),
.Y(n_720)
);

INVx1_ASAP7_75t_SL g721 ( 
.A(n_568),
.Y(n_721)
);

INVx2_ASAP7_75t_L g722 ( 
.A(n_580),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_SL g723 ( 
.A(n_563),
.B(n_526),
.Y(n_723)
);

INVx2_ASAP7_75t_L g724 ( 
.A(n_580),
.Y(n_724)
);

OAI22xp5_ASAP7_75t_L g725 ( 
.A1(n_613),
.A2(n_527),
.B1(n_502),
.B2(n_494),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_L g726 ( 
.A(n_573),
.B(n_527),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_SL g727 ( 
.A(n_609),
.B(n_515),
.Y(n_727)
);

AOI22xp33_ASAP7_75t_L g728 ( 
.A1(n_534),
.A2(n_405),
.B1(n_398),
.B2(n_609),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_573),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_574),
.Y(n_730)
);

BUFx6f_ASAP7_75t_L g731 ( 
.A(n_609),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_574),
.Y(n_732)
);

OAI22xp5_ASAP7_75t_L g733 ( 
.A1(n_613),
.A2(n_473),
.B1(n_444),
.B2(n_403),
.Y(n_733)
);

AND3x2_ASAP7_75t_L g734 ( 
.A(n_584),
.B(n_294),
.C(n_291),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_SL g735 ( 
.A(n_560),
.B(n_459),
.Y(n_735)
);

AOI22xp5_ASAP7_75t_L g736 ( 
.A1(n_534),
.A2(n_500),
.B1(n_215),
.B2(n_219),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_577),
.Y(n_737)
);

INVx2_ASAP7_75t_L g738 ( 
.A(n_581),
.Y(n_738)
);

CKINVDCx20_ASAP7_75t_R g739 ( 
.A(n_550),
.Y(n_739)
);

INVx1_ASAP7_75t_SL g740 ( 
.A(n_572),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_SL g741 ( 
.A(n_562),
.B(n_250),
.Y(n_741)
);

OAI21xp33_ASAP7_75t_SL g742 ( 
.A1(n_588),
.A2(n_317),
.B(n_315),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_L g743 ( 
.A(n_577),
.B(n_287),
.Y(n_743)
);

BUFx8_ASAP7_75t_SL g744 ( 
.A(n_561),
.Y(n_744)
);

AOI22xp33_ASAP7_75t_L g745 ( 
.A1(n_534),
.A2(n_337),
.B1(n_418),
.B2(n_417),
.Y(n_745)
);

INVx3_ASAP7_75t_L g746 ( 
.A(n_542),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_583),
.Y(n_747)
);

INVx2_ASAP7_75t_SL g748 ( 
.A(n_534),
.Y(n_748)
);

INVx2_ASAP7_75t_L g749 ( 
.A(n_581),
.Y(n_749)
);

INVx2_ASAP7_75t_L g750 ( 
.A(n_557),
.Y(n_750)
);

NAND2x1p5_ASAP7_75t_L g751 ( 
.A(n_575),
.B(n_296),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_583),
.Y(n_752)
);

AND2x2_ASAP7_75t_L g753 ( 
.A(n_588),
.B(n_462),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_575),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_575),
.Y(n_755)
);

OR2x6_ASAP7_75t_L g756 ( 
.A(n_596),
.B(n_407),
.Y(n_756)
);

INVx4_ASAP7_75t_L g757 ( 
.A(n_544),
.Y(n_757)
);

INVx2_ASAP7_75t_L g758 ( 
.A(n_557),
.Y(n_758)
);

INVx3_ASAP7_75t_L g759 ( 
.A(n_544),
.Y(n_759)
);

NOR2xp33_ASAP7_75t_L g760 ( 
.A(n_590),
.B(n_379),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_575),
.B(n_328),
.Y(n_761)
);

BUFx3_ASAP7_75t_L g762 ( 
.A(n_544),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_SL g763 ( 
.A(n_571),
.B(n_250),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_SL g764 ( 
.A(n_582),
.B(n_250),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_579),
.Y(n_765)
);

INVx3_ASAP7_75t_L g766 ( 
.A(n_544),
.Y(n_766)
);

NOR2xp33_ASAP7_75t_L g767 ( 
.A(n_619),
.B(n_214),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_L g768 ( 
.A(n_616),
.B(n_579),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_L g769 ( 
.A(n_616),
.B(n_579),
.Y(n_769)
);

INVx2_ASAP7_75t_L g770 ( 
.A(n_750),
.Y(n_770)
);

INVx5_ASAP7_75t_L g771 ( 
.A(n_643),
.Y(n_771)
);

AOI21xp5_ASAP7_75t_L g772 ( 
.A1(n_616),
.A2(n_544),
.B(n_579),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_632),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_L g774 ( 
.A(n_625),
.B(n_544),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_625),
.B(n_302),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_625),
.B(n_306),
.Y(n_776)
);

CKINVDCx5p33_ASAP7_75t_R g777 ( 
.A(n_661),
.Y(n_777)
);

AND2x6_ASAP7_75t_L g778 ( 
.A(n_736),
.B(n_307),
.Y(n_778)
);

INVx2_ASAP7_75t_L g779 ( 
.A(n_750),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_628),
.B(n_310),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_628),
.B(n_312),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_632),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_648),
.Y(n_783)
);

INVx3_ASAP7_75t_L g784 ( 
.A(n_676),
.Y(n_784)
);

NAND3xp33_ASAP7_75t_L g785 ( 
.A(n_614),
.B(n_586),
.C(n_215),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_L g786 ( 
.A(n_628),
.B(n_321),
.Y(n_786)
);

INVx2_ASAP7_75t_L g787 ( 
.A(n_758),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_SL g788 ( 
.A(n_638),
.B(n_214),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_638),
.B(n_620),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_648),
.Y(n_790)
);

AOI22xp33_ASAP7_75t_L g791 ( 
.A1(n_662),
.A2(n_699),
.B1(n_745),
.B2(n_695),
.Y(n_791)
);

OAI22xp5_ASAP7_75t_L g792 ( 
.A1(n_618),
.A2(n_326),
.B1(n_324),
.B2(n_331),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_SL g793 ( 
.A(n_626),
.B(n_219),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_L g794 ( 
.A(n_620),
.B(n_340),
.Y(n_794)
);

OAI22xp33_ASAP7_75t_L g795 ( 
.A1(n_630),
.A2(n_359),
.B1(n_363),
.B2(n_368),
.Y(n_795)
);

NAND2x1_ASAP7_75t_L g796 ( 
.A(n_634),
.B(n_531),
.Y(n_796)
);

HB1xp67_ASAP7_75t_L g797 ( 
.A(n_686),
.Y(n_797)
);

NOR2xp33_ASAP7_75t_L g798 ( 
.A(n_647),
.B(n_222),
.Y(n_798)
);

A2O1A1Ixp33_ASAP7_75t_L g799 ( 
.A1(n_652),
.A2(n_394),
.B(n_391),
.C(n_374),
.Y(n_799)
);

INVxp67_ASAP7_75t_L g800 ( 
.A(n_665),
.Y(n_800)
);

NOR2xp67_ASAP7_75t_L g801 ( 
.A(n_661),
.B(n_645),
.Y(n_801)
);

AOI22xp33_ASAP7_75t_L g802 ( 
.A1(n_662),
.A2(n_365),
.B1(n_377),
.B2(n_386),
.Y(n_802)
);

INVx2_ASAP7_75t_L g803 ( 
.A(n_758),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_670),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_670),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_L g806 ( 
.A(n_621),
.B(n_370),
.Y(n_806)
);

AND2x2_ASAP7_75t_L g807 ( 
.A(n_667),
.B(n_587),
.Y(n_807)
);

NOR2xp33_ASAP7_75t_L g808 ( 
.A(n_647),
.B(n_222),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_L g809 ( 
.A(n_621),
.B(n_531),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_671),
.Y(n_810)
);

INVx3_ASAP7_75t_L g811 ( 
.A(n_676),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_L g812 ( 
.A(n_652),
.B(n_531),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_SL g813 ( 
.A(n_667),
.B(n_223),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_L g814 ( 
.A(n_652),
.B(n_531),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_L g815 ( 
.A(n_634),
.B(n_532),
.Y(n_815)
);

INVxp67_ASAP7_75t_SL g816 ( 
.A(n_646),
.Y(n_816)
);

HB1xp67_ASAP7_75t_L g817 ( 
.A(n_686),
.Y(n_817)
);

INVx2_ASAP7_75t_L g818 ( 
.A(n_622),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_L g819 ( 
.A(n_634),
.B(n_532),
.Y(n_819)
);

INVx2_ASAP7_75t_L g820 ( 
.A(n_622),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_671),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_SL g822 ( 
.A(n_635),
.B(n_223),
.Y(n_822)
);

INVxp67_ASAP7_75t_L g823 ( 
.A(n_665),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_SL g824 ( 
.A(n_636),
.B(n_225),
.Y(n_824)
);

INVxp33_ASAP7_75t_L g825 ( 
.A(n_698),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_627),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_L g827 ( 
.A(n_653),
.B(n_532),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_L g828 ( 
.A(n_653),
.B(n_532),
.Y(n_828)
);

BUFx6f_ASAP7_75t_L g829 ( 
.A(n_678),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_L g830 ( 
.A(n_668),
.B(n_596),
.Y(n_830)
);

AOI22xp5_ASAP7_75t_L g831 ( 
.A1(n_617),
.A2(n_615),
.B1(n_644),
.B2(n_639),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_SL g832 ( 
.A(n_682),
.B(n_248),
.Y(n_832)
);

AOI22xp33_ASAP7_75t_L g833 ( 
.A1(n_677),
.A2(n_339),
.B1(n_416),
.B2(n_414),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_657),
.Y(n_834)
);

INVx2_ASAP7_75t_L g835 ( 
.A(n_631),
.Y(n_835)
);

INVxp67_ASAP7_75t_L g836 ( 
.A(n_655),
.Y(n_836)
);

AOI22xp5_ASAP7_75t_L g837 ( 
.A1(n_617),
.A2(n_615),
.B1(n_623),
.B2(n_656),
.Y(n_837)
);

NOR2xp33_ASAP7_75t_L g838 ( 
.A(n_655),
.B(n_225),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_L g839 ( 
.A(n_629),
.B(n_590),
.Y(n_839)
);

AOI22xp5_ASAP7_75t_L g840 ( 
.A1(n_617),
.A2(n_350),
.B1(n_333),
.B2(n_334),
.Y(n_840)
);

NOR2x1p5_ASAP7_75t_L g841 ( 
.A(n_681),
.B(n_529),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_680),
.Y(n_842)
);

CKINVDCx5p33_ASAP7_75t_R g843 ( 
.A(n_744),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_L g844 ( 
.A(n_629),
.B(n_597),
.Y(n_844)
);

NOR2xp33_ASAP7_75t_L g845 ( 
.A(n_690),
.B(n_226),
.Y(n_845)
);

INVxp33_ASAP7_75t_L g846 ( 
.A(n_698),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_L g847 ( 
.A(n_629),
.B(n_597),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_L g848 ( 
.A(n_708),
.B(n_598),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_SL g849 ( 
.A(n_674),
.B(n_226),
.Y(n_849)
);

CKINVDCx20_ASAP7_75t_R g850 ( 
.A(n_739),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_716),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_L g852 ( 
.A(n_708),
.B(n_598),
.Y(n_852)
);

BUFx3_ASAP7_75t_L g853 ( 
.A(n_615),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_711),
.B(n_682),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_L g855 ( 
.A(n_711),
.B(n_601),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_L g856 ( 
.A(n_694),
.B(n_601),
.Y(n_856)
);

INVx2_ASAP7_75t_L g857 ( 
.A(n_631),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_SL g858 ( 
.A(n_694),
.B(n_248),
.Y(n_858)
);

INVx2_ASAP7_75t_SL g859 ( 
.A(n_656),
.Y(n_859)
);

OAI22xp33_ASAP7_75t_L g860 ( 
.A1(n_756),
.A2(n_392),
.B1(n_242),
.B2(n_309),
.Y(n_860)
);

INVxp67_ASAP7_75t_L g861 ( 
.A(n_707),
.Y(n_861)
);

BUFx5_ASAP7_75t_L g862 ( 
.A(n_643),
.Y(n_862)
);

HB1xp67_ASAP7_75t_L g863 ( 
.A(n_756),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_700),
.B(n_602),
.Y(n_864)
);

NOR2xp33_ASAP7_75t_L g865 ( 
.A(n_691),
.B(n_228),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_L g866 ( 
.A(n_700),
.B(n_602),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_705),
.B(n_714),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_705),
.B(n_341),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_716),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_L g870 ( 
.A(n_714),
.B(n_343),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_L g871 ( 
.A(n_715),
.B(n_344),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_753),
.Y(n_872)
);

OAI22xp5_ASAP7_75t_L g873 ( 
.A1(n_642),
.A2(n_230),
.B1(n_412),
.B2(n_410),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_753),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_715),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_718),
.Y(n_876)
);

AND2x4_ASAP7_75t_L g877 ( 
.A(n_656),
.B(n_318),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_SL g878 ( 
.A(n_693),
.B(n_228),
.Y(n_878)
);

AND2x4_ASAP7_75t_SL g879 ( 
.A(n_640),
.B(n_286),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_SL g880 ( 
.A(n_702),
.B(n_229),
.Y(n_880)
);

NOR2xp33_ASAP7_75t_L g881 ( 
.A(n_703),
.B(n_229),
.Y(n_881)
);

AOI21xp5_ASAP7_75t_L g882 ( 
.A1(n_761),
.A2(n_380),
.B(n_375),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_718),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_L g884 ( 
.A(n_729),
.B(n_355),
.Y(n_884)
);

NOR2xp33_ASAP7_75t_L g885 ( 
.A(n_704),
.B(n_230),
.Y(n_885)
);

NOR2x1p5_ASAP7_75t_L g886 ( 
.A(n_710),
.B(n_227),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_L g887 ( 
.A(n_729),
.B(n_356),
.Y(n_887)
);

INVx2_ASAP7_75t_L g888 ( 
.A(n_641),
.Y(n_888)
);

INVx2_ASAP7_75t_L g889 ( 
.A(n_641),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_730),
.Y(n_890)
);

BUFx6f_ASAP7_75t_SL g891 ( 
.A(n_640),
.Y(n_891)
);

AOI22xp33_ASAP7_75t_L g892 ( 
.A1(n_677),
.A2(n_395),
.B1(n_358),
.B2(n_325),
.Y(n_892)
);

INVx2_ASAP7_75t_L g893 ( 
.A(n_650),
.Y(n_893)
);

INVx2_ASAP7_75t_L g894 ( 
.A(n_650),
.Y(n_894)
);

AND2x2_ASAP7_75t_L g895 ( 
.A(n_651),
.B(n_286),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_L g896 ( 
.A(n_730),
.B(n_357),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_SL g897 ( 
.A(n_678),
.B(n_248),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_SL g898 ( 
.A(n_695),
.B(n_248),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_L g899 ( 
.A(n_732),
.B(n_362),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_L g900 ( 
.A(n_732),
.B(n_367),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_737),
.B(n_372),
.Y(n_901)
);

OAI22xp5_ASAP7_75t_L g902 ( 
.A1(n_728),
.A2(n_415),
.B1(n_412),
.B2(n_410),
.Y(n_902)
);

INVx2_ASAP7_75t_SL g903 ( 
.A(n_669),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_SL g904 ( 
.A(n_646),
.B(n_248),
.Y(n_904)
);

INVx4_ASAP7_75t_L g905 ( 
.A(n_659),
.Y(n_905)
);

INVx5_ASAP7_75t_L g906 ( 
.A(n_643),
.Y(n_906)
);

NOR2xp33_ASAP7_75t_L g907 ( 
.A(n_720),
.B(n_232),
.Y(n_907)
);

OR2x2_ASAP7_75t_L g908 ( 
.A(n_726),
.B(n_689),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_747),
.B(n_373),
.Y(n_909)
);

INVx2_ASAP7_75t_L g910 ( 
.A(n_664),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_752),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_669),
.Y(n_912)
);

BUFx3_ASAP7_75t_L g913 ( 
.A(n_669),
.Y(n_913)
);

INVx2_ASAP7_75t_L g914 ( 
.A(n_664),
.Y(n_914)
);

BUFx6f_ASAP7_75t_SL g915 ( 
.A(n_640),
.Y(n_915)
);

NOR2xp33_ASAP7_75t_L g916 ( 
.A(n_727),
.B(n_232),
.Y(n_916)
);

INVx2_ASAP7_75t_L g917 ( 
.A(n_709),
.Y(n_917)
);

INVx2_ASAP7_75t_L g918 ( 
.A(n_709),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_SL g919 ( 
.A(n_646),
.B(n_248),
.Y(n_919)
);

NAND3xp33_ASAP7_75t_L g920 ( 
.A(n_760),
.B(n_415),
.C(n_409),
.Y(n_920)
);

INVx2_ASAP7_75t_L g921 ( 
.A(n_722),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_L g922 ( 
.A(n_748),
.B(n_235),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_754),
.Y(n_923)
);

BUFx6f_ASAP7_75t_SL g924 ( 
.A(n_649),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_754),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_SL g926 ( 
.A(n_748),
.B(n_248),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_L g927 ( 
.A(n_679),
.B(n_235),
.Y(n_927)
);

INVxp67_ASAP7_75t_L g928 ( 
.A(n_654),
.Y(n_928)
);

BUFx3_ASAP7_75t_L g929 ( 
.A(n_744),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_692),
.B(n_755),
.Y(n_930)
);

AOI22xp33_ASAP7_75t_L g931 ( 
.A1(n_643),
.A2(n_408),
.B1(n_393),
.B2(n_389),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_SL g932 ( 
.A(n_765),
.B(n_378),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_L g933 ( 
.A(n_743),
.B(n_236),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_L g934 ( 
.A(n_717),
.B(n_236),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_L g935 ( 
.A(n_717),
.B(n_238),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_SL g936 ( 
.A(n_751),
.B(n_378),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_L g937 ( 
.A(n_719),
.B(n_697),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_L g938 ( 
.A(n_719),
.B(n_238),
.Y(n_938)
);

INVx2_ASAP7_75t_L g939 ( 
.A(n_818),
.Y(n_939)
);

AOI21xp5_ASAP7_75t_L g940 ( 
.A1(n_789),
.A2(n_684),
.B(n_666),
.Y(n_940)
);

A2O1A1Ixp33_ASAP7_75t_L g941 ( 
.A1(n_767),
.A2(n_802),
.B(n_865),
.C(n_845),
.Y(n_941)
);

AOI21xp5_ASAP7_75t_L g942 ( 
.A1(n_774),
.A2(n_684),
.B(n_666),
.Y(n_942)
);

OAI22xp5_ASAP7_75t_L g943 ( 
.A1(n_791),
.A2(n_751),
.B1(n_756),
.B2(n_735),
.Y(n_943)
);

AOI21xp5_ASAP7_75t_L g944 ( 
.A1(n_839),
.A2(n_684),
.B(n_666),
.Y(n_944)
);

OAI21xp5_ASAP7_75t_L g945 ( 
.A1(n_926),
.A2(n_643),
.B(n_751),
.Y(n_945)
);

A2O1A1Ixp33_ASAP7_75t_L g946 ( 
.A1(n_767),
.A2(n_742),
.B(n_764),
.C(n_763),
.Y(n_946)
);

AOI22xp5_ASAP7_75t_L g947 ( 
.A1(n_831),
.A2(n_791),
.B1(n_802),
.B2(n_907),
.Y(n_947)
);

AOI21xp5_ASAP7_75t_L g948 ( 
.A1(n_844),
.A2(n_757),
.B(n_659),
.Y(n_948)
);

AOI21xp5_ASAP7_75t_L g949 ( 
.A1(n_847),
.A2(n_814),
.B(n_812),
.Y(n_949)
);

INVxp67_ASAP7_75t_L g950 ( 
.A(n_797),
.Y(n_950)
);

INVx3_ASAP7_75t_L g951 ( 
.A(n_829),
.Y(n_951)
);

AOI21xp33_ASAP7_75t_L g952 ( 
.A1(n_907),
.A2(n_673),
.B(n_741),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_SL g953 ( 
.A(n_837),
.B(n_649),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_L g954 ( 
.A(n_845),
.B(n_643),
.Y(n_954)
);

AOI21xp33_ASAP7_75t_L g955 ( 
.A1(n_865),
.A2(n_633),
.B(n_637),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_SL g956 ( 
.A(n_853),
.B(n_829),
.Y(n_956)
);

AOI21xp5_ASAP7_75t_L g957 ( 
.A1(n_768),
.A2(n_757),
.B(n_659),
.Y(n_957)
);

AOI21xp5_ASAP7_75t_L g958 ( 
.A1(n_769),
.A2(n_819),
.B(n_815),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_L g959 ( 
.A(n_881),
.B(n_885),
.Y(n_959)
);

AOI21xp5_ASAP7_75t_L g960 ( 
.A1(n_937),
.A2(n_757),
.B(n_659),
.Y(n_960)
);

NOR2xp33_ASAP7_75t_L g961 ( 
.A(n_928),
.B(n_713),
.Y(n_961)
);

O2A1O1Ixp33_ASAP7_75t_L g962 ( 
.A1(n_788),
.A2(n_688),
.B(n_733),
.C(n_725),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_L g963 ( 
.A(n_881),
.B(n_756),
.Y(n_963)
);

AND2x4_ASAP7_75t_L g964 ( 
.A(n_853),
.B(n_712),
.Y(n_964)
);

AOI33xp33_ASAP7_75t_L g965 ( 
.A1(n_860),
.A2(n_696),
.A3(n_366),
.B1(n_740),
.B2(n_721),
.B3(n_734),
.Y(n_965)
);

INVx3_ASAP7_75t_L g966 ( 
.A(n_829),
.Y(n_966)
);

NAND2x1_ASAP7_75t_L g967 ( 
.A(n_905),
.B(n_784),
.Y(n_967)
);

O2A1O1Ixp33_ASAP7_75t_L g968 ( 
.A1(n_851),
.A2(n_724),
.B(n_722),
.C(n_738),
.Y(n_968)
);

AOI21xp5_ASAP7_75t_L g969 ( 
.A1(n_775),
.A2(n_731),
.B(n_659),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_L g970 ( 
.A(n_885),
.B(n_724),
.Y(n_970)
);

HB1xp67_ASAP7_75t_L g971 ( 
.A(n_817),
.Y(n_971)
);

NAND2x1_ASAP7_75t_L g972 ( 
.A(n_905),
.B(n_697),
.Y(n_972)
);

INVx1_ASAP7_75t_L g973 ( 
.A(n_773),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_782),
.Y(n_974)
);

AOI21xp5_ASAP7_75t_L g975 ( 
.A1(n_776),
.A2(n_781),
.B(n_780),
.Y(n_975)
);

INVx2_ASAP7_75t_L g976 ( 
.A(n_818),
.Y(n_976)
);

AOI21xp5_ASAP7_75t_L g977 ( 
.A1(n_786),
.A2(n_926),
.B(n_898),
.Y(n_977)
);

AOI21xp5_ASAP7_75t_L g978 ( 
.A1(n_898),
.A2(n_731),
.B(n_762),
.Y(n_978)
);

NAND2xp5_ASAP7_75t_L g979 ( 
.A(n_875),
.B(n_738),
.Y(n_979)
);

OAI21xp5_ASAP7_75t_L g980 ( 
.A1(n_922),
.A2(n_746),
.B(n_701),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_L g981 ( 
.A(n_876),
.B(n_749),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_L g982 ( 
.A(n_883),
.B(n_890),
.Y(n_982)
);

INVx4_ASAP7_75t_L g983 ( 
.A(n_829),
.Y(n_983)
);

NOR2xp33_ASAP7_75t_L g984 ( 
.A(n_836),
.B(n_713),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_783),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_L g986 ( 
.A(n_790),
.B(n_749),
.Y(n_986)
);

AND2x2_ASAP7_75t_L g987 ( 
.A(n_895),
.B(n_649),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_L g988 ( 
.A(n_804),
.B(n_697),
.Y(n_988)
);

NOR2x1_ASAP7_75t_L g989 ( 
.A(n_801),
.B(n_658),
.Y(n_989)
);

INVx1_ASAP7_75t_SL g990 ( 
.A(n_807),
.Y(n_990)
);

AOI21xp5_ASAP7_75t_L g991 ( 
.A1(n_930),
.A2(n_731),
.B(n_762),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_SL g992 ( 
.A(n_908),
.B(n_913),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_L g993 ( 
.A(n_805),
.B(n_701),
.Y(n_993)
);

AND2x2_ASAP7_75t_L g994 ( 
.A(n_798),
.B(n_685),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_L g995 ( 
.A(n_810),
.B(n_701),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_SL g996 ( 
.A(n_913),
.B(n_685),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_821),
.Y(n_997)
);

INVx1_ASAP7_75t_L g998 ( 
.A(n_923),
.Y(n_998)
);

NOR2xp33_ASAP7_75t_L g999 ( 
.A(n_800),
.B(n_672),
.Y(n_999)
);

AOI21xp5_ASAP7_75t_L g1000 ( 
.A1(n_809),
.A2(n_731),
.B(n_759),
.Y(n_1000)
);

BUFx6f_ASAP7_75t_L g1001 ( 
.A(n_784),
.Y(n_1001)
);

AOI21xp5_ASAP7_75t_L g1002 ( 
.A1(n_816),
.A2(n_731),
.B(n_759),
.Y(n_1002)
);

AOI21xp5_ASAP7_75t_L g1003 ( 
.A1(n_771),
.A2(n_766),
.B(n_759),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_L g1004 ( 
.A(n_811),
.B(n_706),
.Y(n_1004)
);

OAI21xp5_ASAP7_75t_L g1005 ( 
.A1(n_854),
.A2(n_766),
.B(n_746),
.Y(n_1005)
);

INVxp67_ASAP7_75t_SL g1006 ( 
.A(n_811),
.Y(n_1006)
);

NOR3xp33_ASAP7_75t_L g1007 ( 
.A(n_823),
.B(n_687),
.C(n_723),
.Y(n_1007)
);

INVx1_ASAP7_75t_L g1008 ( 
.A(n_925),
.Y(n_1008)
);

OAI22xp5_ASAP7_75t_L g1009 ( 
.A1(n_833),
.A2(n_660),
.B1(n_675),
.B2(n_376),
.Y(n_1009)
);

AOI21xp5_ASAP7_75t_L g1010 ( 
.A1(n_771),
.A2(n_766),
.B(n_746),
.Y(n_1010)
);

O2A1O1Ixp33_ASAP7_75t_L g1011 ( 
.A1(n_869),
.A2(n_624),
.B(n_706),
.C(n_314),
.Y(n_1011)
);

NAND2x1p5_ASAP7_75t_L g1012 ( 
.A(n_771),
.B(n_663),
.Y(n_1012)
);

AOI21xp5_ASAP7_75t_L g1013 ( 
.A1(n_771),
.A2(n_706),
.B(n_663),
.Y(n_1013)
);

AOI21xp5_ASAP7_75t_L g1014 ( 
.A1(n_906),
.A2(n_830),
.B(n_828),
.Y(n_1014)
);

AOI21xp5_ASAP7_75t_L g1015 ( 
.A1(n_906),
.A2(n_663),
.B(n_683),
.Y(n_1015)
);

INVx1_ASAP7_75t_L g1016 ( 
.A(n_770),
.Y(n_1016)
);

INVxp67_ASAP7_75t_L g1017 ( 
.A(n_798),
.Y(n_1017)
);

NAND2xp33_ASAP7_75t_L g1018 ( 
.A(n_862),
.B(n_378),
.Y(n_1018)
);

OAI22xp5_ASAP7_75t_L g1019 ( 
.A1(n_833),
.A2(n_892),
.B1(n_859),
.B2(n_912),
.Y(n_1019)
);

AOI21xp5_ASAP7_75t_L g1020 ( 
.A1(n_906),
.A2(n_663),
.B(n_683),
.Y(n_1020)
);

HB1xp67_ASAP7_75t_L g1021 ( 
.A(n_872),
.Y(n_1021)
);

AO21x1_ASAP7_75t_L g1022 ( 
.A1(n_936),
.A2(n_378),
.B(n_17),
.Y(n_1022)
);

INVx2_ASAP7_75t_SL g1023 ( 
.A(n_877),
.Y(n_1023)
);

AOI21xp5_ASAP7_75t_L g1024 ( 
.A1(n_906),
.A2(n_663),
.B(n_683),
.Y(n_1024)
);

AOI21xp5_ASAP7_75t_L g1025 ( 
.A1(n_827),
.A2(n_683),
.B(n_397),
.Y(n_1025)
);

O2A1O1Ixp33_ASAP7_75t_SL g1026 ( 
.A1(n_897),
.A2(n_378),
.B(n_244),
.C(n_245),
.Y(n_1026)
);

AOI21xp5_ASAP7_75t_L g1027 ( 
.A1(n_867),
.A2(n_683),
.B(n_397),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_L g1028 ( 
.A(n_826),
.B(n_241),
.Y(n_1028)
);

AOI21xp5_ASAP7_75t_L g1029 ( 
.A1(n_897),
.A2(n_257),
.B(n_409),
.Y(n_1029)
);

INVx1_ASAP7_75t_L g1030 ( 
.A(n_770),
.Y(n_1030)
);

AOI21xp5_ASAP7_75t_L g1031 ( 
.A1(n_796),
.A2(n_868),
.B(n_806),
.Y(n_1031)
);

AOI21xp5_ASAP7_75t_L g1032 ( 
.A1(n_794),
.A2(n_390),
.B(n_241),
.Y(n_1032)
);

INVx2_ASAP7_75t_SL g1033 ( 
.A(n_877),
.Y(n_1033)
);

OAI22xp5_ASAP7_75t_L g1034 ( 
.A1(n_892),
.A2(n_258),
.B1(n_244),
.B2(n_245),
.Y(n_1034)
);

INVx1_ASAP7_75t_L g1035 ( 
.A(n_779),
.Y(n_1035)
);

INVx1_ASAP7_75t_L g1036 ( 
.A(n_779),
.Y(n_1036)
);

O2A1O1Ixp33_ASAP7_75t_SL g1037 ( 
.A1(n_936),
.A2(n_378),
.B(n_257),
.C(n_258),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_L g1038 ( 
.A(n_834),
.B(n_254),
.Y(n_1038)
);

AND2x2_ASAP7_75t_L g1039 ( 
.A(n_808),
.B(n_739),
.Y(n_1039)
);

OAI22xp5_ASAP7_75t_L g1040 ( 
.A1(n_874),
.A2(n_254),
.B1(n_259),
.B2(n_402),
.Y(n_1040)
);

OAI21xp5_ASAP7_75t_L g1041 ( 
.A1(n_772),
.A2(n_384),
.B(n_259),
.Y(n_1041)
);

OAI22xp5_ASAP7_75t_L g1042 ( 
.A1(n_903),
.A2(n_384),
.B1(n_316),
.B2(n_402),
.Y(n_1042)
);

NAND2xp5_ASAP7_75t_SL g1043 ( 
.A(n_933),
.B(n_316),
.Y(n_1043)
);

BUFx4f_ASAP7_75t_L g1044 ( 
.A(n_778),
.Y(n_1044)
);

INVxp67_ASAP7_75t_L g1045 ( 
.A(n_808),
.Y(n_1045)
);

AOI21xp5_ASAP7_75t_L g1046 ( 
.A1(n_856),
.A2(n_387),
.B(n_388),
.Y(n_1046)
);

A2O1A1Ixp33_ASAP7_75t_L g1047 ( 
.A1(n_916),
.A2(n_387),
.B(n_388),
.C(n_390),
.Y(n_1047)
);

NAND2xp33_ASAP7_75t_L g1048 ( 
.A(n_862),
.B(n_378),
.Y(n_1048)
);

OAI21xp5_ASAP7_75t_L g1049 ( 
.A1(n_864),
.A2(n_406),
.B(n_404),
.Y(n_1049)
);

INVx1_ASAP7_75t_L g1050 ( 
.A(n_787),
.Y(n_1050)
);

BUFx3_ASAP7_75t_L g1051 ( 
.A(n_850),
.Y(n_1051)
);

AND2x2_ASAP7_75t_L g1052 ( 
.A(n_838),
.B(n_233),
.Y(n_1052)
);

O2A1O1Ixp33_ASAP7_75t_L g1053 ( 
.A1(n_813),
.A2(n_406),
.B(n_404),
.C(n_400),
.Y(n_1053)
);

AND2x2_ASAP7_75t_L g1054 ( 
.A(n_838),
.B(n_233),
.Y(n_1054)
);

INVxp67_ASAP7_75t_L g1055 ( 
.A(n_916),
.Y(n_1055)
);

AND2x2_ASAP7_75t_L g1056 ( 
.A(n_861),
.B(n_879),
.Y(n_1056)
);

HB1xp67_ASAP7_75t_L g1057 ( 
.A(n_863),
.Y(n_1057)
);

AOI21xp5_ASAP7_75t_L g1058 ( 
.A1(n_866),
.A2(n_400),
.B(n_399),
.Y(n_1058)
);

AOI21xp5_ASAP7_75t_L g1059 ( 
.A1(n_934),
.A2(n_399),
.B(n_396),
.Y(n_1059)
);

AOI22xp5_ASAP7_75t_L g1060 ( 
.A1(n_778),
.A2(n_378),
.B1(n_396),
.B2(n_383),
.Y(n_1060)
);

O2A1O1Ixp5_ASAP7_75t_L g1061 ( 
.A1(n_832),
.A2(n_385),
.B(n_383),
.C(n_381),
.Y(n_1061)
);

NOR2x1_ASAP7_75t_L g1062 ( 
.A(n_785),
.B(n_385),
.Y(n_1062)
);

NAND2xp5_ASAP7_75t_SL g1063 ( 
.A(n_927),
.B(n_381),
.Y(n_1063)
);

NAND2xp5_ASAP7_75t_SL g1064 ( 
.A(n_870),
.B(n_255),
.Y(n_1064)
);

INVx2_ASAP7_75t_L g1065 ( 
.A(n_820),
.Y(n_1065)
);

OAI22xp5_ASAP7_75t_L g1066 ( 
.A1(n_842),
.A2(n_911),
.B1(n_931),
.B2(n_793),
.Y(n_1066)
);

AOI21xp5_ASAP7_75t_L g1067 ( 
.A1(n_935),
.A2(n_255),
.B(n_253),
.Y(n_1067)
);

NAND2xp5_ASAP7_75t_L g1068 ( 
.A(n_848),
.B(n_253),
.Y(n_1068)
);

AND2x6_ASAP7_75t_L g1069 ( 
.A(n_787),
.B(n_204),
.Y(n_1069)
);

AOI21xp5_ASAP7_75t_L g1070 ( 
.A1(n_938),
.A2(n_243),
.B(n_239),
.Y(n_1070)
);

NAND2xp5_ASAP7_75t_L g1071 ( 
.A(n_852),
.B(n_243),
.Y(n_1071)
);

NOR2xp33_ASAP7_75t_L g1072 ( 
.A(n_873),
.B(n_239),
.Y(n_1072)
);

BUFx6f_ASAP7_75t_L g1073 ( 
.A(n_803),
.Y(n_1073)
);

OAI21xp5_ASAP7_75t_L g1074 ( 
.A1(n_820),
.A2(n_199),
.B(n_197),
.Y(n_1074)
);

AOI21xp5_ASAP7_75t_L g1075 ( 
.A1(n_871),
.A2(n_185),
.B(n_184),
.Y(n_1075)
);

NOR2xp33_ASAP7_75t_L g1076 ( 
.A(n_849),
.B(n_16),
.Y(n_1076)
);

HB1xp67_ASAP7_75t_L g1077 ( 
.A(n_855),
.Y(n_1077)
);

O2A1O1Ixp33_ASAP7_75t_SL g1078 ( 
.A1(n_799),
.A2(n_16),
.B(n_17),
.C(n_19),
.Y(n_1078)
);

BUFx12f_ASAP7_75t_L g1079 ( 
.A(n_843),
.Y(n_1079)
);

AOI22xp33_ASAP7_75t_SL g1080 ( 
.A1(n_879),
.A2(n_19),
.B1(n_21),
.B2(n_23),
.Y(n_1080)
);

OAI21xp5_ASAP7_75t_L g1081 ( 
.A1(n_835),
.A2(n_179),
.B(n_172),
.Y(n_1081)
);

NAND2xp5_ASAP7_75t_SL g1082 ( 
.A(n_884),
.B(n_162),
.Y(n_1082)
);

OAI22xp5_ASAP7_75t_L g1083 ( 
.A1(n_931),
.A2(n_160),
.B1(n_152),
.B2(n_145),
.Y(n_1083)
);

NAND2xp5_ASAP7_75t_L g1084 ( 
.A(n_887),
.B(n_25),
.Y(n_1084)
);

OAI21xp33_ASAP7_75t_L g1085 ( 
.A1(n_878),
.A2(n_26),
.B(n_29),
.Y(n_1085)
);

NOR2x1_ASAP7_75t_L g1086 ( 
.A(n_841),
.B(n_141),
.Y(n_1086)
);

AOI22xp33_ASAP7_75t_L g1087 ( 
.A1(n_778),
.A2(n_30),
.B1(n_31),
.B2(n_36),
.Y(n_1087)
);

INVx2_ASAP7_75t_L g1088 ( 
.A(n_835),
.Y(n_1088)
);

AOI21xp5_ASAP7_75t_L g1089 ( 
.A1(n_896),
.A2(n_136),
.B(n_118),
.Y(n_1089)
);

OAI22xp5_ASAP7_75t_L g1090 ( 
.A1(n_899),
.A2(n_113),
.B1(n_111),
.B2(n_109),
.Y(n_1090)
);

AOI21xp5_ASAP7_75t_L g1091 ( 
.A1(n_900),
.A2(n_103),
.B(n_94),
.Y(n_1091)
);

INVx2_ASAP7_75t_L g1092 ( 
.A(n_857),
.Y(n_1092)
);

NAND2xp5_ASAP7_75t_L g1093 ( 
.A(n_921),
.B(n_889),
.Y(n_1093)
);

AOI21xp5_ASAP7_75t_L g1094 ( 
.A1(n_901),
.A2(n_85),
.B(n_81),
.Y(n_1094)
);

AOI21xp5_ASAP7_75t_L g1095 ( 
.A1(n_909),
.A2(n_79),
.B(n_38),
.Y(n_1095)
);

OAI22xp5_ASAP7_75t_L g1096 ( 
.A1(n_822),
.A2(n_72),
.B1(n_41),
.B2(n_42),
.Y(n_1096)
);

AOI21xp5_ASAP7_75t_L g1097 ( 
.A1(n_932),
.A2(n_31),
.B(n_41),
.Y(n_1097)
);

NAND2xp5_ASAP7_75t_L g1098 ( 
.A(n_921),
.B(n_889),
.Y(n_1098)
);

BUFx2_ASAP7_75t_L g1099 ( 
.A(n_777),
.Y(n_1099)
);

INVx4_ASAP7_75t_L g1100 ( 
.A(n_891),
.Y(n_1100)
);

NAND2xp5_ASAP7_75t_L g1101 ( 
.A(n_857),
.B(n_893),
.Y(n_1101)
);

INVxp67_ASAP7_75t_L g1102 ( 
.A(n_824),
.Y(n_1102)
);

NAND2xp5_ASAP7_75t_L g1103 ( 
.A(n_888),
.B(n_43),
.Y(n_1103)
);

O2A1O1Ixp33_ASAP7_75t_L g1104 ( 
.A1(n_792),
.A2(n_44),
.B(n_45),
.C(n_48),
.Y(n_1104)
);

AND2x2_ASAP7_75t_L g1105 ( 
.A(n_886),
.B(n_72),
.Y(n_1105)
);

AND2x2_ASAP7_75t_L g1106 ( 
.A(n_880),
.B(n_48),
.Y(n_1106)
);

AOI21xp5_ASAP7_75t_L g1107 ( 
.A1(n_932),
.A2(n_49),
.B(n_50),
.Y(n_1107)
);

AOI21xp5_ASAP7_75t_L g1108 ( 
.A1(n_904),
.A2(n_919),
.B(n_858),
.Y(n_1108)
);

AOI21xp5_ASAP7_75t_L g1109 ( 
.A1(n_904),
.A2(n_50),
.B(n_55),
.Y(n_1109)
);

A2O1A1Ixp33_ASAP7_75t_L g1110 ( 
.A1(n_920),
.A2(n_56),
.B(n_57),
.C(n_61),
.Y(n_1110)
);

AOI21xp5_ASAP7_75t_L g1111 ( 
.A1(n_919),
.A2(n_63),
.B(n_64),
.Y(n_1111)
);

NAND2xp5_ASAP7_75t_L g1112 ( 
.A(n_894),
.B(n_67),
.Y(n_1112)
);

INVx2_ASAP7_75t_SL g1113 ( 
.A(n_929),
.Y(n_1113)
);

AOI21xp5_ASAP7_75t_L g1114 ( 
.A1(n_832),
.A2(n_67),
.B(n_68),
.Y(n_1114)
);

HB1xp67_ASAP7_75t_L g1115 ( 
.A(n_894),
.Y(n_1115)
);

OAI22xp5_ASAP7_75t_L g1116 ( 
.A1(n_840),
.A2(n_69),
.B1(n_70),
.B2(n_71),
.Y(n_1116)
);

OR2x2_ASAP7_75t_L g1117 ( 
.A(n_825),
.B(n_69),
.Y(n_1117)
);

NOR2xp33_ASAP7_75t_SL g1118 ( 
.A(n_891),
.B(n_70),
.Y(n_1118)
);

NAND2xp5_ASAP7_75t_L g1119 ( 
.A(n_910),
.B(n_918),
.Y(n_1119)
);

AOI21xp5_ASAP7_75t_L g1120 ( 
.A1(n_858),
.A2(n_910),
.B(n_917),
.Y(n_1120)
);

OA22x2_ASAP7_75t_L g1121 ( 
.A1(n_902),
.A2(n_914),
.B1(n_918),
.B2(n_917),
.Y(n_1121)
);

NOR2xp33_ASAP7_75t_R g1122 ( 
.A(n_929),
.B(n_924),
.Y(n_1122)
);

NAND2xp5_ASAP7_75t_L g1123 ( 
.A(n_914),
.B(n_778),
.Y(n_1123)
);

INVx2_ASAP7_75t_L g1124 ( 
.A(n_778),
.Y(n_1124)
);

AOI21xp5_ASAP7_75t_L g1125 ( 
.A1(n_882),
.A2(n_862),
.B(n_795),
.Y(n_1125)
);

NOR2xp33_ASAP7_75t_L g1126 ( 
.A(n_915),
.B(n_924),
.Y(n_1126)
);

AND2x2_ASAP7_75t_L g1127 ( 
.A(n_846),
.B(n_915),
.Y(n_1127)
);

NAND2xp5_ASAP7_75t_SL g1128 ( 
.A(n_862),
.B(n_837),
.Y(n_1128)
);

AOI21xp5_ASAP7_75t_L g1129 ( 
.A1(n_862),
.A2(n_625),
.B(n_616),
.Y(n_1129)
);

AOI21xp5_ASAP7_75t_L g1130 ( 
.A1(n_1129),
.A2(n_862),
.B(n_975),
.Y(n_1130)
);

AND2x2_ASAP7_75t_L g1131 ( 
.A(n_994),
.B(n_1052),
.Y(n_1131)
);

NAND2xp5_ASAP7_75t_SL g1132 ( 
.A(n_941),
.B(n_959),
.Y(n_1132)
);

AOI21x1_ASAP7_75t_L g1133 ( 
.A1(n_949),
.A2(n_958),
.B(n_1128),
.Y(n_1133)
);

AOI21x1_ASAP7_75t_L g1134 ( 
.A1(n_1123),
.A2(n_940),
.B(n_970),
.Y(n_1134)
);

AOI21xp5_ASAP7_75t_L g1135 ( 
.A1(n_945),
.A2(n_977),
.B(n_954),
.Y(n_1135)
);

NAND2xp5_ASAP7_75t_L g1136 ( 
.A(n_1077),
.B(n_1017),
.Y(n_1136)
);

AO21x2_ASAP7_75t_L g1137 ( 
.A1(n_980),
.A2(n_1005),
.B(n_947),
.Y(n_1137)
);

BUFx6f_ASAP7_75t_L g1138 ( 
.A(n_1001),
.Y(n_1138)
);

NAND2xp5_ASAP7_75t_SL g1139 ( 
.A(n_1055),
.B(n_943),
.Y(n_1139)
);

AOI21xp33_ASAP7_75t_L g1140 ( 
.A1(n_1072),
.A2(n_962),
.B(n_1055),
.Y(n_1140)
);

NAND2xp5_ASAP7_75t_L g1141 ( 
.A(n_1077),
.B(n_1017),
.Y(n_1141)
);

INVx1_ASAP7_75t_L g1142 ( 
.A(n_1115),
.Y(n_1142)
);

INVx1_ASAP7_75t_L g1143 ( 
.A(n_1115),
.Y(n_1143)
);

NAND2xp5_ASAP7_75t_L g1144 ( 
.A(n_1045),
.B(n_1054),
.Y(n_1144)
);

BUFx3_ASAP7_75t_L g1145 ( 
.A(n_1099),
.Y(n_1145)
);

NAND2xp5_ASAP7_75t_L g1146 ( 
.A(n_1045),
.B(n_973),
.Y(n_1146)
);

AO31x2_ASAP7_75t_L g1147 ( 
.A1(n_1022),
.A2(n_1019),
.A3(n_1066),
.B(n_1076),
.Y(n_1147)
);

AND2x2_ASAP7_75t_L g1148 ( 
.A(n_987),
.B(n_1039),
.Y(n_1148)
);

BUFx6f_ASAP7_75t_L g1149 ( 
.A(n_1001),
.Y(n_1149)
);

INVx1_ASAP7_75t_L g1150 ( 
.A(n_1021),
.Y(n_1150)
);

AOI21x1_ASAP7_75t_L g1151 ( 
.A1(n_960),
.A2(n_948),
.B(n_944),
.Y(n_1151)
);

AND2x4_ASAP7_75t_L g1152 ( 
.A(n_964),
.B(n_983),
.Y(n_1152)
);

CKINVDCx5p33_ASAP7_75t_R g1153 ( 
.A(n_1079),
.Y(n_1153)
);

OR2x2_ASAP7_75t_L g1154 ( 
.A(n_990),
.B(n_971),
.Y(n_1154)
);

OAI21xp5_ASAP7_75t_L g1155 ( 
.A1(n_1108),
.A2(n_1121),
.B(n_1120),
.Y(n_1155)
);

AOI221xp5_ASAP7_75t_L g1156 ( 
.A1(n_1072),
.A2(n_1009),
.B1(n_1076),
.B2(n_952),
.C(n_1034),
.Y(n_1156)
);

INVxp67_ASAP7_75t_L g1157 ( 
.A(n_971),
.Y(n_1157)
);

OR2x2_ASAP7_75t_L g1158 ( 
.A(n_1068),
.B(n_1071),
.Y(n_1158)
);

AND2x2_ASAP7_75t_L g1159 ( 
.A(n_961),
.B(n_984),
.Y(n_1159)
);

OAI21x1_ASAP7_75t_L g1160 ( 
.A1(n_1121),
.A2(n_957),
.B(n_942),
.Y(n_1160)
);

NAND2xp5_ASAP7_75t_L g1161 ( 
.A(n_974),
.B(n_985),
.Y(n_1161)
);

NAND2xp5_ASAP7_75t_L g1162 ( 
.A(n_997),
.B(n_982),
.Y(n_1162)
);

AOI21xp5_ASAP7_75t_L g1163 ( 
.A1(n_1031),
.A2(n_1014),
.B(n_1125),
.Y(n_1163)
);

AOI21xp5_ASAP7_75t_L g1164 ( 
.A1(n_1018),
.A2(n_1048),
.B(n_1006),
.Y(n_1164)
);

INVx2_ASAP7_75t_L g1165 ( 
.A(n_939),
.Y(n_1165)
);

BUFx4f_ASAP7_75t_SL g1166 ( 
.A(n_1051),
.Y(n_1166)
);

NAND2xp5_ASAP7_75t_L g1167 ( 
.A(n_963),
.B(n_1021),
.Y(n_1167)
);

OAI21xp5_ASAP7_75t_L g1168 ( 
.A1(n_978),
.A2(n_991),
.B(n_1093),
.Y(n_1168)
);

NAND2xp5_ASAP7_75t_L g1169 ( 
.A(n_1006),
.B(n_998),
.Y(n_1169)
);

AOI21xp5_ASAP7_75t_L g1170 ( 
.A1(n_1004),
.A2(n_969),
.B(n_967),
.Y(n_1170)
);

INVx1_ASAP7_75t_L g1171 ( 
.A(n_1016),
.Y(n_1171)
);

OAI21x1_ASAP7_75t_L g1172 ( 
.A1(n_1000),
.A2(n_1002),
.B(n_968),
.Y(n_1172)
);

INVx3_ASAP7_75t_L g1173 ( 
.A(n_1001),
.Y(n_1173)
);

NOR2xp67_ASAP7_75t_L g1174 ( 
.A(n_1100),
.B(n_1102),
.Y(n_1174)
);

OAI21x1_ASAP7_75t_L g1175 ( 
.A1(n_1124),
.A2(n_1010),
.B(n_1003),
.Y(n_1175)
);

NAND2xp5_ASAP7_75t_L g1176 ( 
.A(n_1008),
.B(n_946),
.Y(n_1176)
);

OAI21x1_ASAP7_75t_L g1177 ( 
.A1(n_1013),
.A2(n_1101),
.B(n_1098),
.Y(n_1177)
);

BUFx2_ASAP7_75t_L g1178 ( 
.A(n_950),
.Y(n_1178)
);

INVx4_ASAP7_75t_L g1179 ( 
.A(n_983),
.Y(n_1179)
);

AOI21xp5_ASAP7_75t_L g1180 ( 
.A1(n_1119),
.A2(n_956),
.B(n_992),
.Y(n_1180)
);

OAI21xp5_ASAP7_75t_L g1181 ( 
.A1(n_1084),
.A2(n_1061),
.B(n_988),
.Y(n_1181)
);

AOI21xp5_ASAP7_75t_SL g1182 ( 
.A1(n_1074),
.A2(n_1081),
.B(n_1001),
.Y(n_1182)
);

BUFx6f_ASAP7_75t_L g1183 ( 
.A(n_1073),
.Y(n_1183)
);

NAND2xp5_ASAP7_75t_L g1184 ( 
.A(n_1049),
.B(n_1102),
.Y(n_1184)
);

BUFx3_ASAP7_75t_L g1185 ( 
.A(n_964),
.Y(n_1185)
);

OAI21xp5_ASAP7_75t_L g1186 ( 
.A1(n_1061),
.A2(n_993),
.B(n_995),
.Y(n_1186)
);

OAI22xp5_ASAP7_75t_L g1187 ( 
.A1(n_1044),
.A2(n_961),
.B1(n_1087),
.B2(n_953),
.Y(n_1187)
);

OAI21x1_ASAP7_75t_L g1188 ( 
.A1(n_972),
.A2(n_1103),
.B(n_1112),
.Y(n_1188)
);

AND2x2_ASAP7_75t_L g1189 ( 
.A(n_984),
.B(n_1056),
.Y(n_1189)
);

INVx1_ASAP7_75t_L g1190 ( 
.A(n_1030),
.Y(n_1190)
);

NAND2xp5_ASAP7_75t_L g1191 ( 
.A(n_955),
.B(n_1106),
.Y(n_1191)
);

AO31x2_ASAP7_75t_L g1192 ( 
.A1(n_1110),
.A2(n_1047),
.A3(n_1096),
.B(n_1116),
.Y(n_1192)
);

INVx2_ASAP7_75t_L g1193 ( 
.A(n_976),
.Y(n_1193)
);

AOI21xp5_ASAP7_75t_L g1194 ( 
.A1(n_986),
.A2(n_981),
.B(n_979),
.Y(n_1194)
);

OAI21xp5_ASAP7_75t_L g1195 ( 
.A1(n_1035),
.A2(n_1036),
.B(n_1050),
.Y(n_1195)
);

AOI21xp5_ASAP7_75t_L g1196 ( 
.A1(n_1082),
.A2(n_1012),
.B(n_1044),
.Y(n_1196)
);

CKINVDCx20_ASAP7_75t_R g1197 ( 
.A(n_1122),
.Y(n_1197)
);

NAND2xp5_ASAP7_75t_L g1198 ( 
.A(n_951),
.B(n_966),
.Y(n_1198)
);

BUFx10_ASAP7_75t_L g1199 ( 
.A(n_1126),
.Y(n_1199)
);

NAND2xp5_ASAP7_75t_L g1200 ( 
.A(n_999),
.B(n_1065),
.Y(n_1200)
);

AOI21xp5_ASAP7_75t_L g1201 ( 
.A1(n_1012),
.A2(n_1073),
.B(n_1088),
.Y(n_1201)
);

AOI21xp5_ASAP7_75t_L g1202 ( 
.A1(n_1073),
.A2(n_1092),
.B(n_1025),
.Y(n_1202)
);

OAI21x1_ASAP7_75t_L g1203 ( 
.A1(n_1015),
.A2(n_1024),
.B(n_1020),
.Y(n_1203)
);

OA21x2_ASAP7_75t_L g1204 ( 
.A1(n_1041),
.A2(n_1095),
.B(n_1089),
.Y(n_1204)
);

AND2x2_ASAP7_75t_L g1205 ( 
.A(n_950),
.B(n_999),
.Y(n_1205)
);

AOI21xp5_ASAP7_75t_L g1206 ( 
.A1(n_1073),
.A2(n_1033),
.B(n_1023),
.Y(n_1206)
);

A2O1A1Ixp33_ASAP7_75t_L g1207 ( 
.A1(n_1085),
.A2(n_1087),
.B(n_1011),
.C(n_1104),
.Y(n_1207)
);

NAND2xp5_ASAP7_75t_L g1208 ( 
.A(n_1028),
.B(n_1038),
.Y(n_1208)
);

CKINVDCx8_ASAP7_75t_R g1209 ( 
.A(n_1126),
.Y(n_1209)
);

OAI21x1_ASAP7_75t_L g1210 ( 
.A1(n_1075),
.A2(n_1091),
.B(n_1094),
.Y(n_1210)
);

AOI21xp5_ASAP7_75t_L g1211 ( 
.A1(n_1027),
.A2(n_1043),
.B(n_1083),
.Y(n_1211)
);

INVx2_ASAP7_75t_L g1212 ( 
.A(n_1069),
.Y(n_1212)
);

AND2x2_ASAP7_75t_L g1213 ( 
.A(n_1057),
.B(n_1105),
.Y(n_1213)
);

OAI21xp5_ASAP7_75t_L g1214 ( 
.A1(n_1063),
.A2(n_1064),
.B(n_1029),
.Y(n_1214)
);

OAI21x1_ASAP7_75t_L g1215 ( 
.A1(n_1090),
.A2(n_1111),
.B(n_1109),
.Y(n_1215)
);

INVx1_ASAP7_75t_SL g1216 ( 
.A(n_1117),
.Y(n_1216)
);

AOI21xp5_ASAP7_75t_L g1217 ( 
.A1(n_996),
.A2(n_1037),
.B(n_1026),
.Y(n_1217)
);

OAI21x1_ASAP7_75t_L g1218 ( 
.A1(n_1114),
.A2(n_1097),
.B(n_1107),
.Y(n_1218)
);

AO21x2_ASAP7_75t_L g1219 ( 
.A1(n_1007),
.A2(n_1046),
.B(n_1032),
.Y(n_1219)
);

OAI21x1_ASAP7_75t_L g1220 ( 
.A1(n_1086),
.A2(n_989),
.B(n_1053),
.Y(n_1220)
);

AND2x2_ASAP7_75t_SL g1221 ( 
.A(n_1007),
.B(n_1060),
.Y(n_1221)
);

NAND2xp5_ASAP7_75t_L g1222 ( 
.A(n_1058),
.B(n_1070),
.Y(n_1222)
);

AOI22xp33_ASAP7_75t_L g1223 ( 
.A1(n_1080),
.A2(n_1069),
.B1(n_1062),
.B2(n_1118),
.Y(n_1223)
);

OAI21x1_ASAP7_75t_L g1224 ( 
.A1(n_1059),
.A2(n_1067),
.B(n_1042),
.Y(n_1224)
);

BUFx6f_ASAP7_75t_L g1225 ( 
.A(n_1069),
.Y(n_1225)
);

NOR3xp33_ASAP7_75t_L g1226 ( 
.A(n_965),
.B(n_1040),
.C(n_1080),
.Y(n_1226)
);

INVx1_ASAP7_75t_SL g1227 ( 
.A(n_1057),
.Y(n_1227)
);

OAI21x1_ASAP7_75t_L g1228 ( 
.A1(n_1069),
.A2(n_1127),
.B(n_1078),
.Y(n_1228)
);

OAI21x1_ASAP7_75t_L g1229 ( 
.A1(n_1069),
.A2(n_1100),
.B(n_1113),
.Y(n_1229)
);

AO31x2_ASAP7_75t_L g1230 ( 
.A1(n_1122),
.A2(n_941),
.A3(n_1022),
.B(n_943),
.Y(n_1230)
);

OAI21x1_ASAP7_75t_L g1231 ( 
.A1(n_958),
.A2(n_1121),
.B(n_949),
.Y(n_1231)
);

INVx1_ASAP7_75t_L g1232 ( 
.A(n_1115),
.Y(n_1232)
);

AOI21xp5_ASAP7_75t_L g1233 ( 
.A1(n_1129),
.A2(n_625),
.B(n_616),
.Y(n_1233)
);

NOR2xp33_ASAP7_75t_L g1234 ( 
.A(n_1017),
.B(n_1045),
.Y(n_1234)
);

AND2x2_ASAP7_75t_L g1235 ( 
.A(n_994),
.B(n_1052),
.Y(n_1235)
);

AND2x2_ASAP7_75t_L g1236 ( 
.A(n_994),
.B(n_1052),
.Y(n_1236)
);

OAI21x1_ASAP7_75t_L g1237 ( 
.A1(n_958),
.A2(n_1121),
.B(n_949),
.Y(n_1237)
);

OAI21x1_ASAP7_75t_L g1238 ( 
.A1(n_958),
.A2(n_1121),
.B(n_949),
.Y(n_1238)
);

OA22x2_ASAP7_75t_L g1239 ( 
.A1(n_947),
.A2(n_836),
.B1(n_959),
.B2(n_800),
.Y(n_1239)
);

OAI21x1_ASAP7_75t_L g1240 ( 
.A1(n_958),
.A2(n_1121),
.B(n_949),
.Y(n_1240)
);

AOI21xp33_ASAP7_75t_L g1241 ( 
.A1(n_959),
.A2(n_767),
.B(n_941),
.Y(n_1241)
);

INVxp67_ASAP7_75t_L g1242 ( 
.A(n_971),
.Y(n_1242)
);

AOI21xp5_ASAP7_75t_L g1243 ( 
.A1(n_1129),
.A2(n_625),
.B(n_616),
.Y(n_1243)
);

AO21x1_ASAP7_75t_L g1244 ( 
.A1(n_959),
.A2(n_947),
.B(n_943),
.Y(n_1244)
);

OAI21x1_ASAP7_75t_L g1245 ( 
.A1(n_958),
.A2(n_1121),
.B(n_949),
.Y(n_1245)
);

OAI21x1_ASAP7_75t_L g1246 ( 
.A1(n_958),
.A2(n_1121),
.B(n_949),
.Y(n_1246)
);

AOI21x1_ASAP7_75t_L g1247 ( 
.A1(n_949),
.A2(n_926),
.B(n_898),
.Y(n_1247)
);

HB1xp67_ASAP7_75t_L g1248 ( 
.A(n_971),
.Y(n_1248)
);

AOI21xp5_ASAP7_75t_L g1249 ( 
.A1(n_1129),
.A2(n_625),
.B(n_616),
.Y(n_1249)
);

AOI21x1_ASAP7_75t_L g1250 ( 
.A1(n_949),
.A2(n_926),
.B(n_898),
.Y(n_1250)
);

OAI21x1_ASAP7_75t_L g1251 ( 
.A1(n_958),
.A2(n_1121),
.B(n_949),
.Y(n_1251)
);

OAI21xp5_ASAP7_75t_L g1252 ( 
.A1(n_941),
.A2(n_959),
.B(n_791),
.Y(n_1252)
);

BUFx6f_ASAP7_75t_L g1253 ( 
.A(n_1001),
.Y(n_1253)
);

OAI21x1_ASAP7_75t_L g1254 ( 
.A1(n_958),
.A2(n_1121),
.B(n_949),
.Y(n_1254)
);

OAI21x1_ASAP7_75t_L g1255 ( 
.A1(n_958),
.A2(n_1121),
.B(n_949),
.Y(n_1255)
);

AO31x2_ASAP7_75t_L g1256 ( 
.A1(n_941),
.A2(n_1022),
.A3(n_943),
.B(n_1019),
.Y(n_1256)
);

OAI21x1_ASAP7_75t_L g1257 ( 
.A1(n_958),
.A2(n_1121),
.B(n_949),
.Y(n_1257)
);

AOI21xp5_ASAP7_75t_L g1258 ( 
.A1(n_1129),
.A2(n_625),
.B(n_616),
.Y(n_1258)
);

AOI21xp5_ASAP7_75t_L g1259 ( 
.A1(n_1129),
.A2(n_625),
.B(n_616),
.Y(n_1259)
);

BUFx6f_ASAP7_75t_L g1260 ( 
.A(n_1001),
.Y(n_1260)
);

A2O1A1Ixp33_ASAP7_75t_L g1261 ( 
.A1(n_941),
.A2(n_947),
.B(n_959),
.C(n_1076),
.Y(n_1261)
);

OAI21xp5_ASAP7_75t_L g1262 ( 
.A1(n_941),
.A2(n_959),
.B(n_791),
.Y(n_1262)
);

AND2x2_ASAP7_75t_L g1263 ( 
.A(n_994),
.B(n_1052),
.Y(n_1263)
);

AO31x2_ASAP7_75t_L g1264 ( 
.A1(n_941),
.A2(n_1022),
.A3(n_943),
.B(n_1019),
.Y(n_1264)
);

AND2x2_ASAP7_75t_L g1265 ( 
.A(n_994),
.B(n_1052),
.Y(n_1265)
);

INVx1_ASAP7_75t_L g1266 ( 
.A(n_1115),
.Y(n_1266)
);

OAI21x1_ASAP7_75t_L g1267 ( 
.A1(n_958),
.A2(n_1121),
.B(n_949),
.Y(n_1267)
);

AND2x2_ASAP7_75t_L g1268 ( 
.A(n_994),
.B(n_1052),
.Y(n_1268)
);

INVx2_ASAP7_75t_L g1269 ( 
.A(n_939),
.Y(n_1269)
);

AOI21xp5_ASAP7_75t_L g1270 ( 
.A1(n_1129),
.A2(n_625),
.B(n_616),
.Y(n_1270)
);

OAI21x1_ASAP7_75t_L g1271 ( 
.A1(n_958),
.A2(n_1121),
.B(n_949),
.Y(n_1271)
);

NAND2xp5_ASAP7_75t_L g1272 ( 
.A(n_959),
.B(n_1077),
.Y(n_1272)
);

OR2x2_ASAP7_75t_L g1273 ( 
.A(n_990),
.B(n_836),
.Y(n_1273)
);

AO21x1_ASAP7_75t_L g1274 ( 
.A1(n_959),
.A2(n_947),
.B(n_943),
.Y(n_1274)
);

NAND2xp5_ASAP7_75t_L g1275 ( 
.A(n_959),
.B(n_1077),
.Y(n_1275)
);

INVxp67_ASAP7_75t_L g1276 ( 
.A(n_971),
.Y(n_1276)
);

NOR2xp33_ASAP7_75t_L g1277 ( 
.A(n_1017),
.B(n_1045),
.Y(n_1277)
);

OAI21x1_ASAP7_75t_L g1278 ( 
.A1(n_958),
.A2(n_1121),
.B(n_949),
.Y(n_1278)
);

AND2x2_ASAP7_75t_L g1279 ( 
.A(n_994),
.B(n_1052),
.Y(n_1279)
);

OAI21x1_ASAP7_75t_L g1280 ( 
.A1(n_958),
.A2(n_1121),
.B(n_949),
.Y(n_1280)
);

INVxp67_ASAP7_75t_L g1281 ( 
.A(n_971),
.Y(n_1281)
);

NAND2xp5_ASAP7_75t_L g1282 ( 
.A(n_959),
.B(n_1077),
.Y(n_1282)
);

NAND2xp5_ASAP7_75t_L g1283 ( 
.A(n_959),
.B(n_1077),
.Y(n_1283)
);

AOI21x1_ASAP7_75t_L g1284 ( 
.A1(n_949),
.A2(n_926),
.B(n_898),
.Y(n_1284)
);

OAI21x1_ASAP7_75t_L g1285 ( 
.A1(n_957),
.A2(n_960),
.B(n_942),
.Y(n_1285)
);

NAND2xp5_ASAP7_75t_L g1286 ( 
.A(n_959),
.B(n_1077),
.Y(n_1286)
);

NAND2xp5_ASAP7_75t_SL g1287 ( 
.A(n_941),
.B(n_959),
.Y(n_1287)
);

OAI21xp5_ASAP7_75t_L g1288 ( 
.A1(n_941),
.A2(n_959),
.B(n_791),
.Y(n_1288)
);

OAI21x1_ASAP7_75t_L g1289 ( 
.A1(n_958),
.A2(n_1121),
.B(n_949),
.Y(n_1289)
);

AOI22xp5_ASAP7_75t_L g1290 ( 
.A1(n_959),
.A2(n_767),
.B1(n_941),
.B2(n_1017),
.Y(n_1290)
);

OAI21x1_ASAP7_75t_L g1291 ( 
.A1(n_958),
.A2(n_1121),
.B(n_949),
.Y(n_1291)
);

A2O1A1Ixp33_ASAP7_75t_L g1292 ( 
.A1(n_941),
.A2(n_947),
.B(n_959),
.C(n_1076),
.Y(n_1292)
);

AND2x2_ASAP7_75t_L g1293 ( 
.A(n_994),
.B(n_1052),
.Y(n_1293)
);

AND2x4_ASAP7_75t_L g1294 ( 
.A(n_964),
.B(n_853),
.Y(n_1294)
);

NAND2xp5_ASAP7_75t_L g1295 ( 
.A(n_1290),
.B(n_1272),
.Y(n_1295)
);

AOI21xp5_ASAP7_75t_L g1296 ( 
.A1(n_1163),
.A2(n_1182),
.B(n_1130),
.Y(n_1296)
);

CKINVDCx5p33_ASAP7_75t_R g1297 ( 
.A(n_1153),
.Y(n_1297)
);

AND2x2_ASAP7_75t_L g1298 ( 
.A(n_1148),
.B(n_1159),
.Y(n_1298)
);

BUFx6f_ASAP7_75t_L g1299 ( 
.A(n_1138),
.Y(n_1299)
);

INVx4_ASAP7_75t_L g1300 ( 
.A(n_1138),
.Y(n_1300)
);

OAI221xp5_ASAP7_75t_L g1301 ( 
.A1(n_1156),
.A2(n_1140),
.B1(n_1261),
.B2(n_1292),
.C(n_1207),
.Y(n_1301)
);

AND2x4_ASAP7_75t_L g1302 ( 
.A(n_1152),
.B(n_1294),
.Y(n_1302)
);

NOR2xp33_ASAP7_75t_L g1303 ( 
.A(n_1275),
.B(n_1282),
.Y(n_1303)
);

INVx3_ASAP7_75t_L g1304 ( 
.A(n_1138),
.Y(n_1304)
);

INVx1_ASAP7_75t_L g1305 ( 
.A(n_1161),
.Y(n_1305)
);

OAI21xp33_ASAP7_75t_L g1306 ( 
.A1(n_1184),
.A2(n_1286),
.B(n_1283),
.Y(n_1306)
);

INVx2_ASAP7_75t_L g1307 ( 
.A(n_1193),
.Y(n_1307)
);

INVx2_ASAP7_75t_SL g1308 ( 
.A(n_1145),
.Y(n_1308)
);

AND2x2_ASAP7_75t_L g1309 ( 
.A(n_1131),
.B(n_1235),
.Y(n_1309)
);

BUFx10_ASAP7_75t_L g1310 ( 
.A(n_1153),
.Y(n_1310)
);

OAI22xp33_ASAP7_75t_L g1311 ( 
.A1(n_1144),
.A2(n_1191),
.B1(n_1273),
.B2(n_1216),
.Y(n_1311)
);

AOI21xp5_ASAP7_75t_L g1312 ( 
.A1(n_1135),
.A2(n_1287),
.B(n_1132),
.Y(n_1312)
);

BUFx2_ASAP7_75t_L g1313 ( 
.A(n_1248),
.Y(n_1313)
);

AOI22xp33_ASAP7_75t_L g1314 ( 
.A1(n_1221),
.A2(n_1226),
.B1(n_1274),
.B2(n_1244),
.Y(n_1314)
);

NAND2xp5_ASAP7_75t_L g1315 ( 
.A(n_1261),
.B(n_1292),
.Y(n_1315)
);

OR2x2_ASAP7_75t_L g1316 ( 
.A(n_1154),
.B(n_1158),
.Y(n_1316)
);

A2O1A1Ixp33_ASAP7_75t_L g1317 ( 
.A1(n_1241),
.A2(n_1262),
.B(n_1288),
.C(n_1252),
.Y(n_1317)
);

AND2x2_ASAP7_75t_L g1318 ( 
.A(n_1236),
.B(n_1263),
.Y(n_1318)
);

AND2x4_ASAP7_75t_L g1319 ( 
.A(n_1152),
.B(n_1294),
.Y(n_1319)
);

A2O1A1Ixp33_ASAP7_75t_SL g1320 ( 
.A1(n_1181),
.A2(n_1186),
.B(n_1214),
.C(n_1234),
.Y(n_1320)
);

AOI21xp5_ASAP7_75t_L g1321 ( 
.A1(n_1132),
.A2(n_1287),
.B(n_1164),
.Y(n_1321)
);

BUFx2_ASAP7_75t_L g1322 ( 
.A(n_1248),
.Y(n_1322)
);

CKINVDCx6p67_ASAP7_75t_R g1323 ( 
.A(n_1145),
.Y(n_1323)
);

AOI21xp5_ASAP7_75t_L g1324 ( 
.A1(n_1233),
.A2(n_1243),
.B(n_1259),
.Y(n_1324)
);

INVx2_ASAP7_75t_L g1325 ( 
.A(n_1269),
.Y(n_1325)
);

AND2x2_ASAP7_75t_L g1326 ( 
.A(n_1265),
.B(n_1268),
.Y(n_1326)
);

INVx2_ASAP7_75t_L g1327 ( 
.A(n_1142),
.Y(n_1327)
);

AOI21xp5_ASAP7_75t_L g1328 ( 
.A1(n_1249),
.A2(n_1258),
.B(n_1270),
.Y(n_1328)
);

AND2x2_ASAP7_75t_L g1329 ( 
.A(n_1279),
.B(n_1293),
.Y(n_1329)
);

NAND2xp5_ASAP7_75t_L g1330 ( 
.A(n_1234),
.B(n_1277),
.Y(n_1330)
);

AND2x4_ASAP7_75t_L g1331 ( 
.A(n_1152),
.B(n_1294),
.Y(n_1331)
);

BUFx2_ASAP7_75t_L g1332 ( 
.A(n_1178),
.Y(n_1332)
);

AND2x4_ASAP7_75t_L g1333 ( 
.A(n_1185),
.B(n_1174),
.Y(n_1333)
);

AOI22xp33_ASAP7_75t_L g1334 ( 
.A1(n_1221),
.A2(n_1187),
.B1(n_1223),
.B2(n_1139),
.Y(n_1334)
);

HB1xp67_ASAP7_75t_L g1335 ( 
.A(n_1227),
.Y(n_1335)
);

AND2x2_ASAP7_75t_L g1336 ( 
.A(n_1189),
.B(n_1213),
.Y(n_1336)
);

INVx2_ASAP7_75t_L g1337 ( 
.A(n_1143),
.Y(n_1337)
);

AOI22xp33_ASAP7_75t_SL g1338 ( 
.A1(n_1205),
.A2(n_1277),
.B1(n_1166),
.B2(n_1208),
.Y(n_1338)
);

INVx2_ASAP7_75t_L g1339 ( 
.A(n_1232),
.Y(n_1339)
);

OAI21x1_ASAP7_75t_L g1340 ( 
.A1(n_1177),
.A2(n_1175),
.B(n_1203),
.Y(n_1340)
);

INVx1_ASAP7_75t_L g1341 ( 
.A(n_1266),
.Y(n_1341)
);

BUFx6f_ASAP7_75t_L g1342 ( 
.A(n_1149),
.Y(n_1342)
);

AOI21xp5_ASAP7_75t_L g1343 ( 
.A1(n_1176),
.A2(n_1168),
.B(n_1204),
.Y(n_1343)
);

INVx4_ASAP7_75t_L g1344 ( 
.A(n_1149),
.Y(n_1344)
);

INVx3_ASAP7_75t_SL g1345 ( 
.A(n_1197),
.Y(n_1345)
);

AOI22xp33_ASAP7_75t_L g1346 ( 
.A1(n_1223),
.A2(n_1139),
.B1(n_1239),
.B2(n_1167),
.Y(n_1346)
);

BUFx6f_ASAP7_75t_L g1347 ( 
.A(n_1149),
.Y(n_1347)
);

INVx3_ASAP7_75t_L g1348 ( 
.A(n_1253),
.Y(n_1348)
);

BUFx4_ASAP7_75t_SL g1349 ( 
.A(n_1197),
.Y(n_1349)
);

NOR2xp33_ASAP7_75t_SL g1350 ( 
.A(n_1207),
.B(n_1209),
.Y(n_1350)
);

BUFx2_ASAP7_75t_R g1351 ( 
.A(n_1185),
.Y(n_1351)
);

INVx1_ASAP7_75t_SL g1352 ( 
.A(n_1136),
.Y(n_1352)
);

NOR2xp33_ASAP7_75t_L g1353 ( 
.A(n_1141),
.B(n_1157),
.Y(n_1353)
);

O2A1O1Ixp5_ASAP7_75t_L g1354 ( 
.A1(n_1211),
.A2(n_1133),
.B(n_1134),
.C(n_1217),
.Y(n_1354)
);

BUFx2_ASAP7_75t_L g1355 ( 
.A(n_1242),
.Y(n_1355)
);

NAND2xp5_ASAP7_75t_L g1356 ( 
.A(n_1162),
.B(n_1200),
.Y(n_1356)
);

O2A1O1Ixp33_ASAP7_75t_L g1357 ( 
.A1(n_1222),
.A2(n_1146),
.B(n_1276),
.C(n_1281),
.Y(n_1357)
);

NOR2xp67_ASAP7_75t_R g1358 ( 
.A(n_1179),
.B(n_1225),
.Y(n_1358)
);

OAI22xp5_ASAP7_75t_L g1359 ( 
.A1(n_1169),
.A2(n_1239),
.B1(n_1225),
.B2(n_1190),
.Y(n_1359)
);

INVx1_ASAP7_75t_L g1360 ( 
.A(n_1171),
.Y(n_1360)
);

INVx1_ASAP7_75t_L g1361 ( 
.A(n_1150),
.Y(n_1361)
);

OR2x6_ASAP7_75t_L g1362 ( 
.A(n_1225),
.B(n_1179),
.Y(n_1362)
);

NAND2xp5_ASAP7_75t_L g1363 ( 
.A(n_1147),
.B(n_1264),
.Y(n_1363)
);

INVx1_ASAP7_75t_SL g1364 ( 
.A(n_1166),
.Y(n_1364)
);

BUFx2_ASAP7_75t_SL g1365 ( 
.A(n_1199),
.Y(n_1365)
);

AOI21xp33_ASAP7_75t_SL g1366 ( 
.A1(n_1220),
.A2(n_1228),
.B(n_1219),
.Y(n_1366)
);

BUFx6f_ASAP7_75t_L g1367 ( 
.A(n_1253),
.Y(n_1367)
);

AOI21xp5_ASAP7_75t_L g1368 ( 
.A1(n_1204),
.A2(n_1194),
.B(n_1155),
.Y(n_1368)
);

AND2x4_ASAP7_75t_L g1369 ( 
.A(n_1206),
.B(n_1173),
.Y(n_1369)
);

BUFx2_ASAP7_75t_L g1370 ( 
.A(n_1253),
.Y(n_1370)
);

AND2x2_ASAP7_75t_L g1371 ( 
.A(n_1199),
.B(n_1230),
.Y(n_1371)
);

OAI22xp5_ASAP7_75t_L g1372 ( 
.A1(n_1225),
.A2(n_1212),
.B1(n_1195),
.B2(n_1183),
.Y(n_1372)
);

INVx3_ASAP7_75t_SL g1373 ( 
.A(n_1199),
.Y(n_1373)
);

INVx2_ASAP7_75t_L g1374 ( 
.A(n_1173),
.Y(n_1374)
);

OAI22xp33_ASAP7_75t_L g1375 ( 
.A1(n_1212),
.A2(n_1180),
.B1(n_1204),
.B2(n_1198),
.Y(n_1375)
);

AOI22xp33_ASAP7_75t_L g1376 ( 
.A1(n_1219),
.A2(n_1137),
.B1(n_1220),
.B2(n_1228),
.Y(n_1376)
);

NAND2xp5_ASAP7_75t_L g1377 ( 
.A(n_1147),
.B(n_1264),
.Y(n_1377)
);

CKINVDCx11_ASAP7_75t_R g1378 ( 
.A(n_1253),
.Y(n_1378)
);

AND2x4_ASAP7_75t_L g1379 ( 
.A(n_1260),
.B(n_1229),
.Y(n_1379)
);

AOI21xp5_ASAP7_75t_L g1380 ( 
.A1(n_1170),
.A2(n_1137),
.B(n_1196),
.Y(n_1380)
);

NAND3xp33_ASAP7_75t_L g1381 ( 
.A(n_1202),
.B(n_1201),
.C(n_1260),
.Y(n_1381)
);

INVx1_ASAP7_75t_SL g1382 ( 
.A(n_1260),
.Y(n_1382)
);

NAND2xp5_ASAP7_75t_SL g1383 ( 
.A(n_1183),
.B(n_1260),
.Y(n_1383)
);

AOI21xp5_ASAP7_75t_L g1384 ( 
.A1(n_1231),
.A2(n_1245),
.B(n_1289),
.Y(n_1384)
);

OR2x2_ASAP7_75t_L g1385 ( 
.A(n_1147),
.B(n_1230),
.Y(n_1385)
);

NAND2xp5_ASAP7_75t_L g1386 ( 
.A(n_1147),
.B(n_1264),
.Y(n_1386)
);

INVx1_ASAP7_75t_L g1387 ( 
.A(n_1183),
.Y(n_1387)
);

A2O1A1Ixp33_ASAP7_75t_L g1388 ( 
.A1(n_1215),
.A2(n_1224),
.B(n_1218),
.C(n_1229),
.Y(n_1388)
);

OR2x6_ASAP7_75t_L g1389 ( 
.A(n_1183),
.B(n_1224),
.Y(n_1389)
);

A2O1A1Ixp33_ASAP7_75t_SL g1390 ( 
.A1(n_1210),
.A2(n_1264),
.B(n_1256),
.C(n_1230),
.Y(n_1390)
);

CKINVDCx20_ASAP7_75t_R g1391 ( 
.A(n_1230),
.Y(n_1391)
);

NOR2x1_ASAP7_75t_SL g1392 ( 
.A(n_1247),
.B(n_1250),
.Y(n_1392)
);

A2O1A1Ixp33_ASAP7_75t_L g1393 ( 
.A1(n_1215),
.A2(n_1218),
.B(n_1210),
.C(n_1291),
.Y(n_1393)
);

OAI22xp33_ASAP7_75t_L g1394 ( 
.A1(n_1284),
.A2(n_1192),
.B1(n_1256),
.B2(n_1151),
.Y(n_1394)
);

NAND2xp5_ASAP7_75t_L g1395 ( 
.A(n_1256),
.B(n_1192),
.Y(n_1395)
);

O2A1O1Ixp33_ASAP7_75t_L g1396 ( 
.A1(n_1256),
.A2(n_1192),
.B(n_1291),
.C(n_1251),
.Y(n_1396)
);

NOR2xp33_ASAP7_75t_L g1397 ( 
.A(n_1175),
.B(n_1246),
.Y(n_1397)
);

CKINVDCx20_ASAP7_75t_R g1398 ( 
.A(n_1192),
.Y(n_1398)
);

OAI21x1_ASAP7_75t_L g1399 ( 
.A1(n_1177),
.A2(n_1285),
.B(n_1172),
.Y(n_1399)
);

AOI21xp33_ASAP7_75t_SL g1400 ( 
.A1(n_1237),
.A2(n_1254),
.B(n_1280),
.Y(n_1400)
);

AOI22xp33_ASAP7_75t_L g1401 ( 
.A1(n_1237),
.A2(n_1254),
.B1(n_1280),
.B2(n_1278),
.Y(n_1401)
);

CKINVDCx5p33_ASAP7_75t_R g1402 ( 
.A(n_1238),
.Y(n_1402)
);

INVx3_ASAP7_75t_SL g1403 ( 
.A(n_1240),
.Y(n_1403)
);

CKINVDCx11_ASAP7_75t_R g1404 ( 
.A(n_1289),
.Y(n_1404)
);

AOI22xp33_ASAP7_75t_L g1405 ( 
.A1(n_1245),
.A2(n_1255),
.B1(n_1271),
.B2(n_1267),
.Y(n_1405)
);

AOI21xp5_ASAP7_75t_L g1406 ( 
.A1(n_1246),
.A2(n_1257),
.B(n_1267),
.Y(n_1406)
);

AOI22xp33_ASAP7_75t_L g1407 ( 
.A1(n_1257),
.A2(n_1271),
.B1(n_1278),
.B2(n_1160),
.Y(n_1407)
);

AO21x1_ASAP7_75t_L g1408 ( 
.A1(n_1172),
.A2(n_1241),
.B(n_959),
.Y(n_1408)
);

AOI21xp5_ASAP7_75t_L g1409 ( 
.A1(n_1188),
.A2(n_1163),
.B(n_1129),
.Y(n_1409)
);

OAI21xp5_ASAP7_75t_L g1410 ( 
.A1(n_1252),
.A2(n_941),
.B(n_1262),
.Y(n_1410)
);

INVx2_ASAP7_75t_L g1411 ( 
.A(n_1165),
.Y(n_1411)
);

AND2x4_ASAP7_75t_L g1412 ( 
.A(n_1152),
.B(n_1294),
.Y(n_1412)
);

BUFx8_ASAP7_75t_SL g1413 ( 
.A(n_1197),
.Y(n_1413)
);

AOI21xp5_ASAP7_75t_L g1414 ( 
.A1(n_1163),
.A2(n_1129),
.B(n_1182),
.Y(n_1414)
);

OAI22xp5_ASAP7_75t_L g1415 ( 
.A1(n_1261),
.A2(n_941),
.B1(n_947),
.B2(n_802),
.Y(n_1415)
);

INVx3_ASAP7_75t_L g1416 ( 
.A(n_1138),
.Y(n_1416)
);

AOI21xp5_ASAP7_75t_L g1417 ( 
.A1(n_1163),
.A2(n_1129),
.B(n_1182),
.Y(n_1417)
);

NAND2xp5_ASAP7_75t_SL g1418 ( 
.A(n_1131),
.B(n_994),
.Y(n_1418)
);

INVx2_ASAP7_75t_L g1419 ( 
.A(n_1165),
.Y(n_1419)
);

NOR2xp67_ASAP7_75t_L g1420 ( 
.A(n_1273),
.B(n_777),
.Y(n_1420)
);

INVx5_ASAP7_75t_L g1421 ( 
.A(n_1225),
.Y(n_1421)
);

NOR2xp33_ASAP7_75t_L g1422 ( 
.A(n_1159),
.B(n_928),
.Y(n_1422)
);

OR2x2_ASAP7_75t_L g1423 ( 
.A(n_1154),
.B(n_1273),
.Y(n_1423)
);

AND2x2_ASAP7_75t_SL g1424 ( 
.A(n_1156),
.B(n_1223),
.Y(n_1424)
);

AOI21xp5_ASAP7_75t_L g1425 ( 
.A1(n_1163),
.A2(n_1129),
.B(n_1182),
.Y(n_1425)
);

AOI21xp5_ASAP7_75t_L g1426 ( 
.A1(n_1163),
.A2(n_1129),
.B(n_1182),
.Y(n_1426)
);

AOI21xp5_ASAP7_75t_L g1427 ( 
.A1(n_1182),
.A2(n_1129),
.B(n_1163),
.Y(n_1427)
);

AND2x2_ASAP7_75t_L g1428 ( 
.A(n_1148),
.B(n_1159),
.Y(n_1428)
);

AND2x4_ASAP7_75t_L g1429 ( 
.A(n_1152),
.B(n_1294),
.Y(n_1429)
);

INVx5_ASAP7_75t_L g1430 ( 
.A(n_1225),
.Y(n_1430)
);

BUFx6f_ASAP7_75t_L g1431 ( 
.A(n_1138),
.Y(n_1431)
);

INVx2_ASAP7_75t_L g1432 ( 
.A(n_1165),
.Y(n_1432)
);

AND2x2_ASAP7_75t_SL g1433 ( 
.A(n_1156),
.B(n_1223),
.Y(n_1433)
);

AOI22xp33_ASAP7_75t_SL g1434 ( 
.A1(n_1159),
.A2(n_623),
.B1(n_994),
.B2(n_1039),
.Y(n_1434)
);

HB1xp67_ASAP7_75t_L g1435 ( 
.A(n_1248),
.Y(n_1435)
);

INVx3_ASAP7_75t_L g1436 ( 
.A(n_1138),
.Y(n_1436)
);

NOR2xp33_ASAP7_75t_L g1437 ( 
.A(n_1159),
.B(n_928),
.Y(n_1437)
);

INVx1_ASAP7_75t_L g1438 ( 
.A(n_1161),
.Y(n_1438)
);

INVx1_ASAP7_75t_L g1439 ( 
.A(n_1161),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_1161),
.Y(n_1440)
);

INVx1_ASAP7_75t_SL g1441 ( 
.A(n_1154),
.Y(n_1441)
);

INVx1_ASAP7_75t_SL g1442 ( 
.A(n_1154),
.Y(n_1442)
);

INVx8_ASAP7_75t_L g1443 ( 
.A(n_1152),
.Y(n_1443)
);

BUFx2_ASAP7_75t_R g1444 ( 
.A(n_1153),
.Y(n_1444)
);

AOI21xp5_ASAP7_75t_L g1445 ( 
.A1(n_1163),
.A2(n_1129),
.B(n_1182),
.Y(n_1445)
);

CKINVDCx8_ASAP7_75t_R g1446 ( 
.A(n_1153),
.Y(n_1446)
);

AND2x4_ASAP7_75t_L g1447 ( 
.A(n_1152),
.B(n_1294),
.Y(n_1447)
);

INVx1_ASAP7_75t_L g1448 ( 
.A(n_1161),
.Y(n_1448)
);

INVx1_ASAP7_75t_L g1449 ( 
.A(n_1161),
.Y(n_1449)
);

INVx2_ASAP7_75t_L g1450 ( 
.A(n_1165),
.Y(n_1450)
);

AOI21xp5_ASAP7_75t_L g1451 ( 
.A1(n_1163),
.A2(n_1129),
.B(n_1182),
.Y(n_1451)
);

AND2x4_ASAP7_75t_L g1452 ( 
.A(n_1152),
.B(n_1294),
.Y(n_1452)
);

BUFx12f_ASAP7_75t_L g1453 ( 
.A(n_1153),
.Y(n_1453)
);

NAND2xp5_ASAP7_75t_L g1454 ( 
.A(n_1290),
.B(n_959),
.Y(n_1454)
);

NAND2xp5_ASAP7_75t_L g1455 ( 
.A(n_1290),
.B(n_959),
.Y(n_1455)
);

HB1xp67_ASAP7_75t_L g1456 ( 
.A(n_1248),
.Y(n_1456)
);

BUFx2_ASAP7_75t_L g1457 ( 
.A(n_1248),
.Y(n_1457)
);

OA21x2_ASAP7_75t_L g1458 ( 
.A1(n_1393),
.A2(n_1368),
.B(n_1354),
.Y(n_1458)
);

INVx1_ASAP7_75t_L g1459 ( 
.A(n_1360),
.Y(n_1459)
);

NAND2x1p5_ASAP7_75t_L g1460 ( 
.A(n_1421),
.B(n_1430),
.Y(n_1460)
);

NAND2x1p5_ASAP7_75t_L g1461 ( 
.A(n_1421),
.B(n_1430),
.Y(n_1461)
);

INVx2_ASAP7_75t_SL g1462 ( 
.A(n_1349),
.Y(n_1462)
);

INVx1_ASAP7_75t_L g1463 ( 
.A(n_1341),
.Y(n_1463)
);

INVx2_ASAP7_75t_SL g1464 ( 
.A(n_1323),
.Y(n_1464)
);

OR2x2_ASAP7_75t_L g1465 ( 
.A(n_1316),
.B(n_1423),
.Y(n_1465)
);

CKINVDCx20_ASAP7_75t_R g1466 ( 
.A(n_1413),
.Y(n_1466)
);

INVx1_ASAP7_75t_SL g1467 ( 
.A(n_1332),
.Y(n_1467)
);

BUFx3_ASAP7_75t_L g1468 ( 
.A(n_1443),
.Y(n_1468)
);

AND2x4_ASAP7_75t_L g1469 ( 
.A(n_1302),
.B(n_1319),
.Y(n_1469)
);

INVx5_ASAP7_75t_L g1470 ( 
.A(n_1362),
.Y(n_1470)
);

AND2x4_ASAP7_75t_L g1471 ( 
.A(n_1302),
.B(n_1319),
.Y(n_1471)
);

INVx1_ASAP7_75t_L g1472 ( 
.A(n_1361),
.Y(n_1472)
);

INVx1_ASAP7_75t_L g1473 ( 
.A(n_1307),
.Y(n_1473)
);

NAND2x1p5_ASAP7_75t_L g1474 ( 
.A(n_1421),
.B(n_1430),
.Y(n_1474)
);

NAND2xp5_ASAP7_75t_L g1475 ( 
.A(n_1303),
.B(n_1298),
.Y(n_1475)
);

CKINVDCx11_ASAP7_75t_R g1476 ( 
.A(n_1446),
.Y(n_1476)
);

AOI22xp33_ASAP7_75t_L g1477 ( 
.A1(n_1424),
.A2(n_1433),
.B1(n_1301),
.B2(n_1415),
.Y(n_1477)
);

INVx1_ASAP7_75t_L g1478 ( 
.A(n_1325),
.Y(n_1478)
);

CKINVDCx11_ASAP7_75t_R g1479 ( 
.A(n_1453),
.Y(n_1479)
);

INVxp67_ASAP7_75t_L g1480 ( 
.A(n_1335),
.Y(n_1480)
);

OAI21xp5_ASAP7_75t_L g1481 ( 
.A1(n_1434),
.A2(n_1317),
.B(n_1301),
.Y(n_1481)
);

CKINVDCx5p33_ASAP7_75t_R g1482 ( 
.A(n_1297),
.Y(n_1482)
);

HB1xp67_ASAP7_75t_L g1483 ( 
.A(n_1441),
.Y(n_1483)
);

BUFx2_ASAP7_75t_R g1484 ( 
.A(n_1345),
.Y(n_1484)
);

INVx1_ASAP7_75t_L g1485 ( 
.A(n_1411),
.Y(n_1485)
);

INVx1_ASAP7_75t_L g1486 ( 
.A(n_1419),
.Y(n_1486)
);

OAI22xp5_ASAP7_75t_L g1487 ( 
.A1(n_1422),
.A2(n_1437),
.B1(n_1334),
.B2(n_1338),
.Y(n_1487)
);

INVx1_ASAP7_75t_L g1488 ( 
.A(n_1432),
.Y(n_1488)
);

NAND2xp5_ASAP7_75t_L g1489 ( 
.A(n_1428),
.B(n_1306),
.Y(n_1489)
);

INVx1_ASAP7_75t_L g1490 ( 
.A(n_1450),
.Y(n_1490)
);

AND2x2_ASAP7_75t_L g1491 ( 
.A(n_1336),
.B(n_1309),
.Y(n_1491)
);

BUFx2_ASAP7_75t_R g1492 ( 
.A(n_1373),
.Y(n_1492)
);

AO21x1_ASAP7_75t_SL g1493 ( 
.A1(n_1314),
.A2(n_1346),
.B(n_1363),
.Y(n_1493)
);

OAI22xp5_ASAP7_75t_L g1494 ( 
.A1(n_1330),
.A2(n_1352),
.B1(n_1356),
.B2(n_1418),
.Y(n_1494)
);

HB1xp67_ASAP7_75t_L g1495 ( 
.A(n_1441),
.Y(n_1495)
);

OAI22xp5_ASAP7_75t_L g1496 ( 
.A1(n_1330),
.A2(n_1352),
.B1(n_1356),
.B2(n_1438),
.Y(n_1496)
);

INVx1_ASAP7_75t_L g1497 ( 
.A(n_1327),
.Y(n_1497)
);

CKINVDCx20_ASAP7_75t_R g1498 ( 
.A(n_1378),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_1337),
.Y(n_1499)
);

INVx1_ASAP7_75t_L g1500 ( 
.A(n_1339),
.Y(n_1500)
);

INVx2_ASAP7_75t_SL g1501 ( 
.A(n_1308),
.Y(n_1501)
);

CKINVDCx6p67_ASAP7_75t_R g1502 ( 
.A(n_1310),
.Y(n_1502)
);

AO21x1_ASAP7_75t_SL g1503 ( 
.A1(n_1363),
.A2(n_1377),
.B(n_1386),
.Y(n_1503)
);

OAI21x1_ASAP7_75t_L g1504 ( 
.A1(n_1340),
.A2(n_1399),
.B(n_1409),
.Y(n_1504)
);

AND2x4_ASAP7_75t_L g1505 ( 
.A(n_1331),
.B(n_1412),
.Y(n_1505)
);

AOI22xp5_ASAP7_75t_L g1506 ( 
.A1(n_1350),
.A2(n_1420),
.B1(n_1326),
.B2(n_1329),
.Y(n_1506)
);

INVx1_ASAP7_75t_L g1507 ( 
.A(n_1305),
.Y(n_1507)
);

NAND2xp5_ASAP7_75t_L g1508 ( 
.A(n_1439),
.B(n_1440),
.Y(n_1508)
);

AND2x2_ASAP7_75t_L g1509 ( 
.A(n_1318),
.B(n_1442),
.Y(n_1509)
);

AO21x1_ASAP7_75t_SL g1510 ( 
.A1(n_1377),
.A2(n_1386),
.B(n_1315),
.Y(n_1510)
);

AOI22xp33_ASAP7_75t_L g1511 ( 
.A1(n_1415),
.A2(n_1350),
.B1(n_1410),
.B2(n_1454),
.Y(n_1511)
);

INVx5_ASAP7_75t_L g1512 ( 
.A(n_1362),
.Y(n_1512)
);

BUFx6f_ASAP7_75t_L g1513 ( 
.A(n_1443),
.Y(n_1513)
);

AOI222xp33_ASAP7_75t_L g1514 ( 
.A1(n_1410),
.A2(n_1455),
.B1(n_1454),
.B2(n_1315),
.C1(n_1311),
.C2(n_1295),
.Y(n_1514)
);

INVx3_ASAP7_75t_L g1515 ( 
.A(n_1443),
.Y(n_1515)
);

CKINVDCx20_ASAP7_75t_R g1516 ( 
.A(n_1310),
.Y(n_1516)
);

HB1xp67_ASAP7_75t_L g1517 ( 
.A(n_1442),
.Y(n_1517)
);

OAI22xp5_ASAP7_75t_L g1518 ( 
.A1(n_1448),
.A2(n_1449),
.B1(n_1295),
.B2(n_1455),
.Y(n_1518)
);

INVx6_ASAP7_75t_L g1519 ( 
.A(n_1421),
.Y(n_1519)
);

NOR2xp33_ASAP7_75t_L g1520 ( 
.A(n_1355),
.B(n_1353),
.Y(n_1520)
);

NOR2x1_ASAP7_75t_L g1521 ( 
.A(n_1365),
.B(n_1362),
.Y(n_1521)
);

AOI21x1_ASAP7_75t_L g1522 ( 
.A1(n_1414),
.A2(n_1425),
.B(n_1426),
.Y(n_1522)
);

OAI21x1_ASAP7_75t_L g1523 ( 
.A1(n_1409),
.A2(n_1296),
.B(n_1328),
.Y(n_1523)
);

AOI22xp33_ASAP7_75t_SL g1524 ( 
.A1(n_1398),
.A2(n_1391),
.B1(n_1359),
.B2(n_1371),
.Y(n_1524)
);

INVx2_ASAP7_75t_L g1525 ( 
.A(n_1392),
.Y(n_1525)
);

OAI22xp33_ASAP7_75t_L g1526 ( 
.A1(n_1435),
.A2(n_1456),
.B1(n_1313),
.B2(n_1457),
.Y(n_1526)
);

INVx2_ASAP7_75t_L g1527 ( 
.A(n_1389),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_1374),
.Y(n_1528)
);

INVx1_ASAP7_75t_L g1529 ( 
.A(n_1357),
.Y(n_1529)
);

INVx1_ASAP7_75t_L g1530 ( 
.A(n_1322),
.Y(n_1530)
);

BUFx12f_ASAP7_75t_L g1531 ( 
.A(n_1333),
.Y(n_1531)
);

BUFx2_ASAP7_75t_L g1532 ( 
.A(n_1370),
.Y(n_1532)
);

HB1xp67_ASAP7_75t_L g1533 ( 
.A(n_1387),
.Y(n_1533)
);

INVx2_ASAP7_75t_L g1534 ( 
.A(n_1389),
.Y(n_1534)
);

BUFx2_ASAP7_75t_L g1535 ( 
.A(n_1331),
.Y(n_1535)
);

BUFx4f_ASAP7_75t_SL g1536 ( 
.A(n_1364),
.Y(n_1536)
);

HB1xp67_ASAP7_75t_L g1537 ( 
.A(n_1412),
.Y(n_1537)
);

NAND2xp5_ASAP7_75t_L g1538 ( 
.A(n_1452),
.B(n_1429),
.Y(n_1538)
);

AND2x2_ASAP7_75t_L g1539 ( 
.A(n_1429),
.B(n_1447),
.Y(n_1539)
);

OA21x2_ASAP7_75t_L g1540 ( 
.A1(n_1368),
.A2(n_1388),
.B(n_1343),
.Y(n_1540)
);

AOI21x1_ASAP7_75t_L g1541 ( 
.A1(n_1417),
.A2(n_1451),
.B(n_1445),
.Y(n_1541)
);

INVx2_ASAP7_75t_L g1542 ( 
.A(n_1389),
.Y(n_1542)
);

AOI22xp33_ASAP7_75t_L g1543 ( 
.A1(n_1359),
.A2(n_1408),
.B1(n_1321),
.B2(n_1312),
.Y(n_1543)
);

INVx1_ASAP7_75t_L g1544 ( 
.A(n_1304),
.Y(n_1544)
);

OAI21x1_ASAP7_75t_L g1545 ( 
.A1(n_1296),
.A2(n_1328),
.B(n_1324),
.Y(n_1545)
);

CKINVDCx6p67_ASAP7_75t_R g1546 ( 
.A(n_1364),
.Y(n_1546)
);

HB1xp67_ASAP7_75t_L g1547 ( 
.A(n_1447),
.Y(n_1547)
);

AOI21x1_ASAP7_75t_L g1548 ( 
.A1(n_1425),
.A2(n_1426),
.B(n_1451),
.Y(n_1548)
);

BUFx6f_ASAP7_75t_L g1549 ( 
.A(n_1452),
.Y(n_1549)
);

BUFx6f_ASAP7_75t_L g1550 ( 
.A(n_1299),
.Y(n_1550)
);

AOI22xp33_ASAP7_75t_L g1551 ( 
.A1(n_1321),
.A2(n_1312),
.B1(n_1395),
.B2(n_1404),
.Y(n_1551)
);

INVx2_ASAP7_75t_L g1552 ( 
.A(n_1403),
.Y(n_1552)
);

INVx1_ASAP7_75t_L g1553 ( 
.A(n_1348),
.Y(n_1553)
);

AOI22xp33_ASAP7_75t_L g1554 ( 
.A1(n_1395),
.A2(n_1385),
.B1(n_1343),
.B2(n_1402),
.Y(n_1554)
);

CKINVDCx11_ASAP7_75t_R g1555 ( 
.A(n_1444),
.Y(n_1555)
);

OAI22xp33_ASAP7_75t_L g1556 ( 
.A1(n_1430),
.A2(n_1372),
.B1(n_1445),
.B2(n_1427),
.Y(n_1556)
);

OAI22xp5_ASAP7_75t_L g1557 ( 
.A1(n_1351),
.A2(n_1333),
.B1(n_1372),
.B2(n_1376),
.Y(n_1557)
);

CKINVDCx20_ASAP7_75t_R g1558 ( 
.A(n_1444),
.Y(n_1558)
);

BUFx3_ASAP7_75t_L g1559 ( 
.A(n_1299),
.Y(n_1559)
);

AOI22xp33_ASAP7_75t_SL g1560 ( 
.A1(n_1351),
.A2(n_1369),
.B1(n_1381),
.B2(n_1379),
.Y(n_1560)
);

AOI21x1_ASAP7_75t_L g1561 ( 
.A1(n_1380),
.A2(n_1406),
.B(n_1384),
.Y(n_1561)
);

INVx6_ASAP7_75t_L g1562 ( 
.A(n_1300),
.Y(n_1562)
);

AOI21xp33_ASAP7_75t_L g1563 ( 
.A1(n_1320),
.A2(n_1390),
.B(n_1375),
.Y(n_1563)
);

INVx2_ASAP7_75t_L g1564 ( 
.A(n_1379),
.Y(n_1564)
);

INVx1_ASAP7_75t_L g1565 ( 
.A(n_1348),
.Y(n_1565)
);

AOI22xp33_ASAP7_75t_L g1566 ( 
.A1(n_1394),
.A2(n_1397),
.B1(n_1369),
.B2(n_1407),
.Y(n_1566)
);

AOI22xp33_ASAP7_75t_SL g1567 ( 
.A1(n_1382),
.A2(n_1436),
.B1(n_1416),
.B2(n_1300),
.Y(n_1567)
);

AOI22xp33_ASAP7_75t_SL g1568 ( 
.A1(n_1382),
.A2(n_1436),
.B1(n_1416),
.B2(n_1344),
.Y(n_1568)
);

INVx2_ASAP7_75t_L g1569 ( 
.A(n_1299),
.Y(n_1569)
);

AOI22xp33_ASAP7_75t_L g1570 ( 
.A1(n_1401),
.A2(n_1405),
.B1(n_1406),
.B2(n_1324),
.Y(n_1570)
);

AOI22xp33_ASAP7_75t_L g1571 ( 
.A1(n_1383),
.A2(n_1344),
.B1(n_1342),
.B2(n_1347),
.Y(n_1571)
);

AO21x2_ASAP7_75t_L g1572 ( 
.A1(n_1366),
.A2(n_1400),
.B(n_1396),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_1342),
.Y(n_1573)
);

BUFx3_ASAP7_75t_L g1574 ( 
.A(n_1347),
.Y(n_1574)
);

HB1xp67_ASAP7_75t_L g1575 ( 
.A(n_1367),
.Y(n_1575)
);

INVx1_ASAP7_75t_L g1576 ( 
.A(n_1431),
.Y(n_1576)
);

INVx6_ASAP7_75t_L g1577 ( 
.A(n_1367),
.Y(n_1577)
);

AOI22xp33_ASAP7_75t_L g1578 ( 
.A1(n_1367),
.A2(n_1424),
.B1(n_1433),
.B2(n_1156),
.Y(n_1578)
);

INVx1_ASAP7_75t_L g1579 ( 
.A(n_1358),
.Y(n_1579)
);

CKINVDCx5p33_ASAP7_75t_R g1580 ( 
.A(n_1413),
.Y(n_1580)
);

BUFx6f_ASAP7_75t_L g1581 ( 
.A(n_1378),
.Y(n_1581)
);

BUFx3_ASAP7_75t_L g1582 ( 
.A(n_1332),
.Y(n_1582)
);

AOI22xp33_ASAP7_75t_SL g1583 ( 
.A1(n_1350),
.A2(n_1433),
.B1(n_1424),
.B2(n_1118),
.Y(n_1583)
);

NAND2x1p5_ASAP7_75t_L g1584 ( 
.A(n_1421),
.B(n_1430),
.Y(n_1584)
);

HB1xp67_ASAP7_75t_L g1585 ( 
.A(n_1335),
.Y(n_1585)
);

INVx6_ASAP7_75t_L g1586 ( 
.A(n_1443),
.Y(n_1586)
);

INVx3_ASAP7_75t_L g1587 ( 
.A(n_1443),
.Y(n_1587)
);

OA21x2_ASAP7_75t_L g1588 ( 
.A1(n_1393),
.A2(n_1368),
.B(n_1354),
.Y(n_1588)
);

INVx1_ASAP7_75t_L g1589 ( 
.A(n_1360),
.Y(n_1589)
);

CKINVDCx5p33_ASAP7_75t_R g1590 ( 
.A(n_1413),
.Y(n_1590)
);

OAI22xp33_ASAP7_75t_R g1591 ( 
.A1(n_1422),
.A2(n_421),
.B1(n_535),
.B2(n_269),
.Y(n_1591)
);

AOI21xp5_ASAP7_75t_L g1592 ( 
.A1(n_1414),
.A2(n_1425),
.B(n_1417),
.Y(n_1592)
);

BUFx2_ASAP7_75t_L g1593 ( 
.A(n_1332),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_1360),
.Y(n_1594)
);

BUFx4f_ASAP7_75t_L g1595 ( 
.A(n_1453),
.Y(n_1595)
);

AOI22xp33_ASAP7_75t_L g1596 ( 
.A1(n_1424),
.A2(n_1433),
.B1(n_1156),
.B2(n_1140),
.Y(n_1596)
);

OAI22xp5_ASAP7_75t_L g1597 ( 
.A1(n_1434),
.A2(n_941),
.B1(n_959),
.B2(n_767),
.Y(n_1597)
);

NAND3xp33_ASAP7_75t_L g1598 ( 
.A(n_1434),
.B(n_959),
.C(n_1156),
.Y(n_1598)
);

CKINVDCx14_ASAP7_75t_R g1599 ( 
.A(n_1297),
.Y(n_1599)
);

OAI21x1_ASAP7_75t_L g1600 ( 
.A1(n_1340),
.A2(n_1399),
.B(n_1409),
.Y(n_1600)
);

NAND2xp5_ASAP7_75t_L g1601 ( 
.A(n_1303),
.B(n_1298),
.Y(n_1601)
);

INVx1_ASAP7_75t_L g1602 ( 
.A(n_1360),
.Y(n_1602)
);

OAI21xp5_ASAP7_75t_L g1603 ( 
.A1(n_1434),
.A2(n_941),
.B(n_959),
.Y(n_1603)
);

INVx2_ASAP7_75t_SL g1604 ( 
.A(n_1483),
.Y(n_1604)
);

NAND2xp5_ASAP7_75t_L g1605 ( 
.A(n_1465),
.B(n_1494),
.Y(n_1605)
);

AND2x2_ASAP7_75t_L g1606 ( 
.A(n_1510),
.B(n_1564),
.Y(n_1606)
);

HB1xp67_ASAP7_75t_L g1607 ( 
.A(n_1495),
.Y(n_1607)
);

AO21x2_ASAP7_75t_L g1608 ( 
.A1(n_1563),
.A2(n_1592),
.B(n_1541),
.Y(n_1608)
);

HB1xp67_ASAP7_75t_L g1609 ( 
.A(n_1517),
.Y(n_1609)
);

AOI21xp33_ASAP7_75t_L g1610 ( 
.A1(n_1597),
.A2(n_1598),
.B(n_1603),
.Y(n_1610)
);

HB1xp67_ASAP7_75t_L g1611 ( 
.A(n_1585),
.Y(n_1611)
);

OR2x2_ASAP7_75t_L g1612 ( 
.A(n_1554),
.B(n_1527),
.Y(n_1612)
);

AOI221xp5_ASAP7_75t_L g1613 ( 
.A1(n_1596),
.A2(n_1477),
.B1(n_1481),
.B2(n_1487),
.C(n_1583),
.Y(n_1613)
);

INVx2_ASAP7_75t_L g1614 ( 
.A(n_1564),
.Y(n_1614)
);

OAI21x1_ASAP7_75t_L g1615 ( 
.A1(n_1504),
.A2(n_1600),
.B(n_1561),
.Y(n_1615)
);

HB1xp67_ASAP7_75t_L g1616 ( 
.A(n_1530),
.Y(n_1616)
);

AND2x2_ASAP7_75t_L g1617 ( 
.A(n_1477),
.B(n_1503),
.Y(n_1617)
);

OAI21x1_ASAP7_75t_L g1618 ( 
.A1(n_1522),
.A2(n_1548),
.B(n_1523),
.Y(n_1618)
);

OAI21xp5_ASAP7_75t_L g1619 ( 
.A1(n_1596),
.A2(n_1529),
.B(n_1511),
.Y(n_1619)
);

AND2x2_ASAP7_75t_L g1620 ( 
.A(n_1511),
.B(n_1524),
.Y(n_1620)
);

INVx1_ASAP7_75t_L g1621 ( 
.A(n_1527),
.Y(n_1621)
);

NAND2xp5_ASAP7_75t_L g1622 ( 
.A(n_1475),
.B(n_1601),
.Y(n_1622)
);

INVx1_ASAP7_75t_L g1623 ( 
.A(n_1534),
.Y(n_1623)
);

OR2x6_ASAP7_75t_L g1624 ( 
.A(n_1534),
.B(n_1542),
.Y(n_1624)
);

INVx2_ASAP7_75t_SL g1625 ( 
.A(n_1533),
.Y(n_1625)
);

AND2x2_ASAP7_75t_L g1626 ( 
.A(n_1554),
.B(n_1542),
.Y(n_1626)
);

INVx1_ASAP7_75t_L g1627 ( 
.A(n_1525),
.Y(n_1627)
);

HB1xp67_ASAP7_75t_L g1628 ( 
.A(n_1507),
.Y(n_1628)
);

AO21x2_ASAP7_75t_L g1629 ( 
.A1(n_1556),
.A2(n_1545),
.B(n_1572),
.Y(n_1629)
);

AO21x2_ASAP7_75t_L g1630 ( 
.A1(n_1556),
.A2(n_1572),
.B(n_1525),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_1459),
.Y(n_1631)
);

OA21x2_ASAP7_75t_L g1632 ( 
.A1(n_1543),
.A2(n_1570),
.B(n_1566),
.Y(n_1632)
);

AND2x2_ASAP7_75t_L g1633 ( 
.A(n_1578),
.B(n_1493),
.Y(n_1633)
);

OR2x6_ASAP7_75t_L g1634 ( 
.A(n_1552),
.B(n_1540),
.Y(n_1634)
);

AND2x2_ASAP7_75t_L g1635 ( 
.A(n_1578),
.B(n_1551),
.Y(n_1635)
);

AND2x2_ASAP7_75t_L g1636 ( 
.A(n_1551),
.B(n_1514),
.Y(n_1636)
);

AND2x2_ASAP7_75t_L g1637 ( 
.A(n_1552),
.B(n_1509),
.Y(n_1637)
);

OR2x2_ASAP7_75t_L g1638 ( 
.A(n_1518),
.B(n_1496),
.Y(n_1638)
);

OA21x2_ASAP7_75t_L g1639 ( 
.A1(n_1543),
.A2(n_1566),
.B(n_1602),
.Y(n_1639)
);

OAI21x1_ASAP7_75t_L g1640 ( 
.A1(n_1458),
.A2(n_1588),
.B(n_1540),
.Y(n_1640)
);

OR2x6_ASAP7_75t_L g1641 ( 
.A(n_1557),
.B(n_1460),
.Y(n_1641)
);

OAI21x1_ASAP7_75t_L g1642 ( 
.A1(n_1458),
.A2(n_1588),
.B(n_1521),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1589),
.Y(n_1643)
);

OR2x2_ASAP7_75t_L g1644 ( 
.A(n_1489),
.B(n_1526),
.Y(n_1644)
);

AND2x4_ASAP7_75t_L g1645 ( 
.A(n_1470),
.B(n_1512),
.Y(n_1645)
);

INVx1_ASAP7_75t_L g1646 ( 
.A(n_1594),
.Y(n_1646)
);

HB1xp67_ASAP7_75t_L g1647 ( 
.A(n_1480),
.Y(n_1647)
);

OR2x2_ASAP7_75t_L g1648 ( 
.A(n_1526),
.B(n_1458),
.Y(n_1648)
);

BUFx8_ASAP7_75t_SL g1649 ( 
.A(n_1466),
.Y(n_1649)
);

BUFx2_ASAP7_75t_L g1650 ( 
.A(n_1588),
.Y(n_1650)
);

AOI21xp5_ASAP7_75t_L g1651 ( 
.A1(n_1508),
.A2(n_1512),
.B(n_1461),
.Y(n_1651)
);

INVxp67_ASAP7_75t_SL g1652 ( 
.A(n_1497),
.Y(n_1652)
);

INVx2_ASAP7_75t_SL g1653 ( 
.A(n_1512),
.Y(n_1653)
);

NAND2x1p5_ASAP7_75t_L g1654 ( 
.A(n_1579),
.B(n_1515),
.Y(n_1654)
);

AND2x4_ASAP7_75t_L g1655 ( 
.A(n_1515),
.B(n_1587),
.Y(n_1655)
);

INVx6_ASAP7_75t_L g1656 ( 
.A(n_1531),
.Y(n_1656)
);

BUFx3_ASAP7_75t_L g1657 ( 
.A(n_1531),
.Y(n_1657)
);

HB1xp67_ASAP7_75t_L g1658 ( 
.A(n_1532),
.Y(n_1658)
);

BUFx3_ASAP7_75t_L g1659 ( 
.A(n_1586),
.Y(n_1659)
);

HB1xp67_ASAP7_75t_L g1660 ( 
.A(n_1593),
.Y(n_1660)
);

AND2x2_ASAP7_75t_L g1661 ( 
.A(n_1491),
.B(n_1463),
.Y(n_1661)
);

NOR2xp33_ASAP7_75t_L g1662 ( 
.A(n_1506),
.B(n_1520),
.Y(n_1662)
);

INVxp67_ASAP7_75t_L g1663 ( 
.A(n_1520),
.Y(n_1663)
);

BUFx2_ASAP7_75t_R g1664 ( 
.A(n_1580),
.Y(n_1664)
);

NAND2xp5_ASAP7_75t_L g1665 ( 
.A(n_1467),
.B(n_1499),
.Y(n_1665)
);

HB1xp67_ASAP7_75t_L g1666 ( 
.A(n_1582),
.Y(n_1666)
);

INVx2_ASAP7_75t_L g1667 ( 
.A(n_1472),
.Y(n_1667)
);

INVx1_ASAP7_75t_L g1668 ( 
.A(n_1473),
.Y(n_1668)
);

INVx2_ASAP7_75t_L g1669 ( 
.A(n_1478),
.Y(n_1669)
);

INVx1_ASAP7_75t_L g1670 ( 
.A(n_1485),
.Y(n_1670)
);

INVx1_ASAP7_75t_L g1671 ( 
.A(n_1486),
.Y(n_1671)
);

CKINVDCx20_ASAP7_75t_R g1672 ( 
.A(n_1466),
.Y(n_1672)
);

HB1xp67_ASAP7_75t_L g1673 ( 
.A(n_1582),
.Y(n_1673)
);

INVx1_ASAP7_75t_L g1674 ( 
.A(n_1488),
.Y(n_1674)
);

INVx2_ASAP7_75t_L g1675 ( 
.A(n_1490),
.Y(n_1675)
);

INVx1_ASAP7_75t_L g1676 ( 
.A(n_1500),
.Y(n_1676)
);

HB1xp67_ASAP7_75t_L g1677 ( 
.A(n_1575),
.Y(n_1677)
);

NAND2xp5_ASAP7_75t_L g1678 ( 
.A(n_1537),
.B(n_1547),
.Y(n_1678)
);

INVx1_ASAP7_75t_L g1679 ( 
.A(n_1528),
.Y(n_1679)
);

BUFx2_ASAP7_75t_L g1680 ( 
.A(n_1569),
.Y(n_1680)
);

AO21x2_ASAP7_75t_L g1681 ( 
.A1(n_1544),
.A2(n_1553),
.B(n_1565),
.Y(n_1681)
);

BUFx2_ASAP7_75t_L g1682 ( 
.A(n_1569),
.Y(n_1682)
);

INVx5_ASAP7_75t_L g1683 ( 
.A(n_1519),
.Y(n_1683)
);

OR2x2_ASAP7_75t_L g1684 ( 
.A(n_1560),
.B(n_1535),
.Y(n_1684)
);

CKINVDCx11_ASAP7_75t_R g1685 ( 
.A(n_1476),
.Y(n_1685)
);

INVx1_ASAP7_75t_L g1686 ( 
.A(n_1573),
.Y(n_1686)
);

AND2x2_ASAP7_75t_L g1687 ( 
.A(n_1469),
.B(n_1505),
.Y(n_1687)
);

NAND2xp5_ASAP7_75t_L g1688 ( 
.A(n_1469),
.B(n_1505),
.Y(n_1688)
);

INVx1_ASAP7_75t_L g1689 ( 
.A(n_1576),
.Y(n_1689)
);

OR2x2_ASAP7_75t_L g1690 ( 
.A(n_1538),
.B(n_1546),
.Y(n_1690)
);

OA21x2_ASAP7_75t_L g1691 ( 
.A1(n_1571),
.A2(n_1505),
.B(n_1471),
.Y(n_1691)
);

INVx1_ASAP7_75t_L g1692 ( 
.A(n_1474),
.Y(n_1692)
);

INVx1_ASAP7_75t_L g1693 ( 
.A(n_1474),
.Y(n_1693)
);

INVx1_ASAP7_75t_L g1694 ( 
.A(n_1584),
.Y(n_1694)
);

AND2x2_ASAP7_75t_L g1695 ( 
.A(n_1469),
.B(n_1471),
.Y(n_1695)
);

INVx1_ASAP7_75t_L g1696 ( 
.A(n_1584),
.Y(n_1696)
);

NAND2xp33_ASAP7_75t_R g1697 ( 
.A(n_1580),
.B(n_1590),
.Y(n_1697)
);

BUFx3_ASAP7_75t_L g1698 ( 
.A(n_1586),
.Y(n_1698)
);

CKINVDCx11_ASAP7_75t_R g1699 ( 
.A(n_1672),
.Y(n_1699)
);

AOI22xp33_ASAP7_75t_L g1700 ( 
.A1(n_1613),
.A2(n_1591),
.B1(n_1636),
.B2(n_1610),
.Y(n_1700)
);

OR2x2_ASAP7_75t_L g1701 ( 
.A(n_1648),
.B(n_1546),
.Y(n_1701)
);

HB1xp67_ASAP7_75t_L g1702 ( 
.A(n_1607),
.Y(n_1702)
);

HB1xp67_ASAP7_75t_L g1703 ( 
.A(n_1609),
.Y(n_1703)
);

AND2x2_ASAP7_75t_L g1704 ( 
.A(n_1626),
.B(n_1471),
.Y(n_1704)
);

NOR2xp33_ASAP7_75t_L g1705 ( 
.A(n_1622),
.B(n_1484),
.Y(n_1705)
);

AND2x2_ASAP7_75t_L g1706 ( 
.A(n_1626),
.B(n_1549),
.Y(n_1706)
);

BUFx2_ASAP7_75t_L g1707 ( 
.A(n_1634),
.Y(n_1707)
);

BUFx6f_ASAP7_75t_SL g1708 ( 
.A(n_1645),
.Y(n_1708)
);

AO22x1_ASAP7_75t_L g1709 ( 
.A1(n_1636),
.A2(n_1581),
.B1(n_1590),
.B2(n_1482),
.Y(n_1709)
);

AND2x2_ASAP7_75t_L g1710 ( 
.A(n_1621),
.B(n_1623),
.Y(n_1710)
);

HB1xp67_ASAP7_75t_L g1711 ( 
.A(n_1611),
.Y(n_1711)
);

HB1xp67_ASAP7_75t_L g1712 ( 
.A(n_1604),
.Y(n_1712)
);

INVx1_ASAP7_75t_L g1713 ( 
.A(n_1631),
.Y(n_1713)
);

AND2x4_ASAP7_75t_SL g1714 ( 
.A(n_1645),
.B(n_1502),
.Y(n_1714)
);

OR2x2_ASAP7_75t_L g1715 ( 
.A(n_1648),
.B(n_1581),
.Y(n_1715)
);

BUFx3_ASAP7_75t_L g1716 ( 
.A(n_1654),
.Y(n_1716)
);

NOR2x1_ASAP7_75t_SL g1717 ( 
.A(n_1630),
.B(n_1581),
.Y(n_1717)
);

NAND2x1_ASAP7_75t_L g1718 ( 
.A(n_1645),
.B(n_1586),
.Y(n_1718)
);

INVx2_ASAP7_75t_SL g1719 ( 
.A(n_1625),
.Y(n_1719)
);

AND2x4_ASAP7_75t_L g1720 ( 
.A(n_1624),
.B(n_1468),
.Y(n_1720)
);

INVxp67_ASAP7_75t_SL g1721 ( 
.A(n_1625),
.Y(n_1721)
);

AOI22xp33_ASAP7_75t_L g1722 ( 
.A1(n_1619),
.A2(n_1549),
.B1(n_1516),
.B2(n_1462),
.Y(n_1722)
);

NAND2xp5_ASAP7_75t_L g1723 ( 
.A(n_1605),
.B(n_1501),
.Y(n_1723)
);

OR2x2_ASAP7_75t_L g1724 ( 
.A(n_1612),
.B(n_1581),
.Y(n_1724)
);

AND2x2_ASAP7_75t_L g1725 ( 
.A(n_1623),
.B(n_1539),
.Y(n_1725)
);

BUFx2_ASAP7_75t_L g1726 ( 
.A(n_1634),
.Y(n_1726)
);

AND2x2_ASAP7_75t_L g1727 ( 
.A(n_1617),
.B(n_1567),
.Y(n_1727)
);

AND2x2_ASAP7_75t_L g1728 ( 
.A(n_1617),
.B(n_1568),
.Y(n_1728)
);

AND2x2_ASAP7_75t_L g1729 ( 
.A(n_1637),
.B(n_1571),
.Y(n_1729)
);

INVx3_ASAP7_75t_L g1730 ( 
.A(n_1634),
.Y(n_1730)
);

OR2x2_ASAP7_75t_L g1731 ( 
.A(n_1612),
.B(n_1502),
.Y(n_1731)
);

INVx2_ASAP7_75t_L g1732 ( 
.A(n_1667),
.Y(n_1732)
);

HB1xp67_ASAP7_75t_L g1733 ( 
.A(n_1628),
.Y(n_1733)
);

OR2x2_ASAP7_75t_L g1734 ( 
.A(n_1634),
.B(n_1464),
.Y(n_1734)
);

INVx3_ASAP7_75t_L g1735 ( 
.A(n_1634),
.Y(n_1735)
);

AND2x2_ASAP7_75t_L g1736 ( 
.A(n_1637),
.B(n_1550),
.Y(n_1736)
);

NAND2xp5_ASAP7_75t_L g1737 ( 
.A(n_1616),
.B(n_1652),
.Y(n_1737)
);

NAND2xp5_ASAP7_75t_L g1738 ( 
.A(n_1662),
.B(n_1550),
.Y(n_1738)
);

INVx2_ASAP7_75t_L g1739 ( 
.A(n_1643),
.Y(n_1739)
);

NAND2xp5_ASAP7_75t_L g1740 ( 
.A(n_1663),
.B(n_1559),
.Y(n_1740)
);

NOR4xp25_ASAP7_75t_SL g1741 ( 
.A(n_1697),
.B(n_1650),
.C(n_1693),
.D(n_1692),
.Y(n_1741)
);

OR2x2_ASAP7_75t_L g1742 ( 
.A(n_1644),
.B(n_1624),
.Y(n_1742)
);

OR2x2_ASAP7_75t_L g1743 ( 
.A(n_1644),
.B(n_1624),
.Y(n_1743)
);

INVx8_ASAP7_75t_L g1744 ( 
.A(n_1683),
.Y(n_1744)
);

AND2x2_ASAP7_75t_L g1745 ( 
.A(n_1606),
.B(n_1646),
.Y(n_1745)
);

OR2x2_ASAP7_75t_L g1746 ( 
.A(n_1639),
.B(n_1559),
.Y(n_1746)
);

OR2x2_ASAP7_75t_L g1747 ( 
.A(n_1639),
.B(n_1574),
.Y(n_1747)
);

INVxp67_ASAP7_75t_SL g1748 ( 
.A(n_1638),
.Y(n_1748)
);

AND2x2_ASAP7_75t_L g1749 ( 
.A(n_1632),
.B(n_1513),
.Y(n_1749)
);

AND2x2_ASAP7_75t_L g1750 ( 
.A(n_1632),
.B(n_1513),
.Y(n_1750)
);

OR2x2_ASAP7_75t_L g1751 ( 
.A(n_1639),
.B(n_1482),
.Y(n_1751)
);

AND2x4_ASAP7_75t_L g1752 ( 
.A(n_1627),
.B(n_1516),
.Y(n_1752)
);

AND2x2_ASAP7_75t_L g1753 ( 
.A(n_1632),
.B(n_1577),
.Y(n_1753)
);

OR2x2_ASAP7_75t_L g1754 ( 
.A(n_1639),
.B(n_1492),
.Y(n_1754)
);

AND2x2_ASAP7_75t_L g1755 ( 
.A(n_1632),
.B(n_1577),
.Y(n_1755)
);

AOI22xp33_ASAP7_75t_L g1756 ( 
.A1(n_1700),
.A2(n_1620),
.B1(n_1635),
.B2(n_1633),
.Y(n_1756)
);

NAND2xp5_ASAP7_75t_L g1757 ( 
.A(n_1702),
.B(n_1638),
.Y(n_1757)
);

OA21x2_ASAP7_75t_L g1758 ( 
.A1(n_1707),
.A2(n_1640),
.B(n_1642),
.Y(n_1758)
);

NAND2xp5_ASAP7_75t_L g1759 ( 
.A(n_1703),
.B(n_1711),
.Y(n_1759)
);

NAND3xp33_ASAP7_75t_L g1760 ( 
.A(n_1709),
.B(n_1635),
.C(n_1620),
.Y(n_1760)
);

NAND2xp5_ASAP7_75t_L g1761 ( 
.A(n_1733),
.B(n_1660),
.Y(n_1761)
);

NAND3xp33_ASAP7_75t_L g1762 ( 
.A(n_1709),
.B(n_1633),
.C(n_1647),
.Y(n_1762)
);

OAI22xp5_ASAP7_75t_L g1763 ( 
.A1(n_1722),
.A2(n_1641),
.B1(n_1684),
.B2(n_1690),
.Y(n_1763)
);

NAND2xp5_ASAP7_75t_SL g1764 ( 
.A(n_1751),
.B(n_1655),
.Y(n_1764)
);

AND2x2_ASAP7_75t_L g1765 ( 
.A(n_1745),
.B(n_1630),
.Y(n_1765)
);

AND2x2_ASAP7_75t_L g1766 ( 
.A(n_1742),
.B(n_1650),
.Y(n_1766)
);

NAND2xp5_ASAP7_75t_SL g1767 ( 
.A(n_1751),
.B(n_1655),
.Y(n_1767)
);

NOR2xp33_ASAP7_75t_L g1768 ( 
.A(n_1705),
.B(n_1690),
.Y(n_1768)
);

NAND2xp5_ASAP7_75t_L g1769 ( 
.A(n_1737),
.B(n_1658),
.Y(n_1769)
);

NAND2xp5_ASAP7_75t_L g1770 ( 
.A(n_1721),
.B(n_1661),
.Y(n_1770)
);

INVx1_ASAP7_75t_L g1771 ( 
.A(n_1713),
.Y(n_1771)
);

AND2x2_ASAP7_75t_L g1772 ( 
.A(n_1742),
.B(n_1661),
.Y(n_1772)
);

AND2x2_ASAP7_75t_L g1773 ( 
.A(n_1743),
.B(n_1629),
.Y(n_1773)
);

OAI21xp33_ASAP7_75t_L g1774 ( 
.A1(n_1723),
.A2(n_1665),
.B(n_1678),
.Y(n_1774)
);

NAND2xp5_ASAP7_75t_L g1775 ( 
.A(n_1748),
.B(n_1666),
.Y(n_1775)
);

NAND2xp5_ASAP7_75t_L g1776 ( 
.A(n_1712),
.B(n_1673),
.Y(n_1776)
);

AND2x2_ASAP7_75t_L g1777 ( 
.A(n_1749),
.B(n_1629),
.Y(n_1777)
);

NAND3xp33_ASAP7_75t_L g1778 ( 
.A(n_1724),
.B(n_1651),
.C(n_1676),
.Y(n_1778)
);

NAND2xp5_ASAP7_75t_SL g1779 ( 
.A(n_1731),
.B(n_1655),
.Y(n_1779)
);

NAND3xp33_ASAP7_75t_L g1780 ( 
.A(n_1724),
.B(n_1676),
.C(n_1677),
.Y(n_1780)
);

NAND2xp5_ASAP7_75t_L g1781 ( 
.A(n_1719),
.B(n_1704),
.Y(n_1781)
);

OAI21xp33_ASAP7_75t_SL g1782 ( 
.A1(n_1754),
.A2(n_1641),
.B(n_1653),
.Y(n_1782)
);

NAND3xp33_ASAP7_75t_L g1783 ( 
.A(n_1754),
.B(n_1679),
.C(n_1674),
.Y(n_1783)
);

AND2x4_ASAP7_75t_L g1784 ( 
.A(n_1716),
.B(n_1645),
.Y(n_1784)
);

NAND2xp5_ASAP7_75t_L g1785 ( 
.A(n_1719),
.B(n_1668),
.Y(n_1785)
);

NAND3xp33_ASAP7_75t_L g1786 ( 
.A(n_1731),
.B(n_1684),
.C(n_1692),
.Y(n_1786)
);

NAND3xp33_ASAP7_75t_L g1787 ( 
.A(n_1701),
.B(n_1693),
.C(n_1694),
.Y(n_1787)
);

NAND2xp5_ASAP7_75t_L g1788 ( 
.A(n_1704),
.B(n_1668),
.Y(n_1788)
);

OAI221xp5_ASAP7_75t_SL g1789 ( 
.A1(n_1715),
.A2(n_1701),
.B1(n_1641),
.B2(n_1746),
.C(n_1747),
.Y(n_1789)
);

NAND4xp25_ASAP7_75t_L g1790 ( 
.A(n_1738),
.B(n_1686),
.C(n_1689),
.D(n_1679),
.Y(n_1790)
);

AND2x2_ASAP7_75t_L g1791 ( 
.A(n_1750),
.B(n_1681),
.Y(n_1791)
);

NAND3xp33_ASAP7_75t_L g1792 ( 
.A(n_1715),
.B(n_1674),
.C(n_1671),
.Y(n_1792)
);

AND2x2_ASAP7_75t_L g1793 ( 
.A(n_1750),
.B(n_1681),
.Y(n_1793)
);

NAND2xp5_ASAP7_75t_L g1794 ( 
.A(n_1706),
.B(n_1669),
.Y(n_1794)
);

NAND3xp33_ASAP7_75t_L g1795 ( 
.A(n_1734),
.B(n_1694),
.C(n_1696),
.Y(n_1795)
);

OAI21xp5_ASAP7_75t_SL g1796 ( 
.A1(n_1714),
.A2(n_1599),
.B(n_1687),
.Y(n_1796)
);

AND2x2_ASAP7_75t_L g1797 ( 
.A(n_1753),
.B(n_1680),
.Y(n_1797)
);

OAI221xp5_ASAP7_75t_SL g1798 ( 
.A1(n_1746),
.A2(n_1641),
.B1(n_1657),
.B2(n_1688),
.C(n_1599),
.Y(n_1798)
);

NAND2xp5_ASAP7_75t_L g1799 ( 
.A(n_1706),
.B(n_1669),
.Y(n_1799)
);

OAI21xp33_ASAP7_75t_L g1800 ( 
.A1(n_1727),
.A2(n_1641),
.B(n_1664),
.Y(n_1800)
);

OA21x2_ASAP7_75t_L g1801 ( 
.A1(n_1726),
.A2(n_1615),
.B(n_1618),
.Y(n_1801)
);

AOI21xp5_ASAP7_75t_L g1802 ( 
.A1(n_1744),
.A2(n_1683),
.B(n_1608),
.Y(n_1802)
);

AND2x2_ASAP7_75t_L g1803 ( 
.A(n_1755),
.B(n_1682),
.Y(n_1803)
);

AOI22xp33_ASAP7_75t_L g1804 ( 
.A1(n_1752),
.A2(n_1691),
.B1(n_1656),
.B2(n_1687),
.Y(n_1804)
);

NAND2xp5_ASAP7_75t_L g1805 ( 
.A(n_1752),
.B(n_1670),
.Y(n_1805)
);

NAND2xp5_ASAP7_75t_SL g1806 ( 
.A(n_1720),
.B(n_1655),
.Y(n_1806)
);

AOI22xp33_ASAP7_75t_L g1807 ( 
.A1(n_1727),
.A2(n_1728),
.B1(n_1691),
.B2(n_1729),
.Y(n_1807)
);

AND2x2_ASAP7_75t_L g1808 ( 
.A(n_1736),
.B(n_1691),
.Y(n_1808)
);

AND2x2_ASAP7_75t_L g1809 ( 
.A(n_1736),
.B(n_1608),
.Y(n_1809)
);

NAND2xp5_ASAP7_75t_L g1810 ( 
.A(n_1710),
.B(n_1675),
.Y(n_1810)
);

AND2x2_ASAP7_75t_L g1811 ( 
.A(n_1726),
.B(n_1608),
.Y(n_1811)
);

AND2x2_ASAP7_75t_L g1812 ( 
.A(n_1739),
.B(n_1614),
.Y(n_1812)
);

AND2x2_ASAP7_75t_L g1813 ( 
.A(n_1739),
.B(n_1614),
.Y(n_1813)
);

NOR2x1_ASAP7_75t_L g1814 ( 
.A(n_1762),
.B(n_1716),
.Y(n_1814)
);

INVx1_ASAP7_75t_L g1815 ( 
.A(n_1771),
.Y(n_1815)
);

INVx2_ASAP7_75t_L g1816 ( 
.A(n_1771),
.Y(n_1816)
);

INVx1_ASAP7_75t_L g1817 ( 
.A(n_1812),
.Y(n_1817)
);

BUFx3_ASAP7_75t_L g1818 ( 
.A(n_1784),
.Y(n_1818)
);

BUFx2_ASAP7_75t_SL g1819 ( 
.A(n_1784),
.Y(n_1819)
);

AND2x2_ASAP7_75t_L g1820 ( 
.A(n_1808),
.B(n_1730),
.Y(n_1820)
);

INVx1_ASAP7_75t_L g1821 ( 
.A(n_1812),
.Y(n_1821)
);

INVx1_ASAP7_75t_L g1822 ( 
.A(n_1813),
.Y(n_1822)
);

AND2x2_ASAP7_75t_L g1823 ( 
.A(n_1777),
.B(n_1735),
.Y(n_1823)
);

INVx2_ASAP7_75t_SL g1824 ( 
.A(n_1784),
.Y(n_1824)
);

AND2x2_ASAP7_75t_L g1825 ( 
.A(n_1777),
.B(n_1735),
.Y(n_1825)
);

INVx2_ASAP7_75t_L g1826 ( 
.A(n_1791),
.Y(n_1826)
);

INVx3_ASAP7_75t_L g1827 ( 
.A(n_1758),
.Y(n_1827)
);

AND2x4_ASAP7_75t_L g1828 ( 
.A(n_1773),
.B(n_1735),
.Y(n_1828)
);

INVx2_ASAP7_75t_L g1829 ( 
.A(n_1793),
.Y(n_1829)
);

INVx1_ASAP7_75t_L g1830 ( 
.A(n_1813),
.Y(n_1830)
);

AOI22xp33_ASAP7_75t_L g1831 ( 
.A1(n_1756),
.A2(n_1728),
.B1(n_1729),
.B2(n_1699),
.Y(n_1831)
);

INVx1_ASAP7_75t_L g1832 ( 
.A(n_1766),
.Y(n_1832)
);

AND2x2_ASAP7_75t_L g1833 ( 
.A(n_1765),
.B(n_1717),
.Y(n_1833)
);

INVx4_ASAP7_75t_L g1834 ( 
.A(n_1801),
.Y(n_1834)
);

AND2x2_ASAP7_75t_SL g1835 ( 
.A(n_1807),
.B(n_1747),
.Y(n_1835)
);

NAND2xp5_ASAP7_75t_L g1836 ( 
.A(n_1809),
.B(n_1732),
.Y(n_1836)
);

AND2x2_ASAP7_75t_L g1837 ( 
.A(n_1811),
.B(n_1717),
.Y(n_1837)
);

INVx1_ASAP7_75t_L g1838 ( 
.A(n_1766),
.Y(n_1838)
);

AOI22xp5_ASAP7_75t_L g1839 ( 
.A1(n_1760),
.A2(n_1725),
.B1(n_1708),
.B2(n_1695),
.Y(n_1839)
);

BUFx3_ASAP7_75t_L g1840 ( 
.A(n_1780),
.Y(n_1840)
);

INVx1_ASAP7_75t_L g1841 ( 
.A(n_1810),
.Y(n_1841)
);

OAI21xp33_ASAP7_75t_L g1842 ( 
.A1(n_1760),
.A2(n_1740),
.B(n_1725),
.Y(n_1842)
);

INVx1_ASAP7_75t_L g1843 ( 
.A(n_1792),
.Y(n_1843)
);

INVx1_ASAP7_75t_L g1844 ( 
.A(n_1792),
.Y(n_1844)
);

AND2x2_ASAP7_75t_L g1845 ( 
.A(n_1772),
.B(n_1797),
.Y(n_1845)
);

INVx1_ASAP7_75t_L g1846 ( 
.A(n_1785),
.Y(n_1846)
);

OR2x2_ASAP7_75t_L g1847 ( 
.A(n_1757),
.B(n_1713),
.Y(n_1847)
);

INVxp67_ASAP7_75t_SL g1848 ( 
.A(n_1778),
.Y(n_1848)
);

INVx2_ASAP7_75t_L g1849 ( 
.A(n_1758),
.Y(n_1849)
);

INVx2_ASAP7_75t_L g1850 ( 
.A(n_1758),
.Y(n_1850)
);

INVx1_ASAP7_75t_L g1851 ( 
.A(n_1794),
.Y(n_1851)
);

INVxp67_ASAP7_75t_SL g1852 ( 
.A(n_1814),
.Y(n_1852)
);

INVx1_ASAP7_75t_SL g1853 ( 
.A(n_1847),
.Y(n_1853)
);

AND2x2_ASAP7_75t_L g1854 ( 
.A(n_1819),
.B(n_1803),
.Y(n_1854)
);

OR2x2_ASAP7_75t_L g1855 ( 
.A(n_1843),
.B(n_1759),
.Y(n_1855)
);

INVx2_ASAP7_75t_L g1856 ( 
.A(n_1816),
.Y(n_1856)
);

AND2x2_ASAP7_75t_L g1857 ( 
.A(n_1819),
.B(n_1803),
.Y(n_1857)
);

NAND2xp5_ASAP7_75t_L g1858 ( 
.A(n_1848),
.B(n_1776),
.Y(n_1858)
);

INVx1_ASAP7_75t_L g1859 ( 
.A(n_1816),
.Y(n_1859)
);

INVx1_ASAP7_75t_L g1860 ( 
.A(n_1816),
.Y(n_1860)
);

INVx1_ASAP7_75t_L g1861 ( 
.A(n_1815),
.Y(n_1861)
);

AND2x2_ASAP7_75t_L g1862 ( 
.A(n_1824),
.B(n_1818),
.Y(n_1862)
);

AND2x2_ASAP7_75t_L g1863 ( 
.A(n_1824),
.B(n_1818),
.Y(n_1863)
);

NAND2xp5_ASAP7_75t_L g1864 ( 
.A(n_1848),
.B(n_1788),
.Y(n_1864)
);

INVx1_ASAP7_75t_SL g1865 ( 
.A(n_1847),
.Y(n_1865)
);

NOR2x1p5_ASAP7_75t_L g1866 ( 
.A(n_1840),
.B(n_1762),
.Y(n_1866)
);

INVx1_ASAP7_75t_L g1867 ( 
.A(n_1815),
.Y(n_1867)
);

INVx1_ASAP7_75t_L g1868 ( 
.A(n_1817),
.Y(n_1868)
);

AND2x2_ASAP7_75t_L g1869 ( 
.A(n_1824),
.B(n_1806),
.Y(n_1869)
);

INVx1_ASAP7_75t_L g1870 ( 
.A(n_1817),
.Y(n_1870)
);

OR2x2_ASAP7_75t_L g1871 ( 
.A(n_1843),
.B(n_1799),
.Y(n_1871)
);

INVx1_ASAP7_75t_L g1872 ( 
.A(n_1821),
.Y(n_1872)
);

NAND2xp5_ASAP7_75t_L g1873 ( 
.A(n_1842),
.B(n_1770),
.Y(n_1873)
);

AND2x2_ASAP7_75t_L g1874 ( 
.A(n_1818),
.B(n_1781),
.Y(n_1874)
);

OR2x2_ASAP7_75t_L g1875 ( 
.A(n_1844),
.B(n_1761),
.Y(n_1875)
);

AND2x2_ASAP7_75t_L g1876 ( 
.A(n_1833),
.B(n_1804),
.Y(n_1876)
);

NAND2xp5_ASAP7_75t_L g1877 ( 
.A(n_1842),
.B(n_1774),
.Y(n_1877)
);

NAND2xp5_ASAP7_75t_L g1878 ( 
.A(n_1846),
.B(n_1851),
.Y(n_1878)
);

NOR3xp33_ASAP7_75t_L g1879 ( 
.A(n_1814),
.B(n_1778),
.C(n_1798),
.Y(n_1879)
);

AND2x2_ASAP7_75t_L g1880 ( 
.A(n_1833),
.B(n_1764),
.Y(n_1880)
);

INVx2_ASAP7_75t_L g1881 ( 
.A(n_1849),
.Y(n_1881)
);

INVx1_ASAP7_75t_L g1882 ( 
.A(n_1821),
.Y(n_1882)
);

INVx1_ASAP7_75t_SL g1883 ( 
.A(n_1847),
.Y(n_1883)
);

NAND3xp33_ASAP7_75t_L g1884 ( 
.A(n_1840),
.B(n_1783),
.C(n_1774),
.Y(n_1884)
);

OAI21xp33_ASAP7_75t_L g1885 ( 
.A1(n_1840),
.A2(n_1800),
.B(n_1790),
.Y(n_1885)
);

HB1xp67_ASAP7_75t_L g1886 ( 
.A(n_1844),
.Y(n_1886)
);

AOI22xp5_ASAP7_75t_L g1887 ( 
.A1(n_1831),
.A2(n_1800),
.B1(n_1763),
.B2(n_1786),
.Y(n_1887)
);

INVx1_ASAP7_75t_L g1888 ( 
.A(n_1822),
.Y(n_1888)
);

OAI21xp33_ASAP7_75t_L g1889 ( 
.A1(n_1831),
.A2(n_1783),
.B(n_1769),
.Y(n_1889)
);

INVx2_ASAP7_75t_L g1890 ( 
.A(n_1849),
.Y(n_1890)
);

NAND2xp5_ASAP7_75t_L g1891 ( 
.A(n_1846),
.B(n_1775),
.Y(n_1891)
);

INVx1_ASAP7_75t_L g1892 ( 
.A(n_1822),
.Y(n_1892)
);

NAND2xp5_ASAP7_75t_L g1893 ( 
.A(n_1851),
.B(n_1805),
.Y(n_1893)
);

AND2x2_ASAP7_75t_L g1894 ( 
.A(n_1833),
.B(n_1767),
.Y(n_1894)
);

INVx1_ASAP7_75t_L g1895 ( 
.A(n_1830),
.Y(n_1895)
);

INVx2_ASAP7_75t_L g1896 ( 
.A(n_1849),
.Y(n_1896)
);

OR2x2_ASAP7_75t_L g1897 ( 
.A(n_1826),
.B(n_1780),
.Y(n_1897)
);

HB1xp67_ASAP7_75t_L g1898 ( 
.A(n_1886),
.Y(n_1898)
);

OAI31xp33_ASAP7_75t_L g1899 ( 
.A1(n_1866),
.A2(n_1789),
.A3(n_1796),
.B(n_1837),
.Y(n_1899)
);

OAI22xp33_ASAP7_75t_L g1900 ( 
.A1(n_1887),
.A2(n_1839),
.B1(n_1718),
.B2(n_1787),
.Y(n_1900)
);

INVx1_ASAP7_75t_L g1901 ( 
.A(n_1861),
.Y(n_1901)
);

INVx2_ASAP7_75t_L g1902 ( 
.A(n_1881),
.Y(n_1902)
);

NAND2xp5_ASAP7_75t_L g1903 ( 
.A(n_1877),
.B(n_1841),
.Y(n_1903)
);

INVx1_ASAP7_75t_L g1904 ( 
.A(n_1861),
.Y(n_1904)
);

NAND2xp5_ASAP7_75t_L g1905 ( 
.A(n_1889),
.B(n_1841),
.Y(n_1905)
);

INVx1_ASAP7_75t_L g1906 ( 
.A(n_1867),
.Y(n_1906)
);

AND2x2_ASAP7_75t_L g1907 ( 
.A(n_1862),
.B(n_1837),
.Y(n_1907)
);

INVx1_ASAP7_75t_L g1908 ( 
.A(n_1867),
.Y(n_1908)
);

AND2x2_ASAP7_75t_L g1909 ( 
.A(n_1862),
.B(n_1837),
.Y(n_1909)
);

NOR2x1_ASAP7_75t_L g1910 ( 
.A(n_1884),
.B(n_1498),
.Y(n_1910)
);

INVx1_ASAP7_75t_SL g1911 ( 
.A(n_1875),
.Y(n_1911)
);

INVx1_ASAP7_75t_L g1912 ( 
.A(n_1868),
.Y(n_1912)
);

INVxp67_ASAP7_75t_L g1913 ( 
.A(n_1875),
.Y(n_1913)
);

OR2x2_ASAP7_75t_L g1914 ( 
.A(n_1853),
.B(n_1826),
.Y(n_1914)
);

AND2x2_ASAP7_75t_L g1915 ( 
.A(n_1863),
.B(n_1823),
.Y(n_1915)
);

INVx1_ASAP7_75t_L g1916 ( 
.A(n_1868),
.Y(n_1916)
);

NAND2xp5_ASAP7_75t_L g1917 ( 
.A(n_1889),
.B(n_1845),
.Y(n_1917)
);

NAND2xp5_ASAP7_75t_L g1918 ( 
.A(n_1858),
.B(n_1845),
.Y(n_1918)
);

OR2x2_ASAP7_75t_L g1919 ( 
.A(n_1865),
.B(n_1883),
.Y(n_1919)
);

INVx1_ASAP7_75t_L g1920 ( 
.A(n_1870),
.Y(n_1920)
);

INVx1_ASAP7_75t_L g1921 ( 
.A(n_1870),
.Y(n_1921)
);

NAND4xp25_ASAP7_75t_L g1922 ( 
.A(n_1884),
.B(n_1839),
.C(n_1768),
.D(n_1795),
.Y(n_1922)
);

INVx1_ASAP7_75t_L g1923 ( 
.A(n_1872),
.Y(n_1923)
);

INVx1_ASAP7_75t_L g1924 ( 
.A(n_1872),
.Y(n_1924)
);

INVxp67_ASAP7_75t_L g1925 ( 
.A(n_1855),
.Y(n_1925)
);

OR2x2_ASAP7_75t_L g1926 ( 
.A(n_1897),
.B(n_1826),
.Y(n_1926)
);

AND2x2_ASAP7_75t_L g1927 ( 
.A(n_1863),
.B(n_1823),
.Y(n_1927)
);

OAI21xp33_ASAP7_75t_L g1928 ( 
.A1(n_1885),
.A2(n_1835),
.B(n_1782),
.Y(n_1928)
);

INVx1_ASAP7_75t_L g1929 ( 
.A(n_1882),
.Y(n_1929)
);

OR2x2_ASAP7_75t_L g1930 ( 
.A(n_1897),
.B(n_1829),
.Y(n_1930)
);

AND2x2_ASAP7_75t_L g1931 ( 
.A(n_1876),
.B(n_1823),
.Y(n_1931)
);

NAND2xp5_ASAP7_75t_L g1932 ( 
.A(n_1864),
.B(n_1845),
.Y(n_1932)
);

AOI22xp5_ASAP7_75t_L g1933 ( 
.A1(n_1879),
.A2(n_1835),
.B1(n_1782),
.B2(n_1779),
.Y(n_1933)
);

AND2x2_ASAP7_75t_L g1934 ( 
.A(n_1876),
.B(n_1825),
.Y(n_1934)
);

NAND2xp5_ASAP7_75t_L g1935 ( 
.A(n_1855),
.B(n_1836),
.Y(n_1935)
);

INVx2_ASAP7_75t_L g1936 ( 
.A(n_1881),
.Y(n_1936)
);

AND2x2_ASAP7_75t_L g1937 ( 
.A(n_1880),
.B(n_1825),
.Y(n_1937)
);

NAND2xp5_ASAP7_75t_L g1938 ( 
.A(n_1873),
.B(n_1836),
.Y(n_1938)
);

OR2x2_ASAP7_75t_L g1939 ( 
.A(n_1871),
.B(n_1829),
.Y(n_1939)
);

AND2x2_ASAP7_75t_L g1940 ( 
.A(n_1880),
.B(n_1825),
.Y(n_1940)
);

OR2x2_ASAP7_75t_L g1941 ( 
.A(n_1871),
.B(n_1829),
.Y(n_1941)
);

INVx1_ASAP7_75t_L g1942 ( 
.A(n_1882),
.Y(n_1942)
);

AND2x4_ASAP7_75t_L g1943 ( 
.A(n_1866),
.B(n_1828),
.Y(n_1943)
);

INVx1_ASAP7_75t_L g1944 ( 
.A(n_1901),
.Y(n_1944)
);

BUFx4f_ASAP7_75t_SL g1945 ( 
.A(n_1911),
.Y(n_1945)
);

INVx1_ASAP7_75t_L g1946 ( 
.A(n_1904),
.Y(n_1946)
);

INVx1_ASAP7_75t_L g1947 ( 
.A(n_1906),
.Y(n_1947)
);

INVx4_ASAP7_75t_L g1948 ( 
.A(n_1943),
.Y(n_1948)
);

INVx1_ASAP7_75t_L g1949 ( 
.A(n_1908),
.Y(n_1949)
);

NAND2xp5_ASAP7_75t_L g1950 ( 
.A(n_1910),
.B(n_1885),
.Y(n_1950)
);

OR2x2_ASAP7_75t_L g1951 ( 
.A(n_1919),
.B(n_1852),
.Y(n_1951)
);

NAND2xp5_ASAP7_75t_L g1952 ( 
.A(n_1903),
.B(n_1894),
.Y(n_1952)
);

HB1xp67_ASAP7_75t_L g1953 ( 
.A(n_1898),
.Y(n_1953)
);

INVx2_ASAP7_75t_L g1954 ( 
.A(n_1915),
.Y(n_1954)
);

NAND2xp5_ASAP7_75t_L g1955 ( 
.A(n_1925),
.B(n_1894),
.Y(n_1955)
);

OAI22xp5_ASAP7_75t_L g1956 ( 
.A1(n_1933),
.A2(n_1887),
.B1(n_1835),
.B2(n_1869),
.Y(n_1956)
);

HB1xp67_ASAP7_75t_L g1957 ( 
.A(n_1913),
.Y(n_1957)
);

AND2x2_ASAP7_75t_L g1958 ( 
.A(n_1943),
.B(n_1907),
.Y(n_1958)
);

AND2x4_ASAP7_75t_L g1959 ( 
.A(n_1943),
.B(n_1869),
.Y(n_1959)
);

INVx2_ASAP7_75t_L g1960 ( 
.A(n_1915),
.Y(n_1960)
);

INVx1_ASAP7_75t_L g1961 ( 
.A(n_1912),
.Y(n_1961)
);

CKINVDCx16_ASAP7_75t_R g1962 ( 
.A(n_1919),
.Y(n_1962)
);

AND2x2_ASAP7_75t_L g1963 ( 
.A(n_1907),
.B(n_1854),
.Y(n_1963)
);

INVx1_ASAP7_75t_L g1964 ( 
.A(n_1916),
.Y(n_1964)
);

INVx2_ASAP7_75t_SL g1965 ( 
.A(n_1909),
.Y(n_1965)
);

OR2x2_ASAP7_75t_L g1966 ( 
.A(n_1935),
.B(n_1878),
.Y(n_1966)
);

NAND2xp5_ASAP7_75t_L g1967 ( 
.A(n_1905),
.B(n_1891),
.Y(n_1967)
);

INVx1_ASAP7_75t_L g1968 ( 
.A(n_1920),
.Y(n_1968)
);

INVx1_ASAP7_75t_L g1969 ( 
.A(n_1921),
.Y(n_1969)
);

INVx2_ASAP7_75t_SL g1970 ( 
.A(n_1909),
.Y(n_1970)
);

NAND2x1_ASAP7_75t_L g1971 ( 
.A(n_1927),
.B(n_1931),
.Y(n_1971)
);

OR2x2_ASAP7_75t_L g1972 ( 
.A(n_1932),
.B(n_1888),
.Y(n_1972)
);

INVx2_ASAP7_75t_L g1973 ( 
.A(n_1927),
.Y(n_1973)
);

OR2x2_ASAP7_75t_L g1974 ( 
.A(n_1918),
.B(n_1888),
.Y(n_1974)
);

NAND2xp5_ASAP7_75t_L g1975 ( 
.A(n_1917),
.B(n_1928),
.Y(n_1975)
);

INVx1_ASAP7_75t_SL g1976 ( 
.A(n_1931),
.Y(n_1976)
);

INVx1_ASAP7_75t_L g1977 ( 
.A(n_1923),
.Y(n_1977)
);

INVx2_ASAP7_75t_L g1978 ( 
.A(n_1937),
.Y(n_1978)
);

INVx1_ASAP7_75t_SL g1979 ( 
.A(n_1934),
.Y(n_1979)
);

HB1xp67_ASAP7_75t_L g1980 ( 
.A(n_1924),
.Y(n_1980)
);

AND2x4_ASAP7_75t_L g1981 ( 
.A(n_1937),
.B(n_1854),
.Y(n_1981)
);

INVx1_ASAP7_75t_L g1982 ( 
.A(n_1929),
.Y(n_1982)
);

AOI32xp33_ASAP7_75t_L g1983 ( 
.A1(n_1956),
.A2(n_1900),
.A3(n_1934),
.B1(n_1940),
.B2(n_1922),
.Y(n_1983)
);

AOI22xp33_ASAP7_75t_L g1984 ( 
.A1(n_1950),
.A2(n_1835),
.B1(n_1899),
.B2(n_1938),
.Y(n_1984)
);

INVx2_ASAP7_75t_L g1985 ( 
.A(n_1971),
.Y(n_1985)
);

INVx2_ASAP7_75t_L g1986 ( 
.A(n_1971),
.Y(n_1986)
);

OR2x2_ASAP7_75t_L g1987 ( 
.A(n_1962),
.B(n_1914),
.Y(n_1987)
);

NOR2x1_ASAP7_75t_L g1988 ( 
.A(n_1948),
.B(n_1498),
.Y(n_1988)
);

OAI22xp33_ASAP7_75t_L g1989 ( 
.A1(n_1945),
.A2(n_1914),
.B1(n_1558),
.B2(n_1834),
.Y(n_1989)
);

AOI21xp33_ASAP7_75t_L g1990 ( 
.A1(n_1975),
.A2(n_1930),
.B(n_1926),
.Y(n_1990)
);

OAI21xp33_ASAP7_75t_L g1991 ( 
.A1(n_1955),
.A2(n_1930),
.B(n_1926),
.Y(n_1991)
);

NAND2xp5_ASAP7_75t_SL g1992 ( 
.A(n_1948),
.B(n_1942),
.Y(n_1992)
);

NAND3xp33_ASAP7_75t_SL g1993 ( 
.A(n_1951),
.B(n_1741),
.C(n_1558),
.Y(n_1993)
);

AOI22xp5_ASAP7_75t_L g1994 ( 
.A1(n_1948),
.A2(n_1940),
.B1(n_1874),
.B2(n_1857),
.Y(n_1994)
);

NOR3xp33_ASAP7_75t_SL g1995 ( 
.A(n_1967),
.B(n_1893),
.C(n_1802),
.Y(n_1995)
);

NAND2xp5_ASAP7_75t_SL g1996 ( 
.A(n_1951),
.B(n_1939),
.Y(n_1996)
);

OAI21xp33_ASAP7_75t_L g1997 ( 
.A1(n_1957),
.A2(n_1941),
.B(n_1939),
.Y(n_1997)
);

AND2x2_ASAP7_75t_L g1998 ( 
.A(n_1958),
.B(n_1874),
.Y(n_1998)
);

INVx2_ASAP7_75t_L g1999 ( 
.A(n_1981),
.Y(n_1999)
);

OR2x2_ASAP7_75t_L g2000 ( 
.A(n_1976),
.B(n_1941),
.Y(n_2000)
);

INVx2_ASAP7_75t_SL g2001 ( 
.A(n_1959),
.Y(n_2001)
);

AND2x2_ASAP7_75t_L g2002 ( 
.A(n_1958),
.B(n_1857),
.Y(n_2002)
);

NAND4xp25_ASAP7_75t_SL g2003 ( 
.A(n_1979),
.B(n_1838),
.C(n_1832),
.D(n_1820),
.Y(n_2003)
);

INVxp33_ASAP7_75t_L g2004 ( 
.A(n_1953),
.Y(n_2004)
);

AND2x2_ASAP7_75t_L g2005 ( 
.A(n_1959),
.B(n_1828),
.Y(n_2005)
);

OAI21xp33_ASAP7_75t_L g2006 ( 
.A1(n_1952),
.A2(n_1936),
.B(n_1902),
.Y(n_2006)
);

INVx3_ASAP7_75t_L g2007 ( 
.A(n_1959),
.Y(n_2007)
);

INVx1_ASAP7_75t_L g2008 ( 
.A(n_1980),
.Y(n_2008)
);

INVx1_ASAP7_75t_L g2009 ( 
.A(n_1944),
.Y(n_2009)
);

INVxp33_ASAP7_75t_L g2010 ( 
.A(n_1978),
.Y(n_2010)
);

AOI222xp33_ASAP7_75t_L g2011 ( 
.A1(n_1978),
.A2(n_1834),
.B1(n_1827),
.B2(n_1555),
.C1(n_1850),
.C2(n_1685),
.Y(n_2011)
);

INVx2_ASAP7_75t_L g2012 ( 
.A(n_2007),
.Y(n_2012)
);

NAND2xp5_ASAP7_75t_L g2013 ( 
.A(n_2004),
.B(n_1965),
.Y(n_2013)
);

OR2x2_ASAP7_75t_L g2014 ( 
.A(n_1987),
.B(n_1966),
.Y(n_2014)
);

NAND3xp33_ASAP7_75t_L g2015 ( 
.A(n_1984),
.B(n_1961),
.C(n_1949),
.Y(n_2015)
);

NAND2xp5_ASAP7_75t_L g2016 ( 
.A(n_2004),
.B(n_1965),
.Y(n_2016)
);

INVx1_ASAP7_75t_L g2017 ( 
.A(n_1996),
.Y(n_2017)
);

NAND2xp5_ASAP7_75t_L g2018 ( 
.A(n_2001),
.B(n_1970),
.Y(n_2018)
);

HB1xp67_ASAP7_75t_L g2019 ( 
.A(n_1999),
.Y(n_2019)
);

HB1xp67_ASAP7_75t_L g2020 ( 
.A(n_1999),
.Y(n_2020)
);

INVx1_ASAP7_75t_L g2021 ( 
.A(n_2009),
.Y(n_2021)
);

NAND2xp5_ASAP7_75t_L g2022 ( 
.A(n_2008),
.B(n_2007),
.Y(n_2022)
);

INVx1_ASAP7_75t_L g2023 ( 
.A(n_2010),
.Y(n_2023)
);

INVx1_ASAP7_75t_SL g2024 ( 
.A(n_1988),
.Y(n_2024)
);

INVx1_ASAP7_75t_L g2025 ( 
.A(n_1996),
.Y(n_2025)
);

NAND2xp5_ASAP7_75t_L g2026 ( 
.A(n_1984),
.B(n_1970),
.Y(n_2026)
);

AOI22xp33_ASAP7_75t_SL g2027 ( 
.A1(n_1983),
.A2(n_1981),
.B1(n_1954),
.B2(n_1960),
.Y(n_2027)
);

INVx1_ASAP7_75t_L g2028 ( 
.A(n_2010),
.Y(n_2028)
);

INVx1_ASAP7_75t_L g2029 ( 
.A(n_2000),
.Y(n_2029)
);

AND2x2_ASAP7_75t_L g2030 ( 
.A(n_2002),
.B(n_1981),
.Y(n_2030)
);

INVx1_ASAP7_75t_L g2031 ( 
.A(n_1992),
.Y(n_2031)
);

INVx1_ASAP7_75t_L g2032 ( 
.A(n_1992),
.Y(n_2032)
);

HB1xp67_ASAP7_75t_L g2033 ( 
.A(n_1985),
.Y(n_2033)
);

INVx1_ASAP7_75t_L g2034 ( 
.A(n_1985),
.Y(n_2034)
);

AOI211xp5_ASAP7_75t_L g2035 ( 
.A1(n_2024),
.A2(n_1989),
.B(n_1993),
.C(n_1990),
.Y(n_2035)
);

NAND2xp5_ASAP7_75t_L g2036 ( 
.A(n_2012),
.B(n_1997),
.Y(n_2036)
);

OAI22xp5_ASAP7_75t_L g2037 ( 
.A1(n_2027),
.A2(n_1995),
.B1(n_1994),
.B2(n_1989),
.Y(n_2037)
);

NOR2x1_ASAP7_75t_L g2038 ( 
.A(n_2012),
.B(n_1986),
.Y(n_2038)
);

AOI22xp5_ASAP7_75t_L g2039 ( 
.A1(n_2030),
.A2(n_2026),
.B1(n_2015),
.B2(n_2029),
.Y(n_2039)
);

NAND2xp5_ASAP7_75t_L g2040 ( 
.A(n_2023),
.B(n_2028),
.Y(n_2040)
);

NAND3xp33_ASAP7_75t_L g2041 ( 
.A(n_2017),
.B(n_1986),
.C(n_1991),
.Y(n_2041)
);

OAI211xp5_ASAP7_75t_L g2042 ( 
.A1(n_2017),
.A2(n_2011),
.B(n_2006),
.C(n_1555),
.Y(n_2042)
);

AOI21xp5_ASAP7_75t_SL g2043 ( 
.A1(n_2032),
.A2(n_2003),
.B(n_1649),
.Y(n_2043)
);

AOI32xp33_ASAP7_75t_L g2044 ( 
.A1(n_2025),
.A2(n_1998),
.A3(n_1954),
.B1(n_1960),
.B2(n_1973),
.Y(n_2044)
);

NOR2x1_ASAP7_75t_L g2045 ( 
.A(n_2032),
.B(n_2034),
.Y(n_2045)
);

AOI221xp5_ASAP7_75t_L g2046 ( 
.A1(n_2025),
.A2(n_1946),
.B1(n_1968),
.B2(n_1977),
.C(n_1944),
.Y(n_2046)
);

AOI21xp5_ASAP7_75t_L g2047 ( 
.A1(n_2014),
.A2(n_1969),
.B(n_1964),
.Y(n_2047)
);

NAND2xp5_ASAP7_75t_L g2048 ( 
.A(n_2031),
.B(n_1973),
.Y(n_2048)
);

NOR2x1_ASAP7_75t_L g2049 ( 
.A(n_2045),
.B(n_2034),
.Y(n_2049)
);

NAND2xp5_ASAP7_75t_L g2050 ( 
.A(n_2039),
.B(n_2019),
.Y(n_2050)
);

NOR2x1_ASAP7_75t_L g2051 ( 
.A(n_2038),
.B(n_2013),
.Y(n_2051)
);

INVx1_ASAP7_75t_L g2052 ( 
.A(n_2040),
.Y(n_2052)
);

NAND2xp5_ASAP7_75t_SL g2053 ( 
.A(n_2035),
.B(n_2014),
.Y(n_2053)
);

NAND3xp33_ASAP7_75t_L g2054 ( 
.A(n_2041),
.B(n_2022),
.C(n_2020),
.Y(n_2054)
);

XNOR2xp5_ASAP7_75t_L g2055 ( 
.A(n_2042),
.B(n_2016),
.Y(n_2055)
);

INVx1_ASAP7_75t_L g2056 ( 
.A(n_2048),
.Y(n_2056)
);

NOR3xp33_ASAP7_75t_L g2057 ( 
.A(n_2036),
.B(n_2018),
.C(n_2021),
.Y(n_2057)
);

INVxp67_ASAP7_75t_L g2058 ( 
.A(n_2047),
.Y(n_2058)
);

AOI22xp5_ASAP7_75t_L g2059 ( 
.A1(n_2037),
.A2(n_2030),
.B1(n_2033),
.B2(n_2005),
.Y(n_2059)
);

AOI21xp5_ASAP7_75t_L g2060 ( 
.A1(n_2043),
.A2(n_1982),
.B(n_1947),
.Y(n_2060)
);

NOR3x1_ASAP7_75t_L g2061 ( 
.A(n_2044),
.B(n_1947),
.C(n_1946),
.Y(n_2061)
);

NAND3xp33_ASAP7_75t_L g2062 ( 
.A(n_2053),
.B(n_2046),
.C(n_1977),
.Y(n_2062)
);

NAND5xp2_ASAP7_75t_L g2063 ( 
.A(n_2059),
.B(n_1968),
.C(n_1963),
.D(n_1479),
.E(n_1476),
.Y(n_2063)
);

NAND2xp5_ASAP7_75t_SL g2064 ( 
.A(n_2051),
.B(n_1966),
.Y(n_2064)
);

NAND4xp25_ASAP7_75t_SL g2065 ( 
.A(n_2050),
.B(n_1963),
.C(n_1972),
.D(n_1974),
.Y(n_2065)
);

NOR4xp25_ASAP7_75t_L g2066 ( 
.A(n_2054),
.B(n_1974),
.C(n_1972),
.D(n_1936),
.Y(n_2066)
);

NOR4xp25_ASAP7_75t_L g2067 ( 
.A(n_2058),
.B(n_1902),
.C(n_1896),
.D(n_1890),
.Y(n_2067)
);

NAND2xp5_ASAP7_75t_L g2068 ( 
.A(n_2057),
.B(n_1892),
.Y(n_2068)
);

AOI211xp5_ASAP7_75t_L g2069 ( 
.A1(n_2055),
.A2(n_1657),
.B(n_1479),
.C(n_1595),
.Y(n_2069)
);

INVx2_ASAP7_75t_L g2070 ( 
.A(n_2064),
.Y(n_2070)
);

AO22x2_ASAP7_75t_L g2071 ( 
.A1(n_2062),
.A2(n_2052),
.B1(n_2056),
.B2(n_2049),
.Y(n_2071)
);

INVx1_ASAP7_75t_L g2072 ( 
.A(n_2068),
.Y(n_2072)
);

AOI31xp33_ASAP7_75t_L g2073 ( 
.A1(n_2069),
.A2(n_2060),
.A3(n_2061),
.B(n_1595),
.Y(n_2073)
);

INVx1_ASAP7_75t_L g2074 ( 
.A(n_2065),
.Y(n_2074)
);

INVxp67_ASAP7_75t_L g2075 ( 
.A(n_2063),
.Y(n_2075)
);

AOI22xp5_ASAP7_75t_L g2076 ( 
.A1(n_2066),
.A2(n_1536),
.B1(n_1656),
.B2(n_1896),
.Y(n_2076)
);

XNOR2xp5_ASAP7_75t_L g2077 ( 
.A(n_2074),
.B(n_2070),
.Y(n_2077)
);

NOR3xp33_ASAP7_75t_SL g2078 ( 
.A(n_2072),
.B(n_2067),
.C(n_1536),
.Y(n_2078)
);

NAND4xp75_ASAP7_75t_L g2079 ( 
.A(n_2076),
.B(n_1890),
.C(n_1895),
.D(n_1892),
.Y(n_2079)
);

NOR2xp33_ASAP7_75t_R g2080 ( 
.A(n_2075),
.B(n_1657),
.Y(n_2080)
);

AND2x2_ASAP7_75t_L g2081 ( 
.A(n_2071),
.B(n_2073),
.Y(n_2081)
);

NOR2x1_ASAP7_75t_L g2082 ( 
.A(n_2071),
.B(n_1856),
.Y(n_2082)
);

CKINVDCx16_ASAP7_75t_R g2083 ( 
.A(n_2080),
.Y(n_2083)
);

INVx2_ASAP7_75t_L g2084 ( 
.A(n_2082),
.Y(n_2084)
);

INVx2_ASAP7_75t_L g2085 ( 
.A(n_2079),
.Y(n_2085)
);

INVx1_ASAP7_75t_L g2086 ( 
.A(n_2077),
.Y(n_2086)
);

INVx2_ASAP7_75t_L g2087 ( 
.A(n_2084),
.Y(n_2087)
);

XNOR2xp5_ASAP7_75t_L g2088 ( 
.A(n_2087),
.B(n_2086),
.Y(n_2088)
);

INVx1_ASAP7_75t_L g2089 ( 
.A(n_2088),
.Y(n_2089)
);

OAI22x1_ASAP7_75t_L g2090 ( 
.A1(n_2088),
.A2(n_2085),
.B1(n_2081),
.B2(n_2083),
.Y(n_2090)
);

OAI21xp5_ASAP7_75t_L g2091 ( 
.A1(n_2089),
.A2(n_2078),
.B(n_2083),
.Y(n_2091)
);

OAI22xp5_ASAP7_75t_L g2092 ( 
.A1(n_2090),
.A2(n_1656),
.B1(n_1895),
.B2(n_1856),
.Y(n_2092)
);

INVx2_ASAP7_75t_L g2093 ( 
.A(n_2092),
.Y(n_2093)
);

OA21x2_ASAP7_75t_L g2094 ( 
.A1(n_2091),
.A2(n_1856),
.B(n_1859),
.Y(n_2094)
);

AOI21xp5_ASAP7_75t_SL g2095 ( 
.A1(n_2093),
.A2(n_1698),
.B(n_1659),
.Y(n_2095)
);

AOI22xp33_ASAP7_75t_L g2096 ( 
.A1(n_2095),
.A2(n_2094),
.B1(n_1656),
.B2(n_1827),
.Y(n_2096)
);

OAI221xp5_ASAP7_75t_L g2097 ( 
.A1(n_2096),
.A2(n_2094),
.B1(n_1562),
.B2(n_1860),
.C(n_1859),
.Y(n_2097)
);

AOI211xp5_ASAP7_75t_L g2098 ( 
.A1(n_2097),
.A2(n_1659),
.B(n_1698),
.C(n_1860),
.Y(n_2098)
);


endmodule