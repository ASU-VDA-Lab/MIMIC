module fake_jpeg_20527_n_280 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_280);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_280;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_272;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_270;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_265;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_140;
wire n_258;
wire n_96;

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_11),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_2),
.B(n_10),
.Y(n_19)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_12),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_SL g24 ( 
.A(n_6),
.B(n_15),
.Y(n_24)
);

INVx6_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_5),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

BUFx2_ASAP7_75t_R g29 ( 
.A(n_6),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_22),
.Y(n_33)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_28),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_34),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_28),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_35),
.Y(n_53)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_21),
.Y(n_36)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_37),
.Y(n_41)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_28),
.Y(n_39)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g40 ( 
.A(n_24),
.B(n_0),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_40),
.B(n_24),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_SL g42 ( 
.A1(n_36),
.A2(n_29),
.B1(n_25),
.B2(n_20),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_42),
.A2(n_48),
.B1(n_21),
.B2(n_27),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g43 ( 
.A(n_40),
.B(n_24),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_43),
.B(n_49),
.Y(n_67)
);

INVx11_ASAP7_75t_L g45 ( 
.A(n_33),
.Y(n_45)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_45),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_38),
.A2(n_25),
.B1(n_32),
.B2(n_20),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_46),
.A2(n_21),
.B1(n_30),
.B2(n_17),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_33),
.A2(n_25),
.B1(n_29),
.B2(n_20),
.Y(n_48)
);

BUFx5_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_52),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_36),
.B(n_19),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_54),
.B(n_17),
.Y(n_72)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

BUFx2_ASAP7_75t_L g69 ( 
.A(n_55),
.Y(n_69)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_35),
.Y(n_56)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_56),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_37),
.B(n_27),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_58),
.B(n_47),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_59),
.B(n_60),
.Y(n_100)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_51),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_58),
.B(n_38),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_61),
.B(n_63),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_47),
.A2(n_38),
.B1(n_34),
.B2(n_25),
.Y(n_62)
);

OAI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_62),
.A2(n_74),
.B1(n_57),
.B2(n_44),
.Y(n_97)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_51),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_56),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_64),
.B(n_66),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_42),
.B(n_54),
.C(n_46),
.Y(n_65)
);

XNOR2xp5_ASAP7_75t_L g99 ( 
.A(n_65),
.B(n_75),
.Y(n_99)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_51),
.Y(n_66)
);

AOI21xp5_ASAP7_75t_L g70 ( 
.A1(n_42),
.A2(n_34),
.B(n_29),
.Y(n_70)
);

OAI21xp5_ASAP7_75t_SL g93 ( 
.A1(n_70),
.A2(n_76),
.B(n_22),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_45),
.A2(n_17),
.B1(n_23),
.B2(n_32),
.Y(n_71)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_71),
.Y(n_109)
);

CKINVDCx14_ASAP7_75t_R g107 ( 
.A(n_72),
.Y(n_107)
);

OAI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_41),
.A2(n_32),
.B1(n_30),
.B2(n_23),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_46),
.B(n_16),
.C(n_26),
.Y(n_75)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_49),
.B(n_39),
.Y(n_76)
);

CKINVDCx16_ASAP7_75t_R g88 ( 
.A(n_77),
.Y(n_88)
);

CKINVDCx16_ASAP7_75t_R g78 ( 
.A(n_48),
.Y(n_78)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_78),
.Y(n_87)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_51),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_79),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_L g81 ( 
.A1(n_41),
.A2(n_30),
.B1(n_27),
.B2(n_23),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_L g108 ( 
.A1(n_81),
.A2(n_82),
.B1(n_52),
.B2(n_26),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_45),
.A2(n_22),
.B1(n_26),
.B2(n_16),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_83),
.A2(n_55),
.B1(n_50),
.B2(n_57),
.Y(n_96)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_44),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_84),
.Y(n_95)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_57),
.Y(n_85)
);

HB1xp67_ASAP7_75t_L g86 ( 
.A(n_85),
.Y(n_86)
);

AOI32xp33_ASAP7_75t_L g89 ( 
.A1(n_78),
.A2(n_65),
.A3(n_70),
.B1(n_77),
.B2(n_67),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_89),
.B(n_35),
.Y(n_118)
);

A2O1A1Ixp33_ASAP7_75t_L g90 ( 
.A1(n_59),
.A2(n_43),
.B(n_19),
.C(n_50),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_90),
.B(n_67),
.Y(n_115)
);

OA22x2_ASAP7_75t_L g92 ( 
.A1(n_75),
.A2(n_41),
.B1(n_55),
.B2(n_50),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g124 ( 
.A(n_92),
.B(n_105),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_L g117 ( 
.A1(n_93),
.A2(n_98),
.B(n_61),
.Y(n_117)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_76),
.B(n_62),
.Y(n_94)
);

INVx1_ASAP7_75t_SL g128 ( 
.A(n_94),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_96),
.A2(n_68),
.B1(n_80),
.B2(n_69),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_97),
.A2(n_80),
.B1(n_39),
.B2(n_26),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_L g98 ( 
.A1(n_76),
.A2(n_18),
.B(n_31),
.Y(n_98)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_73),
.Y(n_102)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_102),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_73),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_103),
.B(n_104),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_82),
.Y(n_104)
);

OA22x2_ASAP7_75t_L g105 ( 
.A1(n_64),
.A2(n_44),
.B1(n_52),
.B2(n_35),
.Y(n_105)
);

OR2x2_ASAP7_75t_L g113 ( 
.A(n_108),
.B(n_63),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_72),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_110),
.B(n_53),
.Y(n_138)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_69),
.Y(n_111)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_111),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_113),
.A2(n_134),
.B1(n_104),
.B2(n_109),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_86),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_114),
.B(n_122),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_115),
.B(n_123),
.Y(n_139)
);

CKINVDCx9p33_ASAP7_75t_R g116 ( 
.A(n_107),
.Y(n_116)
);

CKINVDCx14_ASAP7_75t_R g147 ( 
.A(n_116),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_SL g167 ( 
.A(n_117),
.B(n_118),
.C(n_119),
.Y(n_167)
);

AND2x4_ASAP7_75t_L g119 ( 
.A(n_93),
.B(n_85),
.Y(n_119)
);

BUFx2_ASAP7_75t_L g120 ( 
.A(n_91),
.Y(n_120)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_120),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_99),
.B(n_53),
.C(n_80),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_121),
.B(n_92),
.C(n_101),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_110),
.B(n_84),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_99),
.B(n_79),
.Y(n_123)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_95),
.Y(n_125)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_125),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_88),
.A2(n_66),
.B1(n_60),
.B2(n_68),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_126),
.A2(n_137),
.B1(n_94),
.B2(n_87),
.Y(n_152)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_129),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_100),
.B(n_69),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_130),
.B(n_138),
.Y(n_148)
);

NAND2xp33_ASAP7_75t_SL g131 ( 
.A(n_94),
.B(n_105),
.Y(n_131)
);

XOR2x2_ASAP7_75t_L g159 ( 
.A(n_131),
.B(n_105),
.Y(n_159)
);

AND2x2_ASAP7_75t_L g133 ( 
.A(n_92),
.B(n_39),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_L g141 ( 
.A(n_133),
.B(n_135),
.Y(n_141)
);

OAI21x1_ASAP7_75t_L g135 ( 
.A1(n_90),
.A2(n_31),
.B(n_18),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_106),
.Y(n_136)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_136),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_88),
.A2(n_53),
.B1(n_31),
.B2(n_18),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_114),
.B(n_107),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_140),
.B(n_146),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_142),
.A2(n_150),
.B1(n_133),
.B2(n_124),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_120),
.Y(n_143)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_143),
.Y(n_180)
);

XOR2xp5_ASAP7_75t_L g145 ( 
.A(n_123),
.B(n_98),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_SL g186 ( 
.A(n_145),
.B(n_7),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_136),
.B(n_103),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_113),
.A2(n_89),
.B1(n_87),
.B2(n_101),
.Y(n_150)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_137),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_151),
.B(n_154),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_152),
.A2(n_160),
.B1(n_0),
.B2(n_1),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_153),
.B(n_150),
.C(n_141),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_130),
.B(n_100),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_115),
.B(n_90),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_156),
.B(n_157),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_112),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_125),
.B(n_106),
.Y(n_158)
);

CKINVDCx14_ASAP7_75t_R g189 ( 
.A(n_158),
.Y(n_189)
);

INVx1_ASAP7_75t_SL g185 ( 
.A(n_159),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_124),
.A2(n_133),
.B1(n_127),
.B2(n_126),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_120),
.Y(n_161)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_161),
.Y(n_193)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_132),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_162),
.B(n_163),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_112),
.Y(n_163)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_132),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_165),
.B(n_53),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_145),
.B(n_121),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_168),
.B(n_170),
.Y(n_195)
);

OA21x2_ASAP7_75t_L g169 ( 
.A1(n_159),
.A2(n_124),
.B(n_131),
.Y(n_169)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_169),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g170 ( 
.A(n_153),
.B(n_117),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_171),
.A2(n_176),
.B1(n_177),
.B2(n_178),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_173),
.B(n_175),
.C(n_186),
.Y(n_199)
);

OAI22xp33_ASAP7_75t_L g174 ( 
.A1(n_151),
.A2(n_144),
.B1(n_142),
.B2(n_160),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_174),
.A2(n_181),
.B1(n_188),
.B2(n_147),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_139),
.B(n_119),
.C(n_128),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_144),
.A2(n_119),
.B1(n_128),
.B2(n_113),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_141),
.A2(n_119),
.B1(n_92),
.B2(n_135),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_156),
.A2(n_167),
.B1(n_149),
.B2(n_139),
.Y(n_178)
);

A2O1A1O1Ixp25_ASAP7_75t_L g179 ( 
.A1(n_167),
.A2(n_119),
.B(n_92),
.C(n_105),
.D(n_129),
.Y(n_179)
);

XNOR2x1_ASAP7_75t_L g205 ( 
.A(n_179),
.B(n_155),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_152),
.A2(n_134),
.B1(n_102),
.B2(n_105),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_148),
.A2(n_111),
.B1(n_95),
.B2(n_91),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_182),
.B(n_166),
.Y(n_200)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_183),
.Y(n_202)
);

OA21x2_ASAP7_75t_L g184 ( 
.A1(n_148),
.A2(n_53),
.B(n_1),
.Y(n_184)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_184),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_165),
.B(n_15),
.C(n_7),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_SL g203 ( 
.A(n_192),
.B(n_9),
.Y(n_203)
);

CKINVDCx16_ASAP7_75t_R g194 ( 
.A(n_187),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_194),
.B(n_200),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_L g196 ( 
.A1(n_172),
.A2(n_164),
.B(n_161),
.Y(n_196)
);

CKINVDCx14_ASAP7_75t_R g225 ( 
.A(n_196),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_197),
.A2(n_214),
.B1(n_184),
.B2(n_171),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_190),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_201),
.B(n_207),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_203),
.B(n_205),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_185),
.A2(n_155),
.B1(n_166),
.B2(n_143),
.Y(n_204)
);

HB1xp67_ASAP7_75t_L g218 ( 
.A(n_204),
.Y(n_218)
);

INVxp33_ASAP7_75t_L g206 ( 
.A(n_191),
.Y(n_206)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_206),
.Y(n_222)
);

INVxp67_ASAP7_75t_L g207 ( 
.A(n_174),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_SL g209 ( 
.A(n_189),
.B(n_7),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_209),
.B(n_212),
.Y(n_221)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_182),
.Y(n_211)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_211),
.Y(n_223)
);

CKINVDCx14_ASAP7_75t_R g212 ( 
.A(n_192),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_193),
.Y(n_213)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_213),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_184),
.B(n_0),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_207),
.A2(n_181),
.B1(n_185),
.B2(n_179),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_216),
.A2(n_231),
.B1(n_198),
.B2(n_200),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_195),
.B(n_173),
.C(n_170),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_217),
.B(n_229),
.C(n_204),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_SL g220 ( 
.A(n_195),
.B(n_168),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_220),
.B(n_226),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_224),
.B(n_2),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_SL g226 ( 
.A(n_199),
.B(n_178),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_199),
.B(n_208),
.C(n_175),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_205),
.B(n_186),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_230),
.B(n_203),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_211),
.A2(n_169),
.B1(n_177),
.B2(n_176),
.Y(n_231)
);

AOI322xp5_ASAP7_75t_L g232 ( 
.A1(n_222),
.A2(n_210),
.A3(n_196),
.B1(n_202),
.B2(n_198),
.C1(n_197),
.C2(n_213),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_232),
.B(n_236),
.Y(n_255)
);

OAI21xp5_ASAP7_75t_SL g234 ( 
.A1(n_218),
.A2(n_201),
.B(n_202),
.Y(n_234)
);

OAI21xp5_ASAP7_75t_SL g245 ( 
.A1(n_234),
.A2(n_221),
.B(n_227),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_235),
.B(n_237),
.C(n_238),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_229),
.B(n_210),
.C(n_169),
.Y(n_237)
);

OAI21xp5_ASAP7_75t_L g239 ( 
.A1(n_225),
.A2(n_214),
.B(n_209),
.Y(n_239)
);

AOI21xp5_ASAP7_75t_L g249 ( 
.A1(n_239),
.A2(n_243),
.B(n_241),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_215),
.B(n_180),
.Y(n_240)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_240),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_216),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_L g246 ( 
.A1(n_241),
.A2(n_223),
.B1(n_231),
.B2(n_228),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_242),
.A2(n_228),
.B1(n_230),
.B2(n_4),
.Y(n_253)
);

OAI21xp5_ASAP7_75t_L g243 ( 
.A1(n_219),
.A2(n_8),
.B(n_14),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_226),
.B(n_8),
.C(n_14),
.Y(n_244)
);

INVxp67_ASAP7_75t_L g247 ( 
.A(n_244),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_245),
.B(n_250),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_246),
.A2(n_251),
.B1(n_253),
.B2(n_247),
.Y(n_257)
);

OR2x2_ASAP7_75t_L g259 ( 
.A(n_249),
.B(n_236),
.Y(n_259)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_243),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_L g251 ( 
.A1(n_239),
.A2(n_237),
.B1(n_244),
.B2(n_235),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_253),
.B(n_10),
.Y(n_263)
);

NAND3xp33_ASAP7_75t_L g254 ( 
.A(n_238),
.B(n_220),
.C(n_217),
.Y(n_254)
);

NOR2xp67_ASAP7_75t_SL g258 ( 
.A(n_254),
.B(n_233),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_257),
.B(n_260),
.Y(n_265)
);

OAI21xp5_ASAP7_75t_L g270 ( 
.A1(n_258),
.A2(n_252),
.B(n_264),
.Y(n_270)
);

AOI21xp5_ASAP7_75t_L g269 ( 
.A1(n_259),
.A2(n_261),
.B(n_264),
.Y(n_269)
);

AO21x1_ASAP7_75t_L g260 ( 
.A1(n_255),
.A2(n_233),
.B(n_8),
.Y(n_260)
);

OAI21xp5_ASAP7_75t_SL g261 ( 
.A1(n_247),
.A2(n_15),
.B(n_12),
.Y(n_261)
);

INVx6_ASAP7_75t_L g262 ( 
.A(n_248),
.Y(n_262)
);

INVx1_ASAP7_75t_SL g267 ( 
.A(n_262),
.Y(n_267)
);

NOR3xp33_ASAP7_75t_L g268 ( 
.A(n_263),
.B(n_2),
.C(n_3),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_249),
.B(n_11),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_256),
.B(n_252),
.C(n_11),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_266),
.B(n_4),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_268),
.Y(n_274)
);

NOR4xp25_ASAP7_75t_L g272 ( 
.A(n_270),
.B(n_3),
.C(n_4),
.D(n_5),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_265),
.A2(n_259),
.B1(n_260),
.B2(n_5),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_271),
.B(n_273),
.Y(n_276)
);

A2O1A1Ixp33_ASAP7_75t_L g275 ( 
.A1(n_272),
.A2(n_269),
.B(n_5),
.C(n_6),
.Y(n_275)
);

OA21x2_ASAP7_75t_SL g277 ( 
.A1(n_275),
.A2(n_274),
.B(n_6),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_277),
.B(n_276),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_278),
.B(n_267),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_279),
.B(n_4),
.Y(n_280)
);


endmodule