module fake_jpeg_10861_n_380 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_380);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_380;

wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_13),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

BUFx4f_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

INVx11_ASAP7_75t_SL g18 ( 
.A(n_14),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_1),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_9),
.Y(n_27)
);

BUFx10_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_10),
.B(n_3),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_10),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_5),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_9),
.Y(n_35)
);

BUFx16f_ASAP7_75t_L g36 ( 
.A(n_6),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_14),
.B(n_13),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_4),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_3),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_1),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_6),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_12),
.Y(n_42)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_26),
.Y(n_43)
);

INVx5_ASAP7_75t_L g122 ( 
.A(n_43),
.Y(n_122)
);

BUFx16f_ASAP7_75t_L g44 ( 
.A(n_28),
.Y(n_44)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_44),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_16),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_45),
.Y(n_92)
);

INVx1_ASAP7_75t_SL g46 ( 
.A(n_28),
.Y(n_46)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_46),
.B(n_66),
.Y(n_110)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_22),
.Y(n_47)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_47),
.Y(n_85)
);

INVx13_ASAP7_75t_L g48 ( 
.A(n_28),
.Y(n_48)
);

BUFx2_ASAP7_75t_L g94 ( 
.A(n_48),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_16),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_49),
.Y(n_100)
);

BUFx10_ASAP7_75t_L g50 ( 
.A(n_28),
.Y(n_50)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_50),
.Y(n_98)
);

INVx5_ASAP7_75t_L g51 ( 
.A(n_23),
.Y(n_51)
);

INVx4_ASAP7_75t_L g116 ( 
.A(n_51),
.Y(n_116)
);

INVx11_ASAP7_75t_L g52 ( 
.A(n_28),
.Y(n_52)
);

INVx11_ASAP7_75t_L g86 ( 
.A(n_52),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_16),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_53),
.Y(n_101)
);

INVx11_ASAP7_75t_L g54 ( 
.A(n_28),
.Y(n_54)
);

INVx4_ASAP7_75t_L g125 ( 
.A(n_54),
.Y(n_125)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_26),
.Y(n_55)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_55),
.Y(n_121)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_26),
.Y(n_56)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_56),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_16),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_57),
.Y(n_112)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_31),
.Y(n_58)
);

INVx6_ASAP7_75t_L g95 ( 
.A(n_58),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_30),
.Y(n_59)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_59),
.Y(n_129)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_31),
.Y(n_60)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_60),
.Y(n_119)
);

BUFx12_ASAP7_75t_L g61 ( 
.A(n_18),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_61),
.Y(n_108)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_31),
.Y(n_62)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_62),
.Y(n_114)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_19),
.Y(n_63)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_63),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_37),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_64),
.B(n_69),
.Y(n_87)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_23),
.Y(n_65)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_65),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_30),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_30),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_67),
.B(n_68),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_37),
.B(n_14),
.Y(n_68)
);

INVx13_ASAP7_75t_L g69 ( 
.A(n_18),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_29),
.B(n_0),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_70),
.B(n_0),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_29),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_71),
.B(n_72),
.Y(n_104)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_40),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_19),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_73),
.B(n_74),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_17),
.Y(n_74)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_22),
.Y(n_75)
);

AO22x1_ASAP7_75t_L g120 ( 
.A1(n_75),
.A2(n_76),
.B1(n_79),
.B2(n_80),
.Y(n_120)
);

INVx2_ASAP7_75t_SL g76 ( 
.A(n_20),
.Y(n_76)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_23),
.Y(n_77)
);

OR2x2_ASAP7_75t_L g106 ( 
.A(n_77),
.B(n_78),
.Y(n_106)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_32),
.Y(n_78)
);

INVx2_ASAP7_75t_SL g79 ( 
.A(n_20),
.Y(n_79)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_35),
.Y(n_80)
);

BUFx5_ASAP7_75t_L g81 ( 
.A(n_36),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_81),
.B(n_1),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_15),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_82),
.B(n_13),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_70),
.A2(n_42),
.B1(n_15),
.B2(n_35),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_83),
.A2(n_89),
.B1(n_115),
.B2(n_120),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_47),
.A2(n_20),
.B1(n_24),
.B2(n_32),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_84),
.A2(n_88),
.B1(n_90),
.B2(n_117),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_L g88 ( 
.A1(n_59),
.A2(n_24),
.B1(n_41),
.B2(n_39),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_66),
.A2(n_42),
.B1(n_24),
.B2(n_21),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_L g90 ( 
.A1(n_67),
.A2(n_41),
.B1(n_21),
.B2(n_39),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_93),
.B(n_11),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_75),
.B(n_25),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_96),
.B(n_103),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_46),
.A2(n_32),
.B1(n_40),
.B2(n_79),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_97),
.A2(n_99),
.B1(n_102),
.B2(n_109),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_76),
.A2(n_40),
.B1(n_25),
.B2(n_33),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_65),
.A2(n_38),
.B1(n_34),
.B2(n_33),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_80),
.B(n_38),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_77),
.B(n_34),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_107),
.B(n_126),
.Y(n_158)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_78),
.A2(n_27),
.B1(n_36),
.B2(n_17),
.Y(n_109)
);

OAI22xp33_ASAP7_75t_L g115 ( 
.A1(n_45),
.A2(n_17),
.B1(n_27),
.B2(n_36),
.Y(n_115)
);

OA22x2_ASAP7_75t_L g117 ( 
.A1(n_50),
.A2(n_17),
.B1(n_36),
.B2(n_2),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_43),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g157 ( 
.A(n_118),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_124),
.B(n_87),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_49),
.B(n_0),
.Y(n_126)
);

INVxp33_ASAP7_75t_L g146 ( 
.A(n_128),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_96),
.B(n_105),
.C(n_103),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_130),
.B(n_135),
.C(n_144),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_SL g208 ( 
.A(n_131),
.B(n_141),
.Y(n_208)
);

BUFx4f_ASAP7_75t_L g132 ( 
.A(n_86),
.Y(n_132)
);

INVx3_ASAP7_75t_L g195 ( 
.A(n_132),
.Y(n_195)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_94),
.Y(n_133)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_133),
.Y(n_183)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_94),
.Y(n_134)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_134),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_107),
.B(n_50),
.C(n_54),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_L g136 ( 
.A1(n_115),
.A2(n_53),
.B1(n_57),
.B2(n_74),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_136),
.A2(n_137),
.B1(n_171),
.B2(n_125),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_L g137 ( 
.A1(n_120),
.A2(n_52),
.B1(n_50),
.B2(n_72),
.Y(n_137)
);

INVx13_ASAP7_75t_L g138 ( 
.A(n_108),
.Y(n_138)
);

INVx11_ASAP7_75t_L g178 ( 
.A(n_138),
.Y(n_178)
);

OAI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_84),
.A2(n_62),
.B1(n_56),
.B2(n_48),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_139),
.A2(n_125),
.B1(n_86),
.B2(n_116),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_93),
.B(n_51),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_140),
.B(n_143),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_104),
.B(n_44),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_111),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_142),
.B(n_162),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_113),
.B(n_12),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_85),
.B(n_126),
.C(n_106),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_85),
.B(n_44),
.C(n_55),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_145),
.B(n_163),
.C(n_154),
.Y(n_212)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_120),
.Y(n_147)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_147),
.Y(n_187)
);

BUFx3_ASAP7_75t_L g148 ( 
.A(n_91),
.Y(n_148)
);

BUFx12f_ASAP7_75t_L g194 ( 
.A(n_148),
.Y(n_194)
);

AND2x2_ASAP7_75t_L g206 ( 
.A(n_149),
.B(n_161),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_106),
.B(n_12),
.Y(n_150)
);

INVxp67_ASAP7_75t_L g191 ( 
.A(n_150),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_114),
.B(n_81),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_151),
.B(n_156),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_110),
.B(n_2),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_154),
.B(n_160),
.Y(n_179)
);

INVx5_ASAP7_75t_L g155 ( 
.A(n_91),
.Y(n_155)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_155),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_114),
.B(n_55),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_117),
.A2(n_60),
.B1(n_58),
.B2(n_69),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_159),
.A2(n_122),
.B1(n_123),
.B2(n_129),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_117),
.B(n_2),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_SL g161 ( 
.A1(n_117),
.A2(n_61),
.B(n_5),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g162 ( 
.A(n_127),
.Y(n_162)
);

OR2x2_ASAP7_75t_L g163 ( 
.A(n_98),
.B(n_61),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_163),
.B(n_167),
.Y(n_198)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_110),
.Y(n_164)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_164),
.Y(n_199)
);

INVx3_ASAP7_75t_L g165 ( 
.A(n_95),
.Y(n_165)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_165),
.Y(n_209)
);

INVx5_ASAP7_75t_L g166 ( 
.A(n_121),
.Y(n_166)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_166),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_SL g167 ( 
.A(n_121),
.B(n_4),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_168),
.B(n_173),
.Y(n_186)
);

OR2x2_ASAP7_75t_L g169 ( 
.A(n_98),
.B(n_11),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_169),
.B(n_172),
.Y(n_192)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_110),
.Y(n_170)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_170),
.Y(n_214)
);

AOI22xp33_ASAP7_75t_L g171 ( 
.A1(n_129),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_119),
.B(n_7),
.Y(n_172)
);

INVx4_ASAP7_75t_L g173 ( 
.A(n_95),
.Y(n_173)
);

INVxp67_ASAP7_75t_L g174 ( 
.A(n_119),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_174),
.B(n_8),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_176),
.A2(n_181),
.B1(n_189),
.B2(n_203),
.Y(n_243)
);

AOI22xp33_ASAP7_75t_SL g177 ( 
.A1(n_157),
.A2(n_123),
.B1(n_122),
.B2(n_116),
.Y(n_177)
);

CKINVDCx14_ASAP7_75t_R g249 ( 
.A(n_177),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_180),
.A2(n_190),
.B1(n_197),
.B2(n_155),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_153),
.A2(n_92),
.B1(n_100),
.B2(n_101),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_147),
.A2(n_92),
.B1(n_100),
.B2(n_101),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_172),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_193),
.B(n_202),
.Y(n_235)
);

AOI22xp33_ASAP7_75t_SL g197 ( 
.A1(n_157),
.A2(n_112),
.B1(n_10),
.B2(n_11),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_158),
.B(n_112),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_200),
.B(n_210),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_138),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_153),
.A2(n_160),
.B1(n_159),
.B2(n_152),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_204),
.B(n_134),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_146),
.B(n_8),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_SL g242 ( 
.A(n_205),
.B(n_185),
.Y(n_242)
);

AOI21xp5_ASAP7_75t_L g207 ( 
.A1(n_175),
.A2(n_8),
.B(n_163),
.Y(n_207)
);

AOI21xp5_ASAP7_75t_SL g241 ( 
.A1(n_207),
.A2(n_198),
.B(n_206),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_158),
.B(n_152),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_212),
.B(n_132),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_138),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_213),
.B(n_148),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_164),
.A2(n_170),
.B1(n_144),
.B2(n_130),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_215),
.B(n_216),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_140),
.B(n_135),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_178),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_217),
.B(n_221),
.Y(n_260)
);

A2O1A1O1Ixp25_ASAP7_75t_L g218 ( 
.A1(n_216),
.A2(n_143),
.B(n_145),
.C(n_142),
.D(n_161),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_SL g267 ( 
.A1(n_218),
.A2(n_219),
.B(n_230),
.Y(n_267)
);

O2A1O1Ixp33_ASAP7_75t_SL g219 ( 
.A1(n_206),
.A2(n_169),
.B(n_175),
.C(n_149),
.Y(n_219)
);

BUFx6f_ASAP7_75t_L g220 ( 
.A(n_194),
.Y(n_220)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_220),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_178),
.Y(n_221)
);

OAI32xp33_ASAP7_75t_L g222 ( 
.A1(n_187),
.A2(n_167),
.A3(n_173),
.B1(n_169),
.B2(n_133),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_222),
.B(n_237),
.Y(n_266)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_183),
.Y(n_224)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_224),
.Y(n_268)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_183),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_226),
.B(n_227),
.Y(n_252)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_184),
.Y(n_227)
);

CKINVDCx14_ASAP7_75t_R g273 ( 
.A(n_228),
.Y(n_273)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_184),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_229),
.B(n_232),
.Y(n_253)
);

A2O1A1O1Ixp25_ASAP7_75t_L g230 ( 
.A1(n_201),
.A2(n_174),
.B(n_162),
.C(n_165),
.D(n_166),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_202),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_SL g257 ( 
.A(n_231),
.B(n_238),
.Y(n_257)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_209),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_209),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_233),
.B(n_236),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_L g256 ( 
.A1(n_234),
.A2(n_207),
.B1(n_176),
.B2(n_189),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_185),
.Y(n_237)
);

BUFx2_ASAP7_75t_R g238 ( 
.A(n_213),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_210),
.B(n_132),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_SL g270 ( 
.A(n_239),
.B(n_211),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_240),
.B(n_248),
.C(n_214),
.Y(n_259)
);

OAI21xp5_ASAP7_75t_SL g269 ( 
.A1(n_241),
.A2(n_188),
.B(n_199),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_242),
.A2(n_247),
.B1(n_194),
.B2(n_217),
.Y(n_277)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_190),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_244),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_193),
.B(n_200),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_245),
.B(n_250),
.Y(n_272)
);

INVx2_ASAP7_75t_SL g246 ( 
.A(n_195),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_246),
.Y(n_278)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_211),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_201),
.B(n_215),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_187),
.B(n_192),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_243),
.A2(n_206),
.B1(n_203),
.B2(n_180),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_L g300 ( 
.A1(n_254),
.A2(n_271),
.B1(n_276),
.B2(n_277),
.Y(n_300)
);

AOI322xp5_ASAP7_75t_L g255 ( 
.A1(n_237),
.A2(n_188),
.A3(n_198),
.B1(n_191),
.B2(n_179),
.C1(n_186),
.C2(n_208),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_SL g284 ( 
.A(n_255),
.B(n_229),
.C(n_224),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_256),
.A2(n_279),
.B1(n_280),
.B2(n_246),
.Y(n_298)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_248),
.B(n_212),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_258),
.B(n_259),
.Y(n_289)
);

AOI21xp5_ASAP7_75t_L g261 ( 
.A1(n_235),
.A2(n_181),
.B(n_182),
.Y(n_261)
);

INVxp67_ASAP7_75t_L g290 ( 
.A(n_261),
.Y(n_290)
);

OAI21xp5_ASAP7_75t_L g263 ( 
.A1(n_241),
.A2(n_179),
.B(n_192),
.Y(n_263)
);

INVxp67_ASAP7_75t_L g294 ( 
.A(n_263),
.Y(n_294)
);

OAI21xp5_ASAP7_75t_L g265 ( 
.A1(n_225),
.A2(n_199),
.B(n_214),
.Y(n_265)
);

INVxp67_ASAP7_75t_L g304 ( 
.A(n_265),
.Y(n_304)
);

OAI21xp33_ASAP7_75t_L g283 ( 
.A1(n_269),
.A2(n_274),
.B(n_275),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_SL g286 ( 
.A(n_270),
.B(n_226),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_243),
.A2(n_208),
.B1(n_191),
.B2(n_196),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_SL g274 ( 
.A(n_225),
.B(n_240),
.Y(n_274)
);

OAI21xp5_ASAP7_75t_L g275 ( 
.A1(n_250),
.A2(n_196),
.B(n_195),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_244),
.A2(n_219),
.B1(n_245),
.B2(n_223),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_219),
.A2(n_194),
.B1(n_223),
.B2(n_234),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_L g280 ( 
.A1(n_218),
.A2(n_249),
.B1(n_222),
.B2(n_230),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_253),
.Y(n_281)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_281),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_253),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_SL g316 ( 
.A(n_282),
.B(n_299),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_L g306 ( 
.A(n_284),
.B(n_286),
.Y(n_306)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_260),
.Y(n_285)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_285),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_252),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_287),
.B(n_288),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_254),
.A2(n_276),
.B1(n_266),
.B2(n_271),
.Y(n_288)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_252),
.Y(n_291)
);

HB1xp67_ASAP7_75t_L g322 ( 
.A(n_291),
.Y(n_322)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_268),
.Y(n_292)
);

BUFx2_ASAP7_75t_L g309 ( 
.A(n_292),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_272),
.B(n_227),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_293),
.Y(n_314)
);

AOI22xp33_ASAP7_75t_SL g295 ( 
.A1(n_279),
.A2(n_247),
.B1(n_220),
.B2(n_232),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_L g307 ( 
.A1(n_295),
.A2(n_297),
.B1(n_298),
.B2(n_301),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_272),
.B(n_233),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_296),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_266),
.A2(n_238),
.B1(n_246),
.B2(n_194),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_273),
.B(n_257),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_251),
.A2(n_263),
.B1(n_265),
.B2(n_261),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_SL g302 ( 
.A(n_257),
.B(n_269),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_L g318 ( 
.A1(n_302),
.A2(n_303),
.B1(n_278),
.B2(n_256),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_SL g303 ( 
.A(n_264),
.B(n_259),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_289),
.B(n_258),
.C(n_274),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_305),
.B(n_315),
.C(n_317),
.Y(n_331)
);

OAI21xp5_ASAP7_75t_L g311 ( 
.A1(n_304),
.A2(n_267),
.B(n_277),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_311),
.B(n_297),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_SL g312 ( 
.A1(n_298),
.A2(n_251),
.B1(n_267),
.B2(n_280),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_312),
.B(n_320),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_289),
.B(n_270),
.C(n_275),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_296),
.B(n_264),
.C(n_268),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_SL g338 ( 
.A(n_318),
.B(n_292),
.Y(n_338)
);

OAI22xp5_ASAP7_75t_SL g320 ( 
.A1(n_304),
.A2(n_262),
.B1(n_278),
.B2(n_294),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_293),
.B(n_262),
.C(n_294),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_321),
.B(n_290),
.C(n_291),
.Y(n_336)
);

XNOR2xp5_ASAP7_75t_L g323 ( 
.A(n_283),
.B(n_301),
.Y(n_323)
);

XOR2xp5_ASAP7_75t_L g329 ( 
.A(n_323),
.B(n_300),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_314),
.B(n_287),
.Y(n_325)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_325),
.Y(n_342)
);

XNOR2xp5_ASAP7_75t_L g340 ( 
.A(n_326),
.B(n_336),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_316),
.B(n_285),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_327),
.B(n_328),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_319),
.B(n_288),
.Y(n_328)
);

XOR2xp5_ASAP7_75t_L g347 ( 
.A(n_329),
.B(n_332),
.Y(n_347)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_319),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_330),
.B(n_333),
.Y(n_345)
);

XOR2xp5_ASAP7_75t_L g332 ( 
.A(n_305),
.B(n_290),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_317),
.B(n_281),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_322),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_334),
.B(n_335),
.Y(n_346)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_310),
.Y(n_335)
);

XOR2xp5_ASAP7_75t_L g337 ( 
.A(n_315),
.B(n_284),
.Y(n_337)
);

XOR2xp5_ASAP7_75t_L g348 ( 
.A(n_337),
.B(n_306),
.Y(n_348)
);

OAI22xp5_ASAP7_75t_L g350 ( 
.A1(n_338),
.A2(n_310),
.B1(n_313),
.B2(n_308),
.Y(n_350)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_321),
.B(n_323),
.C(n_306),
.Y(n_339)
);

HB1xp67_ASAP7_75t_L g349 ( 
.A(n_339),
.Y(n_349)
);

XNOR2xp5_ASAP7_75t_L g343 ( 
.A(n_331),
.B(n_311),
.Y(n_343)
);

XNOR2xp5_ASAP7_75t_L g357 ( 
.A(n_343),
.B(n_344),
.Y(n_357)
);

XNOR2xp5_ASAP7_75t_L g344 ( 
.A(n_331),
.B(n_312),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_348),
.B(n_350),
.Y(n_356)
);

HB1xp67_ASAP7_75t_L g351 ( 
.A(n_336),
.Y(n_351)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_351),
.Y(n_354)
);

OAI22xp5_ASAP7_75t_L g352 ( 
.A1(n_341),
.A2(n_324),
.B1(n_308),
.B2(n_325),
.Y(n_352)
);

XNOR2xp5_ASAP7_75t_L g363 ( 
.A(n_352),
.B(n_353),
.Y(n_363)
);

OAI22xp5_ASAP7_75t_L g353 ( 
.A1(n_342),
.A2(n_324),
.B1(n_345),
.B2(n_346),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_340),
.B(n_314),
.Y(n_355)
);

AOI21x1_ASAP7_75t_SL g365 ( 
.A1(n_355),
.A2(n_358),
.B(n_347),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_340),
.Y(n_358)
);

HB1xp67_ASAP7_75t_L g359 ( 
.A(n_349),
.Y(n_359)
);

AND2x2_ASAP7_75t_L g361 ( 
.A(n_359),
.B(n_360),
.Y(n_361)
);

OAI22xp5_ASAP7_75t_SL g360 ( 
.A1(n_344),
.A2(n_307),
.B1(n_339),
.B2(n_329),
.Y(n_360)
);

OAI22xp5_ASAP7_75t_SL g362 ( 
.A1(n_356),
.A2(n_309),
.B1(n_337),
.B2(n_320),
.Y(n_362)
);

INVxp67_ASAP7_75t_L g371 ( 
.A(n_362),
.Y(n_371)
);

OAI22xp5_ASAP7_75t_L g364 ( 
.A1(n_354),
.A2(n_309),
.B1(n_343),
.B2(n_348),
.Y(n_364)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_364),
.Y(n_370)
);

AOI21xp33_ASAP7_75t_L g368 ( 
.A1(n_365),
.A2(n_357),
.B(n_360),
.Y(n_368)
);

AOI21xp5_ASAP7_75t_L g366 ( 
.A1(n_358),
.A2(n_332),
.B(n_347),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_SL g369 ( 
.A(n_366),
.B(n_361),
.Y(n_369)
);

XOR2x1_ASAP7_75t_L g367 ( 
.A(n_355),
.B(n_357),
.Y(n_367)
);

NOR2xp67_ASAP7_75t_SL g372 ( 
.A(n_367),
.B(n_361),
.Y(n_372)
);

OAI21xp5_ASAP7_75t_L g374 ( 
.A1(n_368),
.A2(n_372),
.B(n_367),
.Y(n_374)
);

INVxp67_ASAP7_75t_L g375 ( 
.A(n_369),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_SL g373 ( 
.A(n_371),
.B(n_363),
.Y(n_373)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_373),
.Y(n_377)
);

HB1xp67_ASAP7_75t_L g376 ( 
.A(n_374),
.Y(n_376)
);

INVxp67_ASAP7_75t_L g378 ( 
.A(n_376),
.Y(n_378)
);

MAJIxp5_ASAP7_75t_L g379 ( 
.A(n_378),
.B(n_375),
.C(n_377),
.Y(n_379)
);

XOR2xp5_ASAP7_75t_L g380 ( 
.A(n_379),
.B(n_370),
.Y(n_380)
);


endmodule