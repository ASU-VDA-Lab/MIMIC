module fake_aes_11090_n_14 (n_1, n_2, n_4, n_3, n_5, n_0, n_14);
input n_1;
input n_2;
input n_4;
input n_3;
input n_5;
input n_0;
output n_14;
wire n_11;
wire n_13;
wire n_12;
wire n_6;
wire n_9;
wire n_7;
wire n_10;
wire n_8;
NOR2xp33_ASAP7_75t_L g6 ( .A(n_4), .B(n_1), .Y(n_6) );
INVx2_ASAP7_75t_L g7 ( .A(n_2), .Y(n_7) );
INVx2_ASAP7_75t_L g8 ( .A(n_5), .Y(n_8) );
AND2x2_ASAP7_75t_L g9 ( .A(n_7), .B(n_0), .Y(n_9) );
INVx2_ASAP7_75t_L g10 ( .A(n_8), .Y(n_10) );
A2O1A1Ixp33_ASAP7_75t_L g11 ( .A1(n_10), .A2(n_6), .B(n_1), .C(n_2), .Y(n_11) );
NAND2xp5_ASAP7_75t_SL g12 ( .A(n_11), .B(n_9), .Y(n_12) );
INVx1_ASAP7_75t_L g13 ( .A(n_12), .Y(n_13) );
AOI22xp33_ASAP7_75t_L g14 ( .A1(n_13), .A2(n_0), .B1(n_3), .B2(n_12), .Y(n_14) );
endmodule