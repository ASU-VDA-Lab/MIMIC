module fake_jpeg_1711_n_19 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_19);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_19;

wire n_13;
wire n_14;
wire n_18;
wire n_16;
wire n_17;
wire n_15;

AOI22xp33_ASAP7_75t_SL g13 ( 
.A1(n_9),
.A2(n_1),
.B1(n_0),
.B2(n_10),
.Y(n_13)
);

AOI22xp33_ASAP7_75t_SL g14 ( 
.A1(n_5),
.A2(n_7),
.B1(n_2),
.B2(n_1),
.Y(n_14)
);

INVx2_ASAP7_75t_L g15 ( 
.A(n_12),
.Y(n_15)
);

OAI22xp5_ASAP7_75t_SL g16 ( 
.A1(n_15),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_16)
);

AOI22xp5_ASAP7_75t_L g18 ( 
.A1(n_16),
.A2(n_17),
.B1(n_13),
.B2(n_14),
.Y(n_18)
);

OAI22xp5_ASAP7_75t_L g17 ( 
.A1(n_15),
.A2(n_4),
.B1(n_6),
.B2(n_8),
.Y(n_17)
);

XOR2xp5_ASAP7_75t_L g19 ( 
.A(n_18),
.B(n_11),
.Y(n_19)
);


endmodule