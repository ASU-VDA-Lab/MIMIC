module fake_jpeg_22911_n_250 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_250);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_250;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_212;
wire n_131;
wire n_56;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

BUFx2_ASAP7_75t_L g15 ( 
.A(n_4),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_0),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_3),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

BUFx10_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_18),
.Y(n_32)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_32),
.Y(n_52)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_18),
.Y(n_33)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_16),
.B(n_8),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_34),
.B(n_38),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g35 ( 
.A1(n_25),
.A2(n_26),
.B1(n_28),
.B2(n_18),
.Y(n_35)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_35),
.A2(n_25),
.B1(n_28),
.B2(n_26),
.Y(n_59)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_23),
.Y(n_36)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_36),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_18),
.Y(n_37)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_37),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_16),
.B(n_8),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_30),
.Y(n_39)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_39),
.Y(n_60)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_40),
.B(n_15),
.Y(n_48)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_23),
.Y(n_41)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_41),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_23),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_42),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_34),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_46),
.B(n_47),
.Y(n_76)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_41),
.Y(n_47)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_48),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_38),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_49),
.B(n_55),
.Y(n_77)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_41),
.Y(n_50)
);

INVx8_ASAP7_75t_L g81 ( 
.A(n_50),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g53 ( 
.A(n_32),
.B(n_9),
.Y(n_53)
);

A2O1A1Ixp33_ASAP7_75t_L g71 ( 
.A1(n_53),
.A2(n_63),
.B(n_31),
.C(n_19),
.Y(n_71)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_35),
.Y(n_54)
);

INVx5_ASAP7_75t_L g78 ( 
.A(n_54),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_33),
.B(n_20),
.Y(n_55)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_32),
.Y(n_56)
);

HB1xp67_ASAP7_75t_L g73 ( 
.A(n_56),
.Y(n_73)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_58),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_59),
.A2(n_22),
.B1(n_29),
.B2(n_27),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_40),
.B(n_20),
.Y(n_62)
);

INVxp67_ASAP7_75t_L g70 ( 
.A(n_62),
.Y(n_70)
);

INVx2_ASAP7_75t_R g63 ( 
.A(n_37),
.Y(n_63)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_42),
.Y(n_64)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_64),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_54),
.A2(n_36),
.B1(n_40),
.B2(n_39),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_65),
.A2(n_79),
.B1(n_17),
.B2(n_24),
.Y(n_99)
);

AND2x2_ASAP7_75t_SL g67 ( 
.A(n_63),
.B(n_36),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_67),
.B(n_49),
.C(n_51),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_46),
.B(n_31),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_69),
.B(n_58),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_71),
.B(n_51),
.Y(n_93)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_60),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_72),
.B(n_74),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g74 ( 
.A(n_56),
.Y(n_74)
);

AO22x1_ASAP7_75t_L g75 ( 
.A1(n_59),
.A2(n_42),
.B1(n_31),
.B2(n_15),
.Y(n_75)
);

AO22x1_ASAP7_75t_L g98 ( 
.A1(n_75),
.A2(n_82),
.B1(n_31),
.B2(n_45),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_L g79 ( 
.A1(n_53),
.A2(n_22),
.B1(n_29),
.B2(n_27),
.Y(n_79)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_57),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_80),
.B(n_64),
.Y(n_92)
);

AO22x1_ASAP7_75t_L g82 ( 
.A1(n_61),
.A2(n_31),
.B1(n_15),
.B2(n_0),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_L g104 ( 
.A1(n_84),
.A2(n_17),
.B1(n_21),
.B2(n_24),
.Y(n_104)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_73),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_85),
.B(n_87),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_82),
.Y(n_87)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_76),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_88),
.B(n_89),
.Y(n_125)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_82),
.Y(n_89)
);

FAx1_ASAP7_75t_L g90 ( 
.A(n_69),
.B(n_53),
.CI(n_61),
.CON(n_90),
.SN(n_90)
);

A2O1A1O1Ixp25_ASAP7_75t_L g111 ( 
.A1(n_90),
.A2(n_106),
.B(n_67),
.C(n_75),
.D(n_78),
.Y(n_111)
);

AOI21xp5_ASAP7_75t_L g113 ( 
.A1(n_91),
.A2(n_83),
.B(n_70),
.Y(n_113)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_92),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_93),
.B(n_105),
.Y(n_109)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_65),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_94),
.B(n_96),
.Y(n_112)
);

BUFx8_ASAP7_75t_L g95 ( 
.A(n_67),
.Y(n_95)
);

INVx1_ASAP7_75t_SL g120 ( 
.A(n_95),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_77),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_84),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_97),
.B(n_99),
.Y(n_118)
);

O2A1O1Ixp33_ASAP7_75t_L g126 ( 
.A1(n_98),
.A2(n_74),
.B(n_44),
.C(n_47),
.Y(n_126)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_77),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_100),
.B(n_101),
.Y(n_121)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_71),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_75),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_102),
.B(n_103),
.Y(n_110)
);

CKINVDCx16_ASAP7_75t_R g107 ( 
.A(n_104),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g105 ( 
.A(n_78),
.B(n_83),
.Y(n_105)
);

AOI32xp33_ASAP7_75t_L g106 ( 
.A1(n_70),
.A2(n_60),
.A3(n_43),
.B1(n_52),
.B2(n_57),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_86),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_108),
.B(n_115),
.Y(n_133)
);

AO21x1_ASAP7_75t_L g147 ( 
.A1(n_111),
.A2(n_21),
.B(n_52),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_L g145 ( 
.A1(n_113),
.A2(n_95),
.B(n_90),
.Y(n_145)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_105),
.Y(n_115)
);

AOI21xp5_ASAP7_75t_L g117 ( 
.A1(n_87),
.A2(n_80),
.B(n_44),
.Y(n_117)
);

AOI21xp5_ASAP7_75t_L g129 ( 
.A1(n_117),
.A2(n_89),
.B(n_98),
.Y(n_129)
);

CKINVDCx14_ASAP7_75t_R g119 ( 
.A(n_93),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_119),
.B(n_122),
.Y(n_141)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_99),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_96),
.B(n_81),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_123),
.B(n_100),
.Y(n_130)
);

INVx13_ASAP7_75t_L g124 ( 
.A(n_85),
.Y(n_124)
);

INVx6_ASAP7_75t_L g134 ( 
.A(n_124),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_126),
.A2(n_128),
.B1(n_68),
.B2(n_81),
.Y(n_131)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_98),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_127),
.B(n_88),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_102),
.A2(n_50),
.B1(n_72),
.B2(n_43),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_SL g171 ( 
.A1(n_129),
.A2(n_142),
.B(n_143),
.Y(n_171)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_130),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_131),
.A2(n_135),
.B1(n_120),
.B2(n_107),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_123),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_132),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_127),
.A2(n_97),
.B1(n_101),
.B2(n_94),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_109),
.B(n_91),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_136),
.B(n_137),
.Y(n_154)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_116),
.Y(n_137)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_116),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_138),
.B(n_140),
.Y(n_151)
);

AO21x2_ASAP7_75t_SL g139 ( 
.A1(n_117),
.A2(n_90),
.B(n_95),
.Y(n_139)
);

AO22x2_ASAP7_75t_L g169 ( 
.A1(n_139),
.A2(n_126),
.B1(n_109),
.B2(n_45),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g140 ( 
.A(n_125),
.Y(n_140)
);

AND2x2_ASAP7_75t_L g142 ( 
.A(n_110),
.B(n_95),
.Y(n_142)
);

CKINVDCx16_ASAP7_75t_R g144 ( 
.A(n_128),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_144),
.B(n_148),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_L g165 ( 
.A1(n_145),
.A2(n_147),
.B(n_139),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_110),
.B(n_112),
.Y(n_146)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_146),
.Y(n_162)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_128),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_112),
.B(n_68),
.Y(n_149)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_149),
.Y(n_168)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_125),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_150),
.B(n_114),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_152),
.A2(n_156),
.B1(n_148),
.B2(n_137),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_144),
.A2(n_122),
.B1(n_118),
.B2(n_111),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_153),
.A2(n_159),
.B1(n_163),
.B2(n_131),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g157 ( 
.A(n_145),
.B(n_113),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_157),
.B(n_158),
.C(n_161),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_132),
.B(n_120),
.C(n_111),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_139),
.A2(n_118),
.B1(n_120),
.B2(n_119),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_139),
.B(n_121),
.C(n_115),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_139),
.A2(n_126),
.B1(n_121),
.B2(n_107),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_133),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_164),
.B(n_166),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_165),
.B(n_135),
.Y(n_182)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_133),
.Y(n_166)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_167),
.Y(n_172)
);

AOI21xp5_ASAP7_75t_L g178 ( 
.A1(n_169),
.A2(n_129),
.B(n_130),
.Y(n_178)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_149),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_170),
.B(n_146),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_173),
.A2(n_181),
.B1(n_185),
.B2(n_189),
.Y(n_191)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_151),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_175),
.B(n_179),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_SL g177 ( 
.A(n_159),
.B(n_141),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_177),
.B(n_182),
.Y(n_197)
);

OAI21xp33_ASAP7_75t_L g198 ( 
.A1(n_178),
.A2(n_184),
.B(n_188),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_154),
.B(n_114),
.Y(n_179)
);

CKINVDCx16_ASAP7_75t_R g200 ( 
.A(n_180),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_161),
.A2(n_136),
.B1(n_141),
.B2(n_150),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_183),
.B(n_186),
.Y(n_192)
);

AOI21xp5_ASAP7_75t_L g184 ( 
.A1(n_171),
.A2(n_143),
.B(n_147),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_169),
.A2(n_147),
.B1(n_142),
.B2(n_134),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_171),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_157),
.B(n_142),
.C(n_134),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_187),
.B(n_158),
.C(n_165),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_162),
.B(n_124),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_169),
.A2(n_134),
.B1(n_124),
.B2(n_66),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_173),
.B(n_160),
.Y(n_193)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_193),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_194),
.B(n_203),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_187),
.B(n_155),
.C(n_170),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_195),
.B(n_196),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_174),
.B(n_155),
.C(n_168),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_174),
.B(n_168),
.C(n_162),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_SL g206 ( 
.A(n_199),
.B(n_201),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_181),
.B(n_153),
.C(n_163),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_L g202 ( 
.A1(n_184),
.A2(n_169),
.B(n_19),
.Y(n_202)
);

AOI21xp5_ASAP7_75t_L g210 ( 
.A1(n_202),
.A2(n_172),
.B(n_185),
.Y(n_210)
);

AOI21x1_ASAP7_75t_SL g203 ( 
.A1(n_177),
.A2(n_0),
.B(n_1),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_178),
.B(n_182),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_204),
.B(n_66),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_190),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_205),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_191),
.A2(n_189),
.B1(n_176),
.B2(n_188),
.Y(n_209)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_209),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_210),
.B(n_213),
.Y(n_226)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_204),
.Y(n_211)
);

AOI21xp5_ASAP7_75t_L g218 ( 
.A1(n_211),
.A2(n_216),
.B(n_203),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_192),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_214)
);

INVxp67_ASAP7_75t_L g220 ( 
.A(n_214),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_197),
.B(n_9),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_215),
.B(n_194),
.C(n_199),
.Y(n_219)
);

AOI21xp5_ASAP7_75t_L g216 ( 
.A1(n_195),
.A2(n_10),
.B(n_4),
.Y(n_216)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_218),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_219),
.B(n_212),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_214),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_221),
.B(n_198),
.Y(n_234)
);

INVxp67_ASAP7_75t_L g222 ( 
.A(n_206),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_222),
.B(n_212),
.Y(n_227)
);

AO221x1_ASAP7_75t_L g223 ( 
.A1(n_213),
.A2(n_200),
.B1(n_198),
.B2(n_196),
.C(n_197),
.Y(n_223)
);

NOR2xp67_ASAP7_75t_SL g230 ( 
.A(n_223),
.B(n_215),
.Y(n_230)
);

HB1xp67_ASAP7_75t_L g225 ( 
.A(n_207),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_225),
.B(n_208),
.Y(n_231)
);

AOI21xp5_ASAP7_75t_L g237 ( 
.A1(n_227),
.A2(n_230),
.B(n_231),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_229),
.B(n_234),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_222),
.B(n_10),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_232),
.B(n_233),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_220),
.B(n_11),
.Y(n_233)
);

AOI322xp5_ASAP7_75t_L g235 ( 
.A1(n_228),
.A2(n_224),
.A3(n_217),
.B1(n_226),
.B2(n_220),
.C1(n_7),
.C2(n_11),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_235),
.B(n_240),
.C(n_5),
.Y(n_242)
);

HB1xp67_ASAP7_75t_L g236 ( 
.A(n_227),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_236),
.B(n_1),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_229),
.B(n_7),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_SL g241 ( 
.A1(n_237),
.A2(n_11),
.B(n_4),
.Y(n_241)
);

AOI21x1_ASAP7_75t_L g245 ( 
.A1(n_241),
.A2(n_244),
.B(n_238),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_242),
.B(n_243),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_SL g244 ( 
.A1(n_239),
.A2(n_5),
.B(n_6),
.Y(n_244)
);

INVxp67_ASAP7_75t_L g247 ( 
.A(n_245),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_247),
.B(n_246),
.C(n_235),
.Y(n_248)
);

OAI321xp33_ASAP7_75t_L g249 ( 
.A1(n_248),
.A2(n_14),
.A3(n_6),
.B1(n_12),
.B2(n_13),
.C(n_1),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_249),
.B(n_14),
.Y(n_250)
);


endmodule