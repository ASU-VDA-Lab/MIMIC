module fake_jpeg_5318_n_69 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_8, n_15, n_7, n_69);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_8;
input n_15;
input n_7;

output n_69;

wire n_61;
wire n_45;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_59;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_65;
wire n_34;
wire n_39;
wire n_42;
wire n_49;
wire n_38;
wire n_56;
wire n_50;
wire n_67;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_40;
wire n_35;
wire n_48;
wire n_46;
wire n_44;
wire n_36;
wire n_62;
wire n_37;
wire n_43;
wire n_32;
wire n_66;

INVx2_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_18),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_26),
.B(n_29),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_31),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_30),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_0),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_9),
.Y(n_39)
);

INVx13_ASAP7_75t_L g40 ( 
.A(n_22),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_7),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_24),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_19),
.Y(n_43)
);

HB1xp67_ASAP7_75t_L g44 ( 
.A(n_39),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_44),
.B(n_40),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_43),
.B(n_1),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_45),
.B(n_46),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g46 ( 
.A1(n_34),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_36),
.B(n_5),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g50 ( 
.A(n_47),
.B(n_35),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_32),
.Y(n_48)
);

INVx4_ASAP7_75t_SL g53 ( 
.A(n_48),
.Y(n_53)
);

AOI22x1_ASAP7_75t_SL g49 ( 
.A1(n_33),
.A2(n_6),
.B1(n_8),
.B2(n_10),
.Y(n_49)
);

AOI21xp5_ASAP7_75t_L g51 ( 
.A1(n_49),
.A2(n_41),
.B(n_38),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_50),
.B(n_51),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g52 ( 
.A(n_49),
.B(n_37),
.Y(n_52)
);

INVx1_ASAP7_75t_SL g59 ( 
.A(n_52),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g54 ( 
.A(n_49),
.B(n_42),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_54),
.B(n_56),
.Y(n_58)
);

CKINVDCx16_ASAP7_75t_R g57 ( 
.A(n_55),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_58),
.B(n_11),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_L g61 ( 
.A1(n_59),
.A2(n_53),
.B1(n_12),
.B2(n_13),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_61),
.B(n_62),
.Y(n_63)
);

OAI21xp5_ASAP7_75t_L g64 ( 
.A1(n_63),
.A2(n_60),
.B(n_57),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_64),
.A2(n_15),
.B1(n_17),
.B2(n_20),
.Y(n_65)
);

OAI21x1_ASAP7_75t_L g66 ( 
.A1(n_65),
.A2(n_21),
.B(n_23),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_66),
.Y(n_67)
);

AOI21xp5_ASAP7_75t_L g68 ( 
.A1(n_67),
.A2(n_25),
.B(n_27),
.Y(n_68)
);

XOR2xp5_ASAP7_75t_L g69 ( 
.A(n_68),
.B(n_28),
.Y(n_69)
);


endmodule