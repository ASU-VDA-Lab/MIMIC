module real_jpeg_25169_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_18;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_330;
wire n_298;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_343;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_299;
wire n_243;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_0),
.A2(n_78),
.B1(n_87),
.B2(n_89),
.Y(n_86)
);

CKINVDCx16_ASAP7_75t_R g89 ( 
.A(n_0),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_0),
.A2(n_33),
.B1(n_34),
.B2(n_89),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_SL g184 ( 
.A1(n_0),
.A2(n_27),
.B1(n_28),
.B2(n_89),
.Y(n_184)
);

AOI22xp33_ASAP7_75t_L g236 ( 
.A1(n_0),
.A2(n_64),
.B1(n_68),
.B2(n_89),
.Y(n_236)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_1),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_2),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_2),
.B(n_55),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_2),
.B(n_28),
.C(n_30),
.Y(n_251)
);

AOI22xp33_ASAP7_75t_L g262 ( 
.A1(n_2),
.A2(n_33),
.B1(n_34),
.B2(n_198),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_2),
.B(n_37),
.Y(n_280)
);

AOI22xp33_ASAP7_75t_L g291 ( 
.A1(n_2),
.A2(n_27),
.B1(n_28),
.B2(n_198),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_2),
.B(n_64),
.C(n_67),
.Y(n_293)
);

OAI21xp5_ASAP7_75t_L g315 ( 
.A1(n_2),
.A2(n_102),
.B(n_285),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_3),
.A2(n_50),
.B1(n_51),
.B2(n_57),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_3),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_3),
.A2(n_33),
.B1(n_34),
.B2(n_57),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_3),
.A2(n_27),
.B1(n_28),
.B2(n_57),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_3),
.A2(n_57),
.B1(n_64),
.B2(n_68),
.Y(n_134)
);

BUFx12f_ASAP7_75t_L g67 ( 
.A(n_4),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_5),
.A2(n_45),
.B1(n_50),
.B2(n_174),
.Y(n_173)
);

CKINVDCx16_ASAP7_75t_R g174 ( 
.A(n_5),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_5),
.A2(n_33),
.B1(n_34),
.B2(n_174),
.Y(n_220)
);

AOI22xp33_ASAP7_75t_L g258 ( 
.A1(n_5),
.A2(n_27),
.B1(n_28),
.B2(n_174),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_5),
.A2(n_64),
.B1(n_68),
.B2(n_174),
.Y(n_298)
);

BUFx10_ASAP7_75t_L g65 ( 
.A(n_6),
.Y(n_65)
);

BUFx10_ASAP7_75t_L g52 ( 
.A(n_7),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_8),
.A2(n_45),
.B1(n_46),
.B2(n_145),
.Y(n_144)
);

CKINVDCx16_ASAP7_75t_R g145 ( 
.A(n_8),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_8),
.A2(n_33),
.B1(n_34),
.B2(n_145),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g259 ( 
.A1(n_8),
.A2(n_27),
.B1(n_28),
.B2(n_145),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_8),
.A2(n_64),
.B1(n_68),
.B2(n_145),
.Y(n_284)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

INVx13_ASAP7_75t_L g46 ( 
.A(n_10),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_11),
.A2(n_46),
.B1(n_78),
.B2(n_79),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_11),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_11),
.A2(n_33),
.B1(n_34),
.B2(n_79),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_11),
.A2(n_27),
.B1(n_28),
.B2(n_79),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_L g203 ( 
.A1(n_11),
.A2(n_64),
.B1(n_68),
.B2(n_79),
.Y(n_203)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

AOI22xp33_ASAP7_75t_SL g43 ( 
.A1(n_13),
.A2(n_44),
.B1(n_45),
.B2(n_47),
.Y(n_43)
);

CKINVDCx16_ASAP7_75t_R g47 ( 
.A(n_13),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_13),
.A2(n_33),
.B1(n_34),
.B2(n_47),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_13),
.A2(n_27),
.B1(n_28),
.B2(n_47),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_13),
.A2(n_47),
.B1(n_64),
.B2(n_68),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_SL g39 ( 
.A1(n_14),
.A2(n_33),
.B1(n_34),
.B2(n_40),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_14),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_14),
.A2(n_27),
.B1(n_28),
.B2(n_40),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_14),
.A2(n_40),
.B1(n_64),
.B2(n_68),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_L g118 ( 
.A1(n_15),
.A2(n_78),
.B1(n_119),
.B2(n_120),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_15),
.Y(n_120)
);

OAI22xp33_ASAP7_75t_SL g178 ( 
.A1(n_15),
.A2(n_33),
.B1(n_34),
.B2(n_120),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_15),
.A2(n_27),
.B1(n_28),
.B2(n_120),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_15),
.A2(n_64),
.B1(n_68),
.B2(n_120),
.Y(n_255)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_16),
.Y(n_103)
);

INVx6_ASAP7_75t_L g106 ( 
.A(n_16),
.Y(n_106)
);

INVx6_ASAP7_75t_L g135 ( 
.A(n_16),
.Y(n_135)
);

INVx3_ASAP7_75t_L g300 ( 
.A(n_16),
.Y(n_300)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_96),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_95),
.Y(n_18)
);

INVxp67_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_80),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_21),
.B(n_80),
.Y(n_95)
);

XNOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_60),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_41),
.B1(n_58),
.B2(n_59),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_23),
.Y(n_58)
);

OAI21xp5_ASAP7_75t_SL g23 ( 
.A1(n_24),
.A2(n_37),
.B(n_38),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_24),
.A2(n_37),
.B1(n_92),
.B2(n_94),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_24),
.B(n_178),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_24),
.A2(n_37),
.B1(n_192),
.B2(n_220),
.Y(n_219)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_25),
.A2(n_26),
.B1(n_39),
.B2(n_74),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_25),
.A2(n_26),
.B1(n_93),
.B2(n_124),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_25),
.A2(n_26),
.B1(n_124),
.B2(n_141),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_SL g190 ( 
.A1(n_25),
.A2(n_191),
.B(n_193),
.Y(n_190)
);

OAI21xp33_ASAP7_75t_L g261 ( 
.A1(n_25),
.A2(n_193),
.B(n_262),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_32),
.Y(n_25)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

OAI21xp5_ASAP7_75t_L g176 ( 
.A1(n_26),
.A2(n_141),
.B(n_177),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_SL g231 ( 
.A1(n_26),
.A2(n_177),
.B(n_232),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_SL g26 ( 
.A1(n_27),
.A2(n_28),
.B1(n_30),
.B2(n_31),
.Y(n_26)
);

OAI22xp33_ASAP7_75t_L g70 ( 
.A1(n_27),
.A2(n_28),
.B1(n_66),
.B2(n_67),
.Y(n_70)
);

INVx3_ASAP7_75t_SL g27 ( 
.A(n_28),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_28),
.B(n_293),
.Y(n_292)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx5_ASAP7_75t_L g31 ( 
.A(n_30),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_L g32 ( 
.A1(n_30),
.A2(n_31),
.B1(n_33),
.B2(n_34),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_L g55 ( 
.A1(n_33),
.A2(n_34),
.B1(n_52),
.B2(n_53),
.Y(n_55)
);

NAND3xp33_ASAP7_75t_SL g199 ( 
.A(n_33),
.B(n_45),
.C(n_53),
.Y(n_199)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

A2O1A1Ixp33_ASAP7_75t_L g196 ( 
.A1(n_34),
.A2(n_52),
.B(n_197),
.C(n_199),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_34),
.B(n_251),
.Y(n_250)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_37),
.B(n_178),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_39),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_41),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g41 ( 
.A1(n_42),
.A2(n_48),
.B1(n_55),
.B2(n_56),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_43),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_43),
.A2(n_54),
.B1(n_76),
.B2(n_77),
.Y(n_75)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

OAI22xp33_ASAP7_75t_L g49 ( 
.A1(n_45),
.A2(n_50),
.B1(n_52),
.B2(n_53),
.Y(n_49)
);

INVx11_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_46),
.Y(n_51)
);

INVx8_ASAP7_75t_L g78 ( 
.A(n_46),
.Y(n_78)
);

INVx6_ASAP7_75t_L g88 ( 
.A(n_46),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_48),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_48),
.B(n_117),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_48),
.A2(n_55),
.B1(n_144),
.B2(n_173),
.Y(n_172)
);

AOI21xp5_ASAP7_75t_L g225 ( 
.A1(n_48),
.A2(n_147),
.B(n_226),
.Y(n_225)
);

AND2x2_ASAP7_75t_L g48 ( 
.A(n_49),
.B(n_54),
.Y(n_48)
);

INVx11_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_52),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_54),
.A2(n_76),
.B1(n_77),
.B2(n_86),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_L g115 ( 
.A1(n_54),
.A2(n_86),
.B(n_116),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_54),
.B(n_118),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_L g188 ( 
.A1(n_54),
.A2(n_116),
.B(n_189),
.Y(n_188)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

MAJIxp5_ASAP7_75t_L g60 ( 
.A(n_61),
.B(n_73),
.C(n_75),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_61),
.A2(n_73),
.B1(n_83),
.B2(n_84),
.Y(n_82)
);

CKINVDCx14_ASAP7_75t_R g84 ( 
.A(n_61),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_61),
.B(n_85),
.C(n_91),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_61),
.A2(n_84),
.B1(n_91),
.B2(n_156),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_L g61 ( 
.A1(n_62),
.A2(n_69),
.B(n_71),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_62),
.A2(n_69),
.B1(n_110),
.B2(n_111),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_62),
.A2(n_69),
.B1(n_110),
.B2(n_138),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_62),
.A2(n_69),
.B1(n_257),
.B2(n_259),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_62),
.B(n_224),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_63),
.Y(n_62)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_63),
.B(n_70),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_63),
.A2(n_72),
.B1(n_126),
.B2(n_127),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_63),
.A2(n_126),
.B1(n_139),
.B2(n_184),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_L g222 ( 
.A1(n_63),
.A2(n_184),
.B(n_223),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_L g282 ( 
.A1(n_63),
.A2(n_223),
.B(n_258),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_63),
.B(n_198),
.Y(n_306)
);

OA22x2_ASAP7_75t_L g63 ( 
.A1(n_64),
.A2(n_66),
.B1(n_67),
.B2(n_68),
.Y(n_63)
);

INVx2_ASAP7_75t_SL g68 ( 
.A(n_64),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_64),
.B(n_103),
.Y(n_102)
);

BUFx4f_ASAP7_75t_SL g64 ( 
.A(n_65),
.Y(n_64)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_68),
.B(n_312),
.Y(n_311)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_69),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_69),
.B(n_224),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_72),
.Y(n_71)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_73),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_74),
.Y(n_94)
);

XNOR2xp5_ASAP7_75t_L g81 ( 
.A(n_75),
.B(n_82),
.Y(n_81)
);

OAI21xp5_ASAP7_75t_L g142 ( 
.A1(n_76),
.A2(n_143),
.B(n_146),
.Y(n_142)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_78),
.Y(n_119)
);

OAI21xp33_ASAP7_75t_SL g226 ( 
.A1(n_78),
.A2(n_197),
.B(n_198),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_85),
.C(n_90),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_81),
.A2(n_85),
.B1(n_157),
.B2(n_162),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_81),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_85),
.A2(n_154),
.B1(n_155),
.B2(n_157),
.Y(n_153)
);

CKINVDCx14_ASAP7_75t_R g157 ( 
.A(n_85),
.Y(n_157)
);

INVx8_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

NAND2xp33_ASAP7_75t_SL g197 ( 
.A(n_88),
.B(n_198),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_90),
.B(n_161),
.Y(n_160)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_91),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_93),
.Y(n_92)
);

OAI31xp33_ASAP7_75t_SL g96 ( 
.A1(n_97),
.A2(n_158),
.A3(n_164),
.B(n_347),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_148),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g348 ( 
.A(n_98),
.B(n_148),
.Y(n_348)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_121),
.C(n_129),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g342 ( 
.A1(n_99),
.A2(n_121),
.B1(n_122),
.B2(n_343),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_99),
.Y(n_343)
);

XOR2xp5_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_112),
.Y(n_99)
);

AOI21xp33_ASAP7_75t_L g149 ( 
.A1(n_100),
.A2(n_101),
.B(n_114),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_108),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_101),
.A2(n_113),
.B1(n_114),
.B2(n_115),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_101),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_101),
.A2(n_108),
.B1(n_109),
.B2(n_113),
.Y(n_207)
);

AOI21xp5_ASAP7_75t_L g101 ( 
.A1(n_102),
.A2(n_104),
.B(n_107),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_102),
.A2(n_107),
.B1(n_134),
.B2(n_135),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_102),
.A2(n_134),
.B1(n_135),
.B2(n_181),
.Y(n_180)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_102),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_102),
.A2(n_135),
.B1(n_203),
.B2(n_236),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_102),
.B(n_255),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_L g283 ( 
.A1(n_102),
.A2(n_284),
.B(n_285),
.Y(n_283)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_103),
.Y(n_286)
);

BUFx2_ASAP7_75t_L g308 ( 
.A(n_103),
.Y(n_308)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

AOI21xp5_ASAP7_75t_L g252 ( 
.A1(n_105),
.A2(n_253),
.B(n_254),
.Y(n_252)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

CKINVDCx16_ASAP7_75t_R g108 ( 
.A(n_109),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_111),
.Y(n_127)
);

CKINVDCx16_ASAP7_75t_R g114 ( 
.A(n_115),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

AOI21xp5_ASAP7_75t_L g122 ( 
.A1(n_123),
.A2(n_125),
.B(n_128),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_123),
.B(n_125),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_SL g271 ( 
.A1(n_126),
.A2(n_272),
.B(n_273),
.Y(n_271)
);

OAI21xp5_ASAP7_75t_SL g290 ( 
.A1(n_126),
.A2(n_273),
.B(n_291),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_128),
.A2(n_151),
.B1(n_152),
.B2(n_153),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_128),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g341 ( 
.A1(n_129),
.A2(n_130),
.B1(n_342),
.B2(n_344),
.Y(n_341)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_140),
.C(n_142),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_131),
.A2(n_132),
.B1(n_209),
.B2(n_210),
.Y(n_208)
);

CKINVDCx14_ASAP7_75t_R g131 ( 
.A(n_132),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_136),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_133),
.A2(n_136),
.B1(n_137),
.B2(n_186),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_133),
.Y(n_186)
);

INVx8_ASAP7_75t_L g204 ( 
.A(n_135),
.Y(n_204)
);

INVx5_ASAP7_75t_L g314 ( 
.A(n_135),
.Y(n_314)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_139),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_SL g210 ( 
.A(n_140),
.B(n_142),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_144),
.Y(n_143)
);

INVxp67_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

XOR2xp5_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_150),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_149),
.B(n_151),
.C(n_153),
.Y(n_163)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVxp67_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

AOI21xp5_ASAP7_75t_L g347 ( 
.A1(n_159),
.A2(n_348),
.B(n_349),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_160),
.B(n_163),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_160),
.B(n_163),
.Y(n_349)
);

AOI21xp5_ASAP7_75t_L g164 ( 
.A1(n_165),
.A2(n_340),
.B(n_346),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_L g165 ( 
.A1(n_166),
.A2(n_212),
.B(n_339),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_205),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_167),
.B(n_205),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_185),
.C(n_187),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g336 ( 
.A1(n_168),
.A2(n_169),
.B1(n_185),
.B2(n_337),
.Y(n_336)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_179),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_171),
.A2(n_172),
.B1(n_175),
.B2(n_176),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_172),
.B(n_175),
.C(n_179),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_173),
.Y(n_189)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_183),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_180),
.B(n_183),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_182),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_182),
.A2(n_201),
.B1(n_202),
.B2(n_204),
.Y(n_200)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_185),
.Y(n_337)
);

XNOR2xp5_ASAP7_75t_L g335 ( 
.A(n_187),
.B(n_336),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_188),
.B(n_190),
.C(n_194),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_188),
.B(n_190),
.Y(n_239)
);

CKINVDCx16_ASAP7_75t_R g191 ( 
.A(n_192),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_SL g238 ( 
.A(n_194),
.B(n_239),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_200),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_195),
.A2(n_196),
.B1(n_200),
.B2(n_229),
.Y(n_228)
);

CKINVDCx16_ASAP7_75t_R g195 ( 
.A(n_196),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_198),
.B(n_313),
.Y(n_312)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_200),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_201),
.A2(n_297),
.B1(n_299),
.B2(n_301),
.Y(n_296)
);

INVxp67_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_211),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_208),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_207),
.B(n_208),
.C(n_211),
.Y(n_345)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

O2A1O1Ixp33_ASAP7_75t_SL g212 ( 
.A1(n_213),
.A2(n_243),
.B(n_333),
.C(n_338),
.Y(n_212)
);

AND2x2_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_237),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_214),
.B(n_237),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_227),
.C(n_230),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g327 ( 
.A1(n_215),
.A2(n_216),
.B1(n_328),
.B2(n_329),
.Y(n_327)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_225),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_218),
.A2(n_219),
.B1(n_221),
.B2(n_222),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_219),
.B(n_221),
.C(n_225),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_220),
.Y(n_232)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g329 ( 
.A1(n_227),
.A2(n_228),
.B1(n_230),
.B2(n_330),
.Y(n_329)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_230),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_233),
.C(n_235),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_231),
.B(n_266),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_233),
.A2(n_234),
.B1(n_235),
.B2(n_267),
.Y(n_266)
);

CKINVDCx16_ASAP7_75t_R g233 ( 
.A(n_234),
.Y(n_233)
);

CKINVDCx16_ASAP7_75t_R g267 ( 
.A(n_235),
.Y(n_267)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_236),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_238),
.B(n_240),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_238),
.B(n_241),
.C(n_242),
.Y(n_334)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_242),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_245),
.Y(n_243)
);

AOI21xp5_ASAP7_75t_SL g245 ( 
.A1(n_246),
.A2(n_326),
.B(n_332),
.Y(n_245)
);

OAI21xp5_ASAP7_75t_L g246 ( 
.A1(n_247),
.A2(n_274),
.B(n_325),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_263),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_248),
.B(n_263),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_256),
.C(n_260),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_249),
.B(n_321),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_SL g249 ( 
.A(n_250),
.B(n_252),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_250),
.B(n_252),
.Y(n_270)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_254),
.Y(n_309)
);

CKINVDCx14_ASAP7_75t_R g287 ( 
.A(n_255),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_256),
.A2(n_260),
.B1(n_261),
.B2(n_322),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_256),
.Y(n_322)
);

INVxp67_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_259),
.Y(n_272)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_264),
.A2(n_265),
.B1(n_268),
.B2(n_269),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_264),
.B(n_270),
.C(n_271),
.Y(n_331)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_270),
.B(n_271),
.Y(n_269)
);

AOI21xp5_ASAP7_75t_L g274 ( 
.A1(n_275),
.A2(n_319),
.B(n_324),
.Y(n_274)
);

OAI21xp5_ASAP7_75t_SL g275 ( 
.A1(n_276),
.A2(n_294),
.B(n_318),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_SL g276 ( 
.A(n_277),
.B(n_288),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_277),
.B(n_288),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_278),
.B(n_283),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_279),
.A2(n_280),
.B1(n_281),
.B2(n_282),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_279),
.B(n_282),
.C(n_283),
.Y(n_323)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

INVxp67_ASAP7_75t_L g301 ( 
.A(n_284),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_286),
.B(n_287),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_SL g288 ( 
.A(n_289),
.B(n_292),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_289),
.A2(n_290),
.B1(n_292),
.B2(n_303),
.Y(n_302)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_292),
.Y(n_303)
);

AOI21xp5_ASAP7_75t_L g294 ( 
.A1(n_295),
.A2(n_304),
.B(n_317),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_296),
.B(n_302),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_296),
.B(n_302),
.Y(n_317)
);

INVxp67_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_L g307 ( 
.A1(n_298),
.A2(n_308),
.B(n_309),
.Y(n_307)
);

INVx3_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

OAI21xp5_ASAP7_75t_SL g304 ( 
.A1(n_305),
.A2(n_310),
.B(n_316),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_306),
.B(n_307),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_306),
.B(n_307),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_311),
.B(n_315),
.Y(n_310)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_SL g319 ( 
.A(n_320),
.B(n_323),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_320),
.B(n_323),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_SL g326 ( 
.A(n_327),
.B(n_331),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_327),
.B(n_331),
.Y(n_332)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_334),
.B(n_335),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_334),
.B(n_335),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_SL g340 ( 
.A(n_341),
.B(n_345),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_341),
.B(n_345),
.Y(n_346)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_342),
.Y(n_344)
);


endmodule