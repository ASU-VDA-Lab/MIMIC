module fake_jpeg_26391_n_325 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_325);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_325;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

INVxp67_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_8),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

CKINVDCx16_ASAP7_75t_R g25 ( 
.A(n_9),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_0),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

BUFx10_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_9),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_0),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_20),
.Y(n_36)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_36),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_20),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_37),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_23),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_SL g47 ( 
.A(n_38),
.B(n_43),
.Y(n_47)
);

INVx5_ASAP7_75t_L g39 ( 
.A(n_20),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_39),
.Y(n_49)
);

BUFx3_ASAP7_75t_SL g40 ( 
.A(n_32),
.Y(n_40)
);

BUFx10_ASAP7_75t_L g61 ( 
.A(n_40),
.Y(n_61)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_32),
.Y(n_41)
);

HAxp5_ASAP7_75t_SL g56 ( 
.A(n_41),
.B(n_33),
.CON(n_56),
.SN(n_56)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_20),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_42),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_20),
.B(n_8),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_23),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_44),
.B(n_45),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_26),
.Y(n_45)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_46),
.B(n_62),
.Y(n_70)
);

HB1xp67_ASAP7_75t_L g48 ( 
.A(n_40),
.Y(n_48)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_48),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_38),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_50),
.Y(n_72)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_53),
.B(n_64),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_44),
.B(n_21),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_54),
.B(n_28),
.Y(n_104)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

INVx4_ASAP7_75t_SL g83 ( 
.A(n_55),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_56),
.B(n_40),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g57 ( 
.A1(n_43),
.A2(n_41),
.B1(n_42),
.B2(n_39),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_57),
.A2(n_40),
.B1(n_25),
.B2(n_17),
.Y(n_77)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_58),
.Y(n_91)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_36),
.Y(n_62)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_36),
.Y(n_63)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_63),
.Y(n_103)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_40),
.Y(n_64)
);

NAND2xp33_ASAP7_75t_SL g65 ( 
.A(n_37),
.B(n_33),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_65),
.A2(n_27),
.B1(n_19),
.B2(n_30),
.Y(n_105)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_37),
.Y(n_66)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_66),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_45),
.B(n_32),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_67),
.B(n_32),
.Y(n_85)
);

HB1xp67_ASAP7_75t_L g68 ( 
.A(n_67),
.Y(n_68)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_68),
.Y(n_113)
);

CKINVDCx16_ASAP7_75t_R g69 ( 
.A(n_57),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_69),
.B(n_74),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_56),
.A2(n_41),
.B1(n_42),
.B2(n_39),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_71),
.A2(n_87),
.B1(n_106),
.B2(n_19),
.Y(n_108)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_52),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_73),
.Y(n_117)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_52),
.Y(n_74)
);

OAI21xp5_ASAP7_75t_L g75 ( 
.A1(n_47),
.A2(n_40),
.B(n_35),
.Y(n_75)
);

CKINVDCx14_ASAP7_75t_R g111 ( 
.A(n_75),
.Y(n_111)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_61),
.Y(n_76)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_76),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_77),
.A2(n_86),
.B1(n_102),
.B2(n_22),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_51),
.B(n_33),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_78),
.B(n_90),
.Y(n_126)
);

INVx5_ASAP7_75t_L g79 ( 
.A(n_60),
.Y(n_79)
);

INVxp33_ASAP7_75t_L g132 ( 
.A(n_79),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_53),
.B(n_64),
.C(n_66),
.Y(n_80)
);

XNOR2xp5_ASAP7_75t_L g121 ( 
.A(n_80),
.B(n_94),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_59),
.B(n_18),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_84),
.B(n_85),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_46),
.A2(n_26),
.B1(n_35),
.B2(n_17),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_59),
.A2(n_40),
.B1(n_34),
.B2(n_18),
.Y(n_87)
);

OR2x2_ASAP7_75t_L g116 ( 
.A(n_88),
.B(n_92),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_60),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_89),
.Y(n_118)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_61),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_60),
.B(n_33),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_60),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_93),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_63),
.B(n_33),
.C(n_31),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_L g95 ( 
.A1(n_62),
.A2(n_34),
.B1(n_32),
.B2(n_31),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_95),
.A2(n_98),
.B1(n_105),
.B2(n_29),
.Y(n_127)
);

BUFx2_ASAP7_75t_L g96 ( 
.A(n_49),
.Y(n_96)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_96),
.Y(n_115)
);

INVx8_ASAP7_75t_L g97 ( 
.A(n_61),
.Y(n_97)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_97),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_49),
.B(n_22),
.Y(n_98)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_55),
.Y(n_99)
);

BUFx2_ASAP7_75t_L g109 ( 
.A(n_99),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_58),
.B(n_27),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_100),
.B(n_28),
.Y(n_112)
);

OAI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_61),
.A2(n_25),
.B1(n_34),
.B2(n_31),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_104),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_56),
.A2(n_34),
.B1(n_16),
.B2(n_30),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_67),
.Y(n_107)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_107),
.Y(n_120)
);

AND2x2_ASAP7_75t_L g141 ( 
.A(n_108),
.B(n_127),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_112),
.B(n_129),
.Y(n_150)
);

BUFx8_ASAP7_75t_L g122 ( 
.A(n_83),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g153 ( 
.A(n_122),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_79),
.A2(n_16),
.B1(n_29),
.B2(n_24),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_123),
.A2(n_83),
.B1(n_91),
.B2(n_103),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_107),
.B(n_31),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_125),
.B(n_128),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_85),
.B(n_28),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_82),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_82),
.B(n_24),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_130),
.B(n_81),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_88),
.A2(n_92),
.B1(n_105),
.B2(n_75),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_SL g160 ( 
.A1(n_133),
.A2(n_10),
.B(n_15),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_134),
.A2(n_106),
.B1(n_87),
.B2(n_73),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_72),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_135),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_71),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_137),
.A2(n_74),
.B1(n_99),
.B2(n_91),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_135),
.B(n_100),
.Y(n_138)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_138),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_140),
.A2(n_145),
.B1(n_147),
.B2(n_169),
.Y(n_199)
);

AND2x2_ASAP7_75t_L g142 ( 
.A(n_133),
.B(n_88),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g176 ( 
.A(n_142),
.Y(n_176)
);

O2A1O1Ixp33_ASAP7_75t_L g143 ( 
.A1(n_111),
.A2(n_97),
.B(n_76),
.C(n_70),
.Y(n_143)
);

OA21x2_ASAP7_75t_L g198 ( 
.A1(n_143),
.A2(n_148),
.B(n_122),
.Y(n_198)
);

AOI21xp5_ASAP7_75t_L g144 ( 
.A1(n_116),
.A2(n_92),
.B(n_101),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g182 ( 
.A(n_144),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_136),
.A2(n_129),
.B1(n_120),
.B2(n_116),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_109),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_146),
.B(n_152),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_120),
.A2(n_113),
.B1(n_125),
.B2(n_134),
.Y(n_147)
);

AOI21xp5_ASAP7_75t_L g148 ( 
.A1(n_121),
.A2(n_81),
.B(n_80),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_149),
.B(n_158),
.Y(n_172)
);

CKINVDCx16_ASAP7_75t_R g185 ( 
.A(n_151),
.Y(n_185)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_109),
.Y(n_152)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_126),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_154),
.B(n_156),
.Y(n_192)
);

BUFx24_ASAP7_75t_SL g155 ( 
.A(n_110),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_155),
.B(n_163),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_121),
.B(n_94),
.C(n_90),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_157),
.B(n_148),
.C(n_142),
.Y(n_184)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_130),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_128),
.B(n_103),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_159),
.B(n_161),
.Y(n_173)
);

XNOR2x1_ASAP7_75t_L g194 ( 
.A(n_160),
.B(n_12),
.Y(n_194)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_112),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_118),
.B(n_10),
.Y(n_162)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_162),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_118),
.B(n_124),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_108),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_164),
.B(n_165),
.Y(n_175)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_124),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_137),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_166),
.B(n_114),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_132),
.B(n_10),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_167),
.Y(n_181)
);

AO21x2_ASAP7_75t_L g169 ( 
.A1(n_113),
.A2(n_114),
.B(n_119),
.Y(n_169)
);

OR2x2_ASAP7_75t_L g170 ( 
.A(n_147),
.B(n_131),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_L g219 ( 
.A1(n_170),
.A2(n_178),
.B(n_198),
.Y(n_219)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_169),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_177),
.B(n_180),
.Y(n_204)
);

OR2x2_ASAP7_75t_L g178 ( 
.A(n_141),
.B(n_131),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_SL g226 ( 
.A1(n_179),
.A2(n_194),
.B(n_201),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_139),
.B(n_110),
.Y(n_180)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_169),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_183),
.B(n_186),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_184),
.B(n_188),
.C(n_193),
.Y(n_208)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_169),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_169),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_187),
.B(n_197),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_157),
.B(n_119),
.C(n_115),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_168),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_189),
.Y(n_220)
);

INVx3_ASAP7_75t_L g190 ( 
.A(n_165),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_190),
.B(n_146),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_142),
.B(n_161),
.C(n_139),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_145),
.B(n_115),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_196),
.B(n_164),
.Y(n_206)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_159),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_150),
.B(n_117),
.C(n_122),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_200),
.B(n_202),
.C(n_149),
.Y(n_211)
);

OR2x2_ASAP7_75t_L g201 ( 
.A(n_141),
.B(n_156),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_144),
.B(n_117),
.C(n_122),
.Y(n_202)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_203),
.Y(n_244)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_174),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_205),
.B(n_209),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_SL g247 ( 
.A(n_206),
.B(n_216),
.Y(n_247)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_179),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_185),
.A2(n_166),
.B1(n_141),
.B2(n_160),
.Y(n_210)
);

INVxp67_ASAP7_75t_L g236 ( 
.A(n_210),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_211),
.B(n_229),
.Y(n_234)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_173),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_213),
.B(n_215),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_184),
.B(n_158),
.C(n_154),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_214),
.B(n_222),
.C(n_202),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_201),
.B(n_152),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_188),
.B(n_143),
.Y(n_216)
);

AND2x2_ASAP7_75t_SL g217 ( 
.A(n_177),
.B(n_153),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_217),
.Y(n_231)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_173),
.Y(n_218)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_218),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_183),
.A2(n_153),
.B1(n_96),
.B2(n_3),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_221),
.A2(n_228),
.B1(n_171),
.B2(n_191),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_193),
.B(n_8),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_175),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_223),
.Y(n_240)
);

INVx1_ASAP7_75t_SL g224 ( 
.A(n_198),
.Y(n_224)
);

INVxp67_ASAP7_75t_SL g250 ( 
.A(n_224),
.Y(n_250)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_175),
.Y(n_225)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_225),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_186),
.A2(n_7),
.B1(n_14),
.B2(n_13),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_227),
.A2(n_190),
.B1(n_170),
.B2(n_199),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_172),
.A2(n_15),
.B1(n_7),
.B2(n_11),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_SL g229 ( 
.A1(n_182),
.A2(n_0),
.B(n_2),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_181),
.B(n_7),
.Y(n_230)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_230),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_233),
.B(n_211),
.Y(n_259)
);

NOR3xp33_ASAP7_75t_SL g235 ( 
.A(n_220),
.B(n_194),
.C(n_192),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_235),
.B(n_219),
.Y(n_256)
);

AOI22x1_ASAP7_75t_SL g237 ( 
.A1(n_224),
.A2(n_198),
.B1(n_182),
.B2(n_178),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_237),
.A2(n_241),
.B1(n_245),
.B2(n_212),
.Y(n_271)
);

CKINVDCx14_ASAP7_75t_R g263 ( 
.A(n_238),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_208),
.B(n_196),
.C(n_197),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_239),
.B(n_243),
.C(n_251),
.Y(n_258)
);

AOI22x1_ASAP7_75t_L g241 ( 
.A1(n_212),
.A2(n_187),
.B1(n_199),
.B2(n_172),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_208),
.B(n_180),
.C(n_200),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_216),
.B(n_176),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_246),
.B(n_222),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_207),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_248),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_214),
.B(n_176),
.C(n_195),
.Y(n_251)
);

INVx6_ASAP7_75t_L g255 ( 
.A(n_241),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_255),
.B(n_266),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_SL g275 ( 
.A1(n_256),
.A2(n_260),
.B(n_236),
.Y(n_275)
);

FAx1_ASAP7_75t_SL g257 ( 
.A(n_247),
.B(n_219),
.CI(n_204),
.CON(n_257),
.SN(n_257)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_257),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_259),
.B(n_252),
.Y(n_287)
);

AOI21xp5_ASAP7_75t_L g260 ( 
.A1(n_236),
.A2(n_226),
.B(n_229),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_240),
.B(n_250),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_261),
.B(n_262),
.Y(n_279)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_232),
.Y(n_262)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_242),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_264),
.B(n_265),
.Y(n_282)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_235),
.Y(n_265)
);

CKINVDCx16_ASAP7_75t_R g266 ( 
.A(n_245),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_234),
.B(n_206),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_267),
.B(n_272),
.Y(n_276)
);

BUFx4f_ASAP7_75t_SL g268 ( 
.A(n_237),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_268),
.Y(n_286)
);

FAx1_ASAP7_75t_SL g269 ( 
.A(n_247),
.B(n_204),
.CI(n_226),
.CON(n_269),
.SN(n_269)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_269),
.B(n_271),
.Y(n_285)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_270),
.B(n_233),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_243),
.B(n_225),
.C(n_209),
.Y(n_272)
);

BUFx12_ASAP7_75t_L g273 ( 
.A(n_268),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_SL g295 ( 
.A(n_273),
.B(n_281),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_274),
.B(n_283),
.Y(n_291)
);

AOI21xp5_ASAP7_75t_L g298 ( 
.A1(n_275),
.A2(n_217),
.B(n_227),
.Y(n_298)
);

A2O1A1O1Ixp25_ASAP7_75t_L g277 ( 
.A1(n_257),
.A2(n_246),
.B(n_234),
.C(n_239),
.D(n_231),
.Y(n_277)
);

NAND3xp33_ASAP7_75t_L g288 ( 
.A(n_277),
.B(n_284),
.C(n_257),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_SL g281 ( 
.A(n_254),
.B(n_253),
.Y(n_281)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_270),
.B(n_251),
.Y(n_283)
);

NAND3xp33_ASAP7_75t_L g284 ( 
.A(n_255),
.B(n_210),
.C(n_217),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_287),
.B(n_244),
.C(n_268),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_L g301 ( 
.A1(n_288),
.A2(n_298),
.B(n_284),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_286),
.B(n_272),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_289),
.B(n_290),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_287),
.B(n_258),
.C(n_259),
.Y(n_290)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_279),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_292),
.B(n_294),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_280),
.A2(n_263),
.B1(n_285),
.B2(n_271),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_L g304 ( 
.A1(n_293),
.A2(n_278),
.B1(n_273),
.B2(n_277),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_276),
.B(n_258),
.C(n_267),
.Y(n_294)
);

BUFx24_ASAP7_75t_SL g296 ( 
.A(n_282),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_296),
.B(n_12),
.Y(n_309)
);

XOR2xp5_ASAP7_75t_L g303 ( 
.A(n_297),
.B(n_269),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_283),
.B(n_249),
.C(n_218),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_299),
.B(n_300),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_274),
.B(n_213),
.C(n_221),
.Y(n_300)
);

AOI21xp5_ASAP7_75t_SL g311 ( 
.A1(n_301),
.A2(n_291),
.B(n_13),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_303),
.B(n_304),
.Y(n_314)
);

AOI21xp5_ASAP7_75t_L g306 ( 
.A1(n_295),
.A2(n_273),
.B(n_269),
.Y(n_306)
);

OAI21xp5_ASAP7_75t_L g310 ( 
.A1(n_306),
.A2(n_288),
.B(n_294),
.Y(n_310)
);

HB1xp67_ASAP7_75t_L g307 ( 
.A(n_290),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_SL g312 ( 
.A1(n_307),
.A2(n_5),
.B1(n_6),
.B2(n_13),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_SL g315 ( 
.A(n_309),
.B(n_6),
.Y(n_315)
);

XOR2xp5_ASAP7_75t_L g316 ( 
.A(n_310),
.B(n_303),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_SL g318 ( 
.A(n_311),
.B(n_315),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_312),
.B(n_313),
.C(n_15),
.Y(n_317)
);

AOI21xp33_ASAP7_75t_L g313 ( 
.A1(n_302),
.A2(n_6),
.B(n_14),
.Y(n_313)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_316),
.Y(n_320)
);

OAI21xp5_ASAP7_75t_L g319 ( 
.A1(n_317),
.A2(n_314),
.B(n_308),
.Y(n_319)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_319),
.Y(n_321)
);

NOR3xp33_ASAP7_75t_L g322 ( 
.A(n_321),
.B(n_320),
.C(n_305),
.Y(n_322)
);

NOR3xp33_ASAP7_75t_SL g323 ( 
.A(n_322),
.B(n_307),
.C(n_318),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_323),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_L g325 ( 
.A(n_324),
.B(n_2),
.Y(n_325)
);


endmodule