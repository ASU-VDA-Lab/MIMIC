module fake_jpeg_21611_n_295 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_295);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_295;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_119;
wire n_23;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_145;
wire n_18;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_212;
wire n_131;
wire n_56;
wire n_240;
wire n_294;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_12;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_6),
.Y(n_12)
);

INVx6_ASAP7_75t_L g13 ( 
.A(n_2),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_8),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_7),
.Y(n_15)
);

BUFx3_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_3),
.Y(n_18)
);

CKINVDCx16_ASAP7_75t_R g19 ( 
.A(n_0),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_3),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_1),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_3),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_2),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_17),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_14),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_27),
.B(n_28),
.Y(n_39)
);

BUFx16f_ASAP7_75t_L g28 ( 
.A(n_19),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_19),
.B(n_12),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_29),
.B(n_30),
.Y(n_41)
);

INVx1_ASAP7_75t_SL g30 ( 
.A(n_17),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

BUFx12_ASAP7_75t_L g32 ( 
.A(n_19),
.Y(n_32)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_32),
.Y(n_38)
);

INVx1_ASAP7_75t_SL g33 ( 
.A(n_17),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_33),
.B(n_34),
.Y(n_44)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_17),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_35),
.B(n_24),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g36 ( 
.A1(n_30),
.A2(n_13),
.B1(n_19),
.B2(n_25),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g61 ( 
.A1(n_36),
.A2(n_42),
.B1(n_33),
.B2(n_30),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g42 ( 
.A1(n_30),
.A2(n_13),
.B1(n_14),
.B2(n_25),
.Y(n_42)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_43),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_30),
.A2(n_13),
.B1(n_15),
.B2(n_12),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_45),
.A2(n_33),
.B1(n_32),
.B2(n_13),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_46),
.B(n_32),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_27),
.B(n_24),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_47),
.B(n_27),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_48),
.B(n_49),
.Y(n_79)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_47),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g50 ( 
.A(n_41),
.B(n_28),
.Y(n_50)
);

OAI21xp33_ASAP7_75t_L g85 ( 
.A1(n_50),
.A2(n_51),
.B(n_66),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g51 ( 
.A(n_41),
.B(n_28),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_47),
.B(n_27),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_52),
.B(n_65),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_53),
.B(n_55),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_54),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_39),
.B(n_29),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

INVx8_ASAP7_75t_L g74 ( 
.A(n_56),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g57 ( 
.A(n_39),
.B(n_29),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_57),
.B(n_62),
.Y(n_82)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_40),
.Y(n_59)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_59),
.Y(n_80)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_60),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_61),
.A2(n_63),
.B1(n_38),
.B2(n_32),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g62 ( 
.A(n_42),
.B(n_12),
.Y(n_62)
);

INVx13_ASAP7_75t_L g64 ( 
.A(n_38),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g86 ( 
.A(n_64),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_46),
.B(n_35),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_42),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_66),
.A2(n_45),
.B1(n_33),
.B2(n_43),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_67),
.A2(n_70),
.B1(n_77),
.B2(n_81),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_58),
.A2(n_38),
.B1(n_43),
.B2(n_33),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_69),
.A2(n_75),
.B1(n_32),
.B2(n_13),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_49),
.A2(n_36),
.B1(n_44),
.B2(n_35),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_72),
.B(n_51),
.Y(n_87)
);

OAI21xp33_ASAP7_75t_SL g73 ( 
.A1(n_61),
.A2(n_32),
.B(n_38),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_73),
.A2(n_60),
.B1(n_28),
.B2(n_64),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_58),
.A2(n_14),
.B1(n_15),
.B2(n_12),
.Y(n_75)
);

HB1xp67_ASAP7_75t_L g76 ( 
.A(n_59),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_76),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_48),
.A2(n_44),
.B1(n_35),
.B2(n_13),
.Y(n_77)
);

NAND3xp33_ASAP7_75t_L g78 ( 
.A(n_52),
.B(n_32),
.C(n_14),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_78),
.B(n_28),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_62),
.A2(n_55),
.B1(n_57),
.B2(n_65),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_87),
.A2(n_105),
.B1(n_69),
.B2(n_75),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_82),
.B(n_53),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_88),
.B(n_89),
.Y(n_113)
);

INVx6_ASAP7_75t_L g90 ( 
.A(n_74),
.Y(n_90)
);

BUFx2_ASAP7_75t_L g128 ( 
.A(n_90),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_91),
.A2(n_84),
.B1(n_80),
.B2(n_68),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_83),
.B(n_51),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_92),
.B(n_93),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_82),
.B(n_50),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_83),
.B(n_79),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_95),
.B(n_97),
.Y(n_124)
);

CKINVDCx6p67_ASAP7_75t_R g96 ( 
.A(n_86),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_96),
.B(n_106),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_81),
.B(n_71),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_79),
.B(n_50),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_98),
.B(n_100),
.Y(n_127)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_68),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_99),
.B(n_74),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_71),
.B(n_50),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_70),
.B(n_51),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_101),
.B(n_28),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_L g102 ( 
.A1(n_73),
.A2(n_60),
.B1(n_59),
.B2(n_36),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_102),
.A2(n_74),
.B1(n_84),
.B2(n_80),
.Y(n_121)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_86),
.Y(n_103)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_103),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_76),
.Y(n_106)
);

XOR2xp5_ASAP7_75t_L g107 ( 
.A(n_92),
.B(n_85),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_107),
.B(n_119),
.C(n_129),
.Y(n_133)
);

AOI21xp5_ASAP7_75t_L g108 ( 
.A1(n_87),
.A2(n_67),
.B(n_72),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_SL g141 ( 
.A1(n_108),
.A2(n_121),
.B(n_126),
.Y(n_141)
);

CKINVDCx16_ASAP7_75t_R g109 ( 
.A(n_88),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_109),
.B(n_117),
.Y(n_151)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_110),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_114),
.A2(n_123),
.B1(n_125),
.B2(n_130),
.Y(n_135)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_103),
.Y(n_115)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_115),
.Y(n_136)
);

NOR2x1_ASAP7_75t_L g116 ( 
.A(n_89),
.B(n_78),
.Y(n_116)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_116),
.Y(n_143)
);

CKINVDCx16_ASAP7_75t_R g117 ( 
.A(n_97),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_103),
.Y(n_118)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_118),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_100),
.B(n_77),
.C(n_28),
.Y(n_119)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_94),
.Y(n_122)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_122),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_101),
.A2(n_37),
.B1(n_26),
.B2(n_20),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_L g129 ( 
.A(n_95),
.B(n_31),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_104),
.A2(n_26),
.B1(n_37),
.B2(n_34),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_122),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_131),
.B(n_134),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_124),
.B(n_104),
.Y(n_134)
);

OAI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_109),
.A2(n_102),
.B1(n_91),
.B2(n_93),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_137),
.A2(n_123),
.B1(n_116),
.B2(n_125),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_117),
.B(n_106),
.Y(n_138)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_138),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g139 ( 
.A(n_111),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_139),
.B(n_144),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_124),
.B(n_98),
.Y(n_140)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_140),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_107),
.B(n_94),
.C(n_40),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_142),
.B(n_150),
.C(n_112),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_129),
.B(n_96),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_127),
.B(n_90),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_145),
.B(n_147),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_114),
.A2(n_90),
.B1(n_99),
.B2(n_96),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_146),
.A2(n_121),
.B1(n_130),
.B2(n_108),
.Y(n_161)
);

INVx4_ASAP7_75t_L g147 ( 
.A(n_128),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_113),
.B(n_96),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g181 ( 
.A(n_148),
.B(n_155),
.Y(n_181)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_128),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_149),
.B(n_153),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_119),
.B(n_40),
.C(n_68),
.Y(n_150)
);

AOI21xp5_ASAP7_75t_L g152 ( 
.A1(n_111),
.A2(n_96),
.B(n_86),
.Y(n_152)
);

INVxp67_ASAP7_75t_L g162 ( 
.A(n_152),
.Y(n_162)
);

INVx4_ASAP7_75t_L g153 ( 
.A(n_128),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_113),
.B(n_64),
.Y(n_155)
);

NOR2xp67_ASAP7_75t_L g157 ( 
.A(n_116),
.B(n_120),
.Y(n_157)
);

NAND2xp67_ASAP7_75t_SL g179 ( 
.A(n_157),
.B(n_16),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g159 ( 
.A(n_133),
.B(n_120),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_159),
.B(n_168),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_160),
.A2(n_163),
.B1(n_172),
.B2(n_146),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_161),
.A2(n_132),
.B1(n_141),
.B2(n_143),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_134),
.A2(n_127),
.B1(n_126),
.B2(n_118),
.Y(n_163)
);

AOI21xp5_ASAP7_75t_L g164 ( 
.A1(n_151),
.A2(n_115),
.B(n_112),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_SL g205 ( 
.A1(n_164),
.A2(n_15),
.B(n_25),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_131),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_165),
.Y(n_194)
);

CKINVDCx16_ASAP7_75t_R g170 ( 
.A(n_151),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_170),
.B(n_176),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_SL g171 ( 
.A(n_157),
.B(n_31),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_SL g201 ( 
.A(n_171),
.B(n_179),
.C(n_184),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_135),
.A2(n_139),
.B1(n_143),
.B2(n_145),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_133),
.B(n_31),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_174),
.B(n_175),
.C(n_178),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g175 ( 
.A(n_142),
.B(n_31),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_156),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_140),
.B(n_34),
.Y(n_178)
);

INVxp67_ASAP7_75t_L g180 ( 
.A(n_152),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_180),
.B(n_182),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_135),
.A2(n_15),
.B1(n_21),
.B2(n_25),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g183 ( 
.A(n_141),
.B(n_34),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_183),
.B(n_168),
.C(n_174),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_SL g184 ( 
.A(n_150),
.B(n_22),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_165),
.Y(n_187)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_187),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_SL g188 ( 
.A(n_169),
.B(n_132),
.Y(n_188)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_188),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_167),
.B(n_156),
.Y(n_189)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_189),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_190),
.A2(n_203),
.B1(n_204),
.B2(n_206),
.Y(n_219)
);

CKINVDCx16_ASAP7_75t_R g191 ( 
.A(n_166),
.Y(n_191)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_191),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_192),
.A2(n_197),
.B1(n_20),
.B2(n_21),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_SL g193 ( 
.A(n_181),
.B(n_154),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_193),
.B(n_205),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_195),
.B(n_175),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_162),
.A2(n_154),
.B1(n_136),
.B2(n_147),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_177),
.Y(n_198)
);

AOI21xp5_ASAP7_75t_L g226 ( 
.A1(n_198),
.A2(n_199),
.B(n_202),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_173),
.B(n_136),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_159),
.B(n_149),
.C(n_153),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_200),
.B(n_184),
.C(n_178),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_158),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_172),
.A2(n_160),
.B1(n_163),
.B2(n_179),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_171),
.Y(n_204)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_183),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_208),
.B(n_218),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_210),
.B(n_213),
.C(n_214),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_195),
.B(n_180),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_212),
.B(n_216),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_200),
.B(n_162),
.C(n_56),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_207),
.B(n_56),
.C(n_54),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_207),
.B(n_54),
.C(n_26),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_215),
.B(n_220),
.C(n_225),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_185),
.B(n_17),
.C(n_26),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_217),
.A2(n_186),
.B1(n_222),
.B2(n_196),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_185),
.B(n_16),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_206),
.B(n_26),
.C(n_17),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_190),
.A2(n_9),
.B1(n_11),
.B2(n_10),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_224),
.A2(n_186),
.B1(n_189),
.B2(n_198),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_197),
.B(n_23),
.C(n_21),
.Y(n_225)
);

AO22x1_ASAP7_75t_SL g227 ( 
.A1(n_219),
.A2(n_194),
.B1(n_203),
.B2(n_192),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_227),
.B(n_233),
.Y(n_245)
);

A2O1A1O1Ixp25_ASAP7_75t_L g228 ( 
.A1(n_226),
.A2(n_201),
.B(n_204),
.C(n_194),
.D(n_199),
.Y(n_228)
);

HB1xp67_ASAP7_75t_L g247 ( 
.A(n_228),
.Y(n_247)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_211),
.Y(n_230)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_230),
.Y(n_251)
);

CKINVDCx16_ASAP7_75t_R g254 ( 
.A(n_231),
.Y(n_254)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_232),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_221),
.A2(n_201),
.B1(n_205),
.B2(n_23),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_SL g234 ( 
.A(n_209),
.B(n_18),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_234),
.B(n_237),
.Y(n_246)
);

AOI22xp33_ASAP7_75t_SL g236 ( 
.A1(n_223),
.A2(n_18),
.B1(n_23),
.B2(n_21),
.Y(n_236)
);

AOI22xp33_ASAP7_75t_SL g250 ( 
.A1(n_236),
.A2(n_6),
.B1(n_11),
.B2(n_9),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_225),
.A2(n_23),
.B1(n_20),
.B2(n_18),
.Y(n_237)
);

AOI21xp5_ASAP7_75t_L g239 ( 
.A1(n_213),
.A2(n_8),
.B(n_11),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_239),
.B(n_240),
.Y(n_248)
);

AO22x1_ASAP7_75t_L g240 ( 
.A1(n_220),
.A2(n_8),
.B1(n_11),
.B2(n_10),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_214),
.A2(n_18),
.B1(n_20),
.B2(n_8),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_242),
.B(n_6),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_227),
.A2(n_210),
.B1(n_218),
.B2(n_215),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_L g258 ( 
.A1(n_243),
.A2(n_250),
.B1(n_241),
.B2(n_236),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_235),
.B(n_208),
.C(n_24),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_244),
.B(n_238),
.C(n_24),
.Y(n_264)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_249),
.Y(n_256)
);

XNOR2x1_ASAP7_75t_L g253 ( 
.A(n_228),
.B(n_6),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_253),
.B(n_232),
.Y(n_257)
);

AOI21x1_ASAP7_75t_L g255 ( 
.A1(n_227),
.A2(n_5),
.B(n_9),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_255),
.B(n_240),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_SL g272 ( 
.A(n_257),
.B(n_258),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_254),
.B(n_229),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_259),
.B(n_260),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_245),
.B(n_241),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_261),
.B(n_262),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_251),
.B(n_235),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_246),
.B(n_238),
.Y(n_263)
);

AOI21xp5_ASAP7_75t_L g273 ( 
.A1(n_263),
.A2(n_266),
.B(n_267),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_264),
.B(n_265),
.C(n_22),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_244),
.B(n_24),
.C(n_22),
.Y(n_265)
);

OAI21xp5_ASAP7_75t_SL g266 ( 
.A1(n_247),
.A2(n_24),
.B(n_22),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_SL g267 ( 
.A(n_253),
.B(n_5),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_264),
.B(n_243),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_268),
.B(n_270),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_257),
.A2(n_252),
.B1(n_248),
.B2(n_265),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_256),
.B(n_250),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_271),
.B(n_275),
.Y(n_279)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_274),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_264),
.B(n_22),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_262),
.B(n_22),
.C(n_16),
.Y(n_277)
);

FAx1_ASAP7_75t_SL g282 ( 
.A(n_277),
.B(n_4),
.CI(n_7),
.CON(n_282),
.SN(n_282)
);

MAJx2_ASAP7_75t_L g281 ( 
.A(n_276),
.B(n_16),
.C(n_4),
.Y(n_281)
);

OAI21xp5_ASAP7_75t_L g284 ( 
.A1(n_281),
.A2(n_283),
.B(n_273),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_SL g285 ( 
.A(n_282),
.B(n_277),
.Y(n_285)
);

OAI321xp33_ASAP7_75t_L g283 ( 
.A1(n_269),
.A2(n_4),
.A3(n_7),
.B1(n_5),
.B2(n_9),
.C(n_3),
.Y(n_283)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_284),
.B(n_272),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_285),
.B(n_286),
.Y(n_288)
);

OAI21xp5_ASAP7_75t_SL g286 ( 
.A1(n_280),
.A2(n_272),
.B(n_274),
.Y(n_286)
);

AOI21xp5_ASAP7_75t_L g289 ( 
.A1(n_287),
.A2(n_288),
.B(n_278),
.Y(n_289)
);

NAND3xp33_ASAP7_75t_L g290 ( 
.A(n_289),
.B(n_279),
.C(n_7),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_290),
.B(n_279),
.C(n_1),
.Y(n_291)
);

A2O1A1O1Ixp25_ASAP7_75t_L g292 ( 
.A1(n_291),
.A2(n_0),
.B(n_1),
.C(n_2),
.D(n_3),
.Y(n_292)
);

AOI21xp5_ASAP7_75t_SL g293 ( 
.A1(n_292),
.A2(n_0),
.B(n_1),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_SL g294 ( 
.A(n_293),
.B(n_0),
.Y(n_294)
);

OAI21xp5_ASAP7_75t_L g295 ( 
.A1(n_294),
.A2(n_0),
.B(n_1),
.Y(n_295)
);


endmodule