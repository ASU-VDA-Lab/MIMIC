module fake_jpeg_10628_n_139 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_139);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_139;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

INVx1_ASAP7_75t_L g13 ( 
.A(n_0),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_4),
.Y(n_14)
);

INVx13_ASAP7_75t_L g15 ( 
.A(n_7),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_0),
.Y(n_17)
);

INVx8_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_6),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_8),
.Y(n_23)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_2),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_5),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_20),
.Y(n_28)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_28),
.Y(n_43)
);

BUFx12_ASAP7_75t_L g29 ( 
.A(n_20),
.Y(n_29)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_29),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_20),
.Y(n_30)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_30),
.Y(n_50)
);

BUFx8_ASAP7_75t_L g31 ( 
.A(n_22),
.Y(n_31)
);

INVx5_ASAP7_75t_L g51 ( 
.A(n_31),
.Y(n_51)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_22),
.Y(n_32)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_32),
.Y(n_38)
);

BUFx2_ASAP7_75t_L g33 ( 
.A(n_22),
.Y(n_33)
);

CKINVDCx16_ASAP7_75t_R g40 ( 
.A(n_33),
.Y(n_40)
);

INVx5_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_23),
.B(n_0),
.Y(n_35)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_35),
.Y(n_39)
);

AND2x2_ASAP7_75t_L g36 ( 
.A(n_15),
.B(n_1),
.Y(n_36)
);

AND2x2_ASAP7_75t_L g46 ( 
.A(n_36),
.B(n_16),
.Y(n_46)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_24),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_37),
.Y(n_49)
);

CKINVDCx16_ASAP7_75t_R g41 ( 
.A(n_36),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_41),
.B(n_16),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_32),
.A2(n_25),
.B1(n_24),
.B2(n_18),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_45),
.A2(n_21),
.B1(n_14),
.B2(n_13),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_46),
.B(n_48),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g47 ( 
.A1(n_34),
.A2(n_18),
.B1(n_25),
.B2(n_24),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_47),
.A2(n_17),
.B1(n_31),
.B2(n_20),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g48 ( 
.A(n_31),
.B(n_15),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_L g52 ( 
.A1(n_41),
.A2(n_25),
.B1(n_18),
.B2(n_26),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_52),
.A2(n_54),
.B1(n_55),
.B2(n_56),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g53 ( 
.A(n_39),
.B(n_46),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_53),
.B(n_57),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_46),
.A2(n_21),
.B1(n_14),
.B2(n_13),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_51),
.A2(n_27),
.B1(n_26),
.B2(n_19),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_48),
.Y(n_57)
);

OAI21xp5_ASAP7_75t_L g58 ( 
.A1(n_47),
.A2(n_27),
.B(n_19),
.Y(n_58)
);

CKINVDCx16_ASAP7_75t_R g82 ( 
.A(n_58),
.Y(n_82)
);

OR2x2_ASAP7_75t_L g70 ( 
.A(n_59),
.B(n_61),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_48),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_60),
.B(n_66),
.Y(n_72)
);

NAND2x1_ASAP7_75t_SL g61 ( 
.A(n_44),
.B(n_33),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_39),
.B(n_23),
.Y(n_62)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_62),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g64 ( 
.A(n_49),
.B(n_30),
.C(n_28),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_64),
.B(n_65),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_49),
.B(n_20),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_44),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_38),
.B(n_17),
.Y(n_67)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_67),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_68),
.Y(n_79)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_66),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_69),
.B(n_50),
.Y(n_89)
);

BUFx2_ASAP7_75t_L g75 ( 
.A(n_61),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_75),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_62),
.B(n_50),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_77),
.B(n_67),
.Y(n_86)
);

O2A1O1Ixp33_ASAP7_75t_SL g80 ( 
.A1(n_60),
.A2(n_38),
.B(n_40),
.C(n_29),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_80),
.A2(n_68),
.B1(n_57),
.B2(n_61),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_54),
.B(n_40),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_81),
.B(n_83),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_65),
.B(n_43),
.Y(n_83)
);

XNOR2xp5_ASAP7_75t_L g84 ( 
.A(n_74),
.B(n_63),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_84),
.B(n_93),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_85),
.A2(n_71),
.B1(n_79),
.B2(n_76),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_86),
.B(n_96),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_78),
.B(n_53),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_87),
.B(n_88),
.Y(n_102)
);

NAND3xp33_ASAP7_75t_L g88 ( 
.A(n_81),
.B(n_63),
.C(n_59),
.Y(n_88)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_89),
.Y(n_97)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_72),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_91),
.B(n_92),
.Y(n_104)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_83),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_74),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_L g94 ( 
.A1(n_82),
.A2(n_58),
.B(n_64),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_94),
.B(n_75),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_73),
.B(n_43),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_90),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_98),
.B(n_101),
.Y(n_111)
);

XNOR2xp5_ASAP7_75t_SL g113 ( 
.A(n_100),
.B(n_84),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_90),
.Y(n_101)
);

AOI221xp5_ASAP7_75t_L g110 ( 
.A1(n_103),
.A2(n_94),
.B1(n_80),
.B2(n_70),
.C(n_91),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_95),
.A2(n_79),
.B1(n_70),
.B2(n_80),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_105),
.A2(n_78),
.B1(n_69),
.B2(n_51),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_85),
.Y(n_106)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_106),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_104),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_108),
.B(n_109),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_98),
.B(n_92),
.Y(n_109)
);

AOI322xp5_ASAP7_75t_L g118 ( 
.A1(n_110),
.A2(n_116),
.A3(n_102),
.B1(n_105),
.B2(n_100),
.C1(n_97),
.C2(n_73),
.Y(n_118)
);

XOR2xp5_ASAP7_75t_L g117 ( 
.A(n_113),
.B(n_99),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_99),
.B(n_93),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_L g121 ( 
.A(n_114),
.B(n_115),
.Y(n_121)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_107),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_117),
.B(n_120),
.C(n_1),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_L g123 ( 
.A1(n_118),
.A2(n_122),
.B(n_115),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_113),
.B(n_97),
.C(n_42),
.Y(n_120)
);

MAJx2_ASAP7_75t_L g122 ( 
.A(n_114),
.B(n_42),
.C(n_29),
.Y(n_122)
);

AOI21xp5_ASAP7_75t_SL g128 ( 
.A1(n_123),
.A2(n_122),
.B(n_117),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_119),
.B(n_111),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_124),
.B(n_125),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_L g125 ( 
.A(n_120),
.B(n_109),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_121),
.A2(n_112),
.B1(n_12),
.B2(n_11),
.Y(n_126)
);

NAND4xp25_ASAP7_75t_L g131 ( 
.A(n_126),
.B(n_10),
.C(n_8),
.D(n_4),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_L g129 ( 
.A1(n_127),
.A2(n_12),
.B(n_10),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_L g133 ( 
.A(n_128),
.B(n_125),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_129),
.B(n_2),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_131),
.B(n_2),
.Y(n_134)
);

OR2x2_ASAP7_75t_L g136 ( 
.A(n_132),
.B(n_134),
.Y(n_136)
);

OAI321xp33_ASAP7_75t_L g135 ( 
.A1(n_133),
.A2(n_130),
.A3(n_127),
.B1(n_6),
.B2(n_5),
.C(n_3),
.Y(n_135)
);

AOI21xp5_ASAP7_75t_SL g137 ( 
.A1(n_135),
.A2(n_3),
.B(n_5),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_SL g138 ( 
.A1(n_137),
.A2(n_136),
.B(n_6),
.Y(n_138)
);

XOR2xp5_ASAP7_75t_L g139 ( 
.A(n_138),
.B(n_133),
.Y(n_139)
);


endmodule