module fake_jpeg_20089_n_320 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_320);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_320;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

INVx2_ASAP7_75t_R g17 ( 
.A(n_11),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_9),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

INVx13_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

CKINVDCx14_ASAP7_75t_R g24 ( 
.A(n_4),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_11),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

INVx11_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_2),
.Y(n_31)
);

BUFx10_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_3),
.Y(n_33)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_28),
.Y(n_34)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_28),
.Y(n_35)
);

INVx11_ASAP7_75t_L g65 ( 
.A(n_35),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_28),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_L g37 ( 
.A1(n_20),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_37),
.A2(n_33),
.B1(n_31),
.B2(n_18),
.Y(n_56)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_26),
.Y(n_38)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_38),
.Y(n_63)
);

INVx1_ASAP7_75t_SL g39 ( 
.A(n_17),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_39),
.B(n_42),
.Y(n_46)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_28),
.Y(n_41)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_41),
.Y(n_69)
);

CKINVDCx16_ASAP7_75t_R g42 ( 
.A(n_17),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_17),
.Y(n_43)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_43),
.Y(n_67)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_17),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_44),
.B(n_32),
.Y(n_60)
);

OR2x2_ASAP7_75t_SL g45 ( 
.A(n_39),
.B(n_17),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_45),
.B(n_47),
.Y(n_71)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

CKINVDCx14_ASAP7_75t_R g48 ( 
.A(n_42),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_48),
.B(n_49),
.Y(n_78)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

AND2x2_ASAP7_75t_SL g51 ( 
.A(n_39),
.B(n_30),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_51),
.B(n_70),
.Y(n_82)
);

OA22x2_ASAP7_75t_L g52 ( 
.A1(n_43),
.A2(n_21),
.B1(n_20),
.B2(n_29),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_52),
.A2(n_56),
.B1(n_66),
.B2(n_34),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_38),
.A2(n_29),
.B1(n_20),
.B2(n_23),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_55),
.A2(n_29),
.B1(n_34),
.B2(n_23),
.Y(n_73)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_57),
.Y(n_81)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_58),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_43),
.B(n_24),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_59),
.B(n_61),
.Y(n_86)
);

CKINVDCx14_ASAP7_75t_R g77 ( 
.A(n_60),
.Y(n_77)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_35),
.Y(n_61)
);

NAND2x1_ASAP7_75t_L g62 ( 
.A(n_43),
.B(n_32),
.Y(n_62)
);

A2O1A1Ixp33_ASAP7_75t_L g74 ( 
.A1(n_62),
.A2(n_44),
.B(n_35),
.C(n_36),
.Y(n_74)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_36),
.Y(n_64)
);

CKINVDCx16_ASAP7_75t_R g79 ( 
.A(n_64),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_34),
.A2(n_37),
.B1(n_38),
.B2(n_23),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g68 ( 
.A(n_43),
.B(n_32),
.Y(n_68)
);

CKINVDCx16_ASAP7_75t_R g90 ( 
.A(n_68),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_43),
.B(n_44),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_72),
.A2(n_73),
.B1(n_83),
.B2(n_69),
.Y(n_117)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_74),
.B(n_52),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_L g75 ( 
.A1(n_66),
.A2(n_23),
.B1(n_41),
.B2(n_36),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_75),
.A2(n_80),
.B1(n_85),
.B2(n_87),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_54),
.Y(n_76)
);

NAND2x1_ASAP7_75t_SL g97 ( 
.A(n_76),
.B(n_45),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_54),
.A2(n_41),
.B1(n_18),
.B2(n_16),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_67),
.A2(n_29),
.B1(n_22),
.B2(n_25),
.Y(n_83)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_53),
.Y(n_84)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_84),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_70),
.A2(n_41),
.B1(n_24),
.B2(n_22),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_57),
.A2(n_16),
.B1(n_22),
.B2(n_25),
.Y(n_87)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_53),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_88),
.B(n_94),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_62),
.B(n_44),
.C(n_35),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_89),
.B(n_68),
.C(n_51),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_58),
.A2(n_16),
.B1(n_25),
.B2(n_27),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_91),
.A2(n_93),
.B1(n_46),
.B2(n_67),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_62),
.A2(n_19),
.B1(n_27),
.B2(n_44),
.Y(n_93)
);

CKINVDCx16_ASAP7_75t_R g94 ( 
.A(n_52),
.Y(n_94)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_53),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_95),
.B(n_69),
.Y(n_119)
);

O2A1O1Ixp33_ASAP7_75t_L g125 ( 
.A1(n_97),
.A2(n_71),
.B(n_86),
.C(n_74),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_81),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_98),
.B(n_106),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_99),
.A2(n_117),
.B1(n_120),
.B2(n_77),
.Y(n_132)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_81),
.Y(n_100)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_100),
.Y(n_129)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_92),
.Y(n_101)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_101),
.Y(n_135)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_79),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_102),
.B(n_107),
.Y(n_124)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_92),
.Y(n_103)
);

INVx1_ASAP7_75t_SL g134 ( 
.A(n_103),
.Y(n_134)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_80),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_105),
.B(n_111),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_87),
.Y(n_106)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_79),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_L g140 ( 
.A1(n_108),
.A2(n_89),
.B(n_74),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g136 ( 
.A(n_109),
.B(n_114),
.Y(n_136)
);

CKINVDCx16_ASAP7_75t_R g110 ( 
.A(n_78),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_110),
.B(n_63),
.Y(n_137)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_78),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_91),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_112),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_82),
.B(n_51),
.C(n_60),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_76),
.B(n_46),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_115),
.B(n_118),
.Y(n_144)
);

OAI21xp33_ASAP7_75t_L g116 ( 
.A1(n_82),
.A2(n_68),
.B(n_44),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_116),
.Y(n_142)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_85),
.Y(n_118)
);

CKINVDCx14_ASAP7_75t_R g148 ( 
.A(n_119),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_72),
.A2(n_64),
.B1(n_56),
.B2(n_52),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_71),
.B(n_47),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_121),
.B(n_99),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_86),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_122),
.B(n_77),
.Y(n_131)
);

NOR2x1_ASAP7_75t_L g123 ( 
.A(n_97),
.B(n_93),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_L g166 ( 
.A1(n_123),
.A2(n_125),
.B(n_140),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_118),
.A2(n_72),
.B1(n_94),
.B2(n_90),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_126),
.A2(n_138),
.B1(n_108),
.B2(n_113),
.Y(n_150)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_104),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_127),
.B(n_104),
.Y(n_162)
);

CKINVDCx14_ASAP7_75t_R g174 ( 
.A(n_131),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_132),
.A2(n_143),
.B1(n_147),
.B2(n_26),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_137),
.B(n_141),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_105),
.A2(n_90),
.B1(n_75),
.B2(n_73),
.Y(n_138)
);

OR2x2_ASAP7_75t_L g139 ( 
.A(n_122),
.B(n_89),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_139),
.B(n_146),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_111),
.B(n_63),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_120),
.A2(n_95),
.B1(n_88),
.B2(n_84),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_102),
.B(n_107),
.Y(n_145)
);

CKINVDCx16_ASAP7_75t_R g160 ( 
.A(n_145),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_108),
.A2(n_83),
.B1(n_49),
.B2(n_61),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g149 ( 
.A(n_109),
.B(n_30),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_149),
.B(n_26),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_150),
.A2(n_157),
.B1(n_170),
.B2(n_143),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g151 ( 
.A(n_136),
.B(n_114),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_151),
.B(n_153),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_SL g153 ( 
.A(n_123),
.B(n_97),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_144),
.B(n_98),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_154),
.B(n_168),
.Y(n_178)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_124),
.Y(n_155)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_155),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_132),
.A2(n_112),
.B1(n_106),
.B2(n_96),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_156),
.A2(n_175),
.B1(n_133),
.B2(n_146),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_126),
.A2(n_96),
.B1(n_115),
.B2(n_121),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_136),
.B(n_103),
.C(n_101),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_158),
.B(n_139),
.C(n_123),
.Y(n_186)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_129),
.Y(n_159)
);

CKINVDCx16_ASAP7_75t_R g190 ( 
.A(n_159),
.Y(n_190)
);

AO32x1_ASAP7_75t_L g161 ( 
.A1(n_131),
.A2(n_100),
.A3(n_26),
.B1(n_30),
.B2(n_21),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_SL g201 ( 
.A(n_161),
.B(n_33),
.Y(n_201)
);

CKINVDCx14_ASAP7_75t_R g193 ( 
.A(n_162),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_149),
.B(n_30),
.Y(n_163)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_163),
.B(n_32),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_129),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_164),
.B(n_165),
.Y(n_179)
);

CKINVDCx16_ASAP7_75t_R g165 ( 
.A(n_135),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_144),
.B(n_32),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_128),
.B(n_32),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_169),
.B(n_173),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_138),
.A2(n_50),
.B1(n_65),
.B2(n_27),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_171),
.B(n_147),
.Y(n_177)
);

AOI21xp5_ASAP7_75t_L g172 ( 
.A1(n_140),
.A2(n_0),
.B(n_1),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_SL g187 ( 
.A1(n_172),
.A2(n_125),
.B(n_142),
.Y(n_187)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_127),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_SL g175 ( 
.A1(n_133),
.A2(n_50),
.B1(n_65),
.B2(n_19),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_176),
.B(n_0),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_177),
.B(n_186),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_SL g180 ( 
.A(n_174),
.B(n_128),
.Y(n_180)
);

CKINVDCx14_ASAP7_75t_R g207 ( 
.A(n_180),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_181),
.A2(n_182),
.B1(n_188),
.B2(n_189),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_SL g183 ( 
.A(n_167),
.B(n_148),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_SL g209 ( 
.A(n_183),
.B(n_185),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_SL g185 ( 
.A(n_154),
.B(n_130),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_SL g211 ( 
.A1(n_187),
.A2(n_201),
.B(n_161),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_157),
.A2(n_139),
.B1(n_142),
.B2(n_135),
.Y(n_188)
);

OAI22xp33_ASAP7_75t_SL g189 ( 
.A1(n_155),
.A2(n_134),
.B1(n_19),
.B2(n_31),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_150),
.A2(n_152),
.B1(n_166),
.B2(n_170),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_191),
.A2(n_8),
.B1(n_14),
.B2(n_13),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_SL g192 ( 
.A(n_152),
.B(n_134),
.Y(n_192)
);

AOI21xp33_ASAP7_75t_L g219 ( 
.A1(n_192),
.A2(n_163),
.B(n_171),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_194),
.B(n_195),
.Y(n_225)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_173),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_151),
.B(n_21),
.Y(n_196)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_196),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_172),
.A2(n_31),
.B1(n_33),
.B2(n_21),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_197),
.A2(n_200),
.B1(n_169),
.B2(n_159),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_166),
.B(n_32),
.Y(n_198)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_198),
.Y(n_213)
);

AOI21xp5_ASAP7_75t_L g204 ( 
.A1(n_187),
.A2(n_153),
.B(n_160),
.Y(n_204)
);

INVxp67_ASAP7_75t_L g242 ( 
.A(n_204),
.Y(n_242)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_179),
.Y(n_205)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_205),
.Y(n_229)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_195),
.Y(n_206)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_206),
.Y(n_234)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_202),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_208),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_178),
.A2(n_176),
.B1(n_168),
.B2(n_158),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_210),
.A2(n_212),
.B1(n_223),
.B2(n_15),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_211),
.B(n_214),
.Y(n_240)
);

INVxp67_ASAP7_75t_L g214 ( 
.A(n_199),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_202),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_215),
.Y(n_235)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_185),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_216),
.Y(n_243)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_192),
.Y(n_217)
);

CKINVDCx16_ASAP7_75t_R g239 ( 
.A(n_217),
.Y(n_239)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_180),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_218),
.B(n_188),
.Y(n_227)
);

AO22x1_ASAP7_75t_L g244 ( 
.A1(n_219),
.A2(n_222),
.B1(n_226),
.B2(n_2),
.Y(n_244)
);

AND2x2_ASAP7_75t_L g222 ( 
.A(n_193),
.B(n_1),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_178),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_224),
.B(n_191),
.C(n_190),
.Y(n_228)
);

AND2x2_ASAP7_75t_L g226 ( 
.A(n_186),
.B(n_1),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_SL g257 ( 
.A(n_227),
.B(n_209),
.Y(n_257)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_228),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_220),
.B(n_184),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_230),
.B(n_233),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_220),
.B(n_184),
.C(n_196),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_231),
.B(n_241),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_204),
.B(n_177),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_SL g236 ( 
.A(n_210),
.B(n_198),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_236),
.B(n_237),
.C(n_238),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_SL g237 ( 
.A(n_225),
.B(n_194),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_225),
.B(n_182),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_213),
.B(n_201),
.C(n_9),
.Y(n_241)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_244),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_245),
.B(n_246),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_221),
.B(n_8),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_213),
.B(n_8),
.C(n_4),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_247),
.B(n_207),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_229),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_250),
.B(n_254),
.Y(n_268)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_234),
.Y(n_252)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_252),
.Y(n_276)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_238),
.Y(n_254)
);

INVxp67_ASAP7_75t_L g255 ( 
.A(n_240),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_255),
.B(n_259),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_256),
.B(n_257),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_242),
.A2(n_203),
.B1(n_221),
.B2(n_226),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_242),
.A2(n_223),
.B1(n_203),
.B2(n_214),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_260),
.B(n_263),
.Y(n_271)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_246),
.Y(n_262)
);

CKINVDCx16_ASAP7_75t_R g279 ( 
.A(n_262),
.Y(n_279)
);

INVxp67_ASAP7_75t_SL g263 ( 
.A(n_243),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_241),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_264),
.B(n_244),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_SL g265 ( 
.A(n_249),
.B(n_248),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_265),
.B(n_269),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_253),
.B(n_230),
.C(n_236),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_SL g286 ( 
.A(n_266),
.B(n_277),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_253),
.B(n_233),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_267),
.B(n_275),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_SL g269 ( 
.A(n_262),
.B(n_247),
.Y(n_269)
);

AOI21xp5_ASAP7_75t_L g270 ( 
.A1(n_255),
.A2(n_239),
.B(n_235),
.Y(n_270)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_270),
.Y(n_280)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_273),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_259),
.B(n_237),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_258),
.B(n_226),
.C(n_232),
.Y(n_277)
);

MAJx2_ASAP7_75t_L g278 ( 
.A(n_258),
.B(n_211),
.C(n_222),
.Y(n_278)
);

OAI21xp5_ASAP7_75t_L g287 ( 
.A1(n_278),
.A2(n_261),
.B(n_251),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_276),
.B(n_252),
.Y(n_281)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_281),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_271),
.B(n_206),
.Y(n_284)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_284),
.Y(n_301)
);

XOR2xp5_ASAP7_75t_L g296 ( 
.A(n_287),
.B(n_286),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_272),
.B(n_254),
.C(n_260),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_288),
.B(n_289),
.Y(n_300)
);

AND2x2_ASAP7_75t_L g289 ( 
.A(n_277),
.B(n_275),
.Y(n_289)
);

AOI21xp5_ASAP7_75t_L g290 ( 
.A1(n_268),
.A2(n_222),
.B(n_5),
.Y(n_290)
);

OAI21xp5_ASAP7_75t_L g293 ( 
.A1(n_290),
.A2(n_278),
.B(n_279),
.Y(n_293)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_274),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_291),
.B(n_284),
.Y(n_292)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_292),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_293),
.B(n_294),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_285),
.B(n_267),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_SL g306 ( 
.A(n_296),
.B(n_7),
.Y(n_306)
);

OAI21xp5_ASAP7_75t_L g297 ( 
.A1(n_289),
.A2(n_266),
.B(n_5),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_297),
.B(n_299),
.Y(n_304)
);

AOI21xp33_ASAP7_75t_L g298 ( 
.A1(n_280),
.A2(n_12),
.B(n_6),
.Y(n_298)
);

AND2x2_ASAP7_75t_L g308 ( 
.A(n_298),
.B(n_10),
.Y(n_308)
);

AND2x2_ASAP7_75t_SL g299 ( 
.A(n_282),
.B(n_7),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_295),
.B(n_281),
.Y(n_302)
);

AOI21xp33_ASAP7_75t_L g311 ( 
.A1(n_302),
.A2(n_305),
.B(n_306),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_292),
.B(n_283),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_301),
.B(n_7),
.Y(n_307)
);

HB1xp67_ASAP7_75t_L g312 ( 
.A(n_307),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_308),
.B(n_10),
.C(n_12),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_303),
.B(n_300),
.C(n_299),
.Y(n_310)
);

CKINVDCx14_ASAP7_75t_R g316 ( 
.A(n_310),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_309),
.B(n_304),
.C(n_10),
.Y(n_313)
);

AOI21xp5_ASAP7_75t_L g315 ( 
.A1(n_313),
.A2(n_314),
.B(n_12),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_315),
.A2(n_312),
.B1(n_13),
.B2(n_14),
.Y(n_317)
);

OAI21xp5_ASAP7_75t_SL g318 ( 
.A1(n_317),
.A2(n_311),
.B(n_316),
.Y(n_318)
);

AO21x1_ASAP7_75t_L g319 ( 
.A1(n_318),
.A2(n_15),
.B(n_3),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_319),
.B(n_15),
.Y(n_320)
);


endmodule