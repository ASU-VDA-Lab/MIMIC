module fake_ariane_264_n_754 (n_83, n_8, n_56, n_60, n_64, n_119, n_124, n_90, n_38, n_47, n_110, n_18, n_86, n_75, n_89, n_67, n_34, n_69, n_95, n_92, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_120, n_106, n_12, n_53, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_49, n_20, n_100, n_17, n_50, n_132, n_62, n_51, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_85, n_130, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_11, n_129, n_126, n_137, n_122, n_52, n_135, n_73, n_77, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_136, n_28, n_80, n_97, n_14, n_88, n_68, n_116, n_104, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_127, n_35, n_54, n_25, n_754);

input n_83;
input n_8;
input n_56;
input n_60;
input n_64;
input n_119;
input n_124;
input n_90;
input n_38;
input n_47;
input n_110;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_34;
input n_69;
input n_95;
input n_92;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_120;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_51;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_85;
input n_130;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_52;
input n_135;
input n_73;
input n_77;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_136;
input n_28;
input n_80;
input n_97;
input n_14;
input n_88;
input n_68;
input n_116;
input n_104;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_127;
input n_35;
input n_54;
input n_25;

output n_754;

wire n_295;
wire n_356;
wire n_556;
wire n_170;
wire n_190;
wire n_698;
wire n_695;
wire n_160;
wire n_180;
wire n_730;
wire n_386;
wire n_307;
wire n_516;
wire n_589;
wire n_332;
wire n_581;
wire n_294;
wire n_646;
wire n_197;
wire n_640;
wire n_463;
wire n_176;
wire n_691;
wire n_404;
wire n_172;
wire n_678;
wire n_651;
wire n_347;
wire n_423;
wire n_183;
wire n_469;
wire n_479;
wire n_726;
wire n_603;
wire n_373;
wire n_299;
wire n_541;
wire n_499;
wire n_564;
wire n_610;
wire n_205;
wire n_752;
wire n_341;
wire n_245;
wire n_421;
wire n_549;
wire n_522;
wire n_319;
wire n_591;
wire n_690;
wire n_416;
wire n_283;
wire n_187;
wire n_525;
wire n_367;
wire n_713;
wire n_649;
wire n_598;
wire n_345;
wire n_374;
wire n_318;
wire n_244;
wire n_643;
wire n_679;
wire n_226;
wire n_220;
wire n_261;
wire n_682;
wire n_663;
wire n_370;
wire n_706;
wire n_189;
wire n_717;
wire n_286;
wire n_443;
wire n_586;
wire n_686;
wire n_605;
wire n_424;
wire n_528;
wire n_584;
wire n_387;
wire n_406;
wire n_524;
wire n_391;
wire n_349;
wire n_634;
wire n_466;
wire n_346;
wire n_214;
wire n_552;
wire n_348;
wire n_462;
wire n_607;
wire n_670;
wire n_410;
wire n_445;
wire n_515;
wire n_379;
wire n_162;
wire n_264;
wire n_737;
wire n_198;
wire n_232;
wire n_441;
wire n_568;
wire n_385;
wire n_637;
wire n_327;
wire n_372;
wire n_377;
wire n_396;
wire n_631;
wire n_399;
wire n_554;
wire n_520;
wire n_714;
wire n_279;
wire n_702;
wire n_207;
wire n_363;
wire n_720;
wire n_354;
wire n_725;
wire n_419;
wire n_151;
wire n_146;
wire n_230;
wire n_270;
wire n_194;
wire n_633;
wire n_154;
wire n_338;
wire n_142;
wire n_285;
wire n_473;
wire n_186;
wire n_202;
wire n_145;
wire n_193;
wire n_733;
wire n_500;
wire n_665;
wire n_336;
wire n_731;
wire n_315;
wire n_594;
wire n_311;
wire n_239;
wire n_402;
wire n_272;
wire n_668;
wire n_339;
wire n_738;
wire n_672;
wire n_487;
wire n_740;
wire n_167;
wire n_422;
wire n_153;
wire n_648;
wire n_269;
wire n_597;
wire n_158;
wire n_259;
wire n_553;
wire n_446;
wire n_143;
wire n_753;
wire n_566;
wire n_578;
wire n_701;
wire n_625;
wire n_152;
wire n_557;
wire n_405;
wire n_169;
wire n_173;
wire n_242;
wire n_645;
wire n_331;
wire n_320;
wire n_309;
wire n_559;
wire n_485;
wire n_401;
wire n_267;
wire n_495;
wire n_504;
wire n_647;
wire n_483;
wire n_335;
wire n_435;
wire n_350;
wire n_291;
wire n_344;
wire n_381;
wire n_426;
wire n_433;
wire n_481;
wire n_600;
wire n_721;
wire n_398;
wire n_210;
wire n_200;
wire n_529;
wire n_502;
wire n_166;
wire n_253;
wire n_561;
wire n_218;
wire n_271;
wire n_465;
wire n_507;
wire n_486;
wire n_247;
wire n_569;
wire n_567;
wire n_732;
wire n_240;
wire n_369;
wire n_224;
wire n_547;
wire n_420;
wire n_562;
wire n_518;
wire n_439;
wire n_604;
wire n_614;
wire n_677;
wire n_222;
wire n_478;
wire n_703;
wire n_748;
wire n_510;
wire n_256;
wire n_326;
wire n_681;
wire n_227;
wire n_188;
wire n_323;
wire n_550;
wire n_635;
wire n_707;
wire n_330;
wire n_400;
wire n_689;
wire n_694;
wire n_282;
wire n_328;
wire n_368;
wire n_590;
wire n_699;
wire n_727;
wire n_277;
wire n_248;
wire n_301;
wire n_467;
wire n_432;
wire n_545;
wire n_536;
wire n_644;
wire n_293;
wire n_620;
wire n_228;
wire n_325;
wire n_276;
wire n_688;
wire n_636;
wire n_427;
wire n_587;
wire n_497;
wire n_693;
wire n_303;
wire n_671;
wire n_442;
wire n_168;
wire n_206;
wire n_352;
wire n_538;
wire n_576;
wire n_511;
wire n_611;
wire n_238;
wire n_455;
wire n_429;
wire n_365;
wire n_654;
wire n_588;
wire n_638;
wire n_334;
wire n_192;
wire n_729;
wire n_661;
wire n_488;
wire n_667;
wire n_300;
wire n_533;
wire n_505;
wire n_163;
wire n_141;
wire n_390;
wire n_498;
wire n_501;
wire n_438;
wire n_314;
wire n_684;
wire n_440;
wire n_627;
wire n_273;
wire n_305;
wire n_539;
wire n_312;
wire n_233;
wire n_728;
wire n_388;
wire n_333;
wire n_449;
wire n_612;
wire n_413;
wire n_392;
wire n_376;
wire n_512;
wire n_715;
wire n_579;
wire n_459;
wire n_685;
wire n_221;
wire n_321;
wire n_458;
wire n_361;
wire n_149;
wire n_383;
wire n_623;
wire n_237;
wire n_175;
wire n_711;
wire n_453;
wire n_734;
wire n_491;
wire n_181;
wire n_723;
wire n_617;
wire n_616;
wire n_658;
wire n_630;
wire n_705;
wire n_570;
wire n_260;
wire n_362;
wire n_543;
wire n_310;
wire n_709;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_281;
wire n_628;
wire n_461;
wire n_209;
wire n_262;
wire n_490;
wire n_743;
wire n_225;
wire n_235;
wire n_660;
wire n_464;
wire n_735;
wire n_575;
wire n_546;
wire n_297;
wire n_662;
wire n_641;
wire n_503;
wire n_700;
wire n_290;
wire n_527;
wire n_741;
wire n_747;
wire n_371;
wire n_199;
wire n_639;
wire n_217;
wire n_452;
wire n_673;
wire n_676;
wire n_178;
wire n_551;
wire n_308;
wire n_708;
wire n_417;
wire n_201;
wire n_572;
wire n_343;
wire n_414;
wire n_571;
wire n_680;
wire n_287;
wire n_302;
wire n_380;
wire n_582;
wire n_284;
wire n_448;
wire n_593;
wire n_710;
wire n_249;
wire n_534;
wire n_212;
wire n_444;
wire n_355;
wire n_609;
wire n_278;
wire n_255;
wire n_560;
wire n_450;
wire n_257;
wire n_148;
wire n_652;
wire n_451;
wire n_613;
wire n_745;
wire n_475;
wire n_409;
wire n_171;
wire n_519;
wire n_384;
wire n_468;
wire n_526;
wire n_716;
wire n_742;
wire n_182;
wire n_696;
wire n_674;
wire n_482;
wire n_316;
wire n_196;
wire n_577;
wire n_407;
wire n_254;
wire n_596;
wire n_476;
wire n_460;
wire n_219;
wire n_535;
wire n_231;
wire n_366;
wire n_744;
wire n_656;
wire n_555;
wire n_234;
wire n_492;
wire n_574;
wire n_280;
wire n_215;
wire n_252;
wire n_629;
wire n_664;
wire n_161;
wire n_454;
wire n_298;
wire n_532;
wire n_415;
wire n_655;
wire n_540;
wire n_216;
wire n_544;
wire n_692;
wire n_599;
wire n_514;
wire n_418;
wire n_537;
wire n_223;
wire n_403;
wire n_750;
wire n_389;
wire n_657;
wire n_513;
wire n_288;
wire n_179;
wire n_395;
wire n_621;
wire n_195;
wire n_606;
wire n_213;
wire n_304;
wire n_659;
wire n_509;
wire n_583;
wire n_724;
wire n_306;
wire n_666;
wire n_313;
wire n_430;
wire n_626;
wire n_493;
wire n_722;
wire n_203;
wire n_378;
wire n_436;
wire n_150;
wire n_375;
wire n_324;
wire n_585;
wire n_669;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_622;
wire n_697;
wire n_472;
wire n_296;
wire n_265;
wire n_746;
wire n_208;
wire n_456;
wire n_156;
wire n_292;
wire n_174;
wire n_275;
wire n_704;
wire n_147;
wire n_204;
wire n_751;
wire n_615;
wire n_521;
wire n_496;
wire n_739;
wire n_342;
wire n_246;
wire n_517;
wire n_530;
wire n_428;
wire n_159;
wire n_358;
wire n_580;
wire n_608;
wire n_494;
wire n_719;
wire n_263;
wire n_434;
wire n_360;
wire n_563;
wire n_229;
wire n_394;
wire n_250;
wire n_165;
wire n_144;
wire n_317;
wire n_243;
wire n_329;
wire n_718;
wire n_185;
wire n_340;
wire n_749;
wire n_289;
wire n_548;
wire n_542;
wire n_523;
wire n_268;
wire n_266;
wire n_470;
wire n_457;
wire n_164;
wire n_157;
wire n_632;
wire n_184;
wire n_177;
wire n_477;
wire n_364;
wire n_258;
wire n_650;
wire n_425;
wire n_431;
wire n_508;
wire n_624;
wire n_618;
wire n_484;
wire n_411;
wire n_712;
wire n_353;
wire n_736;
wire n_241;
wire n_357;
wire n_412;
wire n_687;
wire n_447;
wire n_191;
wire n_382;
wire n_489;
wire n_480;
wire n_211;
wire n_642;
wire n_408;
wire n_595;
wire n_322;
wire n_251;
wire n_506;
wire n_602;
wire n_558;
wire n_592;
wire n_397;
wire n_471;
wire n_351;
wire n_393;
wire n_474;
wire n_653;
wire n_359;
wire n_155;
wire n_573;
wire n_531;
wire n_675;

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_63),
.Y(n_141)
);

CKINVDCx5p33_ASAP7_75t_R g142 ( 
.A(n_0),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_131),
.Y(n_143)
);

CKINVDCx5p33_ASAP7_75t_R g144 ( 
.A(n_105),
.Y(n_144)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_28),
.Y(n_145)
);

CKINVDCx5p33_ASAP7_75t_R g146 ( 
.A(n_23),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_99),
.Y(n_147)
);

CKINVDCx5p33_ASAP7_75t_R g148 ( 
.A(n_7),
.Y(n_148)
);

CKINVDCx5p33_ASAP7_75t_R g149 ( 
.A(n_75),
.Y(n_149)
);

CKINVDCx5p33_ASAP7_75t_R g150 ( 
.A(n_9),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_70),
.Y(n_151)
);

INVx1_ASAP7_75t_SL g152 ( 
.A(n_133),
.Y(n_152)
);

CKINVDCx5p33_ASAP7_75t_R g153 ( 
.A(n_64),
.Y(n_153)
);

INVx2_ASAP7_75t_SL g154 ( 
.A(n_67),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_59),
.Y(n_155)
);

CKINVDCx5p33_ASAP7_75t_R g156 ( 
.A(n_114),
.Y(n_156)
);

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_17),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_41),
.Y(n_158)
);

CKINVDCx5p33_ASAP7_75t_R g159 ( 
.A(n_68),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_134),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_121),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_79),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_107),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_60),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_117),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_101),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_9),
.Y(n_167)
);

INVx1_ASAP7_75t_SL g168 ( 
.A(n_26),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_0),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_73),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_71),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_10),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_84),
.Y(n_173)
);

BUFx10_ASAP7_75t_L g174 ( 
.A(n_98),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_77),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_36),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_11),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_5),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g179 ( 
.A(n_116),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_132),
.Y(n_180)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_5),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_13),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_85),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_109),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_128),
.Y(n_185)
);

CKINVDCx16_ASAP7_75t_R g186 ( 
.A(n_136),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_37),
.Y(n_187)
);

INVx2_ASAP7_75t_SL g188 ( 
.A(n_53),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_135),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_139),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_21),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_126),
.Y(n_192)
);

BUFx6f_ASAP7_75t_L g193 ( 
.A(n_51),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_137),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_143),
.B(n_1),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_147),
.B(n_1),
.Y(n_196)
);

BUFx2_ASAP7_75t_L g197 ( 
.A(n_142),
.Y(n_197)
);

BUFx6f_ASAP7_75t_L g198 ( 
.A(n_179),
.Y(n_198)
);

BUFx6f_ASAP7_75t_L g199 ( 
.A(n_179),
.Y(n_199)
);

BUFx12f_ASAP7_75t_L g200 ( 
.A(n_174),
.Y(n_200)
);

BUFx6f_ASAP7_75t_L g201 ( 
.A(n_179),
.Y(n_201)
);

INVx5_ASAP7_75t_L g202 ( 
.A(n_179),
.Y(n_202)
);

AND2x2_ASAP7_75t_L g203 ( 
.A(n_181),
.B(n_2),
.Y(n_203)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_151),
.Y(n_204)
);

BUFx12f_ASAP7_75t_L g205 ( 
.A(n_174),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_167),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_155),
.B(n_2),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_169),
.Y(n_208)
);

INVx3_ASAP7_75t_L g209 ( 
.A(n_181),
.Y(n_209)
);

CKINVDCx11_ASAP7_75t_R g210 ( 
.A(n_141),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_160),
.B(n_3),
.Y(n_211)
);

BUFx6f_ASAP7_75t_L g212 ( 
.A(n_193),
.Y(n_212)
);

BUFx6f_ASAP7_75t_L g213 ( 
.A(n_193),
.Y(n_213)
);

AND2x6_ASAP7_75t_L g214 ( 
.A(n_145),
.B(n_24),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_SL g215 ( 
.A(n_186),
.B(n_25),
.Y(n_215)
);

BUFx12f_ASAP7_75t_L g216 ( 
.A(n_174),
.Y(n_216)
);

AND2x6_ASAP7_75t_L g217 ( 
.A(n_145),
.B(n_27),
.Y(n_217)
);

INVx5_ASAP7_75t_L g218 ( 
.A(n_193),
.Y(n_218)
);

INVx4_ASAP7_75t_L g219 ( 
.A(n_193),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_162),
.B(n_3),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_163),
.B(n_4),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_141),
.Y(n_222)
);

AND2x4_ASAP7_75t_L g223 ( 
.A(n_154),
.B(n_4),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_165),
.B(n_6),
.Y(n_224)
);

BUFx2_ASAP7_75t_L g225 ( 
.A(n_146),
.Y(n_225)
);

AND2x2_ASAP7_75t_L g226 ( 
.A(n_188),
.B(n_6),
.Y(n_226)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_171),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_176),
.B(n_184),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_148),
.B(n_7),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_144),
.B(n_8),
.Y(n_230)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_149),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_153),
.B(n_8),
.Y(n_232)
);

XNOR2x1_ASAP7_75t_L g233 ( 
.A(n_150),
.B(n_157),
.Y(n_233)
);

INVx5_ASAP7_75t_L g234 ( 
.A(n_156),
.Y(n_234)
);

OAI22xp33_ASAP7_75t_SL g235 ( 
.A1(n_215),
.A2(n_177),
.B1(n_172),
.B2(n_191),
.Y(n_235)
);

OAI22xp33_ASAP7_75t_L g236 ( 
.A1(n_200),
.A2(n_216),
.B1(n_205),
.B2(n_194),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_233),
.A2(n_194),
.B1(n_170),
.B2(n_192),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_206),
.Y(n_238)
);

OAI22xp33_ASAP7_75t_L g239 ( 
.A1(n_200),
.A2(n_170),
.B1(n_185),
.B2(n_178),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_233),
.A2(n_182),
.B1(n_152),
.B2(n_168),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_208),
.Y(n_241)
);

INVx3_ASAP7_75t_L g242 ( 
.A(n_219),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_204),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_204),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_223),
.A2(n_190),
.B1(n_189),
.B2(n_187),
.Y(n_245)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_219),
.Y(n_246)
);

OAI22xp33_ASAP7_75t_SL g247 ( 
.A1(n_229),
.A2(n_183),
.B1(n_180),
.B2(n_175),
.Y(n_247)
);

BUFx6f_ASAP7_75t_L g248 ( 
.A(n_198),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_223),
.A2(n_173),
.B1(n_166),
.B2(n_164),
.Y(n_249)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_219),
.Y(n_250)
);

OAI22xp33_ASAP7_75t_SL g251 ( 
.A1(n_228),
.A2(n_161),
.B1(n_159),
.B2(n_158),
.Y(n_251)
);

INVxp67_ASAP7_75t_SL g252 ( 
.A(n_227),
.Y(n_252)
);

OAI22xp33_ASAP7_75t_L g253 ( 
.A1(n_205),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_253)
);

OAI22xp33_ASAP7_75t_L g254 ( 
.A1(n_216),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_254)
);

OR2x2_ASAP7_75t_L g255 ( 
.A(n_197),
.B(n_14),
.Y(n_255)
);

AND2x2_ASAP7_75t_L g256 ( 
.A(n_225),
.B(n_15),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_231),
.B(n_15),
.Y(n_257)
);

OAI22xp33_ASAP7_75t_L g258 ( 
.A1(n_222),
.A2(n_195),
.B1(n_196),
.B2(n_220),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_223),
.A2(n_16),
.B1(n_17),
.B2(n_18),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_226),
.A2(n_16),
.B1(n_18),
.B2(n_19),
.Y(n_260)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_198),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_227),
.Y(n_262)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_198),
.Y(n_263)
);

OAI22xp33_ASAP7_75t_L g264 ( 
.A1(n_222),
.A2(n_221),
.B1(n_224),
.B2(n_203),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_L g265 ( 
.A1(n_226),
.A2(n_19),
.B1(n_20),
.B2(n_21),
.Y(n_265)
);

NAND3x1_ASAP7_75t_L g266 ( 
.A(n_203),
.B(n_20),
.C(n_22),
.Y(n_266)
);

OAI22xp33_ASAP7_75t_L g267 ( 
.A1(n_230),
.A2(n_22),
.B1(n_23),
.B2(n_29),
.Y(n_267)
);

OAI22xp33_ASAP7_75t_L g268 ( 
.A1(n_232),
.A2(n_30),
.B1(n_31),
.B2(n_32),
.Y(n_268)
);

AND2x4_ASAP7_75t_L g269 ( 
.A(n_231),
.B(n_33),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_207),
.A2(n_34),
.B1(n_35),
.B2(n_38),
.Y(n_270)
);

AND2x2_ASAP7_75t_L g271 ( 
.A(n_209),
.B(n_202),
.Y(n_271)
);

BUFx2_ASAP7_75t_L g272 ( 
.A(n_209),
.Y(n_272)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_198),
.Y(n_273)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_198),
.Y(n_274)
);

OAI22xp33_ASAP7_75t_SL g275 ( 
.A1(n_211),
.A2(n_39),
.B1(n_40),
.B2(n_42),
.Y(n_275)
);

OA22x2_ASAP7_75t_L g276 ( 
.A1(n_209),
.A2(n_43),
.B1(n_44),
.B2(n_45),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_210),
.A2(n_46),
.B1(n_47),
.B2(n_48),
.Y(n_277)
);

AO22x2_ASAP7_75t_L g278 ( 
.A1(n_210),
.A2(n_49),
.B1(n_50),
.B2(n_52),
.Y(n_278)
);

OAI22xp33_ASAP7_75t_SL g279 ( 
.A1(n_234),
.A2(n_218),
.B1(n_202),
.B2(n_214),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_199),
.Y(n_280)
);

AND2x2_ASAP7_75t_L g281 ( 
.A(n_202),
.B(n_54),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_272),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_246),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_250),
.Y(n_284)
);

AND2x2_ASAP7_75t_L g285 ( 
.A(n_240),
.B(n_234),
.Y(n_285)
);

AND2x6_ASAP7_75t_L g286 ( 
.A(n_269),
.B(n_199),
.Y(n_286)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_243),
.Y(n_287)
);

INVx2_ASAP7_75t_L g288 ( 
.A(n_244),
.Y(n_288)
);

CKINVDCx14_ASAP7_75t_R g289 ( 
.A(n_245),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_237),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_242),
.B(n_234),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_SL g292 ( 
.A(n_269),
.B(n_234),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_238),
.Y(n_293)
);

BUFx3_ASAP7_75t_L g294 ( 
.A(n_242),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_241),
.Y(n_295)
);

AND2x4_ASAP7_75t_L g296 ( 
.A(n_252),
.B(n_214),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_262),
.Y(n_297)
);

OR2x6_ASAP7_75t_L g298 ( 
.A(n_278),
.B(n_199),
.Y(n_298)
);

INVx3_ASAP7_75t_R g299 ( 
.A(n_255),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_245),
.B(n_234),
.Y(n_300)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_261),
.Y(n_301)
);

INVxp33_ASAP7_75t_L g302 ( 
.A(n_237),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_249),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_271),
.Y(n_304)
);

INVxp33_ASAP7_75t_L g305 ( 
.A(n_249),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_257),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_251),
.B(n_202),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_277),
.Y(n_308)
);

AND2x6_ASAP7_75t_L g309 ( 
.A(n_281),
.B(n_199),
.Y(n_309)
);

AND2x2_ASAP7_75t_L g310 ( 
.A(n_256),
.B(n_202),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_258),
.B(n_218),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_235),
.B(n_218),
.Y(n_312)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_263),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_280),
.Y(n_314)
);

AND2x2_ASAP7_75t_L g315 ( 
.A(n_278),
.B(n_218),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_273),
.Y(n_316)
);

INVxp33_ASAP7_75t_L g317 ( 
.A(n_259),
.Y(n_317)
);

XOR2xp5_ASAP7_75t_L g318 ( 
.A(n_239),
.B(n_55),
.Y(n_318)
);

AND2x2_ASAP7_75t_L g319 ( 
.A(n_276),
.B(n_218),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_274),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_248),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_248),
.Y(n_322)
);

XOR2xp5_ASAP7_75t_L g323 ( 
.A(n_236),
.B(n_56),
.Y(n_323)
);

XOR2xp5_ASAP7_75t_L g324 ( 
.A(n_277),
.B(n_57),
.Y(n_324)
);

OAI21xp5_ASAP7_75t_L g325 ( 
.A1(n_279),
.A2(n_217),
.B(n_214),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_248),
.Y(n_326)
);

INVx2_ASAP7_75t_SL g327 ( 
.A(n_260),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_247),
.B(n_199),
.Y(n_328)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_270),
.Y(n_329)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_266),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_264),
.B(n_201),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_267),
.B(n_201),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_265),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_259),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_275),
.B(n_201),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_253),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_254),
.B(n_201),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_268),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_272),
.Y(n_339)
);

XNOR2x2_ASAP7_75t_L g340 ( 
.A(n_237),
.B(n_214),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_272),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_SL g342 ( 
.A(n_236),
.B(n_214),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_272),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_272),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_272),
.Y(n_345)
);

NOR2xp67_ASAP7_75t_L g346 ( 
.A(n_306),
.B(n_58),
.Y(n_346)
);

BUFx8_ASAP7_75t_L g347 ( 
.A(n_330),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g348 ( 
.A(n_305),
.B(n_214),
.Y(n_348)
);

INVx3_ASAP7_75t_L g349 ( 
.A(n_294),
.Y(n_349)
);

INVx2_ASAP7_75t_L g350 ( 
.A(n_283),
.Y(n_350)
);

INVx1_ASAP7_75t_SL g351 ( 
.A(n_282),
.Y(n_351)
);

AND2x2_ASAP7_75t_SL g352 ( 
.A(n_342),
.B(n_217),
.Y(n_352)
);

AND2x2_ASAP7_75t_L g353 ( 
.A(n_305),
.B(n_217),
.Y(n_353)
);

AND2x2_ASAP7_75t_L g354 ( 
.A(n_298),
.B(n_217),
.Y(n_354)
);

AND2x4_ASAP7_75t_L g355 ( 
.A(n_327),
.B(n_217),
.Y(n_355)
);

BUFx6f_ASAP7_75t_L g356 ( 
.A(n_294),
.Y(n_356)
);

AND2x2_ASAP7_75t_SL g357 ( 
.A(n_315),
.B(n_217),
.Y(n_357)
);

AND2x2_ASAP7_75t_L g358 ( 
.A(n_298),
.B(n_317),
.Y(n_358)
);

AND2x2_ASAP7_75t_L g359 ( 
.A(n_298),
.B(n_201),
.Y(n_359)
);

AND2x2_ASAP7_75t_SL g360 ( 
.A(n_329),
.B(n_212),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_284),
.Y(n_361)
);

AND2x4_ASAP7_75t_L g362 ( 
.A(n_333),
.B(n_61),
.Y(n_362)
);

INVx2_ASAP7_75t_L g363 ( 
.A(n_301),
.Y(n_363)
);

AND2x2_ASAP7_75t_L g364 ( 
.A(n_317),
.B(n_213),
.Y(n_364)
);

OR2x2_ASAP7_75t_L g365 ( 
.A(n_336),
.B(n_213),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_311),
.B(n_213),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_297),
.Y(n_367)
);

INVx2_ASAP7_75t_L g368 ( 
.A(n_313),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_L g369 ( 
.A(n_285),
.B(n_62),
.Y(n_369)
);

AND2x2_ASAP7_75t_L g370 ( 
.A(n_331),
.B(n_213),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_287),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_288),
.Y(n_372)
);

AND2x2_ASAP7_75t_L g373 ( 
.A(n_331),
.B(n_213),
.Y(n_373)
);

AND2x2_ASAP7_75t_L g374 ( 
.A(n_319),
.B(n_212),
.Y(n_374)
);

BUFx3_ASAP7_75t_L g375 ( 
.A(n_293),
.Y(n_375)
);

BUFx3_ASAP7_75t_L g376 ( 
.A(n_295),
.Y(n_376)
);

HB1xp67_ASAP7_75t_L g377 ( 
.A(n_345),
.Y(n_377)
);

INVx2_ASAP7_75t_L g378 ( 
.A(n_314),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_311),
.B(n_212),
.Y(n_379)
);

INVx2_ASAP7_75t_L g380 ( 
.A(n_316),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_320),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_300),
.B(n_212),
.Y(n_382)
);

AND2x6_ASAP7_75t_L g383 ( 
.A(n_296),
.B(n_212),
.Y(n_383)
);

BUFx3_ASAP7_75t_L g384 ( 
.A(n_296),
.Y(n_384)
);

OR2x2_ASAP7_75t_SL g385 ( 
.A(n_289),
.B(n_65),
.Y(n_385)
);

AND2x2_ASAP7_75t_L g386 ( 
.A(n_337),
.B(n_338),
.Y(n_386)
);

OAI21xp33_ASAP7_75t_L g387 ( 
.A1(n_332),
.A2(n_66),
.B(n_69),
.Y(n_387)
);

INVx1_ASAP7_75t_SL g388 ( 
.A(n_339),
.Y(n_388)
);

BUFx6f_ASAP7_75t_L g389 ( 
.A(n_309),
.Y(n_389)
);

INVx1_ASAP7_75t_SL g390 ( 
.A(n_341),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_300),
.B(n_72),
.Y(n_391)
);

BUFx3_ASAP7_75t_L g392 ( 
.A(n_309),
.Y(n_392)
);

AND2x2_ASAP7_75t_L g393 ( 
.A(n_337),
.B(n_74),
.Y(n_393)
);

INVx2_ASAP7_75t_L g394 ( 
.A(n_304),
.Y(n_394)
);

AND2x4_ASAP7_75t_L g395 ( 
.A(n_343),
.B(n_76),
.Y(n_395)
);

AND2x2_ASAP7_75t_L g396 ( 
.A(n_344),
.B(n_78),
.Y(n_396)
);

INVx2_ASAP7_75t_SL g397 ( 
.A(n_286),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_SL g398 ( 
.A(n_312),
.B(n_80),
.Y(n_398)
);

AND2x2_ASAP7_75t_L g399 ( 
.A(n_289),
.B(n_81),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_286),
.B(n_82),
.Y(n_400)
);

INVxp67_ASAP7_75t_SL g401 ( 
.A(n_292),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_286),
.B(n_140),
.Y(n_402)
);

BUFx2_ASAP7_75t_L g403 ( 
.A(n_340),
.Y(n_403)
);

AND2x2_ASAP7_75t_L g404 ( 
.A(n_302),
.B(n_83),
.Y(n_404)
);

INVx2_ASAP7_75t_L g405 ( 
.A(n_321),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_322),
.Y(n_406)
);

INVx3_ASAP7_75t_L g407 ( 
.A(n_309),
.Y(n_407)
);

INVx6_ASAP7_75t_L g408 ( 
.A(n_309),
.Y(n_408)
);

HB1xp67_ASAP7_75t_L g409 ( 
.A(n_334),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_L g410 ( 
.A(n_302),
.B(n_138),
.Y(n_410)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_326),
.Y(n_411)
);

AND2x2_ASAP7_75t_L g412 ( 
.A(n_292),
.B(n_86),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_335),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_SL g414 ( 
.A(n_312),
.B(n_87),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_394),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_386),
.B(n_286),
.Y(n_416)
);

BUFx6f_ASAP7_75t_L g417 ( 
.A(n_389),
.Y(n_417)
);

OR2x2_ASAP7_75t_L g418 ( 
.A(n_409),
.B(n_290),
.Y(n_418)
);

AND2x2_ASAP7_75t_L g419 ( 
.A(n_386),
.B(n_303),
.Y(n_419)
);

NOR2xp33_ASAP7_75t_SL g420 ( 
.A(n_410),
.B(n_308),
.Y(n_420)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_363),
.Y(n_421)
);

HB1xp67_ASAP7_75t_L g422 ( 
.A(n_351),
.Y(n_422)
);

AND2x2_ASAP7_75t_L g423 ( 
.A(n_358),
.B(n_332),
.Y(n_423)
);

NOR2xp33_ASAP7_75t_L g424 ( 
.A(n_358),
.B(n_299),
.Y(n_424)
);

CKINVDCx20_ASAP7_75t_R g425 ( 
.A(n_347),
.Y(n_425)
);

AND2x2_ASAP7_75t_L g426 ( 
.A(n_403),
.B(n_324),
.Y(n_426)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_363),
.Y(n_427)
);

INVx3_ASAP7_75t_L g428 ( 
.A(n_389),
.Y(n_428)
);

AND2x4_ASAP7_75t_L g429 ( 
.A(n_384),
.B(n_328),
.Y(n_429)
);

BUFx6f_ASAP7_75t_L g430 ( 
.A(n_389),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_394),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_413),
.B(n_364),
.Y(n_432)
);

INVx2_ASAP7_75t_L g433 ( 
.A(n_363),
.Y(n_433)
);

INVx1_ASAP7_75t_SL g434 ( 
.A(n_388),
.Y(n_434)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_368),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_413),
.B(n_286),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_347),
.Y(n_437)
);

BUFx2_ASAP7_75t_L g438 ( 
.A(n_384),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_364),
.B(n_328),
.Y(n_439)
);

AND2x2_ASAP7_75t_L g440 ( 
.A(n_403),
.B(n_325),
.Y(n_440)
);

INVx6_ASAP7_75t_L g441 ( 
.A(n_356),
.Y(n_441)
);

OR2x2_ASAP7_75t_L g442 ( 
.A(n_390),
.B(n_318),
.Y(n_442)
);

BUFx2_ASAP7_75t_L g443 ( 
.A(n_384),
.Y(n_443)
);

AND2x4_ASAP7_75t_L g444 ( 
.A(n_392),
.B(n_307),
.Y(n_444)
);

HB1xp67_ASAP7_75t_L g445 ( 
.A(n_377),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_375),
.B(n_310),
.Y(n_446)
);

BUFx3_ASAP7_75t_L g447 ( 
.A(n_347),
.Y(n_447)
);

OR2x6_ASAP7_75t_L g448 ( 
.A(n_362),
.B(n_323),
.Y(n_448)
);

NOR2x1_ASAP7_75t_L g449 ( 
.A(n_375),
.B(n_291),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_394),
.Y(n_450)
);

INVx3_ASAP7_75t_L g451 ( 
.A(n_389),
.Y(n_451)
);

INVxp67_ASAP7_75t_L g452 ( 
.A(n_396),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_375),
.B(n_309),
.Y(n_453)
);

INVx2_ASAP7_75t_L g454 ( 
.A(n_368),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_367),
.Y(n_455)
);

HB1xp67_ASAP7_75t_L g456 ( 
.A(n_359),
.Y(n_456)
);

AND2x2_ASAP7_75t_L g457 ( 
.A(n_404),
.B(n_291),
.Y(n_457)
);

BUFx8_ASAP7_75t_L g458 ( 
.A(n_404),
.Y(n_458)
);

NAND2x1p5_ASAP7_75t_L g459 ( 
.A(n_392),
.B(n_88),
.Y(n_459)
);

INVx2_ASAP7_75t_L g460 ( 
.A(n_368),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_376),
.B(n_89),
.Y(n_461)
);

BUFx6f_ASAP7_75t_L g462 ( 
.A(n_389),
.Y(n_462)
);

BUFx2_ASAP7_75t_L g463 ( 
.A(n_392),
.Y(n_463)
);

OR2x6_ASAP7_75t_L g464 ( 
.A(n_362),
.B(n_90),
.Y(n_464)
);

AND2x2_ASAP7_75t_L g465 ( 
.A(n_393),
.B(n_91),
.Y(n_465)
);

BUFx6f_ASAP7_75t_L g466 ( 
.A(n_389),
.Y(n_466)
);

AND2x2_ASAP7_75t_L g467 ( 
.A(n_393),
.B(n_92),
.Y(n_467)
);

BUFx2_ASAP7_75t_SL g468 ( 
.A(n_407),
.Y(n_468)
);

INVx5_ASAP7_75t_L g469 ( 
.A(n_408),
.Y(n_469)
);

BUFx3_ASAP7_75t_L g470 ( 
.A(n_347),
.Y(n_470)
);

BUFx5_ASAP7_75t_L g471 ( 
.A(n_465),
.Y(n_471)
);

AND2x2_ASAP7_75t_L g472 ( 
.A(n_419),
.B(n_399),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_455),
.Y(n_473)
);

INVx2_ASAP7_75t_L g474 ( 
.A(n_421),
.Y(n_474)
);

INVx3_ASAP7_75t_SL g475 ( 
.A(n_437),
.Y(n_475)
);

NAND2x1p5_ASAP7_75t_L g476 ( 
.A(n_469),
.B(n_407),
.Y(n_476)
);

BUFx3_ASAP7_75t_L g477 ( 
.A(n_447),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_423),
.B(n_376),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_415),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_423),
.B(n_376),
.Y(n_480)
);

BUFx2_ASAP7_75t_SL g481 ( 
.A(n_425),
.Y(n_481)
);

BUFx6f_ASAP7_75t_SL g482 ( 
.A(n_447),
.Y(n_482)
);

BUFx10_ASAP7_75t_L g483 ( 
.A(n_417),
.Y(n_483)
);

CKINVDCx16_ASAP7_75t_R g484 ( 
.A(n_425),
.Y(n_484)
);

AOI22xp33_ASAP7_75t_L g485 ( 
.A1(n_448),
.A2(n_362),
.B1(n_399),
.B2(n_367),
.Y(n_485)
);

BUFx6f_ASAP7_75t_L g486 ( 
.A(n_469),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_431),
.Y(n_487)
);

INVx5_ASAP7_75t_L g488 ( 
.A(n_469),
.Y(n_488)
);

INVx3_ASAP7_75t_L g489 ( 
.A(n_469),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_450),
.Y(n_490)
);

AND2x4_ASAP7_75t_L g491 ( 
.A(n_469),
.B(n_395),
.Y(n_491)
);

BUFx3_ASAP7_75t_L g492 ( 
.A(n_470),
.Y(n_492)
);

BUFx6f_ASAP7_75t_L g493 ( 
.A(n_417),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_421),
.Y(n_494)
);

CKINVDCx11_ASAP7_75t_R g495 ( 
.A(n_434),
.Y(n_495)
);

INVxp67_ASAP7_75t_SL g496 ( 
.A(n_463),
.Y(n_496)
);

OR2x2_ASAP7_75t_L g497 ( 
.A(n_418),
.B(n_385),
.Y(n_497)
);

BUFx2_ASAP7_75t_L g498 ( 
.A(n_422),
.Y(n_498)
);

NOR2xp33_ASAP7_75t_L g499 ( 
.A(n_420),
.B(n_385),
.Y(n_499)
);

BUFx4_ASAP7_75t_SL g500 ( 
.A(n_437),
.Y(n_500)
);

NAND2x1p5_ASAP7_75t_L g501 ( 
.A(n_463),
.B(n_438),
.Y(n_501)
);

INVx2_ASAP7_75t_L g502 ( 
.A(n_427),
.Y(n_502)
);

CKINVDCx5p33_ASAP7_75t_R g503 ( 
.A(n_470),
.Y(n_503)
);

INVx2_ASAP7_75t_SL g504 ( 
.A(n_417),
.Y(n_504)
);

INVx3_ASAP7_75t_L g505 ( 
.A(n_417),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_427),
.Y(n_506)
);

INVx2_ASAP7_75t_L g507 ( 
.A(n_433),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_433),
.Y(n_508)
);

BUFx12f_ASAP7_75t_L g509 ( 
.A(n_418),
.Y(n_509)
);

BUFx2_ASAP7_75t_SL g510 ( 
.A(n_445),
.Y(n_510)
);

CKINVDCx20_ASAP7_75t_R g511 ( 
.A(n_458),
.Y(n_511)
);

INVx5_ASAP7_75t_L g512 ( 
.A(n_417),
.Y(n_512)
);

BUFx12f_ASAP7_75t_L g513 ( 
.A(n_458),
.Y(n_513)
);

INVx3_ASAP7_75t_L g514 ( 
.A(n_430),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_440),
.B(n_362),
.Y(n_515)
);

AOI22xp33_ASAP7_75t_L g516 ( 
.A1(n_485),
.A2(n_426),
.B1(n_448),
.B2(n_419),
.Y(n_516)
);

INVx4_ASAP7_75t_L g517 ( 
.A(n_488),
.Y(n_517)
);

INVx11_ASAP7_75t_L g518 ( 
.A(n_513),
.Y(n_518)
);

OAI22xp5_ASAP7_75t_L g519 ( 
.A1(n_485),
.A2(n_452),
.B1(n_448),
.B2(n_464),
.Y(n_519)
);

AOI22xp33_ASAP7_75t_L g520 ( 
.A1(n_499),
.A2(n_426),
.B1(n_448),
.B2(n_442),
.Y(n_520)
);

BUFx6f_ASAP7_75t_L g521 ( 
.A(n_488),
.Y(n_521)
);

INVx2_ASAP7_75t_SL g522 ( 
.A(n_500),
.Y(n_522)
);

INVx1_ASAP7_75t_SL g523 ( 
.A(n_510),
.Y(n_523)
);

INVx6_ASAP7_75t_L g524 ( 
.A(n_513),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_473),
.Y(n_525)
);

INVx3_ASAP7_75t_L g526 ( 
.A(n_491),
.Y(n_526)
);

INVx11_ASAP7_75t_L g527 ( 
.A(n_509),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_472),
.B(n_440),
.Y(n_528)
);

INVx4_ASAP7_75t_L g529 ( 
.A(n_488),
.Y(n_529)
);

INVx6_ASAP7_75t_L g530 ( 
.A(n_509),
.Y(n_530)
);

BUFx6f_ASAP7_75t_L g531 ( 
.A(n_488),
.Y(n_531)
);

OAI22xp5_ASAP7_75t_L g532 ( 
.A1(n_515),
.A2(n_464),
.B1(n_467),
.B2(n_465),
.Y(n_532)
);

OAI22xp5_ASAP7_75t_L g533 ( 
.A1(n_496),
.A2(n_464),
.B1(n_467),
.B2(n_395),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_479),
.Y(n_534)
);

AOI22xp33_ASAP7_75t_L g535 ( 
.A1(n_499),
.A2(n_442),
.B1(n_458),
.B2(n_464),
.Y(n_535)
);

OAI22xp5_ASAP7_75t_L g536 ( 
.A1(n_497),
.A2(n_395),
.B1(n_457),
.B2(n_391),
.Y(n_536)
);

CKINVDCx5p33_ASAP7_75t_R g537 ( 
.A(n_495),
.Y(n_537)
);

BUFx2_ASAP7_75t_SL g538 ( 
.A(n_482),
.Y(n_538)
);

OAI22xp33_ASAP7_75t_L g539 ( 
.A1(n_484),
.A2(n_443),
.B1(n_438),
.B2(n_456),
.Y(n_539)
);

INVx2_ASAP7_75t_L g540 ( 
.A(n_487),
.Y(n_540)
);

AOI22xp5_ASAP7_75t_L g541 ( 
.A1(n_478),
.A2(n_387),
.B1(n_429),
.B2(n_424),
.Y(n_541)
);

AOI22xp33_ASAP7_75t_L g542 ( 
.A1(n_480),
.A2(n_429),
.B1(n_369),
.B2(n_444),
.Y(n_542)
);

CKINVDCx11_ASAP7_75t_R g543 ( 
.A(n_495),
.Y(n_543)
);

INVx2_ASAP7_75t_SL g544 ( 
.A(n_503),
.Y(n_544)
);

INVx6_ASAP7_75t_L g545 ( 
.A(n_477),
.Y(n_545)
);

OR2x2_ASAP7_75t_L g546 ( 
.A(n_498),
.B(n_429),
.Y(n_546)
);

OAI22xp5_ASAP7_75t_L g547 ( 
.A1(n_491),
.A2(n_395),
.B1(n_457),
.B2(n_352),
.Y(n_547)
);

OAI21xp5_ASAP7_75t_L g548 ( 
.A1(n_490),
.A2(n_449),
.B(n_346),
.Y(n_548)
);

CKINVDCx20_ASAP7_75t_R g549 ( 
.A(n_511),
.Y(n_549)
);

BUFx2_ASAP7_75t_SL g550 ( 
.A(n_482),
.Y(n_550)
);

INVx2_ASAP7_75t_L g551 ( 
.A(n_474),
.Y(n_551)
);

AOI22xp33_ASAP7_75t_SL g552 ( 
.A1(n_471),
.A2(n_352),
.B1(n_360),
.B2(n_412),
.Y(n_552)
);

OAI22xp5_ASAP7_75t_L g553 ( 
.A1(n_491),
.A2(n_501),
.B1(n_352),
.B2(n_475),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_503),
.B(n_443),
.Y(n_554)
);

INVx2_ASAP7_75t_SL g555 ( 
.A(n_518),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_525),
.Y(n_556)
);

AOI22xp33_ASAP7_75t_L g557 ( 
.A1(n_516),
.A2(n_387),
.B1(n_350),
.B2(n_361),
.Y(n_557)
);

INVx2_ASAP7_75t_L g558 ( 
.A(n_551),
.Y(n_558)
);

BUFx3_ASAP7_75t_L g559 ( 
.A(n_545),
.Y(n_559)
);

BUFx3_ASAP7_75t_L g560 ( 
.A(n_545),
.Y(n_560)
);

AOI22xp33_ASAP7_75t_L g561 ( 
.A1(n_519),
.A2(n_350),
.B1(n_361),
.B2(n_371),
.Y(n_561)
);

AOI22xp33_ASAP7_75t_L g562 ( 
.A1(n_520),
.A2(n_536),
.B1(n_535),
.B2(n_528),
.Y(n_562)
);

INVx2_ASAP7_75t_SL g563 ( 
.A(n_527),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_540),
.Y(n_564)
);

AOI22xp33_ASAP7_75t_SL g565 ( 
.A1(n_533),
.A2(n_471),
.B1(n_360),
.B2(n_511),
.Y(n_565)
);

AOI22xp33_ASAP7_75t_L g566 ( 
.A1(n_552),
.A2(n_371),
.B1(n_372),
.B2(n_471),
.Y(n_566)
);

OAI22xp5_ASAP7_75t_L g567 ( 
.A1(n_532),
.A2(n_475),
.B1(n_481),
.B2(n_501),
.Y(n_567)
);

BUFx6f_ASAP7_75t_L g568 ( 
.A(n_521),
.Y(n_568)
);

CKINVDCx14_ASAP7_75t_R g569 ( 
.A(n_543),
.Y(n_569)
);

AND2x2_ASAP7_75t_L g570 ( 
.A(n_546),
.B(n_477),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_534),
.Y(n_571)
);

AOI22xp33_ASAP7_75t_L g572 ( 
.A1(n_547),
.A2(n_372),
.B1(n_471),
.B2(n_378),
.Y(n_572)
);

AND2x2_ASAP7_75t_L g573 ( 
.A(n_523),
.B(n_544),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_554),
.Y(n_574)
);

AOI222xp33_ASAP7_75t_L g575 ( 
.A1(n_539),
.A2(n_353),
.B1(n_348),
.B2(n_357),
.C1(n_396),
.C2(n_412),
.Y(n_575)
);

AND2x2_ASAP7_75t_L g576 ( 
.A(n_523),
.B(n_492),
.Y(n_576)
);

AOI22xp33_ASAP7_75t_L g577 ( 
.A1(n_542),
.A2(n_471),
.B1(n_378),
.B2(n_444),
.Y(n_577)
);

AOI22xp33_ASAP7_75t_L g578 ( 
.A1(n_541),
.A2(n_471),
.B1(n_444),
.B2(n_439),
.Y(n_578)
);

INVx5_ASAP7_75t_SL g579 ( 
.A(n_521),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_526),
.Y(n_580)
);

AOI22xp33_ASAP7_75t_L g581 ( 
.A1(n_541),
.A2(n_471),
.B1(n_432),
.B2(n_381),
.Y(n_581)
);

BUFx6f_ASAP7_75t_L g582 ( 
.A(n_521),
.Y(n_582)
);

AOI22xp33_ASAP7_75t_SL g583 ( 
.A1(n_553),
.A2(n_360),
.B1(n_459),
.B2(n_357),
.Y(n_583)
);

OAI21xp5_ASAP7_75t_SL g584 ( 
.A1(n_522),
.A2(n_459),
.B(n_354),
.Y(n_584)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_526),
.Y(n_585)
);

INVx2_ASAP7_75t_L g586 ( 
.A(n_531),
.Y(n_586)
);

BUFx2_ASAP7_75t_L g587 ( 
.A(n_530),
.Y(n_587)
);

OAI22xp33_ASAP7_75t_L g588 ( 
.A1(n_530),
.A2(n_492),
.B1(n_416),
.B2(n_446),
.Y(n_588)
);

AOI22xp33_ASAP7_75t_SL g589 ( 
.A1(n_538),
.A2(n_459),
.B1(n_357),
.B2(n_353),
.Y(n_589)
);

INVx4_ASAP7_75t_L g590 ( 
.A(n_524),
.Y(n_590)
);

AOI22xp33_ASAP7_75t_L g591 ( 
.A1(n_524),
.A2(n_381),
.B1(n_414),
.B2(n_398),
.Y(n_591)
);

OAI22xp5_ASAP7_75t_L g592 ( 
.A1(n_549),
.A2(n_346),
.B1(n_349),
.B2(n_356),
.Y(n_592)
);

AOI22xp33_ASAP7_75t_L g593 ( 
.A1(n_548),
.A2(n_380),
.B1(n_508),
.B2(n_506),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_L g594 ( 
.A(n_550),
.B(n_494),
.Y(n_594)
);

OAI22xp5_ASAP7_75t_L g595 ( 
.A1(n_537),
.A2(n_349),
.B1(n_356),
.B2(n_453),
.Y(n_595)
);

OAI222xp33_ASAP7_75t_L g596 ( 
.A1(n_517),
.A2(n_365),
.B1(n_507),
.B2(n_502),
.C1(n_474),
.C2(n_460),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_L g597 ( 
.A(n_531),
.B(n_502),
.Y(n_597)
);

OAI22xp5_ASAP7_75t_L g598 ( 
.A1(n_548),
.A2(n_349),
.B1(n_356),
.B2(n_461),
.Y(n_598)
);

AOI22xp33_ASAP7_75t_L g599 ( 
.A1(n_531),
.A2(n_380),
.B1(n_365),
.B2(n_460),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_L g600 ( 
.A(n_517),
.B(n_507),
.Y(n_600)
);

AOI22xp5_ASAP7_75t_L g601 ( 
.A1(n_575),
.A2(n_354),
.B1(n_359),
.B2(n_401),
.Y(n_601)
);

OAI222xp33_ASAP7_75t_L g602 ( 
.A1(n_562),
.A2(n_565),
.B1(n_561),
.B2(n_557),
.C1(n_566),
.C2(n_583),
.Y(n_602)
);

AOI22xp33_ASAP7_75t_L g603 ( 
.A1(n_562),
.A2(n_380),
.B1(n_454),
.B2(n_435),
.Y(n_603)
);

AOI221xp5_ASAP7_75t_L g604 ( 
.A1(n_574),
.A2(n_406),
.B1(n_374),
.B2(n_405),
.C(n_411),
.Y(n_604)
);

AOI22xp33_ASAP7_75t_SL g605 ( 
.A1(n_567),
.A2(n_373),
.B1(n_370),
.B2(n_529),
.Y(n_605)
);

OAI22xp5_ASAP7_75t_L g606 ( 
.A1(n_581),
.A2(n_441),
.B1(n_356),
.B2(n_512),
.Y(n_606)
);

OAI22xp5_ASAP7_75t_L g607 ( 
.A1(n_581),
.A2(n_441),
.B1(n_356),
.B2(n_512),
.Y(n_607)
);

AOI21xp5_ASAP7_75t_L g608 ( 
.A1(n_584),
.A2(n_512),
.B(n_493),
.Y(n_608)
);

AND2x2_ASAP7_75t_L g609 ( 
.A(n_570),
.B(n_576),
.Y(n_609)
);

AND2x2_ASAP7_75t_L g610 ( 
.A(n_573),
.B(n_505),
.Y(n_610)
);

AOI22xp33_ASAP7_75t_SL g611 ( 
.A1(n_592),
.A2(n_370),
.B1(n_373),
.B2(n_529),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_L g612 ( 
.A(n_556),
.B(n_571),
.Y(n_612)
);

NAND2x1p5_ASAP7_75t_L g613 ( 
.A(n_568),
.B(n_512),
.Y(n_613)
);

OAI22xp5_ASAP7_75t_L g614 ( 
.A1(n_578),
.A2(n_441),
.B1(n_349),
.B2(n_514),
.Y(n_614)
);

OAI22xp5_ASAP7_75t_L g615 ( 
.A1(n_578),
.A2(n_441),
.B1(n_505),
.B2(n_514),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_L g616 ( 
.A(n_564),
.B(n_505),
.Y(n_616)
);

AOI22xp33_ASAP7_75t_L g617 ( 
.A1(n_557),
.A2(n_561),
.B1(n_566),
.B2(n_577),
.Y(n_617)
);

AND2x2_ASAP7_75t_L g618 ( 
.A(n_559),
.B(n_514),
.Y(n_618)
);

OAI211xp5_ASAP7_75t_L g619 ( 
.A1(n_572),
.A2(n_406),
.B(n_411),
.C(n_405),
.Y(n_619)
);

OAI222xp33_ASAP7_75t_L g620 ( 
.A1(n_589),
.A2(n_454),
.B1(n_435),
.B2(n_411),
.C1(n_405),
.C2(n_382),
.Y(n_620)
);

OAI22xp5_ASAP7_75t_L g621 ( 
.A1(n_572),
.A2(n_504),
.B1(n_428),
.B2(n_451),
.Y(n_621)
);

AOI22xp33_ASAP7_75t_L g622 ( 
.A1(n_577),
.A2(n_374),
.B1(n_436),
.B2(n_379),
.Y(n_622)
);

AOI22xp33_ASAP7_75t_L g623 ( 
.A1(n_591),
.A2(n_366),
.B1(n_355),
.B2(n_468),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_558),
.Y(n_624)
);

AOI22xp33_ASAP7_75t_L g625 ( 
.A1(n_588),
.A2(n_468),
.B1(n_355),
.B2(n_383),
.Y(n_625)
);

OAI22xp5_ASAP7_75t_SL g626 ( 
.A1(n_569),
.A2(n_486),
.B1(n_493),
.B2(n_462),
.Y(n_626)
);

AOI22xp33_ASAP7_75t_L g627 ( 
.A1(n_591),
.A2(n_355),
.B1(n_383),
.B2(n_428),
.Y(n_627)
);

AOI221xp5_ASAP7_75t_L g628 ( 
.A1(n_594),
.A2(n_593),
.B1(n_580),
.B2(n_595),
.C(n_587),
.Y(n_628)
);

OAI22xp5_ASAP7_75t_L g629 ( 
.A1(n_590),
.A2(n_504),
.B1(n_428),
.B2(n_451),
.Y(n_629)
);

AOI22xp33_ASAP7_75t_SL g630 ( 
.A1(n_598),
.A2(n_355),
.B1(n_430),
.B2(n_462),
.Y(n_630)
);

NOR2xp33_ASAP7_75t_L g631 ( 
.A(n_559),
.B(n_560),
.Y(n_631)
);

AOI22xp33_ASAP7_75t_L g632 ( 
.A1(n_558),
.A2(n_383),
.B1(n_451),
.B2(n_430),
.Y(n_632)
);

AOI211xp5_ASAP7_75t_L g633 ( 
.A1(n_560),
.A2(n_400),
.B(n_402),
.C(n_493),
.Y(n_633)
);

NAND3xp33_ASAP7_75t_L g634 ( 
.A(n_593),
.B(n_493),
.C(n_462),
.Y(n_634)
);

AND2x2_ASAP7_75t_L g635 ( 
.A(n_585),
.B(n_483),
.Y(n_635)
);

NOR3xp33_ASAP7_75t_L g636 ( 
.A(n_590),
.B(n_586),
.C(n_563),
.Y(n_636)
);

OAI22xp5_ASAP7_75t_L g637 ( 
.A1(n_599),
.A2(n_462),
.B1(n_430),
.B2(n_466),
.Y(n_637)
);

AND2x2_ASAP7_75t_SL g638 ( 
.A(n_617),
.B(n_582),
.Y(n_638)
);

AND2x2_ASAP7_75t_L g639 ( 
.A(n_609),
.B(n_568),
.Y(n_639)
);

AND2x2_ASAP7_75t_L g640 ( 
.A(n_610),
.B(n_568),
.Y(n_640)
);

AND2x2_ASAP7_75t_L g641 ( 
.A(n_612),
.B(n_568),
.Y(n_641)
);

OAI22xp5_ASAP7_75t_L g642 ( 
.A1(n_617),
.A2(n_599),
.B1(n_579),
.B2(n_555),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_L g643 ( 
.A(n_616),
.B(n_600),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_L g644 ( 
.A(n_618),
.B(n_582),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_SL g645 ( 
.A(n_628),
.B(n_633),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_L g646 ( 
.A(n_631),
.B(n_582),
.Y(n_646)
);

AND2x2_ASAP7_75t_SL g647 ( 
.A(n_636),
.B(n_582),
.Y(n_647)
);

NOR3xp33_ASAP7_75t_L g648 ( 
.A(n_602),
.B(n_597),
.C(n_596),
.Y(n_648)
);

NAND4xp25_ASAP7_75t_L g649 ( 
.A(n_605),
.B(n_407),
.C(n_489),
.D(n_579),
.Y(n_649)
);

NAND3xp33_ASAP7_75t_L g650 ( 
.A(n_604),
.B(n_466),
.C(n_430),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_L g651 ( 
.A(n_635),
.B(n_579),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_603),
.B(n_483),
.Y(n_652)
);

OAI221xp5_ASAP7_75t_L g653 ( 
.A1(n_611),
.A2(n_408),
.B1(n_407),
.B2(n_397),
.C(n_489),
.Y(n_653)
);

NAND3xp33_ASAP7_75t_L g654 ( 
.A(n_634),
.B(n_466),
.C(n_462),
.Y(n_654)
);

XNOR2x1_ASAP7_75t_L g655 ( 
.A(n_601),
.B(n_93),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_603),
.B(n_483),
.Y(n_656)
);

OAI21xp5_ASAP7_75t_SL g657 ( 
.A1(n_608),
.A2(n_606),
.B(n_607),
.Y(n_657)
);

AND2x2_ASAP7_75t_L g658 ( 
.A(n_624),
.B(n_466),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_L g659 ( 
.A(n_626),
.B(n_489),
.Y(n_659)
);

AND2x2_ASAP7_75t_L g660 ( 
.A(n_613),
.B(n_615),
.Y(n_660)
);

NAND3xp33_ASAP7_75t_L g661 ( 
.A(n_619),
.B(n_466),
.C(n_486),
.Y(n_661)
);

AND2x2_ASAP7_75t_L g662 ( 
.A(n_623),
.B(n_94),
.Y(n_662)
);

AND2x2_ASAP7_75t_L g663 ( 
.A(n_623),
.B(n_95),
.Y(n_663)
);

AND2x2_ASAP7_75t_L g664 ( 
.A(n_630),
.B(n_96),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_L g665 ( 
.A(n_641),
.B(n_643),
.Y(n_665)
);

AND2x2_ASAP7_75t_L g666 ( 
.A(n_639),
.B(n_637),
.Y(n_666)
);

AND2x4_ASAP7_75t_L g667 ( 
.A(n_641),
.B(n_625),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_639),
.B(n_640),
.Y(n_668)
);

AND2x2_ASAP7_75t_L g669 ( 
.A(n_640),
.B(n_613),
.Y(n_669)
);

NOR3xp33_ASAP7_75t_L g670 ( 
.A(n_645),
.B(n_629),
.C(n_621),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_SL g671 ( 
.A(n_647),
.B(n_638),
.Y(n_671)
);

AND2x2_ASAP7_75t_L g672 ( 
.A(n_644),
.B(n_614),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_658),
.Y(n_673)
);

OR2x2_ASAP7_75t_L g674 ( 
.A(n_646),
.B(n_622),
.Y(n_674)
);

AND2x2_ASAP7_75t_L g675 ( 
.A(n_660),
.B(n_627),
.Y(n_675)
);

AND2x2_ASAP7_75t_L g676 ( 
.A(n_638),
.B(n_632),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_647),
.B(n_622),
.Y(n_677)
);

OA211x2_ASAP7_75t_L g678 ( 
.A1(n_645),
.A2(n_659),
.B(n_661),
.C(n_651),
.Y(n_678)
);

NOR3xp33_ASAP7_75t_L g679 ( 
.A(n_657),
.B(n_620),
.C(n_397),
.Y(n_679)
);

INVx2_ASAP7_75t_L g680 ( 
.A(n_654),
.Y(n_680)
);

NOR2xp33_ASAP7_75t_L g681 ( 
.A(n_665),
.B(n_649),
.Y(n_681)
);

AND2x2_ASAP7_75t_L g682 ( 
.A(n_666),
.B(n_642),
.Y(n_682)
);

XOR2x2_ASAP7_75t_L g683 ( 
.A(n_671),
.B(n_655),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_680),
.B(n_650),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_L g685 ( 
.A(n_680),
.B(n_672),
.Y(n_685)
);

XOR2x2_ASAP7_75t_L g686 ( 
.A(n_671),
.B(n_655),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_673),
.Y(n_687)
);

NAND4xp75_ASAP7_75t_SL g688 ( 
.A(n_678),
.B(n_663),
.C(n_662),
.D(n_664),
.Y(n_688)
);

NAND4xp75_ASAP7_75t_SL g689 ( 
.A(n_666),
.B(n_663),
.C(n_662),
.D(n_664),
.Y(n_689)
);

NAND4xp75_ASAP7_75t_L g690 ( 
.A(n_676),
.B(n_656),
.C(n_652),
.D(n_648),
.Y(n_690)
);

BUFx3_ASAP7_75t_L g691 ( 
.A(n_669),
.Y(n_691)
);

OR2x2_ASAP7_75t_L g692 ( 
.A(n_685),
.B(n_684),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_687),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_L g694 ( 
.A(n_681),
.B(n_672),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_682),
.Y(n_695)
);

XOR2x2_ASAP7_75t_L g696 ( 
.A(n_683),
.B(n_675),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_693),
.Y(n_697)
);

INVx2_ASAP7_75t_SL g698 ( 
.A(n_695),
.Y(n_698)
);

AOI22x1_ASAP7_75t_L g699 ( 
.A1(n_692),
.A2(n_688),
.B1(n_686),
.B2(n_689),
.Y(n_699)
);

HB1xp67_ASAP7_75t_L g700 ( 
.A(n_694),
.Y(n_700)
);

AOI22x1_ASAP7_75t_L g701 ( 
.A1(n_696),
.A2(n_688),
.B1(n_689),
.B2(n_690),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_697),
.Y(n_702)
);

HB1xp67_ASAP7_75t_L g703 ( 
.A(n_700),
.Y(n_703)
);

INVx2_ASAP7_75t_SL g704 ( 
.A(n_701),
.Y(n_704)
);

INVxp67_ASAP7_75t_SL g705 ( 
.A(n_701),
.Y(n_705)
);

NOR4xp25_ASAP7_75t_L g706 ( 
.A(n_704),
.B(n_705),
.C(n_702),
.D(n_694),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_702),
.Y(n_707)
);

INVx2_ASAP7_75t_SL g708 ( 
.A(n_703),
.Y(n_708)
);

AOI311xp33_ASAP7_75t_L g709 ( 
.A1(n_704),
.A2(n_699),
.A3(n_681),
.B(n_670),
.C(n_698),
.Y(n_709)
);

INVx2_ASAP7_75t_L g710 ( 
.A(n_708),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_708),
.Y(n_711)
);

INVxp67_ASAP7_75t_L g712 ( 
.A(n_707),
.Y(n_712)
);

A2O1A1Ixp33_ASAP7_75t_L g713 ( 
.A1(n_706),
.A2(n_699),
.B(n_698),
.C(n_677),
.Y(n_713)
);

AOI22xp33_ASAP7_75t_L g714 ( 
.A1(n_710),
.A2(n_712),
.B1(n_711),
.B2(n_679),
.Y(n_714)
);

AOI22xp5_ASAP7_75t_L g715 ( 
.A1(n_713),
.A2(n_709),
.B1(n_676),
.B2(n_675),
.Y(n_715)
);

OA22x2_ASAP7_75t_L g716 ( 
.A1(n_711),
.A2(n_667),
.B1(n_669),
.B2(n_668),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_L g717 ( 
.A(n_710),
.B(n_691),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_SL g718 ( 
.A(n_713),
.B(n_667),
.Y(n_718)
);

AOI22xp5_ASAP7_75t_L g719 ( 
.A1(n_713),
.A2(n_667),
.B1(n_674),
.B2(n_653),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_711),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_720),
.Y(n_721)
);

INVx2_ASAP7_75t_L g722 ( 
.A(n_716),
.Y(n_722)
);

INVx2_ASAP7_75t_L g723 ( 
.A(n_717),
.Y(n_723)
);

INVx2_ASAP7_75t_L g724 ( 
.A(n_718),
.Y(n_724)
);

INVxp67_ASAP7_75t_L g725 ( 
.A(n_715),
.Y(n_725)
);

AOI22xp5_ASAP7_75t_L g726 ( 
.A1(n_719),
.A2(n_408),
.B1(n_383),
.B2(n_486),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_714),
.Y(n_727)
);

INVx2_ASAP7_75t_L g728 ( 
.A(n_724),
.Y(n_728)
);

OAI22x1_ASAP7_75t_L g729 ( 
.A1(n_725),
.A2(n_476),
.B1(n_408),
.B2(n_486),
.Y(n_729)
);

INVx2_ASAP7_75t_L g730 ( 
.A(n_723),
.Y(n_730)
);

OAI22xp33_ASAP7_75t_L g731 ( 
.A1(n_722),
.A2(n_476),
.B1(n_383),
.B2(n_102),
.Y(n_731)
);

INVx2_ASAP7_75t_L g732 ( 
.A(n_721),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_727),
.Y(n_733)
);

OAI22xp33_ASAP7_75t_L g734 ( 
.A1(n_726),
.A2(n_383),
.B1(n_100),
.B2(n_103),
.Y(n_734)
);

AO22x2_ASAP7_75t_L g735 ( 
.A1(n_724),
.A2(n_97),
.B1(n_104),
.B2(n_106),
.Y(n_735)
);

AND2x2_ASAP7_75t_L g736 ( 
.A(n_728),
.B(n_108),
.Y(n_736)
);

AO22x2_ASAP7_75t_L g737 ( 
.A1(n_733),
.A2(n_110),
.B1(n_111),
.B2(n_112),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_730),
.Y(n_738)
);

BUFx6f_ASAP7_75t_L g739 ( 
.A(n_732),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_735),
.Y(n_740)
);

INVx2_ASAP7_75t_L g741 ( 
.A(n_729),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_731),
.Y(n_742)
);

AOI22xp5_ASAP7_75t_L g743 ( 
.A1(n_738),
.A2(n_734),
.B1(n_383),
.B2(n_118),
.Y(n_743)
);

BUFx2_ASAP7_75t_L g744 ( 
.A(n_739),
.Y(n_744)
);

OA22x2_ASAP7_75t_L g745 ( 
.A1(n_742),
.A2(n_113),
.B1(n_115),
.B2(n_119),
.Y(n_745)
);

OAI22x1_ASAP7_75t_L g746 ( 
.A1(n_740),
.A2(n_120),
.B1(n_122),
.B2(n_123),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_744),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_745),
.Y(n_748)
);

AO22x2_ASAP7_75t_L g749 ( 
.A1(n_748),
.A2(n_736),
.B1(n_741),
.B2(n_739),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_749),
.Y(n_750)
);

AO22x2_ASAP7_75t_L g751 ( 
.A1(n_750),
.A2(n_747),
.B1(n_746),
.B2(n_737),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_751),
.Y(n_752)
);

AOI221xp5_ASAP7_75t_L g753 ( 
.A1(n_752),
.A2(n_737),
.B1(n_743),
.B2(n_127),
.C(n_129),
.Y(n_753)
);

AOI22xp33_ASAP7_75t_L g754 ( 
.A1(n_753),
.A2(n_124),
.B1(n_125),
.B2(n_130),
.Y(n_754)
);


endmodule