module fake_jpeg_11051_n_94 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_2, n_29, n_12, n_8, n_15, n_7, n_94);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_29;
input n_12;
input n_8;
input n_15;
input n_7;

output n_94;

wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_31;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_44;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_20),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_23),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_29),
.Y(n_33)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_11),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_7),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_21),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_14),
.B(n_30),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_6),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_28),
.Y(n_39)
);

INVx1_ASAP7_75t_SL g40 ( 
.A(n_9),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_18),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_39),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_42),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_39),
.Y(n_43)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_43),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_SL g44 ( 
.A(n_37),
.B(n_0),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_44),
.B(n_45),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_40),
.B(n_0),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_31),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_46),
.Y(n_53)
);

HAxp5_ASAP7_75t_SL g47 ( 
.A(n_40),
.B(n_1),
.CON(n_47),
.SN(n_47)
);

OR2x2_ASAP7_75t_SL g54 ( 
.A(n_47),
.B(n_1),
.Y(n_54)
);

BUFx12_ASAP7_75t_L g48 ( 
.A(n_33),
.Y(n_48)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_48),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_49),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_42),
.A2(n_38),
.B1(n_34),
.B2(n_32),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_50),
.A2(n_38),
.B1(n_34),
.B2(n_36),
.Y(n_61)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_46),
.Y(n_51)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_51),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_45),
.B(n_32),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_52),
.B(n_54),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_59),
.B(n_41),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_60),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_61),
.A2(n_65),
.B1(n_71),
.B2(n_57),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_58),
.B(n_49),
.Y(n_62)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_62),
.Y(n_75)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_58),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_63),
.Y(n_78)
);

INVx1_ASAP7_75t_SL g64 ( 
.A(n_56),
.Y(n_64)
);

INVx13_ASAP7_75t_L g73 ( 
.A(n_64),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_57),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_65)
);

OAI21xp5_ASAP7_75t_L g68 ( 
.A1(n_53),
.A2(n_48),
.B(n_3),
.Y(n_68)
);

OAI21xp5_ASAP7_75t_L g74 ( 
.A1(n_68),
.A2(n_53),
.B(n_5),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_55),
.B(n_2),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_69),
.Y(n_80)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_55),
.Y(n_70)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_70),
.B(n_8),
.C(n_10),
.Y(n_77)
);

O2A1O1Ixp33_ASAP7_75t_SL g71 ( 
.A1(n_56),
.A2(n_16),
.B(n_26),
.C(n_25),
.Y(n_71)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_72),
.B(n_74),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_76),
.B(n_77),
.C(n_24),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_68),
.A2(n_12),
.B1(n_13),
.B2(n_15),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_79),
.A2(n_81),
.B1(n_66),
.B2(n_64),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_71),
.A2(n_17),
.B1(n_19),
.B2(n_22),
.Y(n_81)
);

NOR3xp33_ASAP7_75t_L g86 ( 
.A(n_82),
.B(n_83),
.C(n_74),
.Y(n_86)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_78),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_85),
.Y(n_87)
);

A2O1A1O1Ixp25_ASAP7_75t_L g88 ( 
.A1(n_86),
.A2(n_82),
.B(n_75),
.C(n_77),
.D(n_80),
.Y(n_88)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_88),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_89),
.B(n_78),
.Y(n_90)
);

XNOR2xp5_ASAP7_75t_L g91 ( 
.A(n_90),
.B(n_84),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_91),
.B(n_87),
.C(n_67),
.Y(n_92)
);

AOI21xp5_ASAP7_75t_SL g93 ( 
.A1(n_92),
.A2(n_73),
.B(n_27),
.Y(n_93)
);

XOR2xp5_ASAP7_75t_L g94 ( 
.A(n_93),
.B(n_73),
.Y(n_94)
);


endmodule